module tt_um_keszocze_ssmcl (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire a1_1;
 wire bIn;
 wire \c$case_alt_13 ;
 wire \c$case_scrut ;
 wire \c$ds_app_arg_1[0] ;
 wire \c$ds_app_arg_1[10] ;
 wire \c$ds_app_arg_1[11] ;
 wire \c$ds_app_arg_1[12] ;
 wire \c$ds_app_arg_1[13] ;
 wire \c$ds_app_arg_1[14] ;
 wire \c$ds_app_arg_1[16] ;
 wire \c$ds_app_arg_1[17] ;
 wire \c$ds_app_arg_1[18] ;
 wire \c$ds_app_arg_1[19] ;
 wire \c$ds_app_arg_1[20] ;
 wire \c$ds_app_arg_1[21] ;
 wire \c$ds_app_arg_1[22] ;
 wire \c$ds_app_arg_1[23] ;
 wire \c$ds_app_arg_1[2] ;
 wire \c$ds_app_arg_1[3] ;
 wire \c$ds_app_arg_1[5] ;
 wire \c$ds_app_arg_1[6] ;
 wire \c$ds_app_arg_1[7] ;
 wire \c$ds_app_arg_1[8] ;
 wire \c$ds_app_arg_1[9] ;
 wire \c$ds_app_arg_2[0] ;
 wire \c$ds_app_arg_2[10] ;
 wire \c$ds_app_arg_2[11] ;
 wire \c$ds_app_arg_2[12] ;
 wire \c$ds_app_arg_2[1] ;
 wire \c$ds_app_arg_2[2] ;
 wire \c$ds_app_arg_2[3] ;
 wire \c$ds_app_arg_2[4] ;
 wire \c$ds_app_arg_2[5] ;
 wire \c$ds_app_arg_2[6] ;
 wire \c$ds_app_arg_2[7] ;
 wire \c$ds_app_arg_2[8] ;
 wire \c$ds_app_arg_2[9] ;
 wire \result_7[0] ;
 wire \result_7[1] ;
 wire \result_7[2] ;
 wire \result_7[3] ;
 wire \result_7[4] ;
 wire \result_7[5] ;
 wire \s[0] ;
 wire \s[10] ;
 wire \s[1] ;
 wire \s[2] ;
 wire \s[3] ;
 wire \s[4] ;
 wire \s[5] ;
 wire \s[6] ;
 wire \s[7] ;
 wire \s[8] ;
 wire \s_0[0] ;
 wire \s_0[10] ;
 wire \s_0[1] ;
 wire \s_0[2] ;
 wire \s_0[3] ;
 wire \s_0[4] ;
 wire \s_0[7] ;
 wire \s_0[8] ;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire clknet_0_clk;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;

 sg13g2_inv_1 _289_ (.Y(_064_),
    .A(net81));
 sg13g2_inv_1 _290_ (.Y(_065_),
    .A(net53));
 sg13g2_inv_2 _291_ (.Y(_066_),
    .A(\s_0[10] ));
 sg13g2_inv_2 _292_ (.Y(_067_),
    .A(net69));
 sg13g2_inv_1 _293_ (.Y(_068_),
    .A(net57));
 sg13g2_inv_1 _294_ (.Y(_069_),
    .A(net143));
 sg13g2_inv_1 _295_ (.Y(_070_),
    .A(\c$case_alt_13 ));
 sg13g2_inv_1 _296_ (.Y(_071_),
    .A(net121));
 sg13g2_inv_1 _297_ (.Y(_072_),
    .A(net59));
 sg13g2_inv_1 _298_ (.Y(_073_),
    .A(\c$ds_app_arg_1[19] ));
 sg13g2_inv_1 _299_ (.Y(_074_),
    .A(net117));
 sg13g2_inv_1 _300_ (.Y(_075_),
    .A(net52));
 sg13g2_inv_1 _301_ (.Y(_076_),
    .A(net112));
 sg13g2_inv_1 _302_ (.Y(_077_),
    .A(net84));
 sg13g2_inv_1 _303_ (.Y(_078_),
    .A(net115));
 sg13g2_inv_1 _304_ (.Y(_079_),
    .A(net102));
 sg13g2_inv_1 _305_ (.Y(_080_),
    .A(net125));
 sg13g2_inv_1 _306_ (.Y(_081_),
    .A(net76));
 sg13g2_inv_1 _307_ (.Y(_082_),
    .A(net36));
 sg13g2_inv_1 _308_ (.Y(_083_),
    .A(net7));
 sg13g2_inv_1 _309_ (.Y(_084_),
    .A(net4));
 sg13g2_inv_1 _310_ (.Y(_085_),
    .A(\c$ds_app_arg_2[6] ));
 sg13g2_inv_1 _311_ (.Y(_086_),
    .A(net124));
 sg13g2_inv_1 _312_ (.Y(_087_),
    .A(\c$ds_app_arg_2[7] ));
 sg13g2_inv_1 _313_ (.Y(_088_),
    .A(\c$ds_app_arg_2[8] ));
 sg13g2_inv_1 _314_ (.Y(_089_),
    .A(net42));
 sg13g2_inv_1 _315_ (.Y(_090_),
    .A(\c$ds_app_arg_2[10] ));
 sg13g2_inv_1 _316_ (.Y(_091_),
    .A(net26));
 sg13g2_and2_2 _317_ (.A(net57),
    .B(\c$ds_app_arg_1[22] ),
    .X(_092_));
 sg13g2_nand2_2 _318_ (.Y(_093_),
    .A(net56),
    .B(\c$ds_app_arg_1[22] ));
 sg13g2_nor2_2 _319_ (.A(\c$ds_app_arg_2[12] ),
    .B(_092_),
    .Y(_094_));
 sg13g2_and2_1 _320_ (.A(\c$ds_app_arg_2[12] ),
    .B(\c$ds_app_arg_2[1] ),
    .X(_095_));
 sg13g2_a22oi_1 _321_ (.Y(_096_),
    .B1(_095_),
    .B2(\c$ds_app_arg_2[6] ),
    .A2(_094_),
    .A1(\c$ds_app_arg_2[0] ));
 sg13g2_inv_1 _322_ (.Y(\result_7[0] ),
    .A(_096_));
 sg13g2_and2_2 _323_ (.A(\c$ds_app_arg_2[12] ),
    .B(\c$ds_app_arg_2[6] ),
    .X(_097_));
 sg13g2_a22oi_1 _324_ (.Y(_098_),
    .B1(_097_),
    .B2(\c$ds_app_arg_2[2] ),
    .A2(_094_),
    .A1(\c$ds_app_arg_2[1] ));
 sg13g2_inv_1 _325_ (.Y(\result_7[1] ),
    .A(_098_));
 sg13g2_a22oi_1 _326_ (.Y(_099_),
    .B1(_097_),
    .B2(\c$ds_app_arg_2[3] ),
    .A2(_094_),
    .A1(\c$ds_app_arg_2[2] ));
 sg13g2_inv_1 _327_ (.Y(\result_7[2] ),
    .A(_099_));
 sg13g2_a22oi_1 _328_ (.Y(_100_),
    .B1(_097_),
    .B2(\c$ds_app_arg_2[4] ),
    .A2(_094_),
    .A1(\c$ds_app_arg_2[3] ));
 sg13g2_inv_1 _329_ (.Y(\result_7[3] ),
    .A(_100_));
 sg13g2_a22oi_1 _330_ (.Y(_101_),
    .B1(_097_),
    .B2(\c$ds_app_arg_2[5] ),
    .A2(_094_),
    .A1(\c$ds_app_arg_2[4] ));
 sg13g2_inv_1 _331_ (.Y(\result_7[4] ),
    .A(_101_));
 sg13g2_nand3_1 _332_ (.B(_092_),
    .C(_097_),
    .A(bIn),
    .Y(_102_));
 sg13g2_nand2_1 _333_ (.Y(_103_),
    .A(\c$ds_app_arg_2[5] ),
    .B(_094_));
 sg13g2_nand2_1 _334_ (.Y(\result_7[5] ),
    .A(_102_),
    .B(_103_));
 sg13g2_a21o_1 _335_ (.A2(_094_),
    .A1(\c$ds_app_arg_2[11] ),
    .B1(_097_),
    .X(a1_1));
 sg13g2_o21ai_1 _336_ (.B1(_072_),
    .Y(_104_),
    .A1(\s[6] ),
    .A2(\s[5] ));
 sg13g2_or2_1 _337_ (.X(_105_),
    .B(\c$ds_app_arg_1[22] ),
    .A(net56));
 sg13g2_a21oi_2 _338_ (.B1(_105_),
    .Y(_106_),
    .A2(net59),
    .A1(net8));
 sg13g2_and2_1 _339_ (.A(_104_),
    .B(_106_),
    .X(_107_));
 sg13g2_a21oi_2 _340_ (.B1(_067_),
    .Y(_108_),
    .A2(_106_),
    .A1(_104_));
 sg13g2_nand3_1 _341_ (.B(_093_),
    .C(_108_),
    .A(net36),
    .Y(_109_));
 sg13g2_nand3_1 _342_ (.B(\c$ds_app_arg_1[22] ),
    .C(net141),
    .A(net56),
    .Y(_110_));
 sg13g2_a221oi_1 _343_ (.B2(_106_),
    .C1(_067_),
    .B1(_104_),
    .A1(net144),
    .Y(_111_),
    .A2(_092_));
 sg13g2_o21ai_1 _344_ (.B1(_109_),
    .Y(_009_),
    .A1(_073_),
    .A2(_111_));
 sg13g2_nand3_1 _345_ (.B(_093_),
    .C(_108_),
    .A(net88),
    .Y(_112_));
 sg13g2_o21ai_1 _346_ (.B1(_112_),
    .Y(_010_),
    .A1(_082_),
    .A2(_111_));
 sg13g2_nor2b_2 _347_ (.A(\c$ds_app_arg_1[22] ),
    .B_N(net56),
    .Y(_113_));
 sg13g2_nand2_2 _348_ (.Y(_114_),
    .A(net56),
    .B(_069_));
 sg13g2_nand3_1 _349_ (.B(net59),
    .C(net5),
    .A(net8),
    .Y(_115_));
 sg13g2_o21ai_1 _350_ (.B1(_115_),
    .Y(_116_),
    .A1(\s[10] ),
    .A2(net96));
 sg13g2_a22oi_1 _351_ (.Y(_117_),
    .B1(net97),
    .B2(_068_),
    .A2(_113_),
    .A1(\c$ds_app_arg_1[19] ));
 sg13g2_nor2_1 _352_ (.A(net88),
    .B(_111_),
    .Y(_118_));
 sg13g2_a21oi_1 _353_ (.A1(_111_),
    .A2(net98),
    .Y(_011_),
    .B1(_118_));
 sg13g2_o21ai_1 _354_ (.B1(net70),
    .Y(_119_),
    .A1(net8),
    .A2(_072_));
 sg13g2_nor3_2 _355_ (.A(\s[1] ),
    .B(\s[0] ),
    .C(net99),
    .Y(_120_));
 sg13g2_nor2b_1 _356_ (.A(net145),
    .B_N(_120_),
    .Y(_121_));
 sg13g2_nor2_1 _357_ (.A(net59),
    .B(net47),
    .Y(_122_));
 sg13g2_a21o_2 _358_ (.A2(_122_),
    .A1(_121_),
    .B1(_119_),
    .X(_123_));
 sg13g2_o21ai_1 _359_ (.B1(_123_),
    .Y(_012_),
    .A1(_065_),
    .A2(net70));
 sg13g2_nor2_2 _360_ (.A(\c$case_alt_13 ),
    .B(_114_),
    .Y(_124_));
 sg13g2_nand2b_2 _361_ (.Y(_125_),
    .B(_108_),
    .A_N(_124_));
 sg13g2_nor2b_2 _362_ (.A(_124_),
    .B_N(_111_),
    .Y(_126_));
 sg13g2_and2_1 _363_ (.A(net95),
    .B(_093_),
    .X(_127_));
 sg13g2_mux2_1 _364_ (.A0(net138),
    .A1(_127_),
    .S(_126_),
    .X(_013_));
 sg13g2_and2_1 _365_ (.A(net86),
    .B(_093_),
    .X(_128_));
 sg13g2_mux2_1 _366_ (.A0(net95),
    .A1(_128_),
    .S(_126_),
    .X(_014_));
 sg13g2_a21oi_1 _367_ (.A1(net8),
    .A2(net2),
    .Y(_129_),
    .B1(_066_));
 sg13g2_a21oi_1 _368_ (.A1(_066_),
    .A2(_005_),
    .Y(_130_),
    .B1(net57));
 sg13g2_nor2b_1 _369_ (.A(_129_),
    .B_N(_130_),
    .Y(_131_));
 sg13g2_mux2_1 _370_ (.A0(net86),
    .A1(_131_),
    .S(_126_),
    .X(_015_));
 sg13g2_and2_1 _371_ (.A(net69),
    .B(\c$ds_app_arg_2[12] ),
    .X(_132_));
 sg13g2_o21ai_1 _372_ (.B1(net69),
    .Y(_133_),
    .A1(\c$ds_app_arg_2[12] ),
    .A2(_092_));
 sg13g2_nor2_2 _373_ (.A(_067_),
    .B(_094_),
    .Y(_134_));
 sg13g2_a22oi_1 _374_ (.Y(_135_),
    .B1(_133_),
    .B2(net45),
    .A2(_095_),
    .A1(net69));
 sg13g2_inv_1 _375_ (.Y(_016_),
    .A(net46));
 sg13g2_a22oi_1 _376_ (.Y(_136_),
    .B1(_133_),
    .B2(net82),
    .A2(_132_),
    .A1(\c$ds_app_arg_2[2] ));
 sg13g2_inv_1 _377_ (.Y(_017_),
    .A(net83));
 sg13g2_a22oi_1 _378_ (.Y(_137_),
    .B1(_133_),
    .B2(net89),
    .A2(_132_),
    .A1(\c$ds_app_arg_2[3] ));
 sg13g2_inv_1 _379_ (.Y(_018_),
    .A(net90));
 sg13g2_a22oi_1 _380_ (.Y(_138_),
    .B1(_133_),
    .B2(net101),
    .A2(_132_),
    .A1(net91));
 sg13g2_inv_1 _381_ (.Y(_019_),
    .A(_138_));
 sg13g2_a22oi_1 _382_ (.Y(_139_),
    .B1(_133_),
    .B2(net91),
    .A2(_132_),
    .A1(\c$ds_app_arg_2[5] ));
 sg13g2_inv_1 _383_ (.Y(_020_),
    .A(net92));
 sg13g2_nand3_1 _384_ (.B(net117),
    .C(_092_),
    .A(net69),
    .Y(_140_));
 sg13g2_o21ai_1 _385_ (.B1(_140_),
    .Y(_021_),
    .A1(_086_),
    .A2(_134_));
 sg13g2_nor2b_2 _386_ (.A(\c$ds_app_arg_2[6] ),
    .B_N(\c$ds_app_arg_2[12] ),
    .Y(_141_));
 sg13g2_a21oi_1 _387_ (.A1(net107),
    .A2(_141_),
    .Y(_142_),
    .B1(_133_));
 sg13g2_a21oi_1 _388_ (.A1(_085_),
    .A2(_133_),
    .Y(_022_),
    .B1(net108));
 sg13g2_nand3_1 _389_ (.B(_134_),
    .C(_141_),
    .A(net71),
    .Y(_143_));
 sg13g2_o21ai_1 _390_ (.B1(net72),
    .Y(_023_),
    .A1(_087_),
    .A2(_134_));
 sg13g2_nand3_1 _391_ (.B(_134_),
    .C(_141_),
    .A(net42),
    .Y(_144_));
 sg13g2_o21ai_1 _392_ (.B1(net43),
    .Y(_024_),
    .A1(_088_),
    .A2(_134_));
 sg13g2_nand3_1 _393_ (.B(_134_),
    .C(_141_),
    .A(net74),
    .Y(_145_));
 sg13g2_o21ai_1 _394_ (.B1(net75),
    .Y(_025_),
    .A1(_089_),
    .A2(_134_));
 sg13g2_nand3_1 _395_ (.B(net28),
    .C(_092_),
    .A(net69),
    .Y(_146_));
 sg13g2_o21ai_1 _396_ (.B1(_146_),
    .Y(_026_),
    .A1(_090_),
    .A2(_134_));
 sg13g2_a22oi_1 _397_ (.Y(_147_),
    .B1(_133_),
    .B2(net40),
    .A2(_097_),
    .A1(net69));
 sg13g2_inv_1 _398_ (.Y(_027_),
    .A(net41));
 sg13g2_o21ai_1 _399_ (.B1(_105_),
    .Y(_148_),
    .A1(net58),
    .A2(_076_));
 sg13g2_mux2_1 _400_ (.A0(_148_),
    .A1(net119),
    .S(_125_),
    .X(_028_));
 sg13g2_nand2b_1 _401_ (.Y(_149_),
    .B(\c$ds_app_arg_1[22] ),
    .A_N(net56));
 sg13g2_nor2b_2 _402_ (.A(net58),
    .B_N(\c$case_alt_13 ),
    .Y(_150_));
 sg13g2_and2_2 _403_ (.A(_113_),
    .B(_150_),
    .X(_151_));
 sg13g2_nor2_1 _404_ (.A(_069_),
    .B(\c$case_scrut ),
    .Y(_152_));
 sg13g2_nor2_1 _405_ (.A(net58),
    .B(\c$ds_app_arg_1[7] ),
    .Y(_153_));
 sg13g2_o21ai_1 _406_ (.B1(\c$ds_app_arg_1[7] ),
    .Y(_154_),
    .A1(_151_),
    .A2(_152_));
 sg13g2_o21ai_1 _407_ (.B1(_154_),
    .Y(_155_),
    .A1(_149_),
    .A2(_153_));
 sg13g2_mux2_1 _408_ (.A0(_155_),
    .A1(net112),
    .S(_125_),
    .X(_029_));
 sg13g2_nor2b_1 _409_ (.A(net58),
    .B_N(_105_),
    .Y(_156_));
 sg13g2_and2_1 _410_ (.A(net114),
    .B(_156_),
    .X(_157_));
 sg13g2_mux2_1 _411_ (.A0(_157_),
    .A1(net127),
    .S(_125_),
    .X(_030_));
 sg13g2_and2_1 _412_ (.A(net106),
    .B(_156_),
    .X(_158_));
 sg13g2_mux2_1 _413_ (.A0(_158_),
    .A1(net114),
    .S(_125_),
    .X(_031_));
 sg13g2_and2_1 _414_ (.A(\c$case_alt_13 ),
    .B(net58),
    .X(_159_));
 sg13g2_nand2_1 _415_ (.Y(_160_),
    .A(\c$case_alt_13 ),
    .B(net58));
 sg13g2_nor2_2 _416_ (.A(_114_),
    .B(_160_),
    .Y(_161_));
 sg13g2_and2_1 _417_ (.A(_108_),
    .B(_161_),
    .X(_162_));
 sg13g2_a21o_1 _418_ (.A2(_125_),
    .A1(net106),
    .B1(_162_),
    .X(_032_));
 sg13g2_a21o_1 _419_ (.A2(\c$case_scrut ),
    .A1(\c$ds_app_arg_1[22] ),
    .B1(net56),
    .X(_163_));
 sg13g2_nor2_1 _420_ (.A(net141),
    .B(_149_),
    .Y(_164_));
 sg13g2_nand3b_1 _421_ (.B(_163_),
    .C(net70),
    .Y(_165_),
    .A_N(_164_));
 sg13g2_and3_1 _422_ (.X(_166_),
    .A(\c$ds_app_arg_1[16] ),
    .B(\c$ds_app_arg_1[19] ),
    .C(bIn));
 sg13g2_nand3_1 _423_ (.B(\c$ds_app_arg_1[19] ),
    .C(bIn),
    .A(\c$ds_app_arg_1[16] ),
    .Y(_167_));
 sg13g2_a21o_1 _424_ (.A2(\c$ds_app_arg_1[19] ),
    .A1(\c$ds_app_arg_1[16] ),
    .B1(bIn),
    .X(_168_));
 sg13g2_and3_1 _425_ (.X(_169_),
    .A(\c$ds_app_arg_1[0] ),
    .B(_167_),
    .C(_168_));
 sg13g2_a21oi_2 _426_ (.B1(\c$ds_app_arg_1[0] ),
    .Y(_170_),
    .A2(_168_),
    .A1(_167_));
 sg13g2_o21ai_1 _427_ (.B1(_070_),
    .Y(_171_),
    .A1(_169_),
    .A2(_170_));
 sg13g2_a21oi_2 _428_ (.B1(_166_),
    .Y(_172_),
    .A2(_168_),
    .A1(net139));
 sg13g2_a221oi_1 _429_ (.B2(_172_),
    .C1(_114_),
    .B1(_159_),
    .A1(_001_),
    .Y(_173_),
    .A2(_150_));
 sg13g2_nor2_2 _430_ (.A(net58),
    .B(_093_),
    .Y(_174_));
 sg13g2_a221oi_1 _431_ (.B2(bIn),
    .C1(net55),
    .B1(_174_),
    .A1(_171_),
    .Y(_175_),
    .A2(_173_));
 sg13g2_a21oi_1 _432_ (.A1(_078_),
    .A2(net55),
    .Y(_033_),
    .B1(_175_));
 sg13g2_o21ai_1 _433_ (.B1(_159_),
    .Y(_176_),
    .A1(_169_),
    .A2(_170_));
 sg13g2_a221oi_1 _434_ (.B2(_003_),
    .C1(_114_),
    .B1(_150_),
    .A1(_070_),
    .Y(_177_),
    .A2(_002_));
 sg13g2_a221oi_1 _435_ (.B2(_177_),
    .C1(net54),
    .B1(_176_),
    .A1(\c$ds_app_arg_1[10] ),
    .Y(_178_),
    .A2(_174_));
 sg13g2_a21oi_1 _436_ (.A1(_077_),
    .A2(net54),
    .Y(_034_),
    .B1(_178_));
 sg13g2_o21ai_1 _437_ (.B1(net84),
    .Y(_179_),
    .A1(_124_),
    .A2(_174_));
 sg13g2_a221oi_1 _438_ (.B2(\c$ds_app_arg_1[10] ),
    .C1(net54),
    .B1(_161_),
    .A1(\c$ds_app_arg_1[13] ),
    .Y(_180_),
    .A2(_151_));
 sg13g2_a22oi_1 _439_ (.Y(_035_),
    .B1(_179_),
    .B2(_180_),
    .A2(net54),
    .A1(_079_));
 sg13g2_a21oi_1 _440_ (.A1(_070_),
    .A2(_003_),
    .Y(_181_),
    .B1(_114_));
 sg13g2_a22oi_1 _441_ (.Y(_182_),
    .B1(_172_),
    .B2(_150_),
    .A2(_159_),
    .A1(_001_));
 sg13g2_a221oi_1 _442_ (.B2(_182_),
    .C1(net54),
    .B1(_181_),
    .A1(net102),
    .Y(_183_),
    .A2(_174_));
 sg13g2_a21oi_1 _443_ (.A1(_080_),
    .A2(net54),
    .Y(_036_),
    .B1(_183_));
 sg13g2_o21ai_1 _444_ (.B1(_150_),
    .Y(_184_),
    .A1(_169_),
    .A2(_170_));
 sg13g2_a221oi_1 _445_ (.B2(_003_),
    .C1(_114_),
    .B1(_159_),
    .A1(_070_),
    .Y(_185_),
    .A2(_004_));
 sg13g2_a221oi_1 _446_ (.B2(_185_),
    .C1(net55),
    .B1(_184_),
    .A1(\c$ds_app_arg_1[13] ),
    .Y(_186_),
    .A2(_174_));
 sg13g2_a21oi_1 _447_ (.A1(_081_),
    .A2(net54),
    .Y(_037_),
    .B1(_186_));
 sg13g2_o21ai_1 _448_ (.B1(net76),
    .Y(_187_),
    .A1(_124_),
    .A2(_174_));
 sg13g2_a221oi_1 _449_ (.B2(\c$ds_app_arg_1[13] ),
    .C1(net54),
    .B1(_161_),
    .A1(net115),
    .Y(_188_),
    .A2(_151_));
 sg13g2_a22oi_1 _450_ (.Y(_038_),
    .B1(_187_),
    .B2(_188_),
    .A2(net55),
    .A1(_074_));
 sg13g2_nand2_1 _451_ (.Y(_189_),
    .A(_110_),
    .B(_163_));
 sg13g2_nand3_1 _452_ (.B(_110_),
    .C(_163_),
    .A(net70),
    .Y(_190_));
 sg13g2_or2_1 _453_ (.X(_191_),
    .B(_190_),
    .A(_164_));
 sg13g2_nor4_1 _454_ (.A(net120),
    .B(_114_),
    .C(_172_),
    .D(_191_),
    .Y(_192_));
 sg13g2_a21o_1 _455_ (.A2(_191_),
    .A1(net139),
    .B1(_192_),
    .X(_039_));
 sg13g2_nand3_1 _456_ (.B(_113_),
    .C(_160_),
    .A(net50),
    .Y(_193_));
 sg13g2_nand2_1 _457_ (.Y(_194_),
    .A(net120),
    .B(_190_));
 sg13g2_o21ai_1 _458_ (.B1(_194_),
    .Y(_040_),
    .A1(_190_),
    .A2(_193_));
 sg13g2_nand3_1 _459_ (.B(_113_),
    .C(_160_),
    .A(\c$ds_app_arg_1[3] ),
    .Y(_195_));
 sg13g2_nand2_1 _460_ (.Y(_196_),
    .A(net50),
    .B(_190_));
 sg13g2_o21ai_1 _461_ (.B1(_196_),
    .Y(_041_),
    .A1(_190_),
    .A2(_195_));
 sg13g2_nor2_1 _462_ (.A(_151_),
    .B(_191_),
    .Y(_197_));
 sg13g2_a21oi_1 _463_ (.A1(_075_),
    .A2(_190_),
    .Y(_042_),
    .B1(_197_));
 sg13g2_o21ai_1 _464_ (.B1(net1),
    .Y(_198_),
    .A1(_066_),
    .A2(net8));
 sg13g2_nor3_2 _465_ (.A(\s_0[1] ),
    .B(\s_0[0] ),
    .C(net93),
    .Y(_199_));
 sg13g2_nor2b_1 _466_ (.A(\s_0[3] ),
    .B_N(_199_),
    .Y(_200_));
 sg13g2_nor2_1 _467_ (.A(\s_0[10] ),
    .B(net78),
    .Y(_201_));
 sg13g2_a21o_2 _468_ (.A2(_201_),
    .A1(_200_),
    .B1(_198_),
    .X(_202_));
 sg13g2_nand2b_2 _469_ (.Y(_203_),
    .B(_066_),
    .A_N(_202_));
 sg13g2_nand2_1 _470_ (.Y(_204_),
    .A(net136),
    .B(_202_));
 sg13g2_o21ai_1 _471_ (.B1(_204_),
    .Y(_043_),
    .A1(net136),
    .A2(_203_));
 sg13g2_nand2_1 _472_ (.Y(_205_),
    .A(net128),
    .B(_202_));
 sg13g2_xor2_1 _473_ (.B(\s_0[0] ),
    .A(net128),
    .X(_206_));
 sg13g2_o21ai_1 _474_ (.B1(_205_),
    .Y(_044_),
    .A1(_203_),
    .A2(_206_));
 sg13g2_nand2_1 _475_ (.Y(_207_),
    .A(net93),
    .B(_202_));
 sg13g2_o21ai_1 _476_ (.B1(net93),
    .Y(_208_),
    .A1(\s_0[1] ),
    .A2(\s_0[0] ));
 sg13g2_nor2b_1 _477_ (.A(_199_),
    .B_N(_208_),
    .Y(_209_));
 sg13g2_o21ai_1 _478_ (.B1(_207_),
    .Y(_045_),
    .A1(_203_),
    .A2(_209_));
 sg13g2_nand2_1 _479_ (.Y(_210_),
    .A(net110),
    .B(_198_));
 sg13g2_xnor2_1 _480_ (.Y(_211_),
    .A(net110),
    .B(_199_));
 sg13g2_o21ai_1 _481_ (.B1(_210_),
    .Y(_046_),
    .A1(_203_),
    .A2(_211_));
 sg13g2_nand3_1 _482_ (.B(net8),
    .C(net70),
    .A(\s_0[10] ),
    .Y(_212_));
 sg13g2_nand2b_1 _483_ (.Y(_213_),
    .B(_200_),
    .A_N(_198_));
 sg13g2_nand2_1 _484_ (.Y(_214_),
    .A(net78),
    .B(_213_));
 sg13g2_nand2_1 _485_ (.Y(_047_),
    .A(_212_),
    .B(net79));
 sg13g2_or2_1 _486_ (.X(_215_),
    .B(\s_0[8] ),
    .A(\s_0[10] ));
 sg13g2_o21ai_1 _487_ (.B1(_215_),
    .Y(_216_),
    .A1(_066_),
    .A2(net3));
 sg13g2_nand2_1 _488_ (.Y(_217_),
    .A(net30),
    .B(_198_));
 sg13g2_o21ai_1 _489_ (.B1(_217_),
    .Y(_048_),
    .A1(_198_),
    .A2(_216_));
 sg13g2_nand2_1 _490_ (.Y(_218_),
    .A(net34),
    .B(_198_));
 sg13g2_o21ai_1 _491_ (.B1(_218_),
    .Y(_049_),
    .A1(_084_),
    .A2(_212_));
 sg13g2_nor4_1 _492_ (.A(_067_),
    .B(_071_),
    .C(net130),
    .D(net59),
    .Y(_219_));
 sg13g2_a21o_1 _493_ (.A2(_119_),
    .A1(net130),
    .B1(_219_),
    .X(_050_));
 sg13g2_nand3_1 _494_ (.B(net70),
    .C(net59),
    .A(net8),
    .Y(_220_));
 sg13g2_o21ai_1 _495_ (.B1(net121),
    .Y(_221_),
    .A1(\s[5] ),
    .A2(_119_));
 sg13g2_nand2_1 _496_ (.Y(_051_),
    .A(_220_),
    .B(net122));
 sg13g2_nor2b_1 _497_ (.A(net59),
    .B_N(\s[8] ),
    .Y(_222_));
 sg13g2_a21oi_1 _498_ (.A1(net59),
    .A2(net6),
    .Y(_223_),
    .B1(_222_));
 sg13g2_nand2_1 _499_ (.Y(_224_),
    .A(net32),
    .B(_119_));
 sg13g2_o21ai_1 _500_ (.B1(_224_),
    .Y(_052_),
    .A1(_119_),
    .A2(_223_));
 sg13g2_nand2_1 _501_ (.Y(_225_),
    .A(net38),
    .B(_119_));
 sg13g2_o21ai_1 _502_ (.B1(_225_),
    .Y(_053_),
    .A1(_083_),
    .A2(_220_));
 sg13g2_a21oi_1 _503_ (.A1(net69),
    .A2(_092_),
    .Y(_226_),
    .B1(\c$ds_app_arg_2[12] ));
 sg13g2_a21oi_1 _504_ (.A1(_091_),
    .A2(_132_),
    .Y(_054_),
    .B1(_226_));
 sg13g2_o21ai_1 _505_ (.B1(net119),
    .Y(_227_),
    .A1(_151_),
    .A2(_152_));
 sg13g2_nor3_1 _506_ (.A(_067_),
    .B(_107_),
    .C(_227_),
    .Y(_228_));
 sg13g2_a21o_1 _507_ (.A2(_125_),
    .A1(net58),
    .B1(_228_),
    .X(_055_));
 sg13g2_o21ai_1 _508_ (.B1(_108_),
    .Y(_229_),
    .A1(_161_),
    .A2(_189_));
 sg13g2_o21ai_1 _509_ (.B1(_229_),
    .Y(_056_),
    .A1(net1),
    .A2(_069_));
 sg13g2_nor2_1 _510_ (.A(net56),
    .B(_108_),
    .Y(_230_));
 sg13g2_nor2_1 _511_ (.A(_113_),
    .B(_164_),
    .Y(_231_));
 sg13g2_a21oi_1 _512_ (.A1(_111_),
    .A2(_231_),
    .Y(_057_),
    .B1(_230_));
 sg13g2_nand2b_2 _513_ (.Y(_232_),
    .B(_072_),
    .A_N(_123_));
 sg13g2_nand2_1 _514_ (.Y(_233_),
    .A(net134),
    .B(_123_));
 sg13g2_o21ai_1 _515_ (.B1(_233_),
    .Y(_058_),
    .A1(net134),
    .A2(_232_));
 sg13g2_nand2_1 _516_ (.Y(_234_),
    .A(net132),
    .B(_123_));
 sg13g2_xor2_1 _517_ (.B(\s[0] ),
    .A(net132),
    .X(_235_));
 sg13g2_o21ai_1 _518_ (.B1(_234_),
    .Y(_059_),
    .A1(_232_),
    .A2(_235_));
 sg13g2_nand2_1 _519_ (.Y(_236_),
    .A(net99),
    .B(_123_));
 sg13g2_o21ai_1 _520_ (.B1(net99),
    .Y(_237_),
    .A1(\s[1] ),
    .A2(\s[0] ));
 sg13g2_nor2b_1 _521_ (.A(_120_),
    .B_N(_237_),
    .Y(_238_));
 sg13g2_o21ai_1 _522_ (.B1(_236_),
    .Y(_060_),
    .A1(_232_),
    .A2(_238_));
 sg13g2_nand2_1 _523_ (.Y(_239_),
    .A(net104),
    .B(_119_));
 sg13g2_xnor2_1 _524_ (.Y(_240_),
    .A(net104),
    .B(_120_));
 sg13g2_o21ai_1 _525_ (.B1(_239_),
    .Y(_061_),
    .A1(_232_),
    .A2(_240_));
 sg13g2_nand2b_1 _526_ (.Y(_241_),
    .B(_121_),
    .A_N(_119_));
 sg13g2_nand2_1 _527_ (.Y(_242_),
    .A(net47),
    .B(_241_));
 sg13g2_nand2_1 _528_ (.Y(_062_),
    .A(_220_),
    .B(net48));
 sg13g2_o21ai_1 _529_ (.B1(_202_),
    .Y(_063_),
    .A1(_064_),
    .A2(net70));
 sg13g2_dfrbp_1 _530_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net63),
    .D(net37),
    .Q_N(_286_),
    .Q(\c$ds_app_arg_1[19] ));
 sg13g2_dfrbp_1 _531_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net62),
    .D(_010_),
    .Q_N(_285_),
    .Q(\c$ds_app_arg_1[20] ));
 sg13g2_dfrbp_1 _532_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net62),
    .D(_011_),
    .Q_N(_284_),
    .Q(\c$ds_app_arg_1[21] ));
 sg13g2_dfrbp_1 _533_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net67),
    .D(_012_),
    .Q_N(\s[10] ),
    .Q(_287_));
 sg13g2_dfrbp_1 _534_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net65),
    .D(_013_),
    .Q_N(_283_),
    .Q(\c$ds_app_arg_1[16] ));
 sg13g2_dfrbp_1 _535_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net65),
    .D(_014_),
    .Q_N(_282_),
    .Q(\c$ds_app_arg_1[17] ));
 sg13g2_dfrbp_1 _536_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net66),
    .D(net87),
    .Q_N(_281_),
    .Q(\c$ds_app_arg_1[18] ));
 sg13g2_dfrbp_1 _537_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net61),
    .D(_016_),
    .Q_N(_280_),
    .Q(\c$ds_app_arg_2[0] ));
 sg13g2_dfrbp_1 _538_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net61),
    .D(_017_),
    .Q_N(_279_),
    .Q(\c$ds_app_arg_2[1] ));
 sg13g2_dfrbp_1 _539_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net61),
    .D(_018_),
    .Q_N(_278_),
    .Q(\c$ds_app_arg_2[2] ));
 sg13g2_dfrbp_1 _540_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net62),
    .D(_019_),
    .Q_N(_277_),
    .Q(\c$ds_app_arg_2[3] ));
 sg13g2_dfrbp_1 _541_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net61),
    .D(_020_),
    .Q_N(_276_),
    .Q(\c$ds_app_arg_2[4] ));
 sg13g2_dfrbp_1 _542_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net62),
    .D(_021_),
    .Q_N(_275_),
    .Q(\c$ds_app_arg_2[5] ));
 sg13g2_dfrbp_1 _543_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net61),
    .D(net109),
    .Q_N(_008_),
    .Q(\c$ds_app_arg_2[6] ));
 sg13g2_dfrbp_1 _544_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net61),
    .D(net73),
    .Q_N(_274_),
    .Q(\c$ds_app_arg_2[7] ));
 sg13g2_dfrbp_1 _545_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net60),
    .D(net44),
    .Q_N(_273_),
    .Q(\c$ds_app_arg_2[8] ));
 sg13g2_dfrbp_1 _546_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net60),
    .D(_025_),
    .Q_N(_272_),
    .Q(\c$ds_app_arg_2[9] ));
 sg13g2_dfrbp_1 _547_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net60),
    .D(net29),
    .Q_N(_271_),
    .Q(\c$ds_app_arg_2[10] ));
 sg13g2_dfrbp_1 _548_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net61),
    .D(_027_),
    .Q_N(_270_),
    .Q(\c$ds_app_arg_2[11] ));
 sg13g2_dfrbp_1 _549_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net65),
    .D(_028_),
    .Q_N(_269_),
    .Q(\c$ds_app_arg_1[5] ));
 sg13g2_dfrbp_1 _550_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net64),
    .D(net113),
    .Q_N(_268_),
    .Q(\c$ds_app_arg_1[6] ));
 sg13g2_dfrbp_1 _551_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net65),
    .D(_030_),
    .Q_N(_267_),
    .Q(\c$ds_app_arg_1[7] ));
 sg13g2_dfrbp_1 _552_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net64),
    .D(_031_),
    .Q_N(_266_),
    .Q(\c$ds_app_arg_1[8] ));
 sg13g2_dfrbp_1 _553_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net64),
    .D(_032_),
    .Q_N(_265_),
    .Q(\c$ds_app_arg_1[9] ));
 sg13g2_dfrbp_1 _554_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net63),
    .D(net116),
    .Q_N(_002_),
    .Q(\c$ds_app_arg_1[10] ));
 sg13g2_dfrbp_1 _555_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net63),
    .D(net85),
    .Q_N(_001_),
    .Q(\c$ds_app_arg_1[11] ));
 sg13g2_dfrbp_1 _556_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net60),
    .D(net103),
    .Q_N(_003_),
    .Q(\c$ds_app_arg_1[12] ));
 sg13g2_dfrbp_1 _557_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net60),
    .D(net126),
    .Q_N(_004_),
    .Q(\c$ds_app_arg_1[13] ));
 sg13g2_dfrbp_1 _558_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net60),
    .D(net77),
    .Q_N(_264_),
    .Q(\c$ds_app_arg_1[14] ));
 sg13g2_dfrbp_1 _559_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net60),
    .D(net118),
    .Q_N(_263_),
    .Q(bIn));
 sg13g2_dfrbp_1 _560_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net60),
    .D(_039_),
    .Q_N(_262_),
    .Q(\c$ds_app_arg_1[0] ));
 sg13g2_dfrbp_1 _561_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net64),
    .D(_040_),
    .Q_N(_261_),
    .Q(\c$case_alt_13 ));
 sg13g2_dfrbp_1 _562_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net64),
    .D(net51),
    .Q_N(_260_),
    .Q(\c$ds_app_arg_1[2] ));
 sg13g2_dfrbp_1 _563_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net64),
    .D(_042_),
    .Q_N(_259_),
    .Q(\c$ds_app_arg_1[3] ));
 sg13g2_dfrbp_1 _564_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net66),
    .D(net137),
    .Q_N(_258_),
    .Q(\s_0[0] ));
 sg13g2_dfrbp_1 _565_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net66),
    .D(net129),
    .Q_N(_257_),
    .Q(\s_0[1] ));
 sg13g2_dfrbp_1 _566_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net66),
    .D(net94),
    .Q_N(_256_),
    .Q(\s_0[2] ));
 sg13g2_dfrbp_1 _567_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net66),
    .D(net111),
    .Q_N(_255_),
    .Q(\s_0[3] ));
 sg13g2_dfrbp_1 _568_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net66),
    .D(net80),
    .Q_N(_254_),
    .Q(\s_0[4] ));
 sg13g2_dfrbp_1 _569_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net66),
    .D(net31),
    .Q_N(_005_),
    .Q(\s_0[7] ));
 sg13g2_dfrbp_1 _570_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net66),
    .D(net35),
    .Q_N(_253_),
    .Q(\s_0[8] ));
 sg13g2_dfrbp_1 _571_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net67),
    .D(net131),
    .Q_N(_252_),
    .Q(\s[5] ));
 sg13g2_dfrbp_1 _572_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net67),
    .D(net123),
    .Q_N(_251_),
    .Q(\s[6] ));
 sg13g2_dfrbp_1 _573_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net67),
    .D(net33),
    .Q_N(_006_),
    .Q(\s[7] ));
 sg13g2_dfrbp_1 _574_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net67),
    .D(net39),
    .Q_N(_250_),
    .Q(\s[8] ));
 sg13g2_dfrbp_1 _575_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net61),
    .D(net27),
    .Q_N(_007_),
    .Q(\c$ds_app_arg_2[12] ));
 sg13g2_dfrbp_1 _576_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net64),
    .D(_055_),
    .Q_N(_000_),
    .Q(\c$case_scrut ));
 sg13g2_dfrbp_1 _577_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net64),
    .D(_056_),
    .Q_N(_249_),
    .Q(\c$ds_app_arg_1[22] ));
 sg13g2_dfrbp_1 _578_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net67),
    .D(net142),
    .Q_N(_248_),
    .Q(\c$ds_app_arg_1[23] ));
 sg13g2_dfrbp_1 _579_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net62),
    .D(net135),
    .Q_N(_247_),
    .Q(\s[0] ));
 sg13g2_dfrbp_1 _580_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net62),
    .D(net133),
    .Q_N(_246_),
    .Q(\s[1] ));
 sg13g2_dfrbp_1 _581_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net62),
    .D(net100),
    .Q_N(_245_),
    .Q(\s[2] ));
 sg13g2_dfrbp_1 _582_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net67),
    .D(net105),
    .Q_N(_244_),
    .Q(\s[3] ));
 sg13g2_dfrbp_1 _583_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net67),
    .D(net49),
    .Q_N(_243_),
    .Q(\s[4] ));
 sg13g2_dfrbp_1 _584_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net68),
    .D(_063_),
    .Q_N(\s_0[10] ),
    .Q(_288_));
 sg13g2_tielo tt_um_keszocze_ssmcl_10 (.L_LO(net10));
 sg13g2_tielo tt_um_keszocze_ssmcl_11 (.L_LO(net11));
 sg13g2_tielo tt_um_keszocze_ssmcl_12 (.L_LO(net12));
 sg13g2_tielo tt_um_keszocze_ssmcl_13 (.L_LO(net13));
 sg13g2_tielo tt_um_keszocze_ssmcl_14 (.L_LO(net14));
 sg13g2_tielo tt_um_keszocze_ssmcl_15 (.L_LO(net15));
 sg13g2_tielo tt_um_keszocze_ssmcl_16 (.L_LO(net16));
 sg13g2_tielo tt_um_keszocze_ssmcl_17 (.L_LO(net17));
 sg13g2_tielo tt_um_keszocze_ssmcl_18 (.L_LO(net18));
 sg13g2_tielo tt_um_keszocze_ssmcl_19 (.L_LO(net19));
 sg13g2_tielo tt_um_keszocze_ssmcl_20 (.L_LO(net20));
 sg13g2_tielo tt_um_keszocze_ssmcl_21 (.L_LO(net21));
 sg13g2_tielo tt_um_keszocze_ssmcl_22 (.L_LO(net22));
 sg13g2_tielo tt_um_keszocze_ssmcl_23 (.L_LO(net23));
 sg13g2_tielo tt_um_keszocze_ssmcl_24 (.L_LO(net24));
 sg13g2_tielo tt_um_keszocze_ssmcl_25 (.L_LO(net25));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_1 _602_ (.A(\result_7[0] ),
    .X(uo_out[0]));
 sg13g2_buf_1 _603_ (.A(\result_7[1] ),
    .X(uo_out[1]));
 sg13g2_buf_1 _604_ (.A(\result_7[2] ),
    .X(uo_out[2]));
 sg13g2_buf_1 _605_ (.A(\result_7[3] ),
    .X(uo_out[3]));
 sg13g2_buf_1 _606_ (.A(\result_7[4] ),
    .X(uo_out[4]));
 sg13g2_buf_1 _607_ (.A(\result_7[5] ),
    .X(uo_out[5]));
 sg13g2_buf_1 _608_ (.A(a1_1),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout54 (.A(_165_),
    .X(net54));
 sg13g2_buf_1 fanout55 (.A(_165_),
    .X(net55));
 sg13g2_buf_2 fanout56 (.A(net57),
    .X(net56));
 sg13g2_buf_1 fanout57 (.A(\c$ds_app_arg_1[23] ),
    .X(net57));
 sg13g2_buf_2 fanout58 (.A(net140),
    .X(net58));
 sg13g2_buf_2 fanout59 (.A(\s[10] ),
    .X(net59));
 sg13g2_buf_4 fanout60 (.X(net60),
    .A(net63));
 sg13g2_buf_4 fanout61 (.X(net61),
    .A(net62));
 sg13g2_buf_4 fanout62 (.X(net62),
    .A(net63));
 sg13g2_buf_2 fanout63 (.A(rst_n),
    .X(net63));
 sg13g2_buf_4 fanout64 (.X(net64),
    .A(net68));
 sg13g2_buf_2 fanout65 (.A(net68),
    .X(net65));
 sg13g2_buf_4 fanout66 (.X(net66),
    .A(net68));
 sg13g2_buf_4 fanout67 (.X(net67),
    .A(net68));
 sg13g2_buf_2 fanout68 (.A(rst_n),
    .X(net68));
 sg13g2_buf_2 fanout69 (.A(net70),
    .X(net69));
 sg13g2_buf_2 fanout70 (.A(net1),
    .X(net70));
 sg13g2_buf_1 input1 (.A(ena),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[0]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[1]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[2]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[3]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[4]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[5]),
    .X(net7));
 sg13g2_buf_2 input8 (.A(ui_in[7]),
    .X(net8));
 sg13g2_tielo tt_um_keszocze_ssmcl_9 (.L_LO(net9));
 sg13g2_buf_2 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sg13g2_buf_2 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sg13g2_buf_2 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sg13g2_buf_2 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sg13g2_buf_2 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sg13g2_buf_2 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sg13g2_buf_2 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sg13g2_buf_2 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_3_7__leaf_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(_008_),
    .X(net26));
 sg13g2_dlygate4sd3_1 hold2 (.A(_054_),
    .X(net27));
 sg13g2_dlygate4sd3_1 hold3 (.A(_007_),
    .X(net28));
 sg13g2_dlygate4sd3_1 hold4 (.A(_026_),
    .X(net29));
 sg13g2_dlygate4sd3_1 hold5 (.A(\s_0[7] ),
    .X(net30));
 sg13g2_dlygate4sd3_1 hold6 (.A(_048_),
    .X(net31));
 sg13g2_dlygate4sd3_1 hold7 (.A(\s[7] ),
    .X(net32));
 sg13g2_dlygate4sd3_1 hold8 (.A(_052_),
    .X(net33));
 sg13g2_dlygate4sd3_1 hold9 (.A(\s_0[8] ),
    .X(net34));
 sg13g2_dlygate4sd3_1 hold10 (.A(_049_),
    .X(net35));
 sg13g2_dlygate4sd3_1 hold11 (.A(\c$ds_app_arg_1[20] ),
    .X(net36));
 sg13g2_dlygate4sd3_1 hold12 (.A(_009_),
    .X(net37));
 sg13g2_dlygate4sd3_1 hold13 (.A(\s[8] ),
    .X(net38));
 sg13g2_dlygate4sd3_1 hold14 (.A(_053_),
    .X(net39));
 sg13g2_dlygate4sd3_1 hold15 (.A(\c$ds_app_arg_2[11] ),
    .X(net40));
 sg13g2_dlygate4sd3_1 hold16 (.A(_147_),
    .X(net41));
 sg13g2_dlygate4sd3_1 hold17 (.A(\c$ds_app_arg_2[9] ),
    .X(net42));
 sg13g2_dlygate4sd3_1 hold18 (.A(_144_),
    .X(net43));
 sg13g2_dlygate4sd3_1 hold19 (.A(_024_),
    .X(net44));
 sg13g2_dlygate4sd3_1 hold20 (.A(\c$ds_app_arg_2[0] ),
    .X(net45));
 sg13g2_dlygate4sd3_1 hold21 (.A(_135_),
    .X(net46));
 sg13g2_dlygate4sd3_1 hold22 (.A(\s[4] ),
    .X(net47));
 sg13g2_dlygate4sd3_1 hold23 (.A(_242_),
    .X(net48));
 sg13g2_dlygate4sd3_1 hold24 (.A(_062_),
    .X(net49));
 sg13g2_dlygate4sd3_1 hold25 (.A(\c$ds_app_arg_1[2] ),
    .X(net50));
 sg13g2_dlygate4sd3_1 hold26 (.A(_041_),
    .X(net51));
 sg13g2_dlygate4sd3_1 hold27 (.A(\c$ds_app_arg_1[3] ),
    .X(net52));
 sg13g2_dlygate4sd3_1 hold28 (.A(_287_),
    .X(net53));
 sg13g2_dlygate4sd3_1 hold29 (.A(\c$ds_app_arg_2[8] ),
    .X(net71));
 sg13g2_dlygate4sd3_1 hold30 (.A(_143_),
    .X(net72));
 sg13g2_dlygate4sd3_1 hold31 (.A(_023_),
    .X(net73));
 sg13g2_dlygate4sd3_1 hold32 (.A(\c$ds_app_arg_2[10] ),
    .X(net74));
 sg13g2_dlygate4sd3_1 hold33 (.A(_145_),
    .X(net75));
 sg13g2_dlygate4sd3_1 hold34 (.A(\c$ds_app_arg_1[14] ),
    .X(net76));
 sg13g2_dlygate4sd3_1 hold35 (.A(_037_),
    .X(net77));
 sg13g2_dlygate4sd3_1 hold36 (.A(\s_0[4] ),
    .X(net78));
 sg13g2_dlygate4sd3_1 hold37 (.A(_214_),
    .X(net79));
 sg13g2_dlygate4sd3_1 hold38 (.A(_047_),
    .X(net80));
 sg13g2_dlygate4sd3_1 hold39 (.A(_288_),
    .X(net81));
 sg13g2_dlygate4sd3_1 hold40 (.A(\c$ds_app_arg_2[1] ),
    .X(net82));
 sg13g2_dlygate4sd3_1 hold41 (.A(_136_),
    .X(net83));
 sg13g2_dlygate4sd3_1 hold42 (.A(\c$ds_app_arg_1[11] ),
    .X(net84));
 sg13g2_dlygate4sd3_1 hold43 (.A(_034_),
    .X(net85));
 sg13g2_dlygate4sd3_1 hold44 (.A(\c$ds_app_arg_1[18] ),
    .X(net86));
 sg13g2_dlygate4sd3_1 hold45 (.A(_015_),
    .X(net87));
 sg13g2_dlygate4sd3_1 hold46 (.A(\c$ds_app_arg_1[21] ),
    .X(net88));
 sg13g2_dlygate4sd3_1 hold47 (.A(\c$ds_app_arg_2[2] ),
    .X(net89));
 sg13g2_dlygate4sd3_1 hold48 (.A(_137_),
    .X(net90));
 sg13g2_dlygate4sd3_1 hold49 (.A(\c$ds_app_arg_2[4] ),
    .X(net91));
 sg13g2_dlygate4sd3_1 hold50 (.A(_139_),
    .X(net92));
 sg13g2_dlygate4sd3_1 hold51 (.A(\s_0[2] ),
    .X(net93));
 sg13g2_dlygate4sd3_1 hold52 (.A(_045_),
    .X(net94));
 sg13g2_dlygate4sd3_1 hold53 (.A(\c$ds_app_arg_1[17] ),
    .X(net95));
 sg13g2_dlygate4sd3_1 hold54 (.A(_006_),
    .X(net96));
 sg13g2_dlygate4sd3_1 hold55 (.A(_116_),
    .X(net97));
 sg13g2_dlygate4sd3_1 hold56 (.A(_117_),
    .X(net98));
 sg13g2_dlygate4sd3_1 hold57 (.A(\s[2] ),
    .X(net99));
 sg13g2_dlygate4sd3_1 hold58 (.A(_060_),
    .X(net100));
 sg13g2_dlygate4sd3_1 hold59 (.A(\c$ds_app_arg_2[3] ),
    .X(net101));
 sg13g2_dlygate4sd3_1 hold60 (.A(\c$ds_app_arg_1[12] ),
    .X(net102));
 sg13g2_dlygate4sd3_1 hold61 (.A(_035_),
    .X(net103));
 sg13g2_dlygate4sd3_1 hold62 (.A(\s[3] ),
    .X(net104));
 sg13g2_dlygate4sd3_1 hold63 (.A(_061_),
    .X(net105));
 sg13g2_dlygate4sd3_1 hold64 (.A(\c$ds_app_arg_1[9] ),
    .X(net106));
 sg13g2_dlygate4sd3_1 hold65 (.A(\c$ds_app_arg_2[7] ),
    .X(net107));
 sg13g2_dlygate4sd3_1 hold66 (.A(_142_),
    .X(net108));
 sg13g2_dlygate4sd3_1 hold67 (.A(_022_),
    .X(net109));
 sg13g2_dlygate4sd3_1 hold68 (.A(\s_0[3] ),
    .X(net110));
 sg13g2_dlygate4sd3_1 hold69 (.A(_046_),
    .X(net111));
 sg13g2_dlygate4sd3_1 hold70 (.A(\c$ds_app_arg_1[6] ),
    .X(net112));
 sg13g2_dlygate4sd3_1 hold71 (.A(_029_),
    .X(net113));
 sg13g2_dlygate4sd3_1 hold72 (.A(\c$ds_app_arg_1[8] ),
    .X(net114));
 sg13g2_dlygate4sd3_1 hold73 (.A(\c$ds_app_arg_1[10] ),
    .X(net115));
 sg13g2_dlygate4sd3_1 hold74 (.A(_033_),
    .X(net116));
 sg13g2_dlygate4sd3_1 hold75 (.A(bIn),
    .X(net117));
 sg13g2_dlygate4sd3_1 hold76 (.A(_038_),
    .X(net118));
 sg13g2_dlygate4sd3_1 hold77 (.A(\c$ds_app_arg_1[5] ),
    .X(net119));
 sg13g2_dlygate4sd3_1 hold78 (.A(\c$case_alt_13 ),
    .X(net120));
 sg13g2_dlygate4sd3_1 hold79 (.A(\s[6] ),
    .X(net121));
 sg13g2_dlygate4sd3_1 hold80 (.A(_221_),
    .X(net122));
 sg13g2_dlygate4sd3_1 hold81 (.A(_051_),
    .X(net123));
 sg13g2_dlygate4sd3_1 hold82 (.A(\c$ds_app_arg_2[5] ),
    .X(net124));
 sg13g2_dlygate4sd3_1 hold83 (.A(\c$ds_app_arg_1[13] ),
    .X(net125));
 sg13g2_dlygate4sd3_1 hold84 (.A(_036_),
    .X(net126));
 sg13g2_dlygate4sd3_1 hold85 (.A(\c$ds_app_arg_1[7] ),
    .X(net127));
 sg13g2_dlygate4sd3_1 hold86 (.A(\s_0[1] ),
    .X(net128));
 sg13g2_dlygate4sd3_1 hold87 (.A(_044_),
    .X(net129));
 sg13g2_dlygate4sd3_1 hold88 (.A(\s[5] ),
    .X(net130));
 sg13g2_dlygate4sd3_1 hold89 (.A(_050_),
    .X(net131));
 sg13g2_dlygate4sd3_1 hold90 (.A(\s[1] ),
    .X(net132));
 sg13g2_dlygate4sd3_1 hold91 (.A(_059_),
    .X(net133));
 sg13g2_dlygate4sd3_1 hold92 (.A(\s[0] ),
    .X(net134));
 sg13g2_dlygate4sd3_1 hold93 (.A(_058_),
    .X(net135));
 sg13g2_dlygate4sd3_1 hold94 (.A(\s_0[0] ),
    .X(net136));
 sg13g2_dlygate4sd3_1 hold95 (.A(_043_),
    .X(net137));
 sg13g2_dlygate4sd3_1 hold96 (.A(\c$ds_app_arg_1[16] ),
    .X(net138));
 sg13g2_dlygate4sd3_1 hold97 (.A(\c$ds_app_arg_1[0] ),
    .X(net139));
 sg13g2_dlygate4sd3_1 hold98 (.A(\c$case_scrut ),
    .X(net140));
 sg13g2_dlygate4sd3_1 hold99 (.A(_000_),
    .X(net141));
 sg13g2_dlygate4sd3_1 hold100 (.A(_057_),
    .X(net142));
 sg13g2_dlygate4sd3_1 hold101 (.A(\c$ds_app_arg_1[22] ),
    .X(net143));
 sg13g2_dlygate4sd3_1 hold102 (.A(_000_),
    .X(net144));
 sg13g2_dlygate4sd3_1 hold103 (.A(\s[3] ),
    .X(net145));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_fill_2 FILLER_14_406 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_252 ();
 sg13g2_decap_8 FILLER_15_259 ();
 sg13g2_decap_8 FILLER_15_266 ();
 sg13g2_decap_8 FILLER_15_273 ();
 sg13g2_decap_8 FILLER_15_280 ();
 sg13g2_decap_8 FILLER_15_287 ();
 sg13g2_decap_8 FILLER_15_294 ();
 sg13g2_decap_8 FILLER_15_301 ();
 sg13g2_decap_8 FILLER_15_308 ();
 sg13g2_decap_8 FILLER_15_315 ();
 sg13g2_decap_8 FILLER_15_322 ();
 sg13g2_decap_8 FILLER_15_329 ();
 sg13g2_decap_8 FILLER_15_336 ();
 sg13g2_decap_8 FILLER_15_343 ();
 sg13g2_decap_8 FILLER_15_350 ();
 sg13g2_decap_8 FILLER_15_357 ();
 sg13g2_decap_8 FILLER_15_364 ();
 sg13g2_decap_8 FILLER_15_371 ();
 sg13g2_decap_8 FILLER_15_378 ();
 sg13g2_decap_8 FILLER_15_385 ();
 sg13g2_decap_8 FILLER_15_392 ();
 sg13g2_decap_8 FILLER_15_399 ();
 sg13g2_fill_2 FILLER_15_406 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_decap_8 FILLER_16_217 ();
 sg13g2_decap_8 FILLER_16_224 ();
 sg13g2_decap_8 FILLER_16_231 ();
 sg13g2_decap_8 FILLER_16_238 ();
 sg13g2_decap_8 FILLER_16_245 ();
 sg13g2_decap_8 FILLER_16_252 ();
 sg13g2_decap_8 FILLER_16_259 ();
 sg13g2_decap_8 FILLER_16_266 ();
 sg13g2_decap_8 FILLER_16_273 ();
 sg13g2_decap_8 FILLER_16_280 ();
 sg13g2_decap_8 FILLER_16_287 ();
 sg13g2_decap_8 FILLER_16_294 ();
 sg13g2_decap_8 FILLER_16_301 ();
 sg13g2_decap_8 FILLER_16_308 ();
 sg13g2_decap_8 FILLER_16_315 ();
 sg13g2_decap_8 FILLER_16_322 ();
 sg13g2_decap_8 FILLER_16_329 ();
 sg13g2_decap_8 FILLER_16_336 ();
 sg13g2_decap_8 FILLER_16_343 ();
 sg13g2_decap_8 FILLER_16_350 ();
 sg13g2_decap_8 FILLER_16_357 ();
 sg13g2_decap_8 FILLER_16_364 ();
 sg13g2_decap_8 FILLER_16_371 ();
 sg13g2_decap_8 FILLER_16_378 ();
 sg13g2_decap_8 FILLER_16_385 ();
 sg13g2_decap_8 FILLER_16_392 ();
 sg13g2_decap_8 FILLER_16_399 ();
 sg13g2_fill_2 FILLER_16_406 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_decap_8 FILLER_17_168 ();
 sg13g2_decap_8 FILLER_17_175 ();
 sg13g2_decap_8 FILLER_17_182 ();
 sg13g2_decap_8 FILLER_17_189 ();
 sg13g2_decap_8 FILLER_17_196 ();
 sg13g2_decap_8 FILLER_17_203 ();
 sg13g2_decap_8 FILLER_17_210 ();
 sg13g2_decap_8 FILLER_17_217 ();
 sg13g2_decap_8 FILLER_17_224 ();
 sg13g2_decap_8 FILLER_17_231 ();
 sg13g2_decap_8 FILLER_17_238 ();
 sg13g2_decap_8 FILLER_17_245 ();
 sg13g2_decap_8 FILLER_17_252 ();
 sg13g2_decap_8 FILLER_17_259 ();
 sg13g2_decap_8 FILLER_17_266 ();
 sg13g2_decap_8 FILLER_17_273 ();
 sg13g2_decap_8 FILLER_17_280 ();
 sg13g2_decap_8 FILLER_17_287 ();
 sg13g2_decap_8 FILLER_17_294 ();
 sg13g2_decap_8 FILLER_17_301 ();
 sg13g2_decap_8 FILLER_17_308 ();
 sg13g2_decap_8 FILLER_17_315 ();
 sg13g2_decap_8 FILLER_17_322 ();
 sg13g2_decap_8 FILLER_17_329 ();
 sg13g2_decap_8 FILLER_17_336 ();
 sg13g2_decap_8 FILLER_17_343 ();
 sg13g2_decap_8 FILLER_17_350 ();
 sg13g2_decap_8 FILLER_17_357 ();
 sg13g2_decap_8 FILLER_17_364 ();
 sg13g2_decap_8 FILLER_17_371 ();
 sg13g2_decap_8 FILLER_17_378 ();
 sg13g2_decap_8 FILLER_17_385 ();
 sg13g2_decap_8 FILLER_17_392 ();
 sg13g2_decap_8 FILLER_17_399 ();
 sg13g2_fill_2 FILLER_17_406 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_decap_8 FILLER_18_147 ();
 sg13g2_decap_8 FILLER_18_154 ();
 sg13g2_decap_8 FILLER_18_161 ();
 sg13g2_decap_8 FILLER_18_168 ();
 sg13g2_decap_8 FILLER_18_175 ();
 sg13g2_decap_8 FILLER_18_182 ();
 sg13g2_decap_8 FILLER_18_189 ();
 sg13g2_decap_8 FILLER_18_196 ();
 sg13g2_decap_8 FILLER_18_203 ();
 sg13g2_decap_8 FILLER_18_210 ();
 sg13g2_decap_8 FILLER_18_217 ();
 sg13g2_decap_8 FILLER_18_224 ();
 sg13g2_decap_8 FILLER_18_231 ();
 sg13g2_decap_8 FILLER_18_238 ();
 sg13g2_decap_8 FILLER_18_245 ();
 sg13g2_decap_8 FILLER_18_252 ();
 sg13g2_decap_8 FILLER_18_259 ();
 sg13g2_decap_8 FILLER_18_266 ();
 sg13g2_decap_8 FILLER_18_273 ();
 sg13g2_decap_8 FILLER_18_280 ();
 sg13g2_decap_8 FILLER_18_287 ();
 sg13g2_decap_8 FILLER_18_294 ();
 sg13g2_decap_8 FILLER_18_301 ();
 sg13g2_decap_8 FILLER_18_308 ();
 sg13g2_decap_8 FILLER_18_315 ();
 sg13g2_decap_8 FILLER_18_322 ();
 sg13g2_decap_8 FILLER_18_329 ();
 sg13g2_decap_8 FILLER_18_336 ();
 sg13g2_decap_8 FILLER_18_343 ();
 sg13g2_decap_8 FILLER_18_350 ();
 sg13g2_decap_8 FILLER_18_357 ();
 sg13g2_decap_8 FILLER_18_364 ();
 sg13g2_decap_8 FILLER_18_371 ();
 sg13g2_decap_8 FILLER_18_378 ();
 sg13g2_decap_8 FILLER_18_385 ();
 sg13g2_decap_8 FILLER_18_392 ();
 sg13g2_decap_8 FILLER_18_399 ();
 sg13g2_fill_2 FILLER_18_406 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_decap_8 FILLER_19_140 ();
 sg13g2_decap_8 FILLER_19_147 ();
 sg13g2_decap_8 FILLER_19_154 ();
 sg13g2_decap_8 FILLER_19_161 ();
 sg13g2_decap_8 FILLER_19_168 ();
 sg13g2_decap_8 FILLER_19_175 ();
 sg13g2_decap_8 FILLER_19_182 ();
 sg13g2_decap_8 FILLER_19_189 ();
 sg13g2_decap_8 FILLER_19_196 ();
 sg13g2_decap_8 FILLER_19_203 ();
 sg13g2_decap_8 FILLER_19_210 ();
 sg13g2_decap_8 FILLER_19_217 ();
 sg13g2_decap_8 FILLER_19_224 ();
 sg13g2_decap_8 FILLER_19_231 ();
 sg13g2_decap_8 FILLER_19_238 ();
 sg13g2_decap_8 FILLER_19_245 ();
 sg13g2_decap_8 FILLER_19_252 ();
 sg13g2_decap_8 FILLER_19_259 ();
 sg13g2_decap_8 FILLER_19_266 ();
 sg13g2_decap_8 FILLER_19_273 ();
 sg13g2_decap_8 FILLER_19_280 ();
 sg13g2_decap_8 FILLER_19_287 ();
 sg13g2_decap_8 FILLER_19_294 ();
 sg13g2_decap_8 FILLER_19_301 ();
 sg13g2_decap_8 FILLER_19_308 ();
 sg13g2_decap_8 FILLER_19_315 ();
 sg13g2_decap_8 FILLER_19_322 ();
 sg13g2_decap_8 FILLER_19_329 ();
 sg13g2_decap_8 FILLER_19_336 ();
 sg13g2_decap_8 FILLER_19_343 ();
 sg13g2_decap_8 FILLER_19_350 ();
 sg13g2_decap_8 FILLER_19_357 ();
 sg13g2_decap_8 FILLER_19_364 ();
 sg13g2_decap_8 FILLER_19_371 ();
 sg13g2_decap_8 FILLER_19_378 ();
 sg13g2_decap_8 FILLER_19_385 ();
 sg13g2_decap_8 FILLER_19_392 ();
 sg13g2_decap_8 FILLER_19_399 ();
 sg13g2_fill_2 FILLER_19_406 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_decap_8 FILLER_20_126 ();
 sg13g2_decap_8 FILLER_20_133 ();
 sg13g2_decap_8 FILLER_20_140 ();
 sg13g2_decap_8 FILLER_20_147 ();
 sg13g2_decap_8 FILLER_20_154 ();
 sg13g2_decap_8 FILLER_20_161 ();
 sg13g2_decap_8 FILLER_20_168 ();
 sg13g2_decap_8 FILLER_20_175 ();
 sg13g2_decap_8 FILLER_20_182 ();
 sg13g2_decap_8 FILLER_20_189 ();
 sg13g2_decap_8 FILLER_20_196 ();
 sg13g2_decap_8 FILLER_20_203 ();
 sg13g2_decap_8 FILLER_20_210 ();
 sg13g2_decap_8 FILLER_20_217 ();
 sg13g2_decap_8 FILLER_20_224 ();
 sg13g2_decap_8 FILLER_20_231 ();
 sg13g2_decap_8 FILLER_20_238 ();
 sg13g2_decap_8 FILLER_20_245 ();
 sg13g2_decap_8 FILLER_20_252 ();
 sg13g2_decap_8 FILLER_20_259 ();
 sg13g2_decap_8 FILLER_20_266 ();
 sg13g2_decap_8 FILLER_20_273 ();
 sg13g2_decap_8 FILLER_20_280 ();
 sg13g2_decap_8 FILLER_20_287 ();
 sg13g2_decap_8 FILLER_20_294 ();
 sg13g2_decap_8 FILLER_20_301 ();
 sg13g2_decap_8 FILLER_20_308 ();
 sg13g2_decap_8 FILLER_20_315 ();
 sg13g2_decap_8 FILLER_20_322 ();
 sg13g2_decap_8 FILLER_20_329 ();
 sg13g2_decap_8 FILLER_20_336 ();
 sg13g2_decap_8 FILLER_20_343 ();
 sg13g2_decap_8 FILLER_20_350 ();
 sg13g2_decap_8 FILLER_20_357 ();
 sg13g2_decap_8 FILLER_20_364 ();
 sg13g2_decap_8 FILLER_20_371 ();
 sg13g2_decap_8 FILLER_20_378 ();
 sg13g2_decap_8 FILLER_20_385 ();
 sg13g2_decap_8 FILLER_20_392 ();
 sg13g2_decap_8 FILLER_20_399 ();
 sg13g2_fill_2 FILLER_20_406 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_decap_8 FILLER_21_119 ();
 sg13g2_decap_8 FILLER_21_126 ();
 sg13g2_decap_8 FILLER_21_133 ();
 sg13g2_decap_8 FILLER_21_140 ();
 sg13g2_decap_8 FILLER_21_147 ();
 sg13g2_decap_8 FILLER_21_154 ();
 sg13g2_decap_8 FILLER_21_161 ();
 sg13g2_decap_8 FILLER_21_168 ();
 sg13g2_decap_8 FILLER_21_175 ();
 sg13g2_decap_8 FILLER_21_182 ();
 sg13g2_decap_8 FILLER_21_189 ();
 sg13g2_decap_8 FILLER_21_196 ();
 sg13g2_decap_8 FILLER_21_203 ();
 sg13g2_decap_8 FILLER_21_210 ();
 sg13g2_decap_8 FILLER_21_217 ();
 sg13g2_decap_8 FILLER_21_224 ();
 sg13g2_decap_8 FILLER_21_231 ();
 sg13g2_fill_1 FILLER_21_238 ();
 sg13g2_decap_8 FILLER_21_242 ();
 sg13g2_decap_4 FILLER_21_249 ();
 sg13g2_decap_8 FILLER_21_262 ();
 sg13g2_decap_8 FILLER_21_269 ();
 sg13g2_decap_8 FILLER_21_276 ();
 sg13g2_decap_8 FILLER_21_283 ();
 sg13g2_decap_4 FILLER_21_290 ();
 sg13g2_decap_4 FILLER_21_298 ();
 sg13g2_fill_1 FILLER_21_302 ();
 sg13g2_decap_8 FILLER_21_312 ();
 sg13g2_decap_8 FILLER_21_319 ();
 sg13g2_decap_8 FILLER_21_326 ();
 sg13g2_decap_8 FILLER_21_333 ();
 sg13g2_decap_8 FILLER_21_340 ();
 sg13g2_decap_8 FILLER_21_347 ();
 sg13g2_decap_8 FILLER_21_354 ();
 sg13g2_decap_8 FILLER_21_361 ();
 sg13g2_decap_8 FILLER_21_368 ();
 sg13g2_decap_8 FILLER_21_375 ();
 sg13g2_decap_8 FILLER_21_382 ();
 sg13g2_decap_8 FILLER_21_389 ();
 sg13g2_decap_8 FILLER_21_396 ();
 sg13g2_decap_4 FILLER_21_403 ();
 sg13g2_fill_2 FILLER_21_407 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_8 FILLER_22_105 ();
 sg13g2_decap_8 FILLER_22_112 ();
 sg13g2_decap_8 FILLER_22_119 ();
 sg13g2_decap_8 FILLER_22_126 ();
 sg13g2_decap_8 FILLER_22_133 ();
 sg13g2_decap_8 FILLER_22_140 ();
 sg13g2_decap_8 FILLER_22_147 ();
 sg13g2_decap_8 FILLER_22_154 ();
 sg13g2_decap_8 FILLER_22_161 ();
 sg13g2_decap_8 FILLER_22_168 ();
 sg13g2_decap_8 FILLER_22_175 ();
 sg13g2_decap_8 FILLER_22_182 ();
 sg13g2_decap_8 FILLER_22_189 ();
 sg13g2_decap_4 FILLER_22_196 ();
 sg13g2_fill_2 FILLER_22_209 ();
 sg13g2_fill_1 FILLER_22_211 ();
 sg13g2_fill_1 FILLER_22_293 ();
 sg13g2_decap_8 FILLER_22_320 ();
 sg13g2_decap_8 FILLER_22_327 ();
 sg13g2_decap_8 FILLER_22_334 ();
 sg13g2_decap_8 FILLER_22_341 ();
 sg13g2_decap_8 FILLER_22_348 ();
 sg13g2_decap_8 FILLER_22_355 ();
 sg13g2_decap_8 FILLER_22_362 ();
 sg13g2_decap_8 FILLER_22_369 ();
 sg13g2_decap_8 FILLER_22_376 ();
 sg13g2_decap_8 FILLER_22_383 ();
 sg13g2_decap_8 FILLER_22_390 ();
 sg13g2_decap_8 FILLER_22_397 ();
 sg13g2_decap_4 FILLER_22_404 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_98 ();
 sg13g2_decap_8 FILLER_23_105 ();
 sg13g2_decap_8 FILLER_23_112 ();
 sg13g2_decap_8 FILLER_23_119 ();
 sg13g2_decap_8 FILLER_23_126 ();
 sg13g2_decap_8 FILLER_23_133 ();
 sg13g2_decap_8 FILLER_23_140 ();
 sg13g2_decap_8 FILLER_23_147 ();
 sg13g2_decap_8 FILLER_23_154 ();
 sg13g2_decap_8 FILLER_23_161 ();
 sg13g2_decap_8 FILLER_23_168 ();
 sg13g2_decap_8 FILLER_23_175 ();
 sg13g2_decap_4 FILLER_23_182 ();
 sg13g2_fill_1 FILLER_23_186 ();
 sg13g2_decap_4 FILLER_23_242 ();
 sg13g2_fill_2 FILLER_23_280 ();
 sg13g2_fill_2 FILLER_23_310 ();
 sg13g2_fill_2 FILLER_23_338 ();
 sg13g2_fill_1 FILLER_23_340 ();
 sg13g2_decap_8 FILLER_23_367 ();
 sg13g2_decap_8 FILLER_23_374 ();
 sg13g2_decap_8 FILLER_23_381 ();
 sg13g2_decap_8 FILLER_23_388 ();
 sg13g2_decap_8 FILLER_23_395 ();
 sg13g2_decap_8 FILLER_23_402 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_decap_8 FILLER_24_98 ();
 sg13g2_decap_8 FILLER_24_105 ();
 sg13g2_decap_8 FILLER_24_112 ();
 sg13g2_decap_8 FILLER_24_119 ();
 sg13g2_decap_8 FILLER_24_126 ();
 sg13g2_decap_8 FILLER_24_133 ();
 sg13g2_decap_8 FILLER_24_140 ();
 sg13g2_decap_4 FILLER_24_147 ();
 sg13g2_fill_2 FILLER_24_151 ();
 sg13g2_decap_4 FILLER_24_168 ();
 sg13g2_fill_2 FILLER_24_172 ();
 sg13g2_fill_1 FILLER_24_223 ();
 sg13g2_decap_4 FILLER_24_248 ();
 sg13g2_fill_1 FILLER_24_277 ();
 sg13g2_fill_2 FILLER_24_299 ();
 sg13g2_fill_1 FILLER_24_336 ();
 sg13g2_fill_2 FILLER_24_352 ();
 sg13g2_decap_8 FILLER_24_363 ();
 sg13g2_decap_8 FILLER_24_370 ();
 sg13g2_decap_8 FILLER_24_377 ();
 sg13g2_decap_8 FILLER_24_384 ();
 sg13g2_decap_8 FILLER_24_391 ();
 sg13g2_decap_8 FILLER_24_398 ();
 sg13g2_decap_4 FILLER_24_405 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_8 FILLER_25_91 ();
 sg13g2_decap_8 FILLER_25_98 ();
 sg13g2_decap_8 FILLER_25_105 ();
 sg13g2_decap_8 FILLER_25_112 ();
 sg13g2_decap_8 FILLER_25_119 ();
 sg13g2_decap_8 FILLER_25_126 ();
 sg13g2_decap_8 FILLER_25_133 ();
 sg13g2_fill_2 FILLER_25_140 ();
 sg13g2_fill_1 FILLER_25_142 ();
 sg13g2_decap_4 FILLER_25_182 ();
 sg13g2_fill_1 FILLER_25_186 ();
 sg13g2_fill_1 FILLER_25_225 ();
 sg13g2_fill_2 FILLER_25_242 ();
 sg13g2_fill_1 FILLER_25_276 ();
 sg13g2_fill_1 FILLER_25_304 ();
 sg13g2_decap_4 FILLER_25_321 ();
 sg13g2_fill_2 FILLER_25_334 ();
 sg13g2_fill_1 FILLER_25_346 ();
 sg13g2_fill_2 FILLER_25_357 ();
 sg13g2_fill_1 FILLER_25_359 ();
 sg13g2_decap_8 FILLER_25_386 ();
 sg13g2_decap_8 FILLER_25_393 ();
 sg13g2_decap_8 FILLER_25_400 ();
 sg13g2_fill_2 FILLER_25_407 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_decap_8 FILLER_26_91 ();
 sg13g2_decap_8 FILLER_26_98 ();
 sg13g2_decap_8 FILLER_26_105 ();
 sg13g2_decap_8 FILLER_26_112 ();
 sg13g2_decap_8 FILLER_26_119 ();
 sg13g2_decap_8 FILLER_26_126 ();
 sg13g2_decap_4 FILLER_26_133 ();
 sg13g2_fill_2 FILLER_26_163 ();
 sg13g2_fill_1 FILLER_26_191 ();
 sg13g2_fill_2 FILLER_26_245 ();
 sg13g2_fill_2 FILLER_26_266 ();
 sg13g2_fill_1 FILLER_26_268 ();
 sg13g2_decap_4 FILLER_26_275 ();
 sg13g2_fill_1 FILLER_26_279 ();
 sg13g2_fill_2 FILLER_26_306 ();
 sg13g2_fill_1 FILLER_26_359 ();
 sg13g2_decap_8 FILLER_26_386 ();
 sg13g2_decap_8 FILLER_26_393 ();
 sg13g2_decap_8 FILLER_26_400 ();
 sg13g2_fill_2 FILLER_26_407 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_decap_8 FILLER_27_84 ();
 sg13g2_decap_8 FILLER_27_91 ();
 sg13g2_decap_8 FILLER_27_98 ();
 sg13g2_decap_8 FILLER_27_105 ();
 sg13g2_decap_8 FILLER_27_112 ();
 sg13g2_fill_2 FILLER_27_119 ();
 sg13g2_fill_1 FILLER_27_121 ();
 sg13g2_fill_2 FILLER_27_253 ();
 sg13g2_fill_1 FILLER_27_255 ();
 sg13g2_fill_2 FILLER_27_267 ();
 sg13g2_fill_1 FILLER_27_269 ();
 sg13g2_fill_2 FILLER_27_275 ();
 sg13g2_fill_1 FILLER_27_282 ();
 sg13g2_decap_4 FILLER_27_290 ();
 sg13g2_fill_2 FILLER_27_294 ();
 sg13g2_fill_1 FILLER_27_309 ();
 sg13g2_fill_2 FILLER_27_320 ();
 sg13g2_fill_1 FILLER_27_322 ();
 sg13g2_decap_4 FILLER_27_363 ();
 sg13g2_fill_1 FILLER_27_367 ();
 sg13g2_decap_8 FILLER_27_386 ();
 sg13g2_decap_8 FILLER_27_393 ();
 sg13g2_decap_8 FILLER_27_400 ();
 sg13g2_fill_2 FILLER_27_407 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_decap_8 FILLER_28_84 ();
 sg13g2_decap_8 FILLER_28_91 ();
 sg13g2_decap_8 FILLER_28_98 ();
 sg13g2_decap_8 FILLER_28_105 ();
 sg13g2_decap_8 FILLER_28_112 ();
 sg13g2_fill_2 FILLER_28_119 ();
 sg13g2_fill_1 FILLER_28_121 ();
 sg13g2_fill_1 FILLER_28_187 ();
 sg13g2_decap_8 FILLER_28_207 ();
 sg13g2_decap_4 FILLER_28_214 ();
 sg13g2_fill_2 FILLER_28_218 ();
 sg13g2_fill_2 FILLER_28_310 ();
 sg13g2_fill_2 FILLER_28_335 ();
 sg13g2_decap_8 FILLER_28_387 ();
 sg13g2_decap_8 FILLER_28_394 ();
 sg13g2_decap_8 FILLER_28_401 ();
 sg13g2_fill_1 FILLER_28_408 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_decap_8 FILLER_29_84 ();
 sg13g2_decap_8 FILLER_29_91 ();
 sg13g2_decap_8 FILLER_29_98 ();
 sg13g2_decap_8 FILLER_29_105 ();
 sg13g2_decap_8 FILLER_29_112 ();
 sg13g2_decap_4 FILLER_29_119 ();
 sg13g2_fill_2 FILLER_29_149 ();
 sg13g2_fill_2 FILLER_29_160 ();
 sg13g2_decap_8 FILLER_29_214 ();
 sg13g2_decap_4 FILLER_29_221 ();
 sg13g2_fill_1 FILLER_29_225 ();
 sg13g2_decap_8 FILLER_29_234 ();
 sg13g2_fill_2 FILLER_29_241 ();
 sg13g2_fill_1 FILLER_29_243 ();
 sg13g2_fill_2 FILLER_29_274 ();
 sg13g2_fill_1 FILLER_29_307 ();
 sg13g2_fill_1 FILLER_29_361 ();
 sg13g2_decap_8 FILLER_29_388 ();
 sg13g2_decap_8 FILLER_29_395 ();
 sg13g2_decap_8 FILLER_29_402 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_77 ();
 sg13g2_decap_8 FILLER_30_84 ();
 sg13g2_decap_8 FILLER_30_91 ();
 sg13g2_decap_8 FILLER_30_98 ();
 sg13g2_decap_8 FILLER_30_105 ();
 sg13g2_decap_8 FILLER_30_112 ();
 sg13g2_decap_4 FILLER_30_119 ();
 sg13g2_fill_1 FILLER_30_123 ();
 sg13g2_fill_2 FILLER_30_162 ();
 sg13g2_fill_1 FILLER_30_295 ();
 sg13g2_fill_2 FILLER_30_300 ();
 sg13g2_decap_8 FILLER_30_389 ();
 sg13g2_decap_8 FILLER_30_396 ();
 sg13g2_decap_4 FILLER_30_403 ();
 sg13g2_fill_2 FILLER_30_407 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_decap_8 FILLER_31_84 ();
 sg13g2_decap_8 FILLER_31_91 ();
 sg13g2_decap_8 FILLER_31_98 ();
 sg13g2_decap_8 FILLER_31_105 ();
 sg13g2_decap_4 FILLER_31_112 ();
 sg13g2_fill_1 FILLER_31_175 ();
 sg13g2_fill_2 FILLER_31_199 ();
 sg13g2_decap_8 FILLER_31_209 ();
 sg13g2_fill_1 FILLER_31_216 ();
 sg13g2_fill_1 FILLER_31_221 ();
 sg13g2_decap_8 FILLER_31_227 ();
 sg13g2_decap_4 FILLER_31_234 ();
 sg13g2_fill_1 FILLER_31_238 ();
 sg13g2_fill_2 FILLER_31_249 ();
 sg13g2_fill_1 FILLER_31_251 ();
 sg13g2_fill_2 FILLER_31_266 ();
 sg13g2_fill_2 FILLER_31_321 ();
 sg13g2_decap_4 FILLER_31_405 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_8 FILLER_32_84 ();
 sg13g2_decap_8 FILLER_32_91 ();
 sg13g2_decap_8 FILLER_32_98 ();
 sg13g2_decap_8 FILLER_32_105 ();
 sg13g2_decap_8 FILLER_32_112 ();
 sg13g2_fill_1 FILLER_32_199 ();
 sg13g2_fill_1 FILLER_32_288 ();
 sg13g2_fill_2 FILLER_32_297 ();
 sg13g2_fill_1 FILLER_32_325 ();
 sg13g2_fill_1 FILLER_32_344 ();
 sg13g2_fill_2 FILLER_32_406 ();
 sg13g2_fill_1 FILLER_32_408 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_decap_8 FILLER_33_91 ();
 sg13g2_decap_8 FILLER_33_98 ();
 sg13g2_decap_8 FILLER_33_105 ();
 sg13g2_decap_8 FILLER_33_112 ();
 sg13g2_decap_8 FILLER_33_119 ();
 sg13g2_fill_2 FILLER_33_126 ();
 sg13g2_fill_1 FILLER_33_128 ();
 sg13g2_fill_1 FILLER_33_132 ();
 sg13g2_fill_1 FILLER_33_152 ();
 sg13g2_fill_2 FILLER_33_206 ();
 sg13g2_decap_8 FILLER_33_217 ();
 sg13g2_decap_8 FILLER_33_224 ();
 sg13g2_decap_4 FILLER_33_231 ();
 sg13g2_fill_1 FILLER_33_247 ();
 sg13g2_fill_1 FILLER_33_274 ();
 sg13g2_fill_2 FILLER_33_289 ();
 sg13g2_fill_2 FILLER_33_305 ();
 sg13g2_fill_1 FILLER_33_364 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_decap_8 FILLER_34_91 ();
 sg13g2_decap_8 FILLER_34_98 ();
 sg13g2_decap_8 FILLER_34_105 ();
 sg13g2_decap_8 FILLER_34_112 ();
 sg13g2_decap_8 FILLER_34_119 ();
 sg13g2_fill_2 FILLER_34_152 ();
 sg13g2_decap_8 FILLER_34_220 ();
 sg13g2_fill_1 FILLER_34_227 ();
 sg13g2_fill_1 FILLER_34_367 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_decap_8 FILLER_35_98 ();
 sg13g2_decap_8 FILLER_35_105 ();
 sg13g2_decap_8 FILLER_35_112 ();
 sg13g2_decap_8 FILLER_35_119 ();
 sg13g2_decap_8 FILLER_35_126 ();
 sg13g2_decap_8 FILLER_35_133 ();
 sg13g2_decap_8 FILLER_35_140 ();
 sg13g2_fill_1 FILLER_35_147 ();
 sg13g2_fill_1 FILLER_35_151 ();
 sg13g2_fill_2 FILLER_35_158 ();
 sg13g2_fill_1 FILLER_35_172 ();
 sg13g2_decap_8 FILLER_35_189 ();
 sg13g2_decap_8 FILLER_35_196 ();
 sg13g2_decap_8 FILLER_35_203 ();
 sg13g2_fill_1 FILLER_35_210 ();
 sg13g2_fill_1 FILLER_35_289 ();
 sg13g2_fill_1 FILLER_35_304 ();
 sg13g2_fill_2 FILLER_35_324 ();
 sg13g2_fill_2 FILLER_35_368 ();
 sg13g2_fill_2 FILLER_35_379 ();
 sg13g2_fill_2 FILLER_35_407 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_decap_8 FILLER_36_112 ();
 sg13g2_decap_8 FILLER_36_119 ();
 sg13g2_decap_8 FILLER_36_126 ();
 sg13g2_decap_8 FILLER_36_133 ();
 sg13g2_decap_8 FILLER_36_140 ();
 sg13g2_decap_8 FILLER_36_147 ();
 sg13g2_fill_2 FILLER_36_154 ();
 sg13g2_fill_1 FILLER_36_156 ();
 sg13g2_decap_4 FILLER_36_160 ();
 sg13g2_fill_1 FILLER_36_164 ();
 sg13g2_decap_8 FILLER_36_170 ();
 sg13g2_decap_8 FILLER_36_177 ();
 sg13g2_decap_8 FILLER_36_184 ();
 sg13g2_decap_8 FILLER_36_191 ();
 sg13g2_fill_1 FILLER_36_198 ();
 sg13g2_fill_1 FILLER_36_256 ();
 sg13g2_fill_1 FILLER_36_266 ();
 sg13g2_fill_2 FILLER_36_294 ();
 sg13g2_fill_1 FILLER_36_353 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_8 FILLER_37_112 ();
 sg13g2_decap_8 FILLER_37_119 ();
 sg13g2_decap_8 FILLER_37_126 ();
 sg13g2_decap_8 FILLER_37_133 ();
 sg13g2_decap_8 FILLER_37_140 ();
 sg13g2_decap_8 FILLER_37_147 ();
 sg13g2_decap_8 FILLER_37_154 ();
 sg13g2_decap_8 FILLER_37_161 ();
 sg13g2_decap_8 FILLER_37_168 ();
 sg13g2_decap_8 FILLER_37_175 ();
 sg13g2_decap_8 FILLER_37_182 ();
 sg13g2_decap_8 FILLER_37_189 ();
 sg13g2_decap_8 FILLER_37_196 ();
 sg13g2_decap_4 FILLER_37_203 ();
 sg13g2_fill_2 FILLER_37_295 ();
 sg13g2_fill_2 FILLER_37_357 ();
 sg13g2_fill_2 FILLER_37_396 ();
 sg13g2_fill_2 FILLER_37_407 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_4 FILLER_38_60 ();
 sg13g2_decap_4 FILLER_38_68 ();
 sg13g2_decap_4 FILLER_38_76 ();
 sg13g2_decap_4 FILLER_38_84 ();
 sg13g2_decap_4 FILLER_38_92 ();
 sg13g2_decap_4 FILLER_38_100 ();
 sg13g2_decap_4 FILLER_38_108 ();
 sg13g2_decap_4 FILLER_38_116 ();
 sg13g2_decap_4 FILLER_38_124 ();
 sg13g2_decap_4 FILLER_38_132 ();
 sg13g2_decap_4 FILLER_38_140 ();
 sg13g2_decap_4 FILLER_38_148 ();
 sg13g2_decap_4 FILLER_38_156 ();
 sg13g2_decap_4 FILLER_38_164 ();
 sg13g2_decap_4 FILLER_38_172 ();
 sg13g2_decap_8 FILLER_38_180 ();
 sg13g2_decap_4 FILLER_38_187 ();
 sg13g2_fill_1 FILLER_38_191 ();
 sg13g2_decap_8 FILLER_38_196 ();
 sg13g2_fill_1 FILLER_38_203 ();
 sg13g2_fill_2 FILLER_38_252 ();
 sg13g2_fill_1 FILLER_38_270 ();
 sg13g2_fill_2 FILLER_38_333 ();
 sg13g2_fill_2 FILLER_38_370 ();
 sg13g2_fill_2 FILLER_38_407 ();
 assign uio_oe[0] = net9;
 assign uio_oe[1] = net10;
 assign uio_oe[2] = net11;
 assign uio_oe[3] = net12;
 assign uio_oe[4] = net13;
 assign uio_oe[5] = net14;
 assign uio_oe[6] = net15;
 assign uio_oe[7] = net16;
 assign uio_out[0] = net17;
 assign uio_out[1] = net18;
 assign uio_out[2] = net19;
 assign uio_out[3] = net20;
 assign uio_out[4] = net21;
 assign uio_out[5] = net22;
 assign uio_out[6] = net23;
 assign uio_out[7] = net24;
 assign uo_out[6] = net25;
endmodule

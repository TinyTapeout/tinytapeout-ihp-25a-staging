module tt_um_rebeccargb_intercal_alu (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire clknet_0_clk;
 wire \a[0] ;
 wire \a[10] ;
 wire \a[11] ;
 wire \a[12] ;
 wire \a[13] ;
 wire \a[14] ;
 wire \a[15] ;
 wire \a[16] ;
 wire \a[17] ;
 wire \a[18] ;
 wire \a[19] ;
 wire \a[1] ;
 wire \a[20] ;
 wire \a[21] ;
 wire \a[22] ;
 wire \a[23] ;
 wire \a[24] ;
 wire \a[25] ;
 wire \a[26] ;
 wire \a[27] ;
 wire \a[28] ;
 wire \a[29] ;
 wire \a[2] ;
 wire \a[30] ;
 wire \a[31] ;
 wire \a[3] ;
 wire \a[4] ;
 wire \a[5] ;
 wire \a[6] ;
 wire \a[7] ;
 wire \a[8] ;
 wire \a[9] ;
 wire \ayayayayayaya.b[0] ;
 wire \ayayayayayaya.b[10] ;
 wire \ayayayayayaya.b[11] ;
 wire \ayayayayayaya.b[12] ;
 wire \ayayayayayaya.b[13] ;
 wire \ayayayayayaya.b[14] ;
 wire \ayayayayayaya.b[15] ;
 wire \ayayayayayaya.b[16] ;
 wire \ayayayayayaya.b[17] ;
 wire \ayayayayayaya.b[18] ;
 wire \ayayayayayaya.b[19] ;
 wire \ayayayayayaya.b[1] ;
 wire \ayayayayayaya.b[20] ;
 wire \ayayayayayaya.b[21] ;
 wire \ayayayayayaya.b[22] ;
 wire \ayayayayayaya.b[23] ;
 wire \ayayayayayaya.b[24] ;
 wire \ayayayayayaya.b[25] ;
 wire \ayayayayayaya.b[26] ;
 wire \ayayayayayaya.b[27] ;
 wire \ayayayayayaya.b[28] ;
 wire \ayayayayayaya.b[29] ;
 wire \ayayayayayaya.b[2] ;
 wire \ayayayayayaya.b[30] ;
 wire \ayayayayayaya.b[31] ;
 wire \ayayayayayaya.b[3] ;
 wire \ayayayayayaya.b[4] ;
 wire \ayayayayayaya.b[5] ;
 wire \ayayayayayaya.b[6] ;
 wire \ayayayayayaya.b[7] ;
 wire \ayayayayayaya.b[8] ;
 wire \ayayayayayaya.b[9] ;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;

 sg13g2_inv_1 _1851_ (.Y(_0998_),
    .A(net1));
 sg13g2_inv_1 _1852_ (.Y(_0999_),
    .A(net1106));
 sg13g2_inv_1 _1853_ (.Y(_1000_),
    .A(\a[13] ));
 sg13g2_inv_1 _1854_ (.Y(_1001_),
    .A(net113));
 sg13g2_inv_1 _1855_ (.Y(_1002_),
    .A(\ayayayayayaya.b[28] ));
 sg13g2_inv_2 _1856_ (.Y(_1003_),
    .A(\ayayayayayaya.b[27] ));
 sg13g2_inv_2 _1857_ (.Y(_1004_),
    .A(\ayayayayayaya.b[26] ));
 sg13g2_inv_2 _1858_ (.Y(_1005_),
    .A(net104));
 sg13g2_inv_4 _1859_ (.A(net98),
    .Y(_1006_));
 sg13g2_inv_4 _1860_ (.A(net970),
    .Y(_1007_));
 sg13g2_inv_1 _1861_ (.Y(_1008_),
    .A(net972));
 sg13g2_inv_1 _1862_ (.Y(_1009_),
    .A(net975));
 sg13g2_inv_1 _1863_ (.Y(_1010_),
    .A(net977));
 sg13g2_inv_1 _1864_ (.Y(_1011_),
    .A(net980));
 sg13g2_inv_1 _1865_ (.Y(_1012_),
    .A(net982));
 sg13g2_inv_1 _1866_ (.Y(_1013_),
    .A(net984));
 sg13g2_inv_1 _1867_ (.Y(_1014_),
    .A(net987));
 sg13g2_inv_1 _1868_ (.Y(_1015_),
    .A(net989));
 sg13g2_inv_1 _1869_ (.Y(_1016_),
    .A(net993));
 sg13g2_inv_1 _1870_ (.Y(_1017_),
    .A(net996));
 sg13g2_inv_1 _1871_ (.Y(_1018_),
    .A(net1000));
 sg13g2_inv_1 _1872_ (.Y(_1019_),
    .A(net1003));
 sg13g2_inv_1 _1873_ (.Y(_1020_),
    .A(net1010));
 sg13g2_inv_1 _1874_ (.Y(_1021_),
    .A(net1015));
 sg13g2_inv_1 _1875_ (.Y(_1022_),
    .A(net1020));
 sg13g2_inv_1 _1876_ (.Y(_1023_),
    .A(net1023));
 sg13g2_inv_1 _1877_ (.Y(_1024_),
    .A(net1029));
 sg13g2_inv_1 _1878_ (.Y(_1025_),
    .A(net1036));
 sg13g2_inv_1 _1879_ (.Y(_1026_),
    .A(net1043));
 sg13g2_inv_1 _1880_ (.Y(_1027_),
    .A(net1052));
 sg13g2_inv_1 _1881_ (.Y(_1028_),
    .A(net1059));
 sg13g2_inv_1 _1882_ (.Y(_1029_),
    .A(net1067));
 sg13g2_inv_1 _1883_ (.Y(_1030_),
    .A(net1074));
 sg13g2_inv_1 _1884_ (.Y(_1031_),
    .A(_0053_));
 sg13g2_inv_2 _1885_ (.Y(uio_oe[7]),
    .A(net5));
 sg13g2_nand3_1 _1886_ (.B(\ayayayayayaya.b[31] ),
    .C(\ayayayayayaya.b[30] ),
    .A(net1084),
    .Y(_1032_));
 sg13g2_or2_2 _1887_ (.X(_1033_),
    .B(_1032_),
    .A(_1001_));
 sg13g2_nor2_1 _1888_ (.A(_0059_),
    .B(_1033_),
    .Y(_1034_));
 sg13g2_nor4_2 _1889_ (.A(_0059_),
    .B(_0058_),
    .C(_0057_),
    .Y(_1035_),
    .D(_1033_));
 sg13g2_nand3b_1 _1890_ (.B(\ayayayayayaya.b[31] ),
    .C(net1084),
    .Y(_1036_),
    .A_N(\ayayayayayaya.b[30] ));
 sg13g2_nand2b_1 _1891_ (.Y(_1037_),
    .B(\ayayayayayaya.b[30] ),
    .A_N(_0030_));
 sg13g2_and3_1 _1892_ (.X(_1038_),
    .A(\ayayayayayaya.b[29] ),
    .B(_1036_),
    .C(_1037_));
 sg13g2_and2_1 _1893_ (.A(_1001_),
    .B(_1032_),
    .X(_1039_));
 sg13g2_nor2_1 _1894_ (.A(\ayayayayayaya.b[28] ),
    .B(_1033_),
    .Y(_1040_));
 sg13g2_nor3_2 _1895_ (.A(_1002_),
    .B(_1038_),
    .C(_1039_),
    .Y(_1041_));
 sg13g2_nor3_2 _1896_ (.A(_1003_),
    .B(_1040_),
    .C(_1041_),
    .Y(_1042_));
 sg13g2_nor2_1 _1897_ (.A(\ayayayayayaya.b[27] ),
    .B(_1034_),
    .Y(_1043_));
 sg13g2_nor4_2 _1898_ (.A(\ayayayayayaya.b[26] ),
    .B(_0059_),
    .C(_0058_),
    .Y(_1044_),
    .D(_1033_));
 sg13g2_nor3_2 _1899_ (.A(_1004_),
    .B(_1042_),
    .C(_1043_),
    .Y(_1045_));
 sg13g2_nor3_2 _1900_ (.A(_1005_),
    .B(_1044_),
    .C(_1045_),
    .Y(_1046_));
 sg13g2_nor2_1 _1901_ (.A(\ayayayayayaya.b[25] ),
    .B(_1035_),
    .Y(_1047_));
 sg13g2_nand2b_2 _1902_ (.Y(_1048_),
    .B(_1035_),
    .A_N(_0056_));
 sg13g2_nor2_1 _1903_ (.A(\ayayayayayaya.b[24] ),
    .B(_1048_),
    .Y(_1049_));
 sg13g2_nor3_2 _1904_ (.A(_1006_),
    .B(_1046_),
    .C(_1047_),
    .Y(_1050_));
 sg13g2_and2_1 _1905_ (.A(_0029_),
    .B(\ayayayayayaya.b[29] ),
    .X(_1051_));
 sg13g2_and3_1 _1906_ (.X(_1052_),
    .A(_1001_),
    .B(_1036_),
    .C(_1037_));
 sg13g2_nor3_2 _1907_ (.A(\ayayayayayaya.b[28] ),
    .B(_1038_),
    .C(_1039_),
    .Y(_1053_));
 sg13g2_nor3_2 _1908_ (.A(_1002_),
    .B(_1051_),
    .C(_1052_),
    .Y(_1054_));
 sg13g2_nor3_2 _1909_ (.A(_1003_),
    .B(_1053_),
    .C(_1054_),
    .Y(_1055_));
 sg13g2_nor3_2 _1910_ (.A(\ayayayayayaya.b[27] ),
    .B(_1040_),
    .C(_1041_),
    .Y(_1056_));
 sg13g2_nor3_2 _1911_ (.A(\ayayayayayaya.b[26] ),
    .B(_1042_),
    .C(_1043_),
    .Y(_1057_));
 sg13g2_nor3_2 _1912_ (.A(_1004_),
    .B(_1055_),
    .C(_1056_),
    .Y(_1058_));
 sg13g2_nor3_2 _1913_ (.A(_1005_),
    .B(_1057_),
    .C(_1058_),
    .Y(_1059_));
 sg13g2_nor3_2 _1914_ (.A(net968),
    .B(_1044_),
    .C(_1045_),
    .Y(_1060_));
 sg13g2_nor3_2 _1915_ (.A(net969),
    .B(_1046_),
    .C(_1047_),
    .Y(_1061_));
 sg13g2_nor3_2 _1916_ (.A(_1006_),
    .B(_1059_),
    .C(_1060_),
    .Y(_1062_));
 sg13g2_nor3_2 _1917_ (.A(_1007_),
    .B(_1061_),
    .C(_1062_),
    .Y(_1063_));
 sg13g2_nor3_2 _1918_ (.A(net971),
    .B(_1049_),
    .C(_1050_),
    .Y(_1064_));
 sg13g2_nor2_1 _1919_ (.A(_0055_),
    .B(_1048_),
    .Y(_1065_));
 sg13g2_nor3_2 _1920_ (.A(_1007_),
    .B(_1049_),
    .C(_1050_),
    .Y(_1066_));
 sg13g2_nor2_2 _1921_ (.A(net970),
    .B(_1065_),
    .Y(_1067_));
 sg13g2_nor3_2 _1922_ (.A(net973),
    .B(_1066_),
    .C(_1067_),
    .Y(_1068_));
 sg13g2_nor3_2 _1923_ (.A(net967),
    .B(_1063_),
    .C(_1064_),
    .Y(_1069_));
 sg13g2_nor3_2 _1924_ (.A(\ayayayayayaya.b[28] ),
    .B(_1051_),
    .C(_1052_),
    .Y(_1070_));
 sg13g2_nor2_1 _1925_ (.A(_0028_),
    .B(_1002_),
    .Y(_1071_));
 sg13g2_nor3_2 _1926_ (.A(_1003_),
    .B(_1070_),
    .C(_1071_),
    .Y(_1072_));
 sg13g2_nor3_2 _1927_ (.A(\ayayayayayaya.b[27] ),
    .B(_1053_),
    .C(_1054_),
    .Y(_1073_));
 sg13g2_nor3_2 _1928_ (.A(\ayayayayayaya.b[26] ),
    .B(_1055_),
    .C(_1056_),
    .Y(_1074_));
 sg13g2_nor3_2 _1929_ (.A(_1004_),
    .B(_1072_),
    .C(_1073_),
    .Y(_1075_));
 sg13g2_nor3_2 _1930_ (.A(_1005_),
    .B(_1074_),
    .C(_1075_),
    .Y(_1076_));
 sg13g2_nor3_2 _1931_ (.A(net968),
    .B(_1057_),
    .C(_1058_),
    .Y(_1077_));
 sg13g2_nor3_2 _1932_ (.A(net969),
    .B(_1059_),
    .C(_1060_),
    .Y(_1078_));
 sg13g2_nor3_2 _1933_ (.A(_1006_),
    .B(_1076_),
    .C(_1077_),
    .Y(_1079_));
 sg13g2_nor3_2 _1934_ (.A(_1007_),
    .B(_1078_),
    .C(_1079_),
    .Y(_1080_));
 sg13g2_nor3_2 _1935_ (.A(net970),
    .B(_1061_),
    .C(_1062_),
    .Y(_1081_));
 sg13g2_nor3_2 _1936_ (.A(net972),
    .B(_1063_),
    .C(_1064_),
    .Y(_1082_));
 sg13g2_nor3_2 _1937_ (.A(net967),
    .B(_1080_),
    .C(_1081_),
    .Y(_1083_));
 sg13g2_nor3_2 _1938_ (.A(net966),
    .B(_1082_),
    .C(_1083_),
    .Y(_1084_));
 sg13g2_nor3_2 _1939_ (.A(net974),
    .B(_1068_),
    .C(_1069_),
    .Y(_1085_));
 sg13g2_nor3_2 _1940_ (.A(_0055_),
    .B(_0054_),
    .C(_1048_),
    .Y(_1086_));
 sg13g2_inv_1 _1941_ (.Y(_1087_),
    .A(_1086_));
 sg13g2_nor2_1 _1942_ (.A(net972),
    .B(_1087_),
    .Y(_1088_));
 sg13g2_nor3_2 _1943_ (.A(_1008_),
    .B(_1066_),
    .C(_1067_),
    .Y(_1089_));
 sg13g2_nor3_2 _1944_ (.A(net966),
    .B(_1068_),
    .C(_1069_),
    .Y(_1090_));
 sg13g2_nor3_2 _1945_ (.A(net974),
    .B(_1088_),
    .C(_1089_),
    .Y(_1091_));
 sg13g2_nor3_2 _1946_ (.A(net977),
    .B(_1090_),
    .C(_1091_),
    .Y(_1092_));
 sg13g2_nor3_2 _1947_ (.A(net965),
    .B(_1084_),
    .C(_1085_),
    .Y(_1093_));
 sg13g2_and2_1 _1948_ (.A(_0027_),
    .B(\ayayayayayaya.b[27] ),
    .X(_1094_));
 sg13g2_nor3_2 _1949_ (.A(\ayayayayayaya.b[27] ),
    .B(_1070_),
    .C(_1071_),
    .Y(_1095_));
 sg13g2_nor3_2 _1950_ (.A(\ayayayayayaya.b[26] ),
    .B(_1072_),
    .C(_1073_),
    .Y(_1096_));
 sg13g2_nor3_2 _1951_ (.A(_1004_),
    .B(_1094_),
    .C(_1095_),
    .Y(_1097_));
 sg13g2_nor3_2 _1952_ (.A(_1005_),
    .B(_1096_),
    .C(_1097_),
    .Y(_1098_));
 sg13g2_nor3_2 _1953_ (.A(net968),
    .B(_1074_),
    .C(_1075_),
    .Y(_1099_));
 sg13g2_nor3_2 _1954_ (.A(net969),
    .B(_1076_),
    .C(_1077_),
    .Y(_1100_));
 sg13g2_nor3_2 _1955_ (.A(_1006_),
    .B(_1098_),
    .C(_1099_),
    .Y(_1101_));
 sg13g2_nor3_2 _1956_ (.A(_1007_),
    .B(_1100_),
    .C(_1101_),
    .Y(_1102_));
 sg13g2_nor3_2 _1957_ (.A(net970),
    .B(_1078_),
    .C(_1079_),
    .Y(_1103_));
 sg13g2_nor3_2 _1958_ (.A(net972),
    .B(_1080_),
    .C(_1081_),
    .Y(_1104_));
 sg13g2_nor3_2 _1959_ (.A(net967),
    .B(_1102_),
    .C(_1103_),
    .Y(_1105_));
 sg13g2_nor3_2 _1960_ (.A(_1009_),
    .B(_1104_),
    .C(_1105_),
    .Y(_1106_));
 sg13g2_nor3_2 _1961_ (.A(net975),
    .B(_1082_),
    .C(_1083_),
    .Y(_1107_));
 sg13g2_nor3_2 _1962_ (.A(net978),
    .B(_1084_),
    .C(_1085_),
    .Y(_1108_));
 sg13g2_nor3_2 _1963_ (.A(_1010_),
    .B(_1106_),
    .C(_1107_),
    .Y(_1109_));
 sg13g2_nor3_2 _1964_ (.A(net963),
    .B(_1108_),
    .C(_1109_),
    .Y(_1110_));
 sg13g2_nor3_2 _1965_ (.A(net979),
    .B(_1092_),
    .C(_1093_),
    .Y(_1111_));
 sg13g2_a21oi_1 _1966_ (.A1(_1031_),
    .A2(_1086_),
    .Y(_1112_),
    .B1(net974));
 sg13g2_nor3_2 _1967_ (.A(net966),
    .B(_1088_),
    .C(_1089_),
    .Y(_1113_));
 sg13g2_nor3_2 _1968_ (.A(net977),
    .B(_1112_),
    .C(_1113_),
    .Y(_1114_));
 sg13g2_nor3_2 _1969_ (.A(_1010_),
    .B(_1090_),
    .C(_1091_),
    .Y(_1115_));
 sg13g2_nor3_2 _1970_ (.A(net964),
    .B(_1092_),
    .C(_1093_),
    .Y(_1116_));
 sg13g2_nor3_2 _1971_ (.A(net979),
    .B(_1114_),
    .C(_1115_),
    .Y(_1117_));
 sg13g2_nor3_2 _1972_ (.A(net982),
    .B(_1116_),
    .C(_1117_),
    .Y(_1118_));
 sg13g2_nor3_2 _1973_ (.A(net962),
    .B(_1110_),
    .C(_1111_),
    .Y(_1119_));
 sg13g2_nand2_1 _1974_ (.Y(_1120_),
    .A(_0026_),
    .B(\ayayayayayaya.b[26] ));
 sg13g2_o21ai_1 _1975_ (.B1(_1004_),
    .Y(_1121_),
    .A1(_1094_),
    .A2(_1095_));
 sg13g2_a21oi_1 _1976_ (.A1(_1120_),
    .A2(_1121_),
    .Y(_1122_),
    .B1(_1005_));
 sg13g2_nor3_2 _1977_ (.A(net968),
    .B(_1096_),
    .C(_1097_),
    .Y(_1123_));
 sg13g2_nor3_2 _1978_ (.A(net969),
    .B(_1098_),
    .C(_1099_),
    .Y(_1124_));
 sg13g2_nor3_2 _1979_ (.A(_1006_),
    .B(_1122_),
    .C(_1123_),
    .Y(_1125_));
 sg13g2_nor3_2 _1980_ (.A(_1007_),
    .B(_1124_),
    .C(_1125_),
    .Y(_1126_));
 sg13g2_nor3_2 _1981_ (.A(net970),
    .B(_1100_),
    .C(_1101_),
    .Y(_1127_));
 sg13g2_nor3_2 _1982_ (.A(net972),
    .B(_1102_),
    .C(_1103_),
    .Y(_1128_));
 sg13g2_nor3_2 _1983_ (.A(net967),
    .B(_1126_),
    .C(_1127_),
    .Y(_1129_));
 sg13g2_nor3_2 _1984_ (.A(net966),
    .B(_1128_),
    .C(_1129_),
    .Y(_1130_));
 sg13g2_nor3_2 _1985_ (.A(net975),
    .B(_1104_),
    .C(_1105_),
    .Y(_1131_));
 sg13g2_nor3_2 _1986_ (.A(net978),
    .B(_1106_),
    .C(_1107_),
    .Y(_1132_));
 sg13g2_nor3_2 _1987_ (.A(net965),
    .B(_1130_),
    .C(_1131_),
    .Y(_1133_));
 sg13g2_nor3_2 _1988_ (.A(net963),
    .B(_1132_),
    .C(_1133_),
    .Y(_1134_));
 sg13g2_nor3_2 _1989_ (.A(net979),
    .B(_1108_),
    .C(_1109_),
    .Y(_1135_));
 sg13g2_nor3_2 _1990_ (.A(net981),
    .B(_1110_),
    .C(_1111_),
    .Y(_1136_));
 sg13g2_nor3_2 _1991_ (.A(net962),
    .B(_1134_),
    .C(_1135_),
    .Y(_1137_));
 sg13g2_nor3_2 _1992_ (.A(net960),
    .B(_1136_),
    .C(_1137_),
    .Y(_1138_));
 sg13g2_nor3_2 _1993_ (.A(net984),
    .B(_1118_),
    .C(_1119_),
    .Y(_1139_));
 sg13g2_nor3_1 _1994_ (.A(_0053_),
    .B(_0052_),
    .C(_1087_),
    .Y(_1140_));
 sg13g2_or2_1 _1995_ (.X(_1141_),
    .B(_1140_),
    .A(net977));
 sg13g2_o21ai_1 _1996_ (.B1(net977),
    .Y(_1142_),
    .A1(_1112_),
    .A2(_1113_));
 sg13g2_nor3_2 _1997_ (.A(net964),
    .B(_1114_),
    .C(_1115_),
    .Y(_1143_));
 sg13g2_a21oi_2 _1998_ (.B1(net980),
    .Y(_1144_),
    .A2(_1142_),
    .A1(_1141_));
 sg13g2_nor3_2 _1999_ (.A(net981),
    .B(_1143_),
    .C(_1144_),
    .Y(_1145_));
 sg13g2_nor3_2 _2000_ (.A(net962),
    .B(_1116_),
    .C(_1117_),
    .Y(_1146_));
 sg13g2_nor3_2 _2001_ (.A(net960),
    .B(_1118_),
    .C(_1119_),
    .Y(_1147_));
 sg13g2_nor3_2 _2002_ (.A(net983),
    .B(_1145_),
    .C(_1146_),
    .Y(_1148_));
 sg13g2_nor3_2 _2003_ (.A(net986),
    .B(_1147_),
    .C(_1148_),
    .Y(_1149_));
 sg13g2_nor3_2 _2004_ (.A(net958),
    .B(_1138_),
    .C(_1139_),
    .Y(_1150_));
 sg13g2_and2_1 _2005_ (.A(_0025_),
    .B(net968),
    .X(_1151_));
 sg13g2_a21oi_1 _2006_ (.A1(_1120_),
    .A2(_1121_),
    .Y(_1152_),
    .B1(net968));
 sg13g2_nor3_1 _2007_ (.A(net969),
    .B(_1122_),
    .C(_1123_),
    .Y(_1153_));
 sg13g2_nor3_1 _2008_ (.A(_1006_),
    .B(_1151_),
    .C(_1152_),
    .Y(_1154_));
 sg13g2_nor3_1 _2009_ (.A(_1007_),
    .B(_1153_),
    .C(_1154_),
    .Y(_1155_));
 sg13g2_nor3_1 _2010_ (.A(net970),
    .B(_1124_),
    .C(_1125_),
    .Y(_1156_));
 sg13g2_nor3_2 _2011_ (.A(net972),
    .B(_1126_),
    .C(_1127_),
    .Y(_1157_));
 sg13g2_nor3_2 _2012_ (.A(net967),
    .B(_1155_),
    .C(_1156_),
    .Y(_1158_));
 sg13g2_nor3_2 _2013_ (.A(net966),
    .B(_1157_),
    .C(_1158_),
    .Y(_1159_));
 sg13g2_nor3_2 _2014_ (.A(net975),
    .B(_1128_),
    .C(_1129_),
    .Y(_1160_));
 sg13g2_nor3_2 _2015_ (.A(net977),
    .B(_1130_),
    .C(_1131_),
    .Y(_1161_));
 sg13g2_nor3_2 _2016_ (.A(net965),
    .B(_1159_),
    .C(_1160_),
    .Y(_1162_));
 sg13g2_nor3_2 _2017_ (.A(net963),
    .B(_1161_),
    .C(_1162_),
    .Y(_1163_));
 sg13g2_nor3_2 _2018_ (.A(net979),
    .B(_1132_),
    .C(_1133_),
    .Y(_1164_));
 sg13g2_nor3_2 _2019_ (.A(net982),
    .B(_1134_),
    .C(_1135_),
    .Y(_1165_));
 sg13g2_nor3_2 _2020_ (.A(net962),
    .B(_1163_),
    .C(_1164_),
    .Y(_1166_));
 sg13g2_nor3_2 _2021_ (.A(net960),
    .B(_1165_),
    .C(_1166_),
    .Y(_1167_));
 sg13g2_nor3_2 _2022_ (.A(net984),
    .B(_1136_),
    .C(_1137_),
    .Y(_1168_));
 sg13g2_nor3_2 _2023_ (.A(net987),
    .B(_1138_),
    .C(_1139_),
    .Y(_1169_));
 sg13g2_nor3_2 _2024_ (.A(net958),
    .B(_1167_),
    .C(_1168_),
    .Y(_1170_));
 sg13g2_or2_1 _2025_ (.X(_1171_),
    .B(_1170_),
    .A(_1169_));
 sg13g2_nor3_1 _2026_ (.A(net955),
    .B(_1169_),
    .C(_1170_),
    .Y(_1172_));
 sg13g2_nor3_1 _2027_ (.A(net989),
    .B(_1149_),
    .C(_1150_),
    .Y(_1173_));
 sg13g2_nor2b_1 _2028_ (.A(_0051_),
    .B_N(_1140_),
    .Y(_1174_));
 sg13g2_nor2_1 _2029_ (.A(net979),
    .B(_1174_),
    .Y(_1175_));
 sg13g2_a21oi_1 _2030_ (.A1(_1141_),
    .A2(_1142_),
    .Y(_1176_),
    .B1(net964));
 sg13g2_nor3_2 _2031_ (.A(net981),
    .B(_1175_),
    .C(_1176_),
    .Y(_1177_));
 sg13g2_nor3_2 _2032_ (.A(net962),
    .B(_1143_),
    .C(_1144_),
    .Y(_1178_));
 sg13g2_nor3_2 _2033_ (.A(net959),
    .B(_1145_),
    .C(_1146_),
    .Y(_1179_));
 sg13g2_nor3_2 _2034_ (.A(net984),
    .B(_1177_),
    .C(_1178_),
    .Y(_1180_));
 sg13g2_nor3_2 _2035_ (.A(net987),
    .B(_1179_),
    .C(_1180_),
    .Y(_1181_));
 sg13g2_nor3_2 _2036_ (.A(net958),
    .B(_1147_),
    .C(_1148_),
    .Y(_1182_));
 sg13g2_or2_1 _2037_ (.X(_1183_),
    .B(_1182_),
    .A(_1181_));
 sg13g2_nor3_1 _2038_ (.A(net955),
    .B(_1149_),
    .C(_1150_),
    .Y(_1184_));
 sg13g2_nor3_1 _2039_ (.A(net989),
    .B(_1181_),
    .C(_1182_),
    .Y(_1185_));
 sg13g2_nor3_1 _2040_ (.A(net992),
    .B(_1184_),
    .C(_1185_),
    .Y(_1186_));
 sg13g2_nor3_1 _2041_ (.A(net953),
    .B(_1172_),
    .C(_1173_),
    .Y(_1187_));
 sg13g2_nand2_1 _2042_ (.Y(_1188_),
    .A(_0024_),
    .B(net969));
 sg13g2_o21ai_1 _2043_ (.B1(_1006_),
    .Y(_1189_),
    .A1(_1151_),
    .A2(_1152_));
 sg13g2_a21oi_1 _2044_ (.A1(_1188_),
    .A2(_1189_),
    .Y(_1190_),
    .B1(_1007_));
 sg13g2_nor3_1 _2045_ (.A(net970),
    .B(_1153_),
    .C(_1154_),
    .Y(_1191_));
 sg13g2_nor3_1 _2046_ (.A(net972),
    .B(_1155_),
    .C(_1156_),
    .Y(_1192_));
 sg13g2_nor3_1 _2047_ (.A(net967),
    .B(_1190_),
    .C(_1191_),
    .Y(_1193_));
 sg13g2_nor3_2 _2048_ (.A(net966),
    .B(_1192_),
    .C(_1193_),
    .Y(_1194_));
 sg13g2_nor3_2 _2049_ (.A(net974),
    .B(_1157_),
    .C(_1158_),
    .Y(_1195_));
 sg13g2_nor3_2 _2050_ (.A(net977),
    .B(_1159_),
    .C(_1160_),
    .Y(_1196_));
 sg13g2_nor3_2 _2051_ (.A(net965),
    .B(_1194_),
    .C(_1195_),
    .Y(_1197_));
 sg13g2_nor3_2 _2052_ (.A(net963),
    .B(_1196_),
    .C(_1197_),
    .Y(_1198_));
 sg13g2_nor3_2 _2053_ (.A(net979),
    .B(_1161_),
    .C(_1162_),
    .Y(_1199_));
 sg13g2_nor3_2 _2054_ (.A(net981),
    .B(_1163_),
    .C(_1164_),
    .Y(_1200_));
 sg13g2_nor3_2 _2055_ (.A(net961),
    .B(_1198_),
    .C(_1199_),
    .Y(_1201_));
 sg13g2_nor3_2 _2056_ (.A(net960),
    .B(_1200_),
    .C(_1201_),
    .Y(_1202_));
 sg13g2_nor3_2 _2057_ (.A(net983),
    .B(_1165_),
    .C(_1166_),
    .Y(_1203_));
 sg13g2_nor3_2 _2058_ (.A(net986),
    .B(_1167_),
    .C(_1168_),
    .Y(_1204_));
 sg13g2_nor3_2 _2059_ (.A(_1014_),
    .B(_1202_),
    .C(_1203_),
    .Y(_1205_));
 sg13g2_nor3_1 _2060_ (.A(net955),
    .B(_1204_),
    .C(_1205_),
    .Y(_1206_));
 sg13g2_nor3_1 _2061_ (.A(net988),
    .B(_1169_),
    .C(_1170_),
    .Y(_1207_));
 sg13g2_nor3_1 _2062_ (.A(net992),
    .B(_1172_),
    .C(_1173_),
    .Y(_1208_));
 sg13g2_nor3_1 _2063_ (.A(net953),
    .B(_1206_),
    .C(_1207_),
    .Y(_1209_));
 sg13g2_nor3_1 _2064_ (.A(net952),
    .B(_1208_),
    .C(_1209_),
    .Y(_1210_));
 sg13g2_nor3_1 _2065_ (.A(net996),
    .B(_1186_),
    .C(_1187_),
    .Y(_1211_));
 sg13g2_nand2b_2 _2066_ (.Y(_1212_),
    .B(_1174_),
    .A_N(_0050_));
 sg13g2_nor2_1 _2067_ (.A(net981),
    .B(_1212_),
    .Y(_1213_));
 sg13g2_nor3_1 _2068_ (.A(net961),
    .B(_1175_),
    .C(_1176_),
    .Y(_1214_));
 sg13g2_o21ai_1 _2069_ (.B1(net959),
    .Y(_1215_),
    .A1(_1213_),
    .A2(_1214_));
 sg13g2_o21ai_1 _2070_ (.B1(net983),
    .Y(_1216_),
    .A1(_1177_),
    .A2(_1178_));
 sg13g2_a21oi_2 _2071_ (.B1(net986),
    .Y(_1217_),
    .A2(_1216_),
    .A1(_1215_));
 sg13g2_nor3_2 _2072_ (.A(_1014_),
    .B(_1179_),
    .C(_1180_),
    .Y(_1218_));
 sg13g2_nor3_1 _2073_ (.A(net955),
    .B(_1181_),
    .C(_1182_),
    .Y(_1219_));
 sg13g2_nor3_1 _2074_ (.A(net988),
    .B(_1217_),
    .C(_1218_),
    .Y(_1220_));
 sg13g2_nor3_1 _2075_ (.A(net992),
    .B(_1219_),
    .C(_1220_),
    .Y(_1221_));
 sg13g2_nor3_1 _2076_ (.A(_1016_),
    .B(_1184_),
    .C(_1185_),
    .Y(_1222_));
 sg13g2_nor3_1 _2077_ (.A(net951),
    .B(_1186_),
    .C(_1187_),
    .Y(_1223_));
 sg13g2_nor3_1 _2078_ (.A(net996),
    .B(_1221_),
    .C(_1222_),
    .Y(_1224_));
 sg13g2_nor3_1 _2079_ (.A(net1000),
    .B(_1223_),
    .C(_1224_),
    .Y(_1225_));
 sg13g2_nor3_1 _2080_ (.A(net947),
    .B(_1210_),
    .C(_1211_),
    .Y(_1226_));
 sg13g2_and2_1 _2081_ (.A(_0023_),
    .B(net971),
    .X(_1227_));
 sg13g2_a21oi_1 _2082_ (.A1(_1188_),
    .A2(_1189_),
    .Y(_1228_),
    .B1(net970));
 sg13g2_nor3_1 _2083_ (.A(net972),
    .B(_1190_),
    .C(_1191_),
    .Y(_1229_));
 sg13g2_nor3_1 _2084_ (.A(net967),
    .B(_1227_),
    .C(_1228_),
    .Y(_1230_));
 sg13g2_nor3_1 _2085_ (.A(net966),
    .B(_1229_),
    .C(_1230_),
    .Y(_1231_));
 sg13g2_nor3_1 _2086_ (.A(net974),
    .B(_1192_),
    .C(_1193_),
    .Y(_1232_));
 sg13g2_nor3_2 _2087_ (.A(net977),
    .B(_1194_),
    .C(_1195_),
    .Y(_1233_));
 sg13g2_nor3_2 _2088_ (.A(net965),
    .B(_1231_),
    .C(_1232_),
    .Y(_1234_));
 sg13g2_nor3_2 _2089_ (.A(net963),
    .B(_1233_),
    .C(_1234_),
    .Y(_1235_));
 sg13g2_nor3_2 _2090_ (.A(net979),
    .B(_1196_),
    .C(_1197_),
    .Y(_1236_));
 sg13g2_nor3_2 _2091_ (.A(net981),
    .B(_1198_),
    .C(_1199_),
    .Y(_1237_));
 sg13g2_nor3_2 _2092_ (.A(net961),
    .B(_1235_),
    .C(_1236_),
    .Y(_1238_));
 sg13g2_nor3_2 _2093_ (.A(net959),
    .B(_1237_),
    .C(_1238_),
    .Y(_1239_));
 sg13g2_nor3_2 _2094_ (.A(net983),
    .B(_1200_),
    .C(_1201_),
    .Y(_1240_));
 sg13g2_nor3_2 _2095_ (.A(net986),
    .B(_1202_),
    .C(_1203_),
    .Y(_1241_));
 sg13g2_nor3_2 _2096_ (.A(net958),
    .B(_1239_),
    .C(_1240_),
    .Y(_1242_));
 sg13g2_nor3_1 _2097_ (.A(net955),
    .B(_1241_),
    .C(_1242_),
    .Y(_1243_));
 sg13g2_nor3_1 _2098_ (.A(net988),
    .B(_1204_),
    .C(_1205_),
    .Y(_1244_));
 sg13g2_nor3_1 _2099_ (.A(net992),
    .B(_1206_),
    .C(_1207_),
    .Y(_1245_));
 sg13g2_nor3_1 _2100_ (.A(net953),
    .B(_1243_),
    .C(_1244_),
    .Y(_1246_));
 sg13g2_nor3_1 _2101_ (.A(net951),
    .B(_1245_),
    .C(_1246_),
    .Y(_1247_));
 sg13g2_nor3_1 _2102_ (.A(net996),
    .B(_1208_),
    .C(_1209_),
    .Y(_1248_));
 sg13g2_nor3_1 _2103_ (.A(net1000),
    .B(_1210_),
    .C(_1211_),
    .Y(_1249_));
 sg13g2_nor3_1 _2104_ (.A(net948),
    .B(_1247_),
    .C(_1248_),
    .Y(_1250_));
 sg13g2_nor3_1 _2105_ (.A(net944),
    .B(_1249_),
    .C(_1250_),
    .Y(_1251_));
 sg13g2_nor3_1 _2106_ (.A(net1003),
    .B(_1225_),
    .C(_1226_),
    .Y(_1252_));
 sg13g2_or3_1 _2107_ (.A(net983),
    .B(_0049_),
    .C(_1212_),
    .X(_1253_));
 sg13g2_o21ai_1 _2108_ (.B1(net983),
    .Y(_1254_),
    .A1(_1213_),
    .A2(_1214_));
 sg13g2_a21oi_2 _2109_ (.B1(net986),
    .Y(_1255_),
    .A2(_1254_),
    .A1(_1253_));
 sg13g2_a21oi_2 _2110_ (.B1(net958),
    .Y(_1256_),
    .A2(_1216_),
    .A1(_1215_));
 sg13g2_nor3_1 _2111_ (.A(net955),
    .B(_1217_),
    .C(_1218_),
    .Y(_1257_));
 sg13g2_nor3_1 _2112_ (.A(net988),
    .B(_1255_),
    .C(_1256_),
    .Y(_1258_));
 sg13g2_nor3_1 _2113_ (.A(net992),
    .B(_1257_),
    .C(_1258_),
    .Y(_1259_));
 sg13g2_nor3_1 _2114_ (.A(net953),
    .B(_1219_),
    .C(_1220_),
    .Y(_1260_));
 sg13g2_nor3_1 _2115_ (.A(net951),
    .B(_1221_),
    .C(_1222_),
    .Y(_1261_));
 sg13g2_nor3_1 _2116_ (.A(net996),
    .B(_1259_),
    .C(_1260_),
    .Y(_1262_));
 sg13g2_nor3_1 _2117_ (.A(net1001),
    .B(_1261_),
    .C(_1262_),
    .Y(_1263_));
 sg13g2_nor3_1 _2118_ (.A(net947),
    .B(_1223_),
    .C(_1224_),
    .Y(_1264_));
 sg13g2_nor3_1 _2119_ (.A(net944),
    .B(_1225_),
    .C(_1226_),
    .Y(_1265_));
 sg13g2_nor3_2 _2120_ (.A(net1004),
    .B(_1263_),
    .C(_1264_),
    .Y(_1266_));
 sg13g2_nor3_1 _2121_ (.A(net1009),
    .B(_1265_),
    .C(_1266_),
    .Y(_1267_));
 sg13g2_nor3_1 _2122_ (.A(net939),
    .B(_1251_),
    .C(_1252_),
    .Y(_1268_));
 sg13g2_nand2_1 _2123_ (.Y(_1269_),
    .A(_0022_),
    .B(net973));
 sg13g2_o21ai_1 _2124_ (.B1(net967),
    .Y(_1270_),
    .A1(_1227_),
    .A2(_1228_));
 sg13g2_a21oi_1 _2125_ (.A1(_1269_),
    .A2(_1270_),
    .Y(_1271_),
    .B1(net966));
 sg13g2_nor3_1 _2126_ (.A(net974),
    .B(_1229_),
    .C(_1230_),
    .Y(_1272_));
 sg13g2_nor3_1 _2127_ (.A(net978),
    .B(_1231_),
    .C(_1232_),
    .Y(_1273_));
 sg13g2_nor3_1 _2128_ (.A(net965),
    .B(_1271_),
    .C(_1272_),
    .Y(_1274_));
 sg13g2_nor3_2 _2129_ (.A(net963),
    .B(_1273_),
    .C(_1274_),
    .Y(_1275_));
 sg13g2_nor3_2 _2130_ (.A(net979),
    .B(_1233_),
    .C(_1234_),
    .Y(_1276_));
 sg13g2_nor3_2 _2131_ (.A(net981),
    .B(_1235_),
    .C(_1236_),
    .Y(_1277_));
 sg13g2_nor3_2 _2132_ (.A(net961),
    .B(_1275_),
    .C(_1276_),
    .Y(_1278_));
 sg13g2_nor3_2 _2133_ (.A(net959),
    .B(_1277_),
    .C(_1278_),
    .Y(_1279_));
 sg13g2_nor3_2 _2134_ (.A(net983),
    .B(_1237_),
    .C(_1238_),
    .Y(_1280_));
 sg13g2_nor3_2 _2135_ (.A(net986),
    .B(_1239_),
    .C(_1240_),
    .Y(_1281_));
 sg13g2_nor3_2 _2136_ (.A(net957),
    .B(_1279_),
    .C(_1280_),
    .Y(_1282_));
 sg13g2_nor3_1 _2137_ (.A(net956),
    .B(_1281_),
    .C(_1282_),
    .Y(_1283_));
 sg13g2_nor3_1 _2138_ (.A(net988),
    .B(_1241_),
    .C(_1242_),
    .Y(_1284_));
 sg13g2_nor3_1 _2139_ (.A(net993),
    .B(_1243_),
    .C(_1244_),
    .Y(_1285_));
 sg13g2_nor3_1 _2140_ (.A(net953),
    .B(_1283_),
    .C(_1284_),
    .Y(_1286_));
 sg13g2_nor3_1 _2141_ (.A(net951),
    .B(_1285_),
    .C(_1286_),
    .Y(_1287_));
 sg13g2_nor3_1 _2142_ (.A(net997),
    .B(_1245_),
    .C(_1246_),
    .Y(_1288_));
 sg13g2_nor3_1 _2143_ (.A(net1001),
    .B(_1247_),
    .C(_1248_),
    .Y(_1289_));
 sg13g2_nor3_1 _2144_ (.A(net948),
    .B(_1287_),
    .C(_1288_),
    .Y(_1290_));
 sg13g2_nor3_1 _2145_ (.A(net944),
    .B(_1289_),
    .C(_1290_),
    .Y(_1291_));
 sg13g2_nor3_1 _2146_ (.A(net1003),
    .B(_1249_),
    .C(_1250_),
    .Y(_1292_));
 sg13g2_nor3_1 _2147_ (.A(net1009),
    .B(_1251_),
    .C(_1252_),
    .Y(_1293_));
 sg13g2_nor3_1 _2148_ (.A(net939),
    .B(_1291_),
    .C(_1292_),
    .Y(_1294_));
 sg13g2_nor3_1 _2149_ (.A(net935),
    .B(_1293_),
    .C(_1294_),
    .Y(_1295_));
 sg13g2_nor3_1 _2150_ (.A(net1014),
    .B(_1267_),
    .C(_1268_),
    .Y(_1296_));
 sg13g2_nor3_2 _2151_ (.A(_0049_),
    .B(_0048_),
    .C(_1212_),
    .Y(_1297_));
 sg13g2_and2_1 _2152_ (.A(net958),
    .B(_1297_),
    .X(_1298_));
 sg13g2_a21oi_2 _2153_ (.B1(net958),
    .Y(_1299_),
    .A2(_1254_),
    .A1(_1253_));
 sg13g2_o21ai_1 _2154_ (.B1(net955),
    .Y(_1300_),
    .A1(_1298_),
    .A2(_1299_));
 sg13g2_o21ai_1 _2155_ (.B1(net988),
    .Y(_1301_),
    .A1(_1255_),
    .A2(_1256_));
 sg13g2_a21oi_1 _2156_ (.A1(_1300_),
    .A2(_1301_),
    .Y(_1302_),
    .B1(net992));
 sg13g2_nor3_1 _2157_ (.A(net953),
    .B(_1257_),
    .C(_1258_),
    .Y(_1303_));
 sg13g2_nor3_1 _2158_ (.A(net951),
    .B(_1259_),
    .C(_1260_),
    .Y(_1304_));
 sg13g2_nor3_1 _2159_ (.A(net996),
    .B(_1302_),
    .C(_1303_),
    .Y(_1305_));
 sg13g2_nor3_1 _2160_ (.A(net1000),
    .B(_1304_),
    .C(_1305_),
    .Y(_1306_));
 sg13g2_nor3_1 _2161_ (.A(net947),
    .B(_1261_),
    .C(_1262_),
    .Y(_1307_));
 sg13g2_nor3_1 _2162_ (.A(net945),
    .B(_1263_),
    .C(_1264_),
    .Y(_1308_));
 sg13g2_nor3_1 _2163_ (.A(net1003),
    .B(_1306_),
    .C(_1307_),
    .Y(_1309_));
 sg13g2_nor3_1 _2164_ (.A(net1009),
    .B(_1308_),
    .C(_1309_),
    .Y(_1310_));
 sg13g2_nor3_1 _2165_ (.A(net939),
    .B(_1265_),
    .C(_1266_),
    .Y(_1311_));
 sg13g2_nor3_1 _2166_ (.A(net935),
    .B(_1267_),
    .C(_1268_),
    .Y(_1312_));
 sg13g2_nor3_1 _2167_ (.A(net1015),
    .B(_1310_),
    .C(_1311_),
    .Y(_1313_));
 sg13g2_nor3_1 _2168_ (.A(net1019),
    .B(_1312_),
    .C(_1313_),
    .Y(_1314_));
 sg13g2_nor3_1 _2169_ (.A(net930),
    .B(_1295_),
    .C(_1296_),
    .Y(_1315_));
 sg13g2_and2_1 _2170_ (.A(_0021_),
    .B(net974),
    .X(_1316_));
 sg13g2_a21oi_1 _2171_ (.A1(_1269_),
    .A2(_1270_),
    .Y(_1317_),
    .B1(net974));
 sg13g2_nor3_1 _2172_ (.A(net978),
    .B(_1271_),
    .C(_1272_),
    .Y(_1318_));
 sg13g2_nor3_1 _2173_ (.A(net965),
    .B(_1316_),
    .C(_1317_),
    .Y(_1319_));
 sg13g2_nor3_1 _2174_ (.A(net963),
    .B(_1318_),
    .C(_1319_),
    .Y(_1320_));
 sg13g2_nor3_1 _2175_ (.A(net980),
    .B(_1273_),
    .C(_1274_),
    .Y(_1321_));
 sg13g2_nor3_2 _2176_ (.A(net981),
    .B(_1275_),
    .C(_1276_),
    .Y(_1322_));
 sg13g2_nor3_2 _2177_ (.A(net961),
    .B(_1320_),
    .C(_1321_),
    .Y(_1323_));
 sg13g2_nor3_2 _2178_ (.A(net959),
    .B(_1322_),
    .C(_1323_),
    .Y(_1324_));
 sg13g2_nor3_2 _2179_ (.A(net983),
    .B(_1277_),
    .C(_1278_),
    .Y(_1325_));
 sg13g2_nor3_2 _2180_ (.A(net986),
    .B(_1279_),
    .C(_1280_),
    .Y(_1326_));
 sg13g2_nor3_2 _2181_ (.A(net957),
    .B(_1324_),
    .C(_1325_),
    .Y(_1327_));
 sg13g2_nor3_1 _2182_ (.A(net956),
    .B(_1326_),
    .C(_1327_),
    .Y(_1328_));
 sg13g2_nor3_2 _2183_ (.A(net988),
    .B(_1281_),
    .C(_1282_),
    .Y(_1329_));
 sg13g2_nor3_2 _2184_ (.A(net993),
    .B(_1283_),
    .C(_1284_),
    .Y(_1330_));
 sg13g2_nor3_2 _2185_ (.A(net954),
    .B(_1328_),
    .C(_1329_),
    .Y(_1331_));
 sg13g2_nor3_2 _2186_ (.A(net952),
    .B(_1330_),
    .C(_1331_),
    .Y(_1332_));
 sg13g2_nor3_2 _2187_ (.A(net997),
    .B(_1285_),
    .C(_1286_),
    .Y(_1333_));
 sg13g2_nor3_2 _2188_ (.A(net1001),
    .B(_1287_),
    .C(_1288_),
    .Y(_1334_));
 sg13g2_nor3_2 _2189_ (.A(net948),
    .B(_1332_),
    .C(_1333_),
    .Y(_1335_));
 sg13g2_nor3_2 _2190_ (.A(net945),
    .B(_1334_),
    .C(_1335_),
    .Y(_1336_));
 sg13g2_nor3_1 _2191_ (.A(net1003),
    .B(_1289_),
    .C(_1290_),
    .Y(_1337_));
 sg13g2_nor3_1 _2192_ (.A(net1010),
    .B(_1291_),
    .C(_1292_),
    .Y(_1338_));
 sg13g2_nor3_2 _2193_ (.A(net939),
    .B(_1336_),
    .C(_1337_),
    .Y(_1339_));
 sg13g2_nor3_1 _2194_ (.A(net935),
    .B(_1338_),
    .C(_1339_),
    .Y(_1340_));
 sg13g2_nor3_1 _2195_ (.A(net1014),
    .B(_1293_),
    .C(_1294_),
    .Y(_1341_));
 sg13g2_nor3_1 _2196_ (.A(net1019),
    .B(_1295_),
    .C(_1296_),
    .Y(_1342_));
 sg13g2_nor3_1 _2197_ (.A(net930),
    .B(_1340_),
    .C(_1341_),
    .Y(_1343_));
 sg13g2_nor3_1 _2198_ (.A(net926),
    .B(_1342_),
    .C(_1343_),
    .Y(_1344_));
 sg13g2_nor3_1 _2199_ (.A(net1026),
    .B(_1314_),
    .C(_1315_),
    .Y(_1345_));
 sg13g2_nand2_1 _2200_ (.Y(_1346_),
    .A(_0020_),
    .B(net978));
 sg13g2_o21ai_1 _2201_ (.B1(net965),
    .Y(_1347_),
    .A1(_1316_),
    .A2(_1317_));
 sg13g2_a21oi_1 _2202_ (.A1(_1346_),
    .A2(_1347_),
    .Y(_1348_),
    .B1(net963));
 sg13g2_nor3_1 _2203_ (.A(net980),
    .B(_1318_),
    .C(_1319_),
    .Y(_1349_));
 sg13g2_nor3_1 _2204_ (.A(net982),
    .B(_1320_),
    .C(_1321_),
    .Y(_1350_));
 sg13g2_nor3_2 _2205_ (.A(net961),
    .B(_1348_),
    .C(_1349_),
    .Y(_1351_));
 sg13g2_nor3_2 _2206_ (.A(net959),
    .B(_1350_),
    .C(_1351_),
    .Y(_1352_));
 sg13g2_nor3_1 _2207_ (.A(net985),
    .B(_1322_),
    .C(_1323_),
    .Y(_1353_));
 sg13g2_nor3_2 _2208_ (.A(net986),
    .B(_1324_),
    .C(_1325_),
    .Y(_1354_));
 sg13g2_nor3_2 _2209_ (.A(net957),
    .B(_1352_),
    .C(_1353_),
    .Y(_1355_));
 sg13g2_o21ai_1 _2210_ (.B1(net956),
    .Y(_1356_),
    .A1(_1326_),
    .A2(_1327_));
 sg13g2_o21ai_1 _2211_ (.B1(net990),
    .Y(_1357_),
    .A1(_1354_),
    .A2(_1355_));
 sg13g2_nand3_1 _2212_ (.B(_1356_),
    .C(_1357_),
    .A(net993),
    .Y(_1358_));
 sg13g2_o21ai_1 _2213_ (.B1(net954),
    .Y(_1359_),
    .A1(_1328_),
    .A2(_1329_));
 sg13g2_o21ai_1 _2214_ (.B1(net950),
    .Y(_1360_),
    .A1(_1330_),
    .A2(_1331_));
 sg13g2_nand3_1 _2215_ (.B(_1358_),
    .C(_1359_),
    .A(net995),
    .Y(_1361_));
 sg13g2_nand3_1 _2216_ (.B(_1360_),
    .C(_1361_),
    .A(net1001),
    .Y(_1362_));
 sg13g2_o21ai_1 _2217_ (.B1(net948),
    .Y(_1363_),
    .A1(_1332_),
    .A2(_1333_));
 sg13g2_o21ai_1 _2218_ (.B1(net945),
    .Y(_1364_),
    .A1(_1334_),
    .A2(_1335_));
 sg13g2_nand3_1 _2219_ (.B(_1362_),
    .C(_1363_),
    .A(net1004),
    .Y(_1365_));
 sg13g2_nand3_1 _2220_ (.B(_1364_),
    .C(_1365_),
    .A(net1009),
    .Y(_1366_));
 sg13g2_o21ai_1 _2221_ (.B1(net939),
    .Y(_1367_),
    .A1(_1336_),
    .A2(_1337_));
 sg13g2_o21ai_1 _2222_ (.B1(net935),
    .Y(_1368_),
    .A1(_1338_),
    .A2(_1339_));
 sg13g2_nand3_1 _2223_ (.B(_1366_),
    .C(_1367_),
    .A(net1014),
    .Y(_1369_));
 sg13g2_nand3_1 _2224_ (.B(_1368_),
    .C(_1369_),
    .A(net1019),
    .Y(_1370_));
 sg13g2_o21ai_1 _2225_ (.B1(net930),
    .Y(_1371_),
    .A1(_1340_),
    .A2(_1341_));
 sg13g2_o21ai_1 _2226_ (.B1(net926),
    .Y(_1372_),
    .A1(_1342_),
    .A2(_1343_));
 sg13g2_nand3_1 _2227_ (.B(_1370_),
    .C(_1371_),
    .A(net1026),
    .Y(_1373_));
 sg13g2_nand3_1 _2228_ (.B(_1372_),
    .C(_1373_),
    .A(net1032),
    .Y(_1374_));
 sg13g2_o21ai_1 _2229_ (.B1(net921),
    .Y(_1375_),
    .A1(_1344_),
    .A2(_1345_));
 sg13g2_nand2b_2 _2230_ (.Y(_1376_),
    .B(_1297_),
    .A_N(_0047_));
 sg13g2_nand2b_1 _2231_ (.Y(_1377_),
    .B(_1015_),
    .A_N(_1376_));
 sg13g2_o21ai_1 _2232_ (.B1(net988),
    .Y(_1378_),
    .A1(_1298_),
    .A2(_1299_));
 sg13g2_nor3_1 _2233_ (.A(net951),
    .B(_1302_),
    .C(_1303_),
    .Y(_1379_));
 sg13g2_a21oi_1 _2234_ (.A1(_1377_),
    .A2(_1378_),
    .Y(_1380_),
    .B1(net992));
 sg13g2_a21oi_1 _2235_ (.A1(_1300_),
    .A2(_1301_),
    .Y(_1381_),
    .B1(net953));
 sg13g2_nor3_1 _2236_ (.A(net997),
    .B(_1380_),
    .C(_1381_),
    .Y(_1382_));
 sg13g2_nor3_1 _2237_ (.A(net1000),
    .B(_1379_),
    .C(_1382_),
    .Y(_1383_));
 sg13g2_nor3_1 _2238_ (.A(net947),
    .B(_1304_),
    .C(_1305_),
    .Y(_1384_));
 sg13g2_nor3_1 _2239_ (.A(net946),
    .B(_1306_),
    .C(_1307_),
    .Y(_1385_));
 sg13g2_nor3_1 _2240_ (.A(net1006),
    .B(_1383_),
    .C(_1384_),
    .Y(_1386_));
 sg13g2_nor3_1 _2241_ (.A(net1010),
    .B(_1385_),
    .C(_1386_),
    .Y(_1387_));
 sg13g2_nor3_1 _2242_ (.A(net940),
    .B(_1308_),
    .C(_1309_),
    .Y(_1388_));
 sg13g2_nor3_1 _2243_ (.A(net936),
    .B(_1310_),
    .C(_1311_),
    .Y(_1389_));
 sg13g2_nor3_1 _2244_ (.A(net1015),
    .B(_1387_),
    .C(_1388_),
    .Y(_1390_));
 sg13g2_nor3_1 _2245_ (.A(net1019),
    .B(_1389_),
    .C(_1390_),
    .Y(_1391_));
 sg13g2_nor3_1 _2246_ (.A(net930),
    .B(_1312_),
    .C(_1313_),
    .Y(_1392_));
 sg13g2_nor3_1 _2247_ (.A(net926),
    .B(_1314_),
    .C(_1315_),
    .Y(_1393_));
 sg13g2_nor3_1 _2248_ (.A(net1026),
    .B(_1391_),
    .C(_1392_),
    .Y(_1394_));
 sg13g2_nor3_1 _2249_ (.A(net1032),
    .B(_1393_),
    .C(_1394_),
    .Y(_1395_));
 sg13g2_nor3_1 _2250_ (.A(net921),
    .B(_1344_),
    .C(_1345_),
    .Y(_1396_));
 sg13g2_o21ai_1 _2251_ (.B1(net916),
    .Y(_1397_),
    .A1(_1395_),
    .A2(_1396_));
 sg13g2_nand3_1 _2252_ (.B(_1374_),
    .C(_1375_),
    .A(net1040),
    .Y(_1398_));
 sg13g2_and2_1 _2253_ (.A(_0019_),
    .B(net980),
    .X(_1399_));
 sg13g2_a21oi_1 _2254_ (.A1(_1346_),
    .A2(_1347_),
    .Y(_1400_),
    .B1(net980));
 sg13g2_nor3_1 _2255_ (.A(net982),
    .B(_1348_),
    .C(_1349_),
    .Y(_1401_));
 sg13g2_nor3_1 _2256_ (.A(net961),
    .B(_1399_),
    .C(_1400_),
    .Y(_1402_));
 sg13g2_nor3_1 _2257_ (.A(net959),
    .B(_1401_),
    .C(_1402_),
    .Y(_1403_));
 sg13g2_nor3_1 _2258_ (.A(net985),
    .B(_1350_),
    .C(_1351_),
    .Y(_1404_));
 sg13g2_o21ai_1 _2259_ (.B1(net987),
    .Y(_1405_),
    .A1(_1403_),
    .A2(_1404_));
 sg13g2_o21ai_1 _2260_ (.B1(net957),
    .Y(_1406_),
    .A1(_1352_),
    .A2(_1353_));
 sg13g2_o21ai_1 _2261_ (.B1(net956),
    .Y(_1407_),
    .A1(_1354_),
    .A2(_1355_));
 sg13g2_nand3_1 _2262_ (.B(_1405_),
    .C(_1406_),
    .A(net990),
    .Y(_1408_));
 sg13g2_nand3_1 _2263_ (.B(_1407_),
    .C(_1408_),
    .A(net993),
    .Y(_1409_));
 sg13g2_nand3_1 _2264_ (.B(_1356_),
    .C(_1357_),
    .A(net954),
    .Y(_1410_));
 sg13g2_nand3_1 _2265_ (.B(_1358_),
    .C(_1359_),
    .A(net952),
    .Y(_1411_));
 sg13g2_nand3_1 _2266_ (.B(_1409_),
    .C(_1410_),
    .A(net998),
    .Y(_1412_));
 sg13g2_nand3_1 _2267_ (.B(_1411_),
    .C(_1412_),
    .A(net1001),
    .Y(_1413_));
 sg13g2_nand3_1 _2268_ (.B(_1360_),
    .C(_1361_),
    .A(net948),
    .Y(_1414_));
 sg13g2_nand3_1 _2269_ (.B(_1362_),
    .C(_1363_),
    .A(net945),
    .Y(_1415_));
 sg13g2_nand3_1 _2270_ (.B(_1413_),
    .C(_1414_),
    .A(net1004),
    .Y(_1416_));
 sg13g2_nand3_1 _2271_ (.B(_1415_),
    .C(_1416_),
    .A(net1009),
    .Y(_1417_));
 sg13g2_nand3_1 _2272_ (.B(_1364_),
    .C(_1365_),
    .A(net941),
    .Y(_1418_));
 sg13g2_nand3_1 _2273_ (.B(_1366_),
    .C(_1367_),
    .A(net935),
    .Y(_1419_));
 sg13g2_nand3_1 _2274_ (.B(_1417_),
    .C(_1418_),
    .A(net1014),
    .Y(_1420_));
 sg13g2_nand3_1 _2275_ (.B(_1419_),
    .C(_1420_),
    .A(net1019),
    .Y(_1421_));
 sg13g2_nand3_1 _2276_ (.B(_1368_),
    .C(_1369_),
    .A(net930),
    .Y(_1422_));
 sg13g2_nand3_1 _2277_ (.B(_1370_),
    .C(_1371_),
    .A(net926),
    .Y(_1423_));
 sg13g2_nand3_1 _2278_ (.B(_1421_),
    .C(_1422_),
    .A(net1026),
    .Y(_1424_));
 sg13g2_nand3_1 _2279_ (.B(_1423_),
    .C(_1424_),
    .A(net1032),
    .Y(_1425_));
 sg13g2_nand3_1 _2280_ (.B(_1372_),
    .C(_1373_),
    .A(net921),
    .Y(_1426_));
 sg13g2_nand3_1 _2281_ (.B(_1374_),
    .C(_1375_),
    .A(net916),
    .Y(_1427_));
 sg13g2_nand3_1 _2282_ (.B(_1425_),
    .C(_1426_),
    .A(net1040),
    .Y(_1428_));
 sg13g2_nand3_1 _2283_ (.B(_1427_),
    .C(_1428_),
    .A(net1047),
    .Y(_1429_));
 sg13g2_nand3_1 _2284_ (.B(_1397_),
    .C(_1398_),
    .A(net910),
    .Y(_1430_));
 sg13g2_o21ai_1 _2285_ (.B1(net953),
    .Y(_1431_),
    .A1(_0046_),
    .A2(_1376_));
 sg13g2_nand3_1 _2286_ (.B(_1377_),
    .C(_1378_),
    .A(net992),
    .Y(_1432_));
 sg13g2_nor3_1 _2287_ (.A(net951),
    .B(_1380_),
    .C(_1381_),
    .Y(_1433_));
 sg13g2_a21oi_1 _2288_ (.A1(_1431_),
    .A2(_1432_),
    .Y(_1434_),
    .B1(net996));
 sg13g2_nor3_1 _2289_ (.A(net1000),
    .B(_1433_),
    .C(_1434_),
    .Y(_1435_));
 sg13g2_nor3_1 _2290_ (.A(net947),
    .B(_1379_),
    .C(_1382_),
    .Y(_1436_));
 sg13g2_nor3_1 _2291_ (.A(net944),
    .B(_1383_),
    .C(_1384_),
    .Y(_1437_));
 sg13g2_nor3_1 _2292_ (.A(net1006),
    .B(_1435_),
    .C(_1436_),
    .Y(_1438_));
 sg13g2_nor3_1 _2293_ (.A(net1010),
    .B(_1437_),
    .C(_1438_),
    .Y(_1439_));
 sg13g2_nor3_1 _2294_ (.A(net940),
    .B(_1385_),
    .C(_1386_),
    .Y(_1440_));
 sg13g2_nor3_1 _2295_ (.A(net936),
    .B(_1387_),
    .C(_1388_),
    .Y(_1441_));
 sg13g2_nor3_1 _2296_ (.A(net1015),
    .B(_1439_),
    .C(_1440_),
    .Y(_1442_));
 sg13g2_nor3_1 _2297_ (.A(net1020),
    .B(_1441_),
    .C(_1442_),
    .Y(_1443_));
 sg13g2_nor3_1 _2298_ (.A(net931),
    .B(_1389_),
    .C(_1390_),
    .Y(_1444_));
 sg13g2_nor3_1 _2299_ (.A(net926),
    .B(_1391_),
    .C(_1392_),
    .Y(_1445_));
 sg13g2_nor3_1 _2300_ (.A(net1027),
    .B(_1443_),
    .C(_1444_),
    .Y(_1446_));
 sg13g2_nor3_1 _2301_ (.A(net1032),
    .B(_1445_),
    .C(_1446_),
    .Y(_1447_));
 sg13g2_nor3_1 _2302_ (.A(net921),
    .B(_1393_),
    .C(_1394_),
    .Y(_1448_));
 sg13g2_nor3_1 _2303_ (.A(net916),
    .B(_1395_),
    .C(_1396_),
    .Y(_1449_));
 sg13g2_nor3_1 _2304_ (.A(net1040),
    .B(_1447_),
    .C(_1448_),
    .Y(_1450_));
 sg13g2_nand3_1 _2305_ (.B(_1397_),
    .C(_1398_),
    .A(net1047),
    .Y(_1451_));
 sg13g2_o21ai_1 _2306_ (.B1(net910),
    .Y(_1452_),
    .A1(_1449_),
    .A2(_1450_));
 sg13g2_nand3_1 _2307_ (.B(_1451_),
    .C(_1452_),
    .A(net905),
    .Y(_1453_));
 sg13g2_nand3_1 _2308_ (.B(_1429_),
    .C(_1430_),
    .A(net1055),
    .Y(_1454_));
 sg13g2_nand2_1 _2309_ (.Y(_1455_),
    .A(_0018_),
    .B(net982));
 sg13g2_o21ai_1 _2310_ (.B1(net961),
    .Y(_1456_),
    .A1(_1399_),
    .A2(_1400_));
 sg13g2_a21oi_1 _2311_ (.A1(_1455_),
    .A2(_1456_),
    .Y(_1457_),
    .B1(net959));
 sg13g2_nor3_1 _2312_ (.A(net985),
    .B(_1401_),
    .C(_1402_),
    .Y(_1458_));
 sg13g2_o21ai_1 _2313_ (.B1(net987),
    .Y(_1459_),
    .A1(_1457_),
    .A2(_1458_));
 sg13g2_o21ai_1 _2314_ (.B1(net957),
    .Y(_1460_),
    .A1(_1403_),
    .A2(_1404_));
 sg13g2_nand3_1 _2315_ (.B(_1405_),
    .C(_1406_),
    .A(net956),
    .Y(_1461_));
 sg13g2_nand3_1 _2316_ (.B(_1459_),
    .C(_1460_),
    .A(net990),
    .Y(_1462_));
 sg13g2_nand3_1 _2317_ (.B(_1461_),
    .C(_1462_),
    .A(net993),
    .Y(_1463_));
 sg13g2_nand3_1 _2318_ (.B(_1407_),
    .C(_1408_),
    .A(net954),
    .Y(_1464_));
 sg13g2_nand3_1 _2319_ (.B(_1409_),
    .C(_1410_),
    .A(net950),
    .Y(_1465_));
 sg13g2_nand3_1 _2320_ (.B(_1463_),
    .C(_1464_),
    .A(net995),
    .Y(_1466_));
 sg13g2_nand3_1 _2321_ (.B(_1465_),
    .C(_1466_),
    .A(net1001),
    .Y(_1467_));
 sg13g2_nand3_1 _2322_ (.B(_1411_),
    .C(_1412_),
    .A(net949),
    .Y(_1468_));
 sg13g2_nand3_1 _2323_ (.B(_1413_),
    .C(_1414_),
    .A(net945),
    .Y(_1469_));
 sg13g2_nand3_1 _2324_ (.B(_1467_),
    .C(_1468_),
    .A(net1004),
    .Y(_1470_));
 sg13g2_nand3_1 _2325_ (.B(_1469_),
    .C(_1470_),
    .A(net1011),
    .Y(_1471_));
 sg13g2_nand3_1 _2326_ (.B(_1415_),
    .C(_1416_),
    .A(net941),
    .Y(_1472_));
 sg13g2_nand3_1 _2327_ (.B(_1417_),
    .C(_1418_),
    .A(net935),
    .Y(_1473_));
 sg13g2_nand3_1 _2328_ (.B(_1471_),
    .C(_1472_),
    .A(net1014),
    .Y(_1474_));
 sg13g2_nand3_1 _2329_ (.B(_1473_),
    .C(_1474_),
    .A(net1019),
    .Y(_1475_));
 sg13g2_nand3_1 _2330_ (.B(_1419_),
    .C(_1420_),
    .A(net931),
    .Y(_1476_));
 sg13g2_nand3_1 _2331_ (.B(_1421_),
    .C(_1422_),
    .A(net927),
    .Y(_1477_));
 sg13g2_nand3_1 _2332_ (.B(_1475_),
    .C(_1476_),
    .A(net1026),
    .Y(_1478_));
 sg13g2_nand3_1 _2333_ (.B(_1477_),
    .C(_1478_),
    .A(net1032),
    .Y(_1479_));
 sg13g2_nand3_1 _2334_ (.B(_1423_),
    .C(_1424_),
    .A(net921),
    .Y(_1480_));
 sg13g2_nand3_1 _2335_ (.B(_1425_),
    .C(_1426_),
    .A(net916),
    .Y(_1481_));
 sg13g2_nand3_1 _2336_ (.B(_1479_),
    .C(_1480_),
    .A(net1040),
    .Y(_1482_));
 sg13g2_nand3_1 _2337_ (.B(_1481_),
    .C(_1482_),
    .A(net1047),
    .Y(_1483_));
 sg13g2_nand3_1 _2338_ (.B(_1427_),
    .C(_1428_),
    .A(net910),
    .Y(_1484_));
 sg13g2_nand3_1 _2339_ (.B(_1429_),
    .C(_1430_),
    .A(net905),
    .Y(_1485_));
 sg13g2_nand3_1 _2340_ (.B(_1483_),
    .C(_1484_),
    .A(net1055),
    .Y(_1486_));
 sg13g2_nand3_1 _2341_ (.B(_1485_),
    .C(_1486_),
    .A(net1063),
    .Y(_1487_));
 sg13g2_nand3_1 _2342_ (.B(_1453_),
    .C(_1454_),
    .A(net899),
    .Y(_1488_));
 sg13g2_and2_1 _2343_ (.A(_0017_),
    .B(net985),
    .X(_1489_));
 sg13g2_a21oi_1 _2344_ (.A1(_1455_),
    .A2(_1456_),
    .Y(_1490_),
    .B1(net985));
 sg13g2_o21ai_1 _2345_ (.B1(net987),
    .Y(_1491_),
    .A1(_1489_),
    .A2(_1490_));
 sg13g2_o21ai_1 _2346_ (.B1(net957),
    .Y(_1492_),
    .A1(_1457_),
    .A2(_1458_));
 sg13g2_nand3_1 _2347_ (.B(_1459_),
    .C(_1460_),
    .A(net956),
    .Y(_1493_));
 sg13g2_nand3_1 _2348_ (.B(_1491_),
    .C(_1492_),
    .A(net990),
    .Y(_1494_));
 sg13g2_nand3_1 _2349_ (.B(_1493_),
    .C(_1494_),
    .A(net994),
    .Y(_1495_));
 sg13g2_nand3_1 _2350_ (.B(_1461_),
    .C(_1462_),
    .A(net954),
    .Y(_1496_));
 sg13g2_nand3_1 _2351_ (.B(_1463_),
    .C(_1464_),
    .A(net950),
    .Y(_1497_));
 sg13g2_nand3_1 _2352_ (.B(_1495_),
    .C(_1496_),
    .A(net995),
    .Y(_1498_));
 sg13g2_nand3_1 _2353_ (.B(_1497_),
    .C(_1498_),
    .A(net999),
    .Y(_1499_));
 sg13g2_nand3_1 _2354_ (.B(_1465_),
    .C(_1466_),
    .A(net949),
    .Y(_1500_));
 sg13g2_nand3_1 _2355_ (.B(_1467_),
    .C(_1468_),
    .A(net946),
    .Y(_1501_));
 sg13g2_nand3_1 _2356_ (.B(_1499_),
    .C(_1500_),
    .A(net1005),
    .Y(_1502_));
 sg13g2_nand3_1 _2357_ (.B(_1501_),
    .C(_1502_),
    .A(net1011),
    .Y(_1503_));
 sg13g2_nand3_1 _2358_ (.B(_1469_),
    .C(_1470_),
    .A(net941),
    .Y(_1504_));
 sg13g2_nand3_1 _2359_ (.B(_1471_),
    .C(_1472_),
    .A(net935),
    .Y(_1505_));
 sg13g2_nand3_1 _2360_ (.B(_1503_),
    .C(_1504_),
    .A(net1016),
    .Y(_1506_));
 sg13g2_nand3_1 _2361_ (.B(_1505_),
    .C(_1506_),
    .A(net1019),
    .Y(_1507_));
 sg13g2_nand3_1 _2362_ (.B(_1473_),
    .C(_1474_),
    .A(net930),
    .Y(_1508_));
 sg13g2_nand3_1 _2363_ (.B(_1475_),
    .C(_1476_),
    .A(net926),
    .Y(_1509_));
 sg13g2_nand3_1 _2364_ (.B(_1507_),
    .C(_1508_),
    .A(net1026),
    .Y(_1510_));
 sg13g2_nand3_1 _2365_ (.B(_1509_),
    .C(_1510_),
    .A(net1032),
    .Y(_1511_));
 sg13g2_nand3_1 _2366_ (.B(_1477_),
    .C(_1478_),
    .A(net921),
    .Y(_1512_));
 sg13g2_nand3_1 _2367_ (.B(_1479_),
    .C(_1480_),
    .A(net917),
    .Y(_1513_));
 sg13g2_nand3_1 _2368_ (.B(_1511_),
    .C(_1512_),
    .A(net1040),
    .Y(_1514_));
 sg13g2_nand3_1 _2369_ (.B(_1513_),
    .C(_1514_),
    .A(net1047),
    .Y(_1515_));
 sg13g2_nand3_1 _2370_ (.B(_1481_),
    .C(_1482_),
    .A(net910),
    .Y(_1516_));
 sg13g2_nand3_1 _2371_ (.B(_1483_),
    .C(_1484_),
    .A(net905),
    .Y(_1517_));
 sg13g2_nand3_1 _2372_ (.B(_1515_),
    .C(_1516_),
    .A(net1055),
    .Y(_1518_));
 sg13g2_nand3_1 _2373_ (.B(_1517_),
    .C(_1518_),
    .A(net1063),
    .Y(_1519_));
 sg13g2_nand3_1 _2374_ (.B(_1485_),
    .C(_1486_),
    .A(net899),
    .Y(_1520_));
 sg13g2_a21oi_1 _2375_ (.A1(_1519_),
    .A2(_1520_),
    .Y(_1521_),
    .B1(net893));
 sg13g2_a21oi_1 _2376_ (.A1(_1487_),
    .A2(_1488_),
    .Y(_1522_),
    .B1(net1071));
 sg13g2_o21ai_1 _2377_ (.B1(net886),
    .Y(_1523_),
    .A1(_1521_),
    .A2(_1522_));
 sg13g2_nor2b_2 _2378_ (.A(net3),
    .B_N(net4),
    .Y(_1524_));
 sg13g2_and3_1 _2379_ (.X(_1525_),
    .A(net1098),
    .B(net2),
    .C(_1524_));
 sg13g2_nand3_1 _2380_ (.B(net2),
    .C(_1524_),
    .A(net1099),
    .Y(_1526_));
 sg13g2_nand2_1 _2381_ (.Y(_1527_),
    .A(_0016_),
    .B(net987));
 sg13g2_o21ai_1 _2382_ (.B1(net957),
    .Y(_1528_),
    .A1(_1489_),
    .A2(_1490_));
 sg13g2_nand3_1 _2383_ (.B(_1491_),
    .C(_1492_),
    .A(net956),
    .Y(_1529_));
 sg13g2_nand3_1 _2384_ (.B(_1527_),
    .C(_1528_),
    .A(net990),
    .Y(_1530_));
 sg13g2_nand3_1 _2385_ (.B(_1529_),
    .C(_1530_),
    .A(net994),
    .Y(_1531_));
 sg13g2_nand3_1 _2386_ (.B(_1493_),
    .C(_1494_),
    .A(net954),
    .Y(_1532_));
 sg13g2_nand3_1 _2387_ (.B(_1495_),
    .C(_1496_),
    .A(net950),
    .Y(_1533_));
 sg13g2_nand3_1 _2388_ (.B(_1531_),
    .C(_1532_),
    .A(net995),
    .Y(_1534_));
 sg13g2_nand3_1 _2389_ (.B(_1533_),
    .C(_1534_),
    .A(net999),
    .Y(_1535_));
 sg13g2_nand3_1 _2390_ (.B(_1497_),
    .C(_1498_),
    .A(net949),
    .Y(_1536_));
 sg13g2_nand3_1 _2391_ (.B(_1499_),
    .C(_1500_),
    .A(net943),
    .Y(_1537_));
 sg13g2_nand3_1 _2392_ (.B(_1535_),
    .C(_1536_),
    .A(net1005),
    .Y(_1538_));
 sg13g2_nand3_1 _2393_ (.B(_1537_),
    .C(_1538_),
    .A(net1011),
    .Y(_1539_));
 sg13g2_nand3_1 _2394_ (.B(_1501_),
    .C(_1502_),
    .A(net942),
    .Y(_1540_));
 sg13g2_nand3_1 _2395_ (.B(_1503_),
    .C(_1504_),
    .A(net937),
    .Y(_1541_));
 sg13g2_nand3_1 _2396_ (.B(_1539_),
    .C(_1540_),
    .A(net1016),
    .Y(_1542_));
 sg13g2_nand3_1 _2397_ (.B(_1541_),
    .C(_1542_),
    .A(net1021),
    .Y(_1543_));
 sg13g2_nand3_1 _2398_ (.B(_1505_),
    .C(_1506_),
    .A(net930),
    .Y(_1544_));
 sg13g2_nand3_1 _2399_ (.B(_1507_),
    .C(_1508_),
    .A(net926),
    .Y(_1545_));
 sg13g2_nand3_1 _2400_ (.B(_1543_),
    .C(_1544_),
    .A(net1028),
    .Y(_1546_));
 sg13g2_nand3_1 _2401_ (.B(_1545_),
    .C(_1546_),
    .A(net1034),
    .Y(_1547_));
 sg13g2_nand3_1 _2402_ (.B(_1509_),
    .C(_1510_),
    .A(net921),
    .Y(_1548_));
 sg13g2_nand3_1 _2403_ (.B(_1511_),
    .C(_1512_),
    .A(net916),
    .Y(_1549_));
 sg13g2_nand3_1 _2404_ (.B(_1547_),
    .C(_1548_),
    .A(net1040),
    .Y(_1550_));
 sg13g2_nand3_1 _2405_ (.B(_1549_),
    .C(_1550_),
    .A(net1047),
    .Y(_1551_));
 sg13g2_nand3_1 _2406_ (.B(_1513_),
    .C(_1514_),
    .A(net910),
    .Y(_1552_));
 sg13g2_nand3_1 _2407_ (.B(_1515_),
    .C(_1516_),
    .A(net905),
    .Y(_1553_));
 sg13g2_nand3_1 _2408_ (.B(_1551_),
    .C(_1552_),
    .A(net1055),
    .Y(_1554_));
 sg13g2_nand3_1 _2409_ (.B(_1553_),
    .C(_1554_),
    .A(net1063),
    .Y(_1555_));
 sg13g2_nand3_1 _2410_ (.B(_1517_),
    .C(_1518_),
    .A(net899),
    .Y(_1556_));
 sg13g2_a21oi_1 _2411_ (.A1(_1555_),
    .A2(_1556_),
    .Y(_1557_),
    .B1(net893));
 sg13g2_a21oi_1 _2412_ (.A1(_1519_),
    .A2(_1520_),
    .Y(_1558_),
    .B1(net1070));
 sg13g2_o21ai_1 _2413_ (.B1(net1078),
    .Y(_1559_),
    .A1(_1557_),
    .A2(_1558_));
 sg13g2_nand3_1 _2414_ (.B(net879),
    .C(_1559_),
    .A(_1523_),
    .Y(_1560_));
 sg13g2_nor2b_2 _2415_ (.A(net2),
    .B_N(net1099),
    .Y(_1561_));
 sg13g2_and2_1 _2416_ (.A(_1524_),
    .B(_1561_),
    .X(_1562_));
 sg13g2_nand2_1 _2417_ (.Y(_1563_),
    .A(_1524_),
    .B(_1561_));
 sg13g2_nand3_1 _2418_ (.B(_1528_),
    .C(net875),
    .A(_1527_),
    .Y(_1564_));
 sg13g2_nor2_2 _2419_ (.A(net1099),
    .B(net2),
    .Y(_1565_));
 sg13g2_and2_1 _2420_ (.A(_1524_),
    .B(_1565_),
    .X(_1566_));
 sg13g2_nor2b_2 _2421_ (.A(net1099),
    .B_N(net2),
    .Y(_1567_));
 sg13g2_and2_1 _2422_ (.A(_1524_),
    .B(_1567_),
    .X(_1568_));
 sg13g2_nand3_1 _2423_ (.B(\a[16] ),
    .C(\a[17] ),
    .A(net1101),
    .Y(_1569_));
 sg13g2_nor2b_1 _2424_ (.A(net4),
    .B_N(net3),
    .Y(_1570_));
 sg13g2_nand2b_1 _2425_ (.Y(_1571_),
    .B(net3),
    .A_N(net4));
 sg13g2_o21ai_1 _2426_ (.B1(_1569_),
    .Y(_1572_),
    .A1(net1085),
    .A2(\a[17] ));
 sg13g2_nor2_1 _2427_ (.A(net1090),
    .B(_1572_),
    .Y(_1573_));
 sg13g2_a221oi_1 _2428_ (.B2(net969),
    .C1(_1573_),
    .B1(net864),
    .A1(net1022),
    .Y(_1574_),
    .A2(net870));
 sg13g2_nor2_1 _2429_ (.A(net3),
    .B(net4),
    .Y(_1575_));
 sg13g2_or2_2 _2430_ (.X(_1576_),
    .B(net4),
    .A(net3));
 sg13g2_and2_1 _2431_ (.A(_1565_),
    .B(net1086),
    .X(_1577_));
 sg13g2_nand2_1 _2432_ (.Y(_1578_),
    .A(_1565_),
    .B(net1086));
 sg13g2_and2_1 _2433_ (.A(net1100),
    .B(net1086),
    .X(_1579_));
 sg13g2_and2_1 _2434_ (.A(\a[17] ),
    .B(net856),
    .X(_1580_));
 sg13g2_o21ai_1 _2435_ (.B1(\a[16] ),
    .Y(_1581_),
    .A1(net860),
    .A2(_1580_));
 sg13g2_and2_1 _2436_ (.A(_1567_),
    .B(net1086),
    .X(_1582_));
 sg13g2_nand2_2 _2437_ (.Y(_1583_),
    .A(_1567_),
    .B(net1086));
 sg13g2_a21oi_1 _2438_ (.A1(\ayayayayayaya.b[16] ),
    .A2(net853),
    .Y(_1584_),
    .B1(net1105));
 sg13g2_and4_1 _2439_ (.A(_1564_),
    .B(_1574_),
    .C(_1581_),
    .D(_1584_),
    .X(_1585_));
 sg13g2_o21ai_1 _2440_ (.B1(net874),
    .Y(_1586_),
    .A1(_1204_),
    .A2(_1205_));
 sg13g2_a21oi_1 _2441_ (.A1(\ayayayayayaya.b[28] ),
    .A2(net865),
    .Y(_1587_),
    .B1(net1095));
 sg13g2_a22oi_1 _2442_ (.Y(_1588_),
    .B1(net852),
    .B2(net969),
    .A2(net870),
    .A1(net1002));
 sg13g2_and2_1 _2443_ (.A(\a[24] ),
    .B(net856),
    .X(_1589_));
 sg13g2_a21oi_1 _2444_ (.A1(net1102),
    .A2(\a[24] ),
    .Y(_1590_),
    .B1(net1091));
 sg13g2_or2_1 _2445_ (.X(_1591_),
    .B(_1590_),
    .A(_1589_));
 sg13g2_o21ai_1 _2446_ (.B1(net857),
    .Y(_1592_),
    .A1(\a[25] ),
    .A2(net1091));
 sg13g2_a22oi_1 _2447_ (.Y(_1593_),
    .B1(_1592_),
    .B2(\a[24] ),
    .A2(_1591_),
    .A1(\a[25] ));
 sg13g2_and4_1 _2448_ (.A(_1586_),
    .B(_1587_),
    .C(_1588_),
    .D(_1593_),
    .X(_1594_));
 sg13g2_nor3_2 _2449_ (.A(_0046_),
    .B(_0045_),
    .C(_1376_),
    .Y(_1595_));
 sg13g2_nand2b_2 _2450_ (.Y(_1596_),
    .B(_1595_),
    .A_N(_0044_));
 sg13g2_nor2_1 _2451_ (.A(_0043_),
    .B(_1596_),
    .Y(_1597_));
 sg13g2_nor4_2 _2452_ (.A(net1009),
    .B(_0043_),
    .C(_0042_),
    .Y(_1598_),
    .D(_1596_));
 sg13g2_nor2_1 _2453_ (.A(net996),
    .B(_1595_),
    .Y(_1599_));
 sg13g2_a21oi_1 _2454_ (.A1(_1431_),
    .A2(_1432_),
    .Y(_1600_),
    .B1(net951));
 sg13g2_nand2_1 _2455_ (.Y(_1601_),
    .A(net947),
    .B(_1596_));
 sg13g2_o21ai_1 _2456_ (.B1(net1000),
    .Y(_1602_),
    .A1(_1599_),
    .A2(_1600_));
 sg13g2_nor2_1 _2457_ (.A(net1003),
    .B(_1597_),
    .Y(_1603_));
 sg13g2_a21oi_2 _2458_ (.B1(net944),
    .Y(_1604_),
    .A2(_1602_),
    .A1(_1601_));
 sg13g2_nor3_2 _2459_ (.A(net939),
    .B(_1603_),
    .C(_1604_),
    .Y(_1605_));
 sg13g2_nor3_1 _2460_ (.A(net1000),
    .B(_1599_),
    .C(_1600_),
    .Y(_1606_));
 sg13g2_nor3_1 _2461_ (.A(net947),
    .B(_1433_),
    .C(_1434_),
    .Y(_1607_));
 sg13g2_nor3_1 _2462_ (.A(net944),
    .B(_1606_),
    .C(_1607_),
    .Y(_1608_));
 sg13g2_a21oi_1 _2463_ (.A1(_1601_),
    .A2(_1602_),
    .Y(_1609_),
    .B1(net1003));
 sg13g2_nor3_2 _2464_ (.A(net1010),
    .B(_1603_),
    .C(_1604_),
    .Y(_1610_));
 sg13g2_nor3_2 _2465_ (.A(net939),
    .B(_1608_),
    .C(_1609_),
    .Y(_1611_));
 sg13g2_nor3_2 _2466_ (.A(net935),
    .B(_1610_),
    .C(_1611_),
    .Y(_1612_));
 sg13g2_nor3_2 _2467_ (.A(net1014),
    .B(_1598_),
    .C(_1605_),
    .Y(_1613_));
 sg13g2_or4_2 _2468_ (.A(_0043_),
    .B(_0042_),
    .C(_0041_),
    .D(_1596_),
    .X(_1614_));
 sg13g2_nand2b_1 _2469_ (.Y(_1615_),
    .B(net937),
    .A_N(_1614_));
 sg13g2_o21ai_1 _2470_ (.B1(net1014),
    .Y(_1616_),
    .A1(_1598_),
    .A2(_1605_));
 sg13g2_a21oi_1 _2471_ (.A1(_1615_),
    .A2(_1616_),
    .Y(_1617_),
    .B1(net1021));
 sg13g2_nor3_2 _2472_ (.A(net930),
    .B(_1612_),
    .C(_1613_),
    .Y(_1618_));
 sg13g2_nor3_1 _2473_ (.A(net944),
    .B(_1435_),
    .C(_1436_),
    .Y(_1619_));
 sg13g2_nor3_1 _2474_ (.A(net1003),
    .B(_1606_),
    .C(_1607_),
    .Y(_1620_));
 sg13g2_nor3_1 _2475_ (.A(net1010),
    .B(_1608_),
    .C(_1609_),
    .Y(_1621_));
 sg13g2_nor3_1 _2476_ (.A(net940),
    .B(_1619_),
    .C(_1620_),
    .Y(_1622_));
 sg13g2_nor3_2 _2477_ (.A(net1019),
    .B(_1612_),
    .C(_1613_),
    .Y(_1623_));
 sg13g2_nor3_2 _2478_ (.A(net936),
    .B(_1621_),
    .C(_1622_),
    .Y(_1624_));
 sg13g2_nor3_2 _2479_ (.A(net1014),
    .B(_1610_),
    .C(_1611_),
    .Y(_1625_));
 sg13g2_nor3_2 _2480_ (.A(net931),
    .B(_1624_),
    .C(_1625_),
    .Y(_1626_));
 sg13g2_nor3_2 _2481_ (.A(net927),
    .B(_1623_),
    .C(_1626_),
    .Y(_1627_));
 sg13g2_nor3_2 _2482_ (.A(net1026),
    .B(_1617_),
    .C(_1618_),
    .Y(_1628_));
 sg13g2_nor3_1 _2483_ (.A(net1021),
    .B(_0040_),
    .C(_1614_),
    .Y(_1629_));
 sg13g2_a21oi_1 _2484_ (.A1(_1615_),
    .A2(_1616_),
    .Y(_1630_),
    .B1(net932));
 sg13g2_nor3_2 _2485_ (.A(net926),
    .B(_1617_),
    .C(_1618_),
    .Y(_1631_));
 sg13g2_nor3_1 _2486_ (.A(net1028),
    .B(_1629_),
    .C(_1630_),
    .Y(_1632_));
 sg13g2_nor3_1 _2487_ (.A(net1032),
    .B(_1631_),
    .C(_1632_),
    .Y(_1633_));
 sg13g2_nor3_2 _2488_ (.A(net921),
    .B(_1627_),
    .C(_1628_),
    .Y(_1634_));
 sg13g2_nor3_1 _2489_ (.A(net1010),
    .B(_1619_),
    .C(_1620_),
    .Y(_1635_));
 sg13g2_nor3_1 _2490_ (.A(net940),
    .B(_1437_),
    .C(_1438_),
    .Y(_1636_));
 sg13g2_nor3_1 _2491_ (.A(net936),
    .B(_1635_),
    .C(_1636_),
    .Y(_1637_));
 sg13g2_nor3_1 _2492_ (.A(net1015),
    .B(_1621_),
    .C(_1622_),
    .Y(_1638_));
 sg13g2_nor3_1 _2493_ (.A(net1020),
    .B(_1624_),
    .C(_1625_),
    .Y(_1639_));
 sg13g2_nor3_1 _2494_ (.A(net931),
    .B(_1637_),
    .C(_1638_),
    .Y(_1640_));
 sg13g2_nor3_2 _2495_ (.A(net1032),
    .B(_1627_),
    .C(_1628_),
    .Y(_1641_));
 sg13g2_nor3_1 _2496_ (.A(net927),
    .B(_1639_),
    .C(_1640_),
    .Y(_1642_));
 sg13g2_nor3_2 _2497_ (.A(net1026),
    .B(_1623_),
    .C(_1626_),
    .Y(_1643_));
 sg13g2_nor3_1 _2498_ (.A(net922),
    .B(_1642_),
    .C(_1643_),
    .Y(_1644_));
 sg13g2_nor3_1 _2499_ (.A(net917),
    .B(_1641_),
    .C(_1644_),
    .Y(_1645_));
 sg13g2_nor3_1 _2500_ (.A(net1040),
    .B(_1633_),
    .C(_1634_),
    .Y(_1646_));
 sg13g2_nor3_2 _2501_ (.A(_0040_),
    .B(_0039_),
    .C(_1614_),
    .Y(_1647_));
 sg13g2_nor2_1 _2502_ (.A(net1023),
    .B(_1647_),
    .Y(_1648_));
 sg13g2_nor3_2 _2503_ (.A(net928),
    .B(_1629_),
    .C(_1630_),
    .Y(_1649_));
 sg13g2_nor3_2 _2504_ (.A(net1031),
    .B(_1648_),
    .C(_1649_),
    .Y(_1650_));
 sg13g2_nor3_2 _2505_ (.A(net923),
    .B(_1631_),
    .C(_1632_),
    .Y(_1651_));
 sg13g2_nor3_2 _2506_ (.A(net916),
    .B(_1633_),
    .C(_1634_),
    .Y(_1652_));
 sg13g2_nor3_1 _2507_ (.A(net1038),
    .B(_1650_),
    .C(_1651_),
    .Y(_1653_));
 sg13g2_nor3_1 _2508_ (.A(net1049),
    .B(_1652_),
    .C(_1653_),
    .Y(_1654_));
 sg13g2_nor3_1 _2509_ (.A(net910),
    .B(_1645_),
    .C(_1646_),
    .Y(_1655_));
 sg13g2_nor3_1 _2510_ (.A(net936),
    .B(_1439_),
    .C(_1440_),
    .Y(_1656_));
 sg13g2_nor3_1 _2511_ (.A(net1015),
    .B(_1635_),
    .C(_1636_),
    .Y(_1657_));
 sg13g2_nor3_1 _2512_ (.A(net1020),
    .B(_1637_),
    .C(_1638_),
    .Y(_1658_));
 sg13g2_nor3_1 _2513_ (.A(net931),
    .B(_1656_),
    .C(_1657_),
    .Y(_1659_));
 sg13g2_nor3_1 _2514_ (.A(net927),
    .B(_1658_),
    .C(_1659_),
    .Y(_1660_));
 sg13g2_nor3_1 _2515_ (.A(net1027),
    .B(_1639_),
    .C(_1640_),
    .Y(_1661_));
 sg13g2_nor3_1 _2516_ (.A(net1033),
    .B(_1642_),
    .C(_1643_),
    .Y(_1662_));
 sg13g2_nor3_1 _2517_ (.A(net922),
    .B(_1660_),
    .C(_1661_),
    .Y(_1663_));
 sg13g2_nand2b_2 _2518_ (.Y(_1664_),
    .B(_1647_),
    .A_N(_0038_));
 sg13g2_nand2_1 _2519_ (.Y(_1665_),
    .A(net919),
    .B(_1664_));
 sg13g2_o21ai_1 _2520_ (.B1(net1031),
    .Y(_1666_),
    .A1(_1648_),
    .A2(_1649_));
 sg13g2_nor3_2 _2521_ (.A(net915),
    .B(_1650_),
    .C(_1651_),
    .Y(_1667_));
 sg13g2_a21oi_2 _2522_ (.B1(net1038),
    .Y(_1668_),
    .A2(_1666_),
    .A1(_1665_));
 sg13g2_nor3_1 _2523_ (.A(net1045),
    .B(_1667_),
    .C(_1668_),
    .Y(_1669_));
 sg13g2_nor3_1 _2524_ (.A(net912),
    .B(_1652_),
    .C(_1653_),
    .Y(_1670_));
 sg13g2_nor3_1 _2525_ (.A(net907),
    .B(_1654_),
    .C(_1655_),
    .Y(_1671_));
 sg13g2_nor3_1 _2526_ (.A(net1056),
    .B(_1669_),
    .C(_1670_),
    .Y(_1672_));
 sg13g2_nor3_1 _2527_ (.A(net1020),
    .B(_1656_),
    .C(_1657_),
    .Y(_1673_));
 sg13g2_nor3_1 _2528_ (.A(net931),
    .B(_1441_),
    .C(_1442_),
    .Y(_1674_));
 sg13g2_nor3_1 _2529_ (.A(net927),
    .B(_1673_),
    .C(_1674_),
    .Y(_1675_));
 sg13g2_nor3_1 _2530_ (.A(net1027),
    .B(_1658_),
    .C(_1659_),
    .Y(_1676_));
 sg13g2_nor3_1 _2531_ (.A(net1033),
    .B(_1660_),
    .C(_1661_),
    .Y(_1677_));
 sg13g2_nor3_1 _2532_ (.A(net922),
    .B(_1675_),
    .C(_1676_),
    .Y(_1678_));
 sg13g2_nor3_1 _2533_ (.A(net917),
    .B(_1677_),
    .C(_1678_),
    .Y(_1679_));
 sg13g2_nor3_1 _2534_ (.A(net1041),
    .B(_1662_),
    .C(_1663_),
    .Y(_1680_));
 sg13g2_nor3_2 _2535_ (.A(net917),
    .B(_1662_),
    .C(_1663_),
    .Y(_1681_));
 sg13g2_nor3_2 _2536_ (.A(net1041),
    .B(_1641_),
    .C(_1644_),
    .Y(_1682_));
 sg13g2_nor3_2 _2537_ (.A(net1048),
    .B(_1681_),
    .C(_1682_),
    .Y(_1683_));
 sg13g2_nor3_2 _2538_ (.A(net911),
    .B(_1679_),
    .C(_1680_),
    .Y(_1684_));
 sg13g2_nor3_1 _2539_ (.A(net906),
    .B(_1683_),
    .C(_1684_),
    .Y(_1685_));
 sg13g2_nor3_1 _2540_ (.A(net1047),
    .B(_1645_),
    .C(_1646_),
    .Y(_1686_));
 sg13g2_nor3_2 _2541_ (.A(net911),
    .B(_1681_),
    .C(_1682_),
    .Y(_1687_));
 sg13g2_nor3_1 _2542_ (.A(net1056),
    .B(_1686_),
    .C(_1687_),
    .Y(_1688_));
 sg13g2_nor3_1 _2543_ (.A(net906),
    .B(_1686_),
    .C(_1687_),
    .Y(_1689_));
 sg13g2_nor3_1 _2544_ (.A(net1056),
    .B(_1654_),
    .C(_1655_),
    .Y(_1690_));
 sg13g2_nor3_1 _2545_ (.A(net1063),
    .B(_1689_),
    .C(_1690_),
    .Y(_1691_));
 sg13g2_nor3_1 _2546_ (.A(net901),
    .B(_1685_),
    .C(_1688_),
    .Y(_1692_));
 sg13g2_nor3_1 _2547_ (.A(net894),
    .B(_1691_),
    .C(_1692_),
    .Y(_1693_));
 sg13g2_nor3_1 _2548_ (.A(net1065),
    .B(_1671_),
    .C(_1672_),
    .Y(_1694_));
 sg13g2_nor3_1 _2549_ (.A(net901),
    .B(_1689_),
    .C(_1690_),
    .Y(_1695_));
 sg13g2_nor3_1 _2550_ (.A(net1070),
    .B(_1694_),
    .C(_1695_),
    .Y(_1696_));
 sg13g2_o21ai_1 _2551_ (.B1(net887),
    .Y(_1697_),
    .A1(_1693_),
    .A2(_1696_));
 sg13g2_nor3_1 _2552_ (.A(net927),
    .B(_1443_),
    .C(_1444_),
    .Y(_1698_));
 sg13g2_nor3_1 _2553_ (.A(net1027),
    .B(_1673_),
    .C(_1674_),
    .Y(_1699_));
 sg13g2_nor3_1 _2554_ (.A(net1033),
    .B(_1675_),
    .C(_1676_),
    .Y(_1700_));
 sg13g2_nor3_1 _2555_ (.A(net922),
    .B(_1698_),
    .C(_1699_),
    .Y(_1701_));
 sg13g2_nor3_1 _2556_ (.A(net917),
    .B(_1700_),
    .C(_1701_),
    .Y(_1702_));
 sg13g2_nor3_1 _2557_ (.A(net1041),
    .B(_1677_),
    .C(_1678_),
    .Y(_1703_));
 sg13g2_nor3_1 _2558_ (.A(net1048),
    .B(_1679_),
    .C(_1680_),
    .Y(_1704_));
 sg13g2_nor3_1 _2559_ (.A(net911),
    .B(_1702_),
    .C(_1703_),
    .Y(_1705_));
 sg13g2_nor3_1 _2560_ (.A(net906),
    .B(_1704_),
    .C(_1705_),
    .Y(_1706_));
 sg13g2_nor3_1 _2561_ (.A(net1057),
    .B(_1683_),
    .C(_1684_),
    .Y(_1707_));
 sg13g2_nor3_1 _2562_ (.A(net1064),
    .B(_1685_),
    .C(_1688_),
    .Y(_1708_));
 sg13g2_nor3_1 _2563_ (.A(net901),
    .B(_1706_),
    .C(_1707_),
    .Y(_1709_));
 sg13g2_nor3_1 _2564_ (.A(net894),
    .B(_1708_),
    .C(_1709_),
    .Y(_1710_));
 sg13g2_nor3_1 _2565_ (.A(net1071),
    .B(_1691_),
    .C(_1692_),
    .Y(_1711_));
 sg13g2_o21ai_1 _2566_ (.B1(net1079),
    .Y(_1712_),
    .A1(_1710_),
    .A2(_1711_));
 sg13g2_nand3_1 _2567_ (.B(_1697_),
    .C(_1712_),
    .A(net879),
    .Y(_1713_));
 sg13g2_a221oi_1 _2568_ (.B2(_1713_),
    .C1(_0998_),
    .B1(_1594_),
    .A1(_1560_),
    .Y(_1714_),
    .A2(_1585_));
 sg13g2_and2_1 _2569_ (.A(_0015_),
    .B(net990),
    .X(_1715_));
 sg13g2_a21oi_1 _2570_ (.A1(_1527_),
    .A2(_1528_),
    .Y(_1716_),
    .B1(net990));
 sg13g2_o21ai_1 _2571_ (.B1(net994),
    .Y(_1717_),
    .A1(_1715_),
    .A2(_1716_));
 sg13g2_nand3_1 _2572_ (.B(_1529_),
    .C(_1530_),
    .A(net954),
    .Y(_1718_));
 sg13g2_nand3_1 _2573_ (.B(_1531_),
    .C(_1532_),
    .A(net950),
    .Y(_1719_));
 sg13g2_nand3_1 _2574_ (.B(_1717_),
    .C(_1718_),
    .A(net995),
    .Y(_1720_));
 sg13g2_nand3_1 _2575_ (.B(_1719_),
    .C(_1720_),
    .A(net999),
    .Y(_1721_));
 sg13g2_nand3_1 _2576_ (.B(_1533_),
    .C(_1534_),
    .A(net949),
    .Y(_1722_));
 sg13g2_nand3_1 _2577_ (.B(_1535_),
    .C(_1536_),
    .A(net943),
    .Y(_1723_));
 sg13g2_nand3_1 _2578_ (.B(_1721_),
    .C(_1722_),
    .A(net1005),
    .Y(_1724_));
 sg13g2_nand2_1 _2579_ (.Y(_1725_),
    .A(_0014_),
    .B(net994));
 sg13g2_o21ai_1 _2580_ (.B1(net954),
    .Y(_1726_),
    .A1(_1715_),
    .A2(_1716_));
 sg13g2_nand3_1 _2581_ (.B(_1717_),
    .C(_1718_),
    .A(net950),
    .Y(_1727_));
 sg13g2_nand3_1 _2582_ (.B(_1725_),
    .C(_1726_),
    .A(net995),
    .Y(_1728_));
 sg13g2_nand3_1 _2583_ (.B(_1727_),
    .C(_1728_),
    .A(net999),
    .Y(_1729_));
 sg13g2_nand3_1 _2584_ (.B(_1719_),
    .C(_1720_),
    .A(net949),
    .Y(_1730_));
 sg13g2_nand3_1 _2585_ (.B(_1721_),
    .C(_1722_),
    .A(net943),
    .Y(_1731_));
 sg13g2_nand3_1 _2586_ (.B(_1729_),
    .C(_1730_),
    .A(net1005),
    .Y(_1732_));
 sg13g2_nand3_1 _2587_ (.B(_1731_),
    .C(_1732_),
    .A(net1008),
    .Y(_1733_));
 sg13g2_nand3_1 _2588_ (.B(_1723_),
    .C(_1724_),
    .A(net942),
    .Y(_1734_));
 sg13g2_nand3_1 _2589_ (.B(_1723_),
    .C(_1724_),
    .A(net1007),
    .Y(_1735_));
 sg13g2_nand3_1 _2590_ (.B(_1537_),
    .C(_1538_),
    .A(net942),
    .Y(_1736_));
 sg13g2_nand3_1 _2591_ (.B(_1735_),
    .C(_1736_),
    .A(net937),
    .Y(_1737_));
 sg13g2_nand3_1 _2592_ (.B(_1733_),
    .C(_1734_),
    .A(net1013),
    .Y(_1738_));
 sg13g2_and2_1 _2593_ (.A(_0013_),
    .B(net998),
    .X(_1739_));
 sg13g2_a21oi_1 _2594_ (.A1(_1725_),
    .A2(_1726_),
    .Y(_1740_),
    .B1(net995));
 sg13g2_o21ai_1 _2595_ (.B1(net999),
    .Y(_1741_),
    .A1(_1739_),
    .A2(_1740_));
 sg13g2_nand3_1 _2596_ (.B(_1727_),
    .C(_1728_),
    .A(net949),
    .Y(_1742_));
 sg13g2_nand3_1 _2597_ (.B(_1729_),
    .C(_1730_),
    .A(net943),
    .Y(_1743_));
 sg13g2_nand3_1 _2598_ (.B(_1741_),
    .C(_1742_),
    .A(net1005),
    .Y(_1744_));
 sg13g2_nand3_1 _2599_ (.B(_1743_),
    .C(_1744_),
    .A(net1007),
    .Y(_1745_));
 sg13g2_nand3_1 _2600_ (.B(_1731_),
    .C(_1732_),
    .A(net942),
    .Y(_1746_));
 sg13g2_nand3_1 _2601_ (.B(_1733_),
    .C(_1734_),
    .A(net938),
    .Y(_1747_));
 sg13g2_nand3_1 _2602_ (.B(_1745_),
    .C(_1746_),
    .A(net1013),
    .Y(_1748_));
 sg13g2_nand3_1 _2603_ (.B(_1747_),
    .C(_1748_),
    .A(net1018),
    .Y(_1749_));
 sg13g2_nand3_1 _2604_ (.B(_1737_),
    .C(_1738_),
    .A(net933),
    .Y(_1750_));
 sg13g2_nand3_1 _2605_ (.B(_1539_),
    .C(_1540_),
    .A(net937),
    .Y(_1751_));
 sg13g2_nand3_1 _2606_ (.B(_1735_),
    .C(_1736_),
    .A(net1016),
    .Y(_1752_));
 sg13g2_nand3_1 _2607_ (.B(_1737_),
    .C(_1738_),
    .A(net1018),
    .Y(_1753_));
 sg13g2_nand3_1 _2608_ (.B(_1751_),
    .C(_1752_),
    .A(net932),
    .Y(_1754_));
 sg13g2_nand3_1 _2609_ (.B(_1753_),
    .C(_1754_),
    .A(net928),
    .Y(_1755_));
 sg13g2_nand3_1 _2610_ (.B(_1749_),
    .C(_1750_),
    .A(net1024),
    .Y(_1756_));
 sg13g2_nand2_1 _2611_ (.Y(_1757_),
    .A(_0012_),
    .B(net999));
 sg13g2_o21ai_1 _2612_ (.B1(net949),
    .Y(_1758_),
    .A1(_1739_),
    .A2(_1740_));
 sg13g2_nand3_1 _2613_ (.B(_1741_),
    .C(_1742_),
    .A(net943),
    .Y(_1759_));
 sg13g2_nand3_1 _2614_ (.B(_1757_),
    .C(_1758_),
    .A(net1005),
    .Y(_1760_));
 sg13g2_nand3_1 _2615_ (.B(_1759_),
    .C(_1760_),
    .A(net1007),
    .Y(_1761_));
 sg13g2_nand3_1 _2616_ (.B(_1743_),
    .C(_1744_),
    .A(net942),
    .Y(_1762_));
 sg13g2_nand3_1 _2617_ (.B(_1745_),
    .C(_1746_),
    .A(net934),
    .Y(_1763_));
 sg13g2_nand3_1 _2618_ (.B(_1761_),
    .C(_1762_),
    .A(net1013),
    .Y(_1764_));
 sg13g2_nand3_1 _2619_ (.B(_1763_),
    .C(_1764_),
    .A(net1018),
    .Y(_1765_));
 sg13g2_nand3_1 _2620_ (.B(_1747_),
    .C(_1748_),
    .A(net929),
    .Y(_1766_));
 sg13g2_nand3_1 _2621_ (.B(_1749_),
    .C(_1750_),
    .A(net925),
    .Y(_1767_));
 sg13g2_nand3_1 _2622_ (.B(_1765_),
    .C(_1766_),
    .A(net1024),
    .Y(_1768_));
 sg13g2_nand3_1 _2623_ (.B(_1767_),
    .C(_1768_),
    .A(net1031),
    .Y(_1769_));
 sg13g2_nand3_1 _2624_ (.B(_1755_),
    .C(_1756_),
    .A(net923),
    .Y(_1770_));
 sg13g2_nand3_1 _2625_ (.B(_1751_),
    .C(_1752_),
    .A(net1021),
    .Y(_1771_));
 sg13g2_nand3_1 _2626_ (.B(_1541_),
    .C(_1542_),
    .A(net932),
    .Y(_1772_));
 sg13g2_nand3_1 _2627_ (.B(_1771_),
    .C(_1772_),
    .A(net928),
    .Y(_1773_));
 sg13g2_nand3_1 _2628_ (.B(_1753_),
    .C(_1754_),
    .A(net1028),
    .Y(_1774_));
 sg13g2_nand3_1 _2629_ (.B(_1755_),
    .C(_1756_),
    .A(net1034),
    .Y(_1775_));
 sg13g2_nand3_1 _2630_ (.B(_1773_),
    .C(_1774_),
    .A(net923),
    .Y(_1776_));
 sg13g2_nand3_1 _2631_ (.B(_1775_),
    .C(_1776_),
    .A(net918),
    .Y(_1777_));
 sg13g2_nand3_1 _2632_ (.B(_1769_),
    .C(_1770_),
    .A(net1042),
    .Y(_1778_));
 sg13g2_and2_1 _2633_ (.A(_0011_),
    .B(net1005),
    .X(_1779_));
 sg13g2_a21oi_2 _2634_ (.B1(net1005),
    .Y(_1780_),
    .A2(_1758_),
    .A1(_1757_));
 sg13g2_o21ai_1 _2635_ (.B1(net1007),
    .Y(_1781_),
    .A1(_1779_),
    .A2(_1780_));
 sg13g2_nand3_1 _2636_ (.B(_1759_),
    .C(_1760_),
    .A(net942),
    .Y(_1782_));
 sg13g2_nand3_1 _2637_ (.B(_1761_),
    .C(_1762_),
    .A(net938),
    .Y(_0124_));
 sg13g2_nand3_1 _2638_ (.B(_1781_),
    .C(_1782_),
    .A(net1012),
    .Y(_0125_));
 sg13g2_nand3_1 _2639_ (.B(_0124_),
    .C(_0125_),
    .A(net1018),
    .Y(_0126_));
 sg13g2_nand3_1 _2640_ (.B(_1763_),
    .C(_1764_),
    .A(net929),
    .Y(_0127_));
 sg13g2_nand3_1 _2641_ (.B(_1765_),
    .C(_1766_),
    .A(net925),
    .Y(_0128_));
 sg13g2_nand3_1 _2642_ (.B(_0126_),
    .C(_0127_),
    .A(net1024),
    .Y(_0129_));
 sg13g2_nand3_1 _2643_ (.B(_0128_),
    .C(_0129_),
    .A(net1031),
    .Y(_0130_));
 sg13g2_nand3_1 _2644_ (.B(_1767_),
    .C(_1768_),
    .A(net920),
    .Y(_0131_));
 sg13g2_nand3_1 _2645_ (.B(_1769_),
    .C(_1770_),
    .A(net918),
    .Y(_0132_));
 sg13g2_nand3_1 _2646_ (.B(_0130_),
    .C(_0131_),
    .A(net1038),
    .Y(_0133_));
 sg13g2_nand3_1 _2647_ (.B(_0132_),
    .C(_0133_),
    .A(net1045),
    .Y(_0134_));
 sg13g2_nand3_1 _2648_ (.B(_1777_),
    .C(_1778_),
    .A(net912),
    .Y(_0135_));
 sg13g2_nand3_1 _2649_ (.B(_1543_),
    .C(_1544_),
    .A(net928),
    .Y(_0136_));
 sg13g2_nand3_1 _2650_ (.B(_1771_),
    .C(_1772_),
    .A(net1028),
    .Y(_0137_));
 sg13g2_nand3_1 _2651_ (.B(_1773_),
    .C(_1774_),
    .A(net1034),
    .Y(_0138_));
 sg13g2_nand3_1 _2652_ (.B(_0136_),
    .C(_0137_),
    .A(net923),
    .Y(_0139_));
 sg13g2_nand3_1 _2653_ (.B(_0138_),
    .C(_0139_),
    .A(net918),
    .Y(_0140_));
 sg13g2_nand3_1 _2654_ (.B(_1775_),
    .C(_1776_),
    .A(net1042),
    .Y(_0141_));
 sg13g2_nand3_1 _2655_ (.B(_1777_),
    .C(_1778_),
    .A(net1049),
    .Y(_0142_));
 sg13g2_nand3_1 _2656_ (.B(_0140_),
    .C(_0141_),
    .A(net912),
    .Y(_0143_));
 sg13g2_nand3_1 _2657_ (.B(_0142_),
    .C(_0143_),
    .A(net907),
    .Y(_0144_));
 sg13g2_nand3_1 _2658_ (.B(_0134_),
    .C(_0135_),
    .A(net1056),
    .Y(_0145_));
 sg13g2_nand2_2 _2659_ (.Y(_0146_),
    .A(_0010_),
    .B(net1008));
 sg13g2_o21ai_1 _2660_ (.B1(net942),
    .Y(_0147_),
    .A1(_1779_),
    .A2(_1780_));
 sg13g2_nand3_1 _2661_ (.B(_1781_),
    .C(_1782_),
    .A(net934),
    .Y(_0148_));
 sg13g2_nand3_1 _2662_ (.B(_0146_),
    .C(_0147_),
    .A(net1012),
    .Y(_0149_));
 sg13g2_nand3_1 _2663_ (.B(_0148_),
    .C(_0149_),
    .A(net1018),
    .Y(_0150_));
 sg13g2_nand3_1 _2664_ (.B(_0124_),
    .C(_0125_),
    .A(net933),
    .Y(_0151_));
 sg13g2_nand3_1 _2665_ (.B(_0126_),
    .C(_0127_),
    .A(net925),
    .Y(_0152_));
 sg13g2_nand3_1 _2666_ (.B(_0150_),
    .C(_0151_),
    .A(net1024),
    .Y(_0153_));
 sg13g2_nand3_1 _2667_ (.B(_0152_),
    .C(_0153_),
    .A(net1031),
    .Y(_0154_));
 sg13g2_nand3_1 _2668_ (.B(_0128_),
    .C(_0129_),
    .A(net920),
    .Y(_0155_));
 sg13g2_nand3_1 _2669_ (.B(_0130_),
    .C(_0131_),
    .A(net915),
    .Y(_0156_));
 sg13g2_nand3_1 _2670_ (.B(_0154_),
    .C(_0155_),
    .A(net1038),
    .Y(_0157_));
 sg13g2_nand3_1 _2671_ (.B(_0156_),
    .C(_0157_),
    .A(net1045),
    .Y(_0158_));
 sg13g2_nand3_1 _2672_ (.B(_0132_),
    .C(_0133_),
    .A(net909),
    .Y(_0159_));
 sg13g2_nand3_1 _2673_ (.B(_0134_),
    .C(_0135_),
    .A(net907),
    .Y(_0160_));
 sg13g2_nand3_1 _2674_ (.B(_0158_),
    .C(_0159_),
    .A(net1053),
    .Y(_0161_));
 sg13g2_nand3_1 _2675_ (.B(_0160_),
    .C(_0161_),
    .A(net1060),
    .Y(_0162_));
 sg13g2_nand3_1 _2676_ (.B(_0144_),
    .C(_0145_),
    .A(net900),
    .Y(_0163_));
 sg13g2_and2_1 _2677_ (.A(_0009_),
    .B(net1013),
    .X(_0164_));
 sg13g2_a21oi_1 _2678_ (.A1(_0146_),
    .A2(_0147_),
    .Y(_0165_),
    .B1(net1012));
 sg13g2_o21ai_1 _2679_ (.B1(net1018),
    .Y(_0166_),
    .A1(_0164_),
    .A2(_0165_));
 sg13g2_nand3_1 _2680_ (.B(_0148_),
    .C(_0149_),
    .A(net929),
    .Y(_0167_));
 sg13g2_nand3_1 _2681_ (.B(_0150_),
    .C(_0151_),
    .A(net925),
    .Y(_0168_));
 sg13g2_nand3_1 _2682_ (.B(_0166_),
    .C(_0167_),
    .A(net1024),
    .Y(_0169_));
 sg13g2_nand3_1 _2683_ (.B(_0168_),
    .C(_0169_),
    .A(net1030),
    .Y(_0170_));
 sg13g2_nand3_1 _2684_ (.B(_0152_),
    .C(_0153_),
    .A(net920),
    .Y(_0171_));
 sg13g2_nand3_1 _2685_ (.B(_0154_),
    .C(_0155_),
    .A(net915),
    .Y(_0172_));
 sg13g2_nand3_1 _2686_ (.B(_0170_),
    .C(_0171_),
    .A(net1038),
    .Y(_0173_));
 sg13g2_nand3_1 _2687_ (.B(_0172_),
    .C(_0173_),
    .A(net1045),
    .Y(_0174_));
 sg13g2_nand3_1 _2688_ (.B(_0156_),
    .C(_0157_),
    .A(net909),
    .Y(_0175_));
 sg13g2_nand3_1 _2689_ (.B(_0158_),
    .C(_0159_),
    .A(net904),
    .Y(_0176_));
 sg13g2_nand3_1 _2690_ (.B(_0174_),
    .C(_0175_),
    .A(net1053),
    .Y(_0177_));
 sg13g2_nand3_1 _2691_ (.B(_0176_),
    .C(_0177_),
    .A(net1060),
    .Y(_0178_));
 sg13g2_nand3_1 _2692_ (.B(_0160_),
    .C(_0161_),
    .A(net900),
    .Y(_0179_));
 sg13g2_a21oi_1 _2693_ (.A1(_0178_),
    .A2(_0179_),
    .Y(_0180_),
    .B1(net892));
 sg13g2_a21oi_1 _2694_ (.A1(_0162_),
    .A2(_0163_),
    .Y(_0181_),
    .B1(net1066));
 sg13g2_o21ai_1 _2695_ (.B1(net885),
    .Y(_0182_),
    .A1(_0180_),
    .A2(_0181_));
 sg13g2_nand2_1 _2696_ (.Y(_0183_),
    .A(_0008_),
    .B(net1022));
 sg13g2_o21ai_1 _2697_ (.B1(net929),
    .Y(_0184_),
    .A1(_0164_),
    .A2(_0165_));
 sg13g2_nand3_1 _2698_ (.B(_0166_),
    .C(_0167_),
    .A(net925),
    .Y(_0185_));
 sg13g2_nand3_1 _2699_ (.B(_0183_),
    .C(_0184_),
    .A(net1024),
    .Y(_0186_));
 sg13g2_nand3_1 _2700_ (.B(_0185_),
    .C(_0186_),
    .A(net1030),
    .Y(_0187_));
 sg13g2_nand3_1 _2701_ (.B(_0168_),
    .C(_0169_),
    .A(net920),
    .Y(_0188_));
 sg13g2_nand3_1 _2702_ (.B(_0170_),
    .C(_0171_),
    .A(net915),
    .Y(_0189_));
 sg13g2_nand3_1 _2703_ (.B(_0187_),
    .C(_0188_),
    .A(net1037),
    .Y(_0190_));
 sg13g2_nand3_1 _2704_ (.B(_0189_),
    .C(_0190_),
    .A(net1045),
    .Y(_0191_));
 sg13g2_nand3_1 _2705_ (.B(_0172_),
    .C(_0173_),
    .A(net909),
    .Y(_0192_));
 sg13g2_nand3_1 _2706_ (.B(_0174_),
    .C(_0175_),
    .A(net904),
    .Y(_0193_));
 sg13g2_nand3_1 _2707_ (.B(_0191_),
    .C(_0192_),
    .A(net1053),
    .Y(_0194_));
 sg13g2_nand3_1 _2708_ (.B(_0193_),
    .C(_0194_),
    .A(net1060),
    .Y(_0195_));
 sg13g2_nand3_1 _2709_ (.B(_0176_),
    .C(_0177_),
    .A(net898),
    .Y(_0196_));
 sg13g2_a21oi_1 _2710_ (.A1(_0195_),
    .A2(_0196_),
    .Y(_0197_),
    .B1(net892));
 sg13g2_a21oi_1 _2711_ (.A1(_0178_),
    .A2(_0179_),
    .Y(_0198_),
    .B1(net1066));
 sg13g2_o21ai_1 _2712_ (.B1(net1073),
    .Y(_0199_),
    .A1(_0197_),
    .A2(_0198_));
 sg13g2_nand3_1 _2713_ (.B(_0182_),
    .C(_0199_),
    .A(net877),
    .Y(_0200_));
 sg13g2_and2_1 _2714_ (.A(\a[15] ),
    .B(net990),
    .X(_0201_));
 sg13g2_nand2_2 _2715_ (.Y(_0202_),
    .A(net993),
    .B(_0201_));
 sg13g2_o21ai_1 _2716_ (.B1(_1725_),
    .Y(_0203_),
    .A1(net994),
    .A2(_0201_));
 sg13g2_and2_1 _2717_ (.A(net995),
    .B(_0203_),
    .X(_0204_));
 sg13g2_a21oi_1 _2718_ (.A1(net950),
    .A2(_0202_),
    .Y(_0205_),
    .B1(_0204_));
 sg13g2_o21ai_1 _2719_ (.B1(net948),
    .Y(_0206_),
    .A1(_0044_),
    .A2(_0202_));
 sg13g2_o21ai_1 _2720_ (.B1(_0206_),
    .Y(_0207_),
    .A1(net949),
    .A2(_0205_));
 sg13g2_a21oi_1 _2721_ (.A1(net950),
    .A2(_0203_),
    .Y(_0208_),
    .B1(_1739_));
 sg13g2_mux2_1 _2722_ (.A0(_0205_),
    .A1(_0208_),
    .S(net999),
    .X(_0209_));
 sg13g2_nand2_1 _2723_ (.Y(_0210_),
    .A(net1004),
    .B(_0209_));
 sg13g2_o21ai_1 _2724_ (.B1(_0210_),
    .Y(_0211_),
    .A1(net1004),
    .A2(_0207_));
 sg13g2_nor3_2 _2725_ (.A(_0044_),
    .B(_0043_),
    .C(_0202_),
    .Y(_0212_));
 sg13g2_nor2_1 _2726_ (.A(net945),
    .B(_0207_),
    .Y(_0213_));
 sg13g2_a21oi_2 _2727_ (.B1(_0213_),
    .Y(_0214_),
    .A2(_0212_),
    .A1(net945));
 sg13g2_nor2_1 _2728_ (.A(net1011),
    .B(_0214_),
    .Y(_0215_));
 sg13g2_a21oi_2 _2729_ (.B1(_0215_),
    .Y(_0216_),
    .A2(_0211_),
    .A1(net1011));
 sg13g2_nor2_1 _2730_ (.A(net1012),
    .B(_0216_),
    .Y(_0217_));
 sg13g2_o21ai_1 _2731_ (.B1(_1757_),
    .Y(_0218_),
    .A1(net999),
    .A2(_0208_));
 sg13g2_nor2_1 _2732_ (.A(net943),
    .B(_0218_),
    .Y(_0219_));
 sg13g2_a21oi_2 _2733_ (.B1(_0219_),
    .Y(_0220_),
    .A2(_0209_),
    .A1(net943));
 sg13g2_nor2_1 _2734_ (.A(net1011),
    .B(_0211_),
    .Y(_0221_));
 sg13g2_a21oi_1 _2735_ (.A1(net1007),
    .A2(_0220_),
    .Y(_0222_),
    .B1(_0221_));
 sg13g2_a21oi_1 _2736_ (.A1(net1012),
    .A2(_0222_),
    .Y(_0223_),
    .B1(_0217_));
 sg13g2_nand2_1 _2737_ (.Y(_0224_),
    .A(net1017),
    .B(_0223_));
 sg13g2_nor2b_1 _2738_ (.A(_0042_),
    .B_N(_0212_),
    .Y(_0225_));
 sg13g2_nor2_1 _2739_ (.A(net1009),
    .B(_0225_),
    .Y(_0226_));
 sg13g2_a21oi_2 _2740_ (.B1(_0226_),
    .Y(_0227_),
    .A2(_0214_),
    .A1(net1009));
 sg13g2_nand2_1 _2741_ (.Y(_0228_),
    .A(net934),
    .B(_0227_));
 sg13g2_o21ai_1 _2742_ (.B1(_0228_),
    .Y(_0229_),
    .A1(net934),
    .A2(_0216_));
 sg13g2_o21ai_1 _2743_ (.B1(_0224_),
    .Y(_0230_),
    .A1(net1017),
    .A2(_0229_));
 sg13g2_nor2_1 _2744_ (.A(net1023),
    .B(_0230_),
    .Y(_0231_));
 sg13g2_a21oi_2 _2745_ (.B1(_1779_),
    .Y(_0232_),
    .A2(_0218_),
    .A1(net943));
 sg13g2_nand2_1 _2746_ (.Y(_0233_),
    .A(net1007),
    .B(_0232_));
 sg13g2_o21ai_1 _2747_ (.B1(_0233_),
    .Y(_0234_),
    .A1(net1007),
    .A2(_0220_));
 sg13g2_and2_1 _2748_ (.A(net1012),
    .B(_0234_),
    .X(_0235_));
 sg13g2_a21oi_1 _2749_ (.A1(net934),
    .A2(_0222_),
    .Y(_0236_),
    .B1(_0235_));
 sg13g2_and2_1 _2750_ (.A(net1017),
    .B(_0236_),
    .X(_0237_));
 sg13g2_a21oi_1 _2751_ (.A1(net929),
    .A2(_0223_),
    .Y(_0238_),
    .B1(_0237_));
 sg13g2_a21oi_1 _2752_ (.A1(net1023),
    .A2(_0238_),
    .Y(_0239_),
    .B1(_0231_));
 sg13g2_nand2_1 _2753_ (.Y(_0240_),
    .A(net1029),
    .B(_0239_));
 sg13g2_nand2b_2 _2754_ (.Y(_0241_),
    .B(_0225_),
    .A_N(_0041_));
 sg13g2_nor2_1 _2755_ (.A(net1012),
    .B(_0241_),
    .Y(_0242_));
 sg13g2_a21oi_1 _2756_ (.A1(net1012),
    .A2(_0227_),
    .Y(_0243_),
    .B1(_0242_));
 sg13g2_nand2_1 _2757_ (.Y(_0244_),
    .A(net929),
    .B(_0243_));
 sg13g2_o21ai_1 _2758_ (.B1(_0244_),
    .Y(_0245_),
    .A1(net929),
    .A2(_0229_));
 sg13g2_nand2b_1 _2759_ (.Y(_0246_),
    .B(net924),
    .A_N(_0245_));
 sg13g2_o21ai_1 _2760_ (.B1(_0246_),
    .Y(_0247_),
    .A1(net924),
    .A2(_0230_));
 sg13g2_o21ai_1 _2761_ (.B1(_0240_),
    .Y(_0248_),
    .A1(net1029),
    .A2(_0247_));
 sg13g2_nor2_1 _2762_ (.A(net1036),
    .B(_0248_),
    .Y(_0249_));
 sg13g2_o21ai_1 _2763_ (.B1(_0146_),
    .Y(_0250_),
    .A1(net1007),
    .A2(_0232_));
 sg13g2_nor2_1 _2764_ (.A(net934),
    .B(_0250_),
    .Y(_0251_));
 sg13g2_a21oi_1 _2765_ (.A1(net934),
    .A2(_0234_),
    .Y(_0252_),
    .B1(_0251_));
 sg13g2_and2_1 _2766_ (.A(net1017),
    .B(_0252_),
    .X(_0253_));
 sg13g2_a21oi_1 _2767_ (.A1(net929),
    .A2(_0236_),
    .Y(_0254_),
    .B1(_0253_));
 sg13g2_and2_1 _2768_ (.A(net1023),
    .B(_0254_),
    .X(_0255_));
 sg13g2_a21oi_1 _2769_ (.A1(net924),
    .A2(_0238_),
    .Y(_0256_),
    .B1(_0255_));
 sg13g2_and2_1 _2770_ (.A(net1029),
    .B(_0256_),
    .X(_0257_));
 sg13g2_a21oi_1 _2771_ (.A1(net919),
    .A2(_0239_),
    .Y(_0258_),
    .B1(_0257_));
 sg13g2_a21oi_1 _2772_ (.A1(net1036),
    .A2(_0258_),
    .Y(_0259_),
    .B1(_0249_));
 sg13g2_or2_1 _2773_ (.X(_0260_),
    .B(_0247_),
    .A(net919));
 sg13g2_nand2_1 _2774_ (.Y(_0261_),
    .A(net1017),
    .B(_0243_));
 sg13g2_o21ai_1 _2775_ (.B1(net933),
    .Y(_0262_),
    .A1(_0040_),
    .A2(_0241_));
 sg13g2_nand2_1 _2776_ (.Y(_0263_),
    .A(_0261_),
    .B(_0262_));
 sg13g2_nand3_1 _2777_ (.B(_0261_),
    .C(_0262_),
    .A(net924),
    .Y(_0264_));
 sg13g2_o21ai_1 _2778_ (.B1(_0264_),
    .Y(_0265_),
    .A1(net924),
    .A2(_0245_));
 sg13g2_o21ai_1 _2779_ (.B1(_0260_),
    .Y(_0266_),
    .A1(net1029),
    .A2(_0265_));
 sg13g2_or2_1 _2780_ (.X(_0267_),
    .B(_0248_),
    .A(net913));
 sg13g2_o21ai_1 _2781_ (.B1(_0267_),
    .Y(_0268_),
    .A1(net1036),
    .A2(_0266_));
 sg13g2_nor2_1 _2782_ (.A(net1043),
    .B(_0268_),
    .Y(_0269_));
 sg13g2_a21oi_1 _2783_ (.A1(net1043),
    .A2(_0259_),
    .Y(_0270_),
    .B1(_0269_));
 sg13g2_a21oi_1 _2784_ (.A1(net934),
    .A2(_0250_),
    .Y(_0271_),
    .B1(_0164_));
 sg13g2_nand2_1 _2785_ (.Y(_0272_),
    .A(net1017),
    .B(_0271_));
 sg13g2_o21ai_1 _2786_ (.B1(_0272_),
    .Y(_0273_),
    .A1(net1017),
    .A2(_0252_));
 sg13g2_and2_1 _2787_ (.A(net1023),
    .B(_0273_),
    .X(_0274_));
 sg13g2_a21oi_1 _2788_ (.A1(net924),
    .A2(_0254_),
    .Y(_0275_),
    .B1(_0274_));
 sg13g2_mux2_1 _2789_ (.A0(_0256_),
    .A1(_0275_),
    .S(net1029),
    .X(_0276_));
 sg13g2_nor2_1 _2790_ (.A(net913),
    .B(_0276_),
    .Y(_0277_));
 sg13g2_a21oi_1 _2791_ (.A1(net913),
    .A2(_0258_),
    .Y(_0278_),
    .B1(_0277_));
 sg13g2_mux2_1 _2792_ (.A0(_0259_),
    .A1(_0278_),
    .S(net1045),
    .X(_0279_));
 sg13g2_nor2_1 _2793_ (.A(net903),
    .B(_0279_),
    .Y(_0280_));
 sg13g2_a21oi_1 _2794_ (.A1(net902),
    .A2(_0270_),
    .Y(_0281_),
    .B1(_0280_));
 sg13g2_nand2_1 _2795_ (.Y(_0282_),
    .A(net1059),
    .B(_0281_));
 sg13g2_nor3_2 _2796_ (.A(_0040_),
    .B(_0039_),
    .C(_0241_),
    .Y(_0283_));
 sg13g2_nor2_1 _2797_ (.A(net1023),
    .B(_0283_),
    .Y(_0284_));
 sg13g2_a21oi_1 _2798_ (.A1(net1023),
    .A2(_0263_),
    .Y(_0285_),
    .B1(_0284_));
 sg13g2_nand2b_1 _2799_ (.Y(_0286_),
    .B(net919),
    .A_N(_0285_));
 sg13g2_o21ai_1 _2800_ (.B1(_0286_),
    .Y(_0287_),
    .A1(net919),
    .A2(_0265_));
 sg13g2_mux2_1 _2801_ (.A0(_0266_),
    .A1(_0287_),
    .S(net913),
    .X(_0288_));
 sg13g2_nor2_1 _2802_ (.A(net1043),
    .B(_0288_),
    .Y(_0289_));
 sg13g2_a21oi_1 _2803_ (.A1(net1043),
    .A2(_0268_),
    .Y(_0290_),
    .B1(_0289_));
 sg13g2_nand2_1 _2804_ (.Y(_0291_),
    .A(net1051),
    .B(_0270_));
 sg13g2_o21ai_1 _2805_ (.B1(_0291_),
    .Y(_0292_),
    .A1(net1051),
    .A2(_0290_));
 sg13g2_o21ai_1 _2806_ (.B1(_0282_),
    .Y(_0293_),
    .A1(net1058),
    .A2(_0292_));
 sg13g2_nor2_1 _2807_ (.A(net1067),
    .B(_0293_),
    .Y(_0294_));
 sg13g2_o21ai_1 _2808_ (.B1(_0183_),
    .Y(_0295_),
    .A1(net1017),
    .A2(_0271_));
 sg13g2_nor2_1 _2809_ (.A(net924),
    .B(_0295_),
    .Y(_0296_));
 sg13g2_a21oi_1 _2810_ (.A1(net925),
    .A2(_0273_),
    .Y(_0297_),
    .B1(_0296_));
 sg13g2_mux2_1 _2811_ (.A0(_0275_),
    .A1(_0297_),
    .S(net1029),
    .X(_0298_));
 sg13g2_or2_1 _2812_ (.X(_0299_),
    .B(_0298_),
    .A(net914));
 sg13g2_o21ai_1 _2813_ (.B1(_0299_),
    .Y(_0300_),
    .A1(net1036),
    .A2(_0276_));
 sg13g2_nor2_1 _2814_ (.A(net908),
    .B(_0300_),
    .Y(_0301_));
 sg13g2_a21oi_1 _2815_ (.A1(net908),
    .A2(_0278_),
    .Y(_0302_),
    .B1(_0301_));
 sg13g2_nand2_1 _2816_ (.Y(_0303_),
    .A(net1051),
    .B(_0302_));
 sg13g2_o21ai_1 _2817_ (.B1(_0303_),
    .Y(_0304_),
    .A1(net1051),
    .A2(_0279_));
 sg13g2_nor2_1 _2818_ (.A(net896),
    .B(_0304_),
    .Y(_0305_));
 sg13g2_a21oi_2 _2819_ (.B1(_0305_),
    .Y(_0306_),
    .A2(_0281_),
    .A1(net896));
 sg13g2_a21oi_2 _2820_ (.B1(_0294_),
    .Y(_0307_),
    .A2(_0306_),
    .A1(net1067));
 sg13g2_nor2b_1 _2821_ (.A(_0038_),
    .B_N(_0283_),
    .Y(_0308_));
 sg13g2_or2_1 _2822_ (.X(_0309_),
    .B(_0308_),
    .A(net1029));
 sg13g2_o21ai_1 _2823_ (.B1(_0309_),
    .Y(_0310_),
    .A1(net919),
    .A2(_0285_));
 sg13g2_nand2b_1 _2824_ (.Y(_0311_),
    .B(net913),
    .A_N(_0310_));
 sg13g2_o21ai_1 _2825_ (.B1(_0311_),
    .Y(_0312_),
    .A1(net913),
    .A2(_0287_));
 sg13g2_nor2_1 _2826_ (.A(net1043),
    .B(_0312_),
    .Y(_0313_));
 sg13g2_a21oi_1 _2827_ (.A1(net1043),
    .A2(_0288_),
    .Y(_0314_),
    .B1(_0313_));
 sg13g2_nor2_1 _2828_ (.A(net1052),
    .B(_0314_),
    .Y(_0315_));
 sg13g2_a21oi_1 _2829_ (.A1(net1051),
    .A2(_0290_),
    .Y(_0316_),
    .B1(_0315_));
 sg13g2_nand2b_1 _2830_ (.Y(_0317_),
    .B(net896),
    .A_N(_0316_));
 sg13g2_o21ai_1 _2831_ (.B1(_0317_),
    .Y(_0318_),
    .A1(net896),
    .A2(_0292_));
 sg13g2_nand2b_1 _2832_ (.Y(_0319_),
    .B(net891),
    .A_N(_0318_));
 sg13g2_o21ai_1 _2833_ (.B1(_0319_),
    .Y(_0320_),
    .A1(net891),
    .A2(_0293_));
 sg13g2_o21ai_1 _2834_ (.B1(net876),
    .Y(_0321_),
    .A1(net1075),
    .A2(_0320_));
 sg13g2_a21o_1 _2835_ (.A2(_0307_),
    .A1(net1075),
    .B1(_0321_),
    .X(_0322_));
 sg13g2_nand2_1 _2836_ (.Y(_0323_),
    .A(net1098),
    .B(\a[8] ));
 sg13g2_nor2_1 _2837_ (.A(net1086),
    .B(_0323_),
    .Y(_0324_));
 sg13g2_a21oi_1 _2838_ (.A1(net1088),
    .A2(_0323_),
    .Y(_0325_),
    .B1(_0324_));
 sg13g2_nor2_1 _2839_ (.A(\a[9] ),
    .B(net1088),
    .Y(_0326_));
 sg13g2_o21ai_1 _2840_ (.B1(\a[8] ),
    .Y(_0327_),
    .A1(net859),
    .A2(_0326_));
 sg13g2_a22oi_1 _2841_ (.Y(_0328_),
    .B1(_0325_),
    .B2(\a[9] ),
    .A2(net867),
    .A1(net1050));
 sg13g2_a221oi_1 _2842_ (.B2(net1022),
    .C1(net1096),
    .B1(net850),
    .A1(\ayayayayayaya.b[20] ),
    .Y(_0329_),
    .A2(net862));
 sg13g2_and4_1 _2843_ (.A(_0322_),
    .B(_0327_),
    .C(_0328_),
    .D(_0329_),
    .X(_0330_));
 sg13g2_and2_1 _2844_ (.A(_0001_),
    .B(net1068),
    .X(_0331_));
 sg13g2_nand2_1 _2845_ (.Y(_0332_),
    .A(_0002_),
    .B(net1061));
 sg13g2_and2_1 _2846_ (.A(_0003_),
    .B(net1054),
    .X(_0333_));
 sg13g2_nand2_1 _2847_ (.Y(_0334_),
    .A(_0004_),
    .B(net1050));
 sg13g2_and2_2 _2848_ (.A(_0005_),
    .B(net1039),
    .X(_0335_));
 sg13g2_nand2_2 _2849_ (.Y(_0336_),
    .A(_0006_),
    .B(net1035));
 sg13g2_and2_1 _2850_ (.A(_0007_),
    .B(net1025),
    .X(_0337_));
 sg13g2_a21oi_1 _2851_ (.A1(_0183_),
    .A2(_0184_),
    .Y(_0338_),
    .B1(net1024));
 sg13g2_o21ai_1 _2852_ (.B1(net919),
    .Y(_0339_),
    .A1(_0337_),
    .A2(_0338_));
 sg13g2_a21oi_1 _2853_ (.A1(_0336_),
    .A2(_0339_),
    .Y(_0340_),
    .B1(net1037));
 sg13g2_o21ai_1 _2854_ (.B1(net908),
    .Y(_0341_),
    .A1(_0335_),
    .A2(_0340_));
 sg13g2_a21oi_1 _2855_ (.A1(_0334_),
    .A2(_0341_),
    .Y(_0342_),
    .B1(net1054));
 sg13g2_o21ai_1 _2856_ (.B1(net897),
    .Y(_0343_),
    .A1(_0333_),
    .A2(_0342_));
 sg13g2_a21oi_1 _2857_ (.A1(_0332_),
    .A2(_0343_),
    .Y(_0344_),
    .B1(net1067));
 sg13g2_o21ai_1 _2858_ (.B1(net882),
    .Y(_0345_),
    .A1(_0331_),
    .A2(_0344_));
 sg13g2_a21oi_1 _2859_ (.A1(_0000_),
    .A2(net1077),
    .Y(_0346_),
    .B1(_1526_));
 sg13g2_a21oi_1 _2860_ (.A1(net925),
    .A2(_0295_),
    .Y(_0347_),
    .B1(_0337_));
 sg13g2_o21ai_1 _2861_ (.B1(_0336_),
    .Y(_0348_),
    .A1(net1030),
    .A2(_0347_));
 sg13g2_a21oi_1 _2862_ (.A1(net914),
    .A2(_0348_),
    .Y(_0349_),
    .B1(_0335_));
 sg13g2_nor2_1 _2863_ (.A(net1046),
    .B(_0349_),
    .Y(_0350_));
 sg13g2_a21oi_1 _2864_ (.A1(_0004_),
    .A2(net1046),
    .Y(_0351_),
    .B1(_0350_));
 sg13g2_nor2_1 _2865_ (.A(net1054),
    .B(_0351_),
    .Y(_0352_));
 sg13g2_nor2_1 _2866_ (.A(_0333_),
    .B(_0352_),
    .Y(_0353_));
 sg13g2_o21ai_1 _2867_ (.B1(_0332_),
    .Y(_0354_),
    .A1(net1061),
    .A2(_0353_));
 sg13g2_a21oi_1 _2868_ (.A1(net890),
    .A2(_0354_),
    .Y(_0355_),
    .B1(_0331_));
 sg13g2_inv_1 _2869_ (.Y(_0356_),
    .A(_0355_));
 sg13g2_a21oi_1 _2870_ (.A1(_0000_),
    .A2(net1077),
    .Y(_0357_),
    .B1(net873));
 sg13g2_o21ai_1 _2871_ (.B1(_0357_),
    .Y(_0358_),
    .A1(net1074),
    .A2(_0355_));
 sg13g2_nand2b_1 _2872_ (.Y(_0359_),
    .B(_1583_),
    .A_N(net868));
 sg13g2_and2_1 _2873_ (.A(net1099),
    .B(\a[1] ),
    .X(_0360_));
 sg13g2_nor2_1 _2874_ (.A(net1083),
    .B(net1093),
    .Y(_0361_));
 sg13g2_o21ai_1 _2875_ (.B1(net858),
    .Y(_0362_),
    .A1(net1088),
    .A2(_0360_));
 sg13g2_nand2b_1 _2876_ (.Y(_0363_),
    .B(net1083),
    .A_N(net855));
 sg13g2_a22oi_1 _2877_ (.Y(_0364_),
    .B1(_0363_),
    .B2(\a[1] ),
    .A2(_0362_),
    .A1(net1083));
 sg13g2_a221oi_1 _2878_ (.B2(net1076),
    .C1(net1104),
    .B1(_0359_),
    .A1(\ayayayayayaya.b[16] ),
    .Y(_0365_),
    .A2(net862));
 sg13g2_o21ai_1 _2879_ (.B1(_0365_),
    .Y(_0366_),
    .A1(_0361_),
    .A2(_0364_));
 sg13g2_a21oi_1 _2880_ (.A1(_0345_),
    .A2(_0346_),
    .Y(_0367_),
    .B1(_0366_));
 sg13g2_a22oi_1 _2881_ (.Y(_0368_),
    .B1(_0358_),
    .B2(_0367_),
    .A2(_0330_),
    .A1(_0200_));
 sg13g2_a21o_2 _2882_ (.A2(_0368_),
    .A1(_0998_),
    .B1(_1714_),
    .X(uio_out[0]));
 sg13g2_a22oi_1 _2883_ (.Y(_0369_),
    .B1(net865),
    .B2(\a[28] ),
    .A2(net871),
    .A1(\a[12] ));
 sg13g2_a21oi_1 _2884_ (.A1(net968),
    .A2(net853),
    .Y(_0370_),
    .B1(net1095));
 sg13g2_and2_1 _2885_ (.A(net1102),
    .B(\a[26] ),
    .X(_0371_));
 sg13g2_a21oi_1 _2886_ (.A1(\a[25] ),
    .A2(_0371_),
    .Y(_0372_),
    .B1(net1092));
 sg13g2_o21ai_1 _2887_ (.B1(_0372_),
    .Y(_0373_),
    .A1(\a[25] ),
    .A2(\a[26] ));
 sg13g2_nand2_1 _2888_ (.Y(_0374_),
    .A(net1087),
    .B(_0371_));
 sg13g2_nand2_1 _2889_ (.Y(_0375_),
    .A(net857),
    .B(_0374_));
 sg13g2_nand3_1 _2890_ (.B(_0370_),
    .C(_0373_),
    .A(_0369_),
    .Y(_0376_));
 sg13g2_a221oi_1 _2891_ (.B2(\a[25] ),
    .C1(_0376_),
    .B1(_0375_),
    .A1(_1171_),
    .Y(_0377_),
    .A2(net876));
 sg13g2_o21ai_1 _2892_ (.B1(net1079),
    .Y(_0378_),
    .A1(_1693_),
    .A2(_1696_));
 sg13g2_o21ai_1 _2893_ (.B1(net1046),
    .Y(_0379_),
    .A1(_1667_),
    .A2(_1668_));
 sg13g2_nor2_1 _2894_ (.A(_0037_),
    .B(_1664_),
    .Y(_0380_));
 sg13g2_nor2_1 _2895_ (.A(net1036),
    .B(_0380_),
    .Y(_0381_));
 sg13g2_a21oi_2 _2896_ (.B1(net915),
    .Y(_0382_),
    .A2(_1666_),
    .A1(_1665_));
 sg13g2_o21ai_1 _2897_ (.B1(net909),
    .Y(_0383_),
    .A1(_0381_),
    .A2(_0382_));
 sg13g2_nor3_1 _2898_ (.A(net907),
    .B(_1669_),
    .C(_1670_),
    .Y(_0384_));
 sg13g2_nor3_1 _2899_ (.A(net1046),
    .B(_0381_),
    .C(_0382_),
    .Y(_0385_));
 sg13g2_nor3_1 _2900_ (.A(net909),
    .B(_1667_),
    .C(_1668_),
    .Y(_0386_));
 sg13g2_nor3_1 _2901_ (.A(net1053),
    .B(_0385_),
    .C(_0386_),
    .Y(_0387_));
 sg13g2_nor3_1 _2902_ (.A(net1065),
    .B(_0384_),
    .C(_0387_),
    .Y(_0388_));
 sg13g2_nor3_1 _2903_ (.A(net900),
    .B(_1671_),
    .C(_1672_),
    .Y(_0389_));
 sg13g2_nor3_1 _2904_ (.A(net894),
    .B(_1694_),
    .C(_1695_),
    .Y(_0390_));
 sg13g2_nor3_1 _2905_ (.A(net1072),
    .B(_0388_),
    .C(_0389_),
    .Y(_0391_));
 sg13g2_o21ai_1 _2906_ (.B1(net886),
    .Y(_0392_),
    .A1(_0390_),
    .A2(_0391_));
 sg13g2_nand3_1 _2907_ (.B(_0378_),
    .C(_0392_),
    .A(net879),
    .Y(_0393_));
 sg13g2_o21ai_1 _2908_ (.B1(net1078),
    .Y(_0394_),
    .A1(_1521_),
    .A2(_1522_));
 sg13g2_nor3_1 _2909_ (.A(net1033),
    .B(_1698_),
    .C(_1699_),
    .Y(_0395_));
 sg13g2_nor3_1 _2910_ (.A(net922),
    .B(_1445_),
    .C(_1446_),
    .Y(_0396_));
 sg13g2_nor3_1 _2911_ (.A(net916),
    .B(_1447_),
    .C(_1448_),
    .Y(_0397_));
 sg13g2_nor3_1 _2912_ (.A(net1040),
    .B(_0395_),
    .C(_0396_),
    .Y(_0398_));
 sg13g2_nor3_1 _2913_ (.A(net1047),
    .B(_0397_),
    .C(_0398_),
    .Y(_0399_));
 sg13g2_nor3_1 _2914_ (.A(net910),
    .B(_1449_),
    .C(_1450_),
    .Y(_0400_));
 sg13g2_a21oi_1 _2915_ (.A1(_1451_),
    .A2(_1452_),
    .Y(_0401_),
    .B1(net905));
 sg13g2_nor3_1 _2916_ (.A(net1055),
    .B(_0399_),
    .C(_0400_),
    .Y(_0402_));
 sg13g2_nor3_1 _2917_ (.A(net1063),
    .B(_0401_),
    .C(_0402_),
    .Y(_0403_));
 sg13g2_a21oi_1 _2918_ (.A1(_1453_),
    .A2(_1454_),
    .Y(_0404_),
    .B1(net899));
 sg13g2_a21oi_1 _2919_ (.A1(_1487_),
    .A2(_1488_),
    .Y(_0405_),
    .B1(net893));
 sg13g2_nor3_1 _2920_ (.A(net1070),
    .B(_0403_),
    .C(_0404_),
    .Y(_0406_));
 sg13g2_o21ai_1 _2921_ (.B1(net886),
    .Y(_0407_),
    .A1(_0405_),
    .A2(_0406_));
 sg13g2_nand3_1 _2922_ (.B(_0394_),
    .C(_0407_),
    .A(net879),
    .Y(_0408_));
 sg13g2_nand3_1 _2923_ (.B(_1492_),
    .C(net875),
    .A(_1491_),
    .Y(_0409_));
 sg13g2_a21oi_1 _2924_ (.A1(net1101),
    .A2(\a[17] ),
    .Y(_0410_),
    .B1(net1090));
 sg13g2_o21ai_1 _2925_ (.B1(\a[18] ),
    .Y(_0411_),
    .A1(_1580_),
    .A2(_0410_));
 sg13g2_o21ai_1 _2926_ (.B1(net857),
    .Y(_0412_),
    .A1(\a[18] ),
    .A2(net1090));
 sg13g2_a22oi_1 _2927_ (.Y(_0413_),
    .B1(net850),
    .B2(\ayayayayayaya.b[17] ),
    .A2(net867),
    .A1(\a[8] ));
 sg13g2_a22oi_1 _2928_ (.Y(_0414_),
    .B1(_0412_),
    .B2(\a[17] ),
    .A2(net864),
    .A1(\a[24] ));
 sg13g2_and3_1 _2929_ (.X(_0415_),
    .A(_0999_),
    .B(_0411_),
    .C(_0414_));
 sg13g2_nand4_1 _2930_ (.B(_0409_),
    .C(_0413_),
    .A(_0408_),
    .Y(_0416_),
    .D(_0415_));
 sg13g2_a21oi_1 _2931_ (.A1(_0377_),
    .A2(_0393_),
    .Y(_0417_),
    .B1(_0998_));
 sg13g2_o21ai_1 _2932_ (.B1(net1030),
    .Y(_0418_),
    .A1(_0337_),
    .A2(_0338_));
 sg13g2_nand3_1 _2933_ (.B(_0185_),
    .C(_0186_),
    .A(net920),
    .Y(_0419_));
 sg13g2_nand3_1 _2934_ (.B(_0418_),
    .C(_0419_),
    .A(net914),
    .Y(_0420_));
 sg13g2_nand3_1 _2935_ (.B(_0336_),
    .C(_0339_),
    .A(net1037),
    .Y(_0421_));
 sg13g2_o21ai_1 _2936_ (.B1(net1046),
    .Y(_0422_),
    .A1(_0335_),
    .A2(_0340_));
 sg13g2_nand3_1 _2937_ (.B(_0420_),
    .C(_0421_),
    .A(net908),
    .Y(_0423_));
 sg13g2_nand3_1 _2938_ (.B(_0422_),
    .C(_0423_),
    .A(net902),
    .Y(_0424_));
 sg13g2_nand3_1 _2939_ (.B(_0334_),
    .C(_0341_),
    .A(net1054),
    .Y(_0425_));
 sg13g2_o21ai_1 _2940_ (.B1(net1061),
    .Y(_0426_),
    .A1(_0333_),
    .A2(_0342_));
 sg13g2_nand3_1 _2941_ (.B(_0424_),
    .C(_0425_),
    .A(net897),
    .Y(_0427_));
 sg13g2_a21oi_1 _2942_ (.A1(_0332_),
    .A2(_0343_),
    .Y(_0428_),
    .B1(net890));
 sg13g2_a21oi_1 _2943_ (.A1(_0426_),
    .A2(_0427_),
    .Y(_0429_),
    .B1(net1067));
 sg13g2_o21ai_1 _2944_ (.B1(net884),
    .Y(_0430_),
    .A1(_0428_),
    .A2(_0429_));
 sg13g2_o21ai_1 _2945_ (.B1(net1074),
    .Y(_0431_),
    .A1(_0331_),
    .A2(_0344_));
 sg13g2_nand3_1 _2946_ (.B(_0430_),
    .C(_0431_),
    .A(net878),
    .Y(_0432_));
 sg13g2_o21ai_1 _2947_ (.B1(net1061),
    .Y(_0433_),
    .A1(_0333_),
    .A2(_0352_));
 sg13g2_nand2_1 _2948_ (.Y(_0434_),
    .A(net1030),
    .B(_0347_));
 sg13g2_o21ai_1 _2949_ (.B1(_0434_),
    .Y(_0435_),
    .A1(net1030),
    .A2(_0297_));
 sg13g2_nor2_1 _2950_ (.A(net914),
    .B(_0348_),
    .Y(_0436_));
 sg13g2_a21oi_1 _2951_ (.A1(net913),
    .A2(_0435_),
    .Y(_0437_),
    .B1(_0436_));
 sg13g2_nand2_1 _2952_ (.Y(_0438_),
    .A(net1046),
    .B(_0349_));
 sg13g2_o21ai_1 _2953_ (.B1(_0438_),
    .Y(_0439_),
    .A1(net1044),
    .A2(_0437_));
 sg13g2_mux2_1 _2954_ (.A0(_0351_),
    .A1(_0439_),
    .S(net902),
    .X(_0440_));
 sg13g2_o21ai_1 _2955_ (.B1(_0433_),
    .Y(_0441_),
    .A1(net1061),
    .A2(_0440_));
 sg13g2_mux2_1 _2956_ (.A0(_0354_),
    .A1(_0441_),
    .S(net890),
    .X(_0442_));
 sg13g2_nand2_1 _2957_ (.Y(_0443_),
    .A(net882),
    .B(_0442_));
 sg13g2_a21oi_1 _2958_ (.A1(net1074),
    .A2(_0356_),
    .Y(_0444_),
    .B1(net873));
 sg13g2_nand2_1 _2959_ (.Y(_0445_),
    .A(\a[2] ),
    .B(_0360_));
 sg13g2_o21ai_1 _2960_ (.B1(net1093),
    .Y(_0446_),
    .A1(\a[1] ),
    .A2(\a[2] ));
 sg13g2_a21oi_1 _2961_ (.A1(\a[0] ),
    .A2(net868),
    .Y(_0447_),
    .B1(net1106));
 sg13g2_mux2_1 _2962_ (.A0(_1576_),
    .A1(_0446_),
    .S(_0445_),
    .X(_0448_));
 sg13g2_a22oi_1 _2963_ (.Y(_0449_),
    .B1(net850),
    .B2(net1068),
    .A2(net862),
    .A1(net1085));
 sg13g2_nand3_1 _2964_ (.B(_0448_),
    .C(_0449_),
    .A(_0447_),
    .Y(_0450_));
 sg13g2_a221oi_1 _2965_ (.B2(_0444_),
    .C1(_0450_),
    .B1(_0443_),
    .A1(\a[1] ),
    .Y(_0451_),
    .A2(net859));
 sg13g2_nand3_1 _2966_ (.B(_0136_),
    .C(_0137_),
    .A(net1034),
    .Y(_0452_));
 sg13g2_nand3_1 _2967_ (.B(_1545_),
    .C(_1546_),
    .A(net923),
    .Y(_0453_));
 sg13g2_nand3_1 _2968_ (.B(_0452_),
    .C(_0453_),
    .A(net918),
    .Y(_0454_));
 sg13g2_nand3_1 _2969_ (.B(_0138_),
    .C(_0139_),
    .A(net1042),
    .Y(_0455_));
 sg13g2_nand3_1 _2970_ (.B(_0140_),
    .C(_0141_),
    .A(net1049),
    .Y(_0456_));
 sg13g2_nand3_1 _2971_ (.B(_0454_),
    .C(_0455_),
    .A(net912),
    .Y(_0457_));
 sg13g2_nand3_1 _2972_ (.B(_0456_),
    .C(_0457_),
    .A(net907),
    .Y(_0458_));
 sg13g2_nand3_1 _2973_ (.B(_0142_),
    .C(_0143_),
    .A(net1056),
    .Y(_0459_));
 sg13g2_nand3_1 _2974_ (.B(_0144_),
    .C(_0145_),
    .A(net1065),
    .Y(_0460_));
 sg13g2_nand3_1 _2975_ (.B(_0458_),
    .C(_0459_),
    .A(net900),
    .Y(_0461_));
 sg13g2_a21oi_1 _2976_ (.A1(_0162_),
    .A2(_0163_),
    .Y(_0462_),
    .B1(net895));
 sg13g2_a21oi_1 _2977_ (.A1(_0460_),
    .A2(_0461_),
    .Y(_0463_),
    .B1(net1072));
 sg13g2_o21ai_1 _2978_ (.B1(net885),
    .Y(_0464_),
    .A1(_0462_),
    .A2(_0463_));
 sg13g2_o21ai_1 _2979_ (.B1(net1073),
    .Y(_0465_),
    .A1(_0180_),
    .A2(_0181_));
 sg13g2_nand3_1 _2980_ (.B(_0464_),
    .C(_0465_),
    .A(net877),
    .Y(_0466_));
 sg13g2_nor2b_1 _2981_ (.A(_0037_),
    .B_N(_0308_),
    .Y(_0467_));
 sg13g2_nor2_1 _2982_ (.A(net1036),
    .B(_0467_),
    .Y(_0468_));
 sg13g2_a21oi_1 _2983_ (.A1(net1036),
    .A2(_0310_),
    .Y(_0469_),
    .B1(_0468_));
 sg13g2_mux2_1 _2984_ (.A0(_0312_),
    .A1(_0469_),
    .S(net908),
    .X(_0470_));
 sg13g2_and2_1 _2985_ (.A(net902),
    .B(_0470_),
    .X(_0471_));
 sg13g2_a21oi_1 _2986_ (.A1(net1052),
    .A2(_0314_),
    .Y(_0472_),
    .B1(_0471_));
 sg13g2_nand2_1 _2987_ (.Y(_0473_),
    .A(net898),
    .B(_0472_));
 sg13g2_o21ai_1 _2988_ (.B1(_0473_),
    .Y(_0474_),
    .A1(net896),
    .A2(_0316_));
 sg13g2_mux2_1 _2989_ (.A0(_0318_),
    .A1(_0474_),
    .S(net889),
    .X(_0475_));
 sg13g2_or2_1 _2990_ (.X(_0476_),
    .B(_0320_),
    .A(net883));
 sg13g2_a21oi_1 _2991_ (.A1(net883),
    .A2(_0475_),
    .Y(_0477_),
    .B1(net872));
 sg13g2_a22oi_1 _2992_ (.Y(_0478_),
    .B1(net862),
    .B2(\a[20] ),
    .A2(net867),
    .A1(\a[4] ));
 sg13g2_and2_1 _2993_ (.A(\a[10] ),
    .B(net855),
    .X(_0479_));
 sg13g2_o21ai_1 _2994_ (.B1(\a[9] ),
    .Y(_0480_),
    .A1(net859),
    .A2(_0479_));
 sg13g2_or2_1 _2995_ (.X(_0481_),
    .B(\a[10] ),
    .A(\a[9] ));
 sg13g2_a21oi_1 _2996_ (.A1(net1098),
    .A2(\a[10] ),
    .Y(_0482_),
    .B1(net1088));
 sg13g2_o21ai_1 _2997_ (.B1(_0481_),
    .Y(_0483_),
    .A1(_0326_),
    .A2(_0482_));
 sg13g2_nand4_1 _2998_ (.B(_0478_),
    .C(_0480_),
    .A(net1104),
    .Y(_0484_),
    .D(_0483_));
 sg13g2_a221oi_1 _2999_ (.B2(_0477_),
    .C1(_0484_),
    .B1(_0476_),
    .A1(net1013),
    .Y(_0485_),
    .A2(net850));
 sg13g2_a221oi_1 _3000_ (.B2(_0485_),
    .C1(net1103),
    .B1(_0466_),
    .A1(_0432_),
    .Y(_0486_),
    .A2(_0451_));
 sg13g2_a21o_2 _3001_ (.A2(_0417_),
    .A1(_0416_),
    .B1(_0486_),
    .X(uio_out[1]));
 sg13g2_o21ai_1 _3002_ (.B1(net874),
    .Y(_0487_),
    .A1(_1149_),
    .A2(_1150_));
 sg13g2_a21oi_1 _3003_ (.A1(\ayayayayayaya.b[29] ),
    .A2(net864),
    .Y(_0488_),
    .B1(net1095));
 sg13g2_a22oi_1 _3004_ (.Y(_0489_),
    .B1(net852),
    .B2(\ayayayayayaya.b[26] ),
    .A2(net870),
    .A1(net998));
 sg13g2_o21ai_1 _3005_ (.B1(_1578_),
    .Y(_0490_),
    .A1(\a[27] ),
    .A2(net1091));
 sg13g2_o21ai_1 _3006_ (.B1(_0374_),
    .Y(_0491_),
    .A1(net1092),
    .A2(_0371_));
 sg13g2_a22oi_1 _3007_ (.Y(_0492_),
    .B1(_0491_),
    .B2(\a[27] ),
    .A2(_0490_),
    .A1(\a[26] ));
 sg13g2_and4_1 _3008_ (.A(_0487_),
    .B(_0488_),
    .C(_0489_),
    .D(_0492_),
    .X(_0493_));
 sg13g2_nor3_2 _3009_ (.A(_0037_),
    .B(_0036_),
    .C(_1664_),
    .Y(_0494_));
 sg13g2_or2_1 _3010_ (.X(_0495_),
    .B(_0494_),
    .A(net1044));
 sg13g2_o21ai_1 _3011_ (.B1(net1044),
    .Y(_0496_),
    .A1(_0381_),
    .A2(_0382_));
 sg13g2_nand3_1 _3012_ (.B(_0495_),
    .C(_0496_),
    .A(net904),
    .Y(_0497_));
 sg13g2_nand3_1 _3013_ (.B(_0379_),
    .C(_0383_),
    .A(net1053),
    .Y(_0498_));
 sg13g2_nor3_1 _3014_ (.A(_1027_),
    .B(_0385_),
    .C(_0386_),
    .Y(_0499_));
 sg13g2_a21oi_1 _3015_ (.A1(_0495_),
    .A2(_0496_),
    .Y(_0500_),
    .B1(net1052));
 sg13g2_nor3_1 _3016_ (.A(net1060),
    .B(_0499_),
    .C(_0500_),
    .Y(_0501_));
 sg13g2_nor3_1 _3017_ (.A(net900),
    .B(_0384_),
    .C(_0387_),
    .Y(_0502_));
 sg13g2_nor3_1 _3018_ (.A(net895),
    .B(_0388_),
    .C(_0389_),
    .Y(_0503_));
 sg13g2_nor3_1 _3019_ (.A(net1066),
    .B(_0501_),
    .C(_0502_),
    .Y(_0504_));
 sg13g2_o21ai_1 _3020_ (.B1(net888),
    .Y(_0505_),
    .A1(_0503_),
    .A2(_0504_));
 sg13g2_o21ai_1 _3021_ (.B1(net1080),
    .Y(_0506_),
    .A1(_0390_),
    .A2(_0391_));
 sg13g2_nand3_1 _3022_ (.B(_0505_),
    .C(_0506_),
    .A(net880),
    .Y(_0507_));
 sg13g2_o21ai_1 _3023_ (.B1(net1078),
    .Y(_0508_),
    .A1(_0405_),
    .A2(_0406_));
 sg13g2_nor3_1 _3024_ (.A(net917),
    .B(_0395_),
    .C(_0396_),
    .Y(_0509_));
 sg13g2_nor3_1 _3025_ (.A(net1041),
    .B(_1700_),
    .C(_1701_),
    .Y(_0510_));
 sg13g2_nor3_1 _3026_ (.A(net1048),
    .B(_0509_),
    .C(_0510_),
    .Y(_0511_));
 sg13g2_nor3_1 _3027_ (.A(net911),
    .B(_0397_),
    .C(_0398_),
    .Y(_0512_));
 sg13g2_nor3_1 _3028_ (.A(net905),
    .B(_0399_),
    .C(_0400_),
    .Y(_0513_));
 sg13g2_nor3_1 _3029_ (.A(net1055),
    .B(_0511_),
    .C(_0512_),
    .Y(_0514_));
 sg13g2_nor3_1 _3030_ (.A(net1063),
    .B(_0513_),
    .C(_0514_),
    .Y(_0515_));
 sg13g2_nor3_1 _3031_ (.A(net899),
    .B(_0401_),
    .C(_0402_),
    .Y(_0516_));
 sg13g2_nor3_1 _3032_ (.A(net893),
    .B(_0403_),
    .C(_0404_),
    .Y(_0517_));
 sg13g2_nor3_1 _3033_ (.A(net1070),
    .B(_0515_),
    .C(_0516_),
    .Y(_0518_));
 sg13g2_o21ai_1 _3034_ (.B1(net886),
    .Y(_0519_),
    .A1(_0517_),
    .A2(_0518_));
 sg13g2_nand3_1 _3035_ (.B(_0508_),
    .C(_0519_),
    .A(net879),
    .Y(_0520_));
 sg13g2_nand3_1 _3036_ (.B(_1460_),
    .C(net875),
    .A(_1459_),
    .Y(_0521_));
 sg13g2_nand3_1 _3037_ (.B(\a[18] ),
    .C(\a[19] ),
    .A(net1102),
    .Y(_0522_));
 sg13g2_or2_1 _3038_ (.X(_0523_),
    .B(\a[19] ),
    .A(\a[18] ));
 sg13g2_nand3_1 _3039_ (.B(_0522_),
    .C(_0523_),
    .A(net1094),
    .Y(_0524_));
 sg13g2_nor2_1 _3040_ (.A(_1576_),
    .B(_0522_),
    .Y(_0525_));
 sg13g2_a21oi_1 _3041_ (.A1(net968),
    .A2(net866),
    .Y(_0526_),
    .B1(_0525_));
 sg13g2_a21o_1 _3042_ (.A2(net871),
    .A1(net1013),
    .B1(net1105),
    .X(_0527_));
 sg13g2_a221oi_1 _3043_ (.B2(\ayayayayayaya.b[18] ),
    .C1(_0527_),
    .B1(net854),
    .A1(\a[18] ),
    .Y(_0528_),
    .A2(net860));
 sg13g2_and4_1 _3044_ (.A(_0521_),
    .B(_0524_),
    .C(_0526_),
    .D(_0528_),
    .X(_0529_));
 sg13g2_a221oi_1 _3045_ (.B2(_0529_),
    .C1(net1097),
    .B1(_0520_),
    .A1(_0493_),
    .Y(_0530_),
    .A2(_0507_));
 sg13g2_o21ai_1 _3046_ (.B1(net1073),
    .Y(_0531_),
    .A1(_0462_),
    .A2(_0463_));
 sg13g2_nand3_1 _3047_ (.B(_1547_),
    .C(_1548_),
    .A(net916),
    .Y(_0532_));
 sg13g2_nand3_1 _3048_ (.B(_0452_),
    .C(_0453_),
    .A(net1042),
    .Y(_0533_));
 sg13g2_nand3_1 _3049_ (.B(_0454_),
    .C(_0455_),
    .A(net1049),
    .Y(_0534_));
 sg13g2_nand3_1 _3050_ (.B(_0532_),
    .C(_0533_),
    .A(net912),
    .Y(_0535_));
 sg13g2_nand3_1 _3051_ (.B(_0534_),
    .C(_0535_),
    .A(net907),
    .Y(_0536_));
 sg13g2_nand3_1 _3052_ (.B(_0456_),
    .C(_0457_),
    .A(net1056),
    .Y(_0537_));
 sg13g2_nand3_1 _3053_ (.B(_0458_),
    .C(_0459_),
    .A(net1065),
    .Y(_0538_));
 sg13g2_nand3_1 _3054_ (.B(_0536_),
    .C(_0537_),
    .A(net900),
    .Y(_0539_));
 sg13g2_a21oi_1 _3055_ (.A1(_0460_),
    .A2(_0461_),
    .Y(_0540_),
    .B1(net895));
 sg13g2_a21oi_1 _3056_ (.A1(_0538_),
    .A2(_0539_),
    .Y(_0541_),
    .B1(net1072));
 sg13g2_o21ai_1 _3057_ (.B1(net888),
    .Y(_0542_),
    .A1(_0540_),
    .A2(_0541_));
 sg13g2_nand3_1 _3058_ (.B(_0531_),
    .C(_0542_),
    .A(net877),
    .Y(_0543_));
 sg13g2_nor2b_1 _3059_ (.A(_0036_),
    .B_N(_0467_),
    .Y(_0544_));
 sg13g2_and2_1 _3060_ (.A(net908),
    .B(_0544_),
    .X(_0545_));
 sg13g2_a21oi_1 _3061_ (.A1(net1043),
    .A2(_0469_),
    .Y(_0546_),
    .B1(_0545_));
 sg13g2_nor2_1 _3062_ (.A(net1052),
    .B(_0546_),
    .Y(_0547_));
 sg13g2_a21oi_1 _3063_ (.A1(net1052),
    .A2(_0470_),
    .Y(_0548_),
    .B1(_0547_));
 sg13g2_mux2_1 _3064_ (.A0(_0472_),
    .A1(_0548_),
    .S(net898),
    .X(_0549_));
 sg13g2_mux2_1 _3065_ (.A0(_0474_),
    .A1(_0549_),
    .S(net889),
    .X(_0550_));
 sg13g2_nand2_1 _3066_ (.Y(_0551_),
    .A(net883),
    .B(_0550_));
 sg13g2_a21oi_1 _3067_ (.A1(net1075),
    .A2(_0475_),
    .Y(_0552_),
    .B1(net872));
 sg13g2_o21ai_1 _3068_ (.B1(\a[11] ),
    .Y(_0553_),
    .A1(_0479_),
    .A2(_0482_));
 sg13g2_o21ai_1 _3069_ (.B1(net858),
    .Y(_0554_),
    .A1(\a[11] ),
    .A2(net1088));
 sg13g2_a22oi_1 _3070_ (.Y(_0555_),
    .B1(net854),
    .B2(net1008),
    .A2(net866),
    .A1(net976));
 sg13g2_a22oi_1 _3071_ (.Y(_0556_),
    .B1(_0554_),
    .B2(\a[10] ),
    .A2(net867),
    .A1(net1039));
 sg13g2_a21oi_1 _3072_ (.A1(_0551_),
    .A2(_0552_),
    .Y(_0557_),
    .B1(net1096));
 sg13g2_and4_1 _3073_ (.A(_0553_),
    .B(_0555_),
    .C(_0556_),
    .D(_0557_),
    .X(_0558_));
 sg13g2_nand3_1 _3074_ (.B(_0187_),
    .C(_0188_),
    .A(net915),
    .Y(_0559_));
 sg13g2_nand3_1 _3075_ (.B(_0418_),
    .C(_0419_),
    .A(net1037),
    .Y(_0560_));
 sg13g2_nand3_1 _3076_ (.B(_0420_),
    .C(_0421_),
    .A(net1044),
    .Y(_0561_));
 sg13g2_nand3_1 _3077_ (.B(_0559_),
    .C(_0560_),
    .A(net909),
    .Y(_0562_));
 sg13g2_nand3_1 _3078_ (.B(_0561_),
    .C(_0562_),
    .A(net904),
    .Y(_0563_));
 sg13g2_nand3_1 _3079_ (.B(_0422_),
    .C(_0423_),
    .A(net1053),
    .Y(_0564_));
 sg13g2_nand3_1 _3080_ (.B(_0424_),
    .C(_0425_),
    .A(net1061),
    .Y(_0565_));
 sg13g2_nand3_1 _3081_ (.B(_0563_),
    .C(_0564_),
    .A(net896),
    .Y(_0566_));
 sg13g2_a21oi_1 _3082_ (.A1(_0426_),
    .A2(_0427_),
    .Y(_0567_),
    .B1(net889));
 sg13g2_a21oi_1 _3083_ (.A1(_0565_),
    .A2(_0566_),
    .Y(_0568_),
    .B1(net1066));
 sg13g2_o21ai_1 _3084_ (.B1(net882),
    .Y(_0569_),
    .A1(_0567_),
    .A2(_0568_));
 sg13g2_o21ai_1 _3085_ (.B1(net1074),
    .Y(_0570_),
    .A1(_0428_),
    .A2(_0429_));
 sg13g2_nand3_1 _3086_ (.B(_0569_),
    .C(_0570_),
    .A(net878),
    .Y(_0571_));
 sg13g2_nand2_1 _3087_ (.Y(_0572_),
    .A(net1077),
    .B(_0442_));
 sg13g2_nand2_1 _3088_ (.Y(_0573_),
    .A(net1044),
    .B(_0437_));
 sg13g2_nand2_1 _3089_ (.Y(_0574_),
    .A(net1037),
    .B(_0435_));
 sg13g2_o21ai_1 _3090_ (.B1(_0574_),
    .Y(_0575_),
    .A1(net1037),
    .A2(_0298_));
 sg13g2_o21ai_1 _3091_ (.B1(_0573_),
    .Y(_0576_),
    .A1(net1044),
    .A2(_0575_));
 sg13g2_nor2_1 _3092_ (.A(net1051),
    .B(_0576_),
    .Y(_0577_));
 sg13g2_a21oi_1 _3093_ (.A1(net1051),
    .A2(_0439_),
    .Y(_0578_),
    .B1(_0577_));
 sg13g2_nor2_1 _3094_ (.A(net1061),
    .B(_0578_),
    .Y(_0579_));
 sg13g2_a21oi_1 _3095_ (.A1(net1061),
    .A2(_0440_),
    .Y(_0580_),
    .B1(_0579_));
 sg13g2_mux2_1 _3096_ (.A0(_0441_),
    .A1(_0580_),
    .S(net890),
    .X(_0581_));
 sg13g2_a21oi_1 _3097_ (.A1(net884),
    .A2(_0581_),
    .Y(_0582_),
    .B1(net872));
 sg13g2_a22oi_1 _3098_ (.Y(_0583_),
    .B1(net850),
    .B2(net1062),
    .A2(net867),
    .A1(net1068));
 sg13g2_and2_1 _3099_ (.A(\a[3] ),
    .B(net855),
    .X(_0584_));
 sg13g2_o21ai_1 _3100_ (.B1(\a[2] ),
    .Y(_0585_),
    .A1(net859),
    .A2(_0584_));
 sg13g2_nand3_1 _3101_ (.B(\a[2] ),
    .C(\a[3] ),
    .A(net1099),
    .Y(_0586_));
 sg13g2_or2_1 _3102_ (.X(_0587_),
    .B(\a[3] ),
    .A(\a[2] ));
 sg13g2_nand3_1 _3103_ (.B(_0586_),
    .C(_0587_),
    .A(net1093),
    .Y(_0588_));
 sg13g2_a21oi_1 _3104_ (.A1(\ayayayayayaya.b[17] ),
    .A2(net862),
    .Y(_0589_),
    .B1(net1104));
 sg13g2_nand4_1 _3105_ (.B(_0585_),
    .C(_0588_),
    .A(_0583_),
    .Y(_0590_),
    .D(_0589_));
 sg13g2_a21oi_1 _3106_ (.A1(_0572_),
    .A2(_0582_),
    .Y(_0591_),
    .B1(_0590_));
 sg13g2_a22oi_1 _3107_ (.Y(_0592_),
    .B1(_0571_),
    .B2(_0591_),
    .A2(_0558_),
    .A1(_0543_));
 sg13g2_a21o_2 _3108_ (.A2(_0592_),
    .A1(net1097),
    .B1(_0530_),
    .X(uio_out[2]));
 sg13g2_nand3_1 _3109_ (.B(_1406_),
    .C(net875),
    .A(_1405_),
    .Y(_0593_));
 sg13g2_and3_1 _3110_ (.X(_0594_),
    .A(net1100),
    .B(\a[19] ),
    .C(\a[20] ));
 sg13g2_nor2_1 _3111_ (.A(\a[19] ),
    .B(\a[20] ),
    .Y(_0595_));
 sg13g2_nor2_1 _3112_ (.A(_0594_),
    .B(_0595_),
    .Y(_0596_));
 sg13g2_a22oi_1 _3113_ (.Y(_0597_),
    .B1(_0594_),
    .B2(net1087),
    .A2(net851),
    .A1(\ayayayayayaya.b[19] ));
 sg13g2_a22oi_1 _3114_ (.Y(_0598_),
    .B1(net861),
    .B2(\a[19] ),
    .A2(net869),
    .A1(\a[9] ));
 sg13g2_a221oi_1 _3115_ (.B2(_0596_),
    .C1(net1105),
    .B1(net1094),
    .A1(\a[25] ),
    .Y(_0599_),
    .A2(net866));
 sg13g2_and4_1 _3116_ (.A(_0593_),
    .B(_0597_),
    .C(_0598_),
    .D(_0599_),
    .X(_0600_));
 sg13g2_nor3_1 _3117_ (.A(net1048),
    .B(_1702_),
    .C(_1703_),
    .Y(_0601_));
 sg13g2_nor3_1 _3118_ (.A(net911),
    .B(_0509_),
    .C(_0510_),
    .Y(_0602_));
 sg13g2_nor3_1 _3119_ (.A(net906),
    .B(_0511_),
    .C(_0512_),
    .Y(_0603_));
 sg13g2_nor3_1 _3120_ (.A(net1057),
    .B(_0601_),
    .C(_0602_),
    .Y(_0604_));
 sg13g2_nor3_1 _3121_ (.A(net1064),
    .B(_0603_),
    .C(_0604_),
    .Y(_0605_));
 sg13g2_nor3_1 _3122_ (.A(net901),
    .B(_0513_),
    .C(_0514_),
    .Y(_0606_));
 sg13g2_nor3_1 _3123_ (.A(net893),
    .B(_0515_),
    .C(_0516_),
    .Y(_0607_));
 sg13g2_nor3_1 _3124_ (.A(net1070),
    .B(_0605_),
    .C(_0606_),
    .Y(_0608_));
 sg13g2_o21ai_1 _3125_ (.B1(net886),
    .Y(_0609_),
    .A1(_0607_),
    .A2(_0608_));
 sg13g2_o21ai_1 _3126_ (.B1(net1078),
    .Y(_0610_),
    .A1(_0517_),
    .A2(_0518_));
 sg13g2_nand3_1 _3127_ (.B(_0609_),
    .C(_0610_),
    .A(net879),
    .Y(_0611_));
 sg13g2_nand3_1 _3128_ (.B(_0497_),
    .C(_0498_),
    .A(net1060),
    .Y(_0612_));
 sg13g2_nand2b_1 _3129_ (.Y(_0613_),
    .B(_0494_),
    .A_N(_0035_));
 sg13g2_nand2b_1 _3130_ (.Y(_0614_),
    .B(net902),
    .A_N(_0613_));
 sg13g2_nand3_1 _3131_ (.B(_0495_),
    .C(_0496_),
    .A(net1052),
    .Y(_0615_));
 sg13g2_nand3_1 _3132_ (.B(_0614_),
    .C(_0615_),
    .A(net898),
    .Y(_0616_));
 sg13g2_nor3_1 _3133_ (.A(net892),
    .B(_0501_),
    .C(_0502_),
    .Y(_0617_));
 sg13g2_a21oi_1 _3134_ (.A1(_0614_),
    .A2(_0615_),
    .Y(_0618_),
    .B1(net1059));
 sg13g2_nor3_1 _3135_ (.A(net898),
    .B(_0499_),
    .C(_0500_),
    .Y(_0619_));
 sg13g2_nor3_1 _3136_ (.A(net1066),
    .B(_0618_),
    .C(_0619_),
    .Y(_0620_));
 sg13g2_o21ai_1 _3137_ (.B1(net885),
    .Y(_0621_),
    .A1(_0617_),
    .A2(_0620_));
 sg13g2_o21ai_1 _3138_ (.B1(net1080),
    .Y(_0622_),
    .A1(_0503_),
    .A2(_0504_));
 sg13g2_nand3_1 _3139_ (.B(_0621_),
    .C(_0622_),
    .A(net880),
    .Y(_0623_));
 sg13g2_a21oi_1 _3140_ (.A1(\ayayayayayaya.b[27] ),
    .A2(net853),
    .Y(_0624_),
    .B1(net1095));
 sg13g2_a22oi_1 _3141_ (.Y(_0625_),
    .B1(net866),
    .B2(\a[29] ),
    .A2(net871),
    .A1(\a[13] ));
 sg13g2_and2_1 _3142_ (.A(net1102),
    .B(\a[28] ),
    .X(_0626_));
 sg13g2_a21oi_1 _3143_ (.A1(\a[27] ),
    .A2(_0626_),
    .Y(_0627_),
    .B1(net1092));
 sg13g2_o21ai_1 _3144_ (.B1(_0627_),
    .Y(_0628_),
    .A1(\a[27] ),
    .A2(\a[28] ));
 sg13g2_nand2_1 _3145_ (.Y(_0629_),
    .A(net1087),
    .B(_0626_));
 sg13g2_nand2_1 _3146_ (.Y(_0630_),
    .A(net857),
    .B(_0629_));
 sg13g2_nand3_1 _3147_ (.B(_0625_),
    .C(_0628_),
    .A(_0624_),
    .Y(_0631_));
 sg13g2_a221oi_1 _3148_ (.B2(\a[27] ),
    .C1(_0631_),
    .B1(_0630_),
    .A1(_1183_),
    .Y(_0632_),
    .A2(net876));
 sg13g2_a221oi_1 _3149_ (.B2(_0632_),
    .C1(net1097),
    .B1(_0623_),
    .A1(_0600_),
    .Y(_0633_),
    .A2(_0611_));
 sg13g2_o21ai_1 _3150_ (.B1(net1074),
    .Y(_0634_),
    .A1(_0567_),
    .A2(_0568_));
 sg13g2_nand3_1 _3151_ (.B(_0559_),
    .C(_0560_),
    .A(net1044),
    .Y(_0635_));
 sg13g2_nand3_1 _3152_ (.B(_0189_),
    .C(_0190_),
    .A(net909),
    .Y(_0636_));
 sg13g2_nand3_1 _3153_ (.B(_0635_),
    .C(_0636_),
    .A(net904),
    .Y(_0637_));
 sg13g2_nand3_1 _3154_ (.B(_0561_),
    .C(_0562_),
    .A(net1051),
    .Y(_0638_));
 sg13g2_nand3_1 _3155_ (.B(_0563_),
    .C(_0564_),
    .A(net1059),
    .Y(_0639_));
 sg13g2_nand3_1 _3156_ (.B(_0637_),
    .C(_0638_),
    .A(net897),
    .Y(_0640_));
 sg13g2_a21oi_1 _3157_ (.A1(_0565_),
    .A2(_0566_),
    .Y(_0641_),
    .B1(net889));
 sg13g2_a21oi_1 _3158_ (.A1(_0639_),
    .A2(_0640_),
    .Y(_0642_),
    .B1(net1066));
 sg13g2_o21ai_1 _3159_ (.B1(net883),
    .Y(_0643_),
    .A1(_0641_),
    .A2(_0642_));
 sg13g2_nand3_1 _3160_ (.B(_0634_),
    .C(_0643_),
    .A(net877),
    .Y(_0644_));
 sg13g2_or2_1 _3161_ (.X(_0645_),
    .B(_0575_),
    .A(net908));
 sg13g2_o21ai_1 _3162_ (.B1(_0645_),
    .Y(_0646_),
    .A1(net1045),
    .A2(_0300_));
 sg13g2_mux2_1 _3163_ (.A0(_0576_),
    .A1(_0646_),
    .S(net903),
    .X(_0647_));
 sg13g2_mux2_1 _3164_ (.A0(_0578_),
    .A1(_0647_),
    .S(net896),
    .X(_0648_));
 sg13g2_mux2_1 _3165_ (.A0(_0580_),
    .A1(_0648_),
    .S(net890),
    .X(_0649_));
 sg13g2_nand2_1 _3166_ (.Y(_0650_),
    .A(net884),
    .B(_0649_));
 sg13g2_a21oi_1 _3167_ (.A1(net1074),
    .A2(_0581_),
    .Y(_0651_),
    .B1(net872));
 sg13g2_a21oi_1 _3168_ (.A1(net1098),
    .A2(\a[3] ),
    .Y(_0652_),
    .B1(net1089));
 sg13g2_o21ai_1 _3169_ (.B1(\a[4] ),
    .Y(_0653_),
    .A1(_0584_),
    .A2(_0652_));
 sg13g2_nor2_1 _3170_ (.A(\a[4] ),
    .B(net1088),
    .Y(_0654_));
 sg13g2_o21ai_1 _3171_ (.B1(\a[3] ),
    .Y(_0655_),
    .A1(net859),
    .A2(_0654_));
 sg13g2_a22oi_1 _3172_ (.Y(_0656_),
    .B1(net862),
    .B2(\a[17] ),
    .A2(net867),
    .A1(\a[1] ));
 sg13g2_nand4_1 _3173_ (.B(_0653_),
    .C(_0655_),
    .A(net1096),
    .Y(_0657_),
    .D(_0656_));
 sg13g2_a221oi_1 _3174_ (.B2(_0651_),
    .C1(_0657_),
    .B1(_0650_),
    .A1(net1054),
    .Y(_0658_),
    .A2(net850));
 sg13g2_o21ai_1 _3175_ (.B1(net1080),
    .Y(_0659_),
    .A1(_0540_),
    .A2(_0541_));
 sg13g2_nand3_1 _3176_ (.B(_0532_),
    .C(_0533_),
    .A(net1047),
    .Y(_0660_));
 sg13g2_nand3_1 _3177_ (.B(_1549_),
    .C(_1550_),
    .A(net910),
    .Y(_0661_));
 sg13g2_nand3_1 _3178_ (.B(_0660_),
    .C(_0661_),
    .A(net905),
    .Y(_0662_));
 sg13g2_nand3_1 _3179_ (.B(_0534_),
    .C(_0535_),
    .A(net1056),
    .Y(_0663_));
 sg13g2_nand3_1 _3180_ (.B(_0536_),
    .C(_0537_),
    .A(net1065),
    .Y(_0664_));
 sg13g2_nand3_1 _3181_ (.B(_0662_),
    .C(_0663_),
    .A(net899),
    .Y(_0665_));
 sg13g2_a21oi_1 _3182_ (.A1(_0538_),
    .A2(_0539_),
    .Y(_0666_),
    .B1(net895));
 sg13g2_a21oi_1 _3183_ (.A1(_0664_),
    .A2(_0665_),
    .Y(_0667_),
    .B1(net1072));
 sg13g2_o21ai_1 _3184_ (.B1(net888),
    .Y(_0668_),
    .A1(_0666_),
    .A2(_0667_));
 sg13g2_nand3_1 _3185_ (.B(_0659_),
    .C(_0668_),
    .A(net880),
    .Y(_0669_));
 sg13g2_nand2_1 _3186_ (.Y(_0670_),
    .A(net1075),
    .B(_0550_));
 sg13g2_nand2b_1 _3187_ (.Y(_0671_),
    .B(_0544_),
    .A_N(_0035_));
 sg13g2_nand2b_1 _3188_ (.Y(_0672_),
    .B(net902),
    .A_N(_0671_));
 sg13g2_o21ai_1 _3189_ (.B1(_0672_),
    .Y(_0673_),
    .A1(net902),
    .A2(_0546_));
 sg13g2_nor2_1 _3190_ (.A(net1058),
    .B(_0673_),
    .Y(_0674_));
 sg13g2_a21oi_2 _3191_ (.B1(_0674_),
    .Y(_0675_),
    .A2(_0548_),
    .A1(net1058));
 sg13g2_nor2_1 _3192_ (.A(net889),
    .B(_0549_),
    .Y(_0676_));
 sg13g2_a21oi_2 _3193_ (.B1(_0676_),
    .Y(_0677_),
    .A2(_0675_),
    .A1(net891));
 sg13g2_a21oi_1 _3194_ (.A1(net883),
    .A2(_0677_),
    .Y(_0678_),
    .B1(net873));
 sg13g2_and2_1 _3195_ (.A(\a[12] ),
    .B(net855),
    .X(_0679_));
 sg13g2_a21oi_1 _3196_ (.A1(net1101),
    .A2(\a[12] ),
    .Y(_0680_),
    .B1(net1090));
 sg13g2_nand3_1 _3197_ (.B(\a[11] ),
    .C(\a[12] ),
    .A(net1101),
    .Y(_0681_));
 sg13g2_o21ai_1 _3198_ (.B1(_0681_),
    .Y(_0682_),
    .A1(\a[11] ),
    .A2(\a[12] ));
 sg13g2_nor2_1 _3199_ (.A(net1090),
    .B(_0682_),
    .Y(_0683_));
 sg13g2_a22oi_1 _3200_ (.Y(_0684_),
    .B1(_0679_),
    .B2(\a[11] ),
    .A2(net864),
    .A1(\a[21] ));
 sg13g2_a22oi_1 _3201_ (.Y(_0685_),
    .B1(net860),
    .B2(\a[11] ),
    .A2(net871),
    .A1(\a[5] ));
 sg13g2_a21oi_1 _3202_ (.A1(net1006),
    .A2(net852),
    .Y(_0686_),
    .B1(_0683_));
 sg13g2_nand4_1 _3203_ (.B(_0684_),
    .C(_0685_),
    .A(net1105),
    .Y(_0687_),
    .D(_0686_));
 sg13g2_a21oi_1 _3204_ (.A1(_0670_),
    .A2(_0678_),
    .Y(_0688_),
    .B1(_0687_));
 sg13g2_a22oi_1 _3205_ (.Y(_0689_),
    .B1(_0669_),
    .B2(_0688_),
    .A2(_0658_),
    .A1(_0644_));
 sg13g2_a21o_2 _3206_ (.A2(_0689_),
    .A1(net1097),
    .B1(_0633_),
    .X(uio_out[3]));
 sg13g2_o21ai_1 _3207_ (.B1(net874),
    .Y(_0690_),
    .A1(_1354_),
    .A2(_1355_));
 sg13g2_nand3_1 _3208_ (.B(\a[20] ),
    .C(\a[21] ),
    .A(net1101),
    .Y(_0691_));
 sg13g2_o21ai_1 _3209_ (.B1(_0691_),
    .Y(_0692_),
    .A1(\a[20] ),
    .A2(\a[21] ));
 sg13g2_nor2_1 _3210_ (.A(net1090),
    .B(_0692_),
    .Y(_0693_));
 sg13g2_a221oi_1 _3211_ (.B2(\ayayayayayaya.b[20] ),
    .C1(_0693_),
    .B1(net852),
    .A1(\ayayayayayaya.b[26] ),
    .Y(_0694_),
    .A2(net864));
 sg13g2_and2_1 _3212_ (.A(\a[21] ),
    .B(net856),
    .X(_0695_));
 sg13g2_o21ai_1 _3213_ (.B1(\a[20] ),
    .Y(_0696_),
    .A1(net861),
    .A2(_0695_));
 sg13g2_a21oi_1 _3214_ (.A1(net1008),
    .A2(net870),
    .Y(_0697_),
    .B1(net1105));
 sg13g2_and4_1 _3215_ (.A(_0690_),
    .B(_0694_),
    .C(_0696_),
    .D(_0697_),
    .X(_0698_));
 sg13g2_o21ai_1 _3216_ (.B1(net1078),
    .Y(_0699_),
    .A1(_0607_),
    .A2(_0608_));
 sg13g2_nor3_1 _3217_ (.A(net906),
    .B(_0601_),
    .C(_0602_),
    .Y(_0700_));
 sg13g2_nor3_1 _3218_ (.A(net1055),
    .B(_1704_),
    .C(_1705_),
    .Y(_0701_));
 sg13g2_nor3_1 _3219_ (.A(net1064),
    .B(_0700_),
    .C(_0701_),
    .Y(_0702_));
 sg13g2_nor3_1 _3220_ (.A(net900),
    .B(_0603_),
    .C(_0604_),
    .Y(_0703_));
 sg13g2_nor3_1 _3221_ (.A(net894),
    .B(_0605_),
    .C(_0606_),
    .Y(_0704_));
 sg13g2_nor3_1 _3222_ (.A(net1071),
    .B(_0702_),
    .C(_0703_),
    .Y(_0705_));
 sg13g2_o21ai_1 _3223_ (.B1(net887),
    .Y(_0706_),
    .A1(_0704_),
    .A2(_0705_));
 sg13g2_nand3_1 _3224_ (.B(_0699_),
    .C(_0706_),
    .A(net880),
    .Y(_0707_));
 sg13g2_nor3_1 _3225_ (.A(net1058),
    .B(_0034_),
    .C(_0613_),
    .Y(_0708_));
 sg13g2_a21oi_1 _3226_ (.A1(_0614_),
    .A2(_0615_),
    .Y(_0709_),
    .B1(net898));
 sg13g2_o21ai_1 _3227_ (.B1(net892),
    .Y(_0710_),
    .A1(_0708_),
    .A2(_0709_));
 sg13g2_nand3_1 _3228_ (.B(_0612_),
    .C(_0616_),
    .A(net1066),
    .Y(_0711_));
 sg13g2_nand3_1 _3229_ (.B(_0710_),
    .C(_0711_),
    .A(net885),
    .Y(_0712_));
 sg13g2_o21ai_1 _3230_ (.B1(net1073),
    .Y(_0713_),
    .A1(_0617_),
    .A2(_0620_));
 sg13g2_nand3_1 _3231_ (.B(_0712_),
    .C(_0713_),
    .A(net877),
    .Y(_0714_));
 sg13g2_o21ai_1 _3232_ (.B1(net874),
    .Y(_0715_),
    .A1(_1217_),
    .A2(_1218_));
 sg13g2_a21oi_1 _3233_ (.A1(\ayayayayayaya.b[30] ),
    .A2(net866),
    .Y(_0716_),
    .B1(net1095));
 sg13g2_a22oi_1 _3234_ (.Y(_0717_),
    .B1(net852),
    .B2(\ayayayayayaya.b[28] ),
    .A2(net870),
    .A1(net994));
 sg13g2_nor2_1 _3235_ (.A(\a[29] ),
    .B(net1092),
    .Y(_0718_));
 sg13g2_or2_1 _3236_ (.X(_0719_),
    .B(_0718_),
    .A(net860));
 sg13g2_o21ai_1 _3237_ (.B1(_0629_),
    .Y(_0720_),
    .A1(net1092),
    .A2(_0626_));
 sg13g2_a22oi_1 _3238_ (.Y(_0721_),
    .B1(_0720_),
    .B2(\a[29] ),
    .A2(_0719_),
    .A1(\a[28] ));
 sg13g2_and4_1 _3239_ (.A(_0715_),
    .B(_0716_),
    .C(_0717_),
    .D(_0721_),
    .X(_0722_));
 sg13g2_a22oi_1 _3240_ (.Y(_0723_),
    .B1(_0714_),
    .B2(_0722_),
    .A2(_0707_),
    .A1(_0698_));
 sg13g2_nand3_1 _3241_ (.B(_0191_),
    .C(_0192_),
    .A(net904),
    .Y(_0724_));
 sg13g2_nand3_1 _3242_ (.B(_0635_),
    .C(_0636_),
    .A(net1053),
    .Y(_0725_));
 sg13g2_nand3_1 _3243_ (.B(_0637_),
    .C(_0638_),
    .A(net1060),
    .Y(_0726_));
 sg13g2_nand3_1 _3244_ (.B(_0724_),
    .C(_0725_),
    .A(net898),
    .Y(_0727_));
 sg13g2_a21oi_1 _3245_ (.A1(_0639_),
    .A2(_0640_),
    .Y(_0728_),
    .B1(net892));
 sg13g2_a21oi_1 _3246_ (.A1(_0726_),
    .A2(_0727_),
    .Y(_0729_),
    .B1(net1066));
 sg13g2_o21ai_1 _3247_ (.B1(net885),
    .Y(_0730_),
    .A1(_0728_),
    .A2(_0729_));
 sg13g2_o21ai_1 _3248_ (.B1(net1073),
    .Y(_0731_),
    .A1(_0641_),
    .A2(_0642_));
 sg13g2_nand3_1 _3249_ (.B(_0730_),
    .C(_0731_),
    .A(net878),
    .Y(_0732_));
 sg13g2_nor2_1 _3250_ (.A(net903),
    .B(_0646_),
    .Y(_0733_));
 sg13g2_a21oi_1 _3251_ (.A1(net903),
    .A2(_0302_),
    .Y(_0734_),
    .B1(_0733_));
 sg13g2_mux2_1 _3252_ (.A0(_0647_),
    .A1(_0734_),
    .S(net896),
    .X(_0735_));
 sg13g2_mux2_1 _3253_ (.A0(_0648_),
    .A1(_0735_),
    .S(net889),
    .X(_0736_));
 sg13g2_nand2_1 _3254_ (.Y(_0737_),
    .A(net883),
    .B(_0736_));
 sg13g2_a21oi_1 _3255_ (.A1(net1075),
    .A2(_0649_),
    .Y(_0738_),
    .B1(net873));
 sg13g2_a22oi_1 _3256_ (.Y(_0739_),
    .B1(net862),
    .B2(\ayayayayayaya.b[18] ),
    .A2(net867),
    .A1(net1062));
 sg13g2_and2_1 _3257_ (.A(\a[5] ),
    .B(net855),
    .X(_0740_));
 sg13g2_o21ai_1 _3258_ (.B1(\a[4] ),
    .Y(_0741_),
    .A1(net859),
    .A2(_0740_));
 sg13g2_or2_1 _3259_ (.X(_0742_),
    .B(\a[5] ),
    .A(\a[4] ));
 sg13g2_a21oi_1 _3260_ (.A1(net1098),
    .A2(\a[5] ),
    .Y(_0743_),
    .B1(net1088));
 sg13g2_o21ai_1 _3261_ (.B1(_0742_),
    .Y(_0744_),
    .A1(_0654_),
    .A2(_0743_));
 sg13g2_nand4_1 _3262_ (.B(_0739_),
    .C(_0741_),
    .A(net1096),
    .Y(_0745_),
    .D(_0744_));
 sg13g2_a221oi_1 _3263_ (.B2(_0738_),
    .C1(_0745_),
    .B1(_0737_),
    .A1(net1046),
    .Y(_0746_),
    .A2(net850));
 sg13g2_o21ai_1 _3264_ (.B1(net1080),
    .Y(_0747_),
    .A1(_0666_),
    .A2(_0667_));
 sg13g2_nand3_1 _3265_ (.B(_1551_),
    .C(_1552_),
    .A(net905),
    .Y(_0748_));
 sg13g2_nand3_1 _3266_ (.B(_0660_),
    .C(_0661_),
    .A(net1055),
    .Y(_0749_));
 sg13g2_nand3_1 _3267_ (.B(_0662_),
    .C(_0663_),
    .A(net1063),
    .Y(_0750_));
 sg13g2_nand3_1 _3268_ (.B(_0748_),
    .C(_0749_),
    .A(net899),
    .Y(_0751_));
 sg13g2_a21oi_1 _3269_ (.A1(_0664_),
    .A2(_0665_),
    .Y(_0752_),
    .B1(net895));
 sg13g2_a21oi_1 _3270_ (.A1(_0750_),
    .A2(_0751_),
    .Y(_0753_),
    .B1(net1070));
 sg13g2_o21ai_1 _3271_ (.B1(net888),
    .Y(_0754_),
    .A1(_0752_),
    .A2(_0753_));
 sg13g2_nand3_1 _3272_ (.B(_0747_),
    .C(_0754_),
    .A(net880),
    .Y(_0755_));
 sg13g2_nor3_1 _3273_ (.A(net1058),
    .B(_0034_),
    .C(_0671_),
    .Y(_0756_));
 sg13g2_a21o_1 _3274_ (.A2(_0673_),
    .A1(net1058),
    .B1(_0756_),
    .X(_0757_));
 sg13g2_mux2_1 _3275_ (.A0(_0675_),
    .A1(_0757_),
    .S(net889),
    .X(_0758_));
 sg13g2_o21ai_1 _3276_ (.B1(net876),
    .Y(_0759_),
    .A1(net1075),
    .A2(_0758_));
 sg13g2_a21oi_1 _3277_ (.A1(net1076),
    .A2(_0677_),
    .Y(_0760_),
    .B1(_0759_));
 sg13g2_a21oi_1 _3278_ (.A1(net1002),
    .A2(net852),
    .Y(_0761_),
    .B1(_0999_));
 sg13g2_a22oi_1 _3279_ (.Y(_0762_),
    .B1(net864),
    .B2(net973),
    .A2(net870),
    .A1(net1035));
 sg13g2_o21ai_1 _3280_ (.B1(net857),
    .Y(_0763_),
    .A1(\a[13] ),
    .A2(net1090));
 sg13g2_a21o_1 _3281_ (.A2(net855),
    .A1(\a[12] ),
    .B1(_0680_),
    .X(_0764_));
 sg13g2_a22oi_1 _3282_ (.Y(_0765_),
    .B1(_0764_),
    .B2(\a[13] ),
    .A2(_0763_),
    .A1(\a[12] ));
 sg13g2_nand3_1 _3283_ (.B(_0762_),
    .C(_0765_),
    .A(_0761_),
    .Y(_0766_));
 sg13g2_nor2_1 _3284_ (.A(_0760_),
    .B(_0766_),
    .Y(_0767_));
 sg13g2_a221oi_1 _3285_ (.B2(_0767_),
    .C1(net1103),
    .B1(_0755_),
    .A1(_0732_),
    .Y(_0768_),
    .A2(_0746_));
 sg13g2_a21o_2 _3286_ (.A2(_0723_),
    .A1(net1),
    .B1(_0768_),
    .X(uio_out[4]));
 sg13g2_nand3_1 _3287_ (.B(_0748_),
    .C(_0749_),
    .A(net1063),
    .Y(_0769_));
 sg13g2_nand3_1 _3288_ (.B(_1553_),
    .C(_1554_),
    .A(net899),
    .Y(_0770_));
 sg13g2_a21oi_1 _3289_ (.A1(_0750_),
    .A2(_0751_),
    .Y(_0771_),
    .B1(net893));
 sg13g2_a21oi_1 _3290_ (.A1(_0769_),
    .A2(_0770_),
    .Y(_0772_),
    .B1(net1070));
 sg13g2_o21ai_1 _3291_ (.B1(net886),
    .Y(_0773_),
    .A1(_0771_),
    .A2(_0772_));
 sg13g2_o21ai_1 _3292_ (.B1(net1080),
    .Y(_0774_),
    .A1(_0752_),
    .A2(_0753_));
 sg13g2_nand3_1 _3293_ (.B(_0773_),
    .C(_0774_),
    .A(net880),
    .Y(_0775_));
 sg13g2_and2_1 _3294_ (.A(net1100),
    .B(\a[14] ),
    .X(_0776_));
 sg13g2_nand2_1 _3295_ (.Y(_0777_),
    .A(net1087),
    .B(_0776_));
 sg13g2_a21o_1 _3296_ (.A2(_0777_),
    .A1(net858),
    .B1(_1000_),
    .X(_0778_));
 sg13g2_a21oi_1 _3297_ (.A1(\a[13] ),
    .A2(_0776_),
    .Y(_0779_),
    .B1(net1089));
 sg13g2_o21ai_1 _3298_ (.B1(_0779_),
    .Y(_0780_),
    .A1(\a[13] ),
    .A2(\a[14] ));
 sg13g2_a22oi_1 _3299_ (.Y(_0781_),
    .B1(net863),
    .B2(\a[22] ),
    .A2(net869),
    .A1(\a[6] ));
 sg13g2_nand4_1 _3300_ (.B(_0778_),
    .C(_0780_),
    .A(net1104),
    .Y(_0782_),
    .D(_0781_));
 sg13g2_nor3_1 _3301_ (.A(_0034_),
    .B(_0033_),
    .C(_0671_),
    .Y(_0783_));
 sg13g2_inv_1 _3302_ (.Y(_0784_),
    .A(_0783_));
 sg13g2_nand2_1 _3303_ (.Y(_0785_),
    .A(net1067),
    .B(_0757_));
 sg13g2_o21ai_1 _3304_ (.B1(_0785_),
    .Y(_0786_),
    .A1(net1067),
    .A2(_0784_));
 sg13g2_mux2_1 _3305_ (.A0(_0758_),
    .A1(_0786_),
    .S(net882),
    .X(_0787_));
 sg13g2_a221oi_1 _3306_ (.B2(net876),
    .C1(_0782_),
    .B1(_0787_),
    .A1(net998),
    .Y(_0788_),
    .A2(net851));
 sg13g2_o21ai_1 _3307_ (.B1(net1073),
    .Y(_0789_),
    .A1(_0728_),
    .A2(_0729_));
 sg13g2_nand3_1 _3308_ (.B(_0724_),
    .C(_0725_),
    .A(net1060),
    .Y(_0790_));
 sg13g2_nand3_1 _3309_ (.B(_0193_),
    .C(_0194_),
    .A(net898),
    .Y(_0791_));
 sg13g2_a21oi_1 _3310_ (.A1(_0726_),
    .A2(_0727_),
    .Y(_0792_),
    .B1(net892));
 sg13g2_a21oi_1 _3311_ (.A1(_0790_),
    .A2(_0791_),
    .Y(_0793_),
    .B1(net1069));
 sg13g2_o21ai_1 _3312_ (.B1(net885),
    .Y(_0794_),
    .A1(_0792_),
    .A2(_0793_));
 sg13g2_nand3_1 _3313_ (.B(_0789_),
    .C(_0794_),
    .A(net877),
    .Y(_0795_));
 sg13g2_nand2_1 _3314_ (.Y(_0796_),
    .A(net1058),
    .B(_0734_));
 sg13g2_o21ai_1 _3315_ (.B1(_0796_),
    .Y(_0797_),
    .A1(net1058),
    .A2(_0304_));
 sg13g2_mux2_1 _3316_ (.A0(_0735_),
    .A1(_0797_),
    .S(net889),
    .X(_0798_));
 sg13g2_nand2_1 _3317_ (.Y(_0799_),
    .A(net883),
    .B(_0798_));
 sg13g2_a21oi_1 _3318_ (.A1(net1075),
    .A2(_0736_),
    .Y(_0800_),
    .B1(net873));
 sg13g2_o21ai_1 _3319_ (.B1(\a[6] ),
    .Y(_0801_),
    .A1(_0740_),
    .A2(_0743_));
 sg13g2_o21ai_1 _3320_ (.B1(net858),
    .Y(_0802_),
    .A1(\a[6] ),
    .A2(net1088));
 sg13g2_a22oi_1 _3321_ (.Y(_0803_),
    .B1(net851),
    .B2(net1039),
    .A2(net863),
    .A1(\a[18] ));
 sg13g2_a22oi_1 _3322_ (.Y(_0804_),
    .B1(_0802_),
    .B2(\a[5] ),
    .A2(net868),
    .A1(\a[2] ));
 sg13g2_nand4_1 _3323_ (.B(_0801_),
    .C(_0803_),
    .A(net1096),
    .Y(_0805_),
    .D(_0804_));
 sg13g2_a21oi_1 _3324_ (.A1(_0799_),
    .A2(_0800_),
    .Y(_0806_),
    .B1(_0805_));
 sg13g2_a22oi_1 _3325_ (.Y(_0807_),
    .B1(_0795_),
    .B2(_0806_),
    .A2(_0788_),
    .A1(_0775_));
 sg13g2_o21ai_1 _3326_ (.B1(net874),
    .Y(_0808_),
    .A1(_1255_),
    .A2(_1256_));
 sg13g2_o21ai_1 _3327_ (.B1(\a[30] ),
    .Y(_0809_),
    .A1(net866),
    .A2(_0718_));
 sg13g2_a221oi_1 _3328_ (.B2(\ayayayayayaya.b[29] ),
    .C1(net1095),
    .B1(net854),
    .A1(\a[14] ),
    .Y(_0810_),
    .A2(net871));
 sg13g2_nand2_1 _3329_ (.Y(_0811_),
    .A(net1100),
    .B(\a[30] ));
 sg13g2_nand2_1 _3330_ (.Y(_0812_),
    .A(net1094),
    .B(_0811_));
 sg13g2_o21ai_1 _3331_ (.B1(_0812_),
    .Y(_0813_),
    .A1(_1576_),
    .A2(_0811_));
 sg13g2_o21ai_1 _3332_ (.B1(\a[29] ),
    .Y(_0814_),
    .A1(net860),
    .A2(_0813_));
 sg13g2_and4_1 _3333_ (.A(_0808_),
    .B(_0809_),
    .C(_0810_),
    .D(_0814_),
    .X(_0815_));
 sg13g2_nand3_1 _3334_ (.B(_0710_),
    .C(_0711_),
    .A(net1073),
    .Y(_0816_));
 sg13g2_nor3_1 _3335_ (.A(_0034_),
    .B(_0033_),
    .C(_0613_),
    .Y(_0817_));
 sg13g2_inv_1 _3336_ (.Y(_0818_),
    .A(_0817_));
 sg13g2_nor2_1 _3337_ (.A(net1067),
    .B(_0817_),
    .Y(_0819_));
 sg13g2_nor3_1 _3338_ (.A(net892),
    .B(_0708_),
    .C(_0709_),
    .Y(_0820_));
 sg13g2_o21ai_1 _3339_ (.B1(net882),
    .Y(_0821_),
    .A1(_0819_),
    .A2(_0820_));
 sg13g2_nand3_1 _3340_ (.B(_0816_),
    .C(_0821_),
    .A(net878),
    .Y(_0822_));
 sg13g2_o21ai_1 _3341_ (.B1(net874),
    .Y(_0823_),
    .A1(_1326_),
    .A2(_1327_));
 sg13g2_a22oi_1 _3342_ (.Y(_0824_),
    .B1(net852),
    .B2(net976),
    .A2(net870),
    .A1(\a[10] ));
 sg13g2_a21oi_1 _3343_ (.A1(\a[26] ),
    .A2(net865),
    .Y(_0825_),
    .B1(net1105));
 sg13g2_nor2_1 _3344_ (.A(\a[22] ),
    .B(net1091),
    .Y(_0826_));
 sg13g2_o21ai_1 _3345_ (.B1(\a[21] ),
    .Y(_0827_),
    .A1(net860),
    .A2(_0826_));
 sg13g2_a21oi_1 _3346_ (.A1(net1101),
    .A2(\a[21] ),
    .Y(_0828_),
    .B1(net1090));
 sg13g2_o21ai_1 _3347_ (.B1(\a[22] ),
    .Y(_0829_),
    .A1(_0695_),
    .A2(_0828_));
 sg13g2_nand4_1 _3348_ (.B(_0825_),
    .C(_0827_),
    .A(_0824_),
    .Y(_0830_),
    .D(_0829_));
 sg13g2_nor2b_1 _3349_ (.A(_0830_),
    .B_N(_0823_),
    .Y(_0831_));
 sg13g2_nor3_1 _3350_ (.A(net1064),
    .B(_1706_),
    .C(_1707_),
    .Y(_0832_));
 sg13g2_nor3_1 _3351_ (.A(net901),
    .B(_0700_),
    .C(_0701_),
    .Y(_0833_));
 sg13g2_nor3_1 _3352_ (.A(net894),
    .B(_0702_),
    .C(_0703_),
    .Y(_0834_));
 sg13g2_nor3_1 _3353_ (.A(net1071),
    .B(_0832_),
    .C(_0833_),
    .Y(_0835_));
 sg13g2_o21ai_1 _3354_ (.B1(net887),
    .Y(_0836_),
    .A1(_0834_),
    .A2(_0835_));
 sg13g2_o21ai_1 _3355_ (.B1(net1079),
    .Y(_0837_),
    .A1(_0704_),
    .A2(_0705_));
 sg13g2_nand3_1 _3356_ (.B(_0836_),
    .C(_0837_),
    .A(net880),
    .Y(_0838_));
 sg13g2_a221oi_1 _3357_ (.B2(_0838_),
    .C1(net1097),
    .B1(_0831_),
    .A1(_0815_),
    .Y(_0839_),
    .A2(_0822_));
 sg13g2_a21o_2 _3358_ (.A2(_0807_),
    .A1(net1097),
    .B1(_0839_),
    .X(uio_out[5]));
 sg13g2_a21oi_1 _3359_ (.A1(_0769_),
    .A2(_0770_),
    .Y(_0840_),
    .B1(net893));
 sg13g2_a21oi_1 _3360_ (.A1(_1555_),
    .A2(_1556_),
    .Y(_0841_),
    .B1(net1070));
 sg13g2_o21ai_1 _3361_ (.B1(net886),
    .Y(_0842_),
    .A1(_0840_),
    .A2(_0841_));
 sg13g2_o21ai_1 _3362_ (.B1(net1078),
    .Y(_0843_),
    .A1(_0771_),
    .A2(_0772_));
 sg13g2_nand3_1 _3363_ (.B(_0842_),
    .C(_0843_),
    .A(net879),
    .Y(_0844_));
 sg13g2_nand2b_1 _3364_ (.Y(_0845_),
    .B(_0783_),
    .A_N(_0032_));
 sg13g2_a21oi_1 _3365_ (.A1(net882),
    .A2(_0845_),
    .Y(_0846_),
    .B1(net872));
 sg13g2_o21ai_1 _3366_ (.B1(_0846_),
    .Y(_0847_),
    .A1(net882),
    .A2(_0786_));
 sg13g2_and2_1 _3367_ (.A(net1025),
    .B(net869),
    .X(_0848_));
 sg13g2_o21ai_1 _3368_ (.B1(_0777_),
    .Y(_0849_),
    .A1(net1089),
    .A2(_0776_));
 sg13g2_o21ai_1 _3369_ (.B1(net858),
    .Y(_0850_),
    .A1(net1082),
    .A2(net1089));
 sg13g2_a221oi_1 _3370_ (.B2(net994),
    .C1(_0999_),
    .B1(net852),
    .A1(net971),
    .Y(_0851_),
    .A2(net864));
 sg13g2_a221oi_1 _3371_ (.B2(\a[14] ),
    .C1(_0848_),
    .B1(_0850_),
    .A1(net1082),
    .Y(_0852_),
    .A2(_0849_));
 sg13g2_nand4_1 _3372_ (.B(_0847_),
    .C(_0851_),
    .A(_0844_),
    .Y(_0853_),
    .D(_0852_));
 sg13g2_a21oi_1 _3373_ (.A1(_0790_),
    .A2(_0791_),
    .Y(_0854_),
    .B1(net892));
 sg13g2_a21oi_1 _3374_ (.A1(_0195_),
    .A2(_0196_),
    .Y(_0855_),
    .B1(net1069));
 sg13g2_o21ai_1 _3375_ (.B1(net885),
    .Y(_0856_),
    .A1(_0854_),
    .A2(_0855_));
 sg13g2_o21ai_1 _3376_ (.B1(net1073),
    .Y(_0857_),
    .A1(_0792_),
    .A2(_0793_));
 sg13g2_nand3_1 _3377_ (.B(_0856_),
    .C(_0857_),
    .A(net877),
    .Y(_0858_));
 sg13g2_nand2_1 _3378_ (.Y(_0859_),
    .A(net1075),
    .B(_0798_));
 sg13g2_nor2_1 _3379_ (.A(net890),
    .B(_0797_),
    .Y(_0860_));
 sg13g2_a21oi_2 _3380_ (.B1(_0860_),
    .Y(_0861_),
    .A2(_0306_),
    .A1(net891));
 sg13g2_a21oi_1 _3381_ (.A1(net883),
    .A2(_0861_),
    .Y(_0862_),
    .B1(net872));
 sg13g2_nand2_1 _3382_ (.Y(_0863_),
    .A(net1098),
    .B(\a[7] ));
 sg13g2_and3_1 _3383_ (.X(_0864_),
    .A(net1098),
    .B(\a[6] ),
    .C(\a[7] ));
 sg13g2_a221oi_1 _3384_ (.B2(net1035),
    .C1(_0864_),
    .B1(_1567_),
    .A1(\a[6] ),
    .Y(_0865_),
    .A2(_1565_));
 sg13g2_o21ai_1 _3385_ (.B1(net1093),
    .Y(_0866_),
    .A1(\a[6] ),
    .A2(\a[7] ));
 sg13g2_o21ai_1 _3386_ (.B1(net1096),
    .Y(_0867_),
    .A1(_0864_),
    .A2(_0866_));
 sg13g2_a221oi_1 _3387_ (.B2(\ayayayayayaya.b[19] ),
    .C1(_0867_),
    .B1(net862),
    .A1(net1054),
    .Y(_0868_),
    .A2(net868));
 sg13g2_o21ai_1 _3388_ (.B1(_0868_),
    .Y(_0869_),
    .A1(_1576_),
    .A2(_0865_));
 sg13g2_a21oi_1 _3389_ (.A1(_0859_),
    .A2(_0862_),
    .Y(_0870_),
    .B1(_0869_));
 sg13g2_a21oi_1 _3390_ (.A1(_0858_),
    .A2(_0870_),
    .Y(_0871_),
    .B1(net1103));
 sg13g2_o21ai_1 _3391_ (.B1(net874),
    .Y(_0872_),
    .A1(_1281_),
    .A2(_1282_));
 sg13g2_a22oi_1 _3392_ (.Y(_0873_),
    .B1(net864),
    .B2(\ayayayayayaya.b[27] ),
    .A2(net870),
    .A1(net1006));
 sg13g2_a21oi_1 _3393_ (.A1(net973),
    .A2(net853),
    .Y(_0874_),
    .B1(net1105));
 sg13g2_a21oi_1 _3394_ (.A1(net1101),
    .A2(\a[23] ),
    .Y(_0875_),
    .B1(net1091));
 sg13g2_or2_1 _3395_ (.X(_0876_),
    .B(_0875_),
    .A(net860));
 sg13g2_a21o_1 _3396_ (.A2(net856),
    .A1(\a[22] ),
    .B1(_0826_),
    .X(_0877_));
 sg13g2_a22oi_1 _3397_ (.Y(_0878_),
    .B1(_0877_),
    .B2(\a[23] ),
    .A2(_0876_),
    .A1(\a[22] ));
 sg13g2_and4_1 _3398_ (.A(_0872_),
    .B(_0873_),
    .C(_0874_),
    .D(_0878_),
    .X(_0879_));
 sg13g2_nor3_1 _3399_ (.A(net893),
    .B(_0832_),
    .C(_0833_),
    .Y(_0880_));
 sg13g2_nor3_1 _3400_ (.A(net1071),
    .B(_1708_),
    .C(_1709_),
    .Y(_0881_));
 sg13g2_o21ai_1 _3401_ (.B1(net887),
    .Y(_0882_),
    .A1(_0880_),
    .A2(_0881_));
 sg13g2_o21ai_1 _3402_ (.B1(net1079),
    .Y(_0883_),
    .A1(_0834_),
    .A2(_0835_));
 sg13g2_nand3_1 _3403_ (.B(_0882_),
    .C(_0883_),
    .A(net881),
    .Y(_0884_));
 sg13g2_o21ai_1 _3404_ (.B1(net875),
    .Y(_0885_),
    .A1(_1298_),
    .A2(_1299_));
 sg13g2_a21oi_1 _3405_ (.A1(\ayayayayayaya.b[30] ),
    .A2(net854),
    .Y(_0886_),
    .B1(net1095));
 sg13g2_a22oi_1 _3406_ (.Y(_0887_),
    .B1(net866),
    .B2(\ayayayayayaya.b[31] ),
    .A2(net871),
    .A1(net991));
 sg13g2_o21ai_1 _3407_ (.B1(net857),
    .Y(_0888_),
    .A1(\a[31] ),
    .A2(net1092));
 sg13g2_a22oi_1 _3408_ (.Y(_0889_),
    .B1(_0888_),
    .B2(\a[30] ),
    .A2(_0813_),
    .A1(\a[31] ));
 sg13g2_and4_1 _3409_ (.A(_0885_),
    .B(_0886_),
    .C(_0887_),
    .D(_0889_),
    .X(_0890_));
 sg13g2_o21ai_1 _3410_ (.B1(net1074),
    .Y(_0891_),
    .A1(_0819_),
    .A2(_0820_));
 sg13g2_o21ai_1 _3411_ (.B1(net882),
    .Y(_0892_),
    .A1(_0032_),
    .A2(_0818_));
 sg13g2_nand3_1 _3412_ (.B(_0891_),
    .C(_0892_),
    .A(net878),
    .Y(_0893_));
 sg13g2_a221oi_1 _3413_ (.B2(_0893_),
    .C1(net1097),
    .B1(_0890_),
    .A1(_0879_),
    .Y(_0894_),
    .A2(_0884_));
 sg13g2_a21o_2 _3414_ (.A2(_0871_),
    .A1(_0853_),
    .B1(_0894_),
    .X(uio_out[6]));
 sg13g2_o21ai_1 _3415_ (.B1(net874),
    .Y(_0895_),
    .A1(_1241_),
    .A2(_1242_));
 sg13g2_nand3_1 _3416_ (.B(\a[23] ),
    .C(\a[24] ),
    .A(net1101),
    .Y(_0896_));
 sg13g2_o21ai_1 _3417_ (.B1(_0896_),
    .Y(_0897_),
    .A1(\a[23] ),
    .A2(\a[24] ));
 sg13g2_nor2_1 _3418_ (.A(net1091),
    .B(_0897_),
    .Y(_0898_));
 sg13g2_a221oi_1 _3419_ (.B2(net971),
    .C1(_0898_),
    .B1(net853),
    .A1(\a[11] ),
    .Y(_0899_),
    .A2(net871));
 sg13g2_o21ai_1 _3420_ (.B1(\a[23] ),
    .Y(_0900_),
    .A1(net860),
    .A2(_1589_));
 sg13g2_a21oi_1 _3421_ (.A1(\a[27] ),
    .A2(net865),
    .Y(_0901_),
    .B1(net1106));
 sg13g2_and4_1 _3422_ (.A(_0895_),
    .B(_0899_),
    .C(_0900_),
    .D(_0901_),
    .X(_0902_));
 sg13g2_o21ai_1 _3423_ (.B1(net887),
    .Y(_0903_),
    .A1(_1710_),
    .A2(_1711_));
 sg13g2_o21ai_1 _3424_ (.B1(net1078),
    .Y(_0904_),
    .A1(_0880_),
    .A2(_0881_));
 sg13g2_nand3_1 _3425_ (.B(_0903_),
    .C(_0904_),
    .A(net881),
    .Y(_0905_));
 sg13g2_nor4_1 _3426_ (.A(_0032_),
    .B(_0031_),
    .C(_1526_),
    .D(_0818_),
    .Y(_0906_));
 sg13g2_nand3_1 _3427_ (.B(_1561_),
    .C(net1086),
    .A(net1085),
    .Y(_0907_));
 sg13g2_nand3_1 _3428_ (.B(\a[0] ),
    .C(net855),
    .A(net2),
    .Y(_0908_));
 sg13g2_nor2_1 _3429_ (.A(net863),
    .B(net859),
    .Y(_0909_));
 sg13g2_nand3_1 _3430_ (.B(_0908_),
    .C(_0909_),
    .A(_0907_),
    .Y(_0910_));
 sg13g2_nand2_1 _3431_ (.Y(_0911_),
    .A(_1567_),
    .B(net1093));
 sg13g2_nand3_1 _3432_ (.B(net2),
    .C(net1094),
    .A(net1098),
    .Y(_0912_));
 sg13g2_and2_1 _3433_ (.A(\a[0] ),
    .B(net1084),
    .X(_0913_));
 sg13g2_o21ai_1 _3434_ (.B1(_0911_),
    .Y(_0914_),
    .A1(_0912_),
    .A2(_0913_));
 sg13g2_o21ai_1 _3435_ (.B1(_0914_),
    .Y(_0915_),
    .A1(net1083),
    .A2(net1084));
 sg13g2_nand2_1 _3436_ (.Y(_0916_),
    .A(_1565_),
    .B(net1093));
 sg13g2_nand2_1 _3437_ (.Y(_0917_),
    .A(_1561_),
    .B(net1093));
 sg13g2_and2_1 _3438_ (.A(net1085),
    .B(net1084),
    .X(_0918_));
 sg13g2_o21ai_1 _3439_ (.B1(_0916_),
    .Y(_0919_),
    .A1(_0917_),
    .A2(_0918_));
 sg13g2_o21ai_1 _3440_ (.B1(_0919_),
    .Y(_0920_),
    .A1(net1085),
    .A2(net1084));
 sg13g2_a22oi_1 _3441_ (.Y(_0921_),
    .B1(net851),
    .B2(\ayayayayayaya.b[31] ),
    .A2(net868),
    .A1(net1082));
 sg13g2_nand3_1 _3442_ (.B(_0920_),
    .C(_0921_),
    .A(net1104),
    .Y(_0922_));
 sg13g2_a21oi_1 _3443_ (.A1(net1084),
    .A2(_0910_),
    .Y(_0923_),
    .B1(_0922_));
 sg13g2_o21ai_1 _3444_ (.B1(_0923_),
    .Y(_0924_),
    .A1(_1376_),
    .A2(net873));
 sg13g2_nor2_1 _3445_ (.A(_0906_),
    .B(_0924_),
    .Y(_0925_));
 sg13g2_a22oi_1 _3446_ (.Y(_0926_),
    .B1(_0915_),
    .B2(_0925_),
    .A2(_0905_),
    .A1(_0902_));
 sg13g2_o21ai_1 _3447_ (.B1(net885),
    .Y(_0927_),
    .A1(_0197_),
    .A2(_0198_));
 sg13g2_o21ai_1 _3448_ (.B1(net1081),
    .Y(_0928_),
    .A1(_0854_),
    .A2(_0855_));
 sg13g2_nand3_1 _3449_ (.B(_0927_),
    .C(_0928_),
    .A(net877),
    .Y(_0929_));
 sg13g2_nand2_1 _3450_ (.Y(_0930_),
    .A(net1076),
    .B(_0861_));
 sg13g2_a21oi_1 _3451_ (.A1(net884),
    .A2(_0307_),
    .Y(_0931_),
    .B1(net872));
 sg13g2_o21ai_1 _3452_ (.B1(\a[7] ),
    .Y(_0932_),
    .A1(net859),
    .A2(_0325_));
 sg13g2_nand3_1 _3453_ (.B(net1093),
    .C(_0863_),
    .A(\a[8] ),
    .Y(_0933_));
 sg13g2_a22oi_1 _3454_ (.Y(_0934_),
    .B1(net863),
    .B2(\a[19] ),
    .A2(net868),
    .A1(\a[3] ));
 sg13g2_a21oi_1 _3455_ (.A1(net1025),
    .A2(net850),
    .Y(_0935_),
    .B1(net1104));
 sg13g2_nand4_1 _3456_ (.B(_0933_),
    .C(_0934_),
    .A(_0932_),
    .Y(_0936_),
    .D(_0935_));
 sg13g2_a21oi_1 _3457_ (.A1(_0930_),
    .A2(_0931_),
    .Y(_0937_),
    .B1(_0936_));
 sg13g2_o21ai_1 _3458_ (.B1(net1078),
    .Y(_0938_),
    .A1(_0840_),
    .A2(_0841_));
 sg13g2_o21ai_1 _3459_ (.B1(net886),
    .Y(_0939_),
    .A1(_1557_),
    .A2(_1558_));
 sg13g2_nand3_1 _3460_ (.B(_0938_),
    .C(_0939_),
    .A(net879),
    .Y(_0940_));
 sg13g2_nor4_1 _3461_ (.A(_0032_),
    .B(_0031_),
    .C(net872),
    .D(_0784_),
    .Y(_0941_));
 sg13g2_and2_1 _3462_ (.A(net1082),
    .B(net1085),
    .X(_0942_));
 sg13g2_o21ai_1 _3463_ (.B1(_0911_),
    .Y(_0943_),
    .A1(_0912_),
    .A2(_0942_));
 sg13g2_o21ai_1 _3464_ (.B1(_0943_),
    .Y(_0944_),
    .A1(net1082),
    .A2(net1085));
 sg13g2_and2_1 _3465_ (.A(net1083),
    .B(net1082),
    .X(_0945_));
 sg13g2_o21ai_1 _3466_ (.B1(_0916_),
    .Y(_0946_),
    .A1(_0917_),
    .A2(_0945_));
 sg13g2_o21ai_1 _3467_ (.B1(_0946_),
    .Y(_0947_),
    .A1(net1083),
    .A2(net1082));
 sg13g2_a21oi_1 _3468_ (.A1(net991),
    .A2(net851),
    .Y(_0948_),
    .B1(net1096));
 sg13g2_a22oi_1 _3469_ (.Y(_0949_),
    .B1(net863),
    .B2(\a[23] ),
    .A2(net867),
    .A1(\a[7] ));
 sg13g2_nand4_1 _3470_ (.B(_0947_),
    .C(_0948_),
    .A(_0944_),
    .Y(_0950_),
    .D(_0949_));
 sg13g2_nand3_1 _3471_ (.B(net1085),
    .C(net855),
    .A(net2),
    .Y(_0951_));
 sg13g2_nand3_1 _3472_ (.B(_1561_),
    .C(net1086),
    .A(net1083),
    .Y(_0952_));
 sg13g2_nand3_1 _3473_ (.B(_0951_),
    .C(_0952_),
    .A(net858),
    .Y(_0953_));
 sg13g2_and2_1 _3474_ (.A(net1082),
    .B(_0953_),
    .X(_0954_));
 sg13g2_nor3_1 _3475_ (.A(_0941_),
    .B(_0950_),
    .C(_0954_),
    .Y(_0955_));
 sg13g2_a221oi_1 _3476_ (.B2(_0955_),
    .C1(net1103),
    .B1(_0940_),
    .A1(_0929_),
    .Y(_0956_),
    .A2(_0937_));
 sg13g2_a21o_2 _3477_ (.A2(_0926_),
    .A1(net1103),
    .B1(_0956_),
    .X(uio_out[7]));
 sg13g2_nand2_2 _3478_ (.Y(_0957_),
    .A(net1),
    .B(net1095));
 sg13g2_nor3_2 _3479_ (.A(net6),
    .B(net857),
    .C(_0957_),
    .Y(_0958_));
 sg13g2_mux2_1 _3480_ (.A0(net80),
    .A1(net7),
    .S(_0958_),
    .X(_0060_));
 sg13g2_mux2_1 _3481_ (.A0(net106),
    .A1(net8),
    .S(_0958_),
    .X(_0061_));
 sg13g2_mux2_1 _3482_ (.A0(net105),
    .A1(net9),
    .S(_0958_),
    .X(_0062_));
 sg13g2_mux2_1 _3483_ (.A0(net100),
    .A1(net10),
    .S(_0958_),
    .X(_0063_));
 sg13g2_mux2_1 _3484_ (.A0(net112),
    .A1(net11),
    .S(_0958_),
    .X(_0064_));
 sg13g2_mux2_1 _3485_ (.A0(net95),
    .A1(net12),
    .S(_0958_),
    .X(_0065_));
 sg13g2_mux2_1 _3486_ (.A0(net91),
    .A1(net13),
    .S(_0958_),
    .X(_0066_));
 sg13g2_mux2_1 _3487_ (.A0(net109),
    .A1(net14),
    .S(_0958_),
    .X(_0067_));
 sg13g2_nand2_1 _3488_ (.Y(_0959_),
    .A(net1103),
    .B(net1104));
 sg13g2_nor3_2 _3489_ (.A(net6),
    .B(net858),
    .C(_0959_),
    .Y(_0960_));
 sg13g2_mux2_1 _3490_ (.A0(net93),
    .A1(net7),
    .S(_0960_),
    .X(_0068_));
 sg13g2_mux2_1 _3491_ (.A0(net97),
    .A1(net8),
    .S(_0960_),
    .X(_0069_));
 sg13g2_mux2_1 _3492_ (.A0(net81),
    .A1(net9),
    .S(_0960_),
    .X(_0070_));
 sg13g2_mux2_1 _3493_ (.A0(net103),
    .A1(net10),
    .S(_0960_),
    .X(_0071_));
 sg13g2_mux2_1 _3494_ (.A0(net87),
    .A1(net11),
    .S(_0960_),
    .X(_0072_));
 sg13g2_mux2_1 _3495_ (.A0(net88),
    .A1(net12),
    .S(_0960_),
    .X(_0073_));
 sg13g2_mux2_1 _3496_ (.A0(net83),
    .A1(net13),
    .S(_0960_),
    .X(_0074_));
 sg13g2_mux2_1 _3497_ (.A0(net1084),
    .A1(net14),
    .S(_0960_),
    .X(_0075_));
 sg13g2_nor4_2 _3498_ (.A(net6),
    .B(net1103),
    .C(net1106),
    .Y(_0961_),
    .D(net858));
 sg13g2_mux2_1 _3499_ (.A0(net1083),
    .A1(net7),
    .S(_0961_),
    .X(_0076_));
 sg13g2_mux2_1 _3500_ (.A0(net89),
    .A1(net8),
    .S(_0961_),
    .X(_0077_));
 sg13g2_mux2_1 _3501_ (.A0(net99),
    .A1(net9),
    .S(_0961_),
    .X(_0078_));
 sg13g2_mux2_1 _3502_ (.A0(net90),
    .A1(net10),
    .S(_0961_),
    .X(_0079_));
 sg13g2_mux2_1 _3503_ (.A0(net82),
    .A1(net11),
    .S(_0961_),
    .X(_0080_));
 sg13g2_mux2_1 _3504_ (.A0(net96),
    .A1(net12),
    .S(_0961_),
    .X(_0081_));
 sg13g2_mux2_1 _3505_ (.A0(net101),
    .A1(net13),
    .S(_0961_),
    .X(_0082_));
 sg13g2_mux2_1 _3506_ (.A0(net85),
    .A1(net14),
    .S(_0961_),
    .X(_0083_));
 sg13g2_nand2_1 _3507_ (.Y(_0962_),
    .A(net1097),
    .B(net1105));
 sg13g2_nor3_2 _3508_ (.A(net6),
    .B(net857),
    .C(_0962_),
    .Y(_0963_));
 sg13g2_mux2_1 _3509_ (.A0(net84),
    .A1(net7),
    .S(_0963_),
    .X(_0084_));
 sg13g2_mux2_1 _3510_ (.A0(net92),
    .A1(net8),
    .S(_0963_),
    .X(_0085_));
 sg13g2_mux2_1 _3511_ (.A0(net102),
    .A1(net9),
    .S(_0963_),
    .X(_0086_));
 sg13g2_mux2_1 _3512_ (.A0(net111),
    .A1(net10),
    .S(_0963_),
    .X(_0087_));
 sg13g2_mux2_1 _3513_ (.A0(net107),
    .A1(net11),
    .S(_0963_),
    .X(_0088_));
 sg13g2_mux2_1 _3514_ (.A0(net110),
    .A1(net12),
    .S(_0963_),
    .X(_0089_));
 sg13g2_mux2_1 _3515_ (.A0(net86),
    .A1(net13),
    .S(_0963_),
    .X(_0090_));
 sg13g2_mux2_1 _3516_ (.A0(net79),
    .A1(net14),
    .S(_0963_),
    .X(_0091_));
 sg13g2_nor4_2 _3517_ (.A(net6),
    .B(net1103),
    .C(net1104),
    .Y(_0964_),
    .D(_1583_));
 sg13g2_nand2_1 _3518_ (.Y(_0965_),
    .A(net7),
    .B(_0964_));
 sg13g2_o21ai_1 _3519_ (.B1(_0965_),
    .Y(_0092_),
    .A1(net884),
    .A2(net849));
 sg13g2_nand2_1 _3520_ (.Y(_0966_),
    .A(net8),
    .B(net849));
 sg13g2_o21ai_1 _3521_ (.B1(_0966_),
    .Y(_0093_),
    .A1(net890),
    .A2(net849));
 sg13g2_nand2_1 _3522_ (.Y(_0967_),
    .A(net9),
    .B(net849));
 sg13g2_o21ai_1 _3523_ (.B1(_0967_),
    .Y(_0094_),
    .A1(net897),
    .A2(net849));
 sg13g2_nand2_1 _3524_ (.Y(_0968_),
    .A(net10),
    .B(net849));
 sg13g2_o21ai_1 _3525_ (.B1(_0968_),
    .Y(_0095_),
    .A1(net902),
    .A2(net849));
 sg13g2_nand2_1 _3526_ (.Y(_0969_),
    .A(net11),
    .B(net848));
 sg13g2_o21ai_1 _3527_ (.B1(_0969_),
    .Y(_0096_),
    .A1(net908),
    .A2(net848));
 sg13g2_nand2_1 _3528_ (.Y(_0970_),
    .A(net12),
    .B(net848));
 sg13g2_o21ai_1 _3529_ (.B1(_0970_),
    .Y(_0097_),
    .A1(net913),
    .A2(net848));
 sg13g2_nand2_1 _3530_ (.Y(_0971_),
    .A(net13),
    .B(net848));
 sg13g2_o21ai_1 _3531_ (.B1(_0971_),
    .Y(_0098_),
    .A1(net919),
    .A2(net848));
 sg13g2_nand2_1 _3532_ (.Y(_0972_),
    .A(net14),
    .B(net848));
 sg13g2_o21ai_1 _3533_ (.B1(_0972_),
    .Y(_0099_),
    .A1(net924),
    .A2(net848));
 sg13g2_nor3_1 _3534_ (.A(net6),
    .B(_1583_),
    .C(_0962_),
    .Y(_0973_));
 sg13g2_nand2_1 _3535_ (.Y(_0974_),
    .A(net7),
    .B(net847));
 sg13g2_o21ai_1 _3536_ (.B1(_0974_),
    .Y(_0100_),
    .A1(net932),
    .A2(net847));
 sg13g2_nand2_1 _3537_ (.Y(_0975_),
    .A(net8),
    .B(net847));
 sg13g2_o21ai_1 _3538_ (.B1(_0975_),
    .Y(_0101_),
    .A1(net937),
    .A2(net847));
 sg13g2_nand2_1 _3539_ (.Y(_0976_),
    .A(net9),
    .B(net845));
 sg13g2_o21ai_1 _3540_ (.B1(_0976_),
    .Y(_0102_),
    .A1(net939),
    .A2(net845));
 sg13g2_nand2_1 _3541_ (.Y(_0977_),
    .A(net10),
    .B(net845));
 sg13g2_o21ai_1 _3542_ (.B1(_0977_),
    .Y(_0103_),
    .A1(net944),
    .A2(net845));
 sg13g2_nand2_1 _3543_ (.Y(_0978_),
    .A(net11),
    .B(net845));
 sg13g2_o21ai_1 _3544_ (.B1(_0978_),
    .Y(_0104_),
    .A1(net947),
    .A2(net845));
 sg13g2_nand2_1 _3545_ (.Y(_0979_),
    .A(net12),
    .B(net845));
 sg13g2_o21ai_1 _3546_ (.B1(_0979_),
    .Y(_0105_),
    .A1(net952),
    .A2(net845));
 sg13g2_nand2_1 _3547_ (.Y(_0980_),
    .A(net13),
    .B(net846));
 sg13g2_o21ai_1 _3548_ (.B1(_0980_),
    .Y(_0106_),
    .A1(_1016_),
    .A2(net846));
 sg13g2_nand2_1 _3549_ (.Y(_0981_),
    .A(net14),
    .B(net846));
 sg13g2_o21ai_1 _3550_ (.B1(_0981_),
    .Y(_0107_),
    .A1(net955),
    .A2(net846));
 sg13g2_nor3_2 _3551_ (.A(net6),
    .B(_1583_),
    .C(_0957_),
    .Y(_0982_));
 sg13g2_nand2_1 _3552_ (.Y(_0983_),
    .A(net7),
    .B(net843));
 sg13g2_o21ai_1 _3553_ (.B1(_0983_),
    .Y(_0108_),
    .A1(net957),
    .A2(net843));
 sg13g2_nand2_1 _3554_ (.Y(_0984_),
    .A(net8),
    .B(net843));
 sg13g2_o21ai_1 _3555_ (.B1(_0984_),
    .Y(_0109_),
    .A1(net960),
    .A2(net843));
 sg13g2_nand2_1 _3556_ (.Y(_0985_),
    .A(net9),
    .B(net843));
 sg13g2_o21ai_1 _3557_ (.B1(_0985_),
    .Y(_0110_),
    .A1(net962),
    .A2(net843));
 sg13g2_nand2_1 _3558_ (.Y(_0986_),
    .A(net10),
    .B(net843));
 sg13g2_o21ai_1 _3559_ (.B1(_0986_),
    .Y(_0111_),
    .A1(net964),
    .A2(net843));
 sg13g2_nand2_1 _3560_ (.Y(_0987_),
    .A(net11),
    .B(net844));
 sg13g2_o21ai_1 _3561_ (.B1(_0987_),
    .Y(_0112_),
    .A1(_1010_),
    .A2(net844));
 sg13g2_nand2_1 _3562_ (.Y(_0988_),
    .A(net12),
    .B(net844));
 sg13g2_o21ai_1 _3563_ (.B1(_0988_),
    .Y(_0113_),
    .A1(_1009_),
    .A2(net844));
 sg13g2_nand2_1 _3564_ (.Y(_0989_),
    .A(net13),
    .B(net844));
 sg13g2_o21ai_1 _3565_ (.B1(_0989_),
    .Y(_0114_),
    .A1(_1008_),
    .A2(net844));
 sg13g2_nand2_1 _3566_ (.Y(_0990_),
    .A(net14),
    .B(net844));
 sg13g2_o21ai_1 _3567_ (.B1(_0990_),
    .Y(_0115_),
    .A1(_1007_),
    .A2(net844));
 sg13g2_nor3_1 _3568_ (.A(net6),
    .B(_1583_),
    .C(_0959_),
    .Y(_0991_));
 sg13g2_nand2_1 _3569_ (.Y(_0992_),
    .A(net7),
    .B(net841));
 sg13g2_o21ai_1 _3570_ (.B1(_0992_),
    .Y(_0116_),
    .A1(_1006_),
    .A2(net841));
 sg13g2_nand2_1 _3571_ (.Y(_0993_),
    .A(net8),
    .B(net842));
 sg13g2_o21ai_1 _3572_ (.B1(_0993_),
    .Y(_0117_),
    .A1(_1005_),
    .A2(net841));
 sg13g2_nand2_1 _3573_ (.Y(_0994_),
    .A(net9),
    .B(net842));
 sg13g2_o21ai_1 _3574_ (.B1(_0994_),
    .Y(_0118_),
    .A1(_1004_),
    .A2(net841));
 sg13g2_nand2_1 _3575_ (.Y(_0995_),
    .A(net10),
    .B(net841));
 sg13g2_o21ai_1 _3576_ (.B1(_0995_),
    .Y(_0119_),
    .A1(_1003_),
    .A2(net841));
 sg13g2_nand2_1 _3577_ (.Y(_0996_),
    .A(net11),
    .B(net841));
 sg13g2_o21ai_1 _3578_ (.B1(_0996_),
    .Y(_0120_),
    .A1(_1002_),
    .A2(net841));
 sg13g2_nand2_1 _3579_ (.Y(_0997_),
    .A(net12),
    .B(net842));
 sg13g2_o21ai_1 _3580_ (.B1(_0997_),
    .Y(_0121_),
    .A1(_1001_),
    .A2(net842));
 sg13g2_mux2_1 _3581_ (.A0(net108),
    .A1(net13),
    .S(net842),
    .X(_0122_));
 sg13g2_mux2_1 _3582_ (.A0(net94),
    .A1(net14),
    .S(net842),
    .X(_0123_));
 sg13g2_dfrbp_1 _3583_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net69),
    .D(_0060_),
    .Q_N(_0016_),
    .Q(\a[16] ));
 sg13g2_dfrbp_1 _3584_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net68),
    .D(_0061_),
    .Q_N(_0017_),
    .Q(\a[17] ));
 sg13g2_dfrbp_1 _3585_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net67),
    .D(_0062_),
    .Q_N(_0018_),
    .Q(\a[18] ));
 sg13g2_dfrbp_1 _3586_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net66),
    .D(_0063_),
    .Q_N(_0019_),
    .Q(\a[19] ));
 sg13g2_dfrbp_1 _3587_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net65),
    .D(_0064_),
    .Q_N(_0020_),
    .Q(\a[20] ));
 sg13g2_dfrbp_1 _3588_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net64),
    .D(_0065_),
    .Q_N(_0021_),
    .Q(\a[21] ));
 sg13g2_dfrbp_1 _3589_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net63),
    .D(_0066_),
    .Q_N(_0022_),
    .Q(\a[22] ));
 sg13g2_dfrbp_1 _3590_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net62),
    .D(_0067_),
    .Q_N(_0023_),
    .Q(\a[23] ));
 sg13g2_dfrbp_1 _3591_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net61),
    .D(_0068_),
    .Q_N(_0024_),
    .Q(\a[24] ));
 sg13g2_dfrbp_1 _3592_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net60),
    .D(_0069_),
    .Q_N(_0025_),
    .Q(\a[25] ));
 sg13g2_dfrbp_1 _3593_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net59),
    .D(_0070_),
    .Q_N(_0026_),
    .Q(\a[26] ));
 sg13g2_dfrbp_1 _3594_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net58),
    .D(_0071_),
    .Q_N(_0027_),
    .Q(\a[27] ));
 sg13g2_dfrbp_1 _3595_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net57),
    .D(_0072_),
    .Q_N(_0028_),
    .Q(\a[28] ));
 sg13g2_dfrbp_1 _3596_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net56),
    .D(_0073_),
    .Q_N(_0029_),
    .Q(\a[29] ));
 sg13g2_dfrbp_1 _3597_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net55),
    .D(_0074_),
    .Q_N(_0030_),
    .Q(\a[30] ));
 sg13g2_dfrbp_1 _3598_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net54),
    .D(_0075_),
    .Q_N(_1786_),
    .Q(\a[31] ));
 sg13g2_dfrbp_1 _3599_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net53),
    .D(_0076_),
    .Q_N(_0000_),
    .Q(\a[0] ));
 sg13g2_dfrbp_1 _3600_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net52),
    .D(_0077_),
    .Q_N(_0001_),
    .Q(\a[1] ));
 sg13g2_dfrbp_1 _3601_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net51),
    .D(_0078_),
    .Q_N(_0002_),
    .Q(\a[2] ));
 sg13g2_dfrbp_1 _3602_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net50),
    .D(_0079_),
    .Q_N(_0003_),
    .Q(\a[3] ));
 sg13g2_dfrbp_1 _3603_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net49),
    .D(_0080_),
    .Q_N(_0004_),
    .Q(\a[4] ));
 sg13g2_dfrbp_1 _3604_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net48),
    .D(_0081_),
    .Q_N(_0005_),
    .Q(\a[5] ));
 sg13g2_dfrbp_1 _3605_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net47),
    .D(_0082_),
    .Q_N(_0006_),
    .Q(\a[6] ));
 sg13g2_dfrbp_1 _3606_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net46),
    .D(_0083_),
    .Q_N(_0007_),
    .Q(\a[7] ));
 sg13g2_dfrbp_1 _3607_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net45),
    .D(_0084_),
    .Q_N(_0008_),
    .Q(\a[8] ));
 sg13g2_dfrbp_1 _3608_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net44),
    .D(_0085_),
    .Q_N(_0009_),
    .Q(\a[9] ));
 sg13g2_dfrbp_1 _3609_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net43),
    .D(_0086_),
    .Q_N(_0010_),
    .Q(\a[10] ));
 sg13g2_dfrbp_1 _3610_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net42),
    .D(_0087_),
    .Q_N(_0011_),
    .Q(\a[11] ));
 sg13g2_dfrbp_1 _3611_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net41),
    .D(_0088_),
    .Q_N(_0012_),
    .Q(\a[12] ));
 sg13g2_dfrbp_1 _3612_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net40),
    .D(_0089_),
    .Q_N(_0013_),
    .Q(\a[13] ));
 sg13g2_dfrbp_1 _3613_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net39),
    .D(_0090_),
    .Q_N(_0014_),
    .Q(\a[14] ));
 sg13g2_dfrbp_1 _3614_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net38),
    .D(_0091_),
    .Q_N(_0015_),
    .Q(\a[15] ));
 sg13g2_dfrbp_1 _3615_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net37),
    .D(_0092_),
    .Q_N(_0031_),
    .Q(\ayayayayayaya.b[0] ));
 sg13g2_dfrbp_1 _3616_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net36),
    .D(_0093_),
    .Q_N(_0032_),
    .Q(\ayayayayayaya.b[1] ));
 sg13g2_dfrbp_1 _3617_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net35),
    .D(_0094_),
    .Q_N(_0033_),
    .Q(\ayayayayayaya.b[2] ));
 sg13g2_dfrbp_1 _3618_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net34),
    .D(_0095_),
    .Q_N(_0034_),
    .Q(\ayayayayayaya.b[3] ));
 sg13g2_dfrbp_1 _3619_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net33),
    .D(_0096_),
    .Q_N(_0035_),
    .Q(\ayayayayayaya.b[4] ));
 sg13g2_dfrbp_1 _3620_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net32),
    .D(_0097_),
    .Q_N(_0036_),
    .Q(\ayayayayayaya.b[5] ));
 sg13g2_dfrbp_1 _3621_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net31),
    .D(_0098_),
    .Q_N(_0037_),
    .Q(\ayayayayayaya.b[6] ));
 sg13g2_dfrbp_1 _3622_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net30),
    .D(_0099_),
    .Q_N(_0038_),
    .Q(\ayayayayayaya.b[7] ));
 sg13g2_dfrbp_1 _3623_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net29),
    .D(_0100_),
    .Q_N(_0039_),
    .Q(\ayayayayayaya.b[8] ));
 sg13g2_dfrbp_1 _3624_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net28),
    .D(_0101_),
    .Q_N(_0040_),
    .Q(\ayayayayayaya.b[9] ));
 sg13g2_dfrbp_1 _3625_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net27),
    .D(_0102_),
    .Q_N(_0041_),
    .Q(\ayayayayayaya.b[10] ));
 sg13g2_dfrbp_1 _3626_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net26),
    .D(_0103_),
    .Q_N(_0042_),
    .Q(\ayayayayayaya.b[11] ));
 sg13g2_dfrbp_1 _3627_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net25),
    .D(_0104_),
    .Q_N(_0043_),
    .Q(\ayayayayayaya.b[12] ));
 sg13g2_dfrbp_1 _3628_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net24),
    .D(_0105_),
    .Q_N(_0044_),
    .Q(\ayayayayayaya.b[13] ));
 sg13g2_dfrbp_1 _3629_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net23),
    .D(_0106_),
    .Q_N(_0045_),
    .Q(\ayayayayayaya.b[14] ));
 sg13g2_dfrbp_1 _3630_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net22),
    .D(_0107_),
    .Q_N(_0046_),
    .Q(\ayayayayayaya.b[15] ));
 sg13g2_dfrbp_1 _3631_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net21),
    .D(_0108_),
    .Q_N(_0047_),
    .Q(\ayayayayayaya.b[16] ));
 sg13g2_dfrbp_1 _3632_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net20),
    .D(_0109_),
    .Q_N(_0048_),
    .Q(\ayayayayayaya.b[17] ));
 sg13g2_dfrbp_1 _3633_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net19),
    .D(_0110_),
    .Q_N(_0049_),
    .Q(\ayayayayayaya.b[18] ));
 sg13g2_dfrbp_1 _3634_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net18),
    .D(_0111_),
    .Q_N(_0050_),
    .Q(\ayayayayayaya.b[19] ));
 sg13g2_dfrbp_1 _3635_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net17),
    .D(_0112_),
    .Q_N(_0051_),
    .Q(\ayayayayayaya.b[20] ));
 sg13g2_dfrbp_1 _3636_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net16),
    .D(_0113_),
    .Q_N(_0052_),
    .Q(\ayayayayayaya.b[21] ));
 sg13g2_dfrbp_1 _3637_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net15),
    .D(_0114_),
    .Q_N(_0053_),
    .Q(\ayayayayayaya.b[22] ));
 sg13g2_dfrbp_1 _3638_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net78),
    .D(_0115_),
    .Q_N(_0054_),
    .Q(\ayayayayayaya.b[23] ));
 sg13g2_dfrbp_1 _3639_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net77),
    .D(_0116_),
    .Q_N(_0055_),
    .Q(\ayayayayayaya.b[24] ));
 sg13g2_dfrbp_1 _3640_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net76),
    .D(_0117_),
    .Q_N(_0056_),
    .Q(\ayayayayayaya.b[25] ));
 sg13g2_dfrbp_1 _3641_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net75),
    .D(_0118_),
    .Q_N(_0057_),
    .Q(\ayayayayayaya.b[26] ));
 sg13g2_dfrbp_1 _3642_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net74),
    .D(_0119_),
    .Q_N(_0058_),
    .Q(\ayayayayayaya.b[27] ));
 sg13g2_dfrbp_1 _3643_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net73),
    .D(_0120_),
    .Q_N(_0059_),
    .Q(\ayayayayayaya.b[28] ));
 sg13g2_dfrbp_1 _3644_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net72),
    .D(_0121_),
    .Q_N(_1785_),
    .Q(\ayayayayayaya.b[29] ));
 sg13g2_dfrbp_1 _3645_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net71),
    .D(_0122_),
    .Q_N(_1784_),
    .Q(\ayayayayayaya.b[30] ));
 sg13g2_dfrbp_1 _3646_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net70),
    .D(_0123_),
    .Q_N(_1783_),
    .Q(\ayayayayayaya.b[31] ));
 sg13g2_tiehi _3636__16 (.L_HI(net16));
 sg13g2_tiehi _3635__17 (.L_HI(net17));
 sg13g2_tiehi _3634__18 (.L_HI(net18));
 sg13g2_tiehi _3633__19 (.L_HI(net19));
 sg13g2_tiehi _3632__20 (.L_HI(net20));
 sg13g2_tiehi _3631__21 (.L_HI(net21));
 sg13g2_tiehi _3630__22 (.L_HI(net22));
 sg13g2_tiehi _3629__23 (.L_HI(net23));
 sg13g2_tiehi _3628__24 (.L_HI(net24));
 sg13g2_tiehi _3627__25 (.L_HI(net25));
 sg13g2_tiehi _3626__26 (.L_HI(net26));
 sg13g2_tiehi _3625__27 (.L_HI(net27));
 sg13g2_tiehi _3624__28 (.L_HI(net28));
 sg13g2_tiehi _3623__29 (.L_HI(net29));
 sg13g2_tiehi _3622__30 (.L_HI(net30));
 sg13g2_tiehi _3621__31 (.L_HI(net31));
 sg13g2_tiehi _3620__32 (.L_HI(net32));
 sg13g2_tiehi _3619__33 (.L_HI(net33));
 sg13g2_tiehi _3618__34 (.L_HI(net34));
 sg13g2_tiehi _3617__35 (.L_HI(net35));
 sg13g2_tiehi _3616__36 (.L_HI(net36));
 sg13g2_tiehi _3615__37 (.L_HI(net37));
 sg13g2_tiehi _3614__38 (.L_HI(net38));
 sg13g2_tiehi _3613__39 (.L_HI(net39));
 sg13g2_tiehi _3612__40 (.L_HI(net40));
 sg13g2_tiehi _3611__41 (.L_HI(net41));
 sg13g2_tiehi _3610__42 (.L_HI(net42));
 sg13g2_tiehi _3609__43 (.L_HI(net43));
 sg13g2_tiehi _3608__44 (.L_HI(net44));
 sg13g2_tiehi _3607__45 (.L_HI(net45));
 sg13g2_tiehi _3606__46 (.L_HI(net46));
 sg13g2_tiehi _3605__47 (.L_HI(net47));
 sg13g2_tiehi _3604__48 (.L_HI(net48));
 sg13g2_tiehi _3603__49 (.L_HI(net49));
 sg13g2_tiehi _3602__50 (.L_HI(net50));
 sg13g2_tiehi _3601__51 (.L_HI(net51));
 sg13g2_tiehi _3600__52 (.L_HI(net52));
 sg13g2_tiehi _3599__53 (.L_HI(net53));
 sg13g2_tiehi _3598__54 (.L_HI(net54));
 sg13g2_tiehi _3597__55 (.L_HI(net55));
 sg13g2_tiehi _3596__56 (.L_HI(net56));
 sg13g2_tiehi _3595__57 (.L_HI(net57));
 sg13g2_tiehi _3594__58 (.L_HI(net58));
 sg13g2_tiehi _3593__59 (.L_HI(net59));
 sg13g2_tiehi _3592__60 (.L_HI(net60));
 sg13g2_tiehi _3591__61 (.L_HI(net61));
 sg13g2_tiehi _3590__62 (.L_HI(net62));
 sg13g2_tiehi _3589__63 (.L_HI(net63));
 sg13g2_tiehi _3588__64 (.L_HI(net64));
 sg13g2_tiehi _3587__65 (.L_HI(net65));
 sg13g2_tiehi _3586__66 (.L_HI(net66));
 sg13g2_tiehi _3585__67 (.L_HI(net67));
 sg13g2_tiehi _3584__68 (.L_HI(net68));
 sg13g2_tiehi _3583__69 (.L_HI(net69));
 sg13g2_tiehi _3646__70 (.L_HI(net70));
 sg13g2_tiehi _3645__71 (.L_HI(net71));
 sg13g2_tiehi _3644__72 (.L_HI(net72));
 sg13g2_tiehi _3643__73 (.L_HI(net73));
 sg13g2_tiehi _3642__74 (.L_HI(net74));
 sg13g2_tiehi _3641__75 (.L_HI(net75));
 sg13g2_tiehi _3640__76 (.L_HI(net76));
 sg13g2_tiehi _3639__77 (.L_HI(net77));
 sg13g2_tiehi _3638__78 (.L_HI(net78));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_1 _3711_ (.A(uio_oe[7]),
    .X(uio_oe[0]));
 sg13g2_buf_1 _3712_ (.A(uio_oe[7]),
    .X(uio_oe[1]));
 sg13g2_buf_1 _3713_ (.A(uio_oe[7]),
    .X(uio_oe[2]));
 sg13g2_buf_1 _3714_ (.A(uio_oe[7]),
    .X(uio_oe[3]));
 sg13g2_buf_1 _3715_ (.A(uio_oe[7]),
    .X(uio_oe[4]));
 sg13g2_buf_1 _3716_ (.A(uio_oe[7]),
    .X(uio_oe[5]));
 sg13g2_buf_1 _3717_ (.A(uio_oe[7]),
    .X(uio_oe[6]));
 sg13g2_buf_1 _3718_ (.A(uio_out[0]),
    .X(uo_out[0]));
 sg13g2_buf_1 _3719_ (.A(uio_out[1]),
    .X(uo_out[1]));
 sg13g2_buf_2 _3720_ (.A(uio_out[2]),
    .X(uo_out[2]));
 sg13g2_buf_2 _3721_ (.A(uio_out[3]),
    .X(uo_out[3]));
 sg13g2_buf_1 _3722_ (.A(uio_out[4]),
    .X(uo_out[4]));
 sg13g2_buf_1 _3723_ (.A(uio_out[5]),
    .X(uo_out[5]));
 sg13g2_buf_1 _3724_ (.A(uio_out[6]),
    .X(uo_out[6]));
 sg13g2_buf_2 _3725_ (.A(uio_out[7]),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout841 (.A(net842),
    .X(net841));
 sg13g2_buf_2 fanout842 (.A(_0991_),
    .X(net842));
 sg13g2_buf_2 fanout843 (.A(_0982_),
    .X(net843));
 sg13g2_buf_2 fanout844 (.A(_0982_),
    .X(net844));
 sg13g2_buf_2 fanout845 (.A(net847),
    .X(net845));
 sg13g2_buf_1 fanout846 (.A(net847),
    .X(net846));
 sg13g2_buf_4 fanout847 (.X(net847),
    .A(_0973_));
 sg13g2_buf_2 fanout848 (.A(net849),
    .X(net848));
 sg13g2_buf_2 fanout849 (.A(_0964_),
    .X(net849));
 sg13g2_buf_2 fanout850 (.A(net851),
    .X(net850));
 sg13g2_buf_2 fanout851 (.A(_1582_),
    .X(net851));
 sg13g2_buf_2 fanout852 (.A(net853),
    .X(net852));
 sg13g2_buf_2 fanout853 (.A(net854),
    .X(net853));
 sg13g2_buf_2 fanout854 (.A(_1582_),
    .X(net854));
 sg13g2_buf_2 fanout855 (.A(_1579_),
    .X(net855));
 sg13g2_buf_1 fanout856 (.A(_1579_),
    .X(net856));
 sg13g2_buf_4 fanout857 (.X(net857),
    .A(_1578_));
 sg13g2_buf_4 fanout858 (.X(net858),
    .A(_1578_));
 sg13g2_buf_2 fanout859 (.A(net861),
    .X(net859));
 sg13g2_buf_2 fanout860 (.A(net861),
    .X(net860));
 sg13g2_buf_2 fanout861 (.A(_1577_),
    .X(net861));
 sg13g2_buf_2 fanout862 (.A(net863),
    .X(net862));
 sg13g2_buf_2 fanout863 (.A(_1568_),
    .X(net863));
 sg13g2_buf_2 fanout864 (.A(net865),
    .X(net864));
 sg13g2_buf_1 fanout865 (.A(net866),
    .X(net865));
 sg13g2_buf_2 fanout866 (.A(_1568_),
    .X(net866));
 sg13g2_buf_2 fanout867 (.A(net869),
    .X(net867));
 sg13g2_buf_2 fanout868 (.A(net869),
    .X(net868));
 sg13g2_buf_1 fanout869 (.A(_1566_),
    .X(net869));
 sg13g2_buf_2 fanout870 (.A(net871),
    .X(net870));
 sg13g2_buf_2 fanout871 (.A(_1566_),
    .X(net871));
 sg13g2_buf_2 fanout872 (.A(net873),
    .X(net872));
 sg13g2_buf_2 fanout873 (.A(_1563_),
    .X(net873));
 sg13g2_buf_2 fanout874 (.A(net875),
    .X(net874));
 sg13g2_buf_2 fanout875 (.A(net876),
    .X(net875));
 sg13g2_buf_4 fanout876 (.X(net876),
    .A(_1562_));
 sg13g2_buf_2 fanout877 (.A(net881),
    .X(net877));
 sg13g2_buf_1 fanout878 (.A(net881),
    .X(net878));
 sg13g2_buf_2 fanout879 (.A(net880),
    .X(net879));
 sg13g2_buf_2 fanout880 (.A(net881),
    .X(net880));
 sg13g2_buf_2 fanout881 (.A(_1525_),
    .X(net881));
 sg13g2_buf_2 fanout882 (.A(net884),
    .X(net882));
 sg13g2_buf_2 fanout883 (.A(net884),
    .X(net883));
 sg13g2_buf_2 fanout884 (.A(_1030_),
    .X(net884));
 sg13g2_buf_2 fanout885 (.A(_1030_),
    .X(net885));
 sg13g2_buf_2 fanout886 (.A(net888),
    .X(net886));
 sg13g2_buf_1 fanout887 (.A(net888),
    .X(net887));
 sg13g2_buf_2 fanout888 (.A(_1030_),
    .X(net888));
 sg13g2_buf_2 fanout889 (.A(net890),
    .X(net889));
 sg13g2_buf_2 fanout890 (.A(net891),
    .X(net890));
 sg13g2_buf_2 fanout891 (.A(_1029_),
    .X(net891));
 sg13g2_buf_2 fanout892 (.A(_1029_),
    .X(net892));
 sg13g2_buf_2 fanout893 (.A(net895),
    .X(net893));
 sg13g2_buf_1 fanout894 (.A(net895),
    .X(net894));
 sg13g2_buf_2 fanout895 (.A(_1029_),
    .X(net895));
 sg13g2_buf_2 fanout896 (.A(net897),
    .X(net896));
 sg13g2_buf_2 fanout897 (.A(_1028_),
    .X(net897));
 sg13g2_buf_2 fanout898 (.A(_1028_),
    .X(net898));
 sg13g2_buf_2 fanout899 (.A(net900),
    .X(net899));
 sg13g2_buf_2 fanout900 (.A(net901),
    .X(net900));
 sg13g2_buf_2 fanout901 (.A(_1028_),
    .X(net901));
 sg13g2_buf_2 fanout902 (.A(net904),
    .X(net902));
 sg13g2_buf_1 fanout903 (.A(net904),
    .X(net903));
 sg13g2_buf_2 fanout904 (.A(_1027_),
    .X(net904));
 sg13g2_buf_2 fanout905 (.A(net907),
    .X(net905));
 sg13g2_buf_1 fanout906 (.A(net907),
    .X(net906));
 sg13g2_buf_2 fanout907 (.A(_1027_),
    .X(net907));
 sg13g2_buf_2 fanout908 (.A(_1026_),
    .X(net908));
 sg13g2_buf_2 fanout909 (.A(_1026_),
    .X(net909));
 sg13g2_buf_2 fanout910 (.A(net911),
    .X(net910));
 sg13g2_buf_2 fanout911 (.A(net912),
    .X(net911));
 sg13g2_buf_2 fanout912 (.A(_1026_),
    .X(net912));
 sg13g2_buf_2 fanout913 (.A(net915),
    .X(net913));
 sg13g2_buf_1 fanout914 (.A(net915),
    .X(net914));
 sg13g2_buf_2 fanout915 (.A(_1025_),
    .X(net915));
 sg13g2_buf_2 fanout916 (.A(net917),
    .X(net916));
 sg13g2_buf_2 fanout917 (.A(net918),
    .X(net917));
 sg13g2_buf_2 fanout918 (.A(_1025_),
    .X(net918));
 sg13g2_buf_2 fanout919 (.A(net920),
    .X(net919));
 sg13g2_buf_2 fanout920 (.A(_1024_),
    .X(net920));
 sg13g2_buf_2 fanout921 (.A(net923),
    .X(net921));
 sg13g2_buf_1 fanout922 (.A(net923),
    .X(net922));
 sg13g2_buf_2 fanout923 (.A(_1024_),
    .X(net923));
 sg13g2_buf_2 fanout924 (.A(net925),
    .X(net924));
 sg13g2_buf_2 fanout925 (.A(_1023_),
    .X(net925));
 sg13g2_buf_2 fanout926 (.A(net927),
    .X(net926));
 sg13g2_buf_2 fanout927 (.A(net928),
    .X(net927));
 sg13g2_buf_2 fanout928 (.A(_1023_),
    .X(net928));
 sg13g2_buf_2 fanout929 (.A(net933),
    .X(net929));
 sg13g2_buf_2 fanout930 (.A(net931),
    .X(net930));
 sg13g2_buf_2 fanout931 (.A(net932),
    .X(net931));
 sg13g2_buf_2 fanout932 (.A(net933),
    .X(net932));
 sg13g2_buf_2 fanout933 (.A(_1022_),
    .X(net933));
 sg13g2_buf_2 fanout934 (.A(net938),
    .X(net934));
 sg13g2_buf_2 fanout935 (.A(net937),
    .X(net935));
 sg13g2_buf_2 fanout936 (.A(net937),
    .X(net936));
 sg13g2_buf_2 fanout937 (.A(net938),
    .X(net937));
 sg13g2_buf_1 fanout938 (.A(_1021_),
    .X(net938));
 sg13g2_buf_4 fanout939 (.X(net939),
    .A(net941));
 sg13g2_buf_1 fanout940 (.A(net941),
    .X(net940));
 sg13g2_buf_1 fanout941 (.A(net942),
    .X(net941));
 sg13g2_buf_2 fanout942 (.A(_1020_),
    .X(net942));
 sg13g2_buf_2 fanout943 (.A(net946),
    .X(net943));
 sg13g2_buf_2 fanout944 (.A(net945),
    .X(net944));
 sg13g2_buf_2 fanout945 (.A(net946),
    .X(net945));
 sg13g2_buf_1 fanout946 (.A(_1019_),
    .X(net946));
 sg13g2_buf_2 fanout947 (.A(net948),
    .X(net947));
 sg13g2_buf_2 fanout948 (.A(_1018_),
    .X(net948));
 sg13g2_buf_2 fanout949 (.A(_1018_),
    .X(net949));
 sg13g2_buf_2 fanout950 (.A(net952),
    .X(net950));
 sg13g2_buf_2 fanout951 (.A(net952),
    .X(net951));
 sg13g2_buf_2 fanout952 (.A(_1017_),
    .X(net952));
 sg13g2_buf_2 fanout953 (.A(_1016_),
    .X(net953));
 sg13g2_buf_2 fanout954 (.A(_1016_),
    .X(net954));
 sg13g2_buf_2 fanout955 (.A(net956),
    .X(net955));
 sg13g2_buf_2 fanout956 (.A(_1015_),
    .X(net956));
 sg13g2_buf_2 fanout957 (.A(net958),
    .X(net957));
 sg13g2_buf_4 fanout958 (.X(net958),
    .A(_1014_));
 sg13g2_buf_4 fanout959 (.X(net959),
    .A(_1013_));
 sg13g2_buf_2 fanout960 (.A(_1013_),
    .X(net960));
 sg13g2_buf_4 fanout961 (.X(net961),
    .A(_1012_));
 sg13g2_buf_2 fanout962 (.A(_1012_),
    .X(net962));
 sg13g2_buf_4 fanout963 (.X(net963),
    .A(_1011_));
 sg13g2_buf_1 fanout964 (.A(_1011_),
    .X(net964));
 sg13g2_buf_4 fanout965 (.X(net965),
    .A(_1010_));
 sg13g2_buf_4 fanout966 (.X(net966),
    .A(_1009_));
 sg13g2_buf_4 fanout967 (.X(net967),
    .A(_1008_));
 sg13g2_buf_4 fanout968 (.X(net968),
    .A(\ayayayayayaya.b[25] ));
 sg13g2_buf_4 fanout969 (.X(net969),
    .A(\ayayayayayaya.b[24] ));
 sg13g2_buf_4 fanout970 (.X(net970),
    .A(net971));
 sg13g2_buf_2 fanout971 (.A(\ayayayayayaya.b[23] ),
    .X(net971));
 sg13g2_buf_4 fanout972 (.X(net972),
    .A(net973));
 sg13g2_buf_2 fanout973 (.A(\ayayayayayaya.b[22] ),
    .X(net973));
 sg13g2_buf_2 fanout974 (.A(net976),
    .X(net974));
 sg13g2_buf_2 fanout975 (.A(net976),
    .X(net975));
 sg13g2_buf_2 fanout976 (.A(\ayayayayayaya.b[21] ),
    .X(net976));
 sg13g2_buf_4 fanout977 (.X(net977),
    .A(net978));
 sg13g2_buf_2 fanout978 (.A(\ayayayayayaya.b[20] ),
    .X(net978));
 sg13g2_buf_4 fanout979 (.X(net979),
    .A(net980));
 sg13g2_buf_2 fanout980 (.A(\ayayayayayaya.b[19] ),
    .X(net980));
 sg13g2_buf_4 fanout981 (.X(net981),
    .A(net982));
 sg13g2_buf_2 fanout982 (.A(\ayayayayayaya.b[18] ),
    .X(net982));
 sg13g2_buf_4 fanout983 (.X(net983),
    .A(net985));
 sg13g2_buf_2 fanout984 (.A(net985),
    .X(net984));
 sg13g2_buf_2 fanout985 (.A(\ayayayayayaya.b[17] ),
    .X(net985));
 sg13g2_buf_4 fanout986 (.X(net986),
    .A(net987));
 sg13g2_buf_2 fanout987 (.A(\ayayayayayaya.b[16] ),
    .X(net987));
 sg13g2_buf_2 fanout988 (.A(net989),
    .X(net988));
 sg13g2_buf_1 fanout989 (.A(net991),
    .X(net989));
 sg13g2_buf_2 fanout990 (.A(net991),
    .X(net990));
 sg13g2_buf_2 fanout991 (.A(\ayayayayayaya.b[15] ),
    .X(net991));
 sg13g2_buf_2 fanout992 (.A(net993),
    .X(net992));
 sg13g2_buf_2 fanout993 (.A(net994),
    .X(net993));
 sg13g2_buf_2 fanout994 (.A(\ayayayayayaya.b[14] ),
    .X(net994));
 sg13g2_buf_2 fanout995 (.A(net998),
    .X(net995));
 sg13g2_buf_2 fanout996 (.A(net997),
    .X(net996));
 sg13g2_buf_1 fanout997 (.A(net998),
    .X(net997));
 sg13g2_buf_2 fanout998 (.A(\ayayayayayaya.b[13] ),
    .X(net998));
 sg13g2_buf_2 fanout999 (.A(net1002),
    .X(net999));
 sg13g2_buf_2 fanout1000 (.A(net1001),
    .X(net1000));
 sg13g2_buf_2 fanout1001 (.A(net1002),
    .X(net1001));
 sg13g2_buf_2 fanout1002 (.A(\ayayayayayaya.b[12] ),
    .X(net1002));
 sg13g2_buf_2 fanout1003 (.A(net1004),
    .X(net1003));
 sg13g2_buf_2 fanout1004 (.A(net1006),
    .X(net1004));
 sg13g2_buf_2 fanout1005 (.A(net1006),
    .X(net1005));
 sg13g2_buf_2 fanout1006 (.A(\ayayayayayaya.b[11] ),
    .X(net1006));
 sg13g2_buf_2 fanout1007 (.A(net1008),
    .X(net1007));
 sg13g2_buf_2 fanout1008 (.A(\ayayayayayaya.b[10] ),
    .X(net1008));
 sg13g2_buf_2 fanout1009 (.A(net1010),
    .X(net1009));
 sg13g2_buf_2 fanout1010 (.A(net1011),
    .X(net1010));
 sg13g2_buf_2 fanout1011 (.A(\ayayayayayaya.b[10] ),
    .X(net1011));
 sg13g2_buf_2 fanout1012 (.A(net1013),
    .X(net1012));
 sg13g2_buf_4 fanout1013 (.X(net1013),
    .A(\ayayayayayaya.b[9] ));
 sg13g2_buf_2 fanout1014 (.A(net1015),
    .X(net1014));
 sg13g2_buf_2 fanout1015 (.A(net1016),
    .X(net1015));
 sg13g2_buf_1 fanout1016 (.A(\ayayayayayaya.b[9] ),
    .X(net1016));
 sg13g2_buf_2 fanout1017 (.A(net1018),
    .X(net1017));
 sg13g2_buf_2 fanout1018 (.A(net1022),
    .X(net1018));
 sg13g2_buf_2 fanout1019 (.A(net1020),
    .X(net1019));
 sg13g2_buf_2 fanout1020 (.A(net1021),
    .X(net1020));
 sg13g2_buf_1 fanout1021 (.A(net1022),
    .X(net1021));
 sg13g2_buf_4 fanout1022 (.X(net1022),
    .A(\ayayayayayaya.b[8] ));
 sg13g2_buf_2 fanout1023 (.A(net1024),
    .X(net1023));
 sg13g2_buf_2 fanout1024 (.A(net1025),
    .X(net1024));
 sg13g2_buf_2 fanout1025 (.A(\ayayayayayaya.b[7] ),
    .X(net1025));
 sg13g2_buf_2 fanout1026 (.A(net1028),
    .X(net1026));
 sg13g2_buf_1 fanout1027 (.A(net1028),
    .X(net1027));
 sg13g2_buf_2 fanout1028 (.A(\ayayayayayaya.b[7] ),
    .X(net1028));
 sg13g2_buf_2 fanout1029 (.A(net1030),
    .X(net1029));
 sg13g2_buf_2 fanout1030 (.A(net1031),
    .X(net1030));
 sg13g2_buf_2 fanout1031 (.A(net1035),
    .X(net1031));
 sg13g2_buf_2 fanout1032 (.A(net1034),
    .X(net1032));
 sg13g2_buf_1 fanout1033 (.A(net1034),
    .X(net1033));
 sg13g2_buf_2 fanout1034 (.A(net1035),
    .X(net1034));
 sg13g2_buf_4 fanout1035 (.X(net1035),
    .A(\ayayayayayaya.b[6] ));
 sg13g2_buf_2 fanout1036 (.A(net1038),
    .X(net1036));
 sg13g2_buf_2 fanout1037 (.A(net1038),
    .X(net1037));
 sg13g2_buf_2 fanout1038 (.A(net1039),
    .X(net1038));
 sg13g2_buf_2 fanout1039 (.A(\ayayayayayaya.b[5] ),
    .X(net1039));
 sg13g2_buf_2 fanout1040 (.A(net1042),
    .X(net1040));
 sg13g2_buf_1 fanout1041 (.A(net1042),
    .X(net1041));
 sg13g2_buf_2 fanout1042 (.A(\ayayayayayaya.b[5] ),
    .X(net1042));
 sg13g2_buf_2 fanout1043 (.A(net1044),
    .X(net1043));
 sg13g2_buf_2 fanout1044 (.A(net1045),
    .X(net1044));
 sg13g2_buf_2 fanout1045 (.A(net1046),
    .X(net1045));
 sg13g2_buf_2 fanout1046 (.A(net1050),
    .X(net1046));
 sg13g2_buf_2 fanout1047 (.A(net1049),
    .X(net1047));
 sg13g2_buf_1 fanout1048 (.A(net1049),
    .X(net1048));
 sg13g2_buf_2 fanout1049 (.A(net1050),
    .X(net1049));
 sg13g2_buf_2 fanout1050 (.A(\ayayayayayaya.b[4] ),
    .X(net1050));
 sg13g2_buf_2 fanout1051 (.A(net1052),
    .X(net1051));
 sg13g2_buf_2 fanout1052 (.A(net1053),
    .X(net1052));
 sg13g2_buf_2 fanout1053 (.A(net1054),
    .X(net1053));
 sg13g2_buf_4 fanout1054 (.X(net1054),
    .A(net1057));
 sg13g2_buf_2 fanout1055 (.A(net1056),
    .X(net1055));
 sg13g2_buf_2 fanout1056 (.A(net1057),
    .X(net1056));
 sg13g2_buf_2 fanout1057 (.A(\ayayayayayaya.b[3] ),
    .X(net1057));
 sg13g2_buf_2 fanout1058 (.A(net1059),
    .X(net1058));
 sg13g2_buf_2 fanout1059 (.A(net1060),
    .X(net1059));
 sg13g2_buf_2 fanout1060 (.A(net1062),
    .X(net1060));
 sg13g2_buf_2 fanout1061 (.A(net1062),
    .X(net1061));
 sg13g2_buf_2 fanout1062 (.A(\ayayayayayaya.b[2] ),
    .X(net1062));
 sg13g2_buf_2 fanout1063 (.A(net1065),
    .X(net1063));
 sg13g2_buf_1 fanout1064 (.A(net1065),
    .X(net1064));
 sg13g2_buf_2 fanout1065 (.A(\ayayayayayaya.b[2] ),
    .X(net1065));
 sg13g2_buf_2 fanout1066 (.A(net1069),
    .X(net1066));
 sg13g2_buf_2 fanout1067 (.A(net1068),
    .X(net1067));
 sg13g2_buf_2 fanout1068 (.A(net1069),
    .X(net1068));
 sg13g2_buf_2 fanout1069 (.A(\ayayayayayaya.b[1] ),
    .X(net1069));
 sg13g2_buf_2 fanout1070 (.A(net1071),
    .X(net1070));
 sg13g2_buf_2 fanout1071 (.A(net1072),
    .X(net1071));
 sg13g2_buf_1 fanout1072 (.A(\ayayayayayaya.b[1] ),
    .X(net1072));
 sg13g2_buf_2 fanout1073 (.A(net1081),
    .X(net1073));
 sg13g2_buf_2 fanout1074 (.A(net1077),
    .X(net1074));
 sg13g2_buf_2 fanout1075 (.A(net1076),
    .X(net1075));
 sg13g2_buf_1 fanout1076 (.A(net1077),
    .X(net1076));
 sg13g2_buf_1 fanout1077 (.A(net1081),
    .X(net1077));
 sg13g2_buf_2 fanout1078 (.A(net1080),
    .X(net1078));
 sg13g2_buf_1 fanout1079 (.A(net1080),
    .X(net1079));
 sg13g2_buf_2 fanout1080 (.A(net1081),
    .X(net1080));
 sg13g2_buf_2 fanout1081 (.A(\ayayayayayaya.b[0] ),
    .X(net1081));
 sg13g2_buf_2 fanout1082 (.A(\a[15] ),
    .X(net1082));
 sg13g2_buf_2 fanout1083 (.A(net115),
    .X(net1083));
 sg13g2_buf_2 fanout1084 (.A(net114),
    .X(net1084));
 sg13g2_buf_2 fanout1085 (.A(\a[16] ),
    .X(net1085));
 sg13g2_buf_2 fanout1086 (.A(_1575_),
    .X(net1086));
 sg13g2_buf_1 fanout1087 (.A(_1575_),
    .X(net1087));
 sg13g2_buf_2 fanout1088 (.A(net1089),
    .X(net1088));
 sg13g2_buf_2 fanout1089 (.A(_1571_),
    .X(net1089));
 sg13g2_buf_2 fanout1090 (.A(net1092),
    .X(net1090));
 sg13g2_buf_1 fanout1091 (.A(net1092),
    .X(net1091));
 sg13g2_buf_2 fanout1092 (.A(_1571_),
    .X(net1092));
 sg13g2_buf_2 fanout1093 (.A(net1094),
    .X(net1093));
 sg13g2_buf_1 fanout1094 (.A(_1570_),
    .X(net1094));
 sg13g2_buf_2 fanout1095 (.A(net1096),
    .X(net1095));
 sg13g2_buf_2 fanout1096 (.A(_0999_),
    .X(net1096));
 sg13g2_buf_2 fanout1097 (.A(_0998_),
    .X(net1097));
 sg13g2_buf_2 fanout1098 (.A(net1100),
    .X(net1098));
 sg13g2_buf_2 fanout1099 (.A(net1100),
    .X(net1099));
 sg13g2_buf_2 fanout1100 (.A(ui_in[3]),
    .X(net1100));
 sg13g2_buf_2 fanout1101 (.A(net1102),
    .X(net1101));
 sg13g2_buf_1 fanout1102 (.A(ui_in[3]),
    .X(net1102));
 sg13g2_buf_2 fanout1103 (.A(net1),
    .X(net1103));
 sg13g2_buf_2 fanout1104 (.A(net1106),
    .X(net1104));
 sg13g2_buf_2 fanout1105 (.A(net1106),
    .X(net1105));
 sg13g2_buf_2 fanout1106 (.A(ui_in[0]),
    .X(net1106));
 sg13g2_buf_2 input1 (.A(ui_in[1]),
    .X(net1));
 sg13g2_buf_4 input2 (.X(net2),
    .A(ui_in[2]));
 sg13g2_buf_2 input3 (.A(ui_in[4]),
    .X(net3));
 sg13g2_buf_2 input4 (.A(ui_in[5]),
    .X(net4));
 sg13g2_buf_2 input5 (.A(ui_in[6]),
    .X(net5));
 sg13g2_buf_4 input6 (.X(net6),
    .A(ui_in[7]));
 sg13g2_buf_4 input7 (.X(net7),
    .A(uio_in[0]));
 sg13g2_buf_4 input8 (.X(net8),
    .A(uio_in[1]));
 sg13g2_buf_8 input9 (.A(uio_in[2]),
    .X(net9));
 sg13g2_buf_8 input10 (.A(uio_in[3]),
    .X(net10));
 sg13g2_buf_8 input11 (.A(uio_in[4]),
    .X(net11));
 sg13g2_buf_8 input12 (.A(uio_in[5]),
    .X(net12));
 sg13g2_buf_8 input13 (.A(uio_in[6]),
    .X(net13));
 sg13g2_buf_8 input14 (.A(uio_in[7]),
    .X(net14));
 sg13g2_tiehi _3637__15 (.L_HI(net15));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\a[15] ),
    .X(net79));
 sg13g2_dlygate4sd3_1 hold2 (.A(\a[16] ),
    .X(net80));
 sg13g2_dlygate4sd3_1 hold3 (.A(\a[26] ),
    .X(net81));
 sg13g2_dlygate4sd3_1 hold4 (.A(\a[4] ),
    .X(net82));
 sg13g2_dlygate4sd3_1 hold5 (.A(\a[30] ),
    .X(net83));
 sg13g2_dlygate4sd3_1 hold6 (.A(\a[8] ),
    .X(net84));
 sg13g2_dlygate4sd3_1 hold7 (.A(\a[7] ),
    .X(net85));
 sg13g2_dlygate4sd3_1 hold8 (.A(\a[14] ),
    .X(net86));
 sg13g2_dlygate4sd3_1 hold9 (.A(\a[28] ),
    .X(net87));
 sg13g2_dlygate4sd3_1 hold10 (.A(\a[29] ),
    .X(net88));
 sg13g2_dlygate4sd3_1 hold11 (.A(\a[1] ),
    .X(net89));
 sg13g2_dlygate4sd3_1 hold12 (.A(\a[3] ),
    .X(net90));
 sg13g2_dlygate4sd3_1 hold13 (.A(\a[22] ),
    .X(net91));
 sg13g2_dlygate4sd3_1 hold14 (.A(\a[9] ),
    .X(net92));
 sg13g2_dlygate4sd3_1 hold15 (.A(\a[24] ),
    .X(net93));
 sg13g2_dlygate4sd3_1 hold16 (.A(\ayayayayayaya.b[31] ),
    .X(net94));
 sg13g2_dlygate4sd3_1 hold17 (.A(\a[21] ),
    .X(net95));
 sg13g2_dlygate4sd3_1 hold18 (.A(\a[5] ),
    .X(net96));
 sg13g2_dlygate4sd3_1 hold19 (.A(\a[25] ),
    .X(net97));
 sg13g2_dlygate4sd3_1 hold20 (.A(\ayayayayayaya.b[24] ),
    .X(net98));
 sg13g2_dlygate4sd3_1 hold21 (.A(\a[2] ),
    .X(net99));
 sg13g2_dlygate4sd3_1 hold22 (.A(\a[19] ),
    .X(net100));
 sg13g2_dlygate4sd3_1 hold23 (.A(\a[6] ),
    .X(net101));
 sg13g2_dlygate4sd3_1 hold24 (.A(\a[10] ),
    .X(net102));
 sg13g2_dlygate4sd3_1 hold25 (.A(\a[27] ),
    .X(net103));
 sg13g2_dlygate4sd3_1 hold26 (.A(\ayayayayayaya.b[25] ),
    .X(net104));
 sg13g2_dlygate4sd3_1 hold27 (.A(\a[18] ),
    .X(net105));
 sg13g2_dlygate4sd3_1 hold28 (.A(\a[17] ),
    .X(net106));
 sg13g2_dlygate4sd3_1 hold29 (.A(\a[12] ),
    .X(net107));
 sg13g2_dlygate4sd3_1 hold30 (.A(\ayayayayayaya.b[30] ),
    .X(net108));
 sg13g2_dlygate4sd3_1 hold31 (.A(\a[23] ),
    .X(net109));
 sg13g2_dlygate4sd3_1 hold32 (.A(\a[13] ),
    .X(net110));
 sg13g2_dlygate4sd3_1 hold33 (.A(\a[11] ),
    .X(net111));
 sg13g2_dlygate4sd3_1 hold34 (.A(\a[20] ),
    .X(net112));
 sg13g2_dlygate4sd3_1 hold35 (.A(\ayayayayayaya.b[29] ),
    .X(net113));
 sg13g2_dlygate4sd3_1 hold36 (.A(\a[31] ),
    .X(net114));
 sg13g2_dlygate4sd3_1 hold37 (.A(\a[0] ),
    .X(net115));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_fill_2 FILLER_0_77 ();
 sg13g2_decap_4 FILLER_0_105 ();
 sg13g2_fill_2 FILLER_0_114 ();
 sg13g2_fill_1 FILLER_0_116 ();
 sg13g2_fill_1 FILLER_0_130 ();
 sg13g2_decap_4 FILLER_0_144 ();
 sg13g2_fill_2 FILLER_0_148 ();
 sg13g2_decap_8 FILLER_0_177 ();
 sg13g2_decap_4 FILLER_0_210 ();
 sg13g2_fill_2 FILLER_0_214 ();
 sg13g2_decap_8 FILLER_0_225 ();
 sg13g2_decap_4 FILLER_0_232 ();
 sg13g2_fill_2 FILLER_0_244 ();
 sg13g2_decap_8 FILLER_0_251 ();
 sg13g2_fill_2 FILLER_0_258 ();
 sg13g2_fill_1 FILLER_0_260 ();
 sg13g2_fill_2 FILLER_0_271 ();
 sg13g2_fill_1 FILLER_0_273 ();
 sg13g2_fill_2 FILLER_0_279 ();
 sg13g2_fill_1 FILLER_0_281 ();
 sg13g2_fill_2 FILLER_0_285 ();
 sg13g2_decap_8 FILLER_0_292 ();
 sg13g2_decap_4 FILLER_0_299 ();
 sg13g2_decap_8 FILLER_0_323 ();
 sg13g2_decap_8 FILLER_0_360 ();
 sg13g2_decap_8 FILLER_0_367 ();
 sg13g2_decap_8 FILLER_0_374 ();
 sg13g2_decap_8 FILLER_0_381 ();
 sg13g2_decap_8 FILLER_0_388 ();
 sg13g2_decap_8 FILLER_0_395 ();
 sg13g2_decap_8 FILLER_0_402 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_fill_1 FILLER_1_35 ();
 sg13g2_fill_2 FILLER_1_51 ();
 sg13g2_fill_1 FILLER_1_53 ();
 sg13g2_fill_1 FILLER_1_58 ();
 sg13g2_decap_4 FILLER_1_73 ();
 sg13g2_fill_1 FILLER_1_77 ();
 sg13g2_fill_1 FILLER_1_83 ();
 sg13g2_fill_1 FILLER_1_106 ();
 sg13g2_fill_1 FILLER_1_142 ();
 sg13g2_fill_2 FILLER_1_147 ();
 sg13g2_fill_2 FILLER_1_196 ();
 sg13g2_fill_1 FILLER_1_198 ();
 sg13g2_fill_2 FILLER_1_211 ();
 sg13g2_fill_1 FILLER_1_213 ();
 sg13g2_fill_2 FILLER_1_223 ();
 sg13g2_fill_1 FILLER_1_251 ();
 sg13g2_fill_2 FILLER_1_261 ();
 sg13g2_fill_1 FILLER_1_263 ();
 sg13g2_fill_2 FILLER_1_288 ();
 sg13g2_fill_2 FILLER_1_308 ();
 sg13g2_fill_1 FILLER_1_310 ();
 sg13g2_fill_1 FILLER_1_329 ();
 sg13g2_fill_2 FILLER_1_335 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_fill_2 FILLER_2_28 ();
 sg13g2_fill_2 FILLER_2_40 ();
 sg13g2_fill_1 FILLER_2_42 ();
 sg13g2_fill_2 FILLER_2_53 ();
 sg13g2_decap_4 FILLER_2_83 ();
 sg13g2_fill_1 FILLER_2_104 ();
 sg13g2_decap_4 FILLER_2_110 ();
 sg13g2_fill_2 FILLER_2_114 ();
 sg13g2_decap_4 FILLER_2_126 ();
 sg13g2_fill_2 FILLER_2_130 ();
 sg13g2_fill_2 FILLER_2_164 ();
 sg13g2_fill_1 FILLER_2_171 ();
 sg13g2_fill_1 FILLER_2_177 ();
 sg13g2_fill_2 FILLER_2_203 ();
 sg13g2_fill_1 FILLER_2_205 ();
 sg13g2_fill_2 FILLER_2_226 ();
 sg13g2_fill_1 FILLER_2_233 ();
 sg13g2_decap_8 FILLER_2_246 ();
 sg13g2_decap_4 FILLER_2_253 ();
 sg13g2_fill_1 FILLER_2_257 ();
 sg13g2_fill_2 FILLER_2_277 ();
 sg13g2_fill_1 FILLER_2_279 ();
 sg13g2_fill_2 FILLER_2_285 ();
 sg13g2_fill_1 FILLER_2_287 ();
 sg13g2_fill_1 FILLER_2_303 ();
 sg13g2_fill_2 FILLER_2_324 ();
 sg13g2_fill_1 FILLER_2_326 ();
 sg13g2_decap_4 FILLER_2_332 ();
 sg13g2_decap_8 FILLER_2_395 ();
 sg13g2_decap_8 FILLER_2_402 ();
 sg13g2_fill_2 FILLER_3_0 ();
 sg13g2_fill_1 FILLER_3_2 ();
 sg13g2_fill_2 FILLER_3_47 ();
 sg13g2_fill_1 FILLER_3_49 ();
 sg13g2_fill_2 FILLER_3_55 ();
 sg13g2_fill_1 FILLER_3_57 ();
 sg13g2_fill_2 FILLER_3_63 ();
 sg13g2_fill_1 FILLER_3_90 ();
 sg13g2_fill_2 FILLER_3_126 ();
 sg13g2_fill_1 FILLER_3_128 ();
 sg13g2_fill_1 FILLER_3_144 ();
 sg13g2_fill_1 FILLER_3_150 ();
 sg13g2_fill_2 FILLER_3_161 ();
 sg13g2_fill_1 FILLER_3_163 ();
 sg13g2_fill_2 FILLER_3_189 ();
 sg13g2_fill_2 FILLER_3_201 ();
 sg13g2_fill_1 FILLER_3_203 ();
 sg13g2_fill_2 FILLER_3_209 ();
 sg13g2_fill_2 FILLER_3_215 ();
 sg13g2_fill_2 FILLER_3_226 ();
 sg13g2_fill_2 FILLER_3_247 ();
 sg13g2_decap_4 FILLER_3_259 ();
 sg13g2_fill_2 FILLER_3_263 ();
 sg13g2_fill_1 FILLER_3_280 ();
 sg13g2_fill_2 FILLER_3_309 ();
 sg13g2_fill_2 FILLER_3_356 ();
 sg13g2_fill_1 FILLER_3_358 ();
 sg13g2_decap_8 FILLER_3_384 ();
 sg13g2_decap_8 FILLER_3_391 ();
 sg13g2_decap_8 FILLER_3_398 ();
 sg13g2_decap_4 FILLER_3_405 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_fill_1 FILLER_4_12 ();
 sg13g2_fill_1 FILLER_4_21 ();
 sg13g2_fill_2 FILLER_4_45 ();
 sg13g2_fill_2 FILLER_4_52 ();
 sg13g2_fill_1 FILLER_4_54 ();
 sg13g2_fill_2 FILLER_4_83 ();
 sg13g2_fill_1 FILLER_4_85 ();
 sg13g2_fill_1 FILLER_4_90 ();
 sg13g2_fill_1 FILLER_4_96 ();
 sg13g2_fill_2 FILLER_4_101 ();
 sg13g2_fill_2 FILLER_4_123 ();
 sg13g2_fill_1 FILLER_4_125 ();
 sg13g2_fill_1 FILLER_4_141 ();
 sg13g2_decap_4 FILLER_4_177 ();
 sg13g2_fill_2 FILLER_4_186 ();
 sg13g2_fill_2 FILLER_4_283 ();
 sg13g2_fill_1 FILLER_4_285 ();
 sg13g2_fill_1 FILLER_4_311 ();
 sg13g2_decap_4 FILLER_4_352 ();
 sg13g2_fill_1 FILLER_4_371 ();
 sg13g2_decap_4 FILLER_4_377 ();
 sg13g2_decap_8 FILLER_4_390 ();
 sg13g2_decap_8 FILLER_4_397 ();
 sg13g2_decap_4 FILLER_4_404 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_4 FILLER_5_16 ();
 sg13g2_fill_1 FILLER_5_20 ();
 sg13g2_fill_1 FILLER_5_71 ();
 sg13g2_fill_1 FILLER_5_115 ();
 sg13g2_fill_1 FILLER_5_131 ();
 sg13g2_fill_2 FILLER_5_142 ();
 sg13g2_fill_2 FILLER_5_149 ();
 sg13g2_fill_1 FILLER_5_151 ();
 sg13g2_decap_4 FILLER_5_162 ();
 sg13g2_decap_8 FILLER_5_186 ();
 sg13g2_fill_1 FILLER_5_193 ();
 sg13g2_decap_8 FILLER_5_214 ();
 sg13g2_decap_8 FILLER_5_221 ();
 sg13g2_fill_2 FILLER_5_228 ();
 sg13g2_fill_1 FILLER_5_230 ();
 sg13g2_decap_4 FILLER_5_241 ();
 sg13g2_decap_4 FILLER_5_270 ();
 sg13g2_fill_2 FILLER_5_279 ();
 sg13g2_fill_2 FILLER_5_296 ();
 sg13g2_fill_1 FILLER_5_303 ();
 sg13g2_decap_8 FILLER_5_314 ();
 sg13g2_fill_2 FILLER_5_321 ();
 sg13g2_fill_1 FILLER_5_323 ();
 sg13g2_decap_4 FILLER_5_338 ();
 sg13g2_fill_2 FILLER_5_342 ();
 sg13g2_fill_2 FILLER_5_373 ();
 sg13g2_fill_1 FILLER_5_375 ();
 sg13g2_decap_4 FILLER_5_403 ();
 sg13g2_fill_2 FILLER_5_407 ();
 sg13g2_fill_2 FILLER_6_0 ();
 sg13g2_fill_2 FILLER_6_28 ();
 sg13g2_fill_2 FILLER_6_50 ();
 sg13g2_fill_1 FILLER_6_52 ();
 sg13g2_fill_2 FILLER_6_58 ();
 sg13g2_decap_4 FILLER_6_74 ();
 sg13g2_decap_4 FILLER_6_83 ();
 sg13g2_fill_2 FILLER_6_87 ();
 sg13g2_fill_2 FILLER_6_110 ();
 sg13g2_fill_1 FILLER_6_112 ();
 sg13g2_fill_2 FILLER_6_133 ();
 sg13g2_fill_1 FILLER_6_149 ();
 sg13g2_decap_4 FILLER_6_165 ();
 sg13g2_fill_1 FILLER_6_169 ();
 sg13g2_fill_1 FILLER_6_180 ();
 sg13g2_fill_2 FILLER_6_186 ();
 sg13g2_decap_8 FILLER_6_212 ();
 sg13g2_decap_4 FILLER_6_224 ();
 sg13g2_fill_2 FILLER_6_228 ();
 sg13g2_fill_2 FILLER_6_245 ();
 sg13g2_fill_1 FILLER_6_247 ();
 sg13g2_fill_2 FILLER_6_278 ();
 sg13g2_fill_1 FILLER_6_280 ();
 sg13g2_fill_1 FILLER_6_286 ();
 sg13g2_fill_1 FILLER_6_315 ();
 sg13g2_decap_4 FILLER_6_321 ();
 sg13g2_decap_4 FILLER_6_333 ();
 sg13g2_fill_2 FILLER_6_337 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_fill_2 FILLER_7_16 ();
 sg13g2_fill_1 FILLER_7_38 ();
 sg13g2_fill_1 FILLER_7_52 ();
 sg13g2_fill_1 FILLER_7_80 ();
 sg13g2_decap_4 FILLER_7_101 ();
 sg13g2_decap_8 FILLER_7_145 ();
 sg13g2_fill_1 FILLER_7_162 ();
 sg13g2_decap_4 FILLER_7_183 ();
 sg13g2_fill_2 FILLER_7_187 ();
 sg13g2_fill_2 FILLER_7_209 ();
 sg13g2_fill_2 FILLER_7_261 ();
 sg13g2_fill_1 FILLER_7_263 ();
 sg13g2_decap_4 FILLER_7_356 ();
 sg13g2_fill_2 FILLER_7_365 ();
 sg13g2_fill_1 FILLER_7_367 ();
 sg13g2_fill_1 FILLER_7_392 ();
 sg13g2_fill_2 FILLER_8_40 ();
 sg13g2_decap_4 FILLER_8_71 ();
 sg13g2_decap_4 FILLER_8_110 ();
 sg13g2_fill_1 FILLER_8_114 ();
 sg13g2_fill_2 FILLER_8_120 ();
 sg13g2_fill_2 FILLER_8_127 ();
 sg13g2_fill_2 FILLER_8_134 ();
 sg13g2_fill_1 FILLER_8_136 ();
 sg13g2_fill_1 FILLER_8_142 ();
 sg13g2_fill_2 FILLER_8_163 ();
 sg13g2_fill_1 FILLER_8_165 ();
 sg13g2_fill_2 FILLER_8_186 ();
 sg13g2_fill_1 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_209 ();
 sg13g2_decap_4 FILLER_8_216 ();
 sg13g2_decap_4 FILLER_8_225 ();
 sg13g2_decap_4 FILLER_8_234 ();
 sg13g2_decap_4 FILLER_8_243 ();
 sg13g2_fill_2 FILLER_8_282 ();
 sg13g2_fill_2 FILLER_8_298 ();
 sg13g2_fill_1 FILLER_8_329 ();
 sg13g2_decap_4 FILLER_8_380 ();
 sg13g2_decap_4 FILLER_8_403 ();
 sg13g2_fill_2 FILLER_8_407 ();
 sg13g2_decap_4 FILLER_9_0 ();
 sg13g2_fill_1 FILLER_9_4 ();
 sg13g2_fill_2 FILLER_9_13 ();
 sg13g2_fill_2 FILLER_9_24 ();
 sg13g2_fill_1 FILLER_9_26 ();
 sg13g2_fill_2 FILLER_9_37 ();
 sg13g2_fill_1 FILLER_9_39 ();
 sg13g2_fill_2 FILLER_9_66 ();
 sg13g2_fill_1 FILLER_9_68 ();
 sg13g2_fill_2 FILLER_9_74 ();
 sg13g2_fill_2 FILLER_9_80 ();
 sg13g2_fill_2 FILLER_9_109 ();
 sg13g2_fill_2 FILLER_9_141 ();
 sg13g2_fill_1 FILLER_9_143 ();
 sg13g2_decap_4 FILLER_9_149 ();
 sg13g2_fill_1 FILLER_9_178 ();
 sg13g2_fill_1 FILLER_9_257 ();
 sg13g2_fill_1 FILLER_9_278 ();
 sg13g2_fill_1 FILLER_9_325 ();
 sg13g2_fill_1 FILLER_9_346 ();
 sg13g2_fill_2 FILLER_9_357 ();
 sg13g2_fill_1 FILLER_9_359 ();
 sg13g2_decap_4 FILLER_9_365 ();
 sg13g2_fill_2 FILLER_10_29 ();
 sg13g2_fill_2 FILLER_10_44 ();
 sg13g2_fill_1 FILLER_10_46 ();
 sg13g2_fill_2 FILLER_10_61 ();
 sg13g2_fill_1 FILLER_10_63 ();
 sg13g2_decap_4 FILLER_10_89 ();
 sg13g2_fill_1 FILLER_10_113 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_fill_2 FILLER_10_178 ();
 sg13g2_decap_8 FILLER_10_220 ();
 sg13g2_fill_2 FILLER_10_227 ();
 sg13g2_fill_1 FILLER_10_234 ();
 sg13g2_decap_4 FILLER_10_245 ();
 sg13g2_fill_2 FILLER_10_249 ();
 sg13g2_fill_2 FILLER_10_296 ();
 sg13g2_fill_2 FILLER_10_375 ();
 sg13g2_fill_1 FILLER_10_382 ();
 sg13g2_fill_1 FILLER_10_393 ();
 sg13g2_fill_2 FILLER_10_398 ();
 sg13g2_fill_2 FILLER_11_26 ();
 sg13g2_fill_1 FILLER_11_28 ();
 sg13g2_fill_1 FILLER_11_34 ();
 sg13g2_fill_2 FILLER_11_39 ();
 sg13g2_fill_1 FILLER_11_41 ();
 sg13g2_fill_1 FILLER_11_47 ();
 sg13g2_fill_1 FILLER_11_58 ();
 sg13g2_fill_2 FILLER_11_64 ();
 sg13g2_fill_1 FILLER_11_80 ();
 sg13g2_fill_1 FILLER_11_139 ();
 sg13g2_decap_4 FILLER_11_145 ();
 sg13g2_decap_8 FILLER_11_164 ();
 sg13g2_decap_8 FILLER_11_171 ();
 sg13g2_decap_4 FILLER_11_178 ();
 sg13g2_decap_8 FILLER_11_197 ();
 sg13g2_decap_8 FILLER_11_204 ();
 sg13g2_fill_1 FILLER_11_211 ();
 sg13g2_fill_1 FILLER_11_217 ();
 sg13g2_fill_2 FILLER_11_228 ();
 sg13g2_decap_4 FILLER_11_270 ();
 sg13g2_decap_4 FILLER_11_286 ();
 sg13g2_fill_2 FILLER_11_290 ();
 sg13g2_fill_2 FILLER_11_316 ();
 sg13g2_fill_1 FILLER_11_318 ();
 sg13g2_fill_1 FILLER_11_337 ();
 sg13g2_fill_1 FILLER_11_371 ();
 sg13g2_fill_2 FILLER_11_381 ();
 sg13g2_fill_2 FILLER_12_0 ();
 sg13g2_fill_1 FILLER_12_2 ();
 sg13g2_fill_1 FILLER_12_16 ();
 sg13g2_fill_2 FILLER_12_21 ();
 sg13g2_fill_1 FILLER_12_38 ();
 sg13g2_fill_1 FILLER_12_64 ();
 sg13g2_fill_2 FILLER_12_102 ();
 sg13g2_fill_2 FILLER_12_109 ();
 sg13g2_fill_2 FILLER_12_116 ();
 sg13g2_fill_1 FILLER_12_123 ();
 sg13g2_fill_2 FILLER_12_134 ();
 sg13g2_fill_1 FILLER_12_136 ();
 sg13g2_decap_8 FILLER_12_142 ();
 sg13g2_decap_8 FILLER_12_149 ();
 sg13g2_decap_4 FILLER_12_176 ();
 sg13g2_fill_2 FILLER_12_184 ();
 sg13g2_decap_8 FILLER_12_206 ();
 sg13g2_decap_8 FILLER_12_223 ();
 sg13g2_decap_4 FILLER_12_230 ();
 sg13g2_fill_2 FILLER_12_234 ();
 sg13g2_decap_8 FILLER_12_241 ();
 sg13g2_decap_4 FILLER_12_268 ();
 sg13g2_fill_1 FILLER_12_272 ();
 sg13g2_fill_1 FILLER_12_278 ();
 sg13g2_fill_1 FILLER_12_284 ();
 sg13g2_decap_4 FILLER_12_293 ();
 sg13g2_fill_2 FILLER_12_302 ();
 sg13g2_fill_2 FILLER_12_346 ();
 sg13g2_fill_2 FILLER_12_353 ();
 sg13g2_fill_1 FILLER_12_370 ();
 sg13g2_fill_2 FILLER_12_385 ();
 sg13g2_fill_2 FILLER_13_0 ();
 sg13g2_fill_1 FILLER_13_2 ();
 sg13g2_fill_2 FILLER_13_7 ();
 sg13g2_fill_2 FILLER_13_29 ();
 sg13g2_fill_1 FILLER_13_31 ();
 sg13g2_fill_2 FILLER_13_47 ();
 sg13g2_fill_2 FILLER_13_59 ();
 sg13g2_fill_2 FILLER_13_71 ();
 sg13g2_fill_1 FILLER_13_93 ();
 sg13g2_decap_4 FILLER_13_144 ();
 sg13g2_fill_1 FILLER_13_213 ();
 sg13g2_fill_2 FILLER_13_309 ();
 sg13g2_fill_1 FILLER_13_311 ();
 sg13g2_fill_2 FILLER_13_317 ();
 sg13g2_fill_1 FILLER_13_319 ();
 sg13g2_fill_1 FILLER_13_335 ();
 sg13g2_fill_1 FILLER_13_355 ();
 sg13g2_fill_2 FILLER_13_365 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_fill_2 FILLER_14_0 ();
 sg13g2_fill_1 FILLER_14_2 ();
 sg13g2_fill_1 FILLER_14_12 ();
 sg13g2_fill_2 FILLER_14_31 ();
 sg13g2_fill_1 FILLER_14_38 ();
 sg13g2_fill_2 FILLER_14_49 ();
 sg13g2_fill_2 FILLER_14_98 ();
 sg13g2_fill_1 FILLER_14_100 ();
 sg13g2_decap_4 FILLER_14_121 ();
 sg13g2_fill_2 FILLER_14_125 ();
 sg13g2_fill_1 FILLER_14_137 ();
 sg13g2_fill_1 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_179 ();
 sg13g2_decap_4 FILLER_14_186 ();
 sg13g2_fill_2 FILLER_14_190 ();
 sg13g2_fill_1 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_212 ();
 sg13g2_fill_2 FILLER_14_219 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_fill_1 FILLER_14_238 ();
 sg13g2_decap_4 FILLER_14_259 ();
 sg13g2_decap_4 FILLER_14_306 ();
 sg13g2_fill_1 FILLER_14_310 ();
 sg13g2_fill_1 FILLER_14_321 ();
 sg13g2_decap_4 FILLER_14_327 ();
 sg13g2_fill_2 FILLER_14_353 ();
 sg13g2_fill_1 FILLER_14_355 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_fill_1 FILLER_14_378 ();
 sg13g2_fill_2 FILLER_14_389 ();
 sg13g2_fill_2 FILLER_15_63 ();
 sg13g2_decap_4 FILLER_15_91 ();
 sg13g2_fill_2 FILLER_15_150 ();
 sg13g2_fill_1 FILLER_15_152 ();
 sg13g2_fill_1 FILLER_15_218 ();
 sg13g2_fill_2 FILLER_15_264 ();
 sg13g2_fill_1 FILLER_15_291 ();
 sg13g2_fill_1 FILLER_15_391 ();
 sg13g2_fill_2 FILLER_16_0 ();
 sg13g2_fill_2 FILLER_16_26 ();
 sg13g2_fill_1 FILLER_16_28 ();
 sg13g2_fill_2 FILLER_16_53 ();
 sg13g2_fill_2 FILLER_16_70 ();
 sg13g2_fill_1 FILLER_16_72 ();
 sg13g2_fill_2 FILLER_16_78 ();
 sg13g2_fill_1 FILLER_16_80 ();
 sg13g2_decap_4 FILLER_16_86 ();
 sg13g2_decap_4 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_4 FILLER_16_126 ();
 sg13g2_fill_2 FILLER_16_149 ();
 sg13g2_fill_1 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_167 ();
 sg13g2_fill_2 FILLER_16_174 ();
 sg13g2_fill_1 FILLER_16_176 ();
 sg13g2_decap_4 FILLER_16_217 ();
 sg13g2_fill_2 FILLER_16_221 ();
 sg13g2_fill_1 FILLER_16_228 ();
 sg13g2_fill_2 FILLER_16_243 ();
 sg13g2_decap_8 FILLER_16_260 ();
 sg13g2_fill_2 FILLER_16_267 ();
 sg13g2_fill_1 FILLER_16_269 ();
 sg13g2_fill_2 FILLER_16_274 ();
 sg13g2_decap_8 FILLER_16_281 ();
 sg13g2_fill_2 FILLER_16_288 ();
 sg13g2_decap_8 FILLER_16_305 ();
 sg13g2_decap_4 FILLER_16_312 ();
 sg13g2_fill_2 FILLER_16_316 ();
 sg13g2_fill_2 FILLER_16_353 ();
 sg13g2_fill_2 FILLER_16_365 ();
 sg13g2_fill_1 FILLER_16_376 ();
 sg13g2_fill_1 FILLER_16_387 ();
 sg13g2_fill_2 FILLER_16_407 ();
 sg13g2_fill_1 FILLER_17_0 ();
 sg13g2_fill_2 FILLER_17_27 ();
 sg13g2_fill_1 FILLER_17_29 ();
 sg13g2_fill_2 FILLER_17_45 ();
 sg13g2_fill_1 FILLER_17_47 ();
 sg13g2_fill_1 FILLER_17_68 ();
 sg13g2_fill_2 FILLER_17_74 ();
 sg13g2_fill_1 FILLER_17_76 ();
 sg13g2_fill_1 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_118 ();
 sg13g2_decap_4 FILLER_17_125 ();
 sg13g2_fill_1 FILLER_17_148 ();
 sg13g2_decap_8 FILLER_17_159 ();
 sg13g2_fill_2 FILLER_17_166 ();
 sg13g2_fill_2 FILLER_17_173 ();
 sg13g2_fill_2 FILLER_17_180 ();
 sg13g2_fill_1 FILLER_17_190 ();
 sg13g2_fill_2 FILLER_17_201 ();
 sg13g2_fill_1 FILLER_17_203 ();
 sg13g2_fill_1 FILLER_17_219 ();
 sg13g2_fill_2 FILLER_17_230 ();
 sg13g2_fill_1 FILLER_17_232 ();
 sg13g2_fill_1 FILLER_17_261 ();
 sg13g2_fill_2 FILLER_17_321 ();
 sg13g2_fill_2 FILLER_17_337 ();
 sg13g2_fill_2 FILLER_17_359 ();
 sg13g2_decap_4 FILLER_17_379 ();
 sg13g2_decap_4 FILLER_18_0 ();
 sg13g2_fill_1 FILLER_18_4 ();
 sg13g2_fill_2 FILLER_18_34 ();
 sg13g2_fill_2 FILLER_18_46 ();
 sg13g2_fill_1 FILLER_18_48 ();
 sg13g2_fill_2 FILLER_18_54 ();
 sg13g2_fill_2 FILLER_18_66 ();
 sg13g2_fill_2 FILLER_18_96 ();
 sg13g2_fill_2 FILLER_18_103 ();
 sg13g2_fill_1 FILLER_18_105 ();
 sg13g2_fill_1 FILLER_18_118 ();
 sg13g2_fill_2 FILLER_18_154 ();
 sg13g2_fill_2 FILLER_18_182 ();
 sg13g2_decap_8 FILLER_18_220 ();
 sg13g2_fill_1 FILLER_18_284 ();
 sg13g2_decap_8 FILLER_18_300 ();
 sg13g2_fill_1 FILLER_18_307 ();
 sg13g2_fill_2 FILLER_18_328 ();
 sg13g2_fill_1 FILLER_18_348 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_12 ();
 sg13g2_fill_1 FILLER_19_32 ();
 sg13g2_decap_8 FILLER_19_62 ();
 sg13g2_fill_1 FILLER_19_69 ();
 sg13g2_decap_8 FILLER_19_80 ();
 sg13g2_fill_2 FILLER_19_87 ();
 sg13g2_fill_1 FILLER_19_108 ();
 sg13g2_fill_2 FILLER_19_138 ();
 sg13g2_fill_2 FILLER_19_146 ();
 sg13g2_fill_1 FILLER_19_148 ();
 sg13g2_fill_1 FILLER_19_164 ();
 sg13g2_fill_1 FILLER_19_178 ();
 sg13g2_fill_2 FILLER_19_188 ();
 sg13g2_fill_2 FILLER_19_194 ();
 sg13g2_fill_2 FILLER_19_201 ();
 sg13g2_fill_1 FILLER_19_203 ();
 sg13g2_fill_2 FILLER_19_254 ();
 sg13g2_decap_4 FILLER_19_269 ();
 sg13g2_fill_1 FILLER_19_273 ();
 sg13g2_decap_4 FILLER_19_294 ();
 sg13g2_fill_2 FILLER_19_314 ();
 sg13g2_fill_2 FILLER_19_394 ();
 sg13g2_fill_1 FILLER_19_396 ();
 sg13g2_fill_2 FILLER_19_406 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_fill_1 FILLER_20_16 ();
 sg13g2_decap_4 FILLER_20_37 ();
 sg13g2_fill_2 FILLER_20_41 ();
 sg13g2_fill_2 FILLER_20_58 ();
 sg13g2_fill_2 FILLER_20_97 ();
 sg13g2_fill_2 FILLER_20_150 ();
 sg13g2_fill_2 FILLER_20_282 ();
 sg13g2_fill_1 FILLER_20_284 ();
 sg13g2_decap_4 FILLER_20_290 ();
 sg13g2_fill_1 FILLER_20_304 ();
 sg13g2_fill_1 FILLER_20_325 ();
 sg13g2_fill_2 FILLER_20_329 ();
 sg13g2_decap_4 FILLER_20_346 ();
 sg13g2_fill_1 FILLER_20_364 ();
 sg13g2_fill_2 FILLER_20_374 ();
 sg13g2_fill_2 FILLER_20_407 ();
 sg13g2_fill_1 FILLER_21_0 ();
 sg13g2_fill_1 FILLER_21_27 ();
 sg13g2_fill_1 FILLER_21_40 ();
 sg13g2_fill_1 FILLER_21_61 ();
 sg13g2_decap_4 FILLER_21_73 ();
 sg13g2_fill_2 FILLER_21_77 ();
 sg13g2_decap_4 FILLER_21_83 ();
 sg13g2_fill_1 FILLER_21_104 ();
 sg13g2_fill_2 FILLER_21_119 ();
 sg13g2_fill_1 FILLER_21_127 ();
 sg13g2_fill_2 FILLER_21_138 ();
 sg13g2_fill_2 FILLER_21_148 ();
 sg13g2_fill_1 FILLER_21_155 ();
 sg13g2_fill_2 FILLER_21_201 ();
 sg13g2_fill_2 FILLER_21_211 ();
 sg13g2_fill_2 FILLER_21_229 ();
 sg13g2_decap_8 FILLER_21_244 ();
 sg13g2_decap_4 FILLER_21_251 ();
 sg13g2_fill_2 FILLER_21_255 ();
 sg13g2_fill_1 FILLER_21_261 ();
 sg13g2_decap_4 FILLER_21_315 ();
 sg13g2_fill_2 FILLER_21_338 ();
 sg13g2_fill_1 FILLER_21_340 ();
 sg13g2_fill_1 FILLER_21_346 ();
 sg13g2_fill_2 FILLER_21_364 ();
 sg13g2_fill_1 FILLER_21_366 ();
 sg13g2_fill_2 FILLER_21_372 ();
 sg13g2_fill_2 FILLER_21_389 ();
 sg13g2_fill_2 FILLER_21_396 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_fill_1 FILLER_22_14 ();
 sg13g2_fill_2 FILLER_22_39 ();
 sg13g2_fill_1 FILLER_22_41 ();
 sg13g2_fill_2 FILLER_22_47 ();
 sg13g2_fill_2 FILLER_22_71 ();
 sg13g2_fill_1 FILLER_22_73 ();
 sg13g2_decap_8 FILLER_22_103 ();
 sg13g2_decap_4 FILLER_22_110 ();
 sg13g2_fill_1 FILLER_22_133 ();
 sg13g2_fill_1 FILLER_22_148 ();
 sg13g2_fill_2 FILLER_22_169 ();
 sg13g2_fill_1 FILLER_22_171 ();
 sg13g2_decap_8 FILLER_22_176 ();
 sg13g2_decap_4 FILLER_22_199 ();
 sg13g2_fill_2 FILLER_22_209 ();
 sg13g2_fill_1 FILLER_22_211 ();
 sg13g2_decap_4 FILLER_22_220 ();
 sg13g2_fill_2 FILLER_22_240 ();
 sg13g2_decap_8 FILLER_22_288 ();
 sg13g2_fill_1 FILLER_22_295 ();
 sg13g2_fill_2 FILLER_22_306 ();
 sg13g2_fill_1 FILLER_22_308 ();
 sg13g2_decap_8 FILLER_22_319 ();
 sg13g2_fill_1 FILLER_22_326 ();
 sg13g2_fill_1 FILLER_22_382 ();
 sg13g2_fill_2 FILLER_23_39 ();
 sg13g2_fill_1 FILLER_23_41 ();
 sg13g2_fill_1 FILLER_23_54 ();
 sg13g2_fill_2 FILLER_23_84 ();
 sg13g2_fill_1 FILLER_23_86 ();
 sg13g2_decap_4 FILLER_23_101 ();
 sg13g2_fill_1 FILLER_23_117 ();
 sg13g2_decap_8 FILLER_23_146 ();
 sg13g2_decap_4 FILLER_23_153 ();
 sg13g2_fill_2 FILLER_23_157 ();
 sg13g2_fill_1 FILLER_23_164 ();
 sg13g2_decap_4 FILLER_23_179 ();
 sg13g2_fill_1 FILLER_23_213 ();
 sg13g2_decap_8 FILLER_23_255 ();
 sg13g2_fill_1 FILLER_23_262 ();
 sg13g2_decap_8 FILLER_23_272 ();
 sg13g2_decap_4 FILLER_23_279 ();
 sg13g2_fill_2 FILLER_23_283 ();
 sg13g2_decap_8 FILLER_23_290 ();
 sg13g2_fill_1 FILLER_23_297 ();
 sg13g2_decap_4 FILLER_23_324 ();
 sg13g2_fill_2 FILLER_23_328 ();
 sg13g2_decap_8 FILLER_23_335 ();
 sg13g2_decap_4 FILLER_23_342 ();
 sg13g2_fill_2 FILLER_23_346 ();
 sg13g2_fill_1 FILLER_23_356 ();
 sg13g2_fill_1 FILLER_23_362 ();
 sg13g2_fill_2 FILLER_23_377 ();
 sg13g2_fill_1 FILLER_23_379 ();
 sg13g2_fill_1 FILLER_23_385 ();
 sg13g2_fill_1 FILLER_23_394 ();
 sg13g2_fill_2 FILLER_23_407 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_fill_2 FILLER_24_58 ();
 sg13g2_fill_2 FILLER_24_87 ();
 sg13g2_fill_1 FILLER_24_89 ();
 sg13g2_fill_2 FILLER_24_116 ();
 sg13g2_fill_1 FILLER_24_118 ();
 sg13g2_fill_1 FILLER_24_146 ();
 sg13g2_fill_1 FILLER_24_170 ();
 sg13g2_decap_4 FILLER_24_198 ();
 sg13g2_fill_2 FILLER_24_207 ();
 sg13g2_fill_1 FILLER_24_209 ();
 sg13g2_decap_8 FILLER_24_259 ();
 sg13g2_fill_2 FILLER_24_266 ();
 sg13g2_decap_4 FILLER_24_272 ();
 sg13g2_decap_4 FILLER_24_290 ();
 sg13g2_fill_2 FILLER_24_303 ();
 sg13g2_fill_2 FILLER_24_361 ();
 sg13g2_fill_2 FILLER_24_407 ();
 sg13g2_decap_4 FILLER_25_0 ();
 sg13g2_fill_1 FILLER_25_4 ();
 sg13g2_fill_2 FILLER_25_54 ();
 sg13g2_decap_4 FILLER_25_77 ();
 sg13g2_fill_1 FILLER_25_87 ();
 sg13g2_fill_1 FILLER_25_93 ();
 sg13g2_fill_2 FILLER_25_108 ();
 sg13g2_fill_1 FILLER_25_129 ();
 sg13g2_decap_4 FILLER_25_135 ();
 sg13g2_decap_8 FILLER_25_147 ();
 sg13g2_fill_1 FILLER_25_154 ();
 sg13g2_fill_1 FILLER_25_161 ();
 sg13g2_decap_4 FILLER_25_181 ();
 sg13g2_fill_2 FILLER_25_203 ();
 sg13g2_fill_1 FILLER_25_205 ();
 sg13g2_fill_1 FILLER_25_222 ();
 sg13g2_fill_1 FILLER_25_244 ();
 sg13g2_fill_2 FILLER_25_255 ();
 sg13g2_decap_4 FILLER_25_298 ();
 sg13g2_fill_2 FILLER_25_302 ();
 sg13g2_decap_4 FILLER_25_349 ();
 sg13g2_fill_1 FILLER_25_353 ();
 sg13g2_fill_2 FILLER_25_381 ();
 sg13g2_fill_2 FILLER_25_395 ();
 sg13g2_fill_1 FILLER_26_0 ();
 sg13g2_fill_1 FILLER_26_15 ();
 sg13g2_fill_1 FILLER_26_29 ();
 sg13g2_fill_1 FILLER_26_35 ();
 sg13g2_fill_2 FILLER_26_46 ();
 sg13g2_fill_1 FILLER_26_48 ();
 sg13g2_fill_2 FILLER_26_65 ();
 sg13g2_fill_2 FILLER_26_77 ();
 sg13g2_fill_2 FILLER_26_89 ();
 sg13g2_fill_2 FILLER_26_128 ();
 sg13g2_fill_1 FILLER_26_140 ();
 sg13g2_fill_2 FILLER_26_154 ();
 sg13g2_decap_4 FILLER_26_175 ();
 sg13g2_fill_2 FILLER_26_187 ();
 sg13g2_decap_8 FILLER_26_199 ();
 sg13g2_decap_4 FILLER_26_206 ();
 sg13g2_fill_1 FILLER_26_210 ();
 sg13g2_fill_2 FILLER_26_227 ();
 sg13g2_fill_1 FILLER_26_229 ();
 sg13g2_fill_2 FILLER_26_292 ();
 sg13g2_decap_4 FILLER_26_303 ();
 sg13g2_fill_2 FILLER_26_330 ();
 sg13g2_fill_1 FILLER_26_332 ();
 sg13g2_fill_1 FILLER_26_374 ();
 sg13g2_decap_4 FILLER_27_0 ();
 sg13g2_fill_2 FILLER_27_4 ();
 sg13g2_fill_2 FILLER_27_32 ();
 sg13g2_fill_2 FILLER_27_68 ();
 sg13g2_fill_1 FILLER_27_81 ();
 sg13g2_decap_4 FILLER_27_99 ();
 sg13g2_fill_2 FILLER_27_111 ();
 sg13g2_fill_1 FILLER_27_113 ();
 sg13g2_fill_2 FILLER_27_124 ();
 sg13g2_fill_1 FILLER_27_132 ();
 sg13g2_fill_2 FILLER_27_155 ();
 sg13g2_fill_2 FILLER_27_167 ();
 sg13g2_fill_1 FILLER_27_169 ();
 sg13g2_fill_2 FILLER_27_181 ();
 sg13g2_fill_2 FILLER_27_188 ();
 sg13g2_fill_1 FILLER_27_190 ();
 sg13g2_fill_1 FILLER_27_200 ();
 sg13g2_fill_2 FILLER_27_224 ();
 sg13g2_fill_1 FILLER_27_242 ();
 sg13g2_fill_2 FILLER_27_284 ();
 sg13g2_fill_2 FILLER_27_291 ();
 sg13g2_fill_1 FILLER_27_298 ();
 sg13g2_decap_4 FILLER_27_308 ();
 sg13g2_fill_2 FILLER_27_312 ();
 sg13g2_decap_4 FILLER_27_323 ();
 sg13g2_fill_2 FILLER_27_390 ();
 sg13g2_fill_2 FILLER_27_407 ();
 sg13g2_fill_1 FILLER_28_14 ();
 sg13g2_fill_2 FILLER_28_41 ();
 sg13g2_fill_1 FILLER_28_78 ();
 sg13g2_fill_2 FILLER_28_88 ();
 sg13g2_fill_1 FILLER_28_90 ();
 sg13g2_fill_2 FILLER_28_110 ();
 sg13g2_fill_1 FILLER_28_112 ();
 sg13g2_fill_2 FILLER_28_118 ();
 sg13g2_fill_2 FILLER_28_134 ();
 sg13g2_fill_1 FILLER_28_141 ();
 sg13g2_fill_2 FILLER_28_159 ();
 sg13g2_fill_2 FILLER_28_174 ();
 sg13g2_fill_1 FILLER_28_190 ();
 sg13g2_decap_8 FILLER_28_215 ();
 sg13g2_fill_2 FILLER_28_252 ();
 sg13g2_fill_1 FILLER_28_254 ();
 sg13g2_fill_1 FILLER_28_295 ();
 sg13g2_decap_4 FILLER_28_301 ();
 sg13g2_fill_2 FILLER_28_305 ();
 sg13g2_fill_2 FILLER_28_334 ();
 sg13g2_decap_4 FILLER_28_345 ();
 sg13g2_fill_1 FILLER_28_349 ();
 sg13g2_fill_1 FILLER_28_375 ();
 sg13g2_fill_1 FILLER_28_408 ();
 sg13g2_fill_1 FILLER_29_48 ();
 sg13g2_fill_2 FILLER_29_62 ();
 sg13g2_fill_1 FILLER_29_64 ();
 sg13g2_fill_2 FILLER_29_70 ();
 sg13g2_fill_1 FILLER_29_87 ();
 sg13g2_decap_8 FILLER_29_94 ();
 sg13g2_fill_1 FILLER_29_105 ();
 sg13g2_fill_1 FILLER_29_112 ();
 sg13g2_fill_2 FILLER_29_192 ();
 sg13g2_fill_1 FILLER_29_194 ();
 sg13g2_fill_1 FILLER_29_208 ();
 sg13g2_fill_2 FILLER_29_219 ();
 sg13g2_fill_1 FILLER_29_221 ();
 sg13g2_fill_1 FILLER_29_240 ();
 sg13g2_decap_8 FILLER_29_301 ();
 sg13g2_fill_1 FILLER_29_317 ();
 sg13g2_fill_2 FILLER_29_332 ();
 sg13g2_fill_1 FILLER_29_334 ();
 sg13g2_fill_1 FILLER_29_353 ();
 sg13g2_fill_1 FILLER_29_382 ();
 sg13g2_fill_1 FILLER_30_18 ();
 sg13g2_fill_2 FILLER_30_45 ();
 sg13g2_fill_2 FILLER_30_63 ();
 sg13g2_fill_2 FILLER_30_105 ();
 sg13g2_decap_4 FILLER_30_125 ();
 sg13g2_fill_1 FILLER_30_139 ();
 sg13g2_fill_2 FILLER_30_149 ();
 sg13g2_fill_1 FILLER_30_151 ();
 sg13g2_fill_2 FILLER_30_157 ();
 sg13g2_fill_1 FILLER_30_176 ();
 sg13g2_fill_2 FILLER_30_182 ();
 sg13g2_fill_2 FILLER_30_199 ();
 sg13g2_fill_2 FILLER_30_280 ();
 sg13g2_fill_2 FILLER_30_300 ();
 sg13g2_fill_1 FILLER_30_302 ();
 sg13g2_fill_1 FILLER_30_373 ();
 sg13g2_fill_2 FILLER_31_0 ();
 sg13g2_fill_2 FILLER_31_31 ();
 sg13g2_fill_2 FILLER_31_57 ();
 sg13g2_fill_1 FILLER_31_59 ();
 sg13g2_fill_1 FILLER_31_65 ();
 sg13g2_fill_1 FILLER_31_75 ();
 sg13g2_fill_1 FILLER_31_86 ();
 sg13g2_fill_1 FILLER_31_97 ();
 sg13g2_fill_2 FILLER_31_114 ();
 sg13g2_fill_2 FILLER_31_145 ();
 sg13g2_fill_1 FILLER_31_147 ();
 sg13g2_fill_2 FILLER_31_164 ();
 sg13g2_fill_2 FILLER_31_184 ();
 sg13g2_fill_1 FILLER_31_186 ();
 sg13g2_fill_2 FILLER_31_208 ();
 sg13g2_fill_1 FILLER_31_210 ();
 sg13g2_fill_2 FILLER_31_221 ();
 sg13g2_fill_1 FILLER_31_260 ();
 sg13g2_fill_1 FILLER_31_371 ();
 sg13g2_fill_1 FILLER_31_382 ();
 sg13g2_fill_2 FILLER_32_45 ();
 sg13g2_fill_1 FILLER_32_91 ();
 sg13g2_decap_8 FILLER_32_96 ();
 sg13g2_fill_1 FILLER_32_103 ();
 sg13g2_fill_2 FILLER_32_123 ();
 sg13g2_fill_1 FILLER_32_152 ();
 sg13g2_fill_1 FILLER_32_161 ();
 sg13g2_fill_2 FILLER_32_166 ();
 sg13g2_fill_1 FILLER_32_168 ();
 sg13g2_fill_2 FILLER_32_178 ();
 sg13g2_fill_1 FILLER_32_180 ();
 sg13g2_fill_2 FILLER_32_185 ();
 sg13g2_fill_2 FILLER_32_197 ();
 sg13g2_fill_2 FILLER_32_239 ();
 sg13g2_fill_1 FILLER_32_272 ();
 sg13g2_fill_2 FILLER_32_288 ();
 sg13g2_fill_2 FILLER_32_304 ();
 sg13g2_fill_1 FILLER_32_306 ();
 sg13g2_fill_2 FILLER_33_0 ();
 sg13g2_fill_1 FILLER_33_2 ();
 sg13g2_fill_1 FILLER_33_67 ();
 sg13g2_fill_1 FILLER_33_112 ();
 sg13g2_fill_1 FILLER_33_139 ();
 sg13g2_fill_2 FILLER_33_150 ();
 sg13g2_fill_1 FILLER_33_192 ();
 sg13g2_fill_2 FILLER_33_223 ();
 sg13g2_fill_1 FILLER_33_225 ();
 sg13g2_fill_1 FILLER_33_282 ();
 sg13g2_fill_2 FILLER_33_308 ();
 sg13g2_fill_2 FILLER_33_329 ();
 sg13g2_fill_1 FILLER_33_331 ();
 sg13g2_fill_2 FILLER_33_354 ();
 sg13g2_fill_1 FILLER_33_396 ();
 sg13g2_fill_1 FILLER_34_79 ();
 sg13g2_fill_1 FILLER_34_90 ();
 sg13g2_fill_2 FILLER_34_105 ();
 sg13g2_fill_2 FILLER_34_116 ();
 sg13g2_fill_2 FILLER_34_122 ();
 sg13g2_decap_8 FILLER_34_137 ();
 sg13g2_fill_1 FILLER_34_175 ();
 sg13g2_fill_2 FILLER_34_185 ();
 sg13g2_fill_1 FILLER_34_187 ();
 sg13g2_fill_2 FILLER_34_193 ();
 sg13g2_fill_2 FILLER_34_205 ();
 sg13g2_fill_2 FILLER_34_224 ();
 sg13g2_fill_1 FILLER_34_306 ();
 sg13g2_fill_1 FILLER_34_325 ();
 sg13g2_fill_2 FILLER_35_0 ();
 sg13g2_fill_2 FILLER_35_64 ();
 sg13g2_fill_1 FILLER_35_66 ();
 sg13g2_fill_2 FILLER_35_99 ();
 sg13g2_fill_2 FILLER_35_146 ();
 sg13g2_fill_2 FILLER_35_175 ();
 sg13g2_fill_1 FILLER_35_177 ();
 sg13g2_fill_2 FILLER_35_196 ();
 sg13g2_fill_2 FILLER_35_248 ();
 sg13g2_fill_2 FILLER_35_278 ();
 sg13g2_fill_1 FILLER_35_280 ();
 sg13g2_fill_2 FILLER_35_407 ();
 sg13g2_fill_1 FILLER_36_50 ();
 sg13g2_fill_2 FILLER_36_121 ();
 sg13g2_decap_8 FILLER_36_132 ();
 sg13g2_fill_2 FILLER_36_170 ();
 sg13g2_fill_1 FILLER_36_172 ();
 sg13g2_fill_2 FILLER_36_196 ();
 sg13g2_fill_1 FILLER_36_198 ();
 sg13g2_fill_1 FILLER_36_204 ();
 sg13g2_fill_1 FILLER_36_291 ();
 sg13g2_fill_2 FILLER_36_310 ();
 sg13g2_fill_2 FILLER_36_329 ();
 sg13g2_fill_1 FILLER_36_345 ();
 sg13g2_fill_2 FILLER_36_381 ();
 sg13g2_fill_2 FILLER_37_0 ();
 sg13g2_fill_1 FILLER_37_2 ();
 sg13g2_fill_2 FILLER_37_59 ();
 sg13g2_fill_1 FILLER_37_61 ();
 sg13g2_fill_2 FILLER_37_84 ();
 sg13g2_fill_2 FILLER_37_95 ();
 sg13g2_fill_2 FILLER_37_122 ();
 sg13g2_fill_1 FILLER_37_124 ();
 sg13g2_fill_2 FILLER_37_221 ();
 sg13g2_fill_1 FILLER_37_255 ();
 sg13g2_fill_1 FILLER_37_362 ();
 sg13g2_fill_1 FILLER_37_408 ();
 sg13g2_fill_1 FILLER_38_70 ();
 sg13g2_decap_4 FILLER_38_101 ();
 sg13g2_decap_4 FILLER_38_118 ();
 sg13g2_fill_1 FILLER_38_122 ();
 sg13g2_fill_1 FILLER_38_154 ();
 sg13g2_fill_1 FILLER_38_176 ();
 sg13g2_fill_2 FILLER_38_199 ();
 sg13g2_fill_1 FILLER_38_201 ();
 sg13g2_fill_2 FILLER_38_229 ();
 sg13g2_fill_1 FILLER_38_231 ();
 sg13g2_fill_2 FILLER_38_246 ();
endmodule

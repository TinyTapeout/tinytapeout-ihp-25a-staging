module tt_um_dendraws_donut (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire _3093_;
 wire _3094_;
 wire _3095_;
 wire _3096_;
 wire _3097_;
 wire _3098_;
 wire _3099_;
 wire _3100_;
 wire _3101_;
 wire _3102_;
 wire _3103_;
 wire _3104_;
 wire _3105_;
 wire _3106_;
 wire _3107_;
 wire _3108_;
 wire _3109_;
 wire _3110_;
 wire _3111_;
 wire _3112_;
 wire _3113_;
 wire _3114_;
 wire _3115_;
 wire _3116_;
 wire _3117_;
 wire _3118_;
 wire _3119_;
 wire _3120_;
 wire _3121_;
 wire _3122_;
 wire _3123_;
 wire _3124_;
 wire _3125_;
 wire _3126_;
 wire _3127_;
 wire _3128_;
 wire _3129_;
 wire _3130_;
 wire _3131_;
 wire _3132_;
 wire _3133_;
 wire _3134_;
 wire _3135_;
 wire _3136_;
 wire _3137_;
 wire _3138_;
 wire _3139_;
 wire _3140_;
 wire _3141_;
 wire _3142_;
 wire _3143_;
 wire _3144_;
 wire _3145_;
 wire _3146_;
 wire _3147_;
 wire _3148_;
 wire _3149_;
 wire _3150_;
 wire _3151_;
 wire _3152_;
 wire _3153_;
 wire _3154_;
 wire _3155_;
 wire _3156_;
 wire _3157_;
 wire _3158_;
 wire _3159_;
 wire _3160_;
 wire _3161_;
 wire _3162_;
 wire _3163_;
 wire _3164_;
 wire _3165_;
 wire _3166_;
 wire _3167_;
 wire _3168_;
 wire _3169_;
 wire _3170_;
 wire _3171_;
 wire _3172_;
 wire _3173_;
 wire _3174_;
 wire _3175_;
 wire _3176_;
 wire _3177_;
 wire _3178_;
 wire _3179_;
 wire _3180_;
 wire _3181_;
 wire _3182_;
 wire _3183_;
 wire _3184_;
 wire _3185_;
 wire _3186_;
 wire _3187_;
 wire _3188_;
 wire _3189_;
 wire _3190_;
 wire _3191_;
 wire _3192_;
 wire _3193_;
 wire _3194_;
 wire _3195_;
 wire _3196_;
 wire _3197_;
 wire _3198_;
 wire _3199_;
 wire _3200_;
 wire _3201_;
 wire _3202_;
 wire _3203_;
 wire _3204_;
 wire _3205_;
 wire _3206_;
 wire _3207_;
 wire _3208_;
 wire _3209_;
 wire _3210_;
 wire _3211_;
 wire _3212_;
 wire _3213_;
 wire _3214_;
 wire _3215_;
 wire _3216_;
 wire _3217_;
 wire _3218_;
 wire _3219_;
 wire _3220_;
 wire _3221_;
 wire _3222_;
 wire _3223_;
 wire _3224_;
 wire _3225_;
 wire _3226_;
 wire _3227_;
 wire _3228_;
 wire _3229_;
 wire _3230_;
 wire _3231_;
 wire _3232_;
 wire _3233_;
 wire _3234_;
 wire _3235_;
 wire _3236_;
 wire _3237_;
 wire _3238_;
 wire _3239_;
 wire _3240_;
 wire _3241_;
 wire _3242_;
 wire _3243_;
 wire _3244_;
 wire _3245_;
 wire _3246_;
 wire _3247_;
 wire _3248_;
 wire _3249_;
 wire _3250_;
 wire _3251_;
 wire _3252_;
 wire _3253_;
 wire _3254_;
 wire _3255_;
 wire _3256_;
 wire _3257_;
 wire _3258_;
 wire _3259_;
 wire _3260_;
 wire _3261_;
 wire _3262_;
 wire _3263_;
 wire _3264_;
 wire _3265_;
 wire _3266_;
 wire _3267_;
 wire _3268_;
 wire _3269_;
 wire _3270_;
 wire _3271_;
 wire _3272_;
 wire _3273_;
 wire _3274_;
 wire _3275_;
 wire _3276_;
 wire _3277_;
 wire _3278_;
 wire _3279_;
 wire _3280_;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire clknet_0_clk;
 wire hsync;
 wire \hvsync_gen.hpos[0] ;
 wire \hvsync_gen.hpos[1] ;
 wire \hvsync_gen.hpos[2] ;
 wire \hvsync_gen.hpos[3] ;
 wire \hvsync_gen.hpos[4] ;
 wire \hvsync_gen.hpos[5] ;
 wire \hvsync_gen.hpos[6] ;
 wire \hvsync_gen.hpos[7] ;
 wire \hvsync_gen.hpos[8] ;
 wire \hvsync_gen.hpos[9] ;
 wire \hvsync_gen.phase ;
 wire \hvsync_gen.vpos[0] ;
 wire \hvsync_gen.vpos[1] ;
 wire \hvsync_gen.vpos[2] ;
 wire \hvsync_gen.vpos[3] ;
 wire \hvsync_gen.vpos[4] ;
 wire \hvsync_gen.vpos[5] ;
 wire \hvsync_gen.vpos[6] ;
 wire \hvsync_gen.vpos[7] ;
 wire \hvsync_gen.vpos[8] ;
 wire \hvsync_gen.vpos[9] ;
 wire \hvsync_gen.vsync ;
 wire i_phase_0;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net1;
 wire net2;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;

 sg13g2_inv_1 _3303_ (.Y(_2971_),
    .A(\hvsync_gen.vpos[9] ));
 sg13g2_inv_4 _3304_ (.A(net563),
    .Y(_2982_));
 sg13g2_inv_2 _3305_ (.Y(_2993_),
    .A(\hvsync_gen.vpos[7] ));
 sg13g2_inv_4 _3306_ (.A(\hvsync_gen.vpos[6] ),
    .Y(_3004_));
 sg13g2_inv_1 _3307_ (.Y(_3015_),
    .A(net567));
 sg13g2_inv_1 _3308_ (.Y(_3026_),
    .A(net569));
 sg13g2_inv_2 _3309_ (.Y(_3037_),
    .A(net572));
 sg13g2_inv_2 _3310_ (.Y(_3048_),
    .A(net583));
 sg13g2_inv_1 _3311_ (.Y(_3059_),
    .A(net553));
 sg13g2_inv_1 _3312_ (.Y(_3070_),
    .A(net584));
 sg13g2_inv_1 _3313_ (.Y(_3081_),
    .A(net588));
 sg13g2_inv_2 _3314_ (.Y(_3092_),
    .A(net591));
 sg13g2_inv_1 _3315_ (.Y(_3103_),
    .A(net597));
 sg13g2_inv_1 _3316_ (.Y(_3114_),
    .A(\hvsync_gen.hpos[3] ));
 sg13g2_inv_2 _3317_ (.Y(_3125_),
    .A(_0019_));
 sg13g2_inv_2 _3318_ (.Y(_3136_),
    .A(_0003_));
 sg13g2_inv_4 _3319_ (.A(_0002_),
    .Y(_3147_));
 sg13g2_inv_2 _3320_ (.Y(_3158_),
    .A(net562));
 sg13g2_inv_2 _3321_ (.Y(_3169_),
    .A(_0007_));
 sg13g2_inv_1 _3322_ (.Y(_3180_),
    .A(net589));
 sg13g2_inv_2 _3323_ (.Y(_3191_),
    .A(_0015_));
 sg13g2_inv_2 _3324_ (.Y(_3202_),
    .A(_0016_));
 sg13g2_inv_1 _3325_ (.Y(_3213_),
    .A(_0000_));
 sg13g2_inv_2 _3326_ (.Y(_3224_),
    .A(_0001_));
 sg13g2_inv_4 _3327_ (.A(_0010_),
    .Y(_3235_));
 sg13g2_inv_1 _3328_ (.Y(_3246_),
    .A(_0011_));
 sg13g2_inv_2 _3329_ (.Y(_3257_),
    .A(net41));
 sg13g2_inv_1 _3330_ (.Y(_3268_),
    .A(net1));
 sg13g2_nand2_1 _3331_ (.Y(_0042_),
    .A(net582),
    .B(net586));
 sg13g2_nor2_2 _3332_ (.A(net594),
    .B(net597),
    .Y(_0053_));
 sg13g2_or2_2 _3333_ (.X(_0064_),
    .B(\hvsync_gen.hpos[4] ),
    .A(\hvsync_gen.hpos[5] ));
 sg13g2_or3_1 _3334_ (.A(net590),
    .B(net593),
    .C(net596),
    .X(_0075_));
 sg13g2_nand3_1 _3335_ (.B(net587),
    .C(_0075_),
    .A(net582),
    .Y(_0086_));
 sg13g2_nand2_2 _3336_ (.Y(_0097_),
    .A(net595),
    .B(net597));
 sg13g2_nor2_2 _3337_ (.A(net537),
    .B(_3092_),
    .Y(_0108_));
 sg13g2_nand2_1 _3338_ (.Y(_0119_),
    .A(net587),
    .B(net590));
 sg13g2_or2_1 _3339_ (.X(_0130_),
    .B(_0119_),
    .A(_0097_));
 sg13g2_nand3_1 _3340_ (.B(_3070_),
    .C(_0130_),
    .A(net582),
    .Y(_0141_));
 sg13g2_a22oi_1 _3341_ (.Y(hsync),
    .B1(_0141_),
    .B2(_3125_),
    .A2(_0086_),
    .A1(_0042_));
 sg13g2_nor2_2 _3342_ (.A(_2993_),
    .B(_3004_),
    .Y(_0162_));
 sg13g2_nand2_1 _3343_ (.Y(_0173_),
    .A(\hvsync_gen.vpos[6] ),
    .B(net567));
 sg13g2_nor2_2 _3344_ (.A(_2993_),
    .B(_0173_),
    .Y(_0184_));
 sg13g2_nand2_1 _3345_ (.Y(_0195_),
    .A(net565),
    .B(_0162_));
 sg13g2_nor2_1 _3346_ (.A(net569),
    .B(_0195_),
    .Y(_0206_));
 sg13g2_nor2_1 _3347_ (.A(\hvsync_gen.vpos[9] ),
    .B(_2982_),
    .Y(_0217_));
 sg13g2_nor2_1 _3348_ (.A(_3037_),
    .B(net574),
    .Y(_0228_));
 sg13g2_and4_1 _3349_ (.A(net576),
    .B(_0206_),
    .C(_0217_),
    .D(_0228_),
    .X(\hvsync_gen.vsync ));
 sg13g2_nor2_2 _3350_ (.A(\hvsync_gen.vpos[7] ),
    .B(\hvsync_gen.vpos[6] ),
    .Y(_0249_));
 sg13g2_inv_1 _3351_ (.Y(_0260_),
    .A(_0249_));
 sg13g2_o21ai_1 _3352_ (.B1(net571),
    .Y(_0271_),
    .A1(net575),
    .A2(net576));
 sg13g2_o21ai_1 _3353_ (.B1(_0003_),
    .Y(_0282_),
    .A1(net569),
    .A2(net536));
 sg13g2_nor2_1 _3354_ (.A(net566),
    .B(_0282_),
    .Y(_0293_));
 sg13g2_nand3_1 _3355_ (.B(_0249_),
    .C(_0293_),
    .A(_2982_),
    .Y(_0304_));
 sg13g2_nor2_2 _3356_ (.A(net563),
    .B(net557),
    .Y(_0315_));
 sg13g2_nor4_2 _3357_ (.A(net565),
    .B(net556),
    .C(_0260_),
    .Y(_0326_),
    .D(_0282_));
 sg13g2_o21ai_1 _3358_ (.B1(_0304_),
    .Y(_0337_),
    .A1(_0315_),
    .A2(_0326_));
 sg13g2_nor2_2 _3359_ (.A(net565),
    .B(net569),
    .Y(_0348_));
 sg13g2_or2_1 _3360_ (.X(_0359_),
    .B(net568),
    .A(net567));
 sg13g2_nor2_2 _3361_ (.A(net576),
    .B(net581),
    .Y(_0370_));
 sg13g2_or2_1 _3362_ (.X(_0381_),
    .B(net579),
    .A(net576));
 sg13g2_o21ai_1 _3363_ (.B1(net574),
    .Y(_0392_),
    .A1(net577),
    .A2(net581));
 sg13g2_and2_1 _3364_ (.A(net572),
    .B(net575),
    .X(_0403_));
 sg13g2_nand2_2 _3365_ (.Y(_0414_),
    .A(net571),
    .B(net574));
 sg13g2_a21oi_2 _3366_ (.B1(_0359_),
    .Y(_0425_),
    .A2(_0403_),
    .A1(_0381_));
 sg13g2_o21ai_1 _3367_ (.B1(_0348_),
    .Y(_0436_),
    .A1(_0370_),
    .A2(_0414_));
 sg13g2_nand2_1 _3368_ (.Y(_0447_),
    .A(_0162_),
    .B(_0436_));
 sg13g2_xnor2_1 _3369_ (.Y(_0458_),
    .A(_3158_),
    .B(_0447_));
 sg13g2_o21ai_1 _3370_ (.B1(_0337_),
    .Y(_0469_),
    .A1(net544),
    .A2(_0458_));
 sg13g2_a21oi_1 _3371_ (.A1(_0162_),
    .A2(_0436_),
    .Y(_0480_),
    .B1(net564));
 sg13g2_nand2_1 _3372_ (.Y(_0491_),
    .A(net563),
    .B(net556));
 sg13g2_nor3_2 _3373_ (.A(_0315_),
    .B(_0326_),
    .C(_0480_),
    .Y(_0502_));
 sg13g2_xnor2_1 _3374_ (.Y(_0513_),
    .A(_3147_),
    .B(_0502_));
 sg13g2_xnor2_1 _3375_ (.Y(_0524_),
    .A(_0002_),
    .B(_0502_));
 sg13g2_nand2_1 _3376_ (.Y(_0535_),
    .A(_3004_),
    .B(net557));
 sg13g2_nor2b_1 _3377_ (.A(net569),
    .B_N(net556),
    .Y(_0546_));
 sg13g2_o21ai_1 _3378_ (.B1(_0546_),
    .Y(_0557_),
    .A1(_0370_),
    .A2(_0414_));
 sg13g2_nand2_1 _3379_ (.Y(_0568_),
    .A(net556),
    .B(_0425_));
 sg13g2_a22oi_1 _3380_ (.Y(_0579_),
    .B1(_0535_),
    .B2(_0568_),
    .A2(_0425_),
    .A1(_3004_));
 sg13g2_o21ai_1 _3381_ (.B1(_0007_),
    .Y(_0590_),
    .A1(net566),
    .A2(_0282_));
 sg13g2_or3_1 _3382_ (.A(net566),
    .B(_0007_),
    .C(_0282_),
    .X(_0601_));
 sg13g2_and3_1 _3383_ (.X(_0612_),
    .A(net544),
    .B(_0590_),
    .C(_0601_));
 sg13g2_nor2_1 _3384_ (.A(_0579_),
    .B(_0612_),
    .Y(_0623_));
 sg13g2_o21ai_1 _3385_ (.B1(_0557_),
    .Y(_0634_),
    .A1(net556),
    .A2(_0282_));
 sg13g2_xnor2_1 _3386_ (.Y(_0645_),
    .A(_0008_),
    .B(_0634_));
 sg13g2_nand2_2 _3387_ (.Y(_0656_),
    .A(net581),
    .B(net558));
 sg13g2_or2_1 _3388_ (.X(_0667_),
    .B(net558),
    .A(net581));
 sg13g2_nand2_2 _3389_ (.Y(_0678_),
    .A(_0656_),
    .B(_0667_));
 sg13g2_nor2b_2 _3390_ (.A(net576),
    .B_N(net579),
    .Y(_0689_));
 sg13g2_nand2b_1 _3391_ (.Y(_0700_),
    .B(net577),
    .A_N(net581));
 sg13g2_xnor2_1 _3392_ (.Y(_0711_),
    .A(net577),
    .B(net581));
 sg13g2_nor2_1 _3393_ (.A(net577),
    .B(net558),
    .Y(_0722_));
 sg13g2_a21oi_1 _3394_ (.A1(net558),
    .A2(_0711_),
    .Y(_0733_),
    .B1(_0722_));
 sg13g2_a221oi_1 _3395_ (.B2(net558),
    .C1(_0722_),
    .B1(_0711_),
    .A1(_0656_),
    .Y(_0744_),
    .A2(_0667_));
 sg13g2_nor3_2 _3396_ (.A(net574),
    .B(net577),
    .C(net581),
    .Y(_0755_));
 sg13g2_xnor2_1 _3397_ (.Y(_0766_),
    .A(net575),
    .B(_0370_));
 sg13g2_xor2_1 _3398_ (.B(net577),
    .A(net574),
    .X(_0777_));
 sg13g2_nand3b_1 _3399_ (.B(net559),
    .C(_0392_),
    .Y(_0788_),
    .A_N(_0755_));
 sg13g2_or2_1 _3400_ (.X(_0799_),
    .B(_0777_),
    .A(net559));
 sg13g2_nand2_1 _3401_ (.Y(_0810_),
    .A(_0788_),
    .B(_0799_));
 sg13g2_and3_1 _3402_ (.X(_0821_),
    .A(_0744_),
    .B(_0788_),
    .C(_0799_));
 sg13g2_or3_2 _3403_ (.A(net571),
    .B(net574),
    .C(net577),
    .X(_0832_));
 sg13g2_nand2_1 _3404_ (.Y(_0843_),
    .A(net536),
    .B(_0832_));
 sg13g2_xnor2_1 _3405_ (.Y(_0854_),
    .A(_0009_),
    .B(_0392_));
 sg13g2_mux2_2 _3406_ (.A0(_0843_),
    .A1(_0854_),
    .S(net558),
    .X(_0865_));
 sg13g2_nand2_1 _3407_ (.Y(_0876_),
    .A(_3026_),
    .B(_0271_));
 sg13g2_or2_1 _3408_ (.X(_0887_),
    .B(net536),
    .A(_3026_));
 sg13g2_a21o_1 _3409_ (.A2(_0887_),
    .A1(_0876_),
    .B1(net555),
    .X(_0898_));
 sg13g2_nor3_1 _3410_ (.A(_0003_),
    .B(_0370_),
    .C(_0414_),
    .Y(_0909_));
 sg13g2_a21oi_1 _3411_ (.A1(_0381_),
    .A2(_0403_),
    .Y(_0920_),
    .B1(_3136_));
 sg13g2_o21ai_1 _3412_ (.B1(net555),
    .Y(_0931_),
    .A1(_0909_),
    .A2(_0920_));
 sg13g2_and2_1 _3413_ (.A(_0898_),
    .B(_0931_),
    .X(_0942_));
 sg13g2_and4_1 _3414_ (.A(_0821_),
    .B(_0865_),
    .C(_0898_),
    .D(_0931_),
    .X(_0953_));
 sg13g2_nand4_1 _3415_ (.B(_0865_),
    .C(_0898_),
    .A(_0821_),
    .Y(_0964_),
    .D(_0931_));
 sg13g2_nand2b_1 _3416_ (.Y(_0975_),
    .B(_0953_),
    .A_N(_0645_));
 sg13g2_nor4_2 _3417_ (.A(_0579_),
    .B(_0612_),
    .C(_0645_),
    .Y(_0986_),
    .D(_0964_));
 sg13g2_nor2_1 _3418_ (.A(_3004_),
    .B(net557),
    .Y(_0997_));
 sg13g2_xor2_1 _3419_ (.B(net556),
    .A(\hvsync_gen.vpos[6] ),
    .X(_1008_));
 sg13g2_a21oi_1 _3420_ (.A1(net556),
    .A2(_0425_),
    .Y(_1019_),
    .B1(_1008_));
 sg13g2_o21ai_1 _3421_ (.B1(_1019_),
    .Y(_1030_),
    .A1(\hvsync_gen.vpos[6] ),
    .A2(_0293_));
 sg13g2_xor2_1 _3422_ (.B(_1030_),
    .A(_0005_),
    .X(_1041_));
 sg13g2_xnor2_1 _3423_ (.Y(_1052_),
    .A(_0005_),
    .B(_1030_));
 sg13g2_nand2_1 _3424_ (.Y(_1063_),
    .A(_0986_),
    .B(_1052_));
 sg13g2_a21o_1 _3425_ (.A2(_1052_),
    .A1(_0986_),
    .B1(_0524_),
    .X(_1074_));
 sg13g2_mux2_1 _3426_ (.A0(_0513_),
    .A1(_1074_),
    .S(_0469_),
    .X(_1085_));
 sg13g2_inv_2 _3427_ (.Y(_1096_),
    .A(_1085_));
 sg13g2_nand3b_1 _3428_ (.B(_1052_),
    .C(_0513_),
    .Y(_1107_),
    .A_N(_0986_));
 sg13g2_o21ai_1 _3429_ (.B1(_1041_),
    .Y(_1118_),
    .A1(_0524_),
    .A2(_0986_));
 sg13g2_nand2_1 _3430_ (.Y(_1129_),
    .A(_1107_),
    .B(_1118_));
 sg13g2_nand3_1 _3431_ (.B(_0623_),
    .C(_0975_),
    .A(_0513_),
    .Y(_1140_));
 sg13g2_a21o_1 _3432_ (.A2(_0975_),
    .A1(_0513_),
    .B1(_0623_),
    .X(_1151_));
 sg13g2_and2_1 _3433_ (.A(_1140_),
    .B(_1151_),
    .X(_1162_));
 sg13g2_nand4_1 _3434_ (.B(_1118_),
    .C(_1140_),
    .A(_1107_),
    .Y(_1173_),
    .D(_1151_));
 sg13g2_nor2b_2 _3435_ (.A(net520),
    .B_N(_1173_),
    .Y(_1184_));
 sg13g2_nand2_1 _3436_ (.Y(_1195_),
    .A(_1096_),
    .B(_1173_));
 sg13g2_nor2_1 _3437_ (.A(net520),
    .B(_1173_),
    .Y(_1206_));
 sg13g2_nand2_2 _3438_ (.Y(_1217_),
    .A(_1096_),
    .B(_1195_));
 sg13g2_nor2_1 _3439_ (.A(_0524_),
    .B(_0953_),
    .Y(_1228_));
 sg13g2_xnor2_1 _3440_ (.Y(_1239_),
    .A(_0645_),
    .B(_1228_));
 sg13g2_xor2_1 _3441_ (.B(_1228_),
    .A(_0645_),
    .X(_1250_));
 sg13g2_nor2_1 _3442_ (.A(_1217_),
    .B(_1250_),
    .Y(_1261_));
 sg13g2_nand2_2 _3443_ (.Y(_1272_),
    .A(net519),
    .B(_1239_));
 sg13g2_nand2_1 _3444_ (.Y(_1283_),
    .A(_1096_),
    .B(_1129_));
 sg13g2_a21oi_1 _3445_ (.A1(_0821_),
    .A2(_0865_),
    .Y(_1294_),
    .B1(_0524_));
 sg13g2_xnor2_1 _3446_ (.Y(_1305_),
    .A(_0942_),
    .B(_1294_));
 sg13g2_nor2_1 _3447_ (.A(_0524_),
    .B(_0744_),
    .Y(_1316_));
 sg13g2_xnor2_1 _3448_ (.Y(_1327_),
    .A(_0810_),
    .B(_1316_));
 sg13g2_nor2_1 _3449_ (.A(_0524_),
    .B(_0678_),
    .Y(_1338_));
 sg13g2_xnor2_1 _3450_ (.Y(_1349_),
    .A(_0733_),
    .B(_1338_));
 sg13g2_nor2_1 _3451_ (.A(_0524_),
    .B(_0821_),
    .Y(_1360_));
 sg13g2_xnor2_1 _3452_ (.Y(_1371_),
    .A(_0865_),
    .B(_1360_));
 sg13g2_inv_1 _3453_ (.Y(_1382_),
    .A(_1371_));
 sg13g2_a21o_1 _3454_ (.A2(_1349_),
    .A1(_1327_),
    .B1(_1371_),
    .X(_1393_));
 sg13g2_nor3_1 _3455_ (.A(net520),
    .B(_1173_),
    .C(_1305_),
    .Y(_1404_));
 sg13g2_nand2b_1 _3456_ (.Y(_1415_),
    .B(net519),
    .A_N(_1305_));
 sg13g2_nor3_2 _3457_ (.A(_0469_),
    .B(_0524_),
    .C(_1063_),
    .Y(_1426_));
 sg13g2_a221oi_1 _3458_ (.B2(_1404_),
    .C1(_1426_),
    .B1(_1393_),
    .A1(net519),
    .Y(_1437_),
    .A2(_1250_));
 sg13g2_nand2_2 _3459_ (.Y(_1448_),
    .A(net513),
    .B(_1437_));
 sg13g2_mux2_1 _3460_ (.A0(_1239_),
    .A1(_1162_),
    .S(_1448_),
    .X(_1459_));
 sg13g2_nor2_1 _3461_ (.A(_1250_),
    .B(_1305_),
    .Y(_1470_));
 sg13g2_o21ai_1 _3462_ (.B1(net514),
    .Y(_1481_),
    .A1(net520),
    .A2(_1470_));
 sg13g2_o21ai_1 _3463_ (.B1(_1415_),
    .Y(_1492_),
    .A1(_1096_),
    .A2(_1129_));
 sg13g2_a21o_2 _3464_ (.A2(_1459_),
    .A1(_1184_),
    .B1(_1492_),
    .X(_1503_));
 sg13g2_mux2_1 _3465_ (.A0(_1305_),
    .A1(_1250_),
    .S(_1448_),
    .X(_1514_));
 sg13g2_nor2_1 _3466_ (.A(_1217_),
    .B(_1382_),
    .Y(_1525_));
 sg13g2_a21oi_1 _3467_ (.A1(_1327_),
    .A2(_1382_),
    .Y(_1536_),
    .B1(net520));
 sg13g2_nor2_1 _3468_ (.A(_1481_),
    .B(_1536_),
    .Y(_1547_));
 sg13g2_nand2_1 _3469_ (.Y(_1558_),
    .A(_1162_),
    .B(net513));
 sg13g2_a21o_1 _3470_ (.A2(_1558_),
    .A1(_1547_),
    .B1(_1525_),
    .X(_1569_));
 sg13g2_a21oi_2 _3471_ (.B1(_1569_),
    .Y(_1580_),
    .A2(_1514_),
    .A1(_1184_));
 sg13g2_a21o_2 _3472_ (.A2(_1514_),
    .A1(_1184_),
    .B1(_1569_),
    .X(_1591_));
 sg13g2_nor2_1 _3473_ (.A(_1217_),
    .B(_1327_),
    .Y(_1602_));
 sg13g2_a21oi_1 _3474_ (.A1(net513),
    .A2(_1437_),
    .Y(_1613_),
    .B1(_1305_));
 sg13g2_o21ai_1 _3475_ (.B1(_1184_),
    .Y(_1624_),
    .A1(_1371_),
    .A2(_1448_));
 sg13g2_a21oi_1 _3476_ (.A1(net513),
    .A2(_1437_),
    .Y(_1635_),
    .B1(_1327_));
 sg13g2_nand3_1 _3477_ (.B(_1349_),
    .C(_1437_),
    .A(net513),
    .Y(_1646_));
 sg13g2_nand2_1 _3478_ (.Y(_1657_),
    .A(_1481_),
    .B(_1646_));
 sg13g2_a21oi_1 _3479_ (.A1(_1470_),
    .A2(_1536_),
    .Y(_1668_),
    .B1(_1184_));
 sg13g2_o21ai_1 _3480_ (.B1(_1668_),
    .Y(_1679_),
    .A1(_1635_),
    .A2(_1657_));
 sg13g2_o21ai_1 _3481_ (.B1(_1679_),
    .Y(_1690_),
    .A1(_1613_),
    .A2(_1624_));
 sg13g2_a21oi_1 _3482_ (.A1(_1459_),
    .A2(_1547_),
    .Y(_1701_),
    .B1(net519));
 sg13g2_a21oi_2 _3483_ (.B1(_1602_),
    .Y(_1712_),
    .A2(_1701_),
    .A1(_1690_));
 sg13g2_o21ai_1 _3484_ (.B1(_1580_),
    .Y(_1723_),
    .A1(_1503_),
    .A2(net486));
 sg13g2_nand2b_1 _3485_ (.Y(_1734_),
    .B(_1591_),
    .A_N(_1503_));
 sg13g2_xnor2_1 _3486_ (.Y(_1745_),
    .A(_1272_),
    .B(_1734_));
 sg13g2_nand2_1 _3487_ (.Y(_1756_),
    .A(_1723_),
    .B(_1745_));
 sg13g2_a21oi_1 _3488_ (.A1(net513),
    .A2(_1437_),
    .Y(_1767_),
    .B1(_1371_));
 sg13g2_and3_1 _3489_ (.X(_1778_),
    .A(net513),
    .B(_1327_),
    .C(_1437_));
 sg13g2_nor3_1 _3490_ (.A(net514),
    .B(_1767_),
    .C(_1778_),
    .Y(_1789_));
 sg13g2_a221oi_1 _3491_ (.B2(net520),
    .C1(_1789_),
    .B1(_1514_),
    .A1(net519),
    .Y(_1800_),
    .A2(_1349_));
 sg13g2_nor2_1 _3492_ (.A(_1261_),
    .B(net486),
    .Y(_1811_));
 sg13g2_or2_2 _3493_ (.X(_1822_),
    .B(_1800_),
    .A(_1261_));
 sg13g2_nor3_2 _3494_ (.A(_1503_),
    .B(net486),
    .C(_1822_),
    .Y(_1833_));
 sg13g2_nand2_2 _3495_ (.Y(_1844_),
    .A(_0678_),
    .B(net519));
 sg13g2_nand2_1 _3496_ (.Y(_1855_),
    .A(_1272_),
    .B(_1844_));
 sg13g2_nor2b_1 _3497_ (.A(_1503_),
    .B_N(_1844_),
    .Y(_1866_));
 sg13g2_nand2b_1 _3498_ (.Y(_1877_),
    .B(_1866_),
    .A_N(_1822_));
 sg13g2_or2_1 _3499_ (.X(_1888_),
    .B(net486),
    .A(_1580_));
 sg13g2_o21ai_1 _3500_ (.B1(_1855_),
    .Y(_1899_),
    .A1(_1503_),
    .A2(_1800_));
 sg13g2_nand2_1 _3501_ (.Y(_1910_),
    .A(_1877_),
    .B(_1899_));
 sg13g2_o21ai_1 _3502_ (.B1(_1877_),
    .Y(_1921_),
    .A1(_1888_),
    .A2(_1910_));
 sg13g2_inv_1 _3503_ (.Y(_1932_),
    .A(_1921_));
 sg13g2_o21ai_1 _3504_ (.B1(_1822_),
    .Y(_1943_),
    .A1(_1503_),
    .A2(net486));
 sg13g2_nor2b_1 _3505_ (.A(_1833_),
    .B_N(_1943_),
    .Y(_1954_));
 sg13g2_xnor2_1 _3506_ (.Y(_1965_),
    .A(_1921_),
    .B(_1954_));
 sg13g2_or2_1 _3507_ (.X(_1976_),
    .B(_1734_),
    .A(net486));
 sg13g2_nand2_1 _3508_ (.Y(_1987_),
    .A(_1723_),
    .B(_1976_));
 sg13g2_xnor2_1 _3509_ (.Y(_1998_),
    .A(_1822_),
    .B(_1987_));
 sg13g2_nor2_1 _3510_ (.A(_1965_),
    .B(_1998_),
    .Y(_2009_));
 sg13g2_o21ai_1 _3511_ (.B1(_1976_),
    .Y(_2020_),
    .A1(_1822_),
    .A2(_1987_));
 sg13g2_a21oi_1 _3512_ (.A1(_1921_),
    .A2(_1943_),
    .Y(_2031_),
    .B1(_1833_));
 sg13g2_mux2_1 _3513_ (.A0(_2031_),
    .A1(_1833_),
    .S(_2009_),
    .X(_2042_));
 sg13g2_nor2b_1 _3514_ (.A(_2042_),
    .B_N(_2020_),
    .Y(_2053_));
 sg13g2_a21oi_2 _3515_ (.B1(_2053_),
    .Y(_2064_),
    .A2(_2009_),
    .A1(_1833_));
 sg13g2_nand2b_1 _3516_ (.Y(_2075_),
    .B(_1580_),
    .A_N(_1503_));
 sg13g2_xnor2_1 _3517_ (.Y(_2086_),
    .A(_1811_),
    .B(_2075_));
 sg13g2_nor2b_1 _3518_ (.A(_2064_),
    .B_N(_2086_),
    .Y(_2097_));
 sg13g2_xnor2_1 _3519_ (.Y(_2108_),
    .A(_2064_),
    .B(_2086_));
 sg13g2_xor2_1 _3520_ (.B(_1910_),
    .A(_1888_),
    .X(_2119_));
 sg13g2_inv_1 _3521_ (.Y(_2130_),
    .A(_2119_));
 sg13g2_mux2_1 _3522_ (.A0(_1932_),
    .A1(_2130_),
    .S(_1591_),
    .X(_2141_));
 sg13g2_xnor2_1 _3523_ (.Y(_2152_),
    .A(_2020_),
    .B(_2042_));
 sg13g2_nand2b_1 _3524_ (.Y(_2163_),
    .B(_2152_),
    .A_N(_2141_));
 sg13g2_nor2_1 _3525_ (.A(_1580_),
    .B(_1800_),
    .Y(_2174_));
 sg13g2_or2_1 _3526_ (.X(_2185_),
    .B(_2174_),
    .A(_1866_));
 sg13g2_nor2_1 _3527_ (.A(net486),
    .B(_1800_),
    .Y(_2196_));
 sg13g2_nand2_1 _3528_ (.Y(_2207_),
    .A(_1591_),
    .B(_1844_));
 sg13g2_and2_1 _3529_ (.A(_1866_),
    .B(_2174_),
    .X(_2218_));
 sg13g2_xnor2_1 _3530_ (.Y(_2229_),
    .A(_2185_),
    .B(_2196_));
 sg13g2_a22oi_1 _3531_ (.Y(_2240_),
    .B1(_2218_),
    .B2(net486),
    .A2(_2196_),
    .A1(_2185_));
 sg13g2_xnor2_1 _3532_ (.Y(_2251_),
    .A(_1591_),
    .B(_2119_));
 sg13g2_nor2_1 _3533_ (.A(_2240_),
    .B(_2251_),
    .Y(_2262_));
 sg13g2_or2_1 _3534_ (.X(_2273_),
    .B(_2207_),
    .A(_1712_));
 sg13g2_xor2_1 _3535_ (.B(_2229_),
    .A(_2218_),
    .X(_2284_));
 sg13g2_nor2_1 _3536_ (.A(_2273_),
    .B(_2284_),
    .Y(_2295_));
 sg13g2_nand2_1 _3537_ (.Y(_2306_),
    .A(_2240_),
    .B(_2251_));
 sg13g2_nand2b_1 _3538_ (.Y(_2317_),
    .B(_2306_),
    .A_N(_2262_));
 sg13g2_a21oi_1 _3539_ (.A1(_2295_),
    .A2(_2306_),
    .Y(_2328_),
    .B1(_2262_));
 sg13g2_xor2_1 _3540_ (.B(_2152_),
    .A(_2141_),
    .X(_2339_));
 sg13g2_o21ai_1 _3541_ (.B1(_2163_),
    .Y(_2348_),
    .A1(_2328_),
    .A2(_2339_));
 sg13g2_a21oi_1 _3542_ (.A1(_2108_),
    .A2(_2348_),
    .Y(_2356_),
    .B1(_2097_));
 sg13g2_or2_1 _3543_ (.X(_2364_),
    .B(_2356_),
    .A(_1756_));
 sg13g2_a21oi_1 _3544_ (.A1(_1503_),
    .A2(_2364_),
    .Y(_2373_),
    .B1(_1261_));
 sg13g2_inv_1 _3545_ (.Y(_2381_),
    .A(_2373_));
 sg13g2_nor2_1 _3546_ (.A(net519),
    .B(_1448_),
    .Y(_2389_));
 sg13g2_nand2b_2 _3547_ (.Y(_2397_),
    .B(_1217_),
    .A_N(_1448_));
 sg13g2_nor2_1 _3548_ (.A(net514),
    .B(_1448_),
    .Y(_2405_));
 sg13g2_xnor2_1 _3549_ (.Y(_2414_),
    .A(_2328_),
    .B(_2339_));
 sg13g2_xnor2_1 _3550_ (.Y(_2425_),
    .A(_2273_),
    .B(_2284_));
 sg13g2_and2_1 _3551_ (.A(_2397_),
    .B(_2425_),
    .X(_2436_));
 sg13g2_a21oi_1 _3552_ (.A1(_2389_),
    .A2(_2414_),
    .Y(_2447_),
    .B1(_2436_));
 sg13g2_xnor2_1 _3553_ (.Y(_2458_),
    .A(_1756_),
    .B(_2356_));
 sg13g2_inv_1 _3554_ (.Y(_2469_),
    .A(_2458_));
 sg13g2_nor2_1 _3555_ (.A(_1283_),
    .B(_2458_),
    .Y(_2480_));
 sg13g2_a221oi_1 _3556_ (.B2(net520),
    .C1(_2480_),
    .B1(_2447_),
    .A1(_2373_),
    .Y(_2491_),
    .A2(_2405_));
 sg13g2_inv_1 _3557_ (.Y(_2502_),
    .A(_2491_));
 sg13g2_or2_1 _3558_ (.X(_2513_),
    .B(net602),
    .A(net599));
 sg13g2_nor2_1 _3559_ (.A(net605),
    .B(net608),
    .Y(_2524_));
 sg13g2_or2_2 _3560_ (.X(_2535_),
    .B(net607),
    .A(net605));
 sg13g2_nor4_2 _3561_ (.A(net598),
    .B(net601),
    .C(net606),
    .Y(_2546_),
    .D(net608));
 sg13g2_or4_1 _3562_ (.A(net598),
    .B(net601),
    .C(net606),
    .D(net608),
    .X(_2557_));
 sg13g2_nand2_1 _3563_ (.Y(_2568_),
    .A(_0053_),
    .B(net534));
 sg13g2_nor4_2 _3564_ (.A(net587),
    .B(_3092_),
    .C(_0064_),
    .Y(_2579_),
    .D(net533));
 sg13g2_nand4_1 _3565_ (.B(net590),
    .C(_0053_),
    .A(net537),
    .Y(_2585_),
    .D(net534));
 sg13g2_nor2_1 _3566_ (.A(net587),
    .B(net590),
    .Y(_2586_));
 sg13g2_nand2_2 _3567_ (.Y(_2587_),
    .A(net537),
    .B(_3092_));
 sg13g2_o21ai_1 _3568_ (.B1(net585),
    .Y(_2588_),
    .A1(net588),
    .A2(net591));
 sg13g2_xnor2_1 _3569_ (.Y(_2589_),
    .A(net582),
    .B(_2588_));
 sg13g2_xnor2_1 _3570_ (.Y(_2590_),
    .A(_3048_),
    .B(_2588_));
 sg13g2_nor3_2 _3571_ (.A(_0013_),
    .B(_2585_),
    .C(_2589_),
    .Y(_2591_));
 sg13g2_nand3b_1 _3572_ (.B(_2579_),
    .C(net531),
    .Y(_2592_),
    .A_N(_0013_));
 sg13g2_xnor2_1 _3573_ (.Y(_2593_),
    .A(_0013_),
    .B(_2586_));
 sg13g2_nand3b_1 _3574_ (.B(net531),
    .C(_2585_),
    .Y(_2594_),
    .A_N(_2593_));
 sg13g2_o21ai_1 _3575_ (.B1(_2593_),
    .Y(_2595_),
    .A1(_2579_),
    .A2(_2589_));
 sg13g2_nand2_2 _3576_ (.Y(_2596_),
    .A(_2594_),
    .B(_2595_));
 sg13g2_and2_1 _3577_ (.A(_2594_),
    .B(_2595_),
    .X(_2597_));
 sg13g2_nand3_1 _3578_ (.B(_0053_),
    .C(net534),
    .A(_3180_),
    .Y(_2598_));
 sg13g2_and4_1 _3579_ (.A(_0119_),
    .B(_2587_),
    .C(net530),
    .D(_2598_),
    .X(_2599_));
 sg13g2_a22oi_1 _3580_ (.Y(_2600_),
    .B1(net530),
    .B2(_2598_),
    .A2(_2587_),
    .A1(_0119_));
 sg13g2_or2_2 _3581_ (.X(_2601_),
    .B(_2600_),
    .A(_2599_));
 sg13g2_nand2b_2 _3582_ (.Y(_2602_),
    .B(net528),
    .A_N(_2601_));
 sg13g2_or2_1 _3583_ (.X(_2603_),
    .B(_2601_),
    .A(_2591_));
 sg13g2_a21oi_1 _3584_ (.A1(_2594_),
    .A2(_2595_),
    .Y(_2604_),
    .B1(_2591_));
 sg13g2_nand2_1 _3585_ (.Y(_2605_),
    .A(_2601_),
    .B(net527));
 sg13g2_a21oi_2 _3586_ (.B1(_2591_),
    .Y(_2606_),
    .A2(_2601_),
    .A1(_2596_));
 sg13g2_nand2_2 _3587_ (.Y(_2607_),
    .A(_2592_),
    .B(_2605_));
 sg13g2_nor2_1 _3588_ (.A(_2597_),
    .B(_2603_),
    .Y(_2608_));
 sg13g2_nand2_2 _3589_ (.Y(_2609_),
    .A(_2596_),
    .B(_2606_));
 sg13g2_nor3_2 _3590_ (.A(net604),
    .B(net606),
    .C(net607),
    .Y(_2610_));
 sg13g2_or3_2 _3591_ (.A(net603),
    .B(net605),
    .C(net608),
    .X(_2611_));
 sg13g2_o21ai_1 _3592_ (.B1(net603),
    .Y(_2612_),
    .A1(net605),
    .A2(net608));
 sg13g2_inv_1 _3593_ (.Y(_2613_),
    .A(_2612_));
 sg13g2_and2_2 _3594_ (.A(_2611_),
    .B(_2612_),
    .X(_2614_));
 sg13g2_nand2_2 _3595_ (.Y(_2615_),
    .A(_2611_),
    .B(_2612_));
 sg13g2_mux2_2 _3596_ (.A0(net600),
    .A1(_2615_),
    .S(net531),
    .X(_2616_));
 sg13g2_and2_2 _3597_ (.A(net605),
    .B(net608),
    .X(_2617_));
 sg13g2_nor2_1 _3598_ (.A(net535),
    .B(_2617_),
    .Y(_2618_));
 sg13g2_xnor2_1 _3599_ (.Y(_2619_),
    .A(net606),
    .B(net607));
 sg13g2_mux2_1 _3600_ (.A0(_3213_),
    .A1(_2618_),
    .S(net531),
    .X(_2620_));
 sg13g2_nor2_1 _3601_ (.A(_0016_),
    .B(net531),
    .Y(_2621_));
 sg13g2_nand2_1 _3602_ (.Y(_2622_),
    .A(net600),
    .B(net535));
 sg13g2_a21oi_1 _3603_ (.A1(net600),
    .A2(net535),
    .Y(_2623_),
    .B1(net598));
 sg13g2_a21o_1 _3604_ (.A2(net535),
    .A1(net600),
    .B1(net598),
    .X(_2624_));
 sg13g2_and3_1 _3605_ (.X(_2625_),
    .A(net598),
    .B(net600),
    .C(net535));
 sg13g2_nand3_1 _3606_ (.B(net600),
    .C(net535),
    .A(net598),
    .Y(_2626_));
 sg13g2_nand2_2 _3607_ (.Y(_2627_),
    .A(_2624_),
    .B(_2626_));
 sg13g2_a21oi_2 _3608_ (.B1(_2621_),
    .Y(_2628_),
    .A2(_2627_),
    .A1(net530));
 sg13g2_a21o_1 _3609_ (.A2(_2627_),
    .A1(net530),
    .B1(_2621_),
    .X(_2629_));
 sg13g2_a221oi_1 _3610_ (.B2(net531),
    .C1(_2621_),
    .B1(_2627_),
    .A1(_2616_),
    .Y(_2630_),
    .A2(_2620_));
 sg13g2_and3_1 _3611_ (.X(_2631_),
    .A(net590),
    .B(_2568_),
    .C(net530));
 sg13g2_a21oi_1 _3612_ (.A1(_2568_),
    .A2(net530),
    .Y(_2632_),
    .B1(net590));
 sg13g2_or2_1 _3613_ (.X(_2633_),
    .B(_2632_),
    .A(_2631_));
 sg13g2_nor4_2 _3614_ (.A(_2599_),
    .B(_2600_),
    .C(_2631_),
    .Y(_2634_),
    .D(_2632_));
 sg13g2_and2_1 _3615_ (.A(net527),
    .B(_2634_),
    .X(_2635_));
 sg13g2_nand2_2 _3616_ (.Y(_2636_),
    .A(net527),
    .B(_2634_));
 sg13g2_nand2_1 _3617_ (.Y(_2637_),
    .A(net596),
    .B(net533));
 sg13g2_nor3_1 _3618_ (.A(net596),
    .B(net598),
    .C(net601),
    .Y(_2638_));
 sg13g2_or3_2 _3619_ (.A(\hvsync_gen.hpos[4] ),
    .B(\hvsync_gen.hpos[3] ),
    .C(net602),
    .X(_2639_));
 sg13g2_nor2_1 _3620_ (.A(_2535_),
    .B(_2639_),
    .Y(_2640_));
 sg13g2_a22oi_1 _3621_ (.Y(_2641_),
    .B1(_2638_),
    .B2(net535),
    .A2(_2557_),
    .A1(net596));
 sg13g2_o21ai_1 _3622_ (.B1(_2637_),
    .Y(_2642_),
    .A1(_2535_),
    .A2(_2639_));
 sg13g2_nor2_1 _3623_ (.A(_2589_),
    .B(_2641_),
    .Y(_2643_));
 sg13g2_nand2_1 _3624_ (.Y(_2644_),
    .A(_0015_),
    .B(_2589_));
 sg13g2_nor2b_1 _3625_ (.A(_2643_),
    .B_N(_2644_),
    .Y(_2645_));
 sg13g2_nand2b_2 _3626_ (.Y(_2646_),
    .B(_2644_),
    .A_N(_2643_));
 sg13g2_nor2_1 _3627_ (.A(net592),
    .B(net530),
    .Y(_2647_));
 sg13g2_nand2_1 _3628_ (.Y(_2648_),
    .A(_0015_),
    .B(net534));
 sg13g2_o21ai_1 _3629_ (.B1(net593),
    .Y(_2649_),
    .A1(_3191_),
    .A2(net533));
 sg13g2_nand3b_1 _3630_ (.B(_0015_),
    .C(_2546_),
    .Y(_2650_),
    .A_N(net593));
 sg13g2_and2_2 _3631_ (.A(_2649_),
    .B(_2650_),
    .X(_2651_));
 sg13g2_a21oi_2 _3632_ (.B1(_2647_),
    .Y(_2652_),
    .A2(_2651_),
    .A1(net530));
 sg13g2_o21ai_1 _3633_ (.B1(_2652_),
    .Y(_2653_),
    .A1(_2630_),
    .A2(_2645_));
 sg13g2_a21o_2 _3634_ (.A2(_2653_),
    .A1(_2635_),
    .B1(_2603_),
    .X(_2654_));
 sg13g2_nand2_2 _3635_ (.Y(_2655_),
    .A(net528),
    .B(_2654_));
 sg13g2_nand4_1 _3636_ (.B(_2634_),
    .C(_2646_),
    .A(net527),
    .Y(_2656_),
    .D(_2652_));
 sg13g2_and2_1 _3637_ (.A(_2616_),
    .B(_2628_),
    .X(_2657_));
 sg13g2_nand2b_1 _3638_ (.Y(_2658_),
    .B(net527),
    .A_N(_2634_));
 sg13g2_o21ai_1 _3639_ (.B1(_2658_),
    .Y(_2659_),
    .A1(_2656_),
    .A2(_2657_));
 sg13g2_a21o_1 _3640_ (.A2(_2654_),
    .A1(net528),
    .B1(_2659_),
    .X(_2660_));
 sg13g2_and2_1 _3641_ (.A(net527),
    .B(_2656_),
    .X(_2661_));
 sg13g2_a221oi_1 _3642_ (.B2(net527),
    .C1(_2659_),
    .B1(_2656_),
    .A1(net528),
    .Y(_2662_),
    .A2(_2654_));
 sg13g2_a21oi_1 _3643_ (.A1(_2601_),
    .A2(net527),
    .Y(_2663_),
    .B1(_2662_));
 sg13g2_o21ai_1 _3644_ (.B1(_2605_),
    .Y(_2664_),
    .A1(_2660_),
    .A2(_2661_));
 sg13g2_nand3_1 _3645_ (.B(_2654_),
    .C(_2659_),
    .A(net528),
    .Y(_2665_));
 sg13g2_nand3_1 _3646_ (.B(_2661_),
    .C(_2665_),
    .A(_2660_),
    .Y(_2666_));
 sg13g2_nor2_1 _3647_ (.A(_2591_),
    .B(_2608_),
    .Y(_2667_));
 sg13g2_nand2_2 _3648_ (.Y(_2668_),
    .A(_2592_),
    .B(_2602_));
 sg13g2_nor2_1 _3649_ (.A(_2609_),
    .B(_2616_),
    .Y(_2669_));
 sg13g2_mux2_1 _3650_ (.A0(_2628_),
    .A1(_2646_),
    .S(_2655_),
    .X(_2670_));
 sg13g2_a21o_1 _3651_ (.A2(_2654_),
    .A1(net528),
    .B1(_2633_),
    .X(_2671_));
 sg13g2_nand3_1 _3652_ (.B(_2652_),
    .C(_2654_),
    .A(net528),
    .Y(_2672_));
 sg13g2_nand2_1 _3653_ (.Y(_2673_),
    .A(_2671_),
    .B(_2672_));
 sg13g2_nand4_1 _3654_ (.B(_2665_),
    .C(_2671_),
    .A(_2660_),
    .Y(_2674_),
    .D(_2672_));
 sg13g2_nand3_1 _3655_ (.B(_2666_),
    .C(_2674_),
    .A(_2663_),
    .Y(_2675_));
 sg13g2_and2_1 _3656_ (.A(_2591_),
    .B(_2675_),
    .X(_2676_));
 sg13g2_a21oi_1 _3657_ (.A1(_2664_),
    .A2(_2670_),
    .Y(_2677_),
    .B1(net522));
 sg13g2_a21o_2 _3658_ (.A2(_2677_),
    .A1(_2675_),
    .B1(_2669_),
    .X(_2678_));
 sg13g2_mux2_1 _3659_ (.A0(_2646_),
    .A1(_2652_),
    .S(_2655_),
    .X(_2679_));
 sg13g2_a21oi_1 _3660_ (.A1(_2664_),
    .A2(_2679_),
    .Y(_2680_),
    .B1(_2668_));
 sg13g2_a21oi_2 _3661_ (.B1(_2680_),
    .Y(_2681_),
    .A2(_2629_),
    .A1(net522));
 sg13g2_a21o_2 _3662_ (.A2(_2629_),
    .A1(net522),
    .B1(_2680_),
    .X(_2682_));
 sg13g2_nand2_1 _3663_ (.Y(_2683_),
    .A(_2678_),
    .B(_2682_));
 sg13g2_nand3_1 _3664_ (.B(_2633_),
    .C(_2654_),
    .A(net528),
    .Y(_2684_));
 sg13g2_nand2_1 _3665_ (.Y(_2685_),
    .A(_2597_),
    .B(_2601_));
 sg13g2_o21ai_1 _3666_ (.B1(_2685_),
    .Y(_2686_),
    .A1(_2609_),
    .A2(_2652_));
 sg13g2_nor2b_2 _3667_ (.A(_2686_),
    .B_N(_2684_),
    .Y(_2687_));
 sg13g2_inv_1 _3668_ (.Y(_2688_),
    .A(_2687_));
 sg13g2_nand2_1 _3669_ (.Y(_2689_),
    .A(_2608_),
    .B(_2620_));
 sg13g2_mux2_1 _3670_ (.A0(_2616_),
    .A1(_2628_),
    .S(_2655_),
    .X(_2690_));
 sg13g2_a21o_1 _3671_ (.A2(_2690_),
    .A1(_2664_),
    .B1(_2668_),
    .X(_2691_));
 sg13g2_nand2_2 _3672_ (.Y(_2692_),
    .A(_2689_),
    .B(_2691_));
 sg13g2_a21o_2 _3673_ (.A2(_2691_),
    .A1(_2689_),
    .B1(_2687_),
    .X(_2693_));
 sg13g2_nor2_2 _3674_ (.A(_3235_),
    .B(_2609_),
    .Y(_2694_));
 sg13g2_nand2_1 _3675_ (.Y(_2695_),
    .A(_0010_),
    .B(net522));
 sg13g2_nor2_1 _3676_ (.A(_2609_),
    .B(_2646_),
    .Y(_2696_));
 sg13g2_nand3_1 _3677_ (.B(_2660_),
    .C(_2665_),
    .A(_2602_),
    .Y(_2697_));
 sg13g2_nand3_1 _3678_ (.B(_2666_),
    .C(_2697_),
    .A(_2663_),
    .Y(_2698_));
 sg13g2_a21oi_1 _3679_ (.A1(_2664_),
    .A2(_2673_),
    .Y(_2699_),
    .B1(net522));
 sg13g2_a21o_2 _3680_ (.A2(_2699_),
    .A1(_2698_),
    .B1(_2696_),
    .X(_2700_));
 sg13g2_nor2_2 _3681_ (.A(_2687_),
    .B(_2694_),
    .Y(_2701_));
 sg13g2_inv_1 _3682_ (.Y(_2702_),
    .A(_2701_));
 sg13g2_nand2_1 _3683_ (.Y(_2703_),
    .A(_2692_),
    .B(net504));
 sg13g2_nand3_1 _3684_ (.B(net504),
    .C(_2701_),
    .A(_2692_),
    .Y(_2704_));
 sg13g2_a21oi_1 _3685_ (.A1(_2692_),
    .A2(net504),
    .Y(_2705_),
    .B1(_2701_));
 sg13g2_xnor2_1 _3686_ (.Y(_2706_),
    .A(_2701_),
    .B(_2703_));
 sg13g2_xnor2_1 _3687_ (.Y(_2707_),
    .A(_2683_),
    .B(_2706_));
 sg13g2_nand2_1 _3688_ (.Y(_2708_),
    .A(_2682_),
    .B(_2700_));
 sg13g2_nand2_2 _3689_ (.Y(_2709_),
    .A(_2678_),
    .B(net504));
 sg13g2_nand3_1 _3690_ (.B(_2682_),
    .C(_2700_),
    .A(_2678_),
    .Y(_2710_));
 sg13g2_xnor2_1 _3691_ (.Y(_2711_),
    .A(_2681_),
    .B(_2709_));
 sg13g2_xnor2_1 _3692_ (.Y(_2712_),
    .A(_2693_),
    .B(_2711_));
 sg13g2_o21ai_1 _3693_ (.B1(_2704_),
    .Y(_2713_),
    .A1(_2683_),
    .A2(_2705_));
 sg13g2_nand2_2 _3694_ (.Y(_2714_),
    .A(_2636_),
    .B(_2695_));
 sg13g2_a21oi_1 _3695_ (.A1(_2689_),
    .A2(_2691_),
    .Y(_2715_),
    .B1(_2635_));
 sg13g2_nand2_1 _3696_ (.Y(_2716_),
    .A(_2636_),
    .B(_2692_));
 sg13g2_xnor2_1 _3697_ (.Y(_2717_),
    .A(_2693_),
    .B(_2714_));
 sg13g2_or2_1 _3698_ (.X(_2718_),
    .B(_2717_),
    .A(_2709_));
 sg13g2_xor2_1 _3699_ (.B(_2717_),
    .A(_2709_),
    .X(_2719_));
 sg13g2_nand2_1 _3700_ (.Y(_2720_),
    .A(_2713_),
    .B(_2719_));
 sg13g2_xnor2_1 _3701_ (.Y(_2721_),
    .A(_2713_),
    .B(_2719_));
 sg13g2_xor2_1 _3702_ (.B(_2721_),
    .A(_2712_),
    .X(_2722_));
 sg13g2_and2_1 _3703_ (.A(_2707_),
    .B(_2722_),
    .X(_2723_));
 sg13g2_or2_1 _3704_ (.X(_2724_),
    .B(_2722_),
    .A(_2707_));
 sg13g2_xnor2_1 _3705_ (.Y(_2725_),
    .A(_2707_),
    .B(_2722_));
 sg13g2_a21oi_2 _3706_ (.B1(_2723_),
    .Y(_2726_),
    .A2(_2724_),
    .A1(_2713_));
 sg13g2_o21ai_1 _3707_ (.B1(_2710_),
    .Y(_2727_),
    .A1(_2693_),
    .A2(_2711_));
 sg13g2_o21ai_1 _3708_ (.B1(_2720_),
    .Y(_2728_),
    .A1(_2712_),
    .A2(_2721_));
 sg13g2_a21oi_1 _3709_ (.A1(_2702_),
    .A2(_2718_),
    .Y(_2729_),
    .B1(_2716_));
 sg13g2_a21oi_1 _3710_ (.A1(_2716_),
    .A2(_2718_),
    .Y(_2730_),
    .B1(_2729_));
 sg13g2_xnor2_1 _3711_ (.Y(_2731_),
    .A(_2728_),
    .B(_2730_));
 sg13g2_nor2b_1 _3712_ (.A(_2731_),
    .B_N(_2727_),
    .Y(_2732_));
 sg13g2_xor2_1 _3713_ (.B(_2731_),
    .A(_2727_),
    .X(_2733_));
 sg13g2_nor2_1 _3714_ (.A(_2726_),
    .B(_2733_),
    .Y(_2734_));
 sg13g2_xor2_1 _3715_ (.B(_2733_),
    .A(_2726_),
    .X(_2735_));
 sg13g2_a21oi_1 _3716_ (.A1(_2715_),
    .A2(_2735_),
    .Y(_2736_),
    .B1(_2734_));
 sg13g2_nand2_1 _3717_ (.Y(_2737_),
    .A(_2636_),
    .B(_2678_));
 sg13g2_inv_1 _3718_ (.Y(_2738_),
    .A(_2737_));
 sg13g2_a21oi_1 _3719_ (.A1(_2728_),
    .A2(_2730_),
    .Y(_2739_),
    .B1(_2732_));
 sg13g2_nor2_1 _3720_ (.A(_2687_),
    .B(_2715_),
    .Y(_2740_));
 sg13g2_a21oi_2 _3721_ (.B1(_2729_),
    .Y(_2741_),
    .A2(_2740_),
    .A1(_2678_));
 sg13g2_nor2b_1 _3722_ (.A(_2700_),
    .B_N(_2693_),
    .Y(_2742_));
 sg13g2_or2_1 _3723_ (.X(_2743_),
    .B(_2742_),
    .A(_2737_));
 sg13g2_inv_1 _3724_ (.Y(_2744_),
    .A(_2743_));
 sg13g2_nand2_1 _3725_ (.Y(_2745_),
    .A(_2693_),
    .B(_2738_));
 sg13g2_xor2_1 _3726_ (.B(_2745_),
    .A(net504),
    .X(_2746_));
 sg13g2_nor2_1 _3727_ (.A(_2741_),
    .B(_2746_),
    .Y(_2747_));
 sg13g2_xnor2_1 _3728_ (.Y(_2748_),
    .A(_2741_),
    .B(_2746_));
 sg13g2_nor2_1 _3729_ (.A(_2708_),
    .B(_2748_),
    .Y(_2749_));
 sg13g2_xor2_1 _3730_ (.B(_2748_),
    .A(_2708_),
    .X(_2750_));
 sg13g2_nor2b_1 _3731_ (.A(_2739_),
    .B_N(_2750_),
    .Y(_2751_));
 sg13g2_xnor2_1 _3732_ (.Y(_2752_),
    .A(_2739_),
    .B(_2750_));
 sg13g2_xnor2_1 _3733_ (.Y(_2753_),
    .A(_2738_),
    .B(_2752_));
 sg13g2_nor2_1 _3734_ (.A(_2736_),
    .B(_2753_),
    .Y(_2754_));
 sg13g2_xnor2_1 _3735_ (.Y(_2755_),
    .A(_2713_),
    .B(_2725_));
 sg13g2_a22oi_1 _3736_ (.Y(_2756_),
    .B1(_2695_),
    .B2(net504),
    .A2(_2692_),
    .A1(_2682_));
 sg13g2_nor2_2 _3737_ (.A(_2681_),
    .B(_2694_),
    .Y(_2757_));
 sg13g2_nor2b_1 _3738_ (.A(_2703_),
    .B_N(_2757_),
    .Y(_2758_));
 sg13g2_and2_1 _3739_ (.A(_2678_),
    .B(_2692_),
    .X(_2759_));
 sg13g2_nor2_1 _3740_ (.A(_2758_),
    .B(_2759_),
    .Y(_2760_));
 sg13g2_nor2_1 _3741_ (.A(_2756_),
    .B(_2760_),
    .Y(_2761_));
 sg13g2_nand2_1 _3742_ (.Y(_2762_),
    .A(_2755_),
    .B(_2761_));
 sg13g2_nor2_1 _3743_ (.A(_2755_),
    .B(_2761_),
    .Y(_2763_));
 sg13g2_xor2_1 _3744_ (.B(_2761_),
    .A(_2755_),
    .X(_2764_));
 sg13g2_o21ai_1 _3745_ (.B1(_2762_),
    .Y(_2765_),
    .A1(_2714_),
    .A2(_2763_));
 sg13g2_xnor2_1 _3746_ (.Y(_2766_),
    .A(_2716_),
    .B(_2735_));
 sg13g2_nand2_1 _3747_ (.Y(_2767_),
    .A(_2765_),
    .B(_2766_));
 sg13g2_xnor2_1 _3748_ (.Y(_2768_),
    .A(_2714_),
    .B(_2764_));
 sg13g2_nand2_1 _3749_ (.Y(_2769_),
    .A(_2678_),
    .B(_2757_));
 sg13g2_or2_1 _3750_ (.X(_2770_),
    .B(_2758_),
    .A(_2756_));
 sg13g2_xor2_1 _3751_ (.B(_2770_),
    .A(_2759_),
    .X(_2771_));
 sg13g2_or2_1 _3752_ (.X(_2772_),
    .B(_2771_),
    .A(_2769_));
 sg13g2_inv_1 _3753_ (.Y(_2773_),
    .A(_2772_));
 sg13g2_nand2_1 _3754_ (.Y(_2774_),
    .A(_2768_),
    .B(_2773_));
 sg13g2_xnor2_1 _3755_ (.Y(_2775_),
    .A(_2765_),
    .B(_2766_));
 sg13g2_o21ai_1 _3756_ (.B1(_2767_),
    .Y(_2776_),
    .A1(_2774_),
    .A2(_2775_));
 sg13g2_xor2_1 _3757_ (.B(_2753_),
    .A(_2736_),
    .X(_2777_));
 sg13g2_a21oi_1 _3758_ (.A1(_2776_),
    .A2(_2777_),
    .Y(_2778_),
    .B1(_2754_));
 sg13g2_a21oi_2 _3759_ (.B1(_2751_),
    .Y(_2779_),
    .A2(_2752_),
    .A1(_2738_));
 sg13g2_nor2_2 _3760_ (.A(_2635_),
    .B(_2681_),
    .Y(_2780_));
 sg13g2_nor2_1 _3761_ (.A(_2747_),
    .B(_2749_),
    .Y(_2781_));
 sg13g2_nor2_1 _3762_ (.A(_2681_),
    .B(_2687_),
    .Y(_2782_));
 sg13g2_nor2_1 _3763_ (.A(_2744_),
    .B(_2780_),
    .Y(_2783_));
 sg13g2_a21oi_1 _3764_ (.A1(_2682_),
    .A2(_2744_),
    .Y(_2784_),
    .B1(_2783_));
 sg13g2_xnor2_1 _3765_ (.Y(_2785_),
    .A(_2782_),
    .B(_2784_));
 sg13g2_nor2_1 _3766_ (.A(_2781_),
    .B(_2785_),
    .Y(_2786_));
 sg13g2_xor2_1 _3767_ (.B(_2785_),
    .A(_2781_),
    .X(_2787_));
 sg13g2_and2_1 _3768_ (.A(_2780_),
    .B(_2787_),
    .X(_2788_));
 sg13g2_xnor2_1 _3769_ (.Y(_2789_),
    .A(_2780_),
    .B(_2787_));
 sg13g2_or2_1 _3770_ (.X(_2790_),
    .B(_2789_),
    .A(_2779_));
 sg13g2_and2_1 _3771_ (.A(_2779_),
    .B(_2789_),
    .X(_2791_));
 sg13g2_xor2_1 _3772_ (.B(_2789_),
    .A(_2779_),
    .X(_2792_));
 sg13g2_xnor2_1 _3773_ (.Y(_2793_),
    .A(_2778_),
    .B(_2792_));
 sg13g2_nand2_1 _3774_ (.Y(_2794_),
    .A(_2606_),
    .B(_2793_));
 sg13g2_a22oi_1 _3775_ (.Y(_2795_),
    .B1(_2782_),
    .B2(_2784_),
    .A2(_2744_),
    .A1(_2682_));
 sg13g2_nand2b_1 _3776_ (.Y(_2796_),
    .B(_2688_),
    .A_N(net504));
 sg13g2_nor2_1 _3777_ (.A(_2795_),
    .B(_2796_),
    .Y(_2797_));
 sg13g2_xor2_1 _3778_ (.B(_2796_),
    .A(_2795_),
    .X(_2798_));
 sg13g2_o21ai_1 _3779_ (.B1(_2798_),
    .Y(_2799_),
    .A1(_2786_),
    .A2(_2788_));
 sg13g2_inv_1 _3780_ (.Y(_2800_),
    .A(_2799_));
 sg13g2_nor3_1 _3781_ (.A(_2786_),
    .B(_2788_),
    .C(_2798_),
    .Y(_2801_));
 sg13g2_nor2_1 _3782_ (.A(_2800_),
    .B(_2801_),
    .Y(_2802_));
 sg13g2_o21ai_1 _3783_ (.B1(_2790_),
    .Y(_2803_),
    .A1(_2778_),
    .A2(_2791_));
 sg13g2_a21oi_1 _3784_ (.A1(_2802_),
    .A2(_2803_),
    .Y(_2804_),
    .B1(_2800_));
 sg13g2_nand2_1 _3785_ (.Y(_2805_),
    .A(_2636_),
    .B(_2687_));
 sg13g2_o21ai_1 _3786_ (.B1(_2805_),
    .Y(_2806_),
    .A1(_2636_),
    .A2(_2652_));
 sg13g2_a21oi_1 _3787_ (.A1(net504),
    .A2(_2806_),
    .Y(_2807_),
    .B1(_2797_));
 sg13g2_nor2_1 _3788_ (.A(_2804_),
    .B(_2807_),
    .Y(_2808_));
 sg13g2_xnor2_1 _3789_ (.Y(_2809_),
    .A(_2804_),
    .B(_2807_));
 sg13g2_o21ai_1 _3790_ (.B1(_2794_),
    .Y(_2810_),
    .A1(_2606_),
    .A2(_2809_));
 sg13g2_xor2_1 _3791_ (.B(_2775_),
    .A(_2774_),
    .X(_2811_));
 sg13g2_nand2_1 _3792_ (.Y(_2812_),
    .A(_2606_),
    .B(_2772_));
 sg13g2_a21oi_1 _3793_ (.A1(_2769_),
    .A2(_2771_),
    .Y(_2813_),
    .B1(_2812_));
 sg13g2_a21o_1 _3794_ (.A2(_2811_),
    .A1(_2607_),
    .B1(_2813_),
    .X(_2814_));
 sg13g2_o21ai_1 _3795_ (.B1(_2636_),
    .Y(_2815_),
    .A1(_2688_),
    .A2(_2808_));
 sg13g2_nor2_1 _3796_ (.A(_2609_),
    .B(_2815_),
    .Y(_2816_));
 sg13g2_a221oi_1 _3797_ (.B2(_2591_),
    .C1(_2816_),
    .B1(_2811_),
    .A1(_2667_),
    .Y(_2817_),
    .A2(_2810_));
 sg13g2_nand3_1 _3798_ (.B(_2075_),
    .C(_2364_),
    .A(_1272_),
    .Y(_2818_));
 sg13g2_xor2_1 _3799_ (.B(_2348_),
    .A(_2108_),
    .X(_2819_));
 sg13g2_a21oi_1 _3800_ (.A1(_2397_),
    .A2(_2819_),
    .Y(_2820_),
    .B1(net514));
 sg13g2_o21ai_1 _3801_ (.B1(_2820_),
    .Y(_2821_),
    .A1(_2397_),
    .A2(_2818_));
 sg13g2_xnor2_1 _3802_ (.Y(_2822_),
    .A(_2295_),
    .B(_2317_));
 sg13g2_xor2_1 _3803_ (.B(_2207_),
    .A(_1712_),
    .X(_2823_));
 sg13g2_o21ai_1 _3804_ (.B1(_2397_),
    .Y(_2824_),
    .A1(_1800_),
    .A2(_1844_));
 sg13g2_inv_1 _3805_ (.Y(_2825_),
    .A(_2824_));
 sg13g2_a22oi_1 _3806_ (.Y(_2826_),
    .B1(_2823_),
    .B2(_2825_),
    .A2(_2822_),
    .A1(_2389_));
 sg13g2_o21ai_1 _3807_ (.B1(net514),
    .Y(_2827_),
    .A1(_1096_),
    .A2(_2826_));
 sg13g2_nand2_2 _3808_ (.Y(_2828_),
    .A(_2821_),
    .B(_2827_));
 sg13g2_nor2_1 _3809_ (.A(net471),
    .B(_2828_),
    .Y(_2829_));
 sg13g2_nand2_2 _3810_ (.Y(_2830_),
    .A(net471),
    .B(_2828_));
 sg13g2_nand2b_2 _3811_ (.Y(_2831_),
    .B(_2830_),
    .A_N(_2829_));
 sg13g2_xnor2_1 _3812_ (.Y(_2832_),
    .A(_2502_),
    .B(_2831_));
 sg13g2_xnor2_1 _3813_ (.Y(_2833_),
    .A(_2776_),
    .B(_2777_));
 sg13g2_xnor2_1 _3814_ (.Y(_2834_),
    .A(_2802_),
    .B(_2803_));
 sg13g2_mux2_1 _3815_ (.A0(_2833_),
    .A1(_2834_),
    .S(_2607_),
    .X(_2835_));
 sg13g2_nand2_1 _3816_ (.Y(_2836_),
    .A(_2636_),
    .B(_2796_));
 sg13g2_nand2_1 _3817_ (.Y(_2837_),
    .A(_2805_),
    .B(_2808_));
 sg13g2_o21ai_1 _3818_ (.B1(_2837_),
    .Y(_2838_),
    .A1(_2808_),
    .A2(_2836_));
 sg13g2_o21ai_1 _3819_ (.B1(_2609_),
    .Y(_2839_),
    .A1(_2668_),
    .A2(_2835_));
 sg13g2_o21ai_1 _3820_ (.B1(_2839_),
    .Y(_2840_),
    .A1(_2609_),
    .A2(_2838_));
 sg13g2_inv_4 _3821_ (.A(_2840_),
    .Y(_2841_));
 sg13g2_a21oi_1 _3822_ (.A1(_1448_),
    .A2(_2414_),
    .Y(_2842_),
    .B1(net514));
 sg13g2_o21ai_1 _3823_ (.B1(_2842_),
    .Y(_2843_),
    .A1(_2397_),
    .A2(_2469_));
 sg13g2_xnor2_1 _3824_ (.Y(_2844_),
    .A(_1712_),
    .B(_1800_));
 sg13g2_a22oi_1 _3825_ (.Y(_2845_),
    .B1(_2844_),
    .B2(_1448_),
    .A2(_2425_),
    .A1(_2389_));
 sg13g2_a21oi_1 _3826_ (.A1(net514),
    .A2(_2845_),
    .Y(_2846_),
    .B1(_1206_));
 sg13g2_a22oi_1 _3827_ (.Y(_2847_),
    .B1(_2843_),
    .B2(_2846_),
    .A2(_2381_),
    .A1(_1206_));
 sg13g2_nand2_1 _3828_ (.Y(_2848_),
    .A(_2841_),
    .B(_2847_));
 sg13g2_xnor2_1 _3829_ (.Y(_2849_),
    .A(net468),
    .B(_2847_));
 sg13g2_o21ai_1 _3830_ (.B1(_2848_),
    .Y(_2850_),
    .A1(_2828_),
    .A2(_2849_));
 sg13g2_and2_1 _3831_ (.A(_2832_),
    .B(_2850_),
    .X(_2851_));
 sg13g2_nand2b_1 _3832_ (.Y(_2852_),
    .B(_2604_),
    .A_N(_2793_));
 sg13g2_o21ai_1 _3833_ (.B1(_2602_),
    .Y(_2853_),
    .A1(_2607_),
    .A2(_2811_));
 sg13g2_nand2b_1 _3834_ (.Y(_2854_),
    .B(_2852_),
    .A_N(_2853_));
 sg13g2_o21ai_1 _3835_ (.B1(_2854_),
    .Y(_2855_),
    .A1(_2609_),
    .A2(_2809_));
 sg13g2_inv_4 _3836_ (.A(_2855_),
    .Y(_2856_));
 sg13g2_mux2_1 _3837_ (.A0(_2819_),
    .A1(_2822_),
    .S(_2397_),
    .X(_2857_));
 sg13g2_nor2_1 _3838_ (.A(_1096_),
    .B(_1426_),
    .Y(_2858_));
 sg13g2_a22oi_1 _3839_ (.Y(_2859_),
    .B1(_2858_),
    .B2(_2823_),
    .A2(_2857_),
    .A1(_1184_));
 sg13g2_o21ai_1 _3840_ (.B1(_2859_),
    .Y(_2860_),
    .A1(_1217_),
    .A2(_2818_));
 sg13g2_nand2_1 _3841_ (.Y(_2861_),
    .A(_2855_),
    .B(_2860_));
 sg13g2_xnor2_1 _3842_ (.Y(_2862_),
    .A(_2856_),
    .B(_2860_));
 sg13g2_nand2_1 _3843_ (.Y(_2863_),
    .A(_2847_),
    .B(_2862_));
 sg13g2_nand2_1 _3844_ (.Y(_2864_),
    .A(_2861_),
    .B(_2863_));
 sg13g2_xor2_1 _3845_ (.B(_2849_),
    .A(_2828_),
    .X(_2865_));
 sg13g2_nand2_1 _3846_ (.Y(_2866_),
    .A(_2606_),
    .B(_2834_));
 sg13g2_o21ai_1 _3847_ (.B1(_2866_),
    .Y(_2867_),
    .A1(_2606_),
    .A2(_2838_));
 sg13g2_nor3_1 _3848_ (.A(_2597_),
    .B(_2607_),
    .C(_2834_),
    .Y(_2868_));
 sg13g2_xnor2_1 _3849_ (.Y(_2869_),
    .A(_2768_),
    .B(_2773_));
 sg13g2_a21o_1 _3850_ (.A2(_2869_),
    .A1(_2597_),
    .B1(_2668_),
    .X(_2870_));
 sg13g2_a21oi_1 _3851_ (.A1(_2607_),
    .A2(_2833_),
    .Y(_2871_),
    .B1(_2870_));
 sg13g2_nor3_2 _3852_ (.A(_2676_),
    .B(_2868_),
    .C(_2871_),
    .Y(_2872_));
 sg13g2_nor3_1 _3853_ (.A(_1184_),
    .B(_2397_),
    .C(_2844_),
    .Y(_2873_));
 sg13g2_a221oi_1 _3854_ (.B2(_1206_),
    .C1(_2873_),
    .B1(_2469_),
    .A1(_1184_),
    .Y(_2874_),
    .A2(_2447_));
 sg13g2_inv_1 _3855_ (.Y(_2875_),
    .A(_2874_));
 sg13g2_nor2_1 _3856_ (.A(_2872_),
    .B(_2874_),
    .Y(_2876_));
 sg13g2_nand2_1 _3857_ (.Y(_2877_),
    .A(_2872_),
    .B(_2874_));
 sg13g2_nand2b_2 _3858_ (.Y(_2878_),
    .B(_2877_),
    .A_N(_2876_));
 sg13g2_a21oi_2 _3859_ (.B1(_2876_),
    .Y(_2879_),
    .A2(_2877_),
    .A1(_2860_));
 sg13g2_xnor2_1 _3860_ (.Y(_2880_),
    .A(_2847_),
    .B(_2862_));
 sg13g2_xor2_1 _3861_ (.B(_2878_),
    .A(_2860_),
    .X(_2881_));
 sg13g2_a221oi_1 _3862_ (.B2(_2667_),
    .C1(_2676_),
    .B1(_2814_),
    .A1(net522),
    .Y(_2882_),
    .A2(_2810_));
 sg13g2_a21oi_1 _3863_ (.A1(net519),
    .A2(_2819_),
    .Y(_2883_),
    .B1(_1426_));
 sg13g2_o21ai_1 _3864_ (.B1(_2883_),
    .Y(_2884_),
    .A1(net514),
    .A2(_2826_));
 sg13g2_inv_2 _3865_ (.Y(_2885_),
    .A(net474));
 sg13g2_nor2_1 _3866_ (.A(net473),
    .B(_2885_),
    .Y(_2886_));
 sg13g2_xnor2_1 _3867_ (.Y(_2887_),
    .A(net473),
    .B(_2884_));
 sg13g2_a21oi_1 _3868_ (.A1(_2875_),
    .A2(_2887_),
    .Y(_2888_),
    .B1(_2886_));
 sg13g2_or2_1 _3869_ (.X(_2889_),
    .B(_2888_),
    .A(_2881_));
 sg13g2_nand2_1 _3870_ (.Y(_2890_),
    .A(net522),
    .B(_2835_));
 sg13g2_xor2_1 _3871_ (.B(_2757_),
    .A(_2678_),
    .X(_2891_));
 sg13g2_a21oi_1 _3872_ (.A1(_2620_),
    .A2(_2694_),
    .Y(_2892_),
    .B1(_2607_));
 sg13g2_a21oi_1 _3873_ (.A1(_2891_),
    .A2(_2892_),
    .Y(_2893_),
    .B1(_2668_));
 sg13g2_o21ai_1 _3874_ (.B1(_2893_),
    .Y(_2894_),
    .A1(_2606_),
    .A2(_2869_));
 sg13g2_nand3_1 _3875_ (.B(_2890_),
    .C(_2894_),
    .A(_2592_),
    .Y(_2895_));
 sg13g2_xnor2_1 _3876_ (.Y(_2896_),
    .A(_2875_),
    .B(_2887_));
 sg13g2_nor3_1 _3877_ (.A(_2885_),
    .B(_2895_),
    .C(_2896_),
    .Y(_2897_));
 sg13g2_inv_1 _3878_ (.Y(_2898_),
    .A(_2897_));
 sg13g2_xnor2_1 _3879_ (.Y(_2899_),
    .A(_2881_),
    .B(_2888_));
 sg13g2_o21ai_1 _3880_ (.B1(_2889_),
    .Y(_2900_),
    .A1(_2898_),
    .A2(_2899_));
 sg13g2_xnor2_1 _3881_ (.Y(_2901_),
    .A(_2879_),
    .B(_2880_));
 sg13g2_nand2b_1 _3882_ (.Y(_2902_),
    .B(_2900_),
    .A_N(_2901_));
 sg13g2_o21ai_1 _3883_ (.B1(_2902_),
    .Y(_2903_),
    .A1(_2879_),
    .A2(_2880_));
 sg13g2_xnor2_1 _3884_ (.Y(_2904_),
    .A(_2864_),
    .B(_2865_));
 sg13g2_nor2b_1 _3885_ (.A(_2904_),
    .B_N(_2903_),
    .Y(_2905_));
 sg13g2_a21o_1 _3886_ (.A2(_2865_),
    .A1(_2864_),
    .B1(_2905_),
    .X(_2906_));
 sg13g2_xor2_1 _3887_ (.B(_2850_),
    .A(_2832_),
    .X(_2907_));
 sg13g2_a21oi_1 _3888_ (.A1(_2906_),
    .A2(_2907_),
    .Y(_2908_),
    .B1(_2851_));
 sg13g2_nor2_1 _3889_ (.A(net513),
    .B(_2818_),
    .Y(_2909_));
 sg13g2_a21oi_2 _3890_ (.B1(_2909_),
    .Y(_2910_),
    .A2(_2857_),
    .A1(net520));
 sg13g2_a21o_2 _3891_ (.A2(_2833_),
    .A1(_2591_),
    .B1(net522),
    .X(_2911_));
 sg13g2_nor2_2 _3892_ (.A(_2867_),
    .B(_2911_),
    .Y(_2912_));
 sg13g2_nor3_2 _3893_ (.A(_2491_),
    .B(_2867_),
    .C(_2911_),
    .Y(_2913_));
 sg13g2_nor2_1 _3894_ (.A(_2502_),
    .B(_2912_),
    .Y(_2914_));
 sg13g2_mux2_1 _3895_ (.A0(_2914_),
    .A1(_2913_),
    .S(_2910_),
    .X(_2915_));
 sg13g2_a21oi_1 _3896_ (.A1(_2502_),
    .A2(_2830_),
    .Y(_2916_),
    .B1(_2829_));
 sg13g2_nor2_1 _3897_ (.A(_2913_),
    .B(_2914_),
    .Y(_2917_));
 sg13g2_xor2_1 _3898_ (.B(_2917_),
    .A(_2910_),
    .X(_2918_));
 sg13g2_a22oi_1 _3899_ (.Y(_2919_),
    .B1(_2916_),
    .B2(_2918_),
    .A2(_2915_),
    .A1(_2908_));
 sg13g2_o21ai_1 _3900_ (.B1(_2915_),
    .Y(_2920_),
    .A1(_2916_),
    .A2(_2918_));
 sg13g2_nand2_1 _3901_ (.Y(_2921_),
    .A(_2908_),
    .B(_2920_));
 sg13g2_mux2_1 _3902_ (.A0(_2921_),
    .A1(_2920_),
    .S(_2919_),
    .X(_2922_));
 sg13g2_nor2_2 _3903_ (.A(\hvsync_gen.vpos[9] ),
    .B(net563),
    .Y(_2923_));
 sg13g2_nand2_2 _3904_ (.Y(_2924_),
    .A(_2971_),
    .B(_2982_));
 sg13g2_a21oi_1 _3905_ (.A1(_0228_),
    .A2(_0689_),
    .Y(_2925_),
    .B1(_0876_));
 sg13g2_o21ai_1 _3906_ (.B1(_2923_),
    .Y(_2926_),
    .A1(_0195_),
    .A2(_2925_));
 sg13g2_xnor2_1 _3907_ (.Y(_2927_),
    .A(_2906_),
    .B(_2907_));
 sg13g2_xnor2_1 _3908_ (.Y(_2928_),
    .A(_2903_),
    .B(_2904_));
 sg13g2_inv_1 _3909_ (.Y(_2929_),
    .A(_2928_));
 sg13g2_xnor2_1 _3910_ (.Y(_2930_),
    .A(_2900_),
    .B(_2901_));
 sg13g2_o21ai_1 _3911_ (.B1(_2896_),
    .Y(_2931_),
    .A1(_2885_),
    .A2(_2895_));
 sg13g2_nor2_1 _3912_ (.A(_2897_),
    .B(_2899_),
    .Y(_2932_));
 sg13g2_and2_1 _3913_ (.A(_2931_),
    .B(_2932_),
    .X(_2933_));
 sg13g2_a21oi_1 _3914_ (.A1(_2930_),
    .A2(_2933_),
    .Y(_2934_),
    .B1(_2928_));
 sg13g2_and2_1 _3915_ (.A(_2927_),
    .B(_2934_),
    .X(_2935_));
 sg13g2_nand2_1 _3916_ (.Y(_2936_),
    .A(_2926_),
    .B(_2935_));
 sg13g2_nand2_2 _3917_ (.Y(_2937_),
    .A(net567),
    .B(net570));
 sg13g2_nand3_1 _3918_ (.B(net567),
    .C(net568),
    .A(\hvsync_gen.vpos[6] ),
    .Y(_2938_));
 sg13g2_and4_2 _3919_ (.A(\hvsync_gen.vpos[7] ),
    .B(\hvsync_gen.vpos[6] ),
    .C(net567),
    .D(net568),
    .X(_2939_));
 sg13g2_nand4_1 _3920_ (.B(\hvsync_gen.vpos[6] ),
    .C(net567),
    .A(\hvsync_gen.vpos[7] ),
    .Y(_2940_),
    .D(net568));
 sg13g2_xnor2_1 _3921_ (.Y(_2941_),
    .A(net562),
    .B(_2939_));
 sg13g2_nand2_1 _3922_ (.Y(_2942_),
    .A(_3147_),
    .B(_2941_));
 sg13g2_nor4_2 _3923_ (.A(\hvsync_gen.vpos[3] ),
    .B(net573),
    .C(net576),
    .Y(_2943_),
    .D(net579));
 sg13g2_or4_2 _3924_ (.A(net572),
    .B(net573),
    .C(net578),
    .D(net579),
    .X(_2944_));
 sg13g2_nand2_1 _3925_ (.Y(_2945_),
    .A(net568),
    .B(_2943_));
 sg13g2_nor2_1 _3926_ (.A(net532),
    .B(_2944_),
    .Y(_2946_));
 sg13g2_nor2_1 _3927_ (.A(_0007_),
    .B(net532),
    .Y(_2947_));
 sg13g2_nor3_1 _3928_ (.A(_0007_),
    .B(net532),
    .C(_2944_),
    .Y(_2948_));
 sg13g2_nor4_2 _3929_ (.A(_0005_),
    .B(_0007_),
    .C(net532),
    .Y(_2949_),
    .D(_2944_));
 sg13g2_nor3_2 _3930_ (.A(net561),
    .B(_3158_),
    .C(_2939_),
    .Y(_2950_));
 sg13g2_nand3_1 _3931_ (.B(net562),
    .C(_2940_),
    .A(_3147_),
    .Y(_2951_));
 sg13g2_a21oi_2 _3932_ (.B1(_3147_),
    .Y(_2952_),
    .A2(_2940_),
    .A1(net562));
 sg13g2_o21ai_1 _3933_ (.B1(net561),
    .Y(_2953_),
    .A1(_3158_),
    .A2(_2939_));
 sg13g2_nor2_1 _3934_ (.A(_2950_),
    .B(_2952_),
    .Y(_2954_));
 sg13g2_nor3_1 _3935_ (.A(_2949_),
    .B(_2950_),
    .C(_2952_),
    .Y(_2955_));
 sg13g2_mux2_2 _3936_ (.A0(_2955_),
    .A1(net561),
    .S(_2941_),
    .X(_2956_));
 sg13g2_o21ai_1 _3937_ (.B1(_2942_),
    .Y(_2957_),
    .A1(_2941_),
    .A2(_2955_));
 sg13g2_nor3_1 _3938_ (.A(_2948_),
    .B(_2950_),
    .C(_2952_),
    .Y(_2958_));
 sg13g2_xnor2_1 _3939_ (.Y(_2959_),
    .A(_0005_),
    .B(_2947_));
 sg13g2_xnor2_1 _3940_ (.Y(_2960_),
    .A(_2958_),
    .B(_2959_));
 sg13g2_and2_1 _3941_ (.A(_2956_),
    .B(_2960_),
    .X(_2961_));
 sg13g2_nand2_2 _3942_ (.Y(_2962_),
    .A(_2956_),
    .B(_2960_));
 sg13g2_nor2b_1 _3943_ (.A(_2942_),
    .B_N(_2949_),
    .Y(_2963_));
 sg13g2_nand3_1 _3944_ (.B(_2941_),
    .C(_2949_),
    .A(_3147_),
    .Y(_2964_));
 sg13g2_nor2_1 _3945_ (.A(_3037_),
    .B(_0755_),
    .Y(_2965_));
 sg13g2_nor4_2 _3946_ (.A(_2943_),
    .B(_2950_),
    .C(_2952_),
    .Y(_2966_),
    .D(_2965_));
 sg13g2_a21oi_2 _3947_ (.B1(_0009_),
    .Y(_2967_),
    .A2(_2953_),
    .A1(_2951_));
 sg13g2_nor2_2 _3948_ (.A(_2966_),
    .B(_2967_),
    .Y(_2968_));
 sg13g2_a21oi_1 _3949_ (.A1(_2951_),
    .A2(_2953_),
    .Y(_2969_),
    .B1(_3246_));
 sg13g2_nor3_1 _3950_ (.A(_0766_),
    .B(_2950_),
    .C(_2952_),
    .Y(_2970_));
 sg13g2_nor2_1 _3951_ (.A(_2969_),
    .B(_2970_),
    .Y(_2972_));
 sg13g2_nor4_1 _3952_ (.A(_2966_),
    .B(_2967_),
    .C(_2969_),
    .D(_2970_),
    .Y(_2973_));
 sg13g2_a21oi_1 _3953_ (.A1(_2951_),
    .A2(_2953_),
    .Y(_2974_),
    .B1(net568));
 sg13g2_xnor2_1 _3954_ (.Y(_2975_),
    .A(_0003_),
    .B(_2943_));
 sg13g2_a21oi_2 _3955_ (.B1(_2974_),
    .Y(_2976_),
    .A2(_2975_),
    .A1(_2954_));
 sg13g2_a21o_1 _3956_ (.A2(_2975_),
    .A1(_2954_),
    .B1(_2974_),
    .X(_2977_));
 sg13g2_a21oi_1 _3957_ (.A1(_2951_),
    .A2(_2953_),
    .Y(_2978_),
    .B1(_0012_));
 sg13g2_nor3_1 _3958_ (.A(_0711_),
    .B(_2950_),
    .C(_2952_),
    .Y(_2979_));
 sg13g2_nor4_1 _3959_ (.A(_2966_),
    .B(_2967_),
    .C(_2978_),
    .D(_2979_),
    .Y(_2980_));
 sg13g2_nor3_1 _3960_ (.A(_2973_),
    .B(_2977_),
    .C(_2980_),
    .Y(_2981_));
 sg13g2_nand3_1 _3961_ (.B(_2951_),
    .C(_2953_),
    .A(_2945_),
    .Y(_2983_));
 sg13g2_nand2_1 _3962_ (.Y(_2984_),
    .A(_0359_),
    .B(_2937_));
 sg13g2_xnor2_1 _3963_ (.Y(_2985_),
    .A(_2983_),
    .B(_2984_));
 sg13g2_inv_1 _3964_ (.Y(_2986_),
    .A(_2985_));
 sg13g2_xnor2_1 _3965_ (.Y(_2987_),
    .A(_3169_),
    .B(net532));
 sg13g2_nor3_1 _3966_ (.A(_2946_),
    .B(_2950_),
    .C(_2952_),
    .Y(_2988_));
 sg13g2_xnor2_1 _3967_ (.Y(_2989_),
    .A(_2987_),
    .B(_2988_));
 sg13g2_inv_1 _3968_ (.Y(_2990_),
    .A(_2989_));
 sg13g2_o21ai_1 _3969_ (.B1(_2989_),
    .Y(_2991_),
    .A1(_2981_),
    .A2(_2986_));
 sg13g2_a21o_1 _3970_ (.A2(_2991_),
    .A1(_2960_),
    .B1(_2957_),
    .X(_2992_));
 sg13g2_and2_2 _3971_ (.A(_2964_),
    .B(_2992_),
    .X(_2994_));
 sg13g2_nand2_2 _3972_ (.Y(_2995_),
    .A(_2964_),
    .B(_2992_));
 sg13g2_nor2_1 _3973_ (.A(net524),
    .B(_2994_),
    .Y(_2996_));
 sg13g2_nand2_1 _3974_ (.Y(_2997_),
    .A(_2962_),
    .B(net518));
 sg13g2_nand2_1 _3975_ (.Y(_2998_),
    .A(net525),
    .B(_2989_));
 sg13g2_nor2_1 _3976_ (.A(_2960_),
    .B(net518),
    .Y(_2999_));
 sg13g2_a21oi_1 _3977_ (.A1(_2990_),
    .A2(net518),
    .Y(_3000_),
    .B1(_2999_));
 sg13g2_nand2_1 _3978_ (.Y(_3001_),
    .A(_2985_),
    .B(_2994_));
 sg13g2_nand2_1 _3979_ (.Y(_3002_),
    .A(_2976_),
    .B(_2995_));
 sg13g2_nand2_1 _3980_ (.Y(_3003_),
    .A(_2976_),
    .B(_2985_));
 sg13g2_nor3_1 _3981_ (.A(_2968_),
    .B(net521),
    .C(_3003_),
    .Y(_3005_));
 sg13g2_nand3_1 _3982_ (.B(_2976_),
    .C(_2985_),
    .A(_2973_),
    .Y(_3006_));
 sg13g2_nand3_1 _3983_ (.B(_2989_),
    .C(_3006_),
    .A(_2960_),
    .Y(_3007_));
 sg13g2_o21ai_1 _3984_ (.B1(_2956_),
    .Y(_3008_),
    .A1(_3005_),
    .A2(_3007_));
 sg13g2_nand2_1 _3985_ (.Y(_3009_),
    .A(net518),
    .B(_3008_));
 sg13g2_or2_1 _3986_ (.X(_3010_),
    .B(_3008_),
    .A(net518));
 sg13g2_nand2_1 _3987_ (.Y(_3011_),
    .A(_3009_),
    .B(_3010_));
 sg13g2_nand3_1 _3988_ (.B(_3002_),
    .C(_3011_),
    .A(_3001_),
    .Y(_3012_));
 sg13g2_o21ai_1 _3989_ (.B1(_2956_),
    .Y(_3013_),
    .A1(net521),
    .A2(_3003_));
 sg13g2_nand2_1 _3990_ (.Y(_3014_),
    .A(_3008_),
    .B(_3013_));
 sg13g2_o21ai_1 _3991_ (.B1(_3014_),
    .Y(_3016_),
    .A1(_2960_),
    .A2(_2994_));
 sg13g2_a21oi_1 _3992_ (.A1(_3009_),
    .A2(_3010_),
    .Y(_3017_),
    .B1(_3013_));
 sg13g2_a221oi_1 _3993_ (.B2(_3009_),
    .C1(_3017_),
    .B1(_3016_),
    .A1(_3000_),
    .Y(_3018_),
    .A2(_3012_));
 sg13g2_nor2_2 _3994_ (.A(net524),
    .B(_2963_),
    .Y(_3019_));
 sg13g2_and2_1 _3995_ (.A(_2968_),
    .B(_2994_),
    .X(_3020_));
 sg13g2_o21ai_1 _3996_ (.B1(_3019_),
    .Y(_3021_),
    .A1(_2972_),
    .A2(_2994_));
 sg13g2_o21ai_1 _3997_ (.B1(net525),
    .Y(_3022_),
    .A1(_2978_),
    .A2(_2979_));
 sg13g2_o21ai_1 _3998_ (.B1(_3022_),
    .Y(_3023_),
    .A1(_3020_),
    .A2(_3021_));
 sg13g2_or2_1 _3999_ (.X(_3024_),
    .B(_3023_),
    .A(_3018_));
 sg13g2_and2_1 _4000_ (.A(_2998_),
    .B(net490),
    .X(_3025_));
 sg13g2_nand2_1 _4001_ (.Y(_3027_),
    .A(_2998_),
    .B(net490));
 sg13g2_nand2_1 _4002_ (.Y(_3028_),
    .A(_2986_),
    .B(_2995_));
 sg13g2_a21oi_1 _4003_ (.A1(_2990_),
    .A2(_2994_),
    .Y(_3029_),
    .B1(net524));
 sg13g2_a22oi_1 _4004_ (.Y(_3030_),
    .B1(_3028_),
    .B2(_3029_),
    .A2(_2976_),
    .A1(net524));
 sg13g2_nand2_1 _4005_ (.Y(_3031_),
    .A(_2977_),
    .B(_3019_));
 sg13g2_nor2_1 _4006_ (.A(_2962_),
    .B(_2972_),
    .Y(_3032_));
 sg13g2_a221oi_1 _4007_ (.B2(_2957_),
    .C1(_3032_),
    .B1(_3031_),
    .A1(_2968_),
    .Y(_3033_),
    .A2(_2996_));
 sg13g2_nand2_2 _4008_ (.Y(_3034_),
    .A(_3030_),
    .B(_3033_));
 sg13g2_nand3_1 _4009_ (.B(_3002_),
    .C(_3019_),
    .A(_3001_),
    .Y(_3035_));
 sg13g2_o21ai_1 _4010_ (.B1(_3035_),
    .Y(_3036_),
    .A1(_2968_),
    .A2(_3019_));
 sg13g2_nand2_1 _4011_ (.Y(_3038_),
    .A(net503),
    .B(_3036_));
 sg13g2_nand2_2 _4012_ (.Y(_3039_),
    .A(_3033_),
    .B(_3036_));
 sg13g2_inv_1 _4013_ (.Y(_3040_),
    .A(_3039_));
 sg13g2_nor2b_2 _4014_ (.A(_3039_),
    .B_N(net503),
    .Y(_3041_));
 sg13g2_o21ai_1 _4015_ (.B1(_3000_),
    .Y(_3042_),
    .A1(_2962_),
    .A2(_2985_));
 sg13g2_inv_1 _4016_ (.Y(_3043_),
    .A(net499));
 sg13g2_and2_1 _4017_ (.A(_3024_),
    .B(_3042_),
    .X(_3044_));
 sg13g2_nand2_1 _4018_ (.Y(_3045_),
    .A(net490),
    .B(net499));
 sg13g2_xnor2_1 _4019_ (.Y(_3046_),
    .A(_3034_),
    .B(_3036_));
 sg13g2_a21oi_1 _4020_ (.A1(_3044_),
    .A2(_3046_),
    .Y(_3047_),
    .B1(_3041_));
 sg13g2_nor2_1 _4021_ (.A(_3027_),
    .B(_3047_),
    .Y(_3049_));
 sg13g2_nand2_1 _4022_ (.Y(_3050_),
    .A(_3033_),
    .B(net499));
 sg13g2_nand2_1 _4023_ (.Y(_3051_),
    .A(_3038_),
    .B(_3050_));
 sg13g2_nand2_1 _4024_ (.Y(_3052_),
    .A(net503),
    .B(net499));
 sg13g2_nor2_1 _4025_ (.A(_3039_),
    .B(_3052_),
    .Y(_3053_));
 sg13g2_nor2_1 _4026_ (.A(_3025_),
    .B(_3053_),
    .Y(_3054_));
 sg13g2_a21oi_1 _4027_ (.A1(_3051_),
    .A2(_3054_),
    .Y(_3055_),
    .B1(_3049_));
 sg13g2_nand2_1 _4028_ (.Y(_3056_),
    .A(_3036_),
    .B(net499));
 sg13g2_nand3_1 _4029_ (.B(_3036_),
    .C(net499),
    .A(net503),
    .Y(_3057_));
 sg13g2_xor2_1 _4030_ (.B(_3056_),
    .A(net503),
    .X(_3058_));
 sg13g2_nand2_2 _4031_ (.Y(_3060_),
    .A(net521),
    .B(_3033_));
 sg13g2_or2_1 _4032_ (.X(_3061_),
    .B(_3060_),
    .A(_3056_));
 sg13g2_xor2_1 _4033_ (.B(_3060_),
    .A(_3056_),
    .X(_3062_));
 sg13g2_a21oi_1 _4034_ (.A1(_3038_),
    .A2(_3050_),
    .Y(_3063_),
    .B1(_3054_));
 sg13g2_nand2_1 _4035_ (.Y(_3064_),
    .A(_3062_),
    .B(_3063_));
 sg13g2_xnor2_1 _4036_ (.Y(_3065_),
    .A(_3062_),
    .B(_3063_));
 sg13g2_xnor2_1 _4037_ (.Y(_3066_),
    .A(_3058_),
    .B(_3065_));
 sg13g2_xor2_1 _4038_ (.B(_3066_),
    .A(_3055_),
    .X(_3067_));
 sg13g2_nand2_1 _4039_ (.Y(_3068_),
    .A(_3053_),
    .B(_3067_));
 sg13g2_o21ai_1 _4040_ (.B1(_3068_),
    .Y(_3069_),
    .A1(_3055_),
    .A2(_3066_));
 sg13g2_nand2_1 _4041_ (.Y(_3071_),
    .A(net521),
    .B(_3036_));
 sg13g2_nand2b_1 _4042_ (.Y(_3072_),
    .B(_3050_),
    .A_N(_3071_));
 sg13g2_o21ai_1 _4043_ (.B1(_3064_),
    .Y(_3073_),
    .A1(_3058_),
    .A2(_3065_));
 sg13g2_nand2b_1 _4044_ (.Y(_3074_),
    .B(_3073_),
    .A_N(_3072_));
 sg13g2_xor2_1 _4045_ (.B(_3073_),
    .A(_3072_),
    .X(_3075_));
 sg13g2_xor2_1 _4046_ (.B(_3075_),
    .A(_3057_),
    .X(_3076_));
 sg13g2_nand2_1 _4047_ (.Y(_3077_),
    .A(_3069_),
    .B(_3076_));
 sg13g2_xor2_1 _4048_ (.B(_3076_),
    .A(_3069_),
    .X(_3078_));
 sg13g2_inv_1 _4049_ (.Y(_3079_),
    .A(_3078_));
 sg13g2_o21ai_1 _4050_ (.B1(_3077_),
    .Y(_3080_),
    .A1(_3071_),
    .A2(_3079_));
 sg13g2_nand2_1 _4051_ (.Y(_3082_),
    .A(net521),
    .B(net503));
 sg13g2_o21ai_1 _4052_ (.B1(_3074_),
    .Y(_3083_),
    .A1(_3057_),
    .A2(_3075_));
 sg13g2_o21ai_1 _4053_ (.B1(_3082_),
    .Y(_3084_),
    .A1(net503),
    .A2(_3043_));
 sg13g2_nand2_1 _4054_ (.Y(_3085_),
    .A(_3061_),
    .B(_3084_));
 sg13g2_nand2b_1 _4055_ (.Y(_3086_),
    .B(_3083_),
    .A_N(_3085_));
 sg13g2_xor2_1 _4056_ (.B(_3085_),
    .A(_3083_),
    .X(_3087_));
 sg13g2_xor2_1 _4057_ (.B(_3087_),
    .A(_3082_),
    .X(_3088_));
 sg13g2_nand2_1 _4058_ (.Y(_3089_),
    .A(_3080_),
    .B(_3088_));
 sg13g2_xnor2_1 _4059_ (.Y(_3090_),
    .A(_3045_),
    .B(_3046_));
 sg13g2_and2_1 _4060_ (.A(_3040_),
    .B(_3090_),
    .X(_3091_));
 sg13g2_and2_1 _4061_ (.A(_0006_),
    .B(net525),
    .X(_3093_));
 sg13g2_nand2_2 _4062_ (.Y(_3094_),
    .A(_0006_),
    .B(net525));
 sg13g2_nand2_1 _4063_ (.Y(_3095_),
    .A(net503),
    .B(_3094_));
 sg13g2_inv_1 _4064_ (.Y(_3096_),
    .A(_3095_));
 sg13g2_nand2_1 _4065_ (.Y(_3097_),
    .A(net521),
    .B(_3094_));
 sg13g2_inv_1 _4066_ (.Y(_3098_),
    .A(_3097_));
 sg13g2_nor2_1 _4067_ (.A(_3034_),
    .B(_3097_),
    .Y(_3099_));
 sg13g2_xnor2_1 _4068_ (.Y(_3100_),
    .A(_3034_),
    .B(_3098_));
 sg13g2_xnor2_1 _4069_ (.Y(_3101_),
    .A(_3045_),
    .B(_3100_));
 sg13g2_xnor2_1 _4070_ (.Y(_3102_),
    .A(_3039_),
    .B(_3090_));
 sg13g2_a21oi_1 _4071_ (.A1(_3101_),
    .A2(_3102_),
    .Y(_3104_),
    .B1(_3091_));
 sg13g2_xnor2_1 _4072_ (.Y(_3105_),
    .A(_3027_),
    .B(_3047_));
 sg13g2_nor2_1 _4073_ (.A(_3104_),
    .B(_3105_),
    .Y(_3106_));
 sg13g2_a21oi_2 _4074_ (.B1(_3099_),
    .Y(_3107_),
    .A2(_3100_),
    .A1(_3044_));
 sg13g2_inv_1 _4075_ (.Y(_3108_),
    .A(_3107_));
 sg13g2_xor2_1 _4076_ (.B(_3105_),
    .A(_3104_),
    .X(_3109_));
 sg13g2_a21oi_2 _4077_ (.B1(_3106_),
    .Y(_3110_),
    .A2(_3109_),
    .A1(_3108_));
 sg13g2_xnor2_1 _4078_ (.Y(_3111_),
    .A(_3053_),
    .B(_3067_));
 sg13g2_nor2_1 _4079_ (.A(_3110_),
    .B(_3111_),
    .Y(_3112_));
 sg13g2_xor2_1 _4080_ (.B(_3111_),
    .A(_3110_),
    .X(_3113_));
 sg13g2_nor2b_1 _4081_ (.A(_3060_),
    .B_N(_3113_),
    .Y(_3115_));
 sg13g2_nor2_1 _4082_ (.A(_3112_),
    .B(_3115_),
    .Y(_3116_));
 sg13g2_xor2_1 _4083_ (.B(_3078_),
    .A(_3071_),
    .X(_3117_));
 sg13g2_nor2_1 _4084_ (.A(_3116_),
    .B(_3117_),
    .Y(_3118_));
 sg13g2_and2_1 _4085_ (.A(net490),
    .B(_3030_),
    .X(_3119_));
 sg13g2_xor2_1 _4086_ (.B(_3102_),
    .A(_3101_),
    .X(_3120_));
 sg13g2_nand2_1 _4087_ (.Y(_3121_),
    .A(_3119_),
    .B(_3120_));
 sg13g2_nand2_1 _4088_ (.Y(_3122_),
    .A(net499),
    .B(_3094_));
 sg13g2_xnor2_1 _4089_ (.Y(_3123_),
    .A(_3119_),
    .B(_3120_));
 sg13g2_o21ai_1 _4090_ (.B1(_3121_),
    .Y(_3124_),
    .A1(_3122_),
    .A2(_3123_));
 sg13g2_xnor2_1 _4091_ (.Y(_3126_),
    .A(_3107_),
    .B(_3109_));
 sg13g2_and2_1 _4092_ (.A(_3124_),
    .B(_3126_),
    .X(_3127_));
 sg13g2_xor2_1 _4093_ (.B(_3126_),
    .A(_3124_),
    .X(_3128_));
 sg13g2_a21oi_1 _4094_ (.A1(_3025_),
    .A2(_3128_),
    .Y(_3129_),
    .B1(_3127_));
 sg13g2_xnor2_1 _4095_ (.Y(_3130_),
    .A(_3060_),
    .B(_3113_));
 sg13g2_nand2b_1 _4096_ (.Y(_3131_),
    .B(_3130_),
    .A_N(_3129_));
 sg13g2_xor2_1 _4097_ (.B(_3036_),
    .A(_3033_),
    .X(_3132_));
 sg13g2_and2_1 _4098_ (.A(net490),
    .B(_3132_),
    .X(_3133_));
 sg13g2_a22oi_1 _4099_ (.Y(_3134_),
    .B1(_3096_),
    .B2(_3133_),
    .A2(_3040_),
    .A1(net490));
 sg13g2_xnor2_1 _4100_ (.Y(_3135_),
    .A(_3122_),
    .B(_3123_));
 sg13g2_nor2_1 _4101_ (.A(_3134_),
    .B(_3135_),
    .Y(_3137_));
 sg13g2_xor2_1 _4102_ (.B(_3135_),
    .A(_3134_),
    .X(_3138_));
 sg13g2_a21oi_2 _4103_ (.B1(_3137_),
    .Y(_3139_),
    .A2(_3138_),
    .A1(_3098_));
 sg13g2_xnor2_1 _4104_ (.Y(_3140_),
    .A(_3025_),
    .B(_3128_));
 sg13g2_nor2_1 _4105_ (.A(_3139_),
    .B(_3140_),
    .Y(_3141_));
 sg13g2_xnor2_1 _4106_ (.Y(_3142_),
    .A(_3096_),
    .B(_3133_));
 sg13g2_nor3_2 _4107_ (.A(_3039_),
    .B(_3093_),
    .C(_3095_),
    .Y(_3143_));
 sg13g2_xnor2_1 _4108_ (.Y(_3144_),
    .A(_3097_),
    .B(_3138_));
 sg13g2_and2_1 _4109_ (.A(_3143_),
    .B(_3144_),
    .X(_3145_));
 sg13g2_xor2_1 _4110_ (.B(_3140_),
    .A(_3139_),
    .X(_3146_));
 sg13g2_a21oi_1 _4111_ (.A1(_3145_),
    .A2(_3146_),
    .Y(_3148_),
    .B1(_3141_));
 sg13g2_xnor2_1 _4112_ (.Y(_3149_),
    .A(_3129_),
    .B(_3130_));
 sg13g2_nand2b_1 _4113_ (.Y(_3150_),
    .B(_3149_),
    .A_N(_3148_));
 sg13g2_nand2_1 _4114_ (.Y(_3151_),
    .A(_3131_),
    .B(_3150_));
 sg13g2_xor2_1 _4115_ (.B(_3117_),
    .A(_3116_),
    .X(_3152_));
 sg13g2_a21oi_2 _4116_ (.B1(_3118_),
    .Y(_3153_),
    .A2(_3152_),
    .A1(_3151_));
 sg13g2_xnor2_1 _4117_ (.Y(_3154_),
    .A(_3080_),
    .B(_3088_));
 sg13g2_o21ai_1 _4118_ (.B1(_3089_),
    .Y(_3155_),
    .A1(_3153_),
    .A2(_3154_));
 sg13g2_o21ai_1 _4119_ (.B1(_3086_),
    .Y(_3156_),
    .A1(_3082_),
    .A2(_3087_));
 sg13g2_nand2_1 _4120_ (.Y(_3157_),
    .A(_3052_),
    .B(_3061_));
 sg13g2_o21ai_1 _4121_ (.B1(_3157_),
    .Y(_3159_),
    .A1(_3057_),
    .A2(_3060_));
 sg13g2_nand2b_1 _4122_ (.Y(_3160_),
    .B(_3156_),
    .A_N(_3159_));
 sg13g2_xor2_1 _4123_ (.B(_3159_),
    .A(_3156_),
    .X(_3161_));
 sg13g2_nand2b_1 _4124_ (.Y(_3162_),
    .B(_3155_),
    .A_N(_3161_));
 sg13g2_xor2_1 _4125_ (.B(_3161_),
    .A(_3155_),
    .X(_3163_));
 sg13g2_nor2_1 _4126_ (.A(_2997_),
    .B(_3163_),
    .Y(_3164_));
 sg13g2_xnor2_1 _4127_ (.Y(_3165_),
    .A(_3151_),
    .B(_3152_));
 sg13g2_nor2_1 _4128_ (.A(net518),
    .B(_3165_),
    .Y(_3166_));
 sg13g2_nor2_1 _4129_ (.A(_3164_),
    .B(_3166_),
    .Y(_3167_));
 sg13g2_nand2_1 _4130_ (.Y(_3168_),
    .A(_3160_),
    .B(_3162_));
 sg13g2_o21ai_1 _4131_ (.B1(net521),
    .Y(_3170_),
    .A1(_3041_),
    .A2(_3043_));
 sg13g2_nand2b_1 _4132_ (.Y(_3171_),
    .B(_3168_),
    .A_N(_3170_));
 sg13g2_o21ai_1 _4133_ (.B1(net521),
    .Y(_3172_),
    .A1(_2962_),
    .A2(net499));
 sg13g2_a22oi_1 _4134_ (.Y(_3173_),
    .B1(_3171_),
    .B2(_3172_),
    .A2(_3167_),
    .A1(_3019_));
 sg13g2_nand2_1 _4135_ (.Y(_3174_),
    .A(_2912_),
    .B(_3173_));
 sg13g2_xor2_1 _4136_ (.B(_3154_),
    .A(_3153_),
    .X(_3175_));
 sg13g2_nor2_1 _4137_ (.A(_2994_),
    .B(_3175_),
    .Y(_3176_));
 sg13g2_xnor2_1 _4138_ (.Y(_3177_),
    .A(_3148_),
    .B(_3149_));
 sg13g2_o21ai_1 _4139_ (.B1(_2962_),
    .Y(_3178_),
    .A1(net518),
    .A2(_3177_));
 sg13g2_nor2_1 _4140_ (.A(_3176_),
    .B(_3178_),
    .Y(_3179_));
 sg13g2_xnor2_1 _4141_ (.Y(_3181_),
    .A(_3168_),
    .B(_3170_));
 sg13g2_a21oi_1 _4142_ (.A1(net524),
    .A2(_3181_),
    .Y(_3182_),
    .B1(_3179_));
 sg13g2_nor2_1 _4143_ (.A(net470),
    .B(_3182_),
    .Y(_3183_));
 sg13g2_xor2_1 _4144_ (.B(_3146_),
    .A(_3145_),
    .X(_3184_));
 sg13g2_o21ai_1 _4145_ (.B1(_2964_),
    .Y(_3185_),
    .A1(_2956_),
    .A2(_3184_));
 sg13g2_a221oi_1 _4146_ (.B2(_2996_),
    .C1(_3185_),
    .B1(_3165_),
    .A1(net524),
    .Y(_3186_),
    .A2(_3163_));
 sg13g2_nand2_1 _4147_ (.Y(_3187_),
    .A(net468),
    .B(_3186_));
 sg13g2_nor2_1 _4148_ (.A(_2962_),
    .B(_3175_),
    .Y(_3188_));
 sg13g2_xnor2_1 _4149_ (.Y(_3189_),
    .A(_3143_),
    .B(_3144_));
 sg13g2_a21oi_1 _4150_ (.A1(_2957_),
    .A2(_3189_),
    .Y(_3190_),
    .B1(_2963_));
 sg13g2_o21ai_1 _4151_ (.B1(_3190_),
    .Y(_3192_),
    .A1(_2997_),
    .A2(_3177_));
 sg13g2_nor2_1 _4152_ (.A(_3188_),
    .B(_3192_),
    .Y(_3193_));
 sg13g2_nor3_1 _4153_ (.A(_2856_),
    .B(_3188_),
    .C(_3192_),
    .Y(_3194_));
 sg13g2_o21ai_1 _4154_ (.B1(_3142_),
    .Y(_3195_),
    .A1(_3039_),
    .A2(_3093_));
 sg13g2_nor2_1 _4155_ (.A(_2995_),
    .B(_3143_),
    .Y(_3196_));
 sg13g2_a22oi_1 _4156_ (.Y(_3197_),
    .B1(_3195_),
    .B2(_3196_),
    .A2(_3184_),
    .A1(_2996_));
 sg13g2_nand2b_1 _4157_ (.Y(_3198_),
    .B(_3033_),
    .A_N(net490));
 sg13g2_xor2_1 _4158_ (.B(_3033_),
    .A(net490),
    .X(_3199_));
 sg13g2_a21oi_1 _4159_ (.A1(_3094_),
    .A2(_3199_),
    .Y(_3200_),
    .B1(_2964_));
 sg13g2_a221oi_1 _4160_ (.B2(_3019_),
    .C1(_3200_),
    .B1(_3197_),
    .A1(net524),
    .Y(_3201_),
    .A2(_3165_));
 sg13g2_nand2b_1 _4161_ (.Y(_3203_),
    .B(_3201_),
    .A_N(net475));
 sg13g2_o21ai_1 _4162_ (.B1(_2994_),
    .Y(_3204_),
    .A1(_3093_),
    .A2(_3132_));
 sg13g2_a21o_1 _4163_ (.A2(_3198_),
    .A1(_3093_),
    .B1(_3204_),
    .X(_3205_));
 sg13g2_o21ai_1 _4164_ (.B1(_3205_),
    .Y(_3206_),
    .A1(_2997_),
    .A2(_3189_));
 sg13g2_a22oi_1 _4165_ (.Y(_3207_),
    .B1(_3206_),
    .B2(_3019_),
    .A2(_3177_),
    .A1(net524));
 sg13g2_or2_1 _4166_ (.X(_3208_),
    .B(_3207_),
    .A(net472));
 sg13g2_xor2_1 _4167_ (.B(_3201_),
    .A(net475),
    .X(_3209_));
 sg13g2_o21ai_1 _4168_ (.B1(_3203_),
    .Y(_3210_),
    .A1(_3208_),
    .A2(_3209_));
 sg13g2_xnor2_1 _4169_ (.Y(_3211_),
    .A(_2856_),
    .B(_3193_));
 sg13g2_a21o_1 _4170_ (.A2(_3211_),
    .A1(_3210_),
    .B1(_3194_),
    .X(_3212_));
 sg13g2_xnor2_1 _4171_ (.Y(_3214_),
    .A(_2840_),
    .B(_3186_));
 sg13g2_nand2_1 _4172_ (.Y(_3215_),
    .A(_3212_),
    .B(_3214_));
 sg13g2_xnor2_1 _4173_ (.Y(_3216_),
    .A(net470),
    .B(_3182_));
 sg13g2_a21oi_1 _4174_ (.A1(_3187_),
    .A2(_3215_),
    .Y(_3217_),
    .B1(_3216_));
 sg13g2_nor2_1 _4175_ (.A(_3183_),
    .B(_3217_),
    .Y(_3218_));
 sg13g2_xnor2_1 _4176_ (.Y(_3219_),
    .A(_2912_),
    .B(_3173_));
 sg13g2_o21ai_1 _4177_ (.B1(_3174_),
    .Y(_3220_),
    .A1(_3218_),
    .A2(_3219_));
 sg13g2_mux2_1 _4178_ (.A0(_3175_),
    .A1(_3181_),
    .S(net518),
    .X(_3221_));
 sg13g2_a21oi_1 _4179_ (.A1(_3019_),
    .A2(_3221_),
    .Y(_3222_),
    .B1(_3018_));
 sg13g2_xnor2_1 _4180_ (.Y(_3223_),
    .A(_3218_),
    .B(_3219_));
 sg13g2_nand3_1 _4181_ (.B(_3215_),
    .C(_3216_),
    .A(_3187_),
    .Y(_3225_));
 sg13g2_nor2b_1 _4182_ (.A(_3217_),
    .B_N(_3225_),
    .Y(_3226_));
 sg13g2_xnor2_1 _4183_ (.Y(_3227_),
    .A(_3210_),
    .B(_3211_));
 sg13g2_xnor2_1 _4184_ (.Y(_3228_),
    .A(_3212_),
    .B(_3214_));
 sg13g2_a21oi_1 _4185_ (.A1(_3227_),
    .A2(_3228_),
    .Y(_3229_),
    .B1(_3223_));
 sg13g2_xnor2_1 _4186_ (.Y(_3230_),
    .A(_3220_),
    .B(_3222_));
 sg13g2_a21o_2 _4187_ (.A2(_3229_),
    .A1(_3226_),
    .B1(_3230_),
    .X(_3231_));
 sg13g2_nand2b_1 _4188_ (.Y(_3232_),
    .B(_2965_),
    .A_N(_2938_));
 sg13g2_nand3_1 _4189_ (.B(_2993_),
    .C(_3232_),
    .A(_2982_),
    .Y(_3233_));
 sg13g2_o21ai_1 _4190_ (.B1(net599),
    .Y(_3234_),
    .A1(net601),
    .A2(net606));
 sg13g2_nand2_1 _4191_ (.Y(_3236_),
    .A(_3103_),
    .B(_3234_));
 sg13g2_nand2_1 _4192_ (.Y(_3237_),
    .A(net585),
    .B(_0108_));
 sg13g2_nand4_1 _4193_ (.B(net595),
    .C(_0108_),
    .A(net585),
    .Y(_3238_),
    .D(_3236_));
 sg13g2_nor2_1 _4194_ (.A(net568),
    .B(net572),
    .Y(_3239_));
 sg13g2_o21ai_1 _4195_ (.B1(_2993_),
    .Y(_3240_),
    .A1(_0173_),
    .A2(_3239_));
 sg13g2_nand2_1 _4196_ (.Y(_3241_),
    .A(net563),
    .B(_3240_));
 sg13g2_nor2_1 _4197_ (.A(\hvsync_gen.vpos[9] ),
    .B(net583),
    .Y(_3242_));
 sg13g2_nand4_1 _4198_ (.B(_3238_),
    .C(_3241_),
    .A(_3233_),
    .Y(_3243_),
    .D(_3242_));
 sg13g2_a21oi_1 _4199_ (.A1(net601),
    .A2(_2617_),
    .Y(_3244_),
    .B1(net599));
 sg13g2_nor3_1 _4200_ (.A(net537),
    .B(net591),
    .C(net595),
    .Y(_3245_));
 sg13g2_o21ai_1 _4201_ (.B1(_3245_),
    .Y(_3247_),
    .A1(_3103_),
    .A2(_3244_));
 sg13g2_a21oi_1 _4202_ (.A1(_3224_),
    .A2(_3247_),
    .Y(_3248_),
    .B1(net585));
 sg13g2_nor2_1 _4203_ (.A(net583),
    .B(net585),
    .Y(_3249_));
 sg13g2_or3_2 _4204_ (.A(_3231_),
    .B(_3243_),
    .C(_3248_),
    .X(_3250_));
 sg13g2_o21ai_1 _4205_ (.B1(_0015_),
    .Y(_3251_),
    .A1(net597),
    .A2(_3234_));
 sg13g2_and2_1 _4206_ (.A(net591),
    .B(\hvsync_gen.hpos[5] ),
    .X(_3252_));
 sg13g2_a21oi_1 _4207_ (.A1(_3251_),
    .A2(_3252_),
    .Y(_3253_),
    .B1(_3224_));
 sg13g2_xor2_1 _4208_ (.B(_3253_),
    .A(_0013_),
    .X(_3254_));
 sg13g2_nand2_2 _4209_ (.Y(_3255_),
    .A(net578),
    .B(net579));
 sg13g2_a21oi_2 _4210_ (.B1(net573),
    .Y(_3256_),
    .A2(net580),
    .A1(net576));
 sg13g2_a21o_1 _4211_ (.A2(net580),
    .A1(net576),
    .B1(net573),
    .X(_3258_));
 sg13g2_nor2_1 _4212_ (.A(net571),
    .B(_3258_),
    .Y(_3259_));
 sg13g2_a21o_2 _4213_ (.A2(_3256_),
    .A1(_3239_),
    .B1(_3015_),
    .X(_3260_));
 sg13g2_and2_1 _4214_ (.A(_3004_),
    .B(_3260_),
    .X(_3261_));
 sg13g2_nand3_1 _4215_ (.B(_0249_),
    .C(_3260_),
    .A(net562),
    .Y(_3262_));
 sg13g2_a21oi_1 _4216_ (.A1(_0249_),
    .A2(_3260_),
    .Y(_3263_),
    .B1(net562));
 sg13g2_nor2_1 _4217_ (.A(net540),
    .B(_3263_),
    .Y(_3264_));
 sg13g2_a22oi_1 _4218_ (.Y(_3265_),
    .B1(_3262_),
    .B2(_3264_),
    .A2(_3254_),
    .A1(net540));
 sg13g2_a21o_1 _4219_ (.A2(_3252_),
    .A1(_3251_),
    .B1(net587),
    .X(_3266_));
 sg13g2_a21oi_1 _4220_ (.A1(net584),
    .A2(_3266_),
    .Y(_3267_),
    .B1(_3125_));
 sg13g2_a21o_1 _4221_ (.A2(_3266_),
    .A1(net584),
    .B1(_3125_),
    .X(_3269_));
 sg13g2_and3_1 _4222_ (.X(_3270_),
    .A(net584),
    .B(_3125_),
    .C(_3266_));
 sg13g2_nor2_2 _4223_ (.A(net549),
    .B(_3270_),
    .Y(_3271_));
 sg13g2_nor3_2 _4224_ (.A(net550),
    .B(_3267_),
    .C(_3270_),
    .Y(_3272_));
 sg13g2_a21oi_1 _4225_ (.A1(_0249_),
    .A2(_3260_),
    .Y(_3273_),
    .B1(_2982_));
 sg13g2_o21ai_1 _4226_ (.B1(net554),
    .Y(_3274_),
    .A1(\hvsync_gen.vpos[9] ),
    .A2(_3273_));
 sg13g2_a21oi_1 _4227_ (.A1(\hvsync_gen.vpos[9] ),
    .A2(_3273_),
    .Y(_3275_),
    .B1(_3274_));
 sg13g2_nor2_1 _4228_ (.A(_3272_),
    .B(net523),
    .Y(_3276_));
 sg13g2_xnor2_1 _4229_ (.Y(_3277_),
    .A(_0005_),
    .B(_3261_));
 sg13g2_nand3_1 _4230_ (.B(_0108_),
    .C(_3251_),
    .A(net594),
    .Y(_3278_));
 sg13g2_nand3_1 _4231_ (.B(_3266_),
    .C(_3278_),
    .A(net540),
    .Y(_0043_));
 sg13g2_o21ai_1 _4232_ (.B1(_0043_),
    .Y(_0044_),
    .A1(net540),
    .A2(_3277_));
 sg13g2_o21ai_1 _4233_ (.B1(_3234_),
    .Y(_0045_),
    .A1(net606),
    .A2(_2513_));
 sg13g2_nand2_1 _4234_ (.Y(_0046_),
    .A(net541),
    .B(_0045_));
 sg13g2_nand3_1 _4235_ (.B(_0011_),
    .C(_3255_),
    .A(_0009_),
    .Y(_0047_));
 sg13g2_a21o_1 _4236_ (.A2(_3255_),
    .A1(_0011_),
    .B1(_0009_),
    .X(_0048_));
 sg13g2_nand3_1 _4237_ (.B(_0047_),
    .C(_0048_),
    .A(net550),
    .Y(_0049_));
 sg13g2_nand2_2 _4238_ (.Y(_0050_),
    .A(_0046_),
    .B(_0049_));
 sg13g2_nor2b_2 _4239_ (.A(net552),
    .B_N(net605),
    .Y(_0051_));
 sg13g2_a21o_2 _4240_ (.A2(_0711_),
    .A1(net554),
    .B1(_0051_),
    .X(_0052_));
 sg13g2_o21ai_1 _4241_ (.B1(_0656_),
    .Y(_0054_),
    .A1(net549),
    .A2(_3235_));
 sg13g2_xnor2_1 _4242_ (.Y(_0055_),
    .A(net604),
    .B(net606));
 sg13g2_and3_2 _4243_ (.X(_0056_),
    .A(net573),
    .B(net578),
    .C(net579));
 sg13g2_nor2_1 _4244_ (.A(_3256_),
    .B(_0056_),
    .Y(_0057_));
 sg13g2_o21ai_1 _4245_ (.B1(net554),
    .Y(_0058_),
    .A1(_3256_),
    .A2(_0056_));
 sg13g2_nand2_1 _4246_ (.Y(_0059_),
    .A(net541),
    .B(_0055_));
 sg13g2_nand2_1 _4247_ (.Y(_0060_),
    .A(_0058_),
    .B(_0059_));
 sg13g2_and4_1 _4248_ (.A(_0052_),
    .B(_0054_),
    .C(_0058_),
    .D(_0059_),
    .X(_0061_));
 sg13g2_nand4_1 _4249_ (.B(_0054_),
    .C(_0058_),
    .A(_0052_),
    .Y(_0062_),
    .D(_0059_));
 sg13g2_xnor2_1 _4250_ (.Y(_0063_),
    .A(net596),
    .B(_3234_));
 sg13g2_nand2_1 _4251_ (.Y(_0065_),
    .A(net540),
    .B(_0063_));
 sg13g2_nand3_1 _4252_ (.B(_0003_),
    .C(_3256_),
    .A(_3037_),
    .Y(_0066_));
 sg13g2_o21ai_1 _4253_ (.B1(_3136_),
    .Y(_0067_),
    .A1(net572),
    .A2(_3258_));
 sg13g2_nand3_1 _4254_ (.B(_0066_),
    .C(_0067_),
    .A(net554),
    .Y(_0068_));
 sg13g2_nand2_2 _4255_ (.Y(_0069_),
    .A(_0065_),
    .B(_0068_));
 sg13g2_a221oi_1 _4256_ (.B2(_0068_),
    .C1(_0062_),
    .B1(_0065_),
    .A1(_0046_),
    .Y(_0070_),
    .A2(_0049_));
 sg13g2_a21oi_2 _4257_ (.B1(net544),
    .Y(_0071_),
    .A2(_3259_),
    .A1(_0348_));
 sg13g2_xor2_1 _4258_ (.B(_3251_),
    .A(net594),
    .X(_0072_));
 sg13g2_a22oi_1 _4259_ (.Y(_0073_),
    .B1(_0072_),
    .B2(net540),
    .A2(_0071_),
    .A1(_3260_));
 sg13g2_o21ai_1 _4260_ (.B1(net550),
    .Y(_0074_),
    .A1(_3169_),
    .A2(_3260_));
 sg13g2_a21o_1 _4261_ (.A2(_3260_),
    .A1(_3169_),
    .B1(_0074_),
    .X(_0076_));
 sg13g2_a21o_1 _4262_ (.A2(_3251_),
    .A1(net594),
    .B1(_3180_),
    .X(_0077_));
 sg13g2_nand3_1 _4263_ (.B(_3180_),
    .C(_3251_),
    .A(net594),
    .Y(_0078_));
 sg13g2_nand3_1 _4264_ (.B(_0077_),
    .C(_0078_),
    .A(net540),
    .Y(_0079_));
 sg13g2_nand2_1 _4265_ (.Y(_0080_),
    .A(_0076_),
    .B(_0079_));
 sg13g2_and4_1 _4266_ (.A(_0070_),
    .B(_0073_),
    .C(_0076_),
    .D(_0079_),
    .X(_0081_));
 sg13g2_a221oi_1 _4267_ (.B2(_0081_),
    .C1(net523),
    .B1(_0044_),
    .A1(_3269_),
    .Y(_0082_),
    .A2(_3271_));
 sg13g2_xor2_1 _4268_ (.B(_0082_),
    .A(_3265_),
    .X(_0083_));
 sg13g2_xnor2_1 _4269_ (.Y(_0084_),
    .A(_3265_),
    .B(_0082_));
 sg13g2_nand4_1 _4270_ (.B(_3276_),
    .C(_0044_),
    .A(_3265_),
    .Y(_0085_),
    .D(_0081_));
 sg13g2_and2_1 _4271_ (.A(_0083_),
    .B(_0085_),
    .X(_0087_));
 sg13g2_nand2_1 _4272_ (.Y(_0088_),
    .A(_0083_),
    .B(_0085_));
 sg13g2_a221oi_1 _4273_ (.B2(_0073_),
    .C1(_3275_),
    .B1(_0070_),
    .A1(_3269_),
    .Y(_0089_),
    .A2(_3271_));
 sg13g2_xnor2_1 _4274_ (.Y(_0090_),
    .A(_0080_),
    .B(_0089_));
 sg13g2_nor3_1 _4275_ (.A(_3272_),
    .B(net523),
    .C(_0081_),
    .Y(_0091_));
 sg13g2_xor2_1 _4276_ (.B(_0091_),
    .A(_0044_),
    .X(_0092_));
 sg13g2_a21o_1 _4277_ (.A2(_0092_),
    .A1(_0090_),
    .B1(_0088_),
    .X(_0093_));
 sg13g2_inv_2 _4278_ (.Y(_0094_),
    .A(net511));
 sg13g2_and2_1 _4279_ (.A(_0087_),
    .B(net512),
    .X(_0095_));
 sg13g2_nand3_1 _4280_ (.B(_0090_),
    .C(_0092_),
    .A(_0087_),
    .Y(_0096_));
 sg13g2_nor3_2 _4281_ (.A(_3272_),
    .B(net523),
    .C(_0061_),
    .Y(_0098_));
 sg13g2_xnor2_1 _4282_ (.Y(_0099_),
    .A(_0050_),
    .B(_0098_));
 sg13g2_xor2_1 _4283_ (.B(_0098_),
    .A(_0050_),
    .X(_0100_));
 sg13g2_nor3_1 _4284_ (.A(_3272_),
    .B(net523),
    .C(_0054_),
    .Y(_0101_));
 sg13g2_xnor2_1 _4285_ (.Y(_0102_),
    .A(_0052_),
    .B(_0101_));
 sg13g2_a221oi_1 _4286_ (.B2(_0054_),
    .C1(net523),
    .B1(_0052_),
    .A1(_3269_),
    .Y(_0103_),
    .A2(_3271_));
 sg13g2_xnor2_1 _4287_ (.Y(_0104_),
    .A(_0060_),
    .B(_0103_));
 sg13g2_a21oi_1 _4288_ (.A1(_0102_),
    .A2(_0104_),
    .Y(_0105_),
    .B1(_0099_));
 sg13g2_a221oi_1 _4289_ (.B2(_0061_),
    .C1(net523),
    .B1(_0050_),
    .A1(_3269_),
    .Y(_0106_),
    .A2(_3271_));
 sg13g2_xnor2_1 _4290_ (.Y(_0107_),
    .A(_0069_),
    .B(_0106_));
 sg13g2_xor2_1 _4291_ (.B(_0106_),
    .A(_0069_),
    .X(_0109_));
 sg13g2_nor3_1 _4292_ (.A(_3272_),
    .B(net523),
    .C(_0070_),
    .Y(_0110_));
 sg13g2_xor2_1 _4293_ (.B(_0110_),
    .A(_0073_),
    .X(_0111_));
 sg13g2_o21ai_1 _4294_ (.B1(_0111_),
    .Y(_0112_),
    .A1(_0105_),
    .A2(_0107_));
 sg13g2_nand2_1 _4295_ (.Y(_0113_),
    .A(_0085_),
    .B(_0092_));
 sg13g2_a21oi_2 _4296_ (.B1(_0113_),
    .Y(_0114_),
    .A2(_0112_),
    .A1(_0090_));
 sg13g2_a21o_2 _4297_ (.A2(_0112_),
    .A1(_0090_),
    .B1(_0113_),
    .X(_0115_));
 sg13g2_nand2_2 _4298_ (.Y(_0116_),
    .A(_0083_),
    .B(_0115_));
 sg13g2_nand2_1 _4299_ (.Y(_0117_),
    .A(net510),
    .B(_0116_));
 sg13g2_nand2_1 _4300_ (.Y(_0118_),
    .A(_0109_),
    .B(_0111_));
 sg13g2_a21o_1 _4301_ (.A2(_0118_),
    .A1(_0095_),
    .B1(_0094_),
    .X(_0120_));
 sg13g2_or2_1 _4302_ (.X(_0121_),
    .B(_0092_),
    .A(_0087_));
 sg13g2_nand2_1 _4303_ (.Y(_0122_),
    .A(net502),
    .B(_0107_));
 sg13g2_nand3_1 _4304_ (.B(_0090_),
    .C(_0115_),
    .A(_0083_),
    .Y(_0123_));
 sg13g2_o21ai_1 _4305_ (.B1(_0111_),
    .Y(_0124_),
    .A1(_0084_),
    .A2(_0114_));
 sg13g2_nand2_1 _4306_ (.Y(_0125_),
    .A(_0123_),
    .B(_0124_));
 sg13g2_nand3_1 _4307_ (.B(_0123_),
    .C(_0124_),
    .A(_0094_),
    .Y(_0126_));
 sg13g2_o21ai_1 _4308_ (.B1(_0100_),
    .Y(_0127_),
    .A1(_0084_),
    .A2(_0114_));
 sg13g2_nand3_1 _4309_ (.B(_0109_),
    .C(_0115_),
    .A(_0083_),
    .Y(_0128_));
 sg13g2_nand3_1 _4310_ (.B(_0127_),
    .C(_0128_),
    .A(_0120_),
    .Y(_0129_));
 sg13g2_nand2_1 _4311_ (.Y(_0131_),
    .A(_0100_),
    .B(_0104_));
 sg13g2_nor2_1 _4312_ (.A(net510),
    .B(_0118_),
    .Y(_0132_));
 sg13g2_a21oi_1 _4313_ (.A1(_0131_),
    .A2(_0132_),
    .Y(_0133_),
    .B1(_0094_));
 sg13g2_inv_1 _4314_ (.Y(_0134_),
    .A(_0133_));
 sg13g2_and3_2 _4315_ (.X(_0135_),
    .A(_0121_),
    .B(_0122_),
    .C(_0126_));
 sg13g2_nand3_1 _4316_ (.B(_0122_),
    .C(_0126_),
    .A(_0121_),
    .Y(_0136_));
 sg13g2_or2_1 _4317_ (.X(_0137_),
    .B(_0102_),
    .A(net510));
 sg13g2_nand3_1 _4318_ (.B(_0111_),
    .C(_0115_),
    .A(_0083_),
    .Y(_0138_));
 sg13g2_o21ai_1 _4319_ (.B1(_0109_),
    .Y(_0139_),
    .A1(_0084_),
    .A2(_0114_));
 sg13g2_nand2_1 _4320_ (.Y(_0140_),
    .A(_0138_),
    .B(_0139_));
 sg13g2_nand3_1 _4321_ (.B(_0138_),
    .C(_0139_),
    .A(net512),
    .Y(_0142_));
 sg13g2_o21ai_1 _4322_ (.B1(_0104_),
    .Y(_0143_),
    .A1(_0084_),
    .A2(_0114_));
 sg13g2_nand3_1 _4323_ (.B(_0100_),
    .C(_0115_),
    .A(_0083_),
    .Y(_0144_));
 sg13g2_nand3_1 _4324_ (.B(_0143_),
    .C(_0144_),
    .A(_0094_),
    .Y(_0145_));
 sg13g2_nand3_1 _4325_ (.B(_0142_),
    .C(_0145_),
    .A(_0096_),
    .Y(_0146_));
 sg13g2_nand2_2 _4326_ (.Y(_0147_),
    .A(_0137_),
    .B(_0146_));
 sg13g2_nor2_1 _4327_ (.A(_0135_),
    .B(_0147_),
    .Y(_0148_));
 sg13g2_nand3_1 _4328_ (.B(_0137_),
    .C(_0146_),
    .A(_0136_),
    .Y(_0149_));
 sg13g2_nor2b_2 _4329_ (.A(net510),
    .B_N(_0111_),
    .Y(_0150_));
 sg13g2_nor2_1 _4330_ (.A(net510),
    .B(_0104_),
    .Y(_0151_));
 sg13g2_nand3_1 _4331_ (.B(_0129_),
    .C(_0134_),
    .A(_0121_),
    .Y(_0152_));
 sg13g2_nor2b_1 _4332_ (.A(_0120_),
    .B_N(_0133_),
    .Y(_0153_));
 sg13g2_a21oi_1 _4333_ (.A1(_0125_),
    .A2(_0153_),
    .Y(_0154_),
    .B1(_0095_));
 sg13g2_a21oi_2 _4334_ (.B1(_0151_),
    .Y(_0155_),
    .A2(_0154_),
    .A1(_0152_));
 sg13g2_nor2_1 _4335_ (.A(_0150_),
    .B(_0155_),
    .Y(_0156_));
 sg13g2_nor2_2 _4336_ (.A(_0135_),
    .B(_0155_),
    .Y(_0157_));
 sg13g2_inv_1 _4337_ (.Y(_0158_),
    .A(_0157_));
 sg13g2_nor2_2 _4338_ (.A(_0147_),
    .B(_0150_),
    .Y(_0159_));
 sg13g2_or2_1 _4339_ (.X(_0160_),
    .B(_0150_),
    .A(_0147_));
 sg13g2_nor2_1 _4340_ (.A(net512),
    .B(_0114_),
    .Y(_0161_));
 sg13g2_nor2_1 _4341_ (.A(_0094_),
    .B(_0116_),
    .Y(_0163_));
 sg13g2_a221oi_1 _4342_ (.B2(_0140_),
    .C1(_0163_),
    .B1(_0134_),
    .A1(_0090_),
    .Y(_0164_),
    .A2(_0116_));
 sg13g2_a21oi_1 _4343_ (.A1(net502),
    .A2(_0099_),
    .Y(_0165_),
    .B1(_0164_));
 sg13g2_nor2_1 _4344_ (.A(_0155_),
    .B(net484),
    .Y(_0166_));
 sg13g2_nor2_1 _4345_ (.A(_0147_),
    .B(net485),
    .Y(_0167_));
 sg13g2_nor2_1 _4346_ (.A(_0135_),
    .B(net485),
    .Y(_0168_));
 sg13g2_nor3_1 _4347_ (.A(_0149_),
    .B(_0155_),
    .C(net485),
    .Y(_0169_));
 sg13g2_nor2b_1 _4348_ (.A(net510),
    .B_N(_0054_),
    .Y(_0170_));
 sg13g2_nand2_2 _4349_ (.Y(_0171_),
    .A(_0054_),
    .B(net502));
 sg13g2_nor2_1 _4350_ (.A(_0150_),
    .B(_0170_),
    .Y(_0172_));
 sg13g2_o21ai_1 _4351_ (.B1(_0149_),
    .Y(_0174_),
    .A1(_0155_),
    .A2(net485));
 sg13g2_nor2b_1 _4352_ (.A(_0169_),
    .B_N(_0174_),
    .Y(_0175_));
 sg13g2_a21oi_2 _4353_ (.B1(_0169_),
    .Y(_0176_),
    .A2(_0174_),
    .A1(_0172_));
 sg13g2_xnor2_1 _4354_ (.Y(_0177_),
    .A(_0157_),
    .B(_0159_));
 sg13g2_nor2_1 _4355_ (.A(_0176_),
    .B(_0177_),
    .Y(_0178_));
 sg13g2_nand2_1 _4356_ (.Y(_0179_),
    .A(_0176_),
    .B(_0177_));
 sg13g2_nand2_1 _4357_ (.Y(_0180_),
    .A(_0158_),
    .B(net484));
 sg13g2_xnor2_1 _4358_ (.Y(_0181_),
    .A(_0157_),
    .B(net484));
 sg13g2_xnor2_1 _4359_ (.Y(_0182_),
    .A(_0160_),
    .B(_0181_));
 sg13g2_nor4_1 _4360_ (.A(_0158_),
    .B(_0160_),
    .C(net484),
    .D(_0176_),
    .Y(_0183_));
 sg13g2_a22oi_1 _4361_ (.Y(_0185_),
    .B1(_0181_),
    .B2(_0159_),
    .A2(_0166_),
    .A1(_0136_));
 sg13g2_a221oi_1 _4362_ (.B2(_0182_),
    .C1(_0178_),
    .B1(_0179_),
    .A1(_0157_),
    .Y(_0186_),
    .A2(_0159_));
 sg13g2_or2_1 _4363_ (.X(_0187_),
    .B(_0186_),
    .A(_0183_));
 sg13g2_nor2_1 _4364_ (.A(_0185_),
    .B(_0187_),
    .Y(_0188_));
 sg13g2_nor2_1 _4365_ (.A(_0183_),
    .B(_0188_),
    .Y(_0189_));
 sg13g2_and2_1 _4366_ (.A(_0136_),
    .B(net484),
    .X(_0190_));
 sg13g2_xnor2_1 _4367_ (.Y(_0191_),
    .A(_0156_),
    .B(_0190_));
 sg13g2_nor2_1 _4368_ (.A(_0189_),
    .B(_0191_),
    .Y(_0192_));
 sg13g2_xnor2_1 _4369_ (.Y(_0193_),
    .A(_0172_),
    .B(_0175_));
 sg13g2_mux2_1 _4370_ (.A0(_0193_),
    .A1(_0176_),
    .S(net484),
    .X(_0194_));
 sg13g2_xor2_1 _4371_ (.B(_0187_),
    .A(_0185_),
    .X(_0196_));
 sg13g2_nor2b_1 _4372_ (.A(_0194_),
    .B_N(_0196_),
    .Y(_0197_));
 sg13g2_xor2_1 _4373_ (.B(_0193_),
    .A(net484),
    .X(_0198_));
 sg13g2_a21oi_1 _4374_ (.A1(_0136_),
    .A2(_0171_),
    .Y(_0199_),
    .B1(_0167_));
 sg13g2_nor2_1 _4375_ (.A(net484),
    .B(_0170_),
    .Y(_0200_));
 sg13g2_nor2_1 _4376_ (.A(_0147_),
    .B(_0155_),
    .Y(_0201_));
 sg13g2_a21oi_1 _4377_ (.A1(_0148_),
    .A2(_0200_),
    .Y(_0202_),
    .B1(_0201_));
 sg13g2_nor2_1 _4378_ (.A(_0199_),
    .B(_0202_),
    .Y(_0203_));
 sg13g2_nand2_1 _4379_ (.Y(_0204_),
    .A(_0198_),
    .B(_0203_));
 sg13g2_nand2_1 _4380_ (.Y(_0205_),
    .A(_0166_),
    .B(_0171_));
 sg13g2_a21oi_1 _4381_ (.A1(_0148_),
    .A2(_0200_),
    .Y(_0207_),
    .B1(_0199_));
 sg13g2_xnor2_1 _4382_ (.Y(_0208_),
    .A(_0201_),
    .B(_0207_));
 sg13g2_or2_1 _4383_ (.X(_0209_),
    .B(_0208_),
    .A(_0205_));
 sg13g2_xor2_1 _4384_ (.B(_0203_),
    .A(_0198_),
    .X(_0210_));
 sg13g2_inv_1 _4385_ (.Y(_0211_),
    .A(_0210_));
 sg13g2_o21ai_1 _4386_ (.B1(_0204_),
    .Y(_0212_),
    .A1(_0209_),
    .A2(_0211_));
 sg13g2_xnor2_1 _4387_ (.Y(_0213_),
    .A(_0194_),
    .B(_0196_));
 sg13g2_a21oi_1 _4388_ (.A1(_0212_),
    .A2(_0213_),
    .Y(_0214_),
    .B1(_0197_));
 sg13g2_xor2_1 _4389_ (.B(_0191_),
    .A(_0189_),
    .X(_0215_));
 sg13g2_nor2b_1 _4390_ (.A(_0214_),
    .B_N(_0215_),
    .Y(_0216_));
 sg13g2_nor2_1 _4391_ (.A(_0192_),
    .B(_0216_),
    .Y(_0218_));
 sg13g2_xnor2_1 _4392_ (.Y(_0219_),
    .A(_0150_),
    .B(_0168_));
 sg13g2_nand2_1 _4393_ (.Y(_0220_),
    .A(_0180_),
    .B(_0219_));
 sg13g2_or2_1 _4394_ (.X(_0221_),
    .B(_0220_),
    .A(_0218_));
 sg13g2_a21oi_1 _4395_ (.A1(_0135_),
    .A2(_0221_),
    .Y(_0222_),
    .B1(_0150_));
 sg13g2_a21oi_1 _4396_ (.A1(_0135_),
    .A2(_0221_),
    .Y(_0223_),
    .B1(net493));
 sg13g2_xnor2_1 _4397_ (.Y(_0224_),
    .A(_0218_),
    .B(_0220_));
 sg13g2_o21ai_1 _4398_ (.B1(_0094_),
    .Y(_0225_),
    .A1(_0116_),
    .A2(_0224_));
 sg13g2_nor2_1 _4399_ (.A(_0223_),
    .B(_0225_),
    .Y(_0226_));
 sg13g2_xnor2_1 _4400_ (.Y(_0227_),
    .A(_0212_),
    .B(_0213_));
 sg13g2_xnor2_1 _4401_ (.Y(_0229_),
    .A(_0205_),
    .B(_0208_));
 sg13g2_mux2_1 _4402_ (.A0(_0227_),
    .A1(_0229_),
    .S(net493),
    .X(_0230_));
 sg13g2_a21oi_1 _4403_ (.A1(net512),
    .A2(_0230_),
    .Y(_0231_),
    .B1(net502));
 sg13g2_nor2b_2 _4404_ (.A(_0226_),
    .B_N(_0231_),
    .Y(_0232_));
 sg13g2_inv_2 _4405_ (.Y(_0233_),
    .A(_0232_));
 sg13g2_nand2_1 _4406_ (.Y(_0234_),
    .A(net470),
    .B(_0233_));
 sg13g2_xnor2_1 _4407_ (.Y(_0235_),
    .A(_0209_),
    .B(_0210_));
 sg13g2_xnor2_1 _4408_ (.Y(_0236_),
    .A(_0155_),
    .B(_0200_));
 sg13g2_o21ai_1 _4409_ (.B1(_0236_),
    .Y(_0237_),
    .A1(_0147_),
    .A2(_0171_));
 sg13g2_nand2_1 _4410_ (.Y(_0238_),
    .A(net493),
    .B(_0237_));
 sg13g2_o21ai_1 _4411_ (.B1(_0238_),
    .Y(_0239_),
    .A1(net493),
    .A2(_0235_));
 sg13g2_nand2b_1 _4412_ (.Y(_0240_),
    .B(_0221_),
    .A_N(_0190_));
 sg13g2_nor2_1 _4413_ (.A(_0150_),
    .B(_0240_),
    .Y(_0241_));
 sg13g2_xor2_1 _4414_ (.B(_0215_),
    .A(_0214_),
    .X(_0242_));
 sg13g2_nor2_1 _4415_ (.A(_0116_),
    .B(_0242_),
    .Y(_0243_));
 sg13g2_a21oi_1 _4416_ (.A1(net511),
    .A2(_0239_),
    .Y(_0244_),
    .B1(net502));
 sg13g2_nor2_1 _4417_ (.A(net511),
    .B(_0243_),
    .Y(_0245_));
 sg13g2_o21ai_1 _4418_ (.B1(_0245_),
    .Y(_0246_),
    .A1(_0117_),
    .A2(_0240_));
 sg13g2_nand2_2 _4419_ (.Y(_0247_),
    .A(_0244_),
    .B(_0246_));
 sg13g2_inv_2 _4420_ (.Y(_0248_),
    .A(_0247_));
 sg13g2_nand2_1 _4421_ (.Y(_0250_),
    .A(net468),
    .B(_0248_));
 sg13g2_xnor2_1 _4422_ (.Y(_0251_),
    .A(_2840_),
    .B(_0247_));
 sg13g2_mux2_1 _4423_ (.A0(_0224_),
    .A1(_0227_),
    .S(net493),
    .X(_0252_));
 sg13g2_nor2_1 _4424_ (.A(_0084_),
    .B(_0094_),
    .Y(_0253_));
 sg13g2_a221oi_1 _4425_ (.B2(_0094_),
    .C1(_0253_),
    .B1(_0252_),
    .A1(_0084_),
    .Y(_0254_),
    .A2(_0229_));
 sg13g2_a21o_2 _4426_ (.A2(_0222_),
    .A1(net502),
    .B1(_0254_),
    .X(_0255_));
 sg13g2_inv_2 _4427_ (.Y(_0256_),
    .A(_0255_));
 sg13g2_nor2_1 _4428_ (.A(_2856_),
    .B(_0256_),
    .Y(_0257_));
 sg13g2_nand2_1 _4429_ (.Y(_0258_),
    .A(net502),
    .B(_0241_));
 sg13g2_nand2_1 _4430_ (.Y(_0259_),
    .A(net493),
    .B(_0235_));
 sg13g2_o21ai_1 _4431_ (.B1(_0259_),
    .Y(_0261_),
    .A1(net493),
    .A2(_0242_));
 sg13g2_o21ai_1 _4432_ (.B1(net511),
    .Y(_0262_),
    .A1(net493),
    .A2(_0237_));
 sg13g2_o21ai_1 _4433_ (.B1(_0262_),
    .Y(_0263_),
    .A1(net511),
    .A2(_0261_));
 sg13g2_nand2_2 _4434_ (.Y(_0264_),
    .A(_0258_),
    .B(_0263_));
 sg13g2_nand2b_1 _4435_ (.Y(_0265_),
    .B(_0264_),
    .A_N(net475));
 sg13g2_xnor2_1 _4436_ (.Y(_0266_),
    .A(net475),
    .B(_0264_));
 sg13g2_nor2_1 _4437_ (.A(net510),
    .B(_0224_),
    .Y(_0267_));
 sg13g2_xor2_1 _4438_ (.B(_0155_),
    .A(_0147_),
    .X(_0268_));
 sg13g2_nand4_1 _4439_ (.B(_0116_),
    .C(_0171_),
    .A(net511),
    .Y(_0269_),
    .D(_0268_));
 sg13g2_o21ai_1 _4440_ (.B1(_0269_),
    .Y(_0270_),
    .A1(net511),
    .A2(_0230_));
 sg13g2_a21oi_2 _4441_ (.B1(_0267_),
    .Y(_0272_),
    .A2(_0270_),
    .A1(net510));
 sg13g2_nor2_1 _4442_ (.A(net472),
    .B(net469),
    .Y(_0273_));
 sg13g2_nor2_1 _4443_ (.A(net511),
    .B(_0239_),
    .Y(_0274_));
 sg13g2_nor2_1 _4444_ (.A(_0253_),
    .B(_0274_),
    .Y(_0275_));
 sg13g2_a21oi_2 _4445_ (.B1(_0275_),
    .Y(_0276_),
    .A2(_0242_),
    .A1(net502));
 sg13g2_inv_4 _4446_ (.A(_0276_),
    .Y(_0277_));
 sg13g2_nand2b_1 _4447_ (.Y(_0278_),
    .B(_0276_),
    .A_N(_2895_));
 sg13g2_xnor2_1 _4448_ (.Y(_0279_),
    .A(net472),
    .B(net469));
 sg13g2_inv_1 _4449_ (.Y(_0280_),
    .A(_0279_));
 sg13g2_nor2_1 _4450_ (.A(_0278_),
    .B(_0279_),
    .Y(_0281_));
 sg13g2_o21ai_1 _4451_ (.B1(_0266_),
    .Y(_0283_),
    .A1(_0273_),
    .A2(_0281_));
 sg13g2_nand2_1 _4452_ (.Y(_0284_),
    .A(_0265_),
    .B(_0283_));
 sg13g2_xnor2_1 _4453_ (.Y(_0285_),
    .A(_2856_),
    .B(_0255_));
 sg13g2_a21oi_2 _4454_ (.B1(_0257_),
    .Y(_0286_),
    .A2(_0285_),
    .A1(_0284_));
 sg13g2_o21ai_1 _4455_ (.B1(_0250_),
    .Y(_0287_),
    .A1(_0251_),
    .A2(_0286_));
 sg13g2_a22oi_1 _4456_ (.Y(_0288_),
    .B1(_0261_),
    .B2(_0088_),
    .A2(_0241_),
    .A1(_0161_));
 sg13g2_xnor2_1 _4457_ (.Y(_0289_),
    .A(_2912_),
    .B(_0288_));
 sg13g2_nand2b_1 _4458_ (.Y(_0290_),
    .B(_0289_),
    .A_N(_0287_));
 sg13g2_o21ai_1 _4459_ (.B1(_0289_),
    .Y(_0291_),
    .A1(net470),
    .A2(_0233_));
 sg13g2_nand3_1 _4460_ (.B(_0290_),
    .C(_0291_),
    .A(_0234_),
    .Y(_0292_));
 sg13g2_nor2b_1 _4461_ (.A(_0287_),
    .B_N(_0291_),
    .Y(_0294_));
 sg13g2_a21o_1 _4462_ (.A2(_0290_),
    .A1(_0234_),
    .B1(_0294_),
    .X(_0295_));
 sg13g2_nand3b_1 _4463_ (.B(_0292_),
    .C(_0295_),
    .Y(_0296_),
    .A_N(_2926_));
 sg13g2_xnor2_1 _4464_ (.Y(_0297_),
    .A(_0251_),
    .B(_0286_));
 sg13g2_xnor2_1 _4465_ (.Y(_0298_),
    .A(_0284_),
    .B(_0285_));
 sg13g2_nand2_1 _4466_ (.Y(_0299_),
    .A(_2895_),
    .B(_0277_));
 sg13g2_nand4_1 _4467_ (.B(_0278_),
    .C(_0280_),
    .A(_0266_),
    .Y(_0300_),
    .D(_0299_));
 sg13g2_nand2b_1 _4468_ (.Y(_0301_),
    .B(_0299_),
    .A_N(_0297_));
 sg13g2_or3_1 _4469_ (.A(_0266_),
    .B(_0273_),
    .C(_0281_),
    .X(_0302_));
 sg13g2_nand2_1 _4470_ (.Y(_0303_),
    .A(_0283_),
    .B(_0302_));
 sg13g2_a21o_1 _4471_ (.A2(_0300_),
    .A1(_0298_),
    .B1(_0297_),
    .X(_0305_));
 sg13g2_nand2b_2 _4472_ (.Y(_0306_),
    .B(_0305_),
    .A_N(_0296_));
 sg13g2_o21ai_1 _4473_ (.B1(_0306_),
    .Y(_0307_),
    .A1(_2922_),
    .A2(_2936_));
 sg13g2_nor2_1 _4474_ (.A(_3250_),
    .B(_0307_),
    .Y(_0308_));
 sg13g2_o21ai_1 _4475_ (.B1(_0184_),
    .Y(_0309_),
    .A1(net568),
    .A2(_2944_));
 sg13g2_nand2_2 _4476_ (.Y(_0310_),
    .A(_2923_),
    .B(_0309_));
 sg13g2_o21ai_1 _4477_ (.B1(_3048_),
    .Y(_0311_),
    .A1(_2579_),
    .A2(_2588_));
 sg13g2_o21ai_1 _4478_ (.B1(net596),
    .Y(_0312_),
    .A1(net598),
    .A2(net604));
 sg13g2_nand2b_1 _4479_ (.Y(_0313_),
    .B(net597),
    .A_N(net593));
 sg13g2_o21ai_1 _4480_ (.B1(net592),
    .Y(_0314_),
    .A1(net593),
    .A2(_0312_));
 sg13g2_nor2_1 _4481_ (.A(net590),
    .B(_0314_),
    .Y(_0316_));
 sg13g2_nor2_1 _4482_ (.A(_2587_),
    .B(_0314_),
    .Y(_0317_));
 sg13g2_nor2_1 _4483_ (.A(_3070_),
    .B(_0317_),
    .Y(_0318_));
 sg13g2_o21ai_1 _4484_ (.B1(net588),
    .Y(_0319_),
    .A1(_0075_),
    .A2(net533));
 sg13g2_nand2_1 _4485_ (.Y(_0320_),
    .A(_0013_),
    .B(_0319_));
 sg13g2_xnor2_1 _4486_ (.Y(_0321_),
    .A(_3125_),
    .B(_0320_));
 sg13g2_xnor2_1 _4487_ (.Y(_0322_),
    .A(_0019_),
    .B(_0320_));
 sg13g2_xnor2_1 _4488_ (.Y(_0323_),
    .A(net584),
    .B(_0319_));
 sg13g2_xnor2_1 _4489_ (.Y(_0324_),
    .A(_3070_),
    .B(_0319_));
 sg13g2_nand3_1 _4490_ (.B(_0053_),
    .C(net534),
    .A(net589),
    .Y(_0325_));
 sg13g2_nand2_1 _4491_ (.Y(_0327_),
    .A(net537),
    .B(_0325_));
 sg13g2_or2_1 _4492_ (.X(_0328_),
    .B(_0325_),
    .A(net537));
 sg13g2_xnor2_1 _4493_ (.Y(_0329_),
    .A(net587),
    .B(_0325_));
 sg13g2_inv_1 _4494_ (.Y(_0330_),
    .A(_0329_));
 sg13g2_o21ai_1 _4495_ (.B1(net589),
    .Y(_0331_),
    .A1(_0064_),
    .A2(net533));
 sg13g2_and2_2 _4496_ (.A(_2598_),
    .B(_0331_),
    .X(_0332_));
 sg13g2_nand2_2 _4497_ (.Y(_0333_),
    .A(_2598_),
    .B(_0331_));
 sg13g2_nor2_1 _4498_ (.A(_0329_),
    .B(_0333_),
    .Y(_0334_));
 sg13g2_o21ai_1 _4499_ (.B1(net592),
    .Y(_0335_),
    .A1(_3191_),
    .A2(net533));
 sg13g2_nand3b_1 _4500_ (.B(net534),
    .C(_0015_),
    .Y(_0336_),
    .A_N(net592));
 sg13g2_nand2_1 _4501_ (.Y(_0338_),
    .A(_0335_),
    .B(_0336_));
 sg13g2_a221oi_1 _4502_ (.B2(_0336_),
    .C1(_2640_),
    .B1(_0335_),
    .A1(net596),
    .Y(_0339_),
    .A2(net533));
 sg13g2_nand3_1 _4503_ (.B(_2624_),
    .C(_2626_),
    .A(_2615_),
    .Y(_0340_));
 sg13g2_nand2b_1 _4504_ (.Y(_0341_),
    .B(_3202_),
    .A_N(_2612_));
 sg13g2_nand4_1 _4505_ (.B(_2624_),
    .C(_2626_),
    .A(_2615_),
    .Y(_0342_),
    .D(_0341_));
 sg13g2_and2_1 _4506_ (.A(_0339_),
    .B(_0342_),
    .X(_0343_));
 sg13g2_a221oi_1 _4507_ (.B2(_0342_),
    .C1(_0333_),
    .B1(_0339_),
    .A1(_0327_),
    .Y(_0344_),
    .A2(_0328_));
 sg13g2_o21ai_1 _4508_ (.B1(_0322_),
    .Y(_0345_),
    .A1(net529),
    .A2(_0344_));
 sg13g2_nand3b_1 _4509_ (.B(_0323_),
    .C(_0321_),
    .Y(_0346_),
    .A_N(_0344_));
 sg13g2_and2_1 _4510_ (.A(net538),
    .B(_0346_),
    .X(_0347_));
 sg13g2_and3_2 _4511_ (.X(_0349_),
    .A(net538),
    .B(_0345_),
    .C(_0346_));
 sg13g2_o21ai_1 _4512_ (.B1(net546),
    .Y(_0350_),
    .A1(net582),
    .A2(_0318_));
 sg13g2_a21oi_2 _4513_ (.B1(_0350_),
    .Y(_0351_),
    .A2(_0318_),
    .A1(net582));
 sg13g2_or2_1 _4514_ (.X(_0352_),
    .B(_0351_),
    .A(_0349_));
 sg13g2_xnor2_1 _4515_ (.Y(_0353_),
    .A(_0013_),
    .B(_0317_));
 sg13g2_nand2_1 _4516_ (.Y(_0354_),
    .A(net547),
    .B(_0353_));
 sg13g2_xnor2_1 _4517_ (.Y(_0355_),
    .A(_0323_),
    .B(_0344_));
 sg13g2_o21ai_1 _4518_ (.B1(_0354_),
    .Y(_0356_),
    .A1(net546),
    .A2(_0355_));
 sg13g2_nand2b_1 _4519_ (.Y(_0357_),
    .B(_0356_),
    .A_N(_0352_));
 sg13g2_inv_1 _4520_ (.Y(_0358_),
    .A(_0357_));
 sg13g2_nand2_1 _4521_ (.Y(_0360_),
    .A(_3191_),
    .B(net533));
 sg13g2_xnor2_1 _4522_ (.Y(_0361_),
    .A(_3191_),
    .B(net534));
 sg13g2_a21oi_1 _4523_ (.A1(_0342_),
    .A2(_0361_),
    .Y(_0362_),
    .B1(_0338_));
 sg13g2_and2_1 _4524_ (.A(net592),
    .B(_0361_),
    .X(_0363_));
 sg13g2_a21o_1 _4525_ (.A2(_0363_),
    .A1(_0342_),
    .B1(net560),
    .X(_0364_));
 sg13g2_o21ai_1 _4526_ (.B1(net548),
    .Y(_0365_),
    .A1(net593),
    .A2(_0312_));
 sg13g2_a21o_1 _4527_ (.A2(_0312_),
    .A1(net593),
    .B1(_0365_),
    .X(_0366_));
 sg13g2_o21ai_1 _4528_ (.B1(_0366_),
    .Y(_0367_),
    .A1(_0362_),
    .A2(_0364_));
 sg13g2_and2_1 _4529_ (.A(net599),
    .B(net602),
    .X(_0368_));
 sg13g2_nand2_1 _4530_ (.Y(_0369_),
    .A(net599),
    .B(net602));
 sg13g2_o21ai_1 _4531_ (.B1(net551),
    .Y(_0371_),
    .A1(net599),
    .A2(net601));
 sg13g2_nor2_2 _4532_ (.A(_0368_),
    .B(_0371_),
    .Y(_0372_));
 sg13g2_xnor2_1 _4533_ (.Y(_0373_),
    .A(_2610_),
    .B(_2627_));
 sg13g2_a21oi_2 _4534_ (.B1(_0372_),
    .Y(_0374_),
    .A2(_0373_),
    .A1(net538));
 sg13g2_xnor2_1 _4535_ (.Y(_0375_),
    .A(net546),
    .B(net607));
 sg13g2_xor2_1 _4536_ (.B(net607),
    .A(net546),
    .X(_0376_));
 sg13g2_nand2_1 _4537_ (.Y(_0377_),
    .A(net551),
    .B(_0000_));
 sg13g2_nor2b_2 _4538_ (.A(_0051_),
    .B_N(_0377_),
    .Y(_0378_));
 sg13g2_nor2_1 _4539_ (.A(_0375_),
    .B(_0378_),
    .Y(_0379_));
 sg13g2_nand2_2 _4540_ (.Y(_0380_),
    .A(net604),
    .B(_0379_));
 sg13g2_inv_1 _4541_ (.Y(_0382_),
    .A(_0380_));
 sg13g2_nor2_1 _4542_ (.A(_0374_),
    .B(_0380_),
    .Y(_0383_));
 sg13g2_nand3_1 _4543_ (.B(_2639_),
    .C(_0312_),
    .A(net548),
    .Y(_0384_));
 sg13g2_xnor2_1 _4544_ (.Y(_0385_),
    .A(_2641_),
    .B(_0342_));
 sg13g2_o21ai_1 _4545_ (.B1(_0384_),
    .Y(_0386_),
    .A1(net546),
    .A2(_0385_));
 sg13g2_nor3_1 _4546_ (.A(_0374_),
    .B(_0380_),
    .C(_0386_),
    .Y(_0387_));
 sg13g2_nor4_2 _4547_ (.A(_0367_),
    .B(_0374_),
    .C(_0380_),
    .Y(_0388_),
    .D(_0386_));
 sg13g2_xnor2_1 _4548_ (.Y(_0389_),
    .A(_0333_),
    .B(_0343_));
 sg13g2_o21ai_1 _4549_ (.B1(net548),
    .Y(_0390_),
    .A1(net589),
    .A2(_0314_));
 sg13g2_a21oi_1 _4550_ (.A1(net589),
    .A2(_0314_),
    .Y(_0391_),
    .B1(_0390_));
 sg13g2_a21oi_2 _4551_ (.B1(_0391_),
    .Y(_0393_),
    .A2(_0389_),
    .A1(net538));
 sg13g2_nand2_1 _4552_ (.Y(_0394_),
    .A(_0388_),
    .B(_0393_));
 sg13g2_o21ai_1 _4553_ (.B1(_0329_),
    .Y(_0395_),
    .A1(_0333_),
    .A2(_0343_));
 sg13g2_nor2_1 _4554_ (.A(net547),
    .B(_0344_),
    .Y(_0396_));
 sg13g2_xnor2_1 _4555_ (.Y(_0397_),
    .A(_3224_),
    .B(_0316_));
 sg13g2_a22oi_1 _4556_ (.Y(_0398_),
    .B1(_0397_),
    .B2(net547),
    .A2(_0396_),
    .A1(_0395_));
 sg13g2_nor2_1 _4557_ (.A(_0394_),
    .B(_0398_),
    .Y(_0399_));
 sg13g2_nor2_1 _4558_ (.A(_0352_),
    .B(_0399_),
    .Y(_0400_));
 sg13g2_mux2_2 _4559_ (.A0(_0400_),
    .A1(_0352_),
    .S(_0356_),
    .X(_0401_));
 sg13g2_o21ai_1 _4560_ (.B1(_0357_),
    .Y(_0402_),
    .A1(_0356_),
    .A2(_0400_));
 sg13g2_nor3_2 _4561_ (.A(_0349_),
    .B(_0351_),
    .C(_0382_),
    .Y(_0404_));
 sg13g2_xor2_1 _4562_ (.B(_0404_),
    .A(_0374_),
    .X(_0405_));
 sg13g2_xnor2_1 _4563_ (.Y(_0406_),
    .A(_0374_),
    .B(_0404_));
 sg13g2_nor3_2 _4564_ (.A(_0349_),
    .B(_0351_),
    .C(_0379_),
    .Y(_0407_));
 sg13g2_xnor2_1 _4565_ (.Y(_0408_),
    .A(net604),
    .B(_0407_));
 sg13g2_xor2_1 _4566_ (.B(_0407_),
    .A(net604),
    .X(_0409_));
 sg13g2_nor3_1 _4567_ (.A(_0349_),
    .B(_0351_),
    .C(_0387_),
    .Y(_0410_));
 sg13g2_xor2_1 _4568_ (.B(_0410_),
    .A(_0367_),
    .X(_0411_));
 sg13g2_xnor2_1 _4569_ (.Y(_0412_),
    .A(_0367_),
    .B(_0410_));
 sg13g2_nor3_2 _4570_ (.A(_0349_),
    .B(_0351_),
    .C(_0383_),
    .Y(_0413_));
 sg13g2_xor2_1 _4571_ (.B(_0413_),
    .A(_0386_),
    .X(_0415_));
 sg13g2_xnor2_1 _4572_ (.Y(_0416_),
    .A(_0386_),
    .B(_0413_));
 sg13g2_nor2_1 _4573_ (.A(_0411_),
    .B(_0415_),
    .Y(_0417_));
 sg13g2_o21ai_1 _4574_ (.B1(_0417_),
    .Y(_0418_),
    .A1(_0405_),
    .A2(_0408_));
 sg13g2_a221oi_1 _4575_ (.B2(_0393_),
    .C1(_0351_),
    .B1(_0388_),
    .A1(_0345_),
    .Y(_0419_),
    .A2(_0347_));
 sg13g2_xnor2_1 _4576_ (.Y(_0420_),
    .A(_0398_),
    .B(_0419_));
 sg13g2_nor3_1 _4577_ (.A(_0349_),
    .B(_0351_),
    .C(_0388_),
    .Y(_0421_));
 sg13g2_xor2_1 _4578_ (.B(_0421_),
    .A(_0393_),
    .X(_0422_));
 sg13g2_inv_1 _4579_ (.Y(_0423_),
    .A(_0422_));
 sg13g2_and2_1 _4580_ (.A(_0420_),
    .B(_0422_),
    .X(_0424_));
 sg13g2_nand2_1 _4581_ (.Y(_0426_),
    .A(_0420_),
    .B(_0422_));
 sg13g2_mux2_1 _4582_ (.A0(_2618_),
    .A1(_0378_),
    .S(_0352_),
    .X(_0427_));
 sg13g2_a21o_1 _4583_ (.A2(_0427_),
    .A1(_0409_),
    .B1(_0405_),
    .X(_0428_));
 sg13g2_a21oi_1 _4584_ (.A1(_0416_),
    .A2(_0428_),
    .Y(_0429_),
    .B1(_0411_));
 sg13g2_o21ai_1 _4585_ (.B1(_0420_),
    .Y(_0430_),
    .A1(_0423_),
    .A2(_0429_));
 sg13g2_and2_1 _4586_ (.A(net501),
    .B(_0430_),
    .X(_0431_));
 sg13g2_nand2_2 _4587_ (.Y(_0432_),
    .A(net501),
    .B(_0430_));
 sg13g2_a21oi_1 _4588_ (.A1(_0418_),
    .A2(_0424_),
    .Y(_0433_),
    .B1(_0402_));
 sg13g2_and2_1 _4589_ (.A(_0417_),
    .B(_0424_),
    .X(_0434_));
 sg13g2_inv_1 _4590_ (.Y(_0435_),
    .A(_0434_));
 sg13g2_nand3_1 _4591_ (.B(_0433_),
    .C(_0435_),
    .A(_0430_),
    .Y(_0437_));
 sg13g2_and2_1 _4592_ (.A(net501),
    .B(_0437_),
    .X(_0438_));
 sg13g2_nand2_2 _4593_ (.Y(_0439_),
    .A(net501),
    .B(_0437_));
 sg13g2_nor3_2 _4594_ (.A(_0357_),
    .B(_0394_),
    .C(_0398_),
    .Y(_0440_));
 sg13g2_a21oi_1 _4595_ (.A1(net501),
    .A2(_0430_),
    .Y(_0441_),
    .B1(_0440_));
 sg13g2_mux2_1 _4596_ (.A0(_0422_),
    .A1(_0420_),
    .S(_0441_),
    .X(_0442_));
 sg13g2_o21ai_1 _4597_ (.B1(_0442_),
    .Y(_0443_),
    .A1(_0412_),
    .A2(_0439_));
 sg13g2_a221oi_1 _4598_ (.B2(_0430_),
    .C1(_0433_),
    .B1(net501),
    .A1(_0358_),
    .Y(_0444_),
    .A2(_0399_));
 sg13g2_a22oi_1 _4599_ (.Y(_0445_),
    .B1(_0435_),
    .B2(_0401_),
    .A2(_0433_),
    .A1(_0430_));
 sg13g2_a22oi_1 _4600_ (.Y(_0446_),
    .B1(_0444_),
    .B2(_0445_),
    .A2(_0431_),
    .A1(_0426_));
 sg13g2_mux2_1 _4601_ (.A0(_0406_),
    .A1(_0416_),
    .S(net492),
    .X(_0448_));
 sg13g2_or2_1 _4602_ (.X(_0449_),
    .B(_0448_),
    .A(_0446_));
 sg13g2_nand3_1 _4603_ (.B(_0408_),
    .C(_0437_),
    .A(_0401_),
    .Y(_0450_));
 sg13g2_o21ai_1 _4604_ (.B1(_0450_),
    .Y(_0451_),
    .A1(_0446_),
    .A2(_0448_));
 sg13g2_and2_1 _4605_ (.A(_0443_),
    .B(_0451_),
    .X(_0452_));
 sg13g2_nand2_2 _4606_ (.Y(_0453_),
    .A(_0422_),
    .B(net489));
 sg13g2_nor2_1 _4607_ (.A(_0406_),
    .B(_0439_),
    .Y(_0454_));
 sg13g2_nand2_1 _4608_ (.Y(_0455_),
    .A(_0405_),
    .B(_0438_));
 sg13g2_a21oi_2 _4609_ (.B1(_0440_),
    .Y(_0456_),
    .A2(_0437_),
    .A1(net501));
 sg13g2_or2_2 _4610_ (.X(_0457_),
    .B(_0440_),
    .A(net489));
 sg13g2_mux2_1 _4611_ (.A0(_0415_),
    .A1(_0411_),
    .S(net492),
    .X(_0459_));
 sg13g2_or2_1 _4612_ (.X(_0460_),
    .B(_0459_),
    .A(_0446_));
 sg13g2_o21ai_1 _4613_ (.B1(_0456_),
    .Y(_0461_),
    .A1(_0446_),
    .A2(_0459_));
 sg13g2_nand2_2 _4614_ (.Y(_0462_),
    .A(_0455_),
    .B(_0461_));
 sg13g2_nand2_1 _4615_ (.Y(_0463_),
    .A(net483),
    .B(_0462_));
 sg13g2_inv_1 _4616_ (.Y(_0464_),
    .A(_0463_));
 sg13g2_nand2_1 _4617_ (.Y(_0465_),
    .A(_0451_),
    .B(net483));
 sg13g2_inv_1 _4618_ (.Y(_0466_),
    .A(_0465_));
 sg13g2_and2_1 _4619_ (.A(_0443_),
    .B(_0462_),
    .X(_0467_));
 sg13g2_nand2_1 _4620_ (.Y(_0468_),
    .A(_0466_),
    .B(_0467_));
 sg13g2_mux2_1 _4621_ (.A0(_0411_),
    .A1(_0423_),
    .S(net492),
    .X(_0470_));
 sg13g2_nand3_1 _4622_ (.B(_0416_),
    .C(_0437_),
    .A(_0401_),
    .Y(_0471_));
 sg13g2_o21ai_1 _4623_ (.B1(_0471_),
    .Y(_0472_),
    .A1(_0438_),
    .A2(_0470_));
 sg13g2_mux2_1 _4624_ (.A0(_0415_),
    .A1(_0470_),
    .S(_0439_),
    .X(_0473_));
 sg13g2_nand2_1 _4625_ (.Y(_0474_),
    .A(net483),
    .B(net482));
 sg13g2_nand2_1 _4626_ (.Y(_0475_),
    .A(_0443_),
    .B(_0472_));
 sg13g2_nand2_1 _4627_ (.Y(_0476_),
    .A(_0474_),
    .B(_0475_));
 sg13g2_nand2_1 _4628_ (.Y(_0477_),
    .A(_0468_),
    .B(_0476_));
 sg13g2_or2_1 _4629_ (.X(_0478_),
    .B(_0463_),
    .A(_0452_));
 sg13g2_xnor2_1 _4630_ (.Y(_0479_),
    .A(_0466_),
    .B(_0467_));
 sg13g2_a21o_1 _4631_ (.A2(net482),
    .A1(_0462_),
    .B1(_0452_),
    .X(_0481_));
 sg13g2_nand2_1 _4632_ (.Y(_0482_),
    .A(_0443_),
    .B(net482));
 sg13g2_a22oi_1 _4633_ (.Y(_0483_),
    .B1(_0455_),
    .B2(_0461_),
    .A2(_0450_),
    .A1(_0449_));
 sg13g2_nand2_1 _4634_ (.Y(_0484_),
    .A(_0467_),
    .B(net482));
 sg13g2_nor2b_2 _4635_ (.A(_0482_),
    .B_N(net478),
    .Y(_0485_));
 sg13g2_nand3_1 _4636_ (.B(_0427_),
    .C(_0437_),
    .A(net501),
    .Y(_0486_));
 sg13g2_mux2_1 _4637_ (.A0(_0409_),
    .A1(_0406_),
    .S(net492),
    .X(_0487_));
 sg13g2_o21ai_1 _4638_ (.B1(_0486_),
    .Y(_0488_),
    .A1(_0446_),
    .A2(_0487_));
 sg13g2_nand2_2 _4639_ (.Y(_0489_),
    .A(_0453_),
    .B(_0488_));
 sg13g2_inv_1 _4640_ (.Y(_0490_),
    .A(_0489_));
 sg13g2_nor2_1 _4641_ (.A(_0485_),
    .B(_0490_),
    .Y(_0492_));
 sg13g2_a21oi_1 _4642_ (.A1(_0481_),
    .A2(_0490_),
    .Y(_0493_),
    .B1(_0485_));
 sg13g2_or2_1 _4643_ (.X(_0494_),
    .B(_0493_),
    .A(_0479_));
 sg13g2_xnor2_1 _4644_ (.Y(_0495_),
    .A(_0467_),
    .B(_0472_));
 sg13g2_inv_1 _4645_ (.Y(_0496_),
    .A(_0495_));
 sg13g2_xnor2_1 _4646_ (.Y(_0497_),
    .A(_0479_),
    .B(_0493_));
 sg13g2_o21ai_1 _4647_ (.B1(_0494_),
    .Y(_0498_),
    .A1(_0496_),
    .A2(_0497_));
 sg13g2_nand2b_1 _4648_ (.Y(_0499_),
    .B(_0498_),
    .A_N(_0478_));
 sg13g2_xor2_1 _4649_ (.B(_0498_),
    .A(_0478_),
    .X(_0500_));
 sg13g2_o21ai_1 _4650_ (.B1(_0499_),
    .Y(_0501_),
    .A1(_0484_),
    .A2(_0500_));
 sg13g2_nand2b_1 _4651_ (.Y(_0503_),
    .B(_0501_),
    .A_N(_0477_));
 sg13g2_xnor2_1 _4652_ (.Y(_0504_),
    .A(_0477_),
    .B(_0501_));
 sg13g2_nand2b_1 _4653_ (.Y(_0505_),
    .B(_0504_),
    .A_N(_0474_));
 sg13g2_nor2_1 _4654_ (.A(_0468_),
    .B(net482),
    .Y(_0506_));
 sg13g2_a21oi_1 _4655_ (.A1(net483),
    .A2(net478),
    .Y(_0507_),
    .B1(_0482_));
 sg13g2_nor2_1 _4656_ (.A(_0506_),
    .B(_0507_),
    .Y(_0508_));
 sg13g2_a21oi_1 _4657_ (.A1(_0503_),
    .A2(_0505_),
    .Y(_0509_),
    .B1(_0508_));
 sg13g2_nand2_1 _4658_ (.Y(_0510_),
    .A(_0451_),
    .B(_0473_));
 sg13g2_a221oi_1 _4659_ (.B2(_0461_),
    .C1(_0472_),
    .B1(_0455_),
    .A1(_0449_),
    .Y(_0511_),
    .A2(_0450_));
 sg13g2_nand2_1 _4660_ (.Y(_0512_),
    .A(net482),
    .B(net478));
 sg13g2_nand2_2 _4661_ (.Y(_0514_),
    .A(_0443_),
    .B(_0488_));
 sg13g2_a221oi_1 _4662_ (.B2(_0451_),
    .C1(_0454_),
    .B1(net482),
    .A1(_0456_),
    .Y(_0515_),
    .A2(_0460_));
 sg13g2_or3_2 _4663_ (.A(_0511_),
    .B(_0514_),
    .C(_0515_),
    .X(_0516_));
 sg13g2_nand2_1 _4664_ (.Y(_0517_),
    .A(_0512_),
    .B(_0516_));
 sg13g2_and2_1 _4665_ (.A(_0481_),
    .B(_0492_),
    .X(_0518_));
 sg13g2_a21o_1 _4666_ (.A2(_0517_),
    .A1(_0490_),
    .B1(_0518_),
    .X(_0519_));
 sg13g2_xnor2_1 _4667_ (.Y(_0520_),
    .A(_0495_),
    .B(_0497_));
 sg13g2_xor2_1 _4668_ (.B(_0520_),
    .A(_0519_),
    .X(_0521_));
 sg13g2_a22oi_1 _4669_ (.Y(_0522_),
    .B1(_0521_),
    .B2(_0485_),
    .A2(_0520_),
    .A1(_0519_));
 sg13g2_xnor2_1 _4670_ (.Y(_0523_),
    .A(_0484_),
    .B(_0500_));
 sg13g2_nor2_1 _4671_ (.A(_0522_),
    .B(_0523_),
    .Y(_0525_));
 sg13g2_xor2_1 _4672_ (.B(_0523_),
    .A(_0522_),
    .X(_0526_));
 sg13g2_a21oi_1 _4673_ (.A1(_0464_),
    .A2(_0526_),
    .Y(_0527_),
    .B1(_0525_));
 sg13g2_xor2_1 _4674_ (.B(_0504_),
    .A(_0474_),
    .X(_0528_));
 sg13g2_nor2_1 _4675_ (.A(_0527_),
    .B(_0528_),
    .Y(_0529_));
 sg13g2_o21ai_1 _4676_ (.B1(_0514_),
    .Y(_0530_),
    .A1(_0511_),
    .A2(_0515_));
 sg13g2_nand3_1 _4677_ (.B(_0516_),
    .C(_0530_),
    .A(net478),
    .Y(_0531_));
 sg13g2_nand2_2 _4678_ (.Y(_0532_),
    .A(_0376_),
    .B(_0438_));
 sg13g2_nand2_1 _4679_ (.Y(_0533_),
    .A(net482),
    .B(_0532_));
 sg13g2_nand2_2 _4680_ (.Y(_0534_),
    .A(_0453_),
    .B(_0532_));
 sg13g2_xor2_1 _4681_ (.B(_0534_),
    .A(_0510_),
    .X(_0536_));
 sg13g2_nand2b_1 _4682_ (.Y(_0537_),
    .B(_0536_),
    .A_N(_0514_));
 sg13g2_xnor2_1 _4683_ (.Y(_0538_),
    .A(_0514_),
    .B(_0536_));
 sg13g2_xor2_1 _4684_ (.B(_0536_),
    .A(_0514_),
    .X(_0539_));
 sg13g2_a21oi_1 _4685_ (.A1(_0516_),
    .A2(_0530_),
    .Y(_0540_),
    .B1(net478));
 sg13g2_a21o_1 _4686_ (.A2(_0530_),
    .A1(_0516_),
    .B1(net478),
    .X(_0541_));
 sg13g2_and3_1 _4687_ (.X(_0542_),
    .A(_0531_),
    .B(_0538_),
    .C(_0541_));
 sg13g2_o21ai_1 _4688_ (.B1(_0531_),
    .Y(_0543_),
    .A1(_0539_),
    .A2(_0540_));
 sg13g2_xnor2_1 _4689_ (.Y(_0544_),
    .A(_0489_),
    .B(_0517_));
 sg13g2_o21ai_1 _4690_ (.B1(_0537_),
    .Y(_0545_),
    .A1(_0510_),
    .A2(_0534_));
 sg13g2_xnor2_1 _4691_ (.Y(_0547_),
    .A(_0543_),
    .B(_0544_));
 sg13g2_nor2b_1 _4692_ (.A(_0547_),
    .B_N(_0545_),
    .Y(_0548_));
 sg13g2_a21oi_1 _4693_ (.A1(_0543_),
    .A2(_0544_),
    .Y(_0549_),
    .B1(_0548_));
 sg13g2_xnor2_1 _4694_ (.Y(_0550_),
    .A(_0485_),
    .B(_0521_));
 sg13g2_nor2_1 _4695_ (.A(_0549_),
    .B(_0550_),
    .Y(_0551_));
 sg13g2_xor2_1 _4696_ (.B(_0550_),
    .A(_0549_),
    .X(_0552_));
 sg13g2_a21oi_1 _4697_ (.A1(_0466_),
    .A2(_0552_),
    .Y(_0553_),
    .B1(_0551_));
 sg13g2_xnor2_1 _4698_ (.Y(_0554_),
    .A(_0464_),
    .B(_0526_));
 sg13g2_or2_1 _4699_ (.X(_0555_),
    .B(_0554_),
    .A(_0553_));
 sg13g2_nand2_1 _4700_ (.Y(_0556_),
    .A(_0473_),
    .B(_0488_));
 sg13g2_a21oi_1 _4701_ (.A1(_0531_),
    .A2(_0541_),
    .Y(_0558_),
    .B1(_0538_));
 sg13g2_nor3_1 _4702_ (.A(_0542_),
    .B(_0556_),
    .C(_0558_),
    .Y(_0559_));
 sg13g2_or3_1 _4703_ (.A(_0542_),
    .B(_0556_),
    .C(_0558_),
    .X(_0560_));
 sg13g2_and2_1 _4704_ (.A(_0443_),
    .B(_0532_),
    .X(_0561_));
 sg13g2_o21ai_1 _4705_ (.B1(_0556_),
    .Y(_0562_),
    .A1(_0542_),
    .A2(_0558_));
 sg13g2_nand3_1 _4706_ (.B(_0561_),
    .C(_0562_),
    .A(_0560_),
    .Y(_0563_));
 sg13g2_a21oi_1 _4707_ (.A1(_0561_),
    .A2(_0562_),
    .Y(_0564_),
    .B1(_0559_));
 sg13g2_xor2_1 _4708_ (.B(_0547_),
    .A(_0545_),
    .X(_0565_));
 sg13g2_nor2_1 _4709_ (.A(_0564_),
    .B(_0565_),
    .Y(_0566_));
 sg13g2_xor2_1 _4710_ (.B(_0565_),
    .A(_0564_),
    .X(_0567_));
 sg13g2_a21oi_1 _4711_ (.A1(_0490_),
    .A2(_0567_),
    .Y(_0569_),
    .B1(_0566_));
 sg13g2_xnor2_1 _4712_ (.Y(_0570_),
    .A(_0465_),
    .B(_0552_));
 sg13g2_nor2b_1 _4713_ (.A(_0569_),
    .B_N(_0570_),
    .Y(_0571_));
 sg13g2_xor2_1 _4714_ (.B(_0462_),
    .A(_0451_),
    .X(_0572_));
 sg13g2_nand2_1 _4715_ (.Y(_0573_),
    .A(_0488_),
    .B(_0572_));
 sg13g2_nand2_1 _4716_ (.Y(_0574_),
    .A(_0483_),
    .B(_0488_));
 sg13g2_o21ai_1 _4717_ (.B1(_0574_),
    .Y(_0575_),
    .A1(_0533_),
    .A2(_0573_));
 sg13g2_a21o_1 _4718_ (.A2(_0562_),
    .A1(_0560_),
    .B1(_0561_),
    .X(_0576_));
 sg13g2_nand3_1 _4719_ (.B(_0575_),
    .C(_0576_),
    .A(_0563_),
    .Y(_0577_));
 sg13g2_a21oi_1 _4720_ (.A1(_0563_),
    .A2(_0576_),
    .Y(_0578_),
    .B1(_0575_));
 sg13g2_a21o_1 _4721_ (.A2(_0576_),
    .A1(_0563_),
    .B1(_0575_),
    .X(_0580_));
 sg13g2_and4_1 _4722_ (.A(_0453_),
    .B(_0532_),
    .C(_0577_),
    .D(_0580_),
    .X(_0581_));
 sg13g2_o21ai_1 _4723_ (.B1(_0577_),
    .Y(_0582_),
    .A1(_0534_),
    .A2(_0578_));
 sg13g2_xnor2_1 _4724_ (.Y(_0583_),
    .A(_0489_),
    .B(_0567_));
 sg13g2_and2_1 _4725_ (.A(_0582_),
    .B(_0583_),
    .X(_0584_));
 sg13g2_xor2_1 _4726_ (.B(_0573_),
    .A(_0533_),
    .X(_0585_));
 sg13g2_nand2_1 _4727_ (.Y(_0586_),
    .A(net478),
    .B(_0532_));
 sg13g2_and3_1 _4728_ (.X(_0587_),
    .A(net478),
    .B(_0532_),
    .C(_0585_));
 sg13g2_inv_1 _4729_ (.Y(_0588_),
    .A(_0587_));
 sg13g2_a22oi_1 _4730_ (.Y(_0589_),
    .B1(_0577_),
    .B2(_0580_),
    .A2(_0532_),
    .A1(net483));
 sg13g2_nor3_2 _4731_ (.A(_0581_),
    .B(_0588_),
    .C(_0589_),
    .Y(_0591_));
 sg13g2_or2_1 _4732_ (.X(_0592_),
    .B(_0583_),
    .A(_0582_));
 sg13g2_nand2b_1 _4733_ (.Y(_0593_),
    .B(_0592_),
    .A_N(_0584_));
 sg13g2_a21o_1 _4734_ (.A2(_0592_),
    .A1(_0591_),
    .B1(_0584_),
    .X(_0594_));
 sg13g2_xnor2_1 _4735_ (.Y(_0595_),
    .A(_0569_),
    .B(_0570_));
 sg13g2_a21oi_1 _4736_ (.A1(_0594_),
    .A2(_0595_),
    .Y(_0596_),
    .B1(_0571_));
 sg13g2_xor2_1 _4737_ (.B(_0554_),
    .A(_0553_),
    .X(_0597_));
 sg13g2_inv_1 _4738_ (.Y(_0598_),
    .A(_0597_));
 sg13g2_o21ai_1 _4739_ (.B1(_0555_),
    .Y(_0599_),
    .A1(_0596_),
    .A2(_0598_));
 sg13g2_xor2_1 _4740_ (.B(_0528_),
    .A(_0527_),
    .X(_0600_));
 sg13g2_a21o_1 _4741_ (.A2(_0600_),
    .A1(_0599_),
    .B1(_0529_),
    .X(_0602_));
 sg13g2_nand3_1 _4742_ (.B(_0505_),
    .C(_0508_),
    .A(_0503_),
    .Y(_0603_));
 sg13g2_nor2b_1 _4743_ (.A(_0509_),
    .B_N(_0603_),
    .Y(_0604_));
 sg13g2_a21oi_2 _4744_ (.B1(_0509_),
    .Y(_0605_),
    .A2(_0604_),
    .A1(_0602_));
 sg13g2_nand2_1 _4745_ (.Y(_0606_),
    .A(_0443_),
    .B(_0512_));
 sg13g2_nand2_1 _4746_ (.Y(_0607_),
    .A(net483),
    .B(_0606_));
 sg13g2_xor2_1 _4747_ (.B(_0607_),
    .A(_0605_),
    .X(_0608_));
 sg13g2_xnor2_1 _4748_ (.Y(_0609_),
    .A(_0599_),
    .B(_0600_));
 sg13g2_nand2_1 _4749_ (.Y(_0610_),
    .A(_0431_),
    .B(_0609_));
 sg13g2_xnor2_1 _4750_ (.Y(_0611_),
    .A(_0594_),
    .B(_0595_));
 sg13g2_a21oi_1 _4751_ (.A1(_0432_),
    .A2(_0611_),
    .Y(_0613_),
    .B1(_0457_));
 sg13g2_nor2_2 _4752_ (.A(net489),
    .B(net492),
    .Y(_0614_));
 sg13g2_a22oi_1 _4753_ (.Y(_0615_),
    .B1(_0610_),
    .B2(_0613_),
    .A2(_0608_),
    .A1(net489));
 sg13g2_nor2_1 _4754_ (.A(_0256_),
    .B(_0615_),
    .Y(_0616_));
 sg13g2_nand2b_1 _4755_ (.Y(_0617_),
    .B(_0614_),
    .A_N(_0608_));
 sg13g2_a21oi_2 _4756_ (.B1(_0457_),
    .Y(_0618_),
    .A2(_0609_),
    .A1(_0432_));
 sg13g2_nand2_2 _4757_ (.Y(_0619_),
    .A(_0617_),
    .B(_0618_));
 sg13g2_xnor2_1 _4758_ (.Y(_0620_),
    .A(_0255_),
    .B(_0615_));
 sg13g2_a21oi_1 _4759_ (.A1(_0619_),
    .A2(_0620_),
    .Y(_0621_),
    .B1(_0616_));
 sg13g2_nand2b_1 _4760_ (.Y(_0622_),
    .B(_0605_),
    .A_N(_0443_));
 sg13g2_nand2_1 _4761_ (.Y(_0624_),
    .A(net483),
    .B(_0622_));
 sg13g2_xnor2_1 _4762_ (.Y(_0625_),
    .A(_0596_),
    .B(_0597_));
 sg13g2_a21oi_1 _4763_ (.A1(_0432_),
    .A2(_0625_),
    .Y(_0626_),
    .B1(_0457_));
 sg13g2_xor2_1 _4764_ (.B(_0604_),
    .A(_0602_),
    .X(_0627_));
 sg13g2_nand2_1 _4765_ (.Y(_0628_),
    .A(_0614_),
    .B(_0627_));
 sg13g2_a22oi_1 _4766_ (.Y(_0629_),
    .B1(_0626_),
    .B2(_0628_),
    .A2(_0624_),
    .A1(net489));
 sg13g2_xnor2_1 _4767_ (.Y(_0630_),
    .A(_0247_),
    .B(_0629_));
 sg13g2_a21oi_1 _4768_ (.A1(net483),
    .A2(_0622_),
    .Y(_0631_),
    .B1(net492));
 sg13g2_o21ai_1 _4769_ (.B1(_0456_),
    .Y(_0632_),
    .A1(_0431_),
    .A2(_0627_));
 sg13g2_or2_2 _4770_ (.X(_0633_),
    .B(_0632_),
    .A(_0631_));
 sg13g2_and2_1 _4771_ (.A(_0630_),
    .B(_0633_),
    .X(_0635_));
 sg13g2_xor2_1 _4772_ (.B(_0633_),
    .A(_0630_),
    .X(_0636_));
 sg13g2_nand2b_1 _4773_ (.Y(_0637_),
    .B(_0636_),
    .A_N(_0621_));
 sg13g2_nand2_1 _4774_ (.Y(_0638_),
    .A(_0614_),
    .B(_0625_));
 sg13g2_xnor2_1 _4775_ (.Y(_0639_),
    .A(_0591_),
    .B(_0593_));
 sg13g2_a21oi_1 _4776_ (.A1(net492),
    .A2(_0639_),
    .Y(_0640_),
    .B1(_0457_));
 sg13g2_a22oi_1 _4777_ (.Y(_0641_),
    .B1(_0638_),
    .B2(_0640_),
    .A2(_0399_),
    .A1(_0358_));
 sg13g2_o21ai_1 _4778_ (.B1(_0641_),
    .Y(_0642_),
    .A1(_0439_),
    .A2(_0627_));
 sg13g2_nand2b_1 _4779_ (.Y(_0643_),
    .B(_0264_),
    .A_N(_0642_));
 sg13g2_xor2_1 _4780_ (.B(_0642_),
    .A(_0264_),
    .X(_0644_));
 sg13g2_o21ai_1 _4781_ (.B1(_0643_),
    .Y(_0646_),
    .A1(_0629_),
    .A2(_0644_));
 sg13g2_xor2_1 _4782_ (.B(_0620_),
    .A(_0619_),
    .X(_0647_));
 sg13g2_nand2_1 _4783_ (.Y(_0648_),
    .A(_0646_),
    .B(_0647_));
 sg13g2_o21ai_1 _4784_ (.B1(_0588_),
    .Y(_0649_),
    .A1(_0581_),
    .A2(_0589_));
 sg13g2_nor2b_1 _4785_ (.A(_0591_),
    .B_N(_0649_),
    .Y(_0650_));
 sg13g2_nand2_1 _4786_ (.Y(_0651_),
    .A(_0611_),
    .B(_0614_));
 sg13g2_o21ai_1 _4787_ (.B1(_0651_),
    .Y(_0652_),
    .A1(_0614_),
    .A2(_0650_));
 sg13g2_mux2_2 _4788_ (.A0(_0609_),
    .A1(_0652_),
    .S(_0439_),
    .X(_0653_));
 sg13g2_nor2_1 _4789_ (.A(_0272_),
    .B(_0653_),
    .Y(_0654_));
 sg13g2_nand2_1 _4790_ (.Y(_0655_),
    .A(net469),
    .B(_0653_));
 sg13g2_nand2b_1 _4791_ (.Y(_0657_),
    .B(_0655_),
    .A_N(_0654_));
 sg13g2_a21oi_1 _4792_ (.A1(_0615_),
    .A2(_0655_),
    .Y(_0658_),
    .B1(_0654_));
 sg13g2_xnor2_1 _4793_ (.Y(_0659_),
    .A(_0629_),
    .B(_0644_));
 sg13g2_nor2_1 _4794_ (.A(_0658_),
    .B(_0659_),
    .Y(_0660_));
 sg13g2_nand2b_1 _4795_ (.Y(_0661_),
    .B(_0277_),
    .A_N(_0642_));
 sg13g2_xnor2_1 _4796_ (.Y(_0662_),
    .A(_0615_),
    .B(_0657_));
 sg13g2_nand2_1 _4797_ (.Y(_0663_),
    .A(_0661_),
    .B(_0662_));
 sg13g2_xnor2_1 _4798_ (.Y(_0664_),
    .A(_0277_),
    .B(_0642_));
 sg13g2_nand2b_1 _4799_ (.Y(_0665_),
    .B(_0614_),
    .A_N(_0639_));
 sg13g2_xor2_1 _4800_ (.B(_0586_),
    .A(_0585_),
    .X(_0666_));
 sg13g2_a21oi_1 _4801_ (.A1(_0432_),
    .A2(_0666_),
    .Y(_0668_),
    .B1(_0457_));
 sg13g2_a22oi_1 _4802_ (.Y(_0669_),
    .B1(_0665_),
    .B2(_0668_),
    .A2(_0625_),
    .A1(net489));
 sg13g2_or2_1 _4803_ (.X(_0670_),
    .B(_0669_),
    .A(_0664_));
 sg13g2_xnor2_1 _4804_ (.Y(_0671_),
    .A(_0661_),
    .B(_0662_));
 sg13g2_o21ai_1 _4805_ (.B1(_0663_),
    .Y(_0672_),
    .A1(_0670_),
    .A2(_0671_));
 sg13g2_xor2_1 _4806_ (.B(_0659_),
    .A(_0658_),
    .X(_0673_));
 sg13g2_a21oi_1 _4807_ (.A1(_0672_),
    .A2(_0673_),
    .Y(_0674_),
    .B1(_0660_));
 sg13g2_xnor2_1 _4808_ (.Y(_0675_),
    .A(_0646_),
    .B(_0647_));
 sg13g2_o21ai_1 _4809_ (.B1(_0648_),
    .Y(_0676_),
    .A1(_0674_),
    .A2(_0675_));
 sg13g2_xnor2_1 _4810_ (.Y(_0677_),
    .A(_0621_),
    .B(_0636_));
 sg13g2_nand2_1 _4811_ (.Y(_0679_),
    .A(_0676_),
    .B(_0677_));
 sg13g2_a21o_1 _4812_ (.A2(_0629_),
    .A1(_0248_),
    .B1(_0635_),
    .X(_0680_));
 sg13g2_a21oi_1 _4813_ (.A1(_0617_),
    .A2(_0618_),
    .Y(_0681_),
    .B1(_0232_));
 sg13g2_xnor2_1 _4814_ (.Y(_0682_),
    .A(_0233_),
    .B(_0619_));
 sg13g2_xnor2_1 _4815_ (.Y(_0683_),
    .A(_0680_),
    .B(_0682_));
 sg13g2_a21oi_1 _4816_ (.A1(_0637_),
    .A2(_0679_),
    .Y(_0684_),
    .B1(_0683_));
 sg13g2_nand3_1 _4817_ (.B(_0679_),
    .C(_0683_),
    .A(_0637_),
    .Y(_0685_));
 sg13g2_nand2b_1 _4818_ (.Y(_0686_),
    .B(_0685_),
    .A_N(_0684_));
 sg13g2_xnor2_1 _4819_ (.Y(_0687_),
    .A(_0676_),
    .B(_0677_));
 sg13g2_xor2_1 _4820_ (.B(_0675_),
    .A(_0674_),
    .X(_0688_));
 sg13g2_inv_1 _4821_ (.Y(_0690_),
    .A(_0688_));
 sg13g2_xnor2_1 _4822_ (.Y(_0691_),
    .A(_0672_),
    .B(_0673_));
 sg13g2_xnor2_1 _4823_ (.Y(_0692_),
    .A(_0664_),
    .B(_0669_));
 sg13g2_xnor2_1 _4824_ (.Y(_0693_),
    .A(_0670_),
    .B(_0671_));
 sg13g2_nand4_1 _4825_ (.B(_0691_),
    .C(_0692_),
    .A(_0687_),
    .Y(_0694_),
    .D(_0693_));
 sg13g2_nor2_1 _4826_ (.A(_0688_),
    .B(_0694_),
    .Y(_0695_));
 sg13g2_a21oi_1 _4827_ (.A1(_0680_),
    .A2(_0682_),
    .Y(_0696_),
    .B1(_0684_));
 sg13g2_xor2_1 _4828_ (.B(_0633_),
    .A(_0288_),
    .X(_0697_));
 sg13g2_xnor2_1 _4829_ (.Y(_0698_),
    .A(_0681_),
    .B(_0697_));
 sg13g2_nor4_1 _4830_ (.A(_0687_),
    .B(_0690_),
    .C(_0691_),
    .D(_0693_),
    .Y(_0699_));
 sg13g2_xnor2_1 _4831_ (.Y(_0701_),
    .A(_0696_),
    .B(_0698_));
 sg13g2_mux2_1 _4832_ (.A0(_0695_),
    .A1(_0699_),
    .S(_0686_),
    .X(_0702_));
 sg13g2_nand4_1 _4833_ (.B(_0311_),
    .C(_0701_),
    .A(_0310_),
    .Y(_0703_),
    .D(_0702_));
 sg13g2_a21oi_1 _4834_ (.A1(_2641_),
    .A2(_0340_),
    .Y(_0704_),
    .B1(_2651_));
 sg13g2_nand2_1 _4835_ (.Y(_0705_),
    .A(_0332_),
    .B(_0704_));
 sg13g2_a21oi_2 _4836_ (.B1(_2610_),
    .Y(_0706_),
    .A2(_2617_),
    .A1(net601));
 sg13g2_o21ai_1 _4837_ (.B1(_0706_),
    .Y(_0707_),
    .A1(_2623_),
    .A2(_2625_));
 sg13g2_and2_1 _4838_ (.A(_2642_),
    .B(_0707_),
    .X(_0708_));
 sg13g2_a22oi_1 _4839_ (.Y(_0709_),
    .B1(_0707_),
    .B2(_2642_),
    .A2(_0336_),
    .A1(_0335_));
 sg13g2_a21o_1 _4840_ (.A2(_0709_),
    .A1(_0333_),
    .B1(net546),
    .X(_0710_));
 sg13g2_a21oi_2 _4841_ (.B1(_0329_),
    .Y(_0712_),
    .A2(_0710_),
    .A1(_0705_));
 sg13g2_a21o_1 _4842_ (.A2(_0710_),
    .A1(_0705_),
    .B1(_0329_),
    .X(_0713_));
 sg13g2_xnor2_1 _4843_ (.Y(_0714_),
    .A(net529),
    .B(_0712_));
 sg13g2_a21oi_2 _4844_ (.B1(_0322_),
    .Y(_0715_),
    .A2(_0713_),
    .A1(_0323_));
 sg13g2_o21ai_1 _4845_ (.B1(_0321_),
    .Y(_0716_),
    .A1(net529),
    .A2(_0712_));
 sg13g2_nor3_2 _4846_ (.A(_0321_),
    .B(net529),
    .C(_0712_),
    .Y(_0717_));
 sg13g2_nand3_1 _4847_ (.B(_0323_),
    .C(_0713_),
    .A(_0322_),
    .Y(_0718_));
 sg13g2_nor2_1 _4848_ (.A(_0715_),
    .B(_0717_),
    .Y(_0719_));
 sg13g2_nand2_1 _4849_ (.Y(_0720_),
    .A(_0714_),
    .B(_0719_));
 sg13g2_nand3_1 _4850_ (.B(_0705_),
    .C(_0710_),
    .A(_0329_),
    .Y(_0721_));
 sg13g2_and2_1 _4851_ (.A(_0713_),
    .B(_0721_),
    .X(_0723_));
 sg13g2_xnor2_1 _4852_ (.Y(_0724_),
    .A(_0332_),
    .B(_0704_));
 sg13g2_xnor2_1 _4853_ (.Y(_0725_),
    .A(_0332_),
    .B(_0709_));
 sg13g2_a22oi_1 _4854_ (.Y(_0726_),
    .B1(_0725_),
    .B2(_3279_),
    .A2(_0724_),
    .A1(net546));
 sg13g2_xnor2_1 _4855_ (.Y(_0727_),
    .A(_3202_),
    .B(_2622_));
 sg13g2_xnor2_1 _4856_ (.Y(_0728_),
    .A(_2614_),
    .B(_0727_));
 sg13g2_xnor2_1 _4857_ (.Y(_0729_),
    .A(_2615_),
    .B(_0727_));
 sg13g2_nand2b_1 _4858_ (.Y(_0730_),
    .B(_0706_),
    .A_N(_0727_));
 sg13g2_xor2_1 _4859_ (.B(_0727_),
    .A(_0706_),
    .X(_0731_));
 sg13g2_mux2_1 _4860_ (.A0(_0728_),
    .A1(_0731_),
    .S(net538),
    .X(_0732_));
 sg13g2_nor2_1 _4861_ (.A(net546),
    .B(_2619_),
    .Y(_0734_));
 sg13g2_xnor2_1 _4862_ (.Y(_0735_),
    .A(net538),
    .B(_2619_));
 sg13g2_nor2_1 _4863_ (.A(net607),
    .B(_0735_),
    .Y(_0736_));
 sg13g2_mux2_1 _4864_ (.A0(_2614_),
    .A1(net604),
    .S(_0734_),
    .X(_0737_));
 sg13g2_and2_1 _4865_ (.A(_0736_),
    .B(_0737_),
    .X(_0738_));
 sg13g2_and2_1 _4866_ (.A(_0732_),
    .B(_0738_),
    .X(_0739_));
 sg13g2_mux2_1 _4867_ (.A0(_0340_),
    .A1(_0730_),
    .S(net538),
    .X(_0740_));
 sg13g2_xnor2_1 _4868_ (.Y(_0741_),
    .A(_2641_),
    .B(_0740_));
 sg13g2_and2_1 _4869_ (.A(_0739_),
    .B(_0741_),
    .X(_0742_));
 sg13g2_a21o_1 _4870_ (.A2(_0361_),
    .A1(_0340_),
    .B1(net539),
    .X(_0743_));
 sg13g2_o21ai_1 _4871_ (.B1(_0743_),
    .Y(_0745_),
    .A1(net548),
    .A2(_0708_));
 sg13g2_xnor2_1 _4872_ (.Y(_0746_),
    .A(_2651_),
    .B(_0745_));
 sg13g2_nand3_1 _4873_ (.B(_0741_),
    .C(_0746_),
    .A(_0739_),
    .Y(_0747_));
 sg13g2_and4_1 _4874_ (.A(_0726_),
    .B(_0739_),
    .C(_0741_),
    .D(_0746_),
    .X(_0748_));
 sg13g2_nand2_1 _4875_ (.Y(_0749_),
    .A(_0723_),
    .B(_0748_));
 sg13g2_a21o_1 _4876_ (.A2(_0749_),
    .A1(_0719_),
    .B1(_0714_),
    .X(_0750_));
 sg13g2_nand2_2 _4877_ (.Y(_0751_),
    .A(_0720_),
    .B(_0750_));
 sg13g2_or3_1 _4878_ (.A(_0715_),
    .B(_0717_),
    .C(_0748_),
    .X(_0752_));
 sg13g2_xor2_1 _4879_ (.B(_0752_),
    .A(_0723_),
    .X(_0753_));
 sg13g2_nand3_1 _4880_ (.B(_0719_),
    .C(_0749_),
    .A(_0714_),
    .Y(_0754_));
 sg13g2_and3_1 _4881_ (.X(_0756_),
    .A(_0750_),
    .B(_0753_),
    .C(_0754_));
 sg13g2_nor2_1 _4882_ (.A(_0751_),
    .B(_0756_),
    .Y(_0757_));
 sg13g2_inv_2 _4883_ (.Y(_0758_),
    .A(net497));
 sg13g2_nand3_1 _4884_ (.B(_0718_),
    .C(_0747_),
    .A(_0716_),
    .Y(_0759_));
 sg13g2_xor2_1 _4885_ (.B(_0759_),
    .A(_0726_),
    .X(_0760_));
 sg13g2_nor2_2 _4886_ (.A(_0753_),
    .B(_0760_),
    .Y(_0761_));
 sg13g2_nor2b_2 _4887_ (.A(_0751_),
    .B_N(_0761_),
    .Y(_0762_));
 sg13g2_nand2b_2 _4888_ (.Y(_0763_),
    .B(_0761_),
    .A_N(_0751_));
 sg13g2_nor2_1 _4889_ (.A(_0720_),
    .B(_0749_),
    .Y(_0764_));
 sg13g2_nor2_1 _4890_ (.A(_0756_),
    .B(_0764_),
    .Y(_0765_));
 sg13g2_nor3_1 _4891_ (.A(_0715_),
    .B(_0717_),
    .C(_0736_),
    .Y(_0767_));
 sg13g2_xor2_1 _4892_ (.B(_0767_),
    .A(_0737_),
    .X(_0768_));
 sg13g2_inv_1 _4893_ (.Y(_0769_),
    .A(_0768_));
 sg13g2_nand3_1 _4894_ (.B(_0716_),
    .C(_0718_),
    .A(net607),
    .Y(_0770_));
 sg13g2_xnor2_1 _4895_ (.Y(_0771_),
    .A(_0735_),
    .B(_0770_));
 sg13g2_nor3_1 _4896_ (.A(_0715_),
    .B(_0717_),
    .C(_0738_),
    .Y(_0772_));
 sg13g2_xnor2_1 _4897_ (.Y(_0773_),
    .A(_0732_),
    .B(_0772_));
 sg13g2_inv_1 _4898_ (.Y(_0774_),
    .A(_0773_));
 sg13g2_a21o_1 _4899_ (.A2(_0771_),
    .A1(_0768_),
    .B1(_0773_),
    .X(_0775_));
 sg13g2_nor3_1 _4900_ (.A(_0715_),
    .B(_0717_),
    .C(_0739_),
    .Y(_0776_));
 sg13g2_xnor2_1 _4901_ (.Y(_0778_),
    .A(_0741_),
    .B(_0776_));
 sg13g2_inv_1 _4902_ (.Y(_0779_),
    .A(_0778_));
 sg13g2_nor3_1 _4903_ (.A(_0715_),
    .B(_0717_),
    .C(_0742_),
    .Y(_0780_));
 sg13g2_xnor2_1 _4904_ (.Y(_0781_),
    .A(_0746_),
    .B(_0780_));
 sg13g2_a21oi_1 _4905_ (.A1(_0775_),
    .A2(_0779_),
    .Y(_0782_),
    .B1(_0781_));
 sg13g2_o21ai_1 _4906_ (.B1(net496),
    .Y(_0783_),
    .A1(_0763_),
    .A2(_0782_));
 sg13g2_mux2_1 _4907_ (.A0(_0753_),
    .A1(_0760_),
    .S(_0783_),
    .X(_0784_));
 sg13g2_a21o_2 _4908_ (.A2(_0781_),
    .A1(net498),
    .B1(_0784_),
    .X(_0785_));
 sg13g2_inv_1 _4909_ (.Y(_0786_),
    .A(net481));
 sg13g2_nor2_1 _4910_ (.A(_0778_),
    .B(_0781_),
    .Y(_0787_));
 sg13g2_o21ai_1 _4911_ (.B1(_0787_),
    .Y(_0789_),
    .A1(_0769_),
    .A2(_0773_));
 sg13g2_a21o_1 _4912_ (.A2(_0789_),
    .A1(_0761_),
    .B1(_0751_),
    .X(_0790_));
 sg13g2_xnor2_1 _4913_ (.Y(_0791_),
    .A(_0783_),
    .B(_0790_));
 sg13g2_a21oi_1 _4914_ (.A1(_0761_),
    .A2(_0787_),
    .Y(_0792_),
    .B1(_0751_));
 sg13g2_inv_1 _4915_ (.Y(_0793_),
    .A(_0792_));
 sg13g2_a21oi_1 _4916_ (.A1(_0790_),
    .A2(_0793_),
    .Y(_0794_),
    .B1(_0756_));
 sg13g2_mux2_1 _4917_ (.A0(_0774_),
    .A1(_0768_),
    .S(_0783_),
    .X(_0795_));
 sg13g2_nor3_1 _4918_ (.A(_0791_),
    .B(_0794_),
    .C(_0795_),
    .Y(_0796_));
 sg13g2_a21o_2 _4919_ (.A2(_0771_),
    .A1(net497),
    .B1(_0796_),
    .X(_0797_));
 sg13g2_nand2_2 _4920_ (.Y(_0798_),
    .A(_0763_),
    .B(_0797_));
 sg13g2_nand2_1 _4921_ (.Y(_0800_),
    .A(net497),
    .B(_0773_));
 sg13g2_nor2_2 _4922_ (.A(net497),
    .B(_0764_),
    .Y(_0801_));
 sg13g2_or2_2 _4923_ (.X(_0802_),
    .B(_0764_),
    .A(net497));
 sg13g2_mux2_1 _4924_ (.A0(_0781_),
    .A1(_0778_),
    .S(_0783_),
    .X(_0803_));
 sg13g2_nor3_1 _4925_ (.A(_0791_),
    .B(_0794_),
    .C(_0803_),
    .Y(_0804_));
 sg13g2_o21ai_1 _4926_ (.B1(_0800_),
    .Y(_0805_),
    .A1(_0802_),
    .A2(_0804_));
 sg13g2_nor2_1 _4927_ (.A(_0778_),
    .B(_0783_),
    .Y(_0806_));
 sg13g2_and2_1 _4928_ (.A(_0774_),
    .B(_0783_),
    .X(_0807_));
 sg13g2_or4_2 _4929_ (.A(_0791_),
    .B(_0794_),
    .C(_0806_),
    .D(_0807_),
    .X(_0808_));
 sg13g2_nand2_2 _4930_ (.Y(_0809_),
    .A(net498),
    .B(_0769_));
 sg13g2_nand2_2 _4931_ (.Y(_0811_),
    .A(_0808_),
    .B(_0809_));
 sg13g2_nand2_1 _4932_ (.Y(_0812_),
    .A(net498),
    .B(_0778_));
 sg13g2_mux2_1 _4933_ (.A0(_0760_),
    .A1(_0781_),
    .S(_0783_),
    .X(_0813_));
 sg13g2_o21ai_1 _4934_ (.B1(_0801_),
    .Y(_0814_),
    .A1(_0791_),
    .A2(_0813_));
 sg13g2_nand2_2 _4935_ (.Y(_0815_),
    .A(_0812_),
    .B(_0814_));
 sg13g2_a22oi_1 _4936_ (.Y(_0816_),
    .B1(_0812_),
    .B2(_0814_),
    .A2(_0809_),
    .A1(_0808_));
 sg13g2_and2_1 _4937_ (.A(net477),
    .B(_0815_),
    .X(_0817_));
 sg13g2_nand2_1 _4938_ (.Y(_0818_),
    .A(_0805_),
    .B(_0816_));
 sg13g2_nand2_2 _4939_ (.Y(_0819_),
    .A(_0785_),
    .B(_0797_));
 sg13g2_xnor2_1 _4940_ (.Y(_0820_),
    .A(_0805_),
    .B(_0816_));
 sg13g2_o21ai_1 _4941_ (.B1(_0818_),
    .Y(_0822_),
    .A1(_0819_),
    .A2(_0820_));
 sg13g2_nor2_1 _4942_ (.A(_0798_),
    .B(_0822_),
    .Y(_0823_));
 sg13g2_nand2_1 _4943_ (.Y(_0824_),
    .A(net481),
    .B(_0811_));
 sg13g2_nand2_1 _4944_ (.Y(_0825_),
    .A(net481),
    .B(net477));
 sg13g2_nand3_1 _4945_ (.B(net477),
    .C(_0816_),
    .A(_0785_),
    .Y(_0826_));
 sg13g2_nor2b_1 _4946_ (.A(_0817_),
    .B_N(_0824_),
    .Y(_0827_));
 sg13g2_xor2_1 _4947_ (.B(_0824_),
    .A(_0817_),
    .X(_0828_));
 sg13g2_a21oi_1 _4948_ (.A1(_0798_),
    .A2(_0828_),
    .Y(_0829_),
    .B1(_0823_));
 sg13g2_nand2_1 _4949_ (.Y(_0830_),
    .A(net481),
    .B(_0817_));
 sg13g2_xor2_1 _4950_ (.B(_0825_),
    .A(_0815_),
    .X(_0831_));
 sg13g2_a21oi_2 _4951_ (.B1(_0762_),
    .Y(_0833_),
    .A2(_0809_),
    .A1(_0808_));
 sg13g2_nand2_1 _4952_ (.Y(_0834_),
    .A(_0763_),
    .B(net477));
 sg13g2_nand3_1 _4953_ (.B(net477),
    .C(_0833_),
    .A(net481),
    .Y(_0835_));
 sg13g2_xnor2_1 _4954_ (.Y(_0836_),
    .A(_0825_),
    .B(_0833_));
 sg13g2_o21ai_1 _4955_ (.B1(_0826_),
    .Y(_0837_),
    .A1(_0798_),
    .A2(_0827_));
 sg13g2_nand2_1 _4956_ (.Y(_0838_),
    .A(_0836_),
    .B(_0837_));
 sg13g2_xnor2_1 _4957_ (.Y(_0839_),
    .A(_0836_),
    .B(_0837_));
 sg13g2_xor2_1 _4958_ (.B(_0839_),
    .A(_0831_),
    .X(_0840_));
 sg13g2_nand2_1 _4959_ (.Y(_0841_),
    .A(_0829_),
    .B(_0840_));
 sg13g2_xnor2_1 _4960_ (.Y(_0842_),
    .A(_0829_),
    .B(_0840_));
 sg13g2_o21ai_1 _4961_ (.B1(_0841_),
    .Y(_0844_),
    .A1(_0826_),
    .A2(_0842_));
 sg13g2_nor2b_1 _4962_ (.A(_0834_),
    .B_N(_0824_),
    .Y(_0845_));
 sg13g2_o21ai_1 _4963_ (.B1(_0838_),
    .Y(_0846_),
    .A1(_0831_),
    .A2(_0839_));
 sg13g2_nand2_1 _4964_ (.Y(_0847_),
    .A(_0845_),
    .B(_0846_));
 sg13g2_xor2_1 _4965_ (.B(_0846_),
    .A(_0845_),
    .X(_0848_));
 sg13g2_nand2b_1 _4966_ (.Y(_0849_),
    .B(_0848_),
    .A_N(_0830_));
 sg13g2_xnor2_1 _4967_ (.Y(_0850_),
    .A(_0830_),
    .B(_0848_));
 sg13g2_nand2_1 _4968_ (.Y(_0851_),
    .A(_0844_),
    .B(_0850_));
 sg13g2_xnor2_1 _4969_ (.Y(_0852_),
    .A(_0844_),
    .B(_0850_));
 sg13g2_o21ai_1 _4970_ (.B1(_0851_),
    .Y(_0853_),
    .A1(_0834_),
    .A2(_0852_));
 sg13g2_nand2_1 _4971_ (.Y(_0855_),
    .A(_0763_),
    .B(_0815_));
 sg13g2_o21ai_1 _4972_ (.B1(_0855_),
    .Y(_0856_),
    .A1(_0786_),
    .A2(_0815_));
 sg13g2_nand2b_1 _4973_ (.Y(_0857_),
    .B(_0835_),
    .A_N(_0815_));
 sg13g2_nand2_1 _4974_ (.Y(_0858_),
    .A(_0835_),
    .B(_0856_));
 sg13g2_a21o_1 _4975_ (.A2(_0849_),
    .A1(_0847_),
    .B1(_0858_),
    .X(_0859_));
 sg13g2_nand3_1 _4976_ (.B(_0849_),
    .C(_0858_),
    .A(_0847_),
    .Y(_0860_));
 sg13g2_nand2_1 _4977_ (.Y(_0861_),
    .A(_0859_),
    .B(_0860_));
 sg13g2_xor2_1 _4978_ (.B(_0861_),
    .A(_0855_),
    .X(_0862_));
 sg13g2_nand2_1 _4979_ (.Y(_0863_),
    .A(_0853_),
    .B(_0862_));
 sg13g2_nand2_2 _4980_ (.Y(_0864_),
    .A(net477),
    .B(_0811_));
 sg13g2_xnor2_1 _4981_ (.Y(_0866_),
    .A(_0819_),
    .B(_0820_));
 sg13g2_nor2_1 _4982_ (.A(_0864_),
    .B(_0866_),
    .Y(_0867_));
 sg13g2_xor2_1 _4983_ (.B(_0866_),
    .A(_0864_),
    .X(_0868_));
 sg13g2_nor2_2 _4984_ (.A(_3235_),
    .B(_0758_),
    .Y(_0869_));
 sg13g2_nand2_2 _4985_ (.Y(_0870_),
    .A(_0010_),
    .B(net498));
 sg13g2_nor2_1 _4986_ (.A(_0762_),
    .B(_0869_),
    .Y(_0871_));
 sg13g2_inv_1 _4987_ (.Y(_0872_),
    .A(_0871_));
 sg13g2_nand2_2 _4988_ (.Y(_0873_),
    .A(_0815_),
    .B(_0870_));
 sg13g2_nand2_1 _4989_ (.Y(_0874_),
    .A(_0816_),
    .B(_0871_));
 sg13g2_xnor2_1 _4990_ (.Y(_0875_),
    .A(_0816_),
    .B(_0871_));
 sg13g2_xor2_1 _4991_ (.B(_0875_),
    .A(_0819_),
    .X(_0877_));
 sg13g2_a21oi_1 _4992_ (.A1(_0868_),
    .A2(_0877_),
    .Y(_0878_),
    .B1(_0867_));
 sg13g2_xnor2_1 _4993_ (.Y(_0879_),
    .A(_0798_),
    .B(_0822_));
 sg13g2_nand2b_1 _4994_ (.Y(_0880_),
    .B(_0879_),
    .A_N(_0878_));
 sg13g2_o21ai_1 _4995_ (.B1(_0874_),
    .Y(_0881_),
    .A1(_0819_),
    .A2(_0875_));
 sg13g2_xor2_1 _4996_ (.B(_0879_),
    .A(_0878_),
    .X(_0882_));
 sg13g2_nand2b_1 _4997_ (.Y(_0883_),
    .B(_0881_),
    .A_N(_0882_));
 sg13g2_and2_1 _4998_ (.A(_0880_),
    .B(_0883_),
    .X(_0884_));
 sg13g2_xor2_1 _4999_ (.B(_0842_),
    .A(_0826_),
    .X(_0885_));
 sg13g2_nor2b_1 _5000_ (.A(_0884_),
    .B_N(_0885_),
    .Y(_0886_));
 sg13g2_xnor2_1 _5001_ (.Y(_0888_),
    .A(_0884_),
    .B(_0885_));
 sg13g2_a21oi_1 _5002_ (.A1(_0833_),
    .A2(_0888_),
    .Y(_0889_),
    .B1(_0886_));
 sg13g2_xor2_1 _5003_ (.B(_0852_),
    .A(_0834_),
    .X(_0890_));
 sg13g2_nor2b_1 _5004_ (.A(_0889_),
    .B_N(_0890_),
    .Y(_0891_));
 sg13g2_nand2_1 _5005_ (.Y(_0892_),
    .A(_0797_),
    .B(_0815_));
 sg13g2_xor2_1 _5006_ (.B(_0877_),
    .A(_0868_),
    .X(_0893_));
 sg13g2_nand2b_1 _5007_ (.Y(_0894_),
    .B(_0893_),
    .A_N(_0892_));
 sg13g2_nand2_1 _5008_ (.Y(_0895_),
    .A(_0785_),
    .B(_0870_));
 sg13g2_xor2_1 _5009_ (.B(_0893_),
    .A(_0892_),
    .X(_0896_));
 sg13g2_o21ai_1 _5010_ (.B1(_0894_),
    .Y(_0897_),
    .A1(_0895_),
    .A2(_0896_));
 sg13g2_xor2_1 _5011_ (.B(_0882_),
    .A(_0881_),
    .X(_0899_));
 sg13g2_inv_1 _5012_ (.Y(_0900_),
    .A(_0899_));
 sg13g2_xor2_1 _5013_ (.B(_0899_),
    .A(_0897_),
    .X(_0901_));
 sg13g2_nor2_1 _5014_ (.A(_0798_),
    .B(_0901_),
    .Y(_0902_));
 sg13g2_a21oi_1 _5015_ (.A1(_0897_),
    .A2(_0900_),
    .Y(_0903_),
    .B1(_0902_));
 sg13g2_xnor2_1 _5016_ (.Y(_0904_),
    .A(_0833_),
    .B(_0888_));
 sg13g2_nor2_1 _5017_ (.A(_0903_),
    .B(_0904_),
    .Y(_0905_));
 sg13g2_xor2_1 _5018_ (.B(_0811_),
    .A(net477),
    .X(_0906_));
 sg13g2_nand2_1 _5019_ (.Y(_0907_),
    .A(_0797_),
    .B(_0906_));
 sg13g2_nand3_1 _5020_ (.B(net477),
    .C(_0811_),
    .A(_0797_),
    .Y(_0908_));
 sg13g2_o21ai_1 _5021_ (.B1(_0908_),
    .Y(_0910_),
    .A1(_0873_),
    .A2(_0907_));
 sg13g2_xor2_1 _5022_ (.B(_0896_),
    .A(_0895_),
    .X(_0911_));
 sg13g2_nand2_1 _5023_ (.Y(_0912_),
    .A(_0910_),
    .B(_0911_));
 sg13g2_xnor2_1 _5024_ (.Y(_0913_),
    .A(_0910_),
    .B(_0911_));
 sg13g2_o21ai_1 _5025_ (.B1(_0912_),
    .Y(_0914_),
    .A1(_0872_),
    .A2(_0913_));
 sg13g2_xnor2_1 _5026_ (.Y(_0915_),
    .A(_0798_),
    .B(_0901_));
 sg13g2_nor2b_1 _5027_ (.A(_0915_),
    .B_N(_0914_),
    .Y(_0916_));
 sg13g2_xnor2_1 _5028_ (.Y(_0917_),
    .A(_0873_),
    .B(_0907_));
 sg13g2_nor3_1 _5029_ (.A(_0864_),
    .B(_0869_),
    .C(_0873_),
    .Y(_0918_));
 sg13g2_xnor2_1 _5030_ (.Y(_0919_),
    .A(_0872_),
    .B(_0913_));
 sg13g2_nor4_2 _5031_ (.A(_0864_),
    .B(_0869_),
    .C(_0873_),
    .Y(_0921_),
    .D(_0919_));
 sg13g2_xnor2_1 _5032_ (.Y(_0922_),
    .A(_0914_),
    .B(_0915_));
 sg13g2_a21o_1 _5033_ (.A2(_0922_),
    .A1(_0921_),
    .B1(_0916_),
    .X(_0923_));
 sg13g2_xor2_1 _5034_ (.B(_0904_),
    .A(_0903_),
    .X(_0924_));
 sg13g2_a21o_1 _5035_ (.A2(_0924_),
    .A1(_0923_),
    .B1(_0905_),
    .X(_0925_));
 sg13g2_xnor2_1 _5036_ (.Y(_0926_),
    .A(_0889_),
    .B(_0890_));
 sg13g2_a21oi_1 _5037_ (.A1(_0925_),
    .A2(_0926_),
    .Y(_0927_),
    .B1(_0891_));
 sg13g2_xnor2_1 _5038_ (.Y(_0928_),
    .A(_0853_),
    .B(_0862_));
 sg13g2_o21ai_1 _5039_ (.B1(_0863_),
    .Y(_0929_),
    .A1(_0927_),
    .A2(_0928_));
 sg13g2_o21ai_1 _5040_ (.B1(_0859_),
    .Y(_0930_),
    .A1(_0855_),
    .A2(_0861_));
 sg13g2_nand3_1 _5041_ (.B(_0817_),
    .C(_0833_),
    .A(net481),
    .Y(_0932_));
 sg13g2_nand3_1 _5042_ (.B(_0857_),
    .C(_0932_),
    .A(net481),
    .Y(_0933_));
 sg13g2_nor2b_1 _5043_ (.A(_0933_),
    .B_N(_0930_),
    .Y(_0934_));
 sg13g2_xor2_1 _5044_ (.B(_0933_),
    .A(_0930_),
    .X(_0935_));
 sg13g2_inv_1 _5045_ (.Y(_0936_),
    .A(_0935_));
 sg13g2_a21oi_1 _5046_ (.A1(_0929_),
    .A2(_0936_),
    .Y(_0937_),
    .B1(_0934_));
 sg13g2_a21oi_1 _5047_ (.A1(_0786_),
    .A2(_0937_),
    .Y(_0938_),
    .B1(_0762_));
 sg13g2_xnor2_1 _5048_ (.Y(_0939_),
    .A(_0929_),
    .B(_0936_));
 sg13g2_xor2_1 _5049_ (.B(_0926_),
    .A(_0925_),
    .X(_0940_));
 sg13g2_a21oi_1 _5050_ (.A1(net494),
    .A2(_0940_),
    .Y(_0941_),
    .B1(_0802_));
 sg13g2_o21ai_1 _5051_ (.B1(_0941_),
    .Y(_0943_),
    .A1(net494),
    .A2(_0939_));
 sg13g2_o21ai_1 _5052_ (.B1(_0943_),
    .Y(_0944_),
    .A1(_0758_),
    .A2(_0938_));
 sg13g2_a21oi_1 _5053_ (.A1(net494),
    .A2(_0939_),
    .Y(_0945_),
    .B1(_0802_));
 sg13g2_o21ai_1 _5054_ (.B1(_0945_),
    .Y(_0946_),
    .A1(net494),
    .A2(_0938_));
 sg13g2_xnor2_1 _5055_ (.Y(_0947_),
    .A(_0248_),
    .B(_0944_));
 sg13g2_nand2_1 _5056_ (.Y(_0948_),
    .A(_0946_),
    .B(_0947_));
 sg13g2_o21ai_1 _5057_ (.B1(_0948_),
    .Y(_0949_),
    .A1(_0247_),
    .A2(_0944_));
 sg13g2_o21ai_1 _5058_ (.B1(_0932_),
    .Y(_0950_),
    .A1(_0762_),
    .A2(net481));
 sg13g2_xnor2_1 _5059_ (.Y(_0951_),
    .A(_0937_),
    .B(_0950_));
 sg13g2_xor2_1 _5060_ (.B(_0928_),
    .A(_0927_),
    .X(_0952_));
 sg13g2_nand2b_1 _5061_ (.Y(_0954_),
    .B(net494),
    .A_N(_0952_));
 sg13g2_o21ai_1 _5062_ (.B1(_0801_),
    .Y(_0955_),
    .A1(net494),
    .A2(_0951_));
 sg13g2_nand2b_2 _5063_ (.Y(_0956_),
    .B(_0954_),
    .A_N(_0955_));
 sg13g2_nand2_1 _5064_ (.Y(_0957_),
    .A(_0233_),
    .B(_0956_));
 sg13g2_xnor2_1 _5065_ (.Y(_0958_),
    .A(_0233_),
    .B(_0956_));
 sg13g2_nand2_1 _5066_ (.Y(_0959_),
    .A(_0949_),
    .B(_0958_));
 sg13g2_or2_1 _5067_ (.X(_0960_),
    .B(_0952_),
    .A(net494));
 sg13g2_xnor2_1 _5068_ (.Y(_0961_),
    .A(_0923_),
    .B(_0924_));
 sg13g2_inv_1 _5069_ (.Y(_0962_),
    .A(_0961_));
 sg13g2_a21oi_1 _5070_ (.A1(net495),
    .A2(_0961_),
    .Y(_0963_),
    .B1(_0802_));
 sg13g2_a22oi_1 _5071_ (.Y(_0965_),
    .B1(_0960_),
    .B2(_0963_),
    .A2(_0951_),
    .A1(net497));
 sg13g2_inv_1 _5072_ (.Y(_0966_),
    .A(_0965_));
 sg13g2_nor2_1 _5073_ (.A(_0256_),
    .B(_0965_),
    .Y(_0967_));
 sg13g2_xnor2_1 _5074_ (.Y(_0968_),
    .A(_0255_),
    .B(_0965_));
 sg13g2_a21oi_1 _5075_ (.A1(_0956_),
    .A2(_0968_),
    .Y(_0969_),
    .B1(_0967_));
 sg13g2_xnor2_1 _5076_ (.Y(_0970_),
    .A(_0946_),
    .B(_0947_));
 sg13g2_nor2_1 _5077_ (.A(_0969_),
    .B(_0970_),
    .Y(_0971_));
 sg13g2_xnor2_1 _5078_ (.Y(_0972_),
    .A(_0921_),
    .B(_0922_));
 sg13g2_a21oi_1 _5079_ (.A1(net495),
    .A2(_0972_),
    .Y(_0973_),
    .B1(_0802_));
 sg13g2_o21ai_1 _5080_ (.B1(_0973_),
    .Y(_0974_),
    .A1(net494),
    .A2(_0940_));
 sg13g2_o21ai_1 _5081_ (.B1(_0974_),
    .Y(_0976_),
    .A1(_0758_),
    .A2(_0939_));
 sg13g2_and2_1 _5082_ (.A(_0264_),
    .B(_0976_),
    .X(_0977_));
 sg13g2_xor2_1 _5083_ (.B(_0976_),
    .A(_0264_),
    .X(_0978_));
 sg13g2_a21oi_1 _5084_ (.A1(_0944_),
    .A2(_0978_),
    .Y(_0979_),
    .B1(_0977_));
 sg13g2_xnor2_1 _5085_ (.Y(_0980_),
    .A(_0956_),
    .B(_0968_));
 sg13g2_or2_1 _5086_ (.X(_0981_),
    .B(_0980_),
    .A(_0979_));
 sg13g2_xnor2_1 _5087_ (.Y(_0982_),
    .A(_0918_),
    .B(_0919_));
 sg13g2_mux2_1 _5088_ (.A0(_0962_),
    .A1(_0982_),
    .S(net495),
    .X(_0983_));
 sg13g2_a22oi_1 _5089_ (.Y(_0984_),
    .B1(_0983_),
    .B2(_0801_),
    .A2(_0952_),
    .A1(net497));
 sg13g2_nor2_1 _5090_ (.A(net469),
    .B(_0984_),
    .Y(_0985_));
 sg13g2_nand2_1 _5091_ (.Y(_0987_),
    .A(net469),
    .B(_0984_));
 sg13g2_nand2b_1 _5092_ (.Y(_0988_),
    .B(_0987_),
    .A_N(_0985_));
 sg13g2_a21oi_2 _5093_ (.B1(_0985_),
    .Y(_0989_),
    .A2(_0987_),
    .A1(_0965_));
 sg13g2_xnor2_1 _5094_ (.Y(_0990_),
    .A(_0944_),
    .B(_0978_));
 sg13g2_nor2_1 _5095_ (.A(_0989_),
    .B(_0990_),
    .Y(_0991_));
 sg13g2_nand2_1 _5096_ (.Y(_0992_),
    .A(_0277_),
    .B(_0976_));
 sg13g2_xnor2_1 _5097_ (.Y(_0993_),
    .A(_0965_),
    .B(_0988_));
 sg13g2_nand2_1 _5098_ (.Y(_0994_),
    .A(_0992_),
    .B(_0993_));
 sg13g2_xnor2_1 _5099_ (.Y(_0995_),
    .A(_0277_),
    .B(_0976_));
 sg13g2_o21ai_1 _5100_ (.B1(_0917_),
    .Y(_0996_),
    .A1(_0864_),
    .A2(_0869_));
 sg13g2_nand2b_1 _5101_ (.Y(_0998_),
    .B(_0996_),
    .A_N(_0918_));
 sg13g2_mux2_1 _5102_ (.A0(_0972_),
    .A1(_0998_),
    .S(net495),
    .X(_0999_));
 sg13g2_nand2_1 _5103_ (.Y(_1000_),
    .A(net497),
    .B(_0940_));
 sg13g2_o21ai_1 _5104_ (.B1(_1000_),
    .Y(_1001_),
    .A1(_0802_),
    .A2(_0999_));
 sg13g2_nand2_1 _5105_ (.Y(_1002_),
    .A(_0995_),
    .B(_1001_));
 sg13g2_xnor2_1 _5106_ (.Y(_1003_),
    .A(_0992_),
    .B(_0993_));
 sg13g2_o21ai_1 _5107_ (.B1(_0994_),
    .Y(_1004_),
    .A1(_1002_),
    .A2(_1003_));
 sg13g2_xor2_1 _5108_ (.B(_0990_),
    .A(_0989_),
    .X(_1005_));
 sg13g2_a21oi_1 _5109_ (.A1(_1004_),
    .A2(_1005_),
    .Y(_1006_),
    .B1(_0991_));
 sg13g2_and2_1 _5110_ (.A(_0979_),
    .B(_0980_),
    .X(_1007_));
 sg13g2_xor2_1 _5111_ (.B(_0980_),
    .A(_0979_),
    .X(_1009_));
 sg13g2_o21ai_1 _5112_ (.B1(_0981_),
    .Y(_1010_),
    .A1(_1006_),
    .A2(_1007_));
 sg13g2_xor2_1 _5113_ (.B(_0970_),
    .A(_0969_),
    .X(_1011_));
 sg13g2_a21oi_1 _5114_ (.A1(_1010_),
    .A2(_1011_),
    .Y(_1012_),
    .B1(_0971_));
 sg13g2_xor2_1 _5115_ (.B(_0958_),
    .A(_0949_),
    .X(_1013_));
 sg13g2_inv_1 _5116_ (.Y(_1014_),
    .A(_1013_));
 sg13g2_o21ai_1 _5117_ (.B1(_0959_),
    .Y(_1015_),
    .A1(_1012_),
    .A2(_1014_));
 sg13g2_xor2_1 _5118_ (.B(_0946_),
    .A(_0288_),
    .X(_1016_));
 sg13g2_xnor2_1 _5119_ (.Y(_1017_),
    .A(_0957_),
    .B(_1016_));
 sg13g2_xnor2_1 _5120_ (.Y(_1018_),
    .A(_1015_),
    .B(_1017_));
 sg13g2_xnor2_1 _5121_ (.Y(_1020_),
    .A(_1012_),
    .B(_1013_));
 sg13g2_xnor2_1 _5122_ (.Y(_1021_),
    .A(_1010_),
    .B(_1011_));
 sg13g2_xnor2_1 _5123_ (.Y(_1022_),
    .A(_1006_),
    .B(_1009_));
 sg13g2_xor2_1 _5124_ (.B(_1005_),
    .A(_1004_),
    .X(_1023_));
 sg13g2_xor2_1 _5125_ (.B(_1003_),
    .A(_1002_),
    .X(_1024_));
 sg13g2_xor2_1 _5126_ (.B(_1001_),
    .A(_0995_),
    .X(_1025_));
 sg13g2_nor3_1 _5127_ (.A(_1023_),
    .B(_1024_),
    .C(_1025_),
    .Y(_1026_));
 sg13g2_nand2_1 _5128_ (.Y(_1027_),
    .A(_1021_),
    .B(_1026_));
 sg13g2_o21ai_1 _5129_ (.B1(_1020_),
    .Y(_1028_),
    .A1(_1022_),
    .A2(_1027_));
 sg13g2_nand3_1 _5130_ (.B(_1023_),
    .C(_1024_),
    .A(_1022_),
    .Y(_1029_));
 sg13g2_nor2_1 _5131_ (.A(_1021_),
    .B(_1029_),
    .Y(_1031_));
 sg13g2_nor2_1 _5132_ (.A(net529),
    .B(_0334_),
    .Y(_1032_));
 sg13g2_nor2_2 _5133_ (.A(_2651_),
    .B(_0361_),
    .Y(_1033_));
 sg13g2_nand2_1 _5134_ (.Y(_1034_),
    .A(_0727_),
    .B(_1033_));
 sg13g2_nor2_1 _5135_ (.A(net587),
    .B(_0332_),
    .Y(_1035_));
 sg13g2_nand4_1 _5136_ (.B(_0727_),
    .C(_1033_),
    .A(_2610_),
    .Y(_1036_),
    .D(_1035_));
 sg13g2_a21oi_2 _5137_ (.B1(_0321_),
    .Y(_1037_),
    .A2(_1036_),
    .A1(_1032_));
 sg13g2_a21oi_2 _5138_ (.B1(_1037_),
    .Y(_1038_),
    .A2(_0309_),
    .A1(_2923_));
 sg13g2_o21ai_1 _5139_ (.B1(_1038_),
    .Y(_1039_),
    .A1(_1020_),
    .A2(_1031_));
 sg13g2_nand3b_1 _5140_ (.B(_1028_),
    .C(_1018_),
    .Y(_1040_),
    .A_N(_1039_));
 sg13g2_nor2b_1 _5141_ (.A(_0315_),
    .B_N(_0491_),
    .Y(_1042_));
 sg13g2_nand2_1 _5142_ (.Y(_1043_),
    .A(net570),
    .B(net557));
 sg13g2_nor2b_1 _5143_ (.A(net554),
    .B_N(net573),
    .Y(_1044_));
 sg13g2_xnor2_1 _5144_ (.Y(_1045_),
    .A(net573),
    .B(net554));
 sg13g2_a21o_1 _5145_ (.A2(_1045_),
    .A1(_0381_),
    .B1(_1044_),
    .X(_1046_));
 sg13g2_xor2_1 _5146_ (.B(net555),
    .A(net569),
    .X(_1047_));
 sg13g2_o21ai_1 _5147_ (.B1(_1047_),
    .Y(_1048_),
    .A1(\hvsync_gen.vpos[3] ),
    .A2(_1046_));
 sg13g2_a21oi_2 _5148_ (.B1(_0008_),
    .Y(_1049_),
    .A2(_1048_),
    .A1(_1043_));
 sg13g2_xnor2_1 _5149_ (.Y(_1050_),
    .A(_1008_),
    .B(_1049_));
 sg13g2_nand3_1 _5150_ (.B(_1043_),
    .C(_1048_),
    .A(_0008_),
    .Y(_1051_));
 sg13g2_nor2b_2 _5151_ (.A(_1049_),
    .B_N(_1051_),
    .Y(_1053_));
 sg13g2_or3_1 _5152_ (.A(\hvsync_gen.vpos[3] ),
    .B(_1046_),
    .C(_1047_),
    .X(_1054_));
 sg13g2_and2_2 _5153_ (.A(_1048_),
    .B(_1054_),
    .X(_1055_));
 sg13g2_nor3_2 _5154_ (.A(_1050_),
    .B(_1053_),
    .C(_1055_),
    .Y(_1056_));
 sg13g2_inv_1 _5155_ (.Y(_1057_),
    .A(_1056_));
 sg13g2_xor2_1 _5156_ (.B(net554),
    .A(\hvsync_gen.vpos[7] ),
    .X(_1058_));
 sg13g2_a21oi_1 _5157_ (.A1(_0535_),
    .A2(_1049_),
    .Y(_1059_),
    .B1(_0997_));
 sg13g2_xnor2_1 _5158_ (.Y(_1060_),
    .A(_1058_),
    .B(_1059_));
 sg13g2_nand2_1 _5159_ (.Y(_1061_),
    .A(_1056_),
    .B(_1060_));
 sg13g2_nor2_1 _5160_ (.A(_0008_),
    .B(_1043_),
    .Y(_1062_));
 sg13g2_a21oi_1 _5161_ (.A1(_2993_),
    .A2(_3004_),
    .Y(_1064_),
    .B1(net556));
 sg13g2_a221oi_1 _5162_ (.B2(_0162_),
    .C1(_1064_),
    .B1(_1062_),
    .A1(_1056_),
    .Y(_1065_),
    .A2(_1060_));
 sg13g2_xnor2_1 _5163_ (.Y(_1066_),
    .A(_1042_),
    .B(_1065_));
 sg13g2_o21ai_1 _5164_ (.B1(_0491_),
    .Y(_1067_),
    .A1(_0315_),
    .A2(_1065_));
 sg13g2_xnor2_1 _5165_ (.Y(_1068_),
    .A(_3147_),
    .B(_1067_));
 sg13g2_xnor2_1 _5166_ (.Y(_1069_),
    .A(net561),
    .B(_1067_));
 sg13g2_nand2b_1 _5167_ (.Y(_1070_),
    .B(_1068_),
    .A_N(_1066_));
 sg13g2_xor2_1 _5168_ (.B(_1046_),
    .A(_0009_),
    .X(_1071_));
 sg13g2_nand3b_1 _5169_ (.B(_1045_),
    .C(_0689_),
    .Y(_1072_),
    .A_N(_1071_));
 sg13g2_nor2_1 _5170_ (.A(_1061_),
    .B(_1072_),
    .Y(_1073_));
 sg13g2_nand2_1 _5171_ (.Y(_1075_),
    .A(_1068_),
    .B(_1072_));
 sg13g2_o21ai_1 _5172_ (.B1(_1066_),
    .Y(_1076_),
    .A1(_1069_),
    .A2(_1073_));
 sg13g2_and2_2 _5173_ (.A(_1070_),
    .B(_1076_),
    .X(_1077_));
 sg13g2_nand2_2 _5174_ (.Y(_1078_),
    .A(_1070_),
    .B(_1076_));
 sg13g2_nor3_1 _5175_ (.A(_1053_),
    .B(_1055_),
    .C(_1072_),
    .Y(_1079_));
 sg13g2_o21ai_1 _5176_ (.B1(_1068_),
    .Y(_1080_),
    .A1(_1057_),
    .A2(_1072_));
 sg13g2_xnor2_1 _5177_ (.Y(_1081_),
    .A(_1060_),
    .B(_1080_));
 sg13g2_o21ai_1 _5178_ (.B1(_1068_),
    .Y(_1082_),
    .A1(_1055_),
    .A2(_1072_));
 sg13g2_nor2_1 _5179_ (.A(_1069_),
    .B(_1079_),
    .Y(_1083_));
 sg13g2_xnor2_1 _5180_ (.Y(_1084_),
    .A(_1050_),
    .B(_1083_));
 sg13g2_a21oi_2 _5181_ (.B1(_1078_),
    .Y(_1086_),
    .A2(_1084_),
    .A1(_1081_));
 sg13g2_a21o_1 _5182_ (.A2(_1084_),
    .A1(_1081_),
    .B1(_1078_),
    .X(_1087_));
 sg13g2_nor2_1 _5183_ (.A(_1078_),
    .B(_1086_),
    .Y(_1088_));
 sg13g2_nand2_2 _5184_ (.Y(_1089_),
    .A(_1077_),
    .B(net491));
 sg13g2_xnor2_1 _5185_ (.Y(_1090_),
    .A(_1053_),
    .B(_1082_));
 sg13g2_xor2_1 _5186_ (.B(_1082_),
    .A(_1053_),
    .X(_1091_));
 sg13g2_nand4_1 _5187_ (.B(_1081_),
    .C(_1084_),
    .A(_1077_),
    .Y(_1092_),
    .D(_1091_));
 sg13g2_a21o_1 _5188_ (.A2(_1045_),
    .A1(_0689_),
    .B1(_1069_),
    .X(_1093_));
 sg13g2_xor2_1 _5189_ (.B(_1093_),
    .A(_1071_),
    .X(_1094_));
 sg13g2_xnor2_1 _5190_ (.Y(_1095_),
    .A(net555),
    .B(_0766_));
 sg13g2_o21ai_1 _5191_ (.B1(_1095_),
    .Y(_1097_),
    .A1(_0689_),
    .A2(_1069_));
 sg13g2_or3_1 _5192_ (.A(_0689_),
    .B(_1069_),
    .C(_1095_),
    .X(_1098_));
 sg13g2_nand2_1 _5193_ (.Y(_1099_),
    .A(_1097_),
    .B(_1098_));
 sg13g2_and2_1 _5194_ (.A(_1097_),
    .B(_1098_),
    .X(_1100_));
 sg13g2_nand2_1 _5195_ (.Y(_1101_),
    .A(_1094_),
    .B(_1100_));
 sg13g2_nand3_1 _5196_ (.B(_1068_),
    .C(_1072_),
    .A(_1055_),
    .Y(_1102_));
 sg13g2_nand2b_1 _5197_ (.Y(_1103_),
    .B(_1075_),
    .A_N(_1055_));
 sg13g2_xnor2_1 _5198_ (.Y(_1104_),
    .A(_1055_),
    .B(_1075_));
 sg13g2_inv_1 _5199_ (.Y(_1105_),
    .A(_1104_));
 sg13g2_nor2_1 _5200_ (.A(_1092_),
    .B(_1104_),
    .Y(_1106_));
 sg13g2_a21oi_2 _5201_ (.B1(_1086_),
    .Y(_1108_),
    .A2(_1106_),
    .A1(_1101_));
 sg13g2_inv_1 _5202_ (.Y(_1109_),
    .A(_1108_));
 sg13g2_or3_1 _5203_ (.A(_1066_),
    .B(_1069_),
    .C(_1073_),
    .X(_1110_));
 sg13g2_nand2_2 _5204_ (.Y(_1111_),
    .A(_1076_),
    .B(_1110_));
 sg13g2_nand3_1 _5205_ (.B(_0711_),
    .C(_1068_),
    .A(_0006_),
    .Y(_1112_));
 sg13g2_a21o_1 _5206_ (.A2(_1068_),
    .A1(_0006_),
    .B1(_0711_),
    .X(_1113_));
 sg13g2_and2_1 _5207_ (.A(_1112_),
    .B(_1113_),
    .X(_1114_));
 sg13g2_nand4_1 _5208_ (.B(_1098_),
    .C(_1112_),
    .A(_1097_),
    .Y(_1115_),
    .D(_1113_));
 sg13g2_a21oi_1 _5209_ (.A1(_1094_),
    .A2(_1115_),
    .Y(_1116_),
    .B1(_1104_));
 sg13g2_o21ai_1 _5210_ (.B1(_1084_),
    .Y(_1117_),
    .A1(_1090_),
    .A2(_1116_));
 sg13g2_and2_1 _5211_ (.A(_1070_),
    .B(_1081_),
    .X(_1119_));
 sg13g2_a21oi_2 _5212_ (.B1(_1111_),
    .Y(_1120_),
    .A2(_1119_),
    .A1(_1117_));
 sg13g2_a21o_2 _5213_ (.A2(_1119_),
    .A1(_1117_),
    .B1(_1111_),
    .X(_1121_));
 sg13g2_nor2_1 _5214_ (.A(_1081_),
    .B(_1120_),
    .Y(_1122_));
 sg13g2_a221oi_1 _5215_ (.B2(_1119_),
    .C1(_1111_),
    .B1(_1117_),
    .A1(_1102_),
    .Y(_1123_),
    .A2(_1103_));
 sg13g2_o21ai_1 _5216_ (.B1(_1077_),
    .Y(_1124_),
    .A1(_1090_),
    .A2(_1104_));
 sg13g2_or2_1 _5217_ (.X(_1125_),
    .B(_1106_),
    .A(_1094_));
 sg13g2_a221oi_1 _5218_ (.B2(_1121_),
    .C1(_1123_),
    .B1(_1125_),
    .A1(net491),
    .Y(_1126_),
    .A2(_1124_));
 sg13g2_o21ai_1 _5219_ (.B1(_1108_),
    .Y(_1127_),
    .A1(_1122_),
    .A2(_1126_));
 sg13g2_mux2_1 _5220_ (.A0(_1084_),
    .A1(_1091_),
    .S(_1121_),
    .X(_1128_));
 sg13g2_a21o_1 _5221_ (.A2(_1128_),
    .A1(_1086_),
    .B1(_1078_),
    .X(_1130_));
 sg13g2_nor2_1 _5222_ (.A(_1089_),
    .B(_1104_),
    .Y(_1131_));
 sg13g2_a21oi_2 _5223_ (.B1(_1131_),
    .Y(_1132_),
    .A2(_1130_),
    .A1(_1127_));
 sg13g2_a21o_2 _5224_ (.A2(_1130_),
    .A1(_1127_),
    .B1(_1131_),
    .X(_1133_));
 sg13g2_mux2_1 _5225_ (.A0(_1091_),
    .A1(_1105_),
    .S(_1121_),
    .X(_1134_));
 sg13g2_nor2_1 _5226_ (.A(_1078_),
    .B(_1134_),
    .Y(_1135_));
 sg13g2_and3_1 _5227_ (.X(_1136_),
    .A(net491),
    .B(_1108_),
    .C(_1124_));
 sg13g2_nand2_1 _5228_ (.Y(_1137_),
    .A(_1084_),
    .B(_1121_));
 sg13g2_a21o_1 _5229_ (.A2(_1137_),
    .A1(_1136_),
    .B1(net487),
    .X(_1138_));
 sg13g2_nand2_1 _5230_ (.Y(_1139_),
    .A(_1078_),
    .B(_1120_));
 sg13g2_a22oi_1 _5231_ (.Y(_1141_),
    .B1(_1120_),
    .B2(_1078_),
    .A2(_1094_),
    .A1(net487));
 sg13g2_o21ai_1 _5232_ (.B1(_1141_),
    .Y(_1142_),
    .A1(_1135_),
    .A2(_1138_));
 sg13g2_inv_1 _5233_ (.Y(_1143_),
    .A(_1142_));
 sg13g2_nor2_1 _5234_ (.A(_1089_),
    .B(_1100_),
    .Y(_1144_));
 sg13g2_or3_1 _5235_ (.A(_1108_),
    .B(_1122_),
    .C(_1126_),
    .X(_1145_));
 sg13g2_a21oi_1 _5236_ (.A1(_1128_),
    .A2(_1136_),
    .Y(_1146_),
    .B1(net487));
 sg13g2_a21oi_2 _5237_ (.B1(_1144_),
    .Y(_1147_),
    .A2(_1146_),
    .A1(_1145_));
 sg13g2_a21o_2 _5238_ (.A2(_1146_),
    .A1(_1145_),
    .B1(_1144_),
    .X(_1148_));
 sg13g2_nor2_1 _5239_ (.A(_1133_),
    .B(_1147_),
    .Y(_1149_));
 sg13g2_o21ai_1 _5240_ (.B1(_1142_),
    .Y(_1150_),
    .A1(_1133_),
    .A2(_1147_));
 sg13g2_or2_1 _5241_ (.X(_1152_),
    .B(_1142_),
    .A(_1133_));
 sg13g2_xnor2_1 _5242_ (.Y(_1153_),
    .A(_1092_),
    .B(_1152_));
 sg13g2_and2_1 _5243_ (.A(_1150_),
    .B(_1153_),
    .X(_1154_));
 sg13g2_inv_1 _5244_ (.Y(_1155_),
    .A(_1154_));
 sg13g2_o21ai_1 _5245_ (.B1(_1099_),
    .Y(_1156_),
    .A1(_1092_),
    .A2(_1104_));
 sg13g2_mux2_1 _5246_ (.A0(_1125_),
    .A1(_1156_),
    .S(_1121_),
    .X(_1157_));
 sg13g2_a221oi_1 _5247_ (.B2(_1109_),
    .C1(net487),
    .B1(_1157_),
    .A1(_1134_),
    .Y(_1158_),
    .A2(_1136_));
 sg13g2_a21o_2 _5248_ (.A2(_1114_),
    .A1(net487),
    .B1(_1158_),
    .X(_1159_));
 sg13g2_nand2_1 _5249_ (.Y(_1160_),
    .A(_1132_),
    .B(_1159_));
 sg13g2_nand2_1 _5250_ (.Y(_1161_),
    .A(_1092_),
    .B(_1148_));
 sg13g2_and2_2 _5251_ (.A(_1092_),
    .B(_1159_),
    .X(_1163_));
 sg13g2_nor2_1 _5252_ (.A(_1160_),
    .B(_1161_),
    .Y(_1164_));
 sg13g2_nand2_1 _5253_ (.Y(_1165_),
    .A(_1149_),
    .B(_1163_));
 sg13g2_and2_1 _5254_ (.A(\hvsync_gen.vpos[0] ),
    .B(net488),
    .X(_1166_));
 sg13g2_o21ai_1 _5255_ (.B1(net487),
    .Y(_1167_),
    .A1(net581),
    .A2(_1091_));
 sg13g2_nor2_1 _5256_ (.A(_1133_),
    .B(_1166_),
    .Y(_1168_));
 sg13g2_nand3_1 _5257_ (.B(_1159_),
    .C(_1167_),
    .A(_1132_),
    .Y(_1169_));
 sg13g2_nor2_1 _5258_ (.A(_1142_),
    .B(_1147_),
    .Y(_1170_));
 sg13g2_nand2b_1 _5259_ (.Y(_1171_),
    .B(_1148_),
    .A_N(_1142_));
 sg13g2_a21oi_1 _5260_ (.A1(_1132_),
    .A2(_1159_),
    .Y(_1172_),
    .B1(_1167_));
 sg13g2_a21o_1 _5261_ (.A2(_1159_),
    .A1(_1132_),
    .B1(_1167_),
    .X(_1174_));
 sg13g2_o21ai_1 _5262_ (.B1(_1169_),
    .Y(_1175_),
    .A1(_1171_),
    .A2(_1172_));
 sg13g2_xor2_1 _5263_ (.B(_1163_),
    .A(_1149_),
    .X(_1176_));
 sg13g2_xnor2_1 _5264_ (.Y(_1177_),
    .A(_1175_),
    .B(_1176_));
 sg13g2_o21ai_1 _5265_ (.B1(_1150_),
    .Y(_1178_),
    .A1(_1147_),
    .A2(_1152_));
 sg13g2_xor2_1 _5266_ (.B(_1178_),
    .A(_1163_),
    .X(_1179_));
 sg13g2_or3_1 _5267_ (.A(_1165_),
    .B(_1177_),
    .C(_1179_),
    .X(_1180_));
 sg13g2_a22oi_1 _5268_ (.Y(_1181_),
    .B1(_1170_),
    .B2(_1132_),
    .A2(_1163_),
    .A1(_1150_));
 sg13g2_inv_1 _5269_ (.Y(_1182_),
    .A(_1181_));
 sg13g2_a21oi_1 _5270_ (.A1(_1175_),
    .A2(_1176_),
    .Y(_1183_),
    .B1(_1164_));
 sg13g2_o21ai_1 _5271_ (.B1(_1183_),
    .Y(_1185_),
    .A1(_1177_),
    .A2(_1179_));
 sg13g2_nand3_1 _5272_ (.B(_1182_),
    .C(_1185_),
    .A(_1180_),
    .Y(_1186_));
 sg13g2_and2_1 _5273_ (.A(_1180_),
    .B(_1186_),
    .X(_1187_));
 sg13g2_nand2_1 _5274_ (.Y(_1188_),
    .A(_1132_),
    .B(_1142_));
 sg13g2_xor2_1 _5275_ (.B(_1188_),
    .A(_1161_),
    .X(_1189_));
 sg13g2_nor2b_1 _5276_ (.A(_1187_),
    .B_N(_1189_),
    .Y(_1190_));
 sg13g2_a21oi_1 _5277_ (.A1(_1169_),
    .A2(_1174_),
    .Y(_1191_),
    .B1(_1171_));
 sg13g2_nand3_1 _5278_ (.B(_1171_),
    .C(_1174_),
    .A(_1169_),
    .Y(_1192_));
 sg13g2_nand2b_1 _5279_ (.Y(_1193_),
    .B(_1192_),
    .A_N(_1191_));
 sg13g2_mux2_1 _5280_ (.A0(_1175_),
    .A1(_1193_),
    .S(_1143_),
    .X(_1194_));
 sg13g2_a21o_1 _5281_ (.A2(_1185_),
    .A1(_1180_),
    .B1(_1182_),
    .X(_1196_));
 sg13g2_and3_1 _5282_ (.X(_1197_),
    .A(_1186_),
    .B(_1194_),
    .C(_1196_));
 sg13g2_nand3_1 _5283_ (.B(_1194_),
    .C(_1196_),
    .A(_1186_),
    .Y(_1198_));
 sg13g2_xnor2_1 _5284_ (.Y(_1199_),
    .A(_1143_),
    .B(_1193_));
 sg13g2_a21oi_1 _5285_ (.A1(_1143_),
    .A2(_1159_),
    .Y(_1200_),
    .B1(_1168_));
 sg13g2_nor2_1 _5286_ (.A(_1142_),
    .B(_1166_),
    .Y(_1201_));
 sg13g2_nor2b_1 _5287_ (.A(_1160_),
    .B_N(_1201_),
    .Y(_1202_));
 sg13g2_nand2_1 _5288_ (.Y(_1203_),
    .A(_1148_),
    .B(_1159_));
 sg13g2_nor2_1 _5289_ (.A(_1200_),
    .B(_1203_),
    .Y(_1204_));
 sg13g2_nor2_1 _5290_ (.A(_1202_),
    .B(_1204_),
    .Y(_1205_));
 sg13g2_nor2_1 _5291_ (.A(_1199_),
    .B(_1205_),
    .Y(_1207_));
 sg13g2_nor2_1 _5292_ (.A(_1166_),
    .B(_1171_),
    .Y(_1208_));
 sg13g2_nor2_1 _5293_ (.A(_1200_),
    .B(_1202_),
    .Y(_1209_));
 sg13g2_xnor2_1 _5294_ (.Y(_1210_),
    .A(_1203_),
    .B(_1209_));
 sg13g2_and2_1 _5295_ (.A(_1208_),
    .B(_1210_),
    .X(_1211_));
 sg13g2_xor2_1 _5296_ (.B(_1205_),
    .A(_1199_),
    .X(_1212_));
 sg13g2_a21oi_2 _5297_ (.B1(_1207_),
    .Y(_1213_),
    .A2(_1212_),
    .A1(_1211_));
 sg13g2_a21oi_1 _5298_ (.A1(_1186_),
    .A2(_1196_),
    .Y(_1214_),
    .B1(_1194_));
 sg13g2_nor3_1 _5299_ (.A(_1197_),
    .B(_1213_),
    .C(_1214_),
    .Y(_1215_));
 sg13g2_o21ai_1 _5300_ (.B1(_1198_),
    .Y(_1216_),
    .A1(_1213_),
    .A2(_1214_));
 sg13g2_xnor2_1 _5301_ (.Y(_1218_),
    .A(_1187_),
    .B(_1189_));
 sg13g2_a21oi_1 _5302_ (.A1(_1216_),
    .A2(_1218_),
    .Y(_1219_),
    .B1(_1190_));
 sg13g2_o21ai_1 _5303_ (.B1(_1133_),
    .Y(_1220_),
    .A1(_1155_),
    .A2(_1219_));
 sg13g2_nand3_1 _5304_ (.B(_1092_),
    .C(_1220_),
    .A(net487),
    .Y(_1221_));
 sg13g2_nor2_1 _5305_ (.A(net487),
    .B(_1120_),
    .Y(_1222_));
 sg13g2_xnor2_1 _5306_ (.Y(_1223_),
    .A(_1154_),
    .B(_1219_));
 sg13g2_o21ai_1 _5307_ (.B1(_1213_),
    .Y(_1224_),
    .A1(_1197_),
    .A2(_1214_));
 sg13g2_nand2b_1 _5308_ (.Y(_1225_),
    .B(_1224_),
    .A_N(_1215_));
 sg13g2_o21ai_1 _5309_ (.B1(_1086_),
    .Y(_1226_),
    .A1(_1121_),
    .A2(_1225_));
 sg13g2_a21oi_1 _5310_ (.A1(net476),
    .A2(_1223_),
    .Y(_1227_),
    .B1(_1226_));
 sg13g2_xor2_1 _5311_ (.B(_1210_),
    .A(_1208_),
    .X(_1229_));
 sg13g2_xnor2_1 _5312_ (.Y(_1230_),
    .A(_1147_),
    .B(_1159_));
 sg13g2_a22oi_1 _5313_ (.Y(_1231_),
    .B1(_1230_),
    .B2(_1120_),
    .A2(_1229_),
    .A1(net476));
 sg13g2_a21o_1 _5314_ (.A2(_1231_),
    .A1(_1087_),
    .B1(net488),
    .X(_1232_));
 sg13g2_o21ai_1 _5315_ (.B1(_1221_),
    .Y(_1233_),
    .A1(_1227_),
    .A2(_1232_));
 sg13g2_inv_4 _5316_ (.A(net467),
    .Y(_1234_));
 sg13g2_nand2_1 _5317_ (.Y(_1235_),
    .A(_1152_),
    .B(_1220_));
 sg13g2_xor2_1 _5318_ (.B(_1218_),
    .A(_1216_),
    .X(_1236_));
 sg13g2_a221oi_1 _5319_ (.B2(_1120_),
    .C1(net491),
    .B1(_1236_),
    .A1(net476),
    .Y(_1237_),
    .A2(_1235_));
 sg13g2_xnor2_1 _5320_ (.Y(_1238_),
    .A(_1211_),
    .B(_1212_));
 sg13g2_xnor2_1 _5321_ (.Y(_1240_),
    .A(_1148_),
    .B(_1201_));
 sg13g2_a21oi_1 _5322_ (.A1(_1114_),
    .A2(_1166_),
    .Y(_1241_),
    .B1(_1240_));
 sg13g2_nand2_1 _5323_ (.Y(_1242_),
    .A(net476),
    .B(_1238_));
 sg13g2_o21ai_1 _5324_ (.B1(_1242_),
    .Y(_1243_),
    .A1(_1222_),
    .A2(_1241_));
 sg13g2_a21oi_1 _5325_ (.A1(_1078_),
    .A2(_1243_),
    .Y(_1244_),
    .B1(net488));
 sg13g2_nand2b_2 _5326_ (.Y(_1245_),
    .B(_1244_),
    .A_N(_1237_));
 sg13g2_xnor2_1 _5327_ (.Y(_1246_),
    .A(net468),
    .B(net467));
 sg13g2_nor2_1 _5328_ (.A(net466),
    .B(_1246_),
    .Y(_1247_));
 sg13g2_a21oi_1 _5329_ (.A1(net468),
    .A2(net467),
    .Y(_1248_),
    .B1(_1247_));
 sg13g2_nand2_1 _5330_ (.Y(_1249_),
    .A(_1120_),
    .B(_1223_));
 sg13g2_a21oi_1 _5331_ (.A1(_1121_),
    .A2(_1220_),
    .Y(_1251_),
    .B1(net491));
 sg13g2_nand2_1 _5332_ (.Y(_1252_),
    .A(net476),
    .B(_1225_));
 sg13g2_o21ai_1 _5333_ (.B1(_1252_),
    .Y(_1253_),
    .A1(net476),
    .A2(_1229_));
 sg13g2_a22oi_1 _5334_ (.Y(_1254_),
    .B1(_1253_),
    .B2(net491),
    .A2(_1251_),
    .A1(_1249_));
 sg13g2_nand2_1 _5335_ (.Y(_1255_),
    .A(_1089_),
    .B(_1254_));
 sg13g2_xor2_1 _5336_ (.B(net466),
    .A(net470),
    .X(_1256_));
 sg13g2_nand2b_1 _5337_ (.Y(_1257_),
    .B(_1256_),
    .A_N(net464));
 sg13g2_xor2_1 _5338_ (.B(_1256_),
    .A(net464),
    .X(_1258_));
 sg13g2_or2_1 _5339_ (.X(_1259_),
    .B(_1258_),
    .A(_1248_));
 sg13g2_and3_1 _5340_ (.X(_1260_),
    .A(_1092_),
    .B(_1120_),
    .C(_1235_));
 sg13g2_nor2_1 _5341_ (.A(_1077_),
    .B(_1241_),
    .Y(_1262_));
 sg13g2_nor2_1 _5342_ (.A(net476),
    .B(_1238_),
    .Y(_1263_));
 sg13g2_a21oi_1 _5343_ (.A1(net476),
    .A2(_1236_),
    .Y(_1264_),
    .B1(_1263_));
 sg13g2_a21oi_1 _5344_ (.A1(_1086_),
    .A2(_1264_),
    .Y(_1265_),
    .B1(_1262_));
 sg13g2_o21ai_1 _5345_ (.B1(_1265_),
    .Y(_1266_),
    .A1(_1089_),
    .A2(_1260_));
 sg13g2_nand2b_1 _5346_ (.Y(_1267_),
    .B(_2855_),
    .A_N(net462));
 sg13g2_xnor2_1 _5347_ (.Y(_1268_),
    .A(_2856_),
    .B(net461));
 sg13g2_o21ai_1 _5348_ (.B1(_1267_),
    .Y(_1269_),
    .A1(_1234_),
    .A2(_1268_));
 sg13g2_xor2_1 _5349_ (.B(_1246_),
    .A(net466),
    .X(_1270_));
 sg13g2_nand2_1 _5350_ (.Y(_1271_),
    .A(_1111_),
    .B(_1230_));
 sg13g2_o21ai_1 _5351_ (.B1(_1271_),
    .Y(_1273_),
    .A1(net491),
    .A2(_1253_));
 sg13g2_a21oi_2 _5352_ (.B1(_1273_),
    .Y(_1274_),
    .A2(_1223_),
    .A1(net488));
 sg13g2_a21o_2 _5353_ (.A2(_1223_),
    .A1(net488),
    .B1(_1273_),
    .X(_1275_));
 sg13g2_nand2b_1 _5354_ (.Y(_1276_),
    .B(_1275_),
    .A_N(_2872_));
 sg13g2_xnor2_1 _5355_ (.Y(_1277_),
    .A(net475),
    .B(_1274_));
 sg13g2_o21ai_1 _5356_ (.B1(_1276_),
    .Y(_1278_),
    .A1(net462),
    .A2(_1277_));
 sg13g2_xnor2_1 _5357_ (.Y(_1279_),
    .A(net467),
    .B(_1268_));
 sg13g2_nand2_1 _5358_ (.Y(_1280_),
    .A(_1278_),
    .B(_1279_));
 sg13g2_o21ai_1 _5359_ (.B1(_1139_),
    .Y(_1281_),
    .A1(net491),
    .A2(_1243_));
 sg13g2_a21oi_2 _5360_ (.B1(_1281_),
    .Y(_1282_),
    .A2(_1236_),
    .A1(net488));
 sg13g2_inv_1 _5361_ (.Y(_1284_),
    .A(_1282_));
 sg13g2_nor2_1 _5362_ (.A(net473),
    .B(_1282_),
    .Y(_1285_));
 sg13g2_xnor2_1 _5363_ (.Y(_1286_),
    .A(net473),
    .B(_1282_));
 sg13g2_nor2_1 _5364_ (.A(_1274_),
    .B(_1286_),
    .Y(_1287_));
 sg13g2_nor2_1 _5365_ (.A(_1285_),
    .B(_1287_),
    .Y(_1288_));
 sg13g2_xor2_1 _5366_ (.B(_1277_),
    .A(net462),
    .X(_1289_));
 sg13g2_nor2b_1 _5367_ (.A(_1288_),
    .B_N(_1289_),
    .Y(_1290_));
 sg13g2_xnor2_1 _5368_ (.Y(_1291_),
    .A(_1275_),
    .B(_1286_));
 sg13g2_nor2_1 _5369_ (.A(_2895_),
    .B(_1282_),
    .Y(_1292_));
 sg13g2_and2_1 _5370_ (.A(_1291_),
    .B(_1292_),
    .X(_1293_));
 sg13g2_xnor2_1 _5371_ (.Y(_1295_),
    .A(_1288_),
    .B(_1289_));
 sg13g2_a21oi_1 _5372_ (.A1(_1293_),
    .A2(_1295_),
    .Y(_1296_),
    .B1(_1290_));
 sg13g2_xnor2_1 _5373_ (.Y(_1297_),
    .A(_1278_),
    .B(_1279_));
 sg13g2_o21ai_1 _5374_ (.B1(_1280_),
    .Y(_1298_),
    .A1(_1296_),
    .A2(_1297_));
 sg13g2_xnor2_1 _5375_ (.Y(_1299_),
    .A(_1269_),
    .B(_1270_));
 sg13g2_nor2b_1 _5376_ (.A(_1299_),
    .B_N(_1298_),
    .Y(_1300_));
 sg13g2_a21oi_1 _5377_ (.A1(_1269_),
    .A2(_1270_),
    .Y(_1301_),
    .B1(_1300_));
 sg13g2_xnor2_1 _5378_ (.Y(_1302_),
    .A(_1248_),
    .B(_1258_));
 sg13g2_o21ai_1 _5379_ (.B1(_1259_),
    .Y(_1303_),
    .A1(_1301_),
    .A2(_1302_));
 sg13g2_o21ai_1 _5380_ (.B1(_1257_),
    .Y(_1304_),
    .A1(net470),
    .A2(net466));
 sg13g2_nand2_1 _5381_ (.Y(_1306_),
    .A(_1086_),
    .B(_1260_));
 sg13g2_o21ai_1 _5382_ (.B1(_1306_),
    .Y(_1307_),
    .A1(_1077_),
    .A2(_1264_));
 sg13g2_inv_4 _5383_ (.A(_1307_),
    .Y(_1308_));
 sg13g2_xor2_1 _5384_ (.B(_1307_),
    .A(net464),
    .X(_1309_));
 sg13g2_xor2_1 _5385_ (.B(_1309_),
    .A(_2912_),
    .X(_1310_));
 sg13g2_xnor2_1 _5386_ (.Y(_1311_),
    .A(_1304_),
    .B(_1310_));
 sg13g2_xnor2_1 _5387_ (.Y(_1312_),
    .A(_1303_),
    .B(_1311_));
 sg13g2_xor2_1 _5388_ (.B(_1302_),
    .A(_1301_),
    .X(_1313_));
 sg13g2_xor2_1 _5389_ (.B(_1299_),
    .A(_1298_),
    .X(_1314_));
 sg13g2_xnor2_1 _5390_ (.Y(_1315_),
    .A(_1296_),
    .B(_1297_));
 sg13g2_xnor2_1 _5391_ (.Y(_1317_),
    .A(_1293_),
    .B(_1295_));
 sg13g2_nand3_1 _5392_ (.B(_1315_),
    .C(_1317_),
    .A(_1314_),
    .Y(_1318_));
 sg13g2_and2_1 _5393_ (.A(_1313_),
    .B(_1318_),
    .X(_1319_));
 sg13g2_nand2_1 _5394_ (.Y(_1320_),
    .A(_2895_),
    .B(_1282_));
 sg13g2_a21oi_1 _5395_ (.A1(_1291_),
    .A2(_1320_),
    .Y(_1321_),
    .B1(_1295_));
 sg13g2_a21o_1 _5396_ (.A2(_1295_),
    .A1(_1293_),
    .B1(_1321_),
    .X(_1322_));
 sg13g2_nor3_1 _5397_ (.A(_1314_),
    .B(_1315_),
    .C(_1322_),
    .Y(_1323_));
 sg13g2_nor2_1 _5398_ (.A(_1313_),
    .B(_1323_),
    .Y(_1324_));
 sg13g2_or2_1 _5399_ (.X(_1325_),
    .B(_0056_),
    .A(net571));
 sg13g2_nand2_1 _5400_ (.Y(_1326_),
    .A(_2923_),
    .B(_2940_));
 sg13g2_a21oi_1 _5401_ (.A1(_0184_),
    .A2(_1325_),
    .Y(_1328_),
    .B1(_1326_));
 sg13g2_nor4_1 _5402_ (.A(_1312_),
    .B(_1319_),
    .C(_1324_),
    .D(_1328_),
    .Y(_1329_));
 sg13g2_a21oi_1 _5403_ (.A1(_2899_),
    .A2(_2931_),
    .Y(_1330_),
    .B1(_2932_));
 sg13g2_nor2b_1 _5404_ (.A(_2930_),
    .B_N(_1330_),
    .Y(_1331_));
 sg13g2_a21oi_1 _5405_ (.A1(_2927_),
    .A2(_1331_),
    .Y(_1332_),
    .B1(_2929_));
 sg13g2_a21oi_1 _5406_ (.A1(_2885_),
    .A2(_2895_),
    .Y(_1333_),
    .B1(_2896_));
 sg13g2_a21oi_1 _5407_ (.A1(_2899_),
    .A2(_1333_),
    .Y(_1334_),
    .B1(_2932_));
 sg13g2_mux2_1 _5408_ (.A0(_2933_),
    .A1(_1334_),
    .S(_2930_),
    .X(_1335_));
 sg13g2_nor2_1 _5409_ (.A(_2927_),
    .B(_1335_),
    .Y(_1336_));
 sg13g2_nor4_2 _5410_ (.A(_2922_),
    .B(_2935_),
    .C(_1332_),
    .Y(_1337_),
    .D(_1336_));
 sg13g2_xnor2_1 _5411_ (.Y(_1339_),
    .A(_3208_),
    .B(_3209_));
 sg13g2_nor3_1 _5412_ (.A(_3227_),
    .B(_3228_),
    .C(_1339_),
    .Y(_1340_));
 sg13g2_nor2_1 _5413_ (.A(_3226_),
    .B(_1340_),
    .Y(_1341_));
 sg13g2_nor3_2 _5414_ (.A(_3223_),
    .B(_3231_),
    .C(_1341_),
    .Y(_1342_));
 sg13g2_a21oi_1 _5415_ (.A1(_0335_),
    .A2(_0336_),
    .Y(_1343_),
    .B1(_0361_));
 sg13g2_a21o_1 _5416_ (.A2(_1343_),
    .A1(_0340_),
    .B1(_0339_),
    .X(_1344_));
 sg13g2_nand3_1 _5417_ (.B(_2598_),
    .C(_0331_),
    .A(net548),
    .Y(_1345_));
 sg13g2_a221oi_1 _5418_ (.B2(_1343_),
    .C1(_1345_),
    .B1(_0340_),
    .A1(_2641_),
    .Y(_1346_),
    .A2(_0338_));
 sg13g2_nor3_2 _5419_ (.A(net601),
    .B(_3202_),
    .C(net535),
    .Y(_1347_));
 sg13g2_a221oi_1 _5420_ (.B2(_2648_),
    .C1(_1347_),
    .B1(_0360_),
    .A1(_2649_),
    .Y(_1348_),
    .A2(_2650_));
 sg13g2_and3_1 _5421_ (.X(_1350_),
    .A(net543),
    .B(_0332_),
    .C(_1348_));
 sg13g2_or2_1 _5422_ (.X(_1351_),
    .B(_1350_),
    .A(_1346_));
 sg13g2_nor4_2 _5423_ (.A(_0324_),
    .B(_0330_),
    .C(_1346_),
    .Y(_1352_),
    .D(_1350_));
 sg13g2_o21ai_1 _5424_ (.B1(net529),
    .Y(_1353_),
    .A1(_0330_),
    .A2(_1351_));
 sg13g2_nor2b_2 _5425_ (.A(_1352_),
    .B_N(_1353_),
    .Y(_1354_));
 sg13g2_xnor2_1 _5426_ (.Y(_1355_),
    .A(_0329_),
    .B(_1351_));
 sg13g2_xnor2_1 _5427_ (.Y(_1356_),
    .A(_0330_),
    .B(_1351_));
 sg13g2_nor4_2 _5428_ (.A(_2614_),
    .B(_2623_),
    .C(_2625_),
    .Y(_1357_),
    .D(_0361_));
 sg13g2_nor2_1 _5429_ (.A(_2641_),
    .B(_1347_),
    .Y(_1358_));
 sg13g2_nor2b_1 _5430_ (.A(net596),
    .B_N(_1347_),
    .Y(_1359_));
 sg13g2_or3_1 _5431_ (.A(net548),
    .B(_1358_),
    .C(_1359_),
    .X(_1361_));
 sg13g2_o21ai_1 _5432_ (.B1(_1361_),
    .Y(_1362_),
    .A1(_0743_),
    .A2(_1357_));
 sg13g2_and2_1 _5433_ (.A(net542),
    .B(_2513_),
    .X(_1363_));
 sg13g2_a22oi_1 _5434_ (.Y(_1364_),
    .B1(_1363_),
    .B2(_0369_),
    .A2(_0729_),
    .A1(net553));
 sg13g2_nor2_1 _5435_ (.A(net552),
    .B(net602),
    .Y(_1365_));
 sg13g2_a21oi_2 _5436_ (.B1(_1365_),
    .Y(_1366_),
    .A2(_2614_),
    .A1(net552));
 sg13g2_a21oi_2 _5437_ (.B1(_0051_),
    .Y(_1367_),
    .A2(_2619_),
    .A1(net551));
 sg13g2_or2_1 _5438_ (.X(_1368_),
    .B(_1367_),
    .A(_0375_));
 sg13g2_or2_1 _5439_ (.X(_1369_),
    .B(_1368_),
    .A(_1366_));
 sg13g2_a221oi_1 _5440_ (.B2(_0369_),
    .C1(_1369_),
    .B1(_1363_),
    .A1(net553),
    .Y(_1370_),
    .A2(_0729_));
 sg13g2_xor2_1 _5441_ (.B(_1357_),
    .A(_2651_),
    .X(_1372_));
 sg13g2_xnor2_1 _5442_ (.Y(_1373_),
    .A(_0338_),
    .B(_1358_));
 sg13g2_mux2_2 _5443_ (.A0(_1372_),
    .A1(_1373_),
    .S(net539),
    .X(_1374_));
 sg13g2_and3_1 _5444_ (.X(_1375_),
    .A(_1362_),
    .B(_1370_),
    .C(_1374_));
 sg13g2_nor2_1 _5445_ (.A(net543),
    .B(_0332_),
    .Y(_1376_));
 sg13g2_xnor2_1 _5446_ (.Y(_1377_),
    .A(_0332_),
    .B(_1348_));
 sg13g2_a221oi_1 _5447_ (.B2(_3279_),
    .C1(_1346_),
    .B1(_1377_),
    .A1(_1344_),
    .Y(_1378_),
    .A2(_1376_));
 sg13g2_and4_1 _5448_ (.A(_1362_),
    .B(_1370_),
    .C(_1374_),
    .D(_1378_),
    .X(_1379_));
 sg13g2_nand2_1 _5449_ (.Y(_1380_),
    .A(_1356_),
    .B(_1379_));
 sg13g2_xnor2_1 _5450_ (.Y(_1381_),
    .A(_0322_),
    .B(_1352_));
 sg13g2_xnor2_1 _5451_ (.Y(_1383_),
    .A(_0321_),
    .B(_1352_));
 sg13g2_a21oi_2 _5452_ (.B1(_1381_),
    .Y(_1384_),
    .A2(_1379_),
    .A1(_1356_));
 sg13g2_xnor2_1 _5453_ (.Y(_1385_),
    .A(_1354_),
    .B(_1384_));
 sg13g2_xor2_1 _5454_ (.B(_1384_),
    .A(_1354_),
    .X(_1386_));
 sg13g2_a221oi_1 _5455_ (.B2(net543),
    .C1(_1346_),
    .B1(_1377_),
    .A1(_1344_),
    .Y(_1387_),
    .A2(_1376_));
 sg13g2_nand4_1 _5456_ (.B(_1370_),
    .C(_1374_),
    .A(_1362_),
    .Y(_1388_),
    .D(_1387_));
 sg13g2_and2_1 _5457_ (.A(_1383_),
    .B(_1388_),
    .X(_1389_));
 sg13g2_nand3_1 _5458_ (.B(_1383_),
    .C(_1388_),
    .A(_1355_),
    .Y(_1390_));
 sg13g2_a21o_1 _5459_ (.A2(_1388_),
    .A1(_1383_),
    .B1(_1355_),
    .X(_1391_));
 sg13g2_nand2_1 _5460_ (.Y(_1392_),
    .A(_1390_),
    .B(_1391_));
 sg13g2_inv_1 _5461_ (.Y(_1394_),
    .A(_1392_));
 sg13g2_nor3_2 _5462_ (.A(_1354_),
    .B(_1380_),
    .C(_1381_),
    .Y(_1395_));
 sg13g2_mux2_2 _5463_ (.A0(_1381_),
    .A1(_1384_),
    .S(_1354_),
    .X(_1396_));
 sg13g2_nand2b_2 _5464_ (.Y(_1397_),
    .B(_1385_),
    .A_N(_1395_));
 sg13g2_nor2_1 _5465_ (.A(_1378_),
    .B(_1383_),
    .Y(_1398_));
 sg13g2_or2_1 _5466_ (.X(_1399_),
    .B(_1387_),
    .A(_1375_));
 sg13g2_a21oi_2 _5467_ (.B1(_1398_),
    .Y(_1400_),
    .A2(_1399_),
    .A1(_1389_));
 sg13g2_a221oi_1 _5468_ (.B2(_1389_),
    .C1(_1398_),
    .B1(_1399_),
    .A1(_1390_),
    .Y(_1401_),
    .A2(_1391_));
 sg13g2_nand2_2 _5469_ (.Y(_1402_),
    .A(_1392_),
    .B(_1400_));
 sg13g2_nor2_1 _5470_ (.A(_1397_),
    .B(_1402_),
    .Y(_1403_));
 sg13g2_nand2_2 _5471_ (.Y(_1405_),
    .A(_1396_),
    .B(_1401_));
 sg13g2_a21oi_1 _5472_ (.A1(_1362_),
    .A2(_1370_),
    .Y(_1406_),
    .B1(_1381_));
 sg13g2_xor2_1 _5473_ (.B(_1406_),
    .A(_1374_),
    .X(_1407_));
 sg13g2_nand3_1 _5474_ (.B(_0375_),
    .C(_1383_),
    .A(\hvsync_gen.hpos[1] ),
    .Y(_1408_));
 sg13g2_o21ai_1 _5475_ (.B1(_1367_),
    .Y(_1409_),
    .A1(_0376_),
    .A2(_1381_));
 sg13g2_nand3_1 _5476_ (.B(_1368_),
    .C(_1383_),
    .A(_1366_),
    .Y(_1410_));
 sg13g2_a21o_1 _5477_ (.A2(_1383_),
    .A1(_1368_),
    .B1(_1366_),
    .X(_1411_));
 sg13g2_and2_1 _5478_ (.A(_1410_),
    .B(_1411_),
    .X(_1412_));
 sg13g2_a22oi_1 _5479_ (.Y(_1413_),
    .B1(_1410_),
    .B2(_1411_),
    .A2(_1409_),
    .A1(_1408_));
 sg13g2_nand2_1 _5480_ (.Y(_1414_),
    .A(_1369_),
    .B(_1383_));
 sg13g2_xor2_1 _5481_ (.B(_1414_),
    .A(_1364_),
    .X(_1416_));
 sg13g2_inv_1 _5482_ (.Y(_1417_),
    .A(_1416_));
 sg13g2_nor2_1 _5483_ (.A(_1370_),
    .B(_1381_),
    .Y(_1418_));
 sg13g2_xor2_1 _5484_ (.B(_1418_),
    .A(_1362_),
    .X(_1419_));
 sg13g2_o21ai_1 _5485_ (.B1(_1419_),
    .Y(_1420_),
    .A1(_1413_),
    .A2(_1416_));
 sg13g2_a21oi_2 _5486_ (.B1(_1405_),
    .Y(_1421_),
    .A2(_1420_),
    .A1(_1407_));
 sg13g2_nor3_2 _5487_ (.A(_1394_),
    .B(_1395_),
    .C(_1421_),
    .Y(_1422_));
 sg13g2_or3_2 _5488_ (.A(_1394_),
    .B(_1395_),
    .C(_1421_),
    .X(_1423_));
 sg13g2_nor2_1 _5489_ (.A(_1397_),
    .B(_1401_),
    .Y(_1424_));
 sg13g2_nand2_2 _5490_ (.Y(_1425_),
    .A(_1396_),
    .B(_1402_));
 sg13g2_a21oi_2 _5491_ (.B1(_1425_),
    .Y(_1427_),
    .A2(_1423_),
    .A1(_1385_));
 sg13g2_nor2b_1 _5492_ (.A(_1405_),
    .B_N(_1407_),
    .Y(_1428_));
 sg13g2_nand2_2 _5493_ (.Y(_1429_),
    .A(_1403_),
    .B(_1407_));
 sg13g2_nand2_1 _5494_ (.Y(_1430_),
    .A(_1386_),
    .B(_1394_));
 sg13g2_a21oi_1 _5495_ (.A1(_1385_),
    .A2(_1423_),
    .Y(_1431_),
    .B1(_1407_));
 sg13g2_nor3_1 _5496_ (.A(_1386_),
    .B(_1400_),
    .C(_1422_),
    .Y(_1432_));
 sg13g2_or2_1 _5497_ (.X(_1433_),
    .B(_1419_),
    .A(_1405_));
 sg13g2_o21ai_1 _5498_ (.B1(_1396_),
    .Y(_1434_),
    .A1(_1431_),
    .A2(_1432_));
 sg13g2_and3_1 _5499_ (.X(_1435_),
    .A(_1430_),
    .B(_1433_),
    .C(_1434_));
 sg13g2_nand3_1 _5500_ (.B(_1433_),
    .C(_1434_),
    .A(_1430_),
    .Y(_1436_));
 sg13g2_a21o_1 _5501_ (.A2(_1409_),
    .A1(_1408_),
    .B1(_1405_),
    .X(_1438_));
 sg13g2_a21oi_1 _5502_ (.A1(_1385_),
    .A2(_1423_),
    .Y(_1439_),
    .B1(_1419_));
 sg13g2_nor3_1 _5503_ (.A(_1386_),
    .B(_1407_),
    .C(_1422_),
    .Y(_1440_));
 sg13g2_o21ai_1 _5504_ (.B1(_1405_),
    .Y(_1441_),
    .A1(_1386_),
    .A2(_1422_));
 sg13g2_nand2_1 _5505_ (.Y(_1442_),
    .A(_1407_),
    .B(_1419_));
 sg13g2_nor2_1 _5506_ (.A(_1402_),
    .B(_1442_),
    .Y(_1443_));
 sg13g2_o21ai_1 _5507_ (.B1(_1412_),
    .Y(_1444_),
    .A1(_1402_),
    .A2(_1442_));
 sg13g2_a221oi_1 _5508_ (.B2(_1385_),
    .C1(_1444_),
    .B1(_1423_),
    .A1(_1396_),
    .Y(_1445_),
    .A2(_1401_));
 sg13g2_nor4_1 _5509_ (.A(_1386_),
    .B(_1401_),
    .C(_1417_),
    .D(_1422_),
    .Y(_1446_));
 sg13g2_o21ai_1 _5510_ (.B1(_1396_),
    .Y(_1447_),
    .A1(_1445_),
    .A2(_1446_));
 sg13g2_o21ai_1 _5511_ (.B1(_1397_),
    .Y(_1449_),
    .A1(_1439_),
    .A2(_1440_));
 sg13g2_nand3_1 _5512_ (.B(_1447_),
    .C(_1449_),
    .A(_1438_),
    .Y(_1450_));
 sg13g2_inv_1 _5513_ (.Y(_1451_),
    .A(_1450_));
 sg13g2_nand2_1 _5514_ (.Y(_1452_),
    .A(_1436_),
    .B(_1450_));
 sg13g2_nor2b_1 _5515_ (.A(_1405_),
    .B_N(_1412_),
    .Y(_1453_));
 sg13g2_nor2_1 _5516_ (.A(_1412_),
    .B(_1416_),
    .Y(_1454_));
 sg13g2_a21o_1 _5517_ (.A2(_1454_),
    .A1(_1443_),
    .B1(_1397_),
    .X(_1455_));
 sg13g2_inv_1 _5518_ (.Y(_1456_),
    .A(_1455_));
 sg13g2_or3_1 _5519_ (.A(_1431_),
    .B(_1432_),
    .C(_1456_),
    .X(_1457_));
 sg13g2_nand2_1 _5520_ (.Y(_1458_),
    .A(_1394_),
    .B(_1396_));
 sg13g2_inv_1 _5521_ (.Y(_1460_),
    .A(_1458_));
 sg13g2_a221oi_1 _5522_ (.B2(_1419_),
    .C1(net500),
    .B1(_1460_),
    .A1(_1417_),
    .Y(_1461_),
    .A2(_1427_));
 sg13g2_a21oi_1 _5523_ (.A1(_1457_),
    .A2(_1461_),
    .Y(_1462_),
    .B1(_1453_));
 sg13g2_a21o_2 _5524_ (.A2(_1461_),
    .A1(_1457_),
    .B1(_1453_),
    .X(_1463_));
 sg13g2_nand2_1 _5525_ (.Y(_1464_),
    .A(_1429_),
    .B(_1463_));
 sg13g2_nor2_2 _5526_ (.A(_1435_),
    .B(_1462_),
    .Y(_1465_));
 sg13g2_nand2_2 _5527_ (.Y(_1466_),
    .A(_1429_),
    .B(_1450_));
 sg13g2_nor2_1 _5528_ (.A(_1452_),
    .B(_1464_),
    .Y(_1467_));
 sg13g2_o21ai_1 _5529_ (.B1(_1396_),
    .Y(_1468_),
    .A1(_1439_),
    .A2(_1440_));
 sg13g2_or3_1 _5530_ (.A(_1395_),
    .B(_1400_),
    .C(_1421_),
    .X(_1469_));
 sg13g2_o21ai_1 _5531_ (.B1(_1469_),
    .Y(_1471_),
    .A1(_1386_),
    .A2(_1392_));
 sg13g2_a21oi_1 _5532_ (.A1(_1455_),
    .A2(_1471_),
    .Y(_1472_),
    .B1(net500));
 sg13g2_a22oi_1 _5533_ (.Y(_1473_),
    .B1(_1468_),
    .B2(_1472_),
    .A2(_1417_),
    .A1(net500));
 sg13g2_and2_1 _5534_ (.A(_1450_),
    .B(net479),
    .X(_1474_));
 sg13g2_nand4_1 _5535_ (.B(_1450_),
    .C(_1463_),
    .A(_1436_),
    .Y(_1475_),
    .D(net479));
 sg13g2_nand2_2 _5536_ (.Y(_1476_),
    .A(_0376_),
    .B(net500));
 sg13g2_nand2_1 _5537_ (.Y(_1477_),
    .A(_1429_),
    .B(_1476_));
 sg13g2_a22oi_1 _5538_ (.Y(_1478_),
    .B1(_1463_),
    .B2(net479),
    .A2(_1450_),
    .A1(_1436_));
 sg13g2_a21oi_1 _5539_ (.A1(_1465_),
    .A2(_1474_),
    .Y(_1479_),
    .B1(_1478_));
 sg13g2_o21ai_1 _5540_ (.B1(_1475_),
    .Y(_1480_),
    .A1(_1477_),
    .A2(_1478_));
 sg13g2_inv_1 _5541_ (.Y(_1482_),
    .A(_1480_));
 sg13g2_xnor2_1 _5542_ (.Y(_1483_),
    .A(_1465_),
    .B(_1466_));
 sg13g2_xnor2_1 _5543_ (.Y(_1484_),
    .A(_1480_),
    .B(_1483_));
 sg13g2_xnor2_1 _5544_ (.Y(_1485_),
    .A(_1465_),
    .B(net479));
 sg13g2_nor2_1 _5545_ (.A(_1466_),
    .B(_1485_),
    .Y(_1486_));
 sg13g2_xnor2_1 _5546_ (.Y(_1487_),
    .A(_1466_),
    .B(_1485_));
 sg13g2_or4_1 _5547_ (.A(_1452_),
    .B(_1464_),
    .C(_1484_),
    .D(_1487_),
    .X(_1488_));
 sg13g2_a21oi_1 _5548_ (.A1(_1465_),
    .A2(net479),
    .Y(_1489_),
    .B1(_1486_));
 sg13g2_a21oi_1 _5549_ (.A1(_1480_),
    .A2(_1483_),
    .Y(_1490_),
    .B1(_1467_));
 sg13g2_o21ai_1 _5550_ (.B1(_1490_),
    .Y(_1491_),
    .A1(_1484_),
    .A2(_1487_));
 sg13g2_nand2_1 _5551_ (.Y(_1493_),
    .A(_1488_),
    .B(_1491_));
 sg13g2_or2_1 _5552_ (.X(_1494_),
    .B(_1493_),
    .A(_1489_));
 sg13g2_or2_1 _5553_ (.X(_1495_),
    .B(net480),
    .A(_1435_));
 sg13g2_xnor2_1 _5554_ (.Y(_1496_),
    .A(_1464_),
    .B(_1495_));
 sg13g2_a21o_1 _5555_ (.A2(_1494_),
    .A1(_1488_),
    .B1(_1496_),
    .X(_1497_));
 sg13g2_xnor2_1 _5556_ (.Y(_1498_),
    .A(_1477_),
    .B(_1479_));
 sg13g2_inv_1 _5557_ (.Y(_1499_),
    .A(_1498_));
 sg13g2_mux2_1 _5558_ (.A0(_1482_),
    .A1(_1499_),
    .S(net480),
    .X(_1500_));
 sg13g2_xnor2_1 _5559_ (.Y(_1501_),
    .A(_1489_),
    .B(_1493_));
 sg13g2_nor2_1 _5560_ (.A(_1500_),
    .B(_1501_),
    .Y(_1502_));
 sg13g2_nand2_1 _5561_ (.Y(_1504_),
    .A(net480),
    .B(_1476_));
 sg13g2_nor2_1 _5562_ (.A(_1452_),
    .B(_1504_),
    .Y(_1505_));
 sg13g2_a21o_1 _5563_ (.A2(_1476_),
    .A1(_1436_),
    .B1(_1474_),
    .X(_1506_));
 sg13g2_nor2_1 _5564_ (.A(_1451_),
    .B(_1462_),
    .Y(_1507_));
 sg13g2_a21oi_1 _5565_ (.A1(_1506_),
    .A2(_1507_),
    .Y(_1508_),
    .B1(_1505_));
 sg13g2_xor2_1 _5566_ (.B(_1498_),
    .A(net480),
    .X(_1509_));
 sg13g2_nor2b_1 _5567_ (.A(_1508_),
    .B_N(_1509_),
    .Y(_1510_));
 sg13g2_nand3_1 _5568_ (.B(net480),
    .C(_1476_),
    .A(_1463_),
    .Y(_1511_));
 sg13g2_nand2b_1 _5569_ (.Y(_1512_),
    .B(_1506_),
    .A_N(_1505_));
 sg13g2_xnor2_1 _5570_ (.Y(_1513_),
    .A(_1507_),
    .B(_1512_));
 sg13g2_nand2b_1 _5571_ (.Y(_1515_),
    .B(_1513_),
    .A_N(_1511_));
 sg13g2_inv_1 _5572_ (.Y(_1516_),
    .A(_1515_));
 sg13g2_xnor2_1 _5573_ (.Y(_1517_),
    .A(_1508_),
    .B(_1509_));
 sg13g2_a21oi_1 _5574_ (.A1(_1516_),
    .A2(_1517_),
    .Y(_1518_),
    .B1(_1510_));
 sg13g2_xnor2_1 _5575_ (.Y(_1519_),
    .A(_1500_),
    .B(_1501_));
 sg13g2_nor2_1 _5576_ (.A(_1518_),
    .B(_1519_),
    .Y(_1520_));
 sg13g2_nor2_1 _5577_ (.A(_1502_),
    .B(_1520_),
    .Y(_1521_));
 sg13g2_nand3_1 _5578_ (.B(_1494_),
    .C(_1496_),
    .A(_1488_),
    .Y(_1522_));
 sg13g2_nand2_1 _5579_ (.Y(_1523_),
    .A(_1497_),
    .B(_1522_));
 sg13g2_o21ai_1 _5580_ (.B1(_1497_),
    .Y(_1524_),
    .A1(_1521_),
    .A2(_1523_));
 sg13g2_a21oi_1 _5581_ (.A1(_1436_),
    .A2(net479),
    .Y(_1526_),
    .B1(_1429_));
 sg13g2_nand3_1 _5582_ (.B(_1436_),
    .C(net479),
    .A(_1429_),
    .Y(_1527_));
 sg13g2_o21ai_1 _5583_ (.B1(_1527_),
    .Y(_1528_),
    .A1(_1465_),
    .A2(net479));
 sg13g2_nor2_1 _5584_ (.A(_1526_),
    .B(_1528_),
    .Y(_1529_));
 sg13g2_nand2_1 _5585_ (.Y(_1530_),
    .A(_1524_),
    .B(_1529_));
 sg13g2_a21oi_1 _5586_ (.A1(_1435_),
    .A2(_1530_),
    .Y(_1531_),
    .B1(_1428_));
 sg13g2_a21o_1 _5587_ (.A2(_1530_),
    .A1(_1435_),
    .B1(_1428_),
    .X(_1532_));
 sg13g2_xnor2_1 _5588_ (.Y(_1533_),
    .A(_1511_),
    .B(_1513_));
 sg13g2_xor2_1 _5589_ (.B(_1519_),
    .A(_1518_),
    .X(_1534_));
 sg13g2_nor2b_1 _5590_ (.A(_1441_),
    .B_N(_1534_),
    .Y(_1535_));
 sg13g2_a21oi_1 _5591_ (.A1(_1441_),
    .A2(_1533_),
    .Y(_1537_),
    .B1(_1535_));
 sg13g2_nor2_1 _5592_ (.A(_1396_),
    .B(_1537_),
    .Y(_1538_));
 sg13g2_xor2_1 _5593_ (.B(_1529_),
    .A(_1524_),
    .X(_1539_));
 sg13g2_a221oi_1 _5594_ (.B2(_1460_),
    .C1(_1538_),
    .B1(_1539_),
    .A1(_1427_),
    .Y(_1540_),
    .A2(_1531_));
 sg13g2_nor2_2 _5595_ (.A(_2491_),
    .B(_1540_),
    .Y(_1541_));
 sg13g2_xnor2_1 _5596_ (.Y(_1542_),
    .A(_2491_),
    .B(_1540_));
 sg13g2_and3_1 _5597_ (.X(_1543_),
    .A(_1429_),
    .B(_1495_),
    .C(_1530_));
 sg13g2_xor2_1 _5598_ (.B(_1523_),
    .A(_1521_),
    .X(_1544_));
 sg13g2_xnor2_1 _5599_ (.Y(_1545_),
    .A(_1515_),
    .B(_1517_));
 sg13g2_xnor2_1 _5600_ (.Y(_1546_),
    .A(_1463_),
    .B(_1504_));
 sg13g2_o21ai_1 _5601_ (.B1(_1546_),
    .Y(_1548_),
    .A1(_1451_),
    .A2(_1476_));
 sg13g2_nor2_1 _5602_ (.A(_1441_),
    .B(_1545_),
    .Y(_1549_));
 sg13g2_a21oi_1 _5603_ (.A1(_1441_),
    .A2(_1548_),
    .Y(_1550_),
    .B1(_1549_));
 sg13g2_and2_1 _5604_ (.A(_1397_),
    .B(_1550_),
    .X(_1551_));
 sg13g2_a221oi_1 _5605_ (.B2(_1460_),
    .C1(_1551_),
    .B1(_1544_),
    .A1(_1427_),
    .Y(_1552_),
    .A2(_1543_));
 sg13g2_inv_1 _5606_ (.Y(_1553_),
    .A(_1552_));
 sg13g2_nor2_1 _5607_ (.A(_2828_),
    .B(_1552_),
    .Y(_1554_));
 sg13g2_xnor2_1 _5608_ (.Y(_1555_),
    .A(_2828_),
    .B(_1552_));
 sg13g2_inv_1 _5609_ (.Y(_1556_),
    .A(_1555_));
 sg13g2_mux2_1 _5610_ (.A0(_1539_),
    .A1(_1534_),
    .S(_1441_),
    .X(_1557_));
 sg13g2_nor2_1 _5611_ (.A(_1425_),
    .B(_1557_),
    .Y(_1559_));
 sg13g2_nor2b_1 _5612_ (.A(_1441_),
    .B_N(_1533_),
    .Y(_1560_));
 sg13g2_xnor2_1 _5613_ (.Y(_1561_),
    .A(_1450_),
    .B(_1463_));
 sg13g2_nor2b_1 _5614_ (.A(_1561_),
    .B_N(_1441_),
    .Y(_1562_));
 sg13g2_nor2_1 _5615_ (.A(_1560_),
    .B(_1562_),
    .Y(_1563_));
 sg13g2_a221oi_1 _5616_ (.B2(_1397_),
    .C1(_1559_),
    .B1(_1563_),
    .A1(net500),
    .Y(_1564_),
    .A2(_1532_));
 sg13g2_inv_1 _5617_ (.Y(_1565_),
    .A(_1564_));
 sg13g2_nand2_1 _5618_ (.Y(_1566_),
    .A(_2847_),
    .B(_1564_));
 sg13g2_xnor2_1 _5619_ (.Y(_1567_),
    .A(_2847_),
    .B(_1564_));
 sg13g2_inv_1 _5620_ (.Y(_1568_),
    .A(_1567_));
 sg13g2_mux2_1 _5621_ (.A0(_1544_),
    .A1(_1545_),
    .S(_1441_),
    .X(_1570_));
 sg13g2_inv_1 _5622_ (.Y(_1571_),
    .A(_1570_));
 sg13g2_a22oi_1 _5623_ (.Y(_1572_),
    .B1(_1546_),
    .B2(_1386_),
    .A2(_1543_),
    .A1(net500));
 sg13g2_o21ai_1 _5624_ (.B1(_1572_),
    .Y(_1573_),
    .A1(_1425_),
    .A2(_1571_));
 sg13g2_inv_1 _5625_ (.Y(_1574_),
    .A(_1573_));
 sg13g2_and2_1 _5626_ (.A(_2860_),
    .B(_1573_),
    .X(_1575_));
 sg13g2_xor2_1 _5627_ (.B(_1573_),
    .A(_2860_),
    .X(_1576_));
 sg13g2_nor2_1 _5628_ (.A(_1425_),
    .B(_1537_),
    .Y(_1577_));
 sg13g2_a21oi_1 _5629_ (.A1(net500),
    .A2(_1539_),
    .Y(_1578_),
    .B1(_1577_));
 sg13g2_o21ai_1 _5630_ (.B1(_1578_),
    .Y(_1579_),
    .A1(_1385_),
    .A2(_1561_));
 sg13g2_nand2_1 _5631_ (.Y(_1581_),
    .A(_2875_),
    .B(_1579_));
 sg13g2_xnor2_1 _5632_ (.Y(_1582_),
    .A(_2875_),
    .B(_1579_));
 sg13g2_a221oi_1 _5633_ (.B2(_1424_),
    .C1(_1395_),
    .B1(_1550_),
    .A1(net500),
    .Y(_1583_),
    .A2(_1544_));
 sg13g2_inv_1 _5634_ (.Y(_1584_),
    .A(_1583_));
 sg13g2_nand3b_1 _5635_ (.B(_1584_),
    .C(net474),
    .Y(_1585_),
    .A_N(_1582_));
 sg13g2_nand2_1 _5636_ (.Y(_1586_),
    .A(_1581_),
    .B(_1585_));
 sg13g2_a21oi_1 _5637_ (.A1(_1576_),
    .A2(_1586_),
    .Y(_1587_),
    .B1(_1575_));
 sg13g2_o21ai_1 _5638_ (.B1(_1566_),
    .Y(_1588_),
    .A1(_1567_),
    .A2(_1587_));
 sg13g2_a21oi_1 _5639_ (.A1(_1556_),
    .A2(_1588_),
    .Y(_1589_),
    .B1(_1554_));
 sg13g2_xnor2_1 _5640_ (.Y(_1590_),
    .A(_1542_),
    .B(_1589_));
 sg13g2_xnor2_1 _5641_ (.Y(_1592_),
    .A(_1556_),
    .B(_1588_));
 sg13g2_xnor2_1 _5642_ (.Y(_1593_),
    .A(_1567_),
    .B(_1587_));
 sg13g2_xor2_1 _5643_ (.B(_1586_),
    .A(_1576_),
    .X(_1594_));
 sg13g2_a22oi_1 _5644_ (.Y(_1595_),
    .B1(_1570_),
    .B2(_1397_),
    .A2(_1543_),
    .A1(_1460_));
 sg13g2_nand2_1 _5645_ (.Y(_1596_),
    .A(_2910_),
    .B(_1595_));
 sg13g2_xnor2_1 _5646_ (.Y(_1597_),
    .A(_2910_),
    .B(_1595_));
 sg13g2_nor2_1 _5647_ (.A(_1458_),
    .B(_1532_),
    .Y(_1598_));
 sg13g2_a21oi_2 _5648_ (.B1(_1598_),
    .Y(_1599_),
    .A2(_1557_),
    .A1(_1397_));
 sg13g2_nor2b_1 _5649_ (.A(_1599_),
    .B_N(_1595_),
    .Y(_1600_));
 sg13g2_nand2_1 _5650_ (.Y(_1601_),
    .A(net569),
    .B(_0162_));
 sg13g2_nand3_1 _5651_ (.B(net571),
    .C(_0162_),
    .A(net569),
    .Y(_1603_));
 sg13g2_nor3_1 _5652_ (.A(net563),
    .B(_3147_),
    .C(_0184_),
    .Y(_1604_));
 sg13g2_nor3_1 _5653_ (.A(net565),
    .B(net571),
    .C(_1601_),
    .Y(_1605_));
 sg13g2_nand3_1 _5654_ (.B(_0056_),
    .C(_1605_),
    .A(_2923_),
    .Y(_1606_));
 sg13g2_nand3_1 _5655_ (.B(_1604_),
    .C(_1606_),
    .A(_1603_),
    .Y(_1607_));
 sg13g2_a21oi_1 _5656_ (.A1(_1596_),
    .A2(_1599_),
    .Y(_1608_),
    .B1(_1607_));
 sg13g2_xor2_1 _5657_ (.B(_1583_),
    .A(net474),
    .X(_1609_));
 sg13g2_o21ai_1 _5658_ (.B1(_1608_),
    .Y(_1610_),
    .A1(_1541_),
    .A2(_1597_));
 sg13g2_o21ai_1 _5659_ (.B1(_1597_),
    .Y(_1611_),
    .A1(_1541_),
    .A2(_1600_));
 sg13g2_o21ai_1 _5660_ (.B1(_1611_),
    .Y(_1612_),
    .A1(_1582_),
    .A2(_1609_));
 sg13g2_nor3_1 _5661_ (.A(_1594_),
    .B(_1610_),
    .C(_1612_),
    .Y(_1614_));
 sg13g2_nand3_1 _5662_ (.B(_1593_),
    .C(_1614_),
    .A(_1592_),
    .Y(_1615_));
 sg13g2_or2_1 _5663_ (.X(_1616_),
    .B(_1615_),
    .A(_1590_));
 sg13g2_xnor2_1 _5664_ (.Y(_1617_),
    .A(_1555_),
    .B(_1595_));
 sg13g2_nand2_1 _5665_ (.Y(_1618_),
    .A(_1540_),
    .B(_1568_));
 sg13g2_and2_1 _5666_ (.A(_1566_),
    .B(_1618_),
    .X(_1619_));
 sg13g2_nor2b_1 _5667_ (.A(_1619_),
    .B_N(_1617_),
    .Y(_1620_));
 sg13g2_xnor2_1 _5668_ (.Y(_1621_),
    .A(_1617_),
    .B(_1619_));
 sg13g2_a21oi_1 _5669_ (.A1(_1552_),
    .A2(_1576_),
    .Y(_1622_),
    .B1(_1575_));
 sg13g2_xor2_1 _5670_ (.B(_1567_),
    .A(_1540_),
    .X(_1623_));
 sg13g2_nand2_1 _5671_ (.Y(_1625_),
    .A(_1622_),
    .B(_1623_));
 sg13g2_nor2_2 _5672_ (.A(net474),
    .B(_1574_),
    .Y(_1626_));
 sg13g2_or2_1 _5673_ (.X(_1627_),
    .B(_1582_),
    .A(_1564_));
 sg13g2_xnor2_1 _5674_ (.Y(_1628_),
    .A(_1564_),
    .B(_1582_));
 sg13g2_xnor2_1 _5675_ (.Y(_1629_),
    .A(net474),
    .B(_1573_));
 sg13g2_nor2_1 _5676_ (.A(_1583_),
    .B(_1629_),
    .Y(_1630_));
 sg13g2_xor2_1 _5677_ (.B(_1628_),
    .A(_1626_),
    .X(_1631_));
 sg13g2_nand2_1 _5678_ (.Y(_1632_),
    .A(_1630_),
    .B(_1631_));
 sg13g2_o21ai_1 _5679_ (.B1(_1632_),
    .Y(_1633_),
    .A1(_1626_),
    .A2(_1628_));
 sg13g2_xnor2_1 _5680_ (.Y(_1634_),
    .A(_1552_),
    .B(_1576_));
 sg13g2_a21oi_1 _5681_ (.A1(_1581_),
    .A2(_1627_),
    .Y(_1636_),
    .B1(_1634_));
 sg13g2_nor2_1 _5682_ (.A(_1622_),
    .B(_1623_),
    .Y(_1637_));
 sg13g2_or3_1 _5683_ (.A(_1633_),
    .B(_1636_),
    .C(_1637_),
    .X(_1638_));
 sg13g2_a21o_1 _5684_ (.A2(_1638_),
    .A1(_1625_),
    .B1(_1621_),
    .X(_1639_));
 sg13g2_nand2b_1 _5685_ (.Y(_1640_),
    .B(_1599_),
    .A_N(_1542_));
 sg13g2_nand2b_1 _5686_ (.Y(_1641_),
    .B(_1640_),
    .A_N(_1541_));
 sg13g2_xor2_1 _5687_ (.B(_1641_),
    .A(_1597_),
    .X(_1642_));
 sg13g2_xnor2_1 _5688_ (.Y(_1643_),
    .A(_1542_),
    .B(_1599_));
 sg13g2_a21o_1 _5689_ (.A2(_1595_),
    .A1(_1556_),
    .B1(_1554_),
    .X(_1644_));
 sg13g2_and2_1 _5690_ (.A(_1643_),
    .B(_1644_),
    .X(_1645_));
 sg13g2_nor2_1 _5691_ (.A(_1620_),
    .B(_1645_),
    .Y(_1647_));
 sg13g2_and3_1 _5692_ (.X(_1648_),
    .A(_1581_),
    .B(_1627_),
    .C(_1634_));
 sg13g2_o21ai_1 _5693_ (.B1(_1633_),
    .Y(_1649_),
    .A1(_1636_),
    .A2(_1648_));
 sg13g2_o21ai_1 _5694_ (.B1(_1649_),
    .Y(_1650_),
    .A1(_1642_),
    .A2(_1647_));
 sg13g2_nor2_1 _5695_ (.A(_1643_),
    .B(_1644_),
    .Y(_1651_));
 sg13g2_o21ai_1 _5696_ (.B1(_1651_),
    .Y(_1652_),
    .A1(_1541_),
    .A2(_1599_));
 sg13g2_or2_1 _5697_ (.X(_1653_),
    .B(_1652_),
    .A(_1642_));
 sg13g2_a221oi_1 _5698_ (.B2(_1653_),
    .C1(_1650_),
    .B1(_1647_),
    .A1(_1621_),
    .Y(_1654_),
    .A2(_1625_));
 sg13g2_nor2_1 _5699_ (.A(_1621_),
    .B(_1637_),
    .Y(_1655_));
 sg13g2_or2_1 _5700_ (.X(_1656_),
    .B(_1655_),
    .A(_1648_));
 sg13g2_or2_1 _5701_ (.X(_1658_),
    .B(_1631_),
    .A(_1630_));
 sg13g2_o21ai_1 _5702_ (.B1(_1620_),
    .Y(_1659_),
    .A1(_1645_),
    .A2(_1651_));
 sg13g2_nor3_1 _5703_ (.A(_3037_),
    .B(_3256_),
    .C(_1601_),
    .Y(_1660_));
 sg13g2_or2_1 _5704_ (.X(_1661_),
    .B(net574),
    .A(net565));
 sg13g2_nor4_1 _5705_ (.A(net565),
    .B(net574),
    .C(_0700_),
    .D(_1603_),
    .Y(_1662_));
 sg13g2_nor4_2 _5706_ (.A(_0184_),
    .B(_2924_),
    .C(_1660_),
    .Y(_1663_),
    .D(_1662_));
 sg13g2_xnor2_1 _5707_ (.Y(_1664_),
    .A(_1596_),
    .B(_1599_));
 sg13g2_o21ai_1 _5708_ (.B1(_1664_),
    .Y(_1665_),
    .A1(_1597_),
    .A2(_1641_));
 sg13g2_nand3_1 _5709_ (.B(_1663_),
    .C(_1665_),
    .A(_1659_),
    .Y(_1666_));
 sg13g2_a21oi_1 _5710_ (.A1(_1632_),
    .A2(_1658_),
    .Y(_1667_),
    .B1(_1666_));
 sg13g2_nand4_1 _5711_ (.B(_1654_),
    .C(_1656_),
    .A(_1639_),
    .Y(_1669_),
    .D(_1667_));
 sg13g2_xor2_1 _5712_ (.B(_2912_),
    .A(_2849_),
    .X(_1670_));
 sg13g2_nand2_1 _5713_ (.Y(_1671_),
    .A(net471),
    .B(_2862_));
 sg13g2_nand2_1 _5714_ (.Y(_1672_),
    .A(_2861_),
    .B(_1671_));
 sg13g2_nand2_1 _5715_ (.Y(_1673_),
    .A(_1670_),
    .B(_1672_));
 sg13g2_o21ai_1 _5716_ (.B1(_2848_),
    .Y(_1674_),
    .A1(_2849_),
    .A2(_2912_));
 sg13g2_nand2_1 _5717_ (.Y(_1675_),
    .A(_2831_),
    .B(_1674_));
 sg13g2_xnor2_1 _5718_ (.Y(_1676_),
    .A(_2831_),
    .B(_1674_));
 sg13g2_xnor2_1 _5719_ (.Y(_1677_),
    .A(_1673_),
    .B(_1676_));
 sg13g2_xnor2_1 _5720_ (.Y(_1678_),
    .A(_2830_),
    .B(_2917_));
 sg13g2_nor2_1 _5721_ (.A(net565),
    .B(_1325_),
    .Y(_1680_));
 sg13g2_nor3_1 _5722_ (.A(_2993_),
    .B(_0348_),
    .C(_1680_),
    .Y(_1681_));
 sg13g2_nor3_1 _5723_ (.A(_0162_),
    .B(_2924_),
    .C(_1681_),
    .Y(_1682_));
 sg13g2_xnor2_1 _5724_ (.Y(_1683_),
    .A(_1675_),
    .B(_1678_));
 sg13g2_xnor2_1 _5725_ (.Y(_1684_),
    .A(_1670_),
    .B(_1672_));
 sg13g2_xnor2_1 _5726_ (.Y(_1685_),
    .A(net471),
    .B(_2862_));
 sg13g2_nor2_1 _5727_ (.A(net468),
    .B(_2878_),
    .Y(_1686_));
 sg13g2_nor2_1 _5728_ (.A(_2876_),
    .B(_1686_),
    .Y(_1687_));
 sg13g2_or2_1 _5729_ (.X(_1688_),
    .B(_1687_),
    .A(_1685_));
 sg13g2_and2_1 _5730_ (.A(_1684_),
    .B(_1688_),
    .X(_1689_));
 sg13g2_nor4_1 _5731_ (.A(_1677_),
    .B(_1682_),
    .C(_1683_),
    .D(_1689_),
    .Y(_1691_));
 sg13g2_a21oi_1 _5732_ (.A1(_1685_),
    .A2(_1687_),
    .Y(_1692_),
    .B1(_1684_));
 sg13g2_xnor2_1 _5733_ (.Y(_1693_),
    .A(_2840_),
    .B(_2878_));
 sg13g2_nor2_1 _5734_ (.A(_2855_),
    .B(net472),
    .Y(_1694_));
 sg13g2_a21o_1 _5735_ (.A2(_1694_),
    .A1(_1693_),
    .B1(_1692_),
    .X(_1695_));
 sg13g2_and3_1 _5736_ (.X(_1696_),
    .A(_2855_),
    .B(net472),
    .C(_1688_));
 sg13g2_nand2b_1 _5737_ (.Y(_1697_),
    .B(_1696_),
    .A_N(_1693_));
 sg13g2_a21oi_1 _5738_ (.A1(net472),
    .A2(_2885_),
    .Y(_1698_),
    .B1(_2855_));
 sg13g2_or4_1 _5739_ (.A(_2886_),
    .B(_1692_),
    .C(_1693_),
    .D(_1698_),
    .X(_1699_));
 sg13g2_a22oi_1 _5740_ (.Y(_1700_),
    .B1(_1697_),
    .B2(_1692_),
    .A2(_1695_),
    .A1(_2884_));
 sg13g2_nand3_1 _5741_ (.B(_1699_),
    .C(_1700_),
    .A(_1691_),
    .Y(_1702_));
 sg13g2_nor2_2 _5742_ (.A(_0097_),
    .B(_2546_),
    .Y(_1703_));
 sg13g2_o21ai_1 _5743_ (.B1(_2586_),
    .Y(_1704_),
    .A1(_0097_),
    .A2(net534));
 sg13g2_xnor2_1 _5744_ (.Y(_1705_),
    .A(net584),
    .B(_1704_));
 sg13g2_nor2_1 _5745_ (.A(net536),
    .B(net532),
    .Y(_1706_));
 sg13g2_nor3_1 _5746_ (.A(_0005_),
    .B(net536),
    .C(_2938_),
    .Y(_1707_));
 sg13g2_o21ai_1 _5747_ (.B1(net550),
    .Y(_1708_),
    .A1(net564),
    .A2(_1707_));
 sg13g2_a21oi_1 _5748_ (.A1(net564),
    .A2(_1707_),
    .Y(_1709_),
    .B1(_1708_));
 sg13g2_a21oi_2 _5749_ (.B1(_1709_),
    .Y(_1710_),
    .A2(_1705_),
    .A1(net541));
 sg13g2_nand3b_1 _5750_ (.B(_2939_),
    .C(_2982_),
    .Y(_1711_),
    .A_N(net536));
 sg13g2_a21oi_1 _5751_ (.A1(_0004_),
    .A2(_1711_),
    .Y(_1713_),
    .B1(net561));
 sg13g2_and3_1 _5752_ (.X(_1714_),
    .A(net561),
    .B(net562),
    .C(_1711_));
 sg13g2_nor3_2 _5753_ (.A(net541),
    .B(_1713_),
    .C(_1714_),
    .Y(_1715_));
 sg13g2_nand2_1 _5754_ (.Y(_1716_),
    .A(net582),
    .B(net538));
 sg13g2_a21o_1 _5755_ (.A2(_1704_),
    .A1(net584),
    .B1(_1716_),
    .X(_1717_));
 sg13g2_nor2_1 _5756_ (.A(net582),
    .B(_3070_),
    .Y(_1718_));
 sg13g2_nand2_1 _5757_ (.Y(_1719_),
    .A(_1704_),
    .B(_1718_));
 sg13g2_o21ai_1 _5758_ (.B1(_1717_),
    .Y(_1720_),
    .A1(net547),
    .A2(_1719_));
 sg13g2_nor2_2 _5759_ (.A(_1715_),
    .B(_1720_),
    .Y(_1721_));
 sg13g2_or2_2 _5760_ (.X(_1722_),
    .B(_1720_),
    .A(_1715_));
 sg13g2_o21ai_1 _5761_ (.B1(_0005_),
    .Y(_1724_),
    .A1(net536),
    .A2(_2938_));
 sg13g2_nand2b_1 _5762_ (.Y(_1725_),
    .B(_1724_),
    .A_N(_1707_));
 sg13g2_nand2_1 _5763_ (.Y(_1726_),
    .A(net550),
    .B(_1725_));
 sg13g2_nor2_1 _5764_ (.A(_3180_),
    .B(_1703_),
    .Y(_1727_));
 sg13g2_xnor2_1 _5765_ (.Y(_1728_),
    .A(_0001_),
    .B(_1727_));
 sg13g2_o21ai_1 _5766_ (.B1(_1726_),
    .Y(_1729_),
    .A1(net550),
    .A2(_1728_));
 sg13g2_o21ai_1 _5767_ (.B1(net554),
    .Y(_1730_),
    .A1(_0271_),
    .A2(_2937_));
 sg13g2_a21oi_2 _5768_ (.B1(_1730_),
    .Y(_1731_),
    .A2(_0887_),
    .A1(_3015_));
 sg13g2_o21ai_1 _5769_ (.B1(net539),
    .Y(_1732_),
    .A1(net592),
    .A2(_2637_));
 sg13g2_a21oi_1 _5770_ (.A1(net592),
    .A2(_2637_),
    .Y(_1733_),
    .B1(_1732_));
 sg13g2_or2_1 _5771_ (.X(_1735_),
    .B(_1733_),
    .A(_1731_));
 sg13g2_nand2_1 _5772_ (.Y(_1736_),
    .A(net578),
    .B(net549));
 sg13g2_o21ai_1 _5773_ (.B1(_1736_),
    .Y(_1737_),
    .A1(net549),
    .A2(_2619_));
 sg13g2_mux2_2 _5774_ (.A0(net607),
    .A1(_0006_),
    .S(net547),
    .X(_1738_));
 sg13g2_nand2_2 _5775_ (.Y(_1739_),
    .A(_1737_),
    .B(_1738_));
 sg13g2_nand2b_1 _5776_ (.Y(_1740_),
    .B(_2535_),
    .A_N(net600));
 sg13g2_a21oi_1 _5777_ (.A1(net600),
    .A2(_2524_),
    .Y(_1741_),
    .B1(net552));
 sg13g2_a22oi_1 _5778_ (.Y(_1742_),
    .B1(_1740_),
    .B2(_1741_),
    .A2(_0777_),
    .A1(net552));
 sg13g2_or2_1 _5779_ (.X(_1743_),
    .B(_1742_),
    .A(_1739_));
 sg13g2_a21oi_1 _5780_ (.A1(_0271_),
    .A2(_0832_),
    .Y(_1744_),
    .B1(net544));
 sg13g2_xnor2_1 _5781_ (.Y(_1746_),
    .A(_3202_),
    .B(_2610_));
 sg13g2_a21oi_2 _5782_ (.B1(_1744_),
    .Y(_1747_),
    .A2(_1746_),
    .A1(net544));
 sg13g2_xnor2_1 _5783_ (.Y(_1748_),
    .A(_3136_),
    .B(net536));
 sg13g2_mux2_1 _5784_ (.A0(_2641_),
    .A1(_1748_),
    .S(net549),
    .X(_1749_));
 sg13g2_nor4_1 _5785_ (.A(_1739_),
    .B(_1742_),
    .C(_1747_),
    .D(_1749_),
    .Y(_1750_));
 sg13g2_nand2_1 _5786_ (.Y(_1751_),
    .A(_1721_),
    .B(_1739_));
 sg13g2_nand2_1 _5787_ (.Y(_1752_),
    .A(_1721_),
    .B(_1743_));
 sg13g2_o21ai_1 _5788_ (.B1(_1721_),
    .Y(_1753_),
    .A1(_1743_),
    .A2(_1747_));
 sg13g2_nor3_2 _5789_ (.A(_1715_),
    .B(_1720_),
    .C(_1750_),
    .Y(_1754_));
 sg13g2_o21ai_1 _5790_ (.B1(_1721_),
    .Y(_1755_),
    .A1(_1735_),
    .A2(_1754_));
 sg13g2_xnor2_1 _5791_ (.Y(_1757_),
    .A(_3169_),
    .B(_1706_));
 sg13g2_xnor2_1 _5792_ (.Y(_1758_),
    .A(net590),
    .B(_1703_));
 sg13g2_nor2_1 _5793_ (.A(net549),
    .B(_1758_),
    .Y(_1759_));
 sg13g2_a21oi_1 _5794_ (.A1(net549),
    .A2(_1757_),
    .Y(_1760_),
    .B1(_1759_));
 sg13g2_nor3_1 _5795_ (.A(_1735_),
    .B(_1754_),
    .C(_1760_),
    .Y(_1761_));
 sg13g2_a21oi_1 _5796_ (.A1(_1729_),
    .A2(_1761_),
    .Y(_1762_),
    .B1(_1722_));
 sg13g2_nor2_1 _5797_ (.A(_1710_),
    .B(_1722_),
    .Y(_1763_));
 sg13g2_mux2_1 _5798_ (.A0(_1722_),
    .A1(_1762_),
    .S(_1710_),
    .X(_1764_));
 sg13g2_or3_1 _5799_ (.A(_1722_),
    .B(_1729_),
    .C(_1761_),
    .X(_1765_));
 sg13g2_o21ai_1 _5800_ (.B1(_1729_),
    .Y(_1766_),
    .A1(_1722_),
    .A2(_1761_));
 sg13g2_nand2_1 _5801_ (.Y(_1768_),
    .A(_1765_),
    .B(_1766_));
 sg13g2_inv_1 _5802_ (.Y(_1769_),
    .A(_1768_));
 sg13g2_xnor2_1 _5803_ (.Y(_1770_),
    .A(_1755_),
    .B(_1760_));
 sg13g2_a21oi_2 _5804_ (.B1(_1770_),
    .Y(_1771_),
    .A2(_1766_),
    .A1(_1765_));
 sg13g2_and2_1 _5805_ (.A(net516),
    .B(_1771_),
    .X(_1772_));
 sg13g2_inv_1 _5806_ (.Y(_1773_),
    .A(net508));
 sg13g2_nor2b_2 _5807_ (.A(_1771_),
    .B_N(net516),
    .Y(_1774_));
 sg13g2_nand2b_2 _5808_ (.Y(_1775_),
    .B(net516),
    .A_N(_1771_));
 sg13g2_xor2_1 _5809_ (.B(_1762_),
    .A(_1710_),
    .X(_1776_));
 sg13g2_a21oi_2 _5810_ (.B1(_1763_),
    .Y(_1777_),
    .A2(_1766_),
    .A1(_1765_));
 sg13g2_a21oi_1 _5811_ (.A1(_1770_),
    .A2(_1777_),
    .Y(_1779_),
    .B1(_1776_));
 sg13g2_a21o_1 _5812_ (.A2(_1777_),
    .A1(_1770_),
    .B1(_1776_),
    .X(_1780_));
 sg13g2_xor2_1 _5813_ (.B(_1753_),
    .A(_1749_),
    .X(_1781_));
 sg13g2_nor2_1 _5814_ (.A(_1722_),
    .B(_1738_),
    .Y(_1782_));
 sg13g2_xnor2_1 _5815_ (.Y(_1783_),
    .A(_1737_),
    .B(_1782_));
 sg13g2_xor2_1 _5816_ (.B(_1782_),
    .A(_1737_),
    .X(_1784_));
 sg13g2_xnor2_1 _5817_ (.Y(_1785_),
    .A(_1742_),
    .B(_1751_));
 sg13g2_inv_1 _5818_ (.Y(_1786_),
    .A(_1785_));
 sg13g2_xor2_1 _5819_ (.B(_1752_),
    .A(_1747_),
    .X(_1787_));
 sg13g2_inv_1 _5820_ (.Y(_1788_),
    .A(_1787_));
 sg13g2_o21ai_1 _5821_ (.B1(_1787_),
    .Y(_1790_),
    .A1(_1784_),
    .A2(_1785_));
 sg13g2_nand4_1 _5822_ (.B(_1771_),
    .C(_1781_),
    .A(net517),
    .Y(_1791_),
    .D(_1790_));
 sg13g2_xnor2_1 _5823_ (.Y(_1792_),
    .A(_1735_),
    .B(_1754_));
 sg13g2_inv_1 _5824_ (.Y(_1793_),
    .A(_1792_));
 sg13g2_nand3_1 _5825_ (.B(_1771_),
    .C(_1793_),
    .A(net517),
    .Y(_1794_));
 sg13g2_nand3_1 _5826_ (.B(_1791_),
    .C(_1794_),
    .A(_1777_),
    .Y(_1795_));
 sg13g2_and2_1 _5827_ (.A(net507),
    .B(_1795_),
    .X(_1796_));
 sg13g2_nand2_2 _5828_ (.Y(_1797_),
    .A(net507),
    .B(_1795_));
 sg13g2_nand3_1 _5829_ (.B(net507),
    .C(_1795_),
    .A(_1770_),
    .Y(_1798_));
 sg13g2_a21o_1 _5830_ (.A2(_1795_),
    .A1(net507),
    .B1(_1792_),
    .X(_1799_));
 sg13g2_nand3_1 _5831_ (.B(_1798_),
    .C(_1799_),
    .A(_1774_),
    .Y(_1801_));
 sg13g2_a21oi_1 _5832_ (.A1(_1769_),
    .A2(_1776_),
    .Y(_1802_),
    .B1(net516));
 sg13g2_a21oi_1 _5833_ (.A1(net509),
    .A2(_1781_),
    .Y(_1803_),
    .B1(_1802_));
 sg13g2_nand2_2 _5834_ (.Y(_1804_),
    .A(_1801_),
    .B(_1803_));
 sg13g2_inv_1 _5835_ (.Y(_1805_),
    .A(_1804_));
 sg13g2_nand2_2 _5836_ (.Y(_1806_),
    .A(net509),
    .B(_1792_));
 sg13g2_nand2_1 _5837_ (.Y(_1807_),
    .A(net509),
    .B(_1785_));
 sg13g2_nand2_1 _5838_ (.Y(_1808_),
    .A(_1781_),
    .B(_1792_));
 sg13g2_a21oi_1 _5839_ (.A1(_1786_),
    .A2(_1787_),
    .Y(_1809_),
    .B1(_1808_));
 sg13g2_a21o_1 _5840_ (.A2(_1809_),
    .A1(net516),
    .B1(_1774_),
    .X(_1810_));
 sg13g2_inv_1 _5841_ (.Y(_1812_),
    .A(_1810_));
 sg13g2_nor2_1 _5842_ (.A(_1805_),
    .B(_1806_),
    .Y(_1813_));
 sg13g2_nand2_1 _5843_ (.Y(_1814_),
    .A(_1785_),
    .B(_1796_));
 sg13g2_nand2_1 _5844_ (.Y(_1815_),
    .A(net516),
    .B(_1808_));
 sg13g2_a22oi_1 _5845_ (.Y(_1816_),
    .B1(_1815_),
    .B2(_1775_),
    .A2(_1797_),
    .A1(_1783_));
 sg13g2_o21ai_1 _5846_ (.B1(_1816_),
    .Y(_1817_),
    .A1(_1813_),
    .A2(_1814_));
 sg13g2_o21ai_1 _5847_ (.B1(_1797_),
    .Y(_1818_),
    .A1(_1787_),
    .A2(_1813_));
 sg13g2_a21oi_1 _5848_ (.A1(_1781_),
    .A2(_1796_),
    .Y(_1819_),
    .B1(_1775_));
 sg13g2_a22oi_1 _5849_ (.Y(_1820_),
    .B1(_1818_),
    .B2(_1819_),
    .A2(_1817_),
    .A1(_1812_));
 sg13g2_nand4_1 _5850_ (.B(_1799_),
    .C(_1812_),
    .A(_1798_),
    .Y(_1821_),
    .D(_1815_));
 sg13g2_nand2_1 _5851_ (.Y(_1823_),
    .A(_1773_),
    .B(_1821_));
 sg13g2_o21ai_1 _5852_ (.B1(_1807_),
    .Y(_1824_),
    .A1(_1820_),
    .A2(_1823_));
 sg13g2_nor2_1 _5853_ (.A(_1781_),
    .B(_1796_),
    .Y(_1825_));
 sg13g2_a21oi_1 _5854_ (.A1(_1793_),
    .A2(_1796_),
    .Y(_1826_),
    .B1(_1825_));
 sg13g2_nand2_1 _5855_ (.Y(_1827_),
    .A(net516),
    .B(_1769_));
 sg13g2_nand2_1 _5856_ (.Y(_1828_),
    .A(_1770_),
    .B(_1797_));
 sg13g2_a22oi_1 _5857_ (.Y(_1829_),
    .B1(_1827_),
    .B2(_1828_),
    .A2(_1826_),
    .A1(_1810_));
 sg13g2_a21oi_2 _5858_ (.B1(_1829_),
    .Y(_1830_),
    .A2(_1788_),
    .A1(net509));
 sg13g2_inv_1 _5859_ (.Y(_1831_),
    .A(_1830_));
 sg13g2_nand2_2 _5860_ (.Y(_1832_),
    .A(_1824_),
    .B(_1831_));
 sg13g2_nand2_1 _5861_ (.Y(_1834_),
    .A(_1775_),
    .B(_1826_));
 sg13g2_nor3_1 _5862_ (.A(_1771_),
    .B(_1787_),
    .C(_1797_),
    .Y(_1835_));
 sg13g2_o21ai_1 _5863_ (.B1(net516),
    .Y(_1836_),
    .A1(net507),
    .A2(_1786_));
 sg13g2_or2_1 _5864_ (.X(_1837_),
    .B(_1836_),
    .A(_1835_));
 sg13g2_a22oi_1 _5865_ (.Y(_1838_),
    .B1(_1834_),
    .B2(_1837_),
    .A2(_1783_),
    .A1(net509));
 sg13g2_inv_1 _5866_ (.Y(_1839_),
    .A(_1838_));
 sg13g2_a22oi_1 _5867_ (.Y(_1840_),
    .B1(_1839_),
    .B2(_1806_),
    .A2(_1824_),
    .A1(_1805_));
 sg13g2_nor2_1 _5868_ (.A(_1832_),
    .B(_1840_),
    .Y(_1841_));
 sg13g2_nand2_1 _5869_ (.Y(_1842_),
    .A(_1806_),
    .B(_1824_));
 sg13g2_nor2_1 _5870_ (.A(_1804_),
    .B(_1831_),
    .Y(_1843_));
 sg13g2_nor2b_1 _5871_ (.A(_1842_),
    .B_N(_1843_),
    .Y(_1845_));
 sg13g2_xnor2_1 _5872_ (.Y(_1846_),
    .A(_1842_),
    .B(_1843_));
 sg13g2_nor2_2 _5873_ (.A(_1804_),
    .B(_1838_),
    .Y(_1847_));
 sg13g2_nand3_1 _5874_ (.B(_1824_),
    .C(_1847_),
    .A(_1806_),
    .Y(_1848_));
 sg13g2_a21oi_1 _5875_ (.A1(_1839_),
    .A2(_1845_),
    .Y(_1849_),
    .B1(_1841_));
 sg13g2_nand2_1 _5876_ (.Y(_1850_),
    .A(_1841_),
    .B(_1846_));
 sg13g2_and2_1 _5877_ (.A(_1832_),
    .B(_1840_),
    .X(_1851_));
 sg13g2_o21ai_1 _5878_ (.B1(_1848_),
    .Y(_1852_),
    .A1(_1841_),
    .A2(_1851_));
 sg13g2_o21ai_1 _5879_ (.B1(_1852_),
    .Y(_1853_),
    .A1(_1831_),
    .A2(_1848_));
 sg13g2_nor2_1 _5880_ (.A(_1824_),
    .B(_1830_),
    .Y(_1854_));
 sg13g2_nand2_2 _5881_ (.Y(_1856_),
    .A(_1738_),
    .B(net508));
 sg13g2_inv_1 _5882_ (.Y(_1857_),
    .A(_1856_));
 sg13g2_nand2_1 _5883_ (.Y(_1858_),
    .A(_1806_),
    .B(_1856_));
 sg13g2_xor2_1 _5884_ (.B(_1854_),
    .A(_1847_),
    .X(_1859_));
 sg13g2_nor2b_1 _5885_ (.A(_1858_),
    .B_N(_1859_),
    .Y(_1860_));
 sg13g2_a21oi_2 _5886_ (.B1(_1860_),
    .Y(_1861_),
    .A2(_1854_),
    .A1(_1847_));
 sg13g2_or2_1 _5887_ (.X(_1862_),
    .B(_1861_),
    .A(_1853_));
 sg13g2_xnor2_1 _5888_ (.Y(_1863_),
    .A(_1824_),
    .B(_1830_));
 sg13g2_and2_1 _5889_ (.A(_1856_),
    .B(_1863_),
    .X(_1864_));
 sg13g2_nand2_1 _5890_ (.Y(_1865_),
    .A(_1805_),
    .B(_1856_));
 sg13g2_nand2_1 _5891_ (.Y(_1867_),
    .A(_1839_),
    .B(_1863_));
 sg13g2_nand2_1 _5892_ (.Y(_1868_),
    .A(_1847_),
    .B(_1864_));
 sg13g2_o21ai_1 _5893_ (.B1(_1868_),
    .Y(_1869_),
    .A1(_1832_),
    .A2(_1838_));
 sg13g2_xnor2_1 _5894_ (.Y(_1870_),
    .A(_1858_),
    .B(_1859_));
 sg13g2_and2_1 _5895_ (.A(_1869_),
    .B(_1870_),
    .X(_1871_));
 sg13g2_xnor2_1 _5896_ (.Y(_1872_),
    .A(_1865_),
    .B(_1867_));
 sg13g2_nor3_2 _5897_ (.A(_1832_),
    .B(_1857_),
    .C(_1865_),
    .Y(_1873_));
 sg13g2_or2_1 _5898_ (.X(_1874_),
    .B(_1870_),
    .A(_1869_));
 sg13g2_nand2b_1 _5899_ (.Y(_1875_),
    .B(_1874_),
    .A_N(_1871_));
 sg13g2_a21oi_1 _5900_ (.A1(_1873_),
    .A2(_1874_),
    .Y(_1876_),
    .B1(_1871_));
 sg13g2_xnor2_1 _5901_ (.Y(_1878_),
    .A(_1853_),
    .B(_1861_));
 sg13g2_o21ai_1 _5902_ (.B1(_1862_),
    .Y(_1879_),
    .A1(_1876_),
    .A2(_1878_));
 sg13g2_xnor2_1 _5903_ (.Y(_1880_),
    .A(_1846_),
    .B(_1849_));
 sg13g2_nand2_1 _5904_ (.Y(_1881_),
    .A(_1879_),
    .B(_1880_));
 sg13g2_xnor2_1 _5905_ (.Y(_1882_),
    .A(_1804_),
    .B(_1806_));
 sg13g2_a21oi_1 _5906_ (.A1(_1831_),
    .A2(_1882_),
    .Y(_1883_),
    .B1(_1845_));
 sg13g2_a21oi_1 _5907_ (.A1(_1850_),
    .A2(_1881_),
    .Y(_1884_),
    .B1(_1883_));
 sg13g2_a21oi_1 _5908_ (.A1(_1805_),
    .A2(_1806_),
    .Y(_1885_),
    .B1(_1884_));
 sg13g2_nand3_1 _5909_ (.B(_1881_),
    .C(_1883_),
    .A(_1850_),
    .Y(_1886_));
 sg13g2_nand2b_1 _5910_ (.Y(_1887_),
    .B(_1886_),
    .A_N(_1884_));
 sg13g2_xnor2_1 _5911_ (.Y(_1889_),
    .A(_1876_),
    .B(_1878_));
 sg13g2_nor2_1 _5912_ (.A(_1780_),
    .B(_1889_),
    .Y(_1890_));
 sg13g2_o21ai_1 _5913_ (.B1(_1774_),
    .Y(_1891_),
    .A1(net506),
    .A2(_1887_));
 sg13g2_o21ai_1 _5914_ (.B1(_1872_),
    .Y(_1892_),
    .A1(_1832_),
    .A2(_1857_));
 sg13g2_nand2b_1 _5915_ (.Y(_1893_),
    .B(_1892_),
    .A_N(_1873_));
 sg13g2_a22oi_1 _5916_ (.Y(_1894_),
    .B1(_1893_),
    .B2(_1776_),
    .A2(net506),
    .A1(_1775_));
 sg13g2_o21ai_1 _5917_ (.B1(_1894_),
    .Y(_1895_),
    .A1(_1890_),
    .A2(_1891_));
 sg13g2_o21ai_1 _5918_ (.B1(_1895_),
    .Y(_1896_),
    .A1(_1773_),
    .A2(_1885_));
 sg13g2_nand2_1 _5919_ (.Y(_1897_),
    .A(net468),
    .B(_1896_));
 sg13g2_mux2_1 _5920_ (.A0(_1889_),
    .A1(_1893_),
    .S(net506),
    .X(_1898_));
 sg13g2_nor2_1 _5921_ (.A(net507),
    .B(_1885_),
    .Y(_1900_));
 sg13g2_nor2_1 _5922_ (.A(_1797_),
    .B(_1887_),
    .Y(_1901_));
 sg13g2_o21ai_1 _5923_ (.B1(_1774_),
    .Y(_1902_),
    .A1(_1900_),
    .A2(_1901_));
 sg13g2_o21ai_1 _5924_ (.B1(_1902_),
    .Y(_1903_),
    .A1(net517),
    .A2(_1898_));
 sg13g2_xnor2_1 _5925_ (.Y(_1904_),
    .A(_2912_),
    .B(_1903_));
 sg13g2_a221oi_1 _5926_ (.B2(_1830_),
    .C1(_1884_),
    .B1(_1805_),
    .A1(net508),
    .Y(_1905_),
    .A2(_1792_));
 sg13g2_xnor2_1 _5927_ (.Y(_1906_),
    .A(_1879_),
    .B(_1880_));
 sg13g2_inv_1 _5928_ (.Y(_1907_),
    .A(_1906_));
 sg13g2_a21oi_1 _5929_ (.A1(net506),
    .A2(_1906_),
    .Y(_1908_),
    .B1(_1775_));
 sg13g2_o21ai_1 _5930_ (.B1(_1908_),
    .Y(_1909_),
    .A1(net506),
    .A2(_1905_));
 sg13g2_nor2_1 _5931_ (.A(_1739_),
    .B(_1786_),
    .Y(_1911_));
 sg13g2_a21oi_1 _5932_ (.A1(net508),
    .A2(_1911_),
    .Y(_1912_),
    .B1(_1864_));
 sg13g2_nand2b_1 _5933_ (.Y(_1913_),
    .B(net506),
    .A_N(_1912_));
 sg13g2_xor2_1 _5934_ (.B(_1875_),
    .A(_1873_),
    .X(_1914_));
 sg13g2_o21ai_1 _5935_ (.B1(_1913_),
    .Y(_1915_),
    .A1(net506),
    .A2(_1914_));
 sg13g2_nand2b_1 _5936_ (.Y(_1916_),
    .B(_1915_),
    .A_N(net517));
 sg13g2_and2_2 _5937_ (.A(_1909_),
    .B(_1916_),
    .X(_1917_));
 sg13g2_or2_1 _5938_ (.X(_1918_),
    .B(_1917_),
    .A(net470));
 sg13g2_nand2_1 _5939_ (.Y(_1919_),
    .A(net470),
    .B(_1917_));
 sg13g2_nor2_1 _5940_ (.A(_1775_),
    .B(_1915_),
    .Y(_1920_));
 sg13g2_nor3_1 _5941_ (.A(net508),
    .B(_1776_),
    .C(_1920_),
    .Y(_1922_));
 sg13g2_a21oi_2 _5942_ (.B1(_1922_),
    .Y(_1923_),
    .A2(_1907_),
    .A1(net508));
 sg13g2_nor2_1 _5943_ (.A(net472),
    .B(_1923_),
    .Y(_1924_));
 sg13g2_nor3_1 _5944_ (.A(net475),
    .B(net472),
    .C(_1923_),
    .Y(_1925_));
 sg13g2_nor2_1 _5945_ (.A(_1775_),
    .B(_1898_),
    .Y(_1926_));
 sg13g2_xnor2_1 _5946_ (.Y(_1927_),
    .A(_1824_),
    .B(_1838_));
 sg13g2_a21oi_1 _5947_ (.A1(_1776_),
    .A2(_1927_),
    .Y(_1928_),
    .B1(_1926_));
 sg13g2_o21ai_1 _5948_ (.B1(_1928_),
    .Y(_1929_),
    .A1(_1773_),
    .A2(_1887_));
 sg13g2_xnor2_1 _5949_ (.Y(_1930_),
    .A(net468),
    .B(_1896_));
 sg13g2_nor2_1 _5950_ (.A(_1780_),
    .B(_1914_),
    .Y(_1931_));
 sg13g2_a21oi_1 _5951_ (.A1(_1780_),
    .A2(_1907_),
    .Y(_1933_),
    .B1(_1931_));
 sg13g2_nand2_1 _5952_ (.Y(_1934_),
    .A(_1810_),
    .B(_1933_));
 sg13g2_o21ai_1 _5953_ (.B1(_1775_),
    .Y(_1935_),
    .A1(net506),
    .A2(_1912_));
 sg13g2_a22oi_1 _5954_ (.Y(_1936_),
    .B1(_1934_),
    .B2(_1935_),
    .A2(_1905_),
    .A1(net508));
 sg13g2_inv_1 _5955_ (.Y(_1937_),
    .A(_1936_));
 sg13g2_a21oi_1 _5956_ (.A1(_2856_),
    .A2(_1936_),
    .Y(_1938_),
    .B1(_1930_));
 sg13g2_nand2_1 _5957_ (.Y(_1939_),
    .A(_1904_),
    .B(_1919_));
 sg13g2_nor2_1 _5958_ (.A(_3259_),
    .B(_1601_),
    .Y(_1940_));
 sg13g2_nor4_1 _5959_ (.A(net571),
    .B(_0700_),
    .C(_1601_),
    .D(_1661_),
    .Y(_1941_));
 sg13g2_nor4_2 _5960_ (.A(_0184_),
    .B(_2924_),
    .C(_1940_),
    .Y(_1942_),
    .D(_1941_));
 sg13g2_nand2_1 _5961_ (.Y(_1944_),
    .A(_2855_),
    .B(_1937_));
 sg13g2_and2_1 _5962_ (.A(_1930_),
    .B(_1944_),
    .X(_1945_));
 sg13g2_xor2_1 _5963_ (.B(_1924_),
    .A(net475),
    .X(_1946_));
 sg13g2_nand2_1 _5964_ (.Y(_1947_),
    .A(_1929_),
    .B(_1946_));
 sg13g2_nand3b_1 _5965_ (.B(_1944_),
    .C(net475),
    .Y(_1948_),
    .A_N(_1924_));
 sg13g2_nor2_1 _5966_ (.A(_1925_),
    .B(_1929_),
    .Y(_1949_));
 sg13g2_mux2_1 _5967_ (.A0(_1949_),
    .A1(_1948_),
    .S(_1938_),
    .X(_1950_));
 sg13g2_nand3b_1 _5968_ (.B(_1918_),
    .C(_1897_),
    .Y(_1951_),
    .A_N(_1904_));
 sg13g2_a21oi_1 _5969_ (.A1(_1918_),
    .A2(_1919_),
    .Y(_1952_),
    .B1(_1897_));
 sg13g2_nand4_1 _5970_ (.B(_1942_),
    .C(_1947_),
    .A(_1939_),
    .Y(_1953_),
    .D(_1951_));
 sg13g2_or4_2 _5971_ (.A(_1945_),
    .B(_1950_),
    .C(_1952_),
    .D(_1953_),
    .X(_1955_));
 sg13g2_nand3_1 _5972_ (.B(_1702_),
    .C(_1955_),
    .A(_3257_),
    .Y(_1956_));
 sg13g2_a21oi_1 _5973_ (.A1(_2535_),
    .A2(_0368_),
    .Y(_1957_),
    .B1(\hvsync_gen.hpos[4] ));
 sg13g2_a21oi_1 _5974_ (.A1(_2535_),
    .A2(_0368_),
    .Y(_1958_),
    .B1(_0064_));
 sg13g2_and2_1 _5975_ (.A(net595),
    .B(_2639_),
    .X(_1959_));
 sg13g2_a21oi_1 _5976_ (.A1(net595),
    .A2(_2639_),
    .Y(_1960_),
    .B1(net591));
 sg13g2_o21ai_1 _5977_ (.B1(_1960_),
    .Y(_1961_),
    .A1(net551),
    .A2(_1958_));
 sg13g2_nand3_1 _5978_ (.B(net588),
    .C(_1961_),
    .A(net585),
    .Y(_1962_));
 sg13g2_a21o_1 _5979_ (.A2(_1961_),
    .A1(net588),
    .B1(net585),
    .X(_1963_));
 sg13g2_nand2_1 _5980_ (.Y(_1964_),
    .A(_1962_),
    .B(_1963_));
 sg13g2_inv_1 _5981_ (.Y(_1966_),
    .A(_1964_));
 sg13g2_xnor2_1 _5982_ (.Y(_1967_),
    .A(_3081_),
    .B(_1961_));
 sg13g2_o21ai_1 _5983_ (.B1(_0377_),
    .Y(_1968_),
    .A1(net551),
    .A2(_2619_));
 sg13g2_nand2_2 _5984_ (.Y(_1969_),
    .A(_0376_),
    .B(_1968_));
 sg13g2_nand3_1 _5985_ (.B(_2611_),
    .C(_2612_),
    .A(net542),
    .Y(_1970_));
 sg13g2_o21ai_1 _5986_ (.B1(_1970_),
    .Y(_1971_),
    .A1(net542),
    .A2(net603));
 sg13g2_xnor2_1 _5987_ (.Y(_1972_),
    .A(_0016_),
    .B(_2612_));
 sg13g2_a21oi_2 _5988_ (.B1(_0372_),
    .Y(_1973_),
    .A2(_1972_),
    .A1(net542));
 sg13g2_nor3_1 _5989_ (.A(_1969_),
    .B(_1971_),
    .C(_1973_),
    .Y(_1974_));
 sg13g2_o21ai_1 _5990_ (.B1(_0371_),
    .Y(_1975_),
    .A1(_3114_),
    .A2(_2612_));
 sg13g2_xnor2_1 _5991_ (.Y(_1977_),
    .A(_3191_),
    .B(_1975_));
 sg13g2_nor4_2 _5992_ (.A(_1969_),
    .B(_1971_),
    .C(_1973_),
    .Y(_1978_),
    .D(_1977_));
 sg13g2_nor2_1 _5993_ (.A(net595),
    .B(_2639_),
    .Y(_1979_));
 sg13g2_o21ai_1 _5994_ (.B1(net551),
    .Y(_1980_),
    .A1(_1959_),
    .A2(_1979_));
 sg13g2_xnor2_1 _5995_ (.Y(_1981_),
    .A(_0018_),
    .B(_1957_));
 sg13g2_o21ai_1 _5996_ (.B1(_1980_),
    .Y(_1982_),
    .A1(net552),
    .A2(_1981_));
 sg13g2_nand2_1 _5997_ (.Y(_1983_),
    .A(_1978_),
    .B(_1982_));
 sg13g2_or2_1 _5998_ (.X(_1984_),
    .B(_1959_),
    .A(_0014_));
 sg13g2_a21oi_1 _5999_ (.A1(net589),
    .A2(_1959_),
    .Y(_1985_),
    .B1(net543));
 sg13g2_xnor2_1 _6000_ (.Y(_1986_),
    .A(_3092_),
    .B(_1958_));
 sg13g2_a22oi_1 _6001_ (.Y(_1988_),
    .B1(_1986_),
    .B2(net543),
    .A2(_1985_),
    .A1(_1984_));
 sg13g2_and3_1 _6002_ (.X(_1989_),
    .A(_1978_),
    .B(_1982_),
    .C(_1988_));
 sg13g2_nand3_1 _6003_ (.B(_1982_),
    .C(_1988_),
    .A(_1978_),
    .Y(_1990_));
 sg13g2_o21ai_1 _6004_ (.B1(_3048_),
    .Y(_1991_),
    .A1(_1967_),
    .A2(_1990_));
 sg13g2_xnor2_1 _6005_ (.Y(_1992_),
    .A(_3048_),
    .B(_1962_));
 sg13g2_xnor2_1 _6006_ (.Y(_1993_),
    .A(net583),
    .B(_1962_));
 sg13g2_and2_1 _6007_ (.A(_1964_),
    .B(_1992_),
    .X(_1994_));
 sg13g2_a21oi_2 _6008_ (.B1(_1994_),
    .Y(_1995_),
    .A2(_1991_),
    .A1(_1966_));
 sg13g2_a21o_2 _6009_ (.A2(_1991_),
    .A1(_1966_),
    .B1(_1994_),
    .X(_1996_));
 sg13g2_o21ai_1 _6010_ (.B1(_1967_),
    .Y(_1997_),
    .A1(_1989_),
    .A2(_1993_));
 sg13g2_nand3b_1 _6011_ (.B(_1990_),
    .C(_1992_),
    .Y(_1999_),
    .A_N(_1967_));
 sg13g2_and2_1 _6012_ (.A(_1997_),
    .B(_1999_),
    .X(_2000_));
 sg13g2_nand3_1 _6013_ (.B(_1988_),
    .C(_1992_),
    .A(_1983_),
    .Y(_2001_));
 sg13g2_a21o_1 _6014_ (.A2(_1992_),
    .A1(_1983_),
    .B1(_1988_),
    .X(_2002_));
 sg13g2_nand2_1 _6015_ (.Y(_2003_),
    .A(_2001_),
    .B(_2002_));
 sg13g2_nand4_1 _6016_ (.B(_1999_),
    .C(_2001_),
    .A(_1997_),
    .Y(_2004_),
    .D(_2002_));
 sg13g2_nor2_2 _6017_ (.A(_1996_),
    .B(_2000_),
    .Y(_2005_));
 sg13g2_and2_2 _6018_ (.A(_1995_),
    .B(_2004_),
    .X(_2006_));
 sg13g2_nand2_2 _6019_ (.Y(_2007_),
    .A(_1995_),
    .B(_2004_));
 sg13g2_nor2_2 _6020_ (.A(_1996_),
    .B(_2004_),
    .Y(_2008_));
 sg13g2_nand2_2 _6021_ (.Y(_2010_),
    .A(_1995_),
    .B(_2007_));
 sg13g2_o21ai_1 _6022_ (.B1(_1992_),
    .Y(_2011_),
    .A1(_1969_),
    .A2(_1971_));
 sg13g2_xnor2_1 _6023_ (.Y(_2012_),
    .A(_1973_),
    .B(_2011_));
 sg13g2_inv_1 _6024_ (.Y(_2013_),
    .A(_2012_));
 sg13g2_nand2_1 _6025_ (.Y(_2014_),
    .A(_1969_),
    .B(_1992_));
 sg13g2_xor2_1 _6026_ (.B(_2014_),
    .A(_1971_),
    .X(_2015_));
 sg13g2_nor2_1 _6027_ (.A(_0376_),
    .B(_1993_),
    .Y(_2016_));
 sg13g2_xnor2_1 _6028_ (.Y(_2017_),
    .A(_1968_),
    .B(_2016_));
 sg13g2_a21o_1 _6029_ (.A2(_2017_),
    .A1(_2015_),
    .B1(_2012_),
    .X(_2018_));
 sg13g2_nor2_1 _6030_ (.A(_1974_),
    .B(_1993_),
    .Y(_2019_));
 sg13g2_xor2_1 _6031_ (.B(_2019_),
    .A(_1977_),
    .X(_2021_));
 sg13g2_xnor2_1 _6032_ (.Y(_2022_),
    .A(_1977_),
    .B(_2019_));
 sg13g2_nor3_1 _6033_ (.A(_1996_),
    .B(_2004_),
    .C(_2021_),
    .Y(_2023_));
 sg13g2_nor2_1 _6034_ (.A(_1978_),
    .B(_1993_),
    .Y(_2024_));
 sg13g2_xnor2_1 _6035_ (.Y(_2025_),
    .A(_1982_),
    .B(_2024_));
 sg13g2_nand2_1 _6036_ (.Y(_2026_),
    .A(net515),
    .B(_2025_));
 sg13g2_nand3b_1 _6037_ (.B(_1989_),
    .C(_1994_),
    .Y(_2027_),
    .A_N(_1967_));
 sg13g2_o21ai_1 _6038_ (.B1(_2027_),
    .Y(_2028_),
    .A1(_1996_),
    .A2(_2000_));
 sg13g2_a221oi_1 _6039_ (.B2(net515),
    .C1(_2028_),
    .B1(_2025_),
    .A1(_2018_),
    .Y(_2029_),
    .A2(_2023_));
 sg13g2_nand2_2 _6040_ (.Y(_2030_),
    .A(_2010_),
    .B(_2029_));
 sg13g2_inv_2 _6041_ (.Y(_2032_),
    .A(_2030_));
 sg13g2_nand2b_1 _6042_ (.Y(_2033_),
    .B(_2021_),
    .A_N(net505));
 sg13g2_nor3_2 _6043_ (.A(_1996_),
    .B(_2004_),
    .C(_2025_),
    .Y(_2034_));
 sg13g2_nand2_1 _6044_ (.Y(_2035_),
    .A(_2008_),
    .B(_2026_));
 sg13g2_a21oi_1 _6045_ (.A1(_2022_),
    .A2(_2034_),
    .Y(_2036_),
    .B1(_2013_));
 sg13g2_nor2_1 _6046_ (.A(_2010_),
    .B(_2022_),
    .Y(_2037_));
 sg13g2_o21ai_1 _6047_ (.B1(_1995_),
    .Y(_2038_),
    .A1(_2004_),
    .A2(_2021_));
 sg13g2_and2_2 _6048_ (.A(_2026_),
    .B(_2038_),
    .X(_2039_));
 sg13g2_a21oi_1 _6049_ (.A1(net505),
    .A2(_2036_),
    .Y(_2040_),
    .B1(_2039_));
 sg13g2_a22oi_1 _6050_ (.Y(_2041_),
    .B1(_2040_),
    .B2(_2033_),
    .A2(_2039_),
    .A1(_2000_));
 sg13g2_nand2_1 _6051_ (.Y(_2043_),
    .A(_2013_),
    .B(_2015_));
 sg13g2_nand3_1 _6052_ (.B(_2034_),
    .C(_2043_),
    .A(_2022_),
    .Y(_2044_));
 sg13g2_nand2_1 _6053_ (.Y(_2045_),
    .A(_2007_),
    .B(_2044_));
 sg13g2_mux2_1 _6054_ (.A0(_2003_),
    .A1(_2025_),
    .S(net505),
    .X(_2046_));
 sg13g2_a221oi_1 _6055_ (.B2(_2006_),
    .C1(_2037_),
    .B1(_2046_),
    .A1(_1996_),
    .Y(_2047_),
    .A2(_2041_));
 sg13g2_nand2b_1 _6056_ (.Y(_2048_),
    .B(_2036_),
    .A_N(net505));
 sg13g2_a21oi_1 _6057_ (.A1(_2022_),
    .A2(_2034_),
    .Y(_2049_),
    .B1(_2015_));
 sg13g2_a21oi_1 _6058_ (.A1(net505),
    .A2(_2049_),
    .Y(_2050_),
    .B1(_2039_));
 sg13g2_nand3_1 _6059_ (.B(_2048_),
    .C(_2050_),
    .A(_2045_),
    .Y(_2051_));
 sg13g2_nand2_1 _6060_ (.Y(_2052_),
    .A(_2022_),
    .B(net505));
 sg13g2_o21ai_1 _6061_ (.B1(_2052_),
    .Y(_2054_),
    .A1(_2025_),
    .A2(net505));
 sg13g2_o21ai_1 _6062_ (.B1(_2007_),
    .Y(_2055_),
    .A1(_1995_),
    .A2(_2054_));
 sg13g2_a22oi_1 _6063_ (.Y(_2056_),
    .B1(_2051_),
    .B2(_2055_),
    .A2(_2017_),
    .A1(net515));
 sg13g2_nor2_1 _6064_ (.A(_0375_),
    .B(_2010_),
    .Y(_2057_));
 sg13g2_a21oi_1 _6065_ (.A1(_0375_),
    .A2(_2025_),
    .Y(_2058_),
    .B1(_2010_));
 sg13g2_nor2_2 _6066_ (.A(_2034_),
    .B(_2056_),
    .Y(_2059_));
 sg13g2_nor2_2 _6067_ (.A(_2047_),
    .B(_2057_),
    .Y(_2060_));
 sg13g2_nor3_1 _6068_ (.A(_2047_),
    .B(_2056_),
    .C(_2058_),
    .Y(_2061_));
 sg13g2_o21ai_1 _6069_ (.B1(_2045_),
    .Y(_2062_),
    .A1(_2039_),
    .A2(_2054_));
 sg13g2_a21o_1 _6070_ (.A2(net505),
    .A1(_2003_),
    .B1(_2005_),
    .X(_2063_));
 sg13g2_nand2_1 _6071_ (.Y(_2065_),
    .A(_2062_),
    .B(_2063_));
 sg13g2_a22oi_1 _6072_ (.Y(_2066_),
    .B1(_2062_),
    .B2(_2063_),
    .A2(_2012_),
    .A1(net515));
 sg13g2_o21ai_1 _6073_ (.B1(_2065_),
    .Y(_2067_),
    .A1(_2010_),
    .A2(_2013_));
 sg13g2_nor2_1 _6074_ (.A(_2010_),
    .B(_2015_),
    .Y(_2068_));
 sg13g2_a221oi_1 _6075_ (.B2(_2039_),
    .C1(_2068_),
    .B1(_2046_),
    .A1(_2006_),
    .Y(_2069_),
    .A2(_2041_));
 sg13g2_inv_1 _6076_ (.Y(_2070_),
    .A(_2069_));
 sg13g2_nor2_2 _6077_ (.A(_2066_),
    .B(_2069_),
    .Y(_2071_));
 sg13g2_o21ai_1 _6078_ (.B1(_2058_),
    .Y(_2072_),
    .A1(_2047_),
    .A2(_2056_));
 sg13g2_nand2b_1 _6079_ (.Y(_2073_),
    .B(_2072_),
    .A_N(_2061_));
 sg13g2_a22oi_1 _6080_ (.Y(_2074_),
    .B1(_2071_),
    .B2(_2072_),
    .A2(_2060_),
    .A1(_2059_));
 sg13g2_nor2_1 _6081_ (.A(_2034_),
    .B(_2069_),
    .Y(_2076_));
 sg13g2_nor2_2 _6082_ (.A(_2047_),
    .B(_2069_),
    .Y(_2077_));
 sg13g2_xor2_1 _6083_ (.B(_2077_),
    .A(_2059_),
    .X(_2078_));
 sg13g2_nor2b_1 _6084_ (.A(_2074_),
    .B_N(_2078_),
    .Y(_2079_));
 sg13g2_xnor2_1 _6085_ (.Y(_2080_),
    .A(_2074_),
    .B(_2078_));
 sg13g2_nor2_1 _6086_ (.A(_2047_),
    .B(_2066_),
    .Y(_2081_));
 sg13g2_o21ai_1 _6087_ (.B1(_2066_),
    .Y(_2082_),
    .A1(_2047_),
    .A2(_2069_));
 sg13g2_xnor2_1 _6088_ (.Y(_2083_),
    .A(_2067_),
    .B(_2077_));
 sg13g2_xnor2_1 _6089_ (.Y(_2084_),
    .A(_2059_),
    .B(_2083_));
 sg13g2_and2_1 _6090_ (.A(_2080_),
    .B(_2084_),
    .X(_2085_));
 sg13g2_xnor2_1 _6091_ (.Y(_2087_),
    .A(_2071_),
    .B(_2073_));
 sg13g2_inv_1 _6092_ (.Y(_2088_),
    .A(_2087_));
 sg13g2_mux2_1 _6093_ (.A0(_2074_),
    .A1(_2088_),
    .S(_2067_),
    .X(_2089_));
 sg13g2_a22oi_1 _6094_ (.Y(_2090_),
    .B1(_2082_),
    .B2(_2059_),
    .A2(_2081_),
    .A1(_2070_));
 sg13g2_nand4_1 _6095_ (.B(_2067_),
    .C(_2077_),
    .A(_2059_),
    .Y(_2091_),
    .D(_2080_));
 sg13g2_a21o_1 _6096_ (.A2(_2077_),
    .A1(_2059_),
    .B1(_2079_),
    .X(_2092_));
 sg13g2_o21ai_1 _6097_ (.B1(_2091_),
    .Y(_2093_),
    .A1(_2085_),
    .A2(_2092_));
 sg13g2_or2_1 _6098_ (.X(_2094_),
    .B(_2093_),
    .A(_2090_));
 sg13g2_xor2_1 _6099_ (.B(_2093_),
    .A(_2090_),
    .X(_2095_));
 sg13g2_nand2b_1 _6100_ (.Y(_2096_),
    .B(_2095_),
    .A_N(_2089_));
 sg13g2_xnor2_1 _6101_ (.Y(_2098_),
    .A(_2067_),
    .B(_2087_));
 sg13g2_inv_1 _6102_ (.Y(_2099_),
    .A(_2098_));
 sg13g2_nor2_2 _6103_ (.A(_2056_),
    .B(_2066_),
    .Y(_2100_));
 sg13g2_nor2_1 _6104_ (.A(_2060_),
    .B(_2100_),
    .Y(_2101_));
 sg13g2_nor2_2 _6105_ (.A(_2056_),
    .B(_2069_),
    .Y(_2102_));
 sg13g2_a21oi_1 _6106_ (.A1(_2060_),
    .A2(_2100_),
    .Y(_2103_),
    .B1(_2102_));
 sg13g2_nor2_1 _6107_ (.A(_2101_),
    .B(_2103_),
    .Y(_2104_));
 sg13g2_nand2b_2 _6108_ (.Y(_2105_),
    .B(_2071_),
    .A_N(_2057_));
 sg13g2_xor2_1 _6109_ (.B(_2100_),
    .A(_2060_),
    .X(_2106_));
 sg13g2_xnor2_1 _6110_ (.Y(_2107_),
    .A(_2102_),
    .B(_2106_));
 sg13g2_or2_1 _6111_ (.X(_2109_),
    .B(_2107_),
    .A(_2105_));
 sg13g2_xor2_1 _6112_ (.B(_2104_),
    .A(_2098_),
    .X(_2110_));
 sg13g2_nor2_1 _6113_ (.A(_2109_),
    .B(_2110_),
    .Y(_2111_));
 sg13g2_a21oi_1 _6114_ (.A1(_2099_),
    .A2(_2104_),
    .Y(_2112_),
    .B1(_2111_));
 sg13g2_nor2b_1 _6115_ (.A(_2095_),
    .B_N(_2089_),
    .Y(_2113_));
 sg13g2_xnor2_1 _6116_ (.Y(_2114_),
    .A(_2089_),
    .B(_2095_));
 sg13g2_o21ai_1 _6117_ (.B1(_2096_),
    .Y(_2115_),
    .A1(_2112_),
    .A2(_2113_));
 sg13g2_nand2b_1 _6118_ (.Y(_2116_),
    .B(_2066_),
    .A_N(_2047_));
 sg13g2_xor2_1 _6119_ (.B(_2116_),
    .A(_2076_),
    .X(_2117_));
 sg13g2_a21oi_1 _6120_ (.A1(_2091_),
    .A2(_2094_),
    .Y(_2118_),
    .B1(_2117_));
 sg13g2_nand3_1 _6121_ (.B(_2094_),
    .C(_2117_),
    .A(_2091_),
    .Y(_2120_));
 sg13g2_nand2b_1 _6122_ (.Y(_2121_),
    .B(_2120_),
    .A_N(_2118_));
 sg13g2_nor2b_1 _6123_ (.A(_2121_),
    .B_N(_2115_),
    .Y(_2122_));
 sg13g2_xnor2_1 _6124_ (.Y(_2123_),
    .A(_2115_),
    .B(_2121_));
 sg13g2_nand2_1 _6125_ (.Y(_2124_),
    .A(_2032_),
    .B(_2123_));
 sg13g2_xnor2_1 _6126_ (.Y(_2125_),
    .A(_2109_),
    .B(_2110_));
 sg13g2_o21ai_1 _6127_ (.B1(_2124_),
    .Y(_2126_),
    .A1(_2032_),
    .A2(_2125_));
 sg13g2_o21ai_1 _6128_ (.B1(_2082_),
    .Y(_2127_),
    .A1(_2035_),
    .A2(_2081_));
 sg13g2_a21oi_1 _6129_ (.A1(_2035_),
    .A2(_2081_),
    .Y(_2128_),
    .B1(_2127_));
 sg13g2_o21ai_1 _6130_ (.B1(_2128_),
    .Y(_2129_),
    .A1(_2118_),
    .A2(_2122_));
 sg13g2_and3_1 _6131_ (.X(_2131_),
    .A(_2035_),
    .B(_2116_),
    .C(_2129_));
 sg13g2_a22oi_1 _6132_ (.Y(_2132_),
    .B1(_2131_),
    .B2(_2005_),
    .A2(_2126_),
    .A1(_2007_));
 sg13g2_inv_1 _6133_ (.Y(_2133_),
    .A(_2132_));
 sg13g2_nor2_1 _6134_ (.A(net515),
    .B(_2132_),
    .Y(_2134_));
 sg13g2_inv_2 _6135_ (.Y(_2135_),
    .A(_2134_));
 sg13g2_nand2_1 _6136_ (.Y(_2136_),
    .A(_2910_),
    .B(_2135_));
 sg13g2_xnor2_1 _6137_ (.Y(_2137_),
    .A(_2910_),
    .B(_2135_));
 sg13g2_or3_1 _6138_ (.A(_2118_),
    .B(_2122_),
    .C(_2128_),
    .X(_2138_));
 sg13g2_and2_1 _6139_ (.A(_2129_),
    .B(_2138_),
    .X(_2139_));
 sg13g2_or2_1 _6140_ (.X(_2140_),
    .B(_2139_),
    .A(_2032_));
 sg13g2_and2_1 _6141_ (.A(_2047_),
    .B(_2129_),
    .X(_2142_));
 sg13g2_a21oi_1 _6142_ (.A1(_2032_),
    .A2(_2142_),
    .Y(_2143_),
    .B1(_2007_));
 sg13g2_xor2_1 _6143_ (.B(_2107_),
    .A(_2105_),
    .X(_2144_));
 sg13g2_xnor2_1 _6144_ (.Y(_2145_),
    .A(_2112_),
    .B(_2114_));
 sg13g2_mux2_1 _6145_ (.A0(_2144_),
    .A1(_2145_),
    .S(_2032_),
    .X(_2146_));
 sg13g2_a22oi_1 _6146_ (.Y(_2147_),
    .B1(_2146_),
    .B2(_1996_),
    .A2(_2143_),
    .A1(_2140_));
 sg13g2_or2_1 _6147_ (.X(_2148_),
    .B(_2147_),
    .A(_2491_));
 sg13g2_xnor2_1 _6148_ (.Y(_2149_),
    .A(_2491_),
    .B(_2147_));
 sg13g2_nor2_1 _6149_ (.A(_2032_),
    .B(_2123_),
    .Y(_2150_));
 sg13g2_nor2_1 _6150_ (.A(_2007_),
    .B(_2150_),
    .Y(_2151_));
 sg13g2_o21ai_1 _6151_ (.B1(_2151_),
    .Y(_2153_),
    .A1(_2030_),
    .A2(_2131_));
 sg13g2_nor2_1 _6152_ (.A(_2030_),
    .B(_2125_),
    .Y(_2154_));
 sg13g2_o21ai_1 _6153_ (.B1(_2069_),
    .Y(_2155_),
    .A1(_2057_),
    .A2(_2066_));
 sg13g2_nand3_1 _6154_ (.B(net515),
    .C(_2017_),
    .A(_0376_),
    .Y(_2156_));
 sg13g2_and3_1 _6155_ (.X(_2157_),
    .A(_2105_),
    .B(_2155_),
    .C(_2156_));
 sg13g2_a21oi_1 _6156_ (.A1(_2030_),
    .A2(_2157_),
    .Y(_2158_),
    .B1(_2154_));
 sg13g2_o21ai_1 _6157_ (.B1(_2153_),
    .Y(_2159_),
    .A1(_1995_),
    .A2(_2158_));
 sg13g2_nor2b_1 _6158_ (.A(_2828_),
    .B_N(_2159_),
    .Y(_2160_));
 sg13g2_xor2_1 _6159_ (.B(_2159_),
    .A(_2828_),
    .X(_2161_));
 sg13g2_inv_1 _6160_ (.Y(_2162_),
    .A(_2161_));
 sg13g2_mux2_1 _6161_ (.A0(_2139_),
    .A1(_2145_),
    .S(_2030_),
    .X(_2164_));
 sg13g2_nor2_1 _6162_ (.A(_2026_),
    .B(_2142_),
    .Y(_2165_));
 sg13g2_nor2_1 _6163_ (.A(_2006_),
    .B(_2030_),
    .Y(_2166_));
 sg13g2_a221oi_1 _6164_ (.B2(_2144_),
    .C1(_2165_),
    .B1(_2166_),
    .A1(_2006_),
    .Y(_2167_),
    .A2(_2164_));
 sg13g2_nand2b_1 _6165_ (.Y(_2168_),
    .B(_2847_),
    .A_N(_2167_));
 sg13g2_xnor2_1 _6166_ (.Y(_2169_),
    .A(_2847_),
    .B(_2167_));
 sg13g2_nand2_1 _6167_ (.Y(_2170_),
    .A(net515),
    .B(_2131_));
 sg13g2_a22oi_1 _6168_ (.Y(_2171_),
    .B1(_2157_),
    .B2(_2166_),
    .A2(_2126_),
    .A1(_2006_));
 sg13g2_nand2_2 _6169_ (.Y(_2172_),
    .A(_2170_),
    .B(_2171_));
 sg13g2_inv_2 _6170_ (.Y(_2173_),
    .A(_2172_));
 sg13g2_nand2_1 _6171_ (.Y(_2175_),
    .A(_2860_),
    .B(_2172_));
 sg13g2_xnor2_1 _6172_ (.Y(_2176_),
    .A(_2860_),
    .B(_2173_));
 sg13g2_inv_1 _6173_ (.Y(_2177_),
    .A(_2176_));
 sg13g2_a21oi_1 _6174_ (.A1(_2056_),
    .A2(_2069_),
    .Y(_2178_),
    .B1(_1995_));
 sg13g2_nor2b_1 _6175_ (.A(_2102_),
    .B_N(_2178_),
    .Y(_2179_));
 sg13g2_a221oi_1 _6176_ (.B2(_2006_),
    .C1(_2179_),
    .B1(_2146_),
    .A1(_2008_),
    .Y(_2180_),
    .A2(_2139_));
 sg13g2_nor2_2 _6177_ (.A(_2874_),
    .B(_2180_),
    .Y(_2181_));
 sg13g2_o21ai_1 _6178_ (.B1(_2027_),
    .Y(_2182_),
    .A1(_2007_),
    .A2(_2158_));
 sg13g2_a21o_2 _6179_ (.A2(_2123_),
    .A1(net515),
    .B1(_2182_),
    .X(_2183_));
 sg13g2_and2_1 _6180_ (.A(net474),
    .B(_2183_),
    .X(_2184_));
 sg13g2_nand2_2 _6181_ (.Y(_2186_),
    .A(_2874_),
    .B(_2180_));
 sg13g2_nand2b_1 _6182_ (.Y(_2187_),
    .B(_2186_),
    .A_N(_2181_));
 sg13g2_a21oi_2 _6183_ (.B1(_2181_),
    .Y(_2188_),
    .A2(_2186_),
    .A1(_2184_));
 sg13g2_o21ai_1 _6184_ (.B1(_2175_),
    .Y(_2189_),
    .A1(_2177_),
    .A2(_2188_));
 sg13g2_nand2_1 _6185_ (.Y(_2190_),
    .A(_2169_),
    .B(_2189_));
 sg13g2_nand2_1 _6186_ (.Y(_2191_),
    .A(_2168_),
    .B(_2190_));
 sg13g2_a21oi_1 _6187_ (.A1(_2162_),
    .A2(_2191_),
    .Y(_2192_),
    .B1(_2160_));
 sg13g2_nor2_1 _6188_ (.A(_2149_),
    .B(_2192_),
    .Y(_2193_));
 sg13g2_nand2_1 _6189_ (.Y(_2194_),
    .A(_2007_),
    .B(_2164_));
 sg13g2_nand2b_1 _6190_ (.Y(_2195_),
    .B(_2005_),
    .A_N(_2142_));
 sg13g2_a21o_2 _6191_ (.A2(_2195_),
    .A1(_2194_),
    .B1(_2008_),
    .X(_2197_));
 sg13g2_inv_1 _6192_ (.Y(_2198_),
    .A(_2197_));
 sg13g2_o21ai_1 _6193_ (.B1(_2148_),
    .Y(_2199_),
    .A1(_2133_),
    .A2(_2197_));
 sg13g2_o21ai_1 _6194_ (.B1(_2137_),
    .Y(_2200_),
    .A1(_2193_),
    .A2(_2199_));
 sg13g2_xor2_1 _6195_ (.B(_2192_),
    .A(_2149_),
    .X(_2201_));
 sg13g2_xnor2_1 _6196_ (.Y(_2202_),
    .A(_2162_),
    .B(_2191_));
 sg13g2_xor2_1 _6197_ (.B(_2189_),
    .A(_2169_),
    .X(_2203_));
 sg13g2_xnor2_1 _6198_ (.Y(_2204_),
    .A(_2176_),
    .B(_2188_));
 sg13g2_nor2_1 _6199_ (.A(net474),
    .B(_2183_),
    .Y(_2205_));
 sg13g2_nor3_1 _6200_ (.A(_2184_),
    .B(_2187_),
    .C(_2205_),
    .Y(_2206_));
 sg13g2_a21oi_1 _6201_ (.A1(_2136_),
    .A2(_2197_),
    .Y(_2208_),
    .B1(_1607_));
 sg13g2_nand2b_1 _6202_ (.Y(_2209_),
    .B(_2148_),
    .A_N(_2137_));
 sg13g2_nand2_1 _6203_ (.Y(_2210_),
    .A(_2208_),
    .B(_2209_));
 sg13g2_nor4_1 _6204_ (.A(_2203_),
    .B(_2204_),
    .C(_2206_),
    .D(_2210_),
    .Y(_2211_));
 sg13g2_xnor2_1 _6205_ (.Y(_2212_),
    .A(_2135_),
    .B(_2161_));
 sg13g2_nand2_1 _6206_ (.Y(_2213_),
    .A(_2147_),
    .B(_2169_));
 sg13g2_nand2_1 _6207_ (.Y(_2214_),
    .A(_2168_),
    .B(_2213_));
 sg13g2_nand2_1 _6208_ (.Y(_2215_),
    .A(_2212_),
    .B(_2214_));
 sg13g2_xnor2_1 _6209_ (.Y(_2216_),
    .A(_2212_),
    .B(_2214_));
 sg13g2_nand2b_1 _6210_ (.Y(_2217_),
    .B(_2176_),
    .A_N(_2159_));
 sg13g2_and2_1 _6211_ (.A(_2175_),
    .B(_2217_),
    .X(_2219_));
 sg13g2_xnor2_1 _6212_ (.Y(_2220_),
    .A(_2147_),
    .B(_2169_));
 sg13g2_nand2_1 _6213_ (.Y(_2221_),
    .A(_2219_),
    .B(_2220_));
 sg13g2_o21ai_1 _6214_ (.B1(_2148_),
    .Y(_2222_),
    .A1(_2149_),
    .A2(_2198_));
 sg13g2_nor2_1 _6215_ (.A(_2137_),
    .B(_2222_),
    .Y(_2223_));
 sg13g2_xnor2_1 _6216_ (.Y(_2224_),
    .A(_2136_),
    .B(_2198_));
 sg13g2_o21ai_1 _6217_ (.B1(_1663_),
    .Y(_2225_),
    .A1(_2223_),
    .A2(_2224_));
 sg13g2_nor2_1 _6218_ (.A(net474),
    .B(_2173_),
    .Y(_2226_));
 sg13g2_nor2_1 _6219_ (.A(_2885_),
    .B(_2172_),
    .Y(_2227_));
 sg13g2_o21ai_1 _6220_ (.B1(_2183_),
    .Y(_2228_),
    .A1(_2226_),
    .A2(_2227_));
 sg13g2_xor2_1 _6221_ (.B(_2187_),
    .A(_2167_),
    .X(_2230_));
 sg13g2_xor2_1 _6222_ (.B(_2230_),
    .A(_2226_),
    .X(_2231_));
 sg13g2_nand2b_1 _6223_ (.Y(_2232_),
    .B(_2231_),
    .A_N(_2228_));
 sg13g2_xor2_1 _6224_ (.B(_2231_),
    .A(_2228_),
    .X(_2233_));
 sg13g2_o21ai_1 _6225_ (.B1(_2232_),
    .Y(_2234_),
    .A1(_2226_),
    .A2(_2230_));
 sg13g2_a21oi_2 _6226_ (.B1(_2181_),
    .Y(_2235_),
    .A2(_2186_),
    .A1(_2167_));
 sg13g2_xor2_1 _6227_ (.B(_2176_),
    .A(_2159_),
    .X(_2236_));
 sg13g2_nand2_1 _6228_ (.Y(_2237_),
    .A(_2235_),
    .B(_2236_));
 sg13g2_nor2_1 _6229_ (.A(_2235_),
    .B(_2236_),
    .Y(_2238_));
 sg13g2_xnor2_1 _6230_ (.Y(_2239_),
    .A(_2235_),
    .B(_2236_));
 sg13g2_a21o_1 _6231_ (.A2(_2162_),
    .A1(_2135_),
    .B1(_2160_),
    .X(_2241_));
 sg13g2_xor2_1 _6232_ (.B(_2197_),
    .A(_2149_),
    .X(_2242_));
 sg13g2_nor2b_1 _6233_ (.A(_2241_),
    .B_N(_2242_),
    .Y(_2243_));
 sg13g2_xnor2_1 _6234_ (.Y(_2244_),
    .A(_2241_),
    .B(_2242_));
 sg13g2_nand2_1 _6235_ (.Y(_2245_),
    .A(_2137_),
    .B(_2222_));
 sg13g2_nor2b_1 _6236_ (.A(_2223_),
    .B_N(_2245_),
    .Y(_2246_));
 sg13g2_nand2_1 _6237_ (.Y(_2247_),
    .A(_2242_),
    .B(_2246_));
 sg13g2_a21oi_1 _6238_ (.A1(_2215_),
    .A2(_2247_),
    .Y(_2248_),
    .B1(_2244_));
 sg13g2_nand2_1 _6239_ (.Y(_2249_),
    .A(_2224_),
    .B(_2245_));
 sg13g2_nand2_1 _6240_ (.Y(_2250_),
    .A(_2215_),
    .B(_2244_));
 sg13g2_a22oi_1 _6241_ (.Y(_2252_),
    .B1(_2250_),
    .B2(_2246_),
    .A2(_2249_),
    .A1(_2243_));
 sg13g2_o21ai_1 _6242_ (.B1(_2216_),
    .Y(_2253_),
    .A1(_2219_),
    .A2(_2220_));
 sg13g2_nor3_1 _6243_ (.A(_2234_),
    .B(_2238_),
    .C(_2253_),
    .Y(_2254_));
 sg13g2_a21o_1 _6244_ (.A2(_2239_),
    .A1(_2234_),
    .B1(_2254_),
    .X(_2255_));
 sg13g2_a21oi_1 _6245_ (.A1(_2237_),
    .A2(_2253_),
    .Y(_2256_),
    .B1(_2225_));
 sg13g2_xnor2_1 _6246_ (.Y(_2257_),
    .A(_2216_),
    .B(_2221_));
 sg13g2_nand3_1 _6247_ (.B(_2256_),
    .C(_2257_),
    .A(_2233_),
    .Y(_2258_));
 sg13g2_nor4_2 _6248_ (.A(_2248_),
    .B(_2252_),
    .C(_2255_),
    .Y(_2259_),
    .D(_2258_));
 sg13g2_and4_1 _6249_ (.A(_2200_),
    .B(_2201_),
    .C(_2202_),
    .D(_2211_),
    .X(_2260_));
 sg13g2_nor3_1 _6250_ (.A(_1956_),
    .B(_2259_),
    .C(_2260_),
    .Y(_2261_));
 sg13g2_nand3_1 _6251_ (.B(_1669_),
    .C(_2261_),
    .A(_1616_),
    .Y(_2263_));
 sg13g2_or2_1 _6252_ (.X(_2264_),
    .B(_2180_),
    .A(_1274_));
 sg13g2_xnor2_1 _6253_ (.Y(_2265_),
    .A(_1274_),
    .B(_2180_));
 sg13g2_or2_1 _6254_ (.X(_2266_),
    .B(_2265_),
    .A(_2167_));
 sg13g2_xnor2_1 _6255_ (.Y(_2267_),
    .A(_2167_),
    .B(_2265_));
 sg13g2_xor2_1 _6256_ (.B(_2183_),
    .A(_1282_),
    .X(_2268_));
 sg13g2_nor2_1 _6257_ (.A(_2173_),
    .B(_2268_),
    .Y(_2269_));
 sg13g2_a21oi_1 _6258_ (.A1(_1284_),
    .A2(_2183_),
    .Y(_2270_),
    .B1(_2269_));
 sg13g2_nor2_1 _6259_ (.A(_2267_),
    .B(_2270_),
    .Y(_2271_));
 sg13g2_xnor2_1 _6260_ (.Y(_2272_),
    .A(net462),
    .B(_2173_));
 sg13g2_nand2b_1 _6261_ (.Y(_2274_),
    .B(_2159_),
    .A_N(_2272_));
 sg13g2_xor2_1 _6262_ (.B(_2272_),
    .A(_2159_),
    .X(_2275_));
 sg13g2_a21oi_1 _6263_ (.A1(_2264_),
    .A2(_2266_),
    .Y(_2276_),
    .B1(_2275_));
 sg13g2_or2_1 _6264_ (.X(_2277_),
    .B(_2276_),
    .A(_2271_));
 sg13g2_o21ai_1 _6265_ (.B1(_2274_),
    .Y(_2278_),
    .A1(net462),
    .A2(_2173_));
 sg13g2_nor2_1 _6266_ (.A(_1234_),
    .B(_2167_),
    .Y(_2279_));
 sg13g2_xnor2_1 _6267_ (.Y(_2280_),
    .A(_1233_),
    .B(_2167_));
 sg13g2_xnor2_1 _6268_ (.Y(_2281_),
    .A(_2147_),
    .B(_2280_));
 sg13g2_nand2_1 _6269_ (.Y(_2282_),
    .A(_2278_),
    .B(_2281_));
 sg13g2_xnor2_1 _6270_ (.Y(_2283_),
    .A(_2278_),
    .B(_2281_));
 sg13g2_and3_1 _6271_ (.X(_2285_),
    .A(_2264_),
    .B(_2266_),
    .C(_2275_));
 sg13g2_nor2_1 _6272_ (.A(_2283_),
    .B(_2285_),
    .Y(_2286_));
 sg13g2_nand2_1 _6273_ (.Y(_2287_),
    .A(_2271_),
    .B(_2276_));
 sg13g2_nand2b_1 _6274_ (.Y(_2288_),
    .B(_2285_),
    .A_N(_2271_));
 sg13g2_xnor2_1 _6275_ (.Y(_2289_),
    .A(_2267_),
    .B(_2270_));
 sg13g2_and2_1 _6276_ (.A(_2173_),
    .B(_2268_),
    .X(_2290_));
 sg13g2_o21ai_1 _6277_ (.B1(_2289_),
    .Y(_2291_),
    .A1(_2269_),
    .A2(_2290_));
 sg13g2_nand3_1 _6278_ (.B(net464),
    .C(_1308_),
    .A(net466),
    .Y(_2292_));
 sg13g2_a21oi_1 _6279_ (.A1(_0053_),
    .A2(_3244_),
    .Y(_2293_),
    .B1(_3237_));
 sg13g2_nor4_2 _6280_ (.A(net583),
    .B(_0310_),
    .C(_2159_),
    .Y(_2294_),
    .D(_2293_));
 sg13g2_nand4_1 _6281_ (.B(_2147_),
    .C(_2197_),
    .A(_2135_),
    .Y(_2296_),
    .D(_2294_));
 sg13g2_nor3_1 _6282_ (.A(_2279_),
    .B(_2292_),
    .C(_2296_),
    .Y(_2297_));
 sg13g2_nand4_1 _6283_ (.B(_2288_),
    .C(_2291_),
    .A(_2282_),
    .Y(_2298_),
    .D(_2297_));
 sg13g2_a221oi_1 _6284_ (.B2(_2283_),
    .C1(_2298_),
    .B1(_2287_),
    .A1(_2277_),
    .Y(_2299_),
    .A2(_2286_));
 sg13g2_nand2_1 _6285_ (.Y(_2300_),
    .A(_1275_),
    .B(_1579_));
 sg13g2_xnor2_1 _6286_ (.Y(_2301_),
    .A(_1275_),
    .B(_1579_));
 sg13g2_xnor2_1 _6287_ (.Y(_2302_),
    .A(_1565_),
    .B(_2301_));
 sg13g2_nand2_1 _6288_ (.Y(_2303_),
    .A(_1284_),
    .B(_1584_));
 sg13g2_xnor2_1 _6289_ (.Y(_2304_),
    .A(_1282_),
    .B(_1583_));
 sg13g2_nand2b_1 _6290_ (.Y(_2305_),
    .B(_1573_),
    .A_N(_2304_));
 sg13g2_o21ai_1 _6291_ (.B1(_2300_),
    .Y(_2307_),
    .A1(_1565_),
    .A2(_2301_));
 sg13g2_nand2b_1 _6292_ (.Y(_2308_),
    .B(_1573_),
    .A_N(net462));
 sg13g2_xnor2_1 _6293_ (.Y(_2309_),
    .A(net461),
    .B(_1574_));
 sg13g2_xnor2_1 _6294_ (.Y(_2310_),
    .A(_1553_),
    .B(_2309_));
 sg13g2_nor2_1 _6295_ (.A(_2307_),
    .B(_2310_),
    .Y(_2311_));
 sg13g2_o21ai_1 _6296_ (.B1(_2308_),
    .Y(_2312_),
    .A1(_1552_),
    .A2(_2309_));
 sg13g2_nor2_1 _6297_ (.A(_1234_),
    .B(_1565_),
    .Y(_2313_));
 sg13g2_nor2_1 _6298_ (.A(_1233_),
    .B(_1564_),
    .Y(_2314_));
 sg13g2_o21ai_1 _6299_ (.B1(_1540_),
    .Y(_2315_),
    .A1(_2313_),
    .A2(_2314_));
 sg13g2_nor2_1 _6300_ (.A(_2312_),
    .B(_2315_),
    .Y(_2316_));
 sg13g2_nor2_1 _6301_ (.A(_2311_),
    .B(_2316_),
    .Y(_2318_));
 sg13g2_or2_1 _6302_ (.X(_2319_),
    .B(_2316_),
    .A(_2311_));
 sg13g2_xnor2_1 _6303_ (.Y(_2320_),
    .A(_1573_),
    .B(_2304_));
 sg13g2_a221oi_1 _6304_ (.B2(_2320_),
    .C1(_2302_),
    .B1(_2319_),
    .A1(_2303_),
    .Y(_2321_),
    .A2(_2305_));
 sg13g2_nand2_1 _6305_ (.Y(_2322_),
    .A(_2307_),
    .B(_2310_));
 sg13g2_a221oi_1 _6306_ (.B2(_2322_),
    .C1(_2302_),
    .B1(_2316_),
    .A1(_2303_),
    .Y(_2323_),
    .A2(_2305_));
 sg13g2_a21oi_1 _6307_ (.A1(_2318_),
    .A2(_2322_),
    .Y(_2324_),
    .B1(_2323_));
 sg13g2_nand2_1 _6308_ (.Y(_2325_),
    .A(_2312_),
    .B(_2315_));
 sg13g2_nor3_1 _6309_ (.A(net602),
    .B(net605),
    .C(_0016_),
    .Y(_2326_));
 sg13g2_a21oi_1 _6310_ (.A1(net608),
    .A2(_2326_),
    .Y(_2327_),
    .B1(_1034_));
 sg13g2_nor4_2 _6311_ (.A(net537),
    .B(net529),
    .C(_0332_),
    .Y(_2329_),
    .D(_2327_));
 sg13g2_nor4_2 _6312_ (.A(_0310_),
    .B(_0321_),
    .C(_1553_),
    .Y(_2330_),
    .D(_2329_));
 sg13g2_nand4_1 _6313_ (.B(_1595_),
    .C(_1599_),
    .A(_1540_),
    .Y(_2331_),
    .D(_2330_));
 sg13g2_nor3_1 _6314_ (.A(_2292_),
    .B(_2313_),
    .C(_2331_),
    .Y(_2332_));
 sg13g2_nand4_1 _6315_ (.B(_1574_),
    .C(_1583_),
    .A(_1282_),
    .Y(_2333_),
    .D(_2302_));
 sg13g2_nand3_1 _6316_ (.B(_2332_),
    .C(_2333_),
    .A(_2325_),
    .Y(_2334_));
 sg13g2_nand3_1 _6317_ (.B(_0279_),
    .C(_0301_),
    .A(_0278_),
    .Y(_2335_));
 sg13g2_nand2b_1 _6318_ (.Y(_2336_),
    .B(_2335_),
    .A_N(_0281_));
 sg13g2_a21oi_2 _6319_ (.B1(_0298_),
    .Y(_2337_),
    .A2(_2336_),
    .A1(_0303_));
 sg13g2_nor3_1 _6320_ (.A(_2321_),
    .B(_2324_),
    .C(_2334_),
    .Y(_2338_));
 sg13g2_or4_1 _6321_ (.A(_1342_),
    .B(_2263_),
    .C(_2299_),
    .D(_2338_),
    .X(_2340_));
 sg13g2_nor3_2 _6322_ (.A(_0296_),
    .B(_0305_),
    .C(_2337_),
    .Y(_2341_));
 sg13g2_nor4_1 _6323_ (.A(_1329_),
    .B(_1337_),
    .C(_2340_),
    .D(_2341_),
    .Y(_2342_));
 sg13g2_and3_2 _6324_ (.X(_2343_),
    .A(_0703_),
    .B(_1040_),
    .C(_2342_));
 sg13g2_o21ai_1 _6325_ (.B1(net583),
    .Y(_2344_),
    .A1(net585),
    .A2(net588));
 sg13g2_nand3_1 _6326_ (.B(_0217_),
    .C(_2943_),
    .A(_0206_),
    .Y(_2345_));
 sg13g2_or2_1 _6327_ (.X(_2346_),
    .B(_0309_),
    .A(_2982_));
 sg13g2_nand4_1 _6328_ (.B(_2344_),
    .C(_2345_),
    .A(_2971_),
    .Y(_2347_),
    .D(_2346_));
 sg13g2_a21oi_2 _6329_ (.B1(_2347_),
    .Y(uo_out[6]),
    .A2(_2343_),
    .A1(_0308_));
 sg13g2_nor2_2 _6330_ (.A(_3250_),
    .B(_2343_),
    .Y(uo_out[5]));
 sg13g2_a21oi_2 _6331_ (.B1(_3250_),
    .Y(uo_out[2]),
    .A2(_2343_),
    .A1(_0307_));
 sg13g2_nor2_1 _6332_ (.A(net610),
    .B(_0375_),
    .Y(_0020_));
 sg13g2_o21ai_1 _6333_ (.B1(net1),
    .Y(_2349_),
    .A1(net551),
    .A2(net605));
 sg13g2_a21oi_1 _6334_ (.A1(net551),
    .A2(_2619_),
    .Y(_0021_),
    .B1(_2349_));
 sg13g2_nand2_2 _6335_ (.Y(_2350_),
    .A(_2617_),
    .B(_0368_));
 sg13g2_nor4_2 _6336_ (.A(_0042_),
    .B(_2587_),
    .C(_0313_),
    .Y(_2351_),
    .D(_2350_));
 sg13g2_nand2_1 _6337_ (.Y(_2352_),
    .A(net548),
    .B(_2351_));
 sg13g2_inv_1 _6338_ (.Y(_2353_),
    .A(net526));
 sg13g2_nor2b_1 _6339_ (.A(net42),
    .B_N(_2617_),
    .Y(_2354_));
 sg13g2_xnor2_1 _6340_ (.Y(_2355_),
    .A(net42),
    .B(_2617_));
 sg13g2_nor2_1 _6341_ (.A(net542),
    .B(_2355_),
    .Y(_2357_));
 sg13g2_nor4_1 _6342_ (.A(net610),
    .B(_1365_),
    .C(_2353_),
    .D(_2357_),
    .Y(_0022_));
 sg13g2_nor2_2 _6343_ (.A(net539),
    .B(_2351_),
    .Y(_2358_));
 sg13g2_xnor2_1 _6344_ (.Y(_2359_),
    .A(net49),
    .B(_2354_));
 sg13g2_a22oi_1 _6345_ (.Y(_2360_),
    .B1(_2358_),
    .B2(_2359_),
    .A2(net599),
    .A1(net542));
 sg13g2_nor2_1 _6346_ (.A(net610),
    .B(net50),
    .Y(_0023_));
 sg13g2_nor2_1 _6347_ (.A(_0015_),
    .B(_2350_),
    .Y(_2361_));
 sg13g2_xnor2_1 _6348_ (.Y(_2362_),
    .A(_3191_),
    .B(_2350_));
 sg13g2_a22oi_1 _6349_ (.Y(_2363_),
    .B1(_2358_),
    .B2(_2362_),
    .A2(net597),
    .A1(net542));
 sg13g2_nor2_1 _6350_ (.A(net610),
    .B(_2363_),
    .Y(_0024_));
 sg13g2_xnor2_1 _6351_ (.Y(_2365_),
    .A(net592),
    .B(_2361_));
 sg13g2_a22oi_1 _6352_ (.Y(_2366_),
    .B1(_2358_),
    .B2(_2365_),
    .A2(net593),
    .A1(net539));
 sg13g2_nor2_1 _6353_ (.A(net609),
    .B(_2366_),
    .Y(_0025_));
 sg13g2_nor3_2 _6354_ (.A(net589),
    .B(_0097_),
    .C(_2350_),
    .Y(_2367_));
 sg13g2_o21ai_1 _6355_ (.B1(net589),
    .Y(_2368_),
    .A1(_0097_),
    .A2(_2350_));
 sg13g2_nor2b_1 _6356_ (.A(_2367_),
    .B_N(_2368_),
    .Y(_2369_));
 sg13g2_a22oi_1 _6357_ (.Y(_2370_),
    .B1(_2358_),
    .B2(_2369_),
    .A2(net591),
    .A1(net542));
 sg13g2_nor2_1 _6358_ (.A(net610),
    .B(_2370_),
    .Y(_0026_));
 sg13g2_xnor2_1 _6359_ (.Y(_2371_),
    .A(net45),
    .B(_2367_));
 sg13g2_a22oi_1 _6360_ (.Y(_2372_),
    .B1(_2358_),
    .B2(_2371_),
    .A2(net587),
    .A1(net540));
 sg13g2_nor2_1 _6361_ (.A(net609),
    .B(_2372_),
    .Y(_0027_));
 sg13g2_o21ai_1 _6362_ (.B1(_0013_),
    .Y(_2374_),
    .A1(_0130_),
    .A2(_2350_));
 sg13g2_nor3_1 _6363_ (.A(_0013_),
    .B(_0130_),
    .C(_2350_),
    .Y(_2375_));
 sg13g2_nor2b_1 _6364_ (.A(_2375_),
    .B_N(_2358_),
    .Y(_2376_));
 sg13g2_a22oi_1 _6365_ (.Y(_2377_),
    .B1(_2374_),
    .B2(_2376_),
    .A2(net584),
    .A1(net539));
 sg13g2_nor2_1 _6366_ (.A(net609),
    .B(_2377_),
    .Y(_0028_));
 sg13g2_xnor2_1 _6367_ (.Y(_2378_),
    .A(net51),
    .B(_2375_));
 sg13g2_nand2_1 _6368_ (.Y(_2379_),
    .A(_2358_),
    .B(_2378_));
 sg13g2_a21oi_1 _6369_ (.A1(_1716_),
    .A2(_2379_),
    .Y(_0029_),
    .B1(net609));
 sg13g2_nor3_1 _6370_ (.A(_2971_),
    .B(net563),
    .C(_0414_),
    .Y(_2380_));
 sg13g2_nand4_1 _6371_ (.B(_0348_),
    .C(_0370_),
    .A(_0249_),
    .Y(_2382_),
    .D(_2380_));
 sg13g2_nor2b_2 _6372_ (.A(_2352_),
    .B_N(_2382_),
    .Y(_2383_));
 sg13g2_a22oi_1 _6373_ (.Y(_2384_),
    .B1(_2383_),
    .B2(net48),
    .A2(net526),
    .A1(net579));
 sg13g2_nor2_1 _6374_ (.A(net609),
    .B(_2384_),
    .Y(_0030_));
 sg13g2_a21oi_1 _6375_ (.A1(net579),
    .A2(_2353_),
    .Y(_2385_),
    .B1(net578));
 sg13g2_o21ai_1 _6376_ (.B1(net1),
    .Y(_2386_),
    .A1(_3255_),
    .A2(net526));
 sg13g2_nor2_1 _6377_ (.A(_2385_),
    .B(_2386_),
    .Y(_0031_));
 sg13g2_a22oi_1 _6378_ (.Y(_2387_),
    .B1(_2383_),
    .B2(_0057_),
    .A2(net526),
    .A1(net573));
 sg13g2_nor2_1 _6379_ (.A(net610),
    .B(_2387_),
    .Y(_0032_));
 sg13g2_nor2_1 _6380_ (.A(net54),
    .B(_3255_),
    .Y(_2388_));
 sg13g2_xnor2_1 _6381_ (.Y(_2390_),
    .A(_3037_),
    .B(_2388_));
 sg13g2_a22oi_1 _6382_ (.Y(_2391_),
    .B1(_2383_),
    .B2(_2390_),
    .A2(net526),
    .A1(net572));
 sg13g2_nor2_1 _6383_ (.A(net609),
    .B(net55),
    .Y(_0033_));
 sg13g2_nand2_1 _6384_ (.Y(_2392_),
    .A(net572),
    .B(_0056_));
 sg13g2_or2_2 _6385_ (.X(_2393_),
    .B(_2392_),
    .A(net526));
 sg13g2_o21ai_1 _6386_ (.B1(net1),
    .Y(_2394_),
    .A1(_3026_),
    .A2(_2393_));
 sg13g2_a21oi_1 _6387_ (.A1(_3026_),
    .A2(_2393_),
    .Y(_0034_),
    .B1(_2394_));
 sg13g2_nor2_1 _6388_ (.A(net56),
    .B(_2393_),
    .Y(_2395_));
 sg13g2_o21ai_1 _6389_ (.B1(net1),
    .Y(_2396_),
    .A1(net565),
    .A2(_2395_));
 sg13g2_a21oi_1 _6390_ (.A1(net566),
    .A2(_2395_),
    .Y(_0035_),
    .B1(_2396_));
 sg13g2_o21ai_1 _6391_ (.B1(_3004_),
    .Y(_2398_),
    .A1(_2937_),
    .A2(_2393_));
 sg13g2_o21ai_1 _6392_ (.B1(net1),
    .Y(_2399_),
    .A1(_2938_),
    .A2(_2393_));
 sg13g2_nor2b_1 _6393_ (.A(_2399_),
    .B_N(_2398_),
    .Y(_0036_));
 sg13g2_nor3_1 _6394_ (.A(_0007_),
    .B(net532),
    .C(_2392_),
    .Y(_2400_));
 sg13g2_xnor2_1 _6395_ (.Y(_2401_),
    .A(_0005_),
    .B(_2400_));
 sg13g2_a22oi_1 _6396_ (.Y(_2402_),
    .B1(_2383_),
    .B2(_2401_),
    .A2(net526),
    .A1(net46));
 sg13g2_nor2_1 _6397_ (.A(net609),
    .B(_2402_),
    .Y(_0037_));
 sg13g2_nor2_1 _6398_ (.A(_2940_),
    .B(_2393_),
    .Y(_2403_));
 sg13g2_o21ai_1 _6399_ (.B1(net1),
    .Y(_2404_),
    .A1(net564),
    .A2(_2403_));
 sg13g2_a21oi_1 _6400_ (.A1(net564),
    .A2(_2403_),
    .Y(_0038_),
    .B1(_2404_));
 sg13g2_nor3_1 _6401_ (.A(net562),
    .B(_2940_),
    .C(_2392_),
    .Y(_2406_));
 sg13g2_xnor2_1 _6402_ (.Y(_2407_),
    .A(net561),
    .B(_2406_));
 sg13g2_a22oi_1 _6403_ (.Y(_2408_),
    .B1(_2383_),
    .B2(_2407_),
    .A2(net526),
    .A1(net44));
 sg13g2_nor2_1 _6404_ (.A(net609),
    .B(_2408_),
    .Y(_0039_));
 sg13g2_and2_1 _6405_ (.A(net40),
    .B(net1),
    .X(_0040_));
 sg13g2_nor2_1 _6406_ (.A(_1234_),
    .B(net463),
    .Y(_2409_));
 sg13g2_nand2_1 _6407_ (.Y(_2410_),
    .A(net467),
    .B(_1275_));
 sg13g2_xor2_1 _6408_ (.B(net461),
    .A(net465),
    .X(_2411_));
 sg13g2_nand2b_1 _6409_ (.Y(_2412_),
    .B(_2411_),
    .A_N(_2410_));
 sg13g2_o21ai_1 _6410_ (.B1(_2412_),
    .Y(_2413_),
    .A1(net465),
    .A2(net461));
 sg13g2_nand2_1 _6411_ (.Y(_2415_),
    .A(_1234_),
    .B(net463));
 sg13g2_nand2b_1 _6412_ (.Y(_2416_),
    .B(_2415_),
    .A_N(_2409_));
 sg13g2_a21o_1 _6413_ (.A2(_2415_),
    .A1(_2413_),
    .B1(_2409_),
    .X(_2417_));
 sg13g2_xor2_1 _6414_ (.B(_1307_),
    .A(net465),
    .X(_2418_));
 sg13g2_nand2b_1 _6415_ (.Y(_2419_),
    .B(_2417_),
    .A_N(_2418_));
 sg13g2_o21ai_1 _6416_ (.B1(_2419_),
    .Y(_2420_),
    .A1(net465),
    .A2(_1308_));
 sg13g2_xnor2_1 _6417_ (.Y(_2421_),
    .A(net463),
    .B(_2420_));
 sg13g2_nand2_1 _6418_ (.Y(_2422_),
    .A(_0966_),
    .B(_2421_));
 sg13g2_a22oi_1 _6419_ (.Y(_2423_),
    .B1(_2420_),
    .B2(_1309_),
    .A2(_2419_),
    .A1(_1308_));
 sg13g2_xnor2_1 _6420_ (.Y(_2424_),
    .A(_0944_),
    .B(_2423_));
 sg13g2_xor2_1 _6421_ (.B(_2418_),
    .A(_2417_),
    .X(_2426_));
 sg13g2_nor2b_1 _6422_ (.A(_2426_),
    .B_N(_0976_),
    .Y(_2427_));
 sg13g2_xnor2_1 _6423_ (.Y(_2428_),
    .A(_2413_),
    .B(_2416_));
 sg13g2_nor2b_1 _6424_ (.A(_0984_),
    .B_N(_2428_),
    .Y(_2429_));
 sg13g2_nand2b_1 _6425_ (.Y(_2430_),
    .B(_2426_),
    .A_N(_0976_));
 sg13g2_a221oi_1 _6426_ (.B2(_2430_),
    .C1(_2427_),
    .B1(_2429_),
    .A1(_2422_),
    .Y(_2431_),
    .A2(_2424_));
 sg13g2_nor2_1 _6427_ (.A(_0966_),
    .B(_2421_),
    .Y(_2432_));
 sg13g2_nand2_1 _6428_ (.Y(_2433_),
    .A(_2427_),
    .B(_2429_));
 sg13g2_nor2_1 _6429_ (.A(_2432_),
    .B(_2433_),
    .Y(_2434_));
 sg13g2_a21oi_1 _6430_ (.A1(_2422_),
    .A2(_2434_),
    .Y(_2435_),
    .B1(_2431_));
 sg13g2_nor2_1 _6431_ (.A(_2424_),
    .B(_2432_),
    .Y(_2437_));
 sg13g2_nor2_1 _6432_ (.A(_2429_),
    .B(_2430_),
    .Y(_2438_));
 sg13g2_xnor2_1 _6433_ (.Y(_2439_),
    .A(_0984_),
    .B(_2428_));
 sg13g2_xnor2_1 _6434_ (.Y(_2440_),
    .A(_2410_),
    .B(_2411_));
 sg13g2_nor2_1 _6435_ (.A(_1001_),
    .B(_2440_),
    .Y(_2441_));
 sg13g2_xnor2_1 _6436_ (.Y(_2442_),
    .A(net467),
    .B(_1275_));
 sg13g2_nor2_1 _6437_ (.A(net496),
    .B(_0982_),
    .Y(_2443_));
 sg13g2_nor3_1 _6438_ (.A(_0768_),
    .B(_0797_),
    .C(_0870_),
    .Y(_2444_));
 sg13g2_a21oi_1 _6439_ (.A1(_0870_),
    .A2(_0906_),
    .Y(_2445_),
    .B1(_2444_));
 sg13g2_a21oi_1 _6440_ (.A1(net496),
    .A2(_2445_),
    .Y(_2446_),
    .B1(_2443_));
 sg13g2_nor2_1 _6441_ (.A(_0758_),
    .B(_0961_),
    .Y(_2448_));
 sg13g2_a21oi_1 _6442_ (.A1(_0801_),
    .A2(_2446_),
    .Y(_2449_),
    .B1(_2448_));
 sg13g2_nor3_1 _6443_ (.A(_2441_),
    .B(_2442_),
    .C(_2449_),
    .Y(_2450_));
 sg13g2_a21o_1 _6444_ (.A2(_2440_),
    .A1(_1001_),
    .B1(_2450_),
    .X(_2451_));
 sg13g2_xnor2_1 _6445_ (.Y(_2452_),
    .A(_1001_),
    .B(_2440_));
 sg13g2_nand2_1 _6446_ (.Y(_2453_),
    .A(_2442_),
    .B(_2449_));
 sg13g2_nand2b_1 _6447_ (.Y(_2454_),
    .B(_2453_),
    .A_N(_2452_));
 sg13g2_nand2b_1 _6448_ (.Y(_2455_),
    .B(_2452_),
    .A_N(_2453_));
 sg13g2_nor2_1 _6449_ (.A(_0321_),
    .B(_0329_),
    .Y(_2456_));
 sg13g2_nand3_1 _6450_ (.B(_0333_),
    .C(_0363_),
    .A(_2627_),
    .Y(_2457_));
 sg13g2_nand2_2 _6451_ (.Y(_2459_),
    .A(_2456_),
    .B(_2457_));
 sg13g2_nor2_1 _6452_ (.A(_0260_),
    .B(_0832_),
    .Y(_2460_));
 sg13g2_a21oi_1 _6453_ (.A1(net580),
    .A2(_0217_),
    .Y(_2461_),
    .B1(_0832_));
 sg13g2_o21ai_1 _6454_ (.B1(_0249_),
    .Y(_2462_),
    .A1(net532),
    .A2(_2461_));
 sg13g2_o21ai_1 _6455_ (.B1(_2462_),
    .Y(_2463_),
    .A1(net563),
    .A2(_2460_));
 sg13g2_nand2_2 _6456_ (.Y(_2464_),
    .A(net561),
    .B(_2463_));
 sg13g2_a21oi_2 _6457_ (.B1(_2464_),
    .Y(_2465_),
    .A2(net529),
    .A1(_0322_));
 sg13g2_nand4_1 _6458_ (.B(_2455_),
    .C(_2459_),
    .A(_2454_),
    .Y(_2466_),
    .D(_2465_));
 sg13g2_a21oi_1 _6459_ (.A1(_2439_),
    .A2(_2451_),
    .Y(_2467_),
    .B1(_2466_));
 sg13g2_o21ai_1 _6460_ (.B1(_2467_),
    .Y(_2468_),
    .A1(_2439_),
    .A2(_2451_));
 sg13g2_or4_2 _6461_ (.A(_2435_),
    .B(_2437_),
    .C(_2438_),
    .D(_2468_),
    .X(_2470_));
 sg13g2_nand2_1 _6462_ (.Y(_2471_),
    .A(_0256_),
    .B(_2426_));
 sg13g2_nor2_1 _6463_ (.A(_0256_),
    .B(_2426_),
    .Y(_2472_));
 sg13g2_nand2_1 _6464_ (.Y(_2473_),
    .A(_0264_),
    .B(_2428_));
 sg13g2_xnor2_1 _6465_ (.Y(_2474_),
    .A(_0264_),
    .B(_2428_));
 sg13g2_nand2b_1 _6466_ (.Y(_2475_),
    .B(net469),
    .A_N(_2440_));
 sg13g2_nor2b_1 _6467_ (.A(net469),
    .B_N(_2440_),
    .Y(_2476_));
 sg13g2_nor2_1 _6468_ (.A(_0277_),
    .B(_2442_),
    .Y(_2477_));
 sg13g2_a21oi_1 _6469_ (.A1(_2475_),
    .A2(_2477_),
    .Y(_2478_),
    .B1(_2476_));
 sg13g2_nor2_1 _6470_ (.A(_2474_),
    .B(_2478_),
    .Y(_2479_));
 sg13g2_inv_1 _6471_ (.Y(_2481_),
    .A(_2479_));
 sg13g2_nand2_1 _6472_ (.Y(_2482_),
    .A(_2473_),
    .B(_2481_));
 sg13g2_a21oi_1 _6473_ (.A1(_2471_),
    .A2(_2482_),
    .Y(_2483_),
    .B1(_2472_));
 sg13g2_xnor2_1 _6474_ (.Y(_2484_),
    .A(_0232_),
    .B(_2423_));
 sg13g2_nand2_1 _6475_ (.Y(_2485_),
    .A(_0248_),
    .B(_2421_));
 sg13g2_nand3b_1 _6476_ (.B(_2485_),
    .C(_2483_),
    .Y(_2486_),
    .A_N(_2484_));
 sg13g2_or2_1 _6477_ (.X(_2487_),
    .B(_2421_),
    .A(_0248_));
 sg13g2_a21o_1 _6478_ (.A2(_2487_),
    .A1(_2485_),
    .B1(_2483_),
    .X(_2488_));
 sg13g2_xnor2_1 _6479_ (.Y(_2489_),
    .A(_0256_),
    .B(_2426_));
 sg13g2_xnor2_1 _6480_ (.Y(_2490_),
    .A(net469),
    .B(_2440_));
 sg13g2_inv_1 _6481_ (.Y(_2492_),
    .A(_2490_));
 sg13g2_and2_1 _6482_ (.A(_0277_),
    .B(_2442_),
    .X(_2493_));
 sg13g2_nand2b_1 _6483_ (.Y(_2494_),
    .B(_2490_),
    .A_N(_2493_));
 sg13g2_nor3_2 _6484_ (.A(_3092_),
    .B(_3114_),
    .C(_0097_),
    .Y(_2495_));
 sg13g2_o21ai_1 _6485_ (.B1(net586),
    .Y(_2496_),
    .A1(net588),
    .A2(_2495_));
 sg13g2_a221oi_1 _6486_ (.B2(_0019_),
    .C1(_2464_),
    .B1(_2496_),
    .A1(_2492_),
    .Y(_2497_),
    .A2(_2493_));
 sg13g2_nand3_1 _6487_ (.B(_2494_),
    .C(_2497_),
    .A(_2481_),
    .Y(_2498_));
 sg13g2_a21oi_1 _6488_ (.A1(_2474_),
    .A2(_2478_),
    .Y(_2499_),
    .B1(_2498_));
 sg13g2_o21ai_1 _6489_ (.B1(_2499_),
    .Y(_2500_),
    .A1(_2473_),
    .A2(_2489_));
 sg13g2_a21oi_1 _6490_ (.A1(_2473_),
    .A2(_2489_),
    .Y(_2501_),
    .B1(_2500_));
 sg13g2_o21ai_1 _6491_ (.B1(_2484_),
    .Y(_2503_),
    .A1(_0248_),
    .A2(_2421_));
 sg13g2_nand4_1 _6492_ (.B(_2488_),
    .C(_2501_),
    .A(_2486_),
    .Y(_2504_),
    .D(_2503_));
 sg13g2_or2_1 _6493_ (.X(_2505_),
    .B(net463),
    .A(_0615_));
 sg13g2_xor2_1 _6494_ (.B(net463),
    .A(_0615_),
    .X(_2506_));
 sg13g2_nor2_1 _6495_ (.A(_0642_),
    .B(net465),
    .Y(_2507_));
 sg13g2_xnor2_1 _6496_ (.Y(_2508_),
    .A(_0629_),
    .B(_1308_));
 sg13g2_o21ai_1 _6497_ (.B1(_2505_),
    .Y(_2509_),
    .A1(_0619_),
    .A2(_1307_));
 sg13g2_mux2_1 _6498_ (.A0(_2509_),
    .A1(net463),
    .S(_2508_),
    .X(_2510_));
 sg13g2_nor2_1 _6499_ (.A(_2507_),
    .B(_2510_),
    .Y(_2511_));
 sg13g2_o21ai_1 _6500_ (.B1(_0619_),
    .Y(_2512_),
    .A1(_0629_),
    .A2(_1307_));
 sg13g2_a21oi_1 _6501_ (.A1(_2610_),
    .A2(_2627_),
    .Y(_2514_),
    .B1(_0727_));
 sg13g2_nor3_1 _6502_ (.A(_2642_),
    .B(_2651_),
    .C(_2514_),
    .Y(_2515_));
 sg13g2_o21ai_1 _6503_ (.B1(_1035_),
    .Y(_2516_),
    .A1(_1033_),
    .A2(_2515_));
 sg13g2_a21o_1 _6504_ (.A2(_2516_),
    .A1(_1032_),
    .B1(_0321_),
    .X(_2517_));
 sg13g2_nor2_1 _6505_ (.A(_0653_),
    .B(_1234_),
    .Y(_2518_));
 sg13g2_xor2_1 _6506_ (.B(net467),
    .A(_0653_),
    .X(_2519_));
 sg13g2_or2_1 _6507_ (.X(_2520_),
    .B(net461),
    .A(_0669_));
 sg13g2_nand2_1 _6508_ (.Y(_2521_),
    .A(_0614_),
    .B(_0650_));
 sg13g2_a21oi_1 _6509_ (.A1(net492),
    .A2(_0572_),
    .Y(_2522_),
    .B1(net489));
 sg13g2_a22oi_1 _6510_ (.Y(_2523_),
    .B1(_2521_),
    .B2(_2522_),
    .A2(_0611_),
    .A1(net489));
 sg13g2_nand2_1 _6511_ (.Y(_2525_),
    .A(_0669_),
    .B(net461));
 sg13g2_nand3_1 _6512_ (.B(_2523_),
    .C(_2525_),
    .A(_1275_),
    .Y(_2526_));
 sg13g2_nand2_1 _6513_ (.Y(_2527_),
    .A(_2520_),
    .B(_2526_));
 sg13g2_nand3b_1 _6514_ (.B(_1274_),
    .C(_2520_),
    .Y(_2528_),
    .A_N(_2523_));
 sg13g2_a21oi_1 _6515_ (.A1(_2525_),
    .A2(_2528_),
    .Y(_2529_),
    .B1(_2519_));
 sg13g2_a21o_1 _6516_ (.A2(_2527_),
    .A1(_2519_),
    .B1(_2529_),
    .X(_2530_));
 sg13g2_xnor2_1 _6517_ (.Y(_2531_),
    .A(_0642_),
    .B(net465));
 sg13g2_xnor2_1 _6518_ (.Y(_2532_),
    .A(_2518_),
    .B(_2531_));
 sg13g2_nand4_1 _6519_ (.B(_2517_),
    .C(_2530_),
    .A(_2512_),
    .Y(_2533_),
    .D(_2532_));
 sg13g2_nand2_1 _6520_ (.Y(_2534_),
    .A(_2507_),
    .B(_2508_));
 sg13g2_a21oi_1 _6521_ (.A1(_2506_),
    .A2(_2534_),
    .Y(_2536_),
    .B1(_2533_));
 sg13g2_o21ai_1 _6522_ (.B1(_2536_),
    .Y(_2537_),
    .A1(_2506_),
    .A2(_2511_));
 sg13g2_nand3_1 _6523_ (.B(_1582_),
    .C(_1583_),
    .A(_2885_),
    .Y(_2538_));
 sg13g2_nand3_1 _6524_ (.B(_0339_),
    .C(_1347_),
    .A(_0333_),
    .Y(_2539_));
 sg13g2_nand3_1 _6525_ (.B(_2456_),
    .C(_2539_),
    .A(_0323_),
    .Y(_2540_));
 sg13g2_nand4_1 _6526_ (.B(_2465_),
    .C(_2538_),
    .A(_1585_),
    .Y(_2541_),
    .D(_2540_));
 sg13g2_nor2_1 _6527_ (.A(_1593_),
    .B(_2541_),
    .Y(_2542_));
 sg13g2_nand4_1 _6528_ (.B(_1592_),
    .C(_1594_),
    .A(_1590_),
    .Y(_2543_),
    .D(_2542_));
 sg13g2_mux2_1 _6529_ (.A0(_2184_),
    .A1(_2205_),
    .S(_2187_),
    .X(_2544_));
 sg13g2_nand2_1 _6530_ (.Y(_2545_),
    .A(net537),
    .B(_1718_));
 sg13g2_a21oi_1 _6531_ (.A1(_2613_),
    .A2(_2495_),
    .Y(_2547_),
    .B1(_2545_));
 sg13g2_nor4_2 _6532_ (.A(_3249_),
    .B(_2464_),
    .C(_2544_),
    .Y(_2548_),
    .D(_2547_));
 sg13g2_nand3_1 _6533_ (.B(_2204_),
    .C(_2548_),
    .A(_2203_),
    .Y(_2549_));
 sg13g2_nor2_2 _6534_ (.A(_2201_),
    .B(_2549_),
    .Y(_2550_));
 sg13g2_nand2_1 _6535_ (.Y(_2551_),
    .A(net467),
    .B(_1937_));
 sg13g2_nand2b_1 _6536_ (.Y(_2552_),
    .B(_1896_),
    .A_N(net465));
 sg13g2_xor2_1 _6537_ (.B(_1896_),
    .A(net465),
    .X(_2553_));
 sg13g2_nand2b_1 _6538_ (.Y(_2554_),
    .B(_1929_),
    .A_N(net461));
 sg13g2_nand3_1 _6539_ (.B(_1923_),
    .C(_2554_),
    .A(_1274_),
    .Y(_2555_));
 sg13g2_nand2b_1 _6540_ (.Y(_2556_),
    .B(net461),
    .A_N(_1929_));
 sg13g2_nand2_1 _6541_ (.Y(_2558_),
    .A(_1234_),
    .B(_1936_));
 sg13g2_and3_1 _6542_ (.X(_2559_),
    .A(_2555_),
    .B(_2556_),
    .C(_2558_));
 sg13g2_o21ai_1 _6543_ (.B1(_2551_),
    .Y(_2560_),
    .A1(_2553_),
    .A2(_2559_));
 sg13g2_nor2_1 _6544_ (.A(_1307_),
    .B(_1903_),
    .Y(_2561_));
 sg13g2_xor2_1 _6545_ (.B(_1903_),
    .A(_1307_),
    .X(_2562_));
 sg13g2_o21ai_1 _6546_ (.B1(_2562_),
    .Y(_2563_),
    .A1(net463),
    .A2(_1917_));
 sg13g2_nand2_1 _6547_ (.Y(_2564_),
    .A(net464),
    .B(_1917_));
 sg13g2_xor2_1 _6548_ (.B(_1917_),
    .A(net463),
    .X(_2565_));
 sg13g2_mux2_1 _6549_ (.A0(_2565_),
    .A1(_2563_),
    .S(_2552_),
    .X(_2566_));
 sg13g2_o21ai_1 _6550_ (.B1(_2566_),
    .Y(_2567_),
    .A1(_2551_),
    .A2(_2553_));
 sg13g2_nand2_1 _6551_ (.Y(_2569_),
    .A(_1275_),
    .B(_2556_));
 sg13g2_o21ai_1 _6552_ (.B1(_2554_),
    .Y(_2570_),
    .A1(_1923_),
    .A2(_2569_));
 sg13g2_a21oi_1 _6553_ (.A1(_2551_),
    .A2(_2558_),
    .Y(_2571_),
    .B1(_2570_));
 sg13g2_nand2b_1 _6554_ (.Y(_2572_),
    .B(_1812_),
    .A_N(_1933_));
 sg13g2_nand2b_1 _6555_ (.Y(_2573_),
    .B(_1905_),
    .A_N(_1827_));
 sg13g2_a21oi_2 _6556_ (.B1(net508),
    .Y(_2574_),
    .A2(_2573_),
    .A1(_2572_));
 sg13g2_a21oi_1 _6557_ (.A1(_1308_),
    .A2(_2574_),
    .Y(_2575_),
    .B1(_2564_));
 sg13g2_nor2_1 _6558_ (.A(_2562_),
    .B(_2575_),
    .Y(_2576_));
 sg13g2_nand4_1 _6559_ (.B(net597),
    .C(\hvsync_gen.hpos[3] ),
    .A(net591),
    .Y(_2577_),
    .D(_2611_));
 sg13g2_nor2_1 _6560_ (.A(_3252_),
    .B(_2545_),
    .Y(_2578_));
 sg13g2_a21oi_2 _6561_ (.B1(_3249_),
    .Y(_2580_),
    .A2(_2578_),
    .A1(_2577_));
 sg13g2_o21ai_1 _6562_ (.B1(_2580_),
    .Y(_2581_),
    .A1(_2561_),
    .A2(_2574_));
 sg13g2_nor4_1 _6563_ (.A(_2567_),
    .B(_2571_),
    .C(_2576_),
    .D(_2581_),
    .Y(_2582_));
 sg13g2_a221oi_1 _6564_ (.B2(_2582_),
    .C1(net547),
    .B1(_2560_),
    .A1(_2202_),
    .Y(_2583_),
    .A2(_2550_));
 sg13g2_and4_1 _6565_ (.A(_2470_),
    .B(_2537_),
    .C(_2543_),
    .D(_2583_),
    .X(_2584_));
 sg13g2_a22oi_1 _6566_ (.Y(_0041_),
    .B1(_2504_),
    .B2(_2584_),
    .A2(_3257_),
    .A1(net549));
 sg13g2_dfrbp_1 _6567_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net35),
    .D(_0020_),
    .Q_N(_0010_),
    .Q(\hvsync_gen.hpos[0] ));
 sg13g2_dfrbp_1 _6568_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net32),
    .D(_0021_),
    .Q_N(_0000_),
    .Q(\hvsync_gen.hpos[1] ));
 sg13g2_dfrbp_1 _6569_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net30),
    .D(_0022_),
    .Q_N(_0017_),
    .Q(\hvsync_gen.hpos[2] ));
 sg13g2_dfrbp_1 _6570_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net28),
    .D(_0023_),
    .Q_N(_0016_),
    .Q(\hvsync_gen.hpos[3] ));
 sg13g2_dfrbp_1 _6571_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net26),
    .D(_0024_),
    .Q_N(_0015_),
    .Q(\hvsync_gen.hpos[4] ));
 sg13g2_dfrbp_1 _6572_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net24),
    .D(_0025_),
    .Q_N(_0018_),
    .Q(\hvsync_gen.hpos[5] ));
 sg13g2_dfrbp_1 _6573_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net22),
    .D(_0026_),
    .Q_N(_0014_),
    .Q(\hvsync_gen.hpos[6] ));
 sg13g2_dfrbp_1 _6574_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net20),
    .D(_0027_),
    .Q_N(_0001_),
    .Q(\hvsync_gen.hpos[7] ));
 sg13g2_dfrbp_1 _6575_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net18),
    .D(_0028_),
    .Q_N(_0013_),
    .Q(\hvsync_gen.hpos[8] ));
 sg13g2_dfrbp_1 _6576_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net38),
    .D(net52),
    .Q_N(_0019_),
    .Q(\hvsync_gen.hpos[9] ));
 sg13g2_dfrbp_1 _6577_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net36),
    .D(_0030_),
    .Q_N(_0006_),
    .Q(\hvsync_gen.vpos[0] ));
 sg13g2_dfrbp_1 _6578_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net34),
    .D(_0031_),
    .Q_N(_0012_),
    .Q(\hvsync_gen.vpos[1] ));
 sg13g2_dfrbp_1 _6579_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net31),
    .D(_0032_),
    .Q_N(_0011_),
    .Q(\hvsync_gen.vpos[2] ));
 sg13g2_dfrbp_1 _6580_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net27),
    .D(_0033_),
    .Q_N(_0009_),
    .Q(\hvsync_gen.vpos[3] ));
 sg13g2_dfrbp_1 _6581_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net23),
    .D(_0034_),
    .Q_N(_0003_),
    .Q(\hvsync_gen.vpos[4] ));
 sg13g2_dfrbp_1 _6582_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net19),
    .D(net57),
    .Q_N(_0008_),
    .Q(\hvsync_gen.vpos[5] ));
 sg13g2_dfrbp_1 _6583_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net37),
    .D(_0036_),
    .Q_N(_0007_),
    .Q(\hvsync_gen.vpos[6] ));
 sg13g2_dfrbp_1 _6584_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net33),
    .D(_0037_),
    .Q_N(_0005_),
    .Q(\hvsync_gen.vpos[7] ));
 sg13g2_dfrbp_1 _6585_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net25),
    .D(_0038_),
    .Q_N(_0004_),
    .Q(\hvsync_gen.vpos[8] ));
 sg13g2_dfrbp_1 _6586_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net39),
    .D(_0039_),
    .Q_N(_0002_),
    .Q(\hvsync_gen.vpos[9] ));
 sg13g2_dfrbp_1 _6587_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net29),
    .D(_0040_),
    .Q_N(_3279_),
    .Q(\hvsync_gen.phase ));
 sg13g2_dfrbp_1 _6588_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net21),
    .D(_0041_),
    .Q_N(_3280_),
    .Q(i_phase_0));
 sg13g2_tiehi _6582__19 (.L_HI(net19));
 sg13g2_tiehi _6574__20 (.L_HI(net20));
 sg13g2_tiehi _6588__21 (.L_HI(net21));
 sg13g2_tiehi _6573__22 (.L_HI(net22));
 sg13g2_tiehi _6581__23 (.L_HI(net23));
 sg13g2_tiehi _6572__24 (.L_HI(net24));
 sg13g2_tiehi _6585__25 (.L_HI(net25));
 sg13g2_tiehi _6571__26 (.L_HI(net26));
 sg13g2_tiehi _6580__27 (.L_HI(net27));
 sg13g2_tiehi _6570__28 (.L_HI(net28));
 sg13g2_tiehi _6587__29 (.L_HI(net29));
 sg13g2_tiehi _6569__30 (.L_HI(net30));
 sg13g2_tiehi _6579__31 (.L_HI(net31));
 sg13g2_tiehi _6568__32 (.L_HI(net32));
 sg13g2_tiehi _6584__33 (.L_HI(net33));
 sg13g2_tiehi _6578__34 (.L_HI(net34));
 sg13g2_tiehi _6567__35 (.L_HI(net35));
 sg13g2_tiehi _6577__36 (.L_HI(net36));
 sg13g2_tiehi _6583__37 (.L_HI(net37));
 sg13g2_tiehi _6576__38 (.L_HI(net38));
 sg13g2_tiehi _6586__39 (.L_HI(net39));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_dendraws_donut_3 (.L_LO(net3));
 sg13g2_tielo tt_um_dendraws_donut_4 (.L_LO(net4));
 sg13g2_tielo tt_um_dendraws_donut_5 (.L_LO(net5));
 sg13g2_tielo tt_um_dendraws_donut_6 (.L_LO(net6));
 sg13g2_tielo tt_um_dendraws_donut_7 (.L_LO(net7));
 sg13g2_tielo tt_um_dendraws_donut_8 (.L_LO(net8));
 sg13g2_tielo tt_um_dendraws_donut_9 (.L_LO(net9));
 sg13g2_tielo tt_um_dendraws_donut_10 (.L_LO(net10));
 sg13g2_tielo tt_um_dendraws_donut_11 (.L_LO(net11));
 sg13g2_tielo tt_um_dendraws_donut_12 (.L_LO(net12));
 sg13g2_tielo tt_um_dendraws_donut_13 (.L_LO(net13));
 sg13g2_tielo tt_um_dendraws_donut_14 (.L_LO(net14));
 sg13g2_tielo tt_um_dendraws_donut_15 (.L_LO(net15));
 sg13g2_tielo tt_um_dendraws_donut_16 (.L_LO(net16));
 sg13g2_tielo tt_um_dendraws_donut_17 (.L_LO(net17));
 sg13g2_tiehi _6575__18 (.L_HI(net18));
 sg13g2_buf_2 _6627_ (.A(uo_out[5]),
    .X(uo_out[0]));
 sg13g2_buf_2 _6628_ (.A(uo_out[2]),
    .X(uo_out[1]));
 sg13g2_buf_2 _6629_ (.A(\hvsync_gen.vsync ),
    .X(uo_out[3]));
 sg13g2_buf_2 _6630_ (.A(uo_out[5]),
    .X(uo_out[4]));
 sg13g2_buf_4 _6631_ (.X(uo_out[7]),
    .A(hsync));
 sg13g2_buf_4 fanout461 (.X(net461),
    .A(_1266_));
 sg13g2_buf_2 fanout462 (.A(_1266_),
    .X(net462));
 sg13g2_buf_2 fanout463 (.A(net464),
    .X(net463));
 sg13g2_buf_4 fanout464 (.X(net464),
    .A(_1255_));
 sg13g2_buf_4 fanout465 (.X(net465),
    .A(_1245_));
 sg13g2_buf_2 fanout466 (.A(_1245_),
    .X(net466));
 sg13g2_buf_4 fanout467 (.X(net467),
    .A(_1233_));
 sg13g2_buf_4 fanout468 (.X(net468),
    .A(_2841_));
 sg13g2_buf_4 fanout469 (.X(net469),
    .A(_0272_));
 sg13g2_buf_4 fanout470 (.X(net470),
    .A(_2817_));
 sg13g2_buf_2 fanout471 (.A(_2817_),
    .X(net471));
 sg13g2_buf_4 fanout472 (.X(net472),
    .A(_2882_));
 sg13g2_buf_2 fanout473 (.A(_2882_),
    .X(net473));
 sg13g2_buf_2 fanout474 (.A(_2884_),
    .X(net474));
 sg13g2_buf_4 fanout475 (.X(net475),
    .A(_2872_));
 sg13g2_buf_2 fanout476 (.A(_1222_),
    .X(net476));
 sg13g2_buf_2 fanout477 (.A(_0805_),
    .X(net477));
 sg13g2_buf_2 fanout478 (.A(_0483_),
    .X(net478));
 sg13g2_buf_2 fanout479 (.A(net480),
    .X(net479));
 sg13g2_buf_2 fanout480 (.A(_1473_),
    .X(net480));
 sg13g2_buf_2 fanout481 (.A(_0785_),
    .X(net481));
 sg13g2_buf_2 fanout482 (.A(_0473_),
    .X(net482));
 sg13g2_buf_2 fanout483 (.A(_0453_),
    .X(net483));
 sg13g2_buf_2 fanout484 (.A(_0165_),
    .X(net484));
 sg13g2_buf_1 fanout485 (.A(_0165_),
    .X(net485));
 sg13g2_buf_2 fanout486 (.A(_1712_),
    .X(net486));
 sg13g2_buf_2 fanout487 (.A(_1088_),
    .X(net487));
 sg13g2_buf_2 fanout488 (.A(_1088_),
    .X(net488));
 sg13g2_buf_2 fanout489 (.A(_0438_),
    .X(net489));
 sg13g2_buf_2 fanout490 (.A(_3024_),
    .X(net490));
 sg13g2_buf_2 fanout491 (.A(_1087_),
    .X(net491));
 sg13g2_buf_4 fanout492 (.X(net492),
    .A(_0441_));
 sg13g2_buf_2 fanout493 (.A(_0117_),
    .X(net493));
 sg13g2_buf_2 fanout494 (.A(net495),
    .X(net494));
 sg13g2_buf_2 fanout495 (.A(net496),
    .X(net495));
 sg13g2_buf_1 fanout496 (.A(_0765_),
    .X(net496));
 sg13g2_buf_2 fanout497 (.A(_0757_),
    .X(net497));
 sg13g2_buf_1 fanout498 (.A(_0757_),
    .X(net498));
 sg13g2_buf_4 fanout499 (.X(net499),
    .A(_3042_));
 sg13g2_buf_2 fanout500 (.A(_1403_),
    .X(net500));
 sg13g2_buf_2 fanout501 (.A(_0401_),
    .X(net501));
 sg13g2_buf_2 fanout502 (.A(_0095_),
    .X(net502));
 sg13g2_buf_2 fanout503 (.A(_3030_),
    .X(net503));
 sg13g2_buf_4 fanout504 (.X(net504),
    .A(_2700_));
 sg13g2_buf_2 fanout505 (.A(_2029_),
    .X(net505));
 sg13g2_buf_2 fanout506 (.A(net507),
    .X(net506));
 sg13g2_buf_2 fanout507 (.A(_1779_),
    .X(net507));
 sg13g2_buf_4 fanout508 (.X(net508),
    .A(_1772_));
 sg13g2_buf_2 fanout509 (.A(_1772_),
    .X(net509));
 sg13g2_buf_2 fanout510 (.A(_0096_),
    .X(net510));
 sg13g2_buf_2 fanout511 (.A(net512),
    .X(net511));
 sg13g2_buf_1 fanout512 (.A(_0093_),
    .X(net512));
 sg13g2_buf_2 fanout513 (.A(_1283_),
    .X(net513));
 sg13g2_buf_2 fanout514 (.A(_1195_),
    .X(net514));
 sg13g2_buf_2 fanout515 (.A(_2008_),
    .X(net515));
 sg13g2_buf_2 fanout516 (.A(net517),
    .X(net516));
 sg13g2_buf_2 fanout517 (.A(_1764_),
    .X(net517));
 sg13g2_buf_2 fanout518 (.A(_2995_),
    .X(net518));
 sg13g2_buf_2 fanout519 (.A(_1206_),
    .X(net519));
 sg13g2_buf_2 fanout520 (.A(_1085_),
    .X(net520));
 sg13g2_buf_4 fanout521 (.X(net521),
    .A(_2998_));
 sg13g2_buf_2 fanout522 (.A(_2608_),
    .X(net522));
 sg13g2_buf_2 fanout523 (.A(_3275_),
    .X(net523));
 sg13g2_buf_2 fanout524 (.A(_2961_),
    .X(net524));
 sg13g2_buf_1 fanout525 (.A(_2961_),
    .X(net525));
 sg13g2_buf_2 fanout526 (.A(_2352_),
    .X(net526));
 sg13g2_buf_2 fanout527 (.A(_2604_),
    .X(net527));
 sg13g2_buf_2 fanout528 (.A(_2596_),
    .X(net528));
 sg13g2_buf_4 fanout529 (.X(net529),
    .A(_0324_));
 sg13g2_buf_2 fanout530 (.A(_2590_),
    .X(net530));
 sg13g2_buf_2 fanout531 (.A(_2590_),
    .X(net531));
 sg13g2_buf_4 fanout532 (.X(net532),
    .A(_2937_));
 sg13g2_buf_2 fanout533 (.A(_2557_),
    .X(net533));
 sg13g2_buf_4 fanout534 (.X(net534),
    .A(_2546_));
 sg13g2_buf_2 fanout535 (.A(_2524_),
    .X(net535));
 sg13g2_buf_4 fanout536 (.X(net536),
    .A(_0271_));
 sg13g2_buf_4 fanout537 (.X(net537),
    .A(_3081_));
 sg13g2_buf_4 fanout538 (.X(net538),
    .A(net545));
 sg13g2_buf_2 fanout539 (.A(net545),
    .X(net539));
 sg13g2_buf_2 fanout540 (.A(net541),
    .X(net540));
 sg13g2_buf_2 fanout541 (.A(net545),
    .X(net541));
 sg13g2_buf_2 fanout542 (.A(net544),
    .X(net542));
 sg13g2_buf_1 fanout543 (.A(net544),
    .X(net543));
 sg13g2_buf_4 fanout544 (.X(net544),
    .A(net545));
 sg13g2_buf_2 fanout545 (.A(_3059_),
    .X(net545));
 sg13g2_buf_2 fanout546 (.A(net547),
    .X(net546));
 sg13g2_buf_2 fanout547 (.A(net548),
    .X(net547));
 sg13g2_buf_2 fanout548 (.A(net560),
    .X(net548));
 sg13g2_buf_2 fanout549 (.A(net550),
    .X(net549));
 sg13g2_buf_2 fanout550 (.A(net560),
    .X(net550));
 sg13g2_buf_2 fanout551 (.A(net552),
    .X(net551));
 sg13g2_buf_2 fanout552 (.A(net553),
    .X(net552));
 sg13g2_buf_1 fanout553 (.A(net560),
    .X(net553));
 sg13g2_buf_4 fanout554 (.X(net554),
    .A(net559));
 sg13g2_buf_2 fanout555 (.A(net559),
    .X(net555));
 sg13g2_buf_2 fanout556 (.A(net558),
    .X(net556));
 sg13g2_buf_1 fanout557 (.A(net558),
    .X(net557));
 sg13g2_buf_2 fanout558 (.A(net559),
    .X(net558));
 sg13g2_buf_2 fanout559 (.A(net560),
    .X(net559));
 sg13g2_buf_2 fanout560 (.A(\hvsync_gen.phase ),
    .X(net560));
 sg13g2_buf_4 fanout561 (.X(net561),
    .A(_0002_));
 sg13g2_buf_4 fanout562 (.X(net562),
    .A(_0004_));
 sg13g2_buf_4 fanout563 (.X(net563),
    .A(net564));
 sg13g2_buf_2 fanout564 (.A(net47),
    .X(net564));
 sg13g2_buf_2 fanout565 (.A(\hvsync_gen.vpos[5] ),
    .X(net565));
 sg13g2_buf_1 fanout566 (.A(net567),
    .X(net566));
 sg13g2_buf_2 fanout567 (.A(\hvsync_gen.vpos[5] ),
    .X(net567));
 sg13g2_buf_2 fanout568 (.A(net570),
    .X(net568));
 sg13g2_buf_4 fanout569 (.X(net569),
    .A(net570));
 sg13g2_buf_2 fanout570 (.A(\hvsync_gen.vpos[4] ),
    .X(net570));
 sg13g2_buf_2 fanout571 (.A(net572),
    .X(net571));
 sg13g2_buf_2 fanout572 (.A(\hvsync_gen.vpos[3] ),
    .X(net572));
 sg13g2_buf_4 fanout573 (.X(net573),
    .A(net575));
 sg13g2_buf_4 fanout574 (.X(net574),
    .A(net575));
 sg13g2_buf_2 fanout575 (.A(\hvsync_gen.vpos[2] ),
    .X(net575));
 sg13g2_buf_2 fanout576 (.A(net578),
    .X(net576));
 sg13g2_buf_2 fanout577 (.A(net578),
    .X(net577));
 sg13g2_buf_4 fanout578 (.X(net578),
    .A(net43));
 sg13g2_buf_2 fanout579 (.A(net580),
    .X(net579));
 sg13g2_buf_1 fanout580 (.A(\hvsync_gen.vpos[0] ),
    .X(net580));
 sg13g2_buf_4 fanout581 (.X(net581),
    .A(\hvsync_gen.vpos[0] ));
 sg13g2_buf_4 fanout582 (.X(net582),
    .A(\hvsync_gen.hpos[9] ));
 sg13g2_buf_2 fanout583 (.A(\hvsync_gen.hpos[9] ),
    .X(net583));
 sg13g2_buf_2 fanout584 (.A(net586),
    .X(net584));
 sg13g2_buf_4 fanout585 (.X(net585),
    .A(net586));
 sg13g2_buf_2 fanout586 (.A(\hvsync_gen.hpos[8] ),
    .X(net586));
 sg13g2_buf_4 fanout587 (.X(net587),
    .A(net588));
 sg13g2_buf_4 fanout588 (.X(net588),
    .A(\hvsync_gen.hpos[7] ));
 sg13g2_buf_4 fanout589 (.X(net589),
    .A(_0014_));
 sg13g2_buf_4 fanout590 (.X(net590),
    .A(\hvsync_gen.hpos[6] ));
 sg13g2_buf_2 fanout591 (.A(net53),
    .X(net591));
 sg13g2_buf_4 fanout592 (.X(net592),
    .A(net59));
 sg13g2_buf_2 fanout593 (.A(net595),
    .X(net593));
 sg13g2_buf_2 fanout594 (.A(net595),
    .X(net594));
 sg13g2_buf_2 fanout595 (.A(\hvsync_gen.hpos[5] ),
    .X(net595));
 sg13g2_buf_2 fanout596 (.A(net597),
    .X(net596));
 sg13g2_buf_4 fanout597 (.X(net597),
    .A(net58));
 sg13g2_buf_2 fanout598 (.A(net599),
    .X(net598));
 sg13g2_buf_2 fanout599 (.A(\hvsync_gen.hpos[3] ),
    .X(net599));
 sg13g2_buf_2 fanout600 (.A(_0017_),
    .X(net600));
 sg13g2_buf_4 fanout601 (.X(net601),
    .A(net603));
 sg13g2_buf_2 fanout602 (.A(net603),
    .X(net602));
 sg13g2_buf_2 fanout603 (.A(net604),
    .X(net603));
 sg13g2_buf_4 fanout604 (.X(net604),
    .A(\hvsync_gen.hpos[2] ));
 sg13g2_buf_2 fanout605 (.A(net606),
    .X(net605));
 sg13g2_buf_4 fanout606 (.X(net606),
    .A(\hvsync_gen.hpos[1] ));
 sg13g2_buf_4 fanout607 (.X(net607),
    .A(\hvsync_gen.hpos[0] ));
 sg13g2_buf_2 fanout608 (.A(\hvsync_gen.hpos[0] ),
    .X(net608));
 sg13g2_buf_4 fanout609 (.X(net609),
    .A(net610));
 sg13g2_buf_4 fanout610 (.X(net610),
    .A(_3268_));
 sg13g2_buf_4 input1 (.X(net1),
    .A(rst_n));
 sg13g2_tielo tt_um_dendraws_donut_2 (.L_LO(net2));
 sg13g2_buf_2 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .X(clknet_2_0__leaf_clk));
 sg13g2_buf_2 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .X(clknet_2_1__leaf_clk));
 sg13g2_buf_2 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .X(clknet_2_2__leaf_clk));
 sg13g2_buf_2 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .X(clknet_2_3__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_2_1__leaf_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_2_3__leaf_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(_3279_),
    .X(net40));
 sg13g2_dlygate4sd3_1 hold2 (.A(i_phase_0),
    .X(net41));
 sg13g2_dlygate4sd3_1 hold3 (.A(_0017_),
    .X(net42));
 sg13g2_dlygate4sd3_1 hold4 (.A(\hvsync_gen.vpos[1] ),
    .X(net43));
 sg13g2_dlygate4sd3_1 hold5 (.A(\hvsync_gen.vpos[9] ),
    .X(net44));
 sg13g2_dlygate4sd3_1 hold6 (.A(_0001_),
    .X(net45));
 sg13g2_dlygate4sd3_1 hold7 (.A(\hvsync_gen.vpos[7] ),
    .X(net46));
 sg13g2_dlygate4sd3_1 hold8 (.A(\hvsync_gen.vpos[8] ),
    .X(net47));
 sg13g2_dlygate4sd3_1 hold9 (.A(_0006_),
    .X(net48));
 sg13g2_dlygate4sd3_1 hold10 (.A(_0016_),
    .X(net49));
 sg13g2_dlygate4sd3_1 hold11 (.A(_2360_),
    .X(net50));
 sg13g2_dlygate4sd3_1 hold12 (.A(_0019_),
    .X(net51));
 sg13g2_dlygate4sd3_1 hold13 (.A(_0029_),
    .X(net52));
 sg13g2_dlygate4sd3_1 hold14 (.A(\hvsync_gen.hpos[6] ),
    .X(net53));
 sg13g2_dlygate4sd3_1 hold15 (.A(_0011_),
    .X(net54));
 sg13g2_dlygate4sd3_1 hold16 (.A(_2391_),
    .X(net55));
 sg13g2_dlygate4sd3_1 hold17 (.A(_0003_),
    .X(net56));
 sg13g2_dlygate4sd3_1 hold18 (.A(_0035_),
    .X(net57));
 sg13g2_dlygate4sd3_1 hold19 (.A(\hvsync_gen.hpos[4] ),
    .X(net58));
 sg13g2_dlygate4sd3_1 hold20 (.A(_0018_),
    .X(net59));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_4 FILLER_0_117 ();
 sg13g2_fill_1 FILLER_0_121 ();
 sg13g2_decap_4 FILLER_0_126 ();
 sg13g2_fill_1 FILLER_0_130 ();
 sg13g2_fill_2 FILLER_0_136 ();
 sg13g2_fill_1 FILLER_0_138 ();
 sg13g2_fill_1 FILLER_0_153 ();
 sg13g2_decap_4 FILLER_0_159 ();
 sg13g2_fill_2 FILLER_0_163 ();
 sg13g2_fill_2 FILLER_0_170 ();
 sg13g2_fill_1 FILLER_0_172 ();
 sg13g2_decap_8 FILLER_0_176 ();
 sg13g2_decap_8 FILLER_0_183 ();
 sg13g2_decap_4 FILLER_0_190 ();
 sg13g2_fill_1 FILLER_0_194 ();
 sg13g2_decap_8 FILLER_0_199 ();
 sg13g2_decap_8 FILLER_0_206 ();
 sg13g2_decap_8 FILLER_0_213 ();
 sg13g2_decap_8 FILLER_0_220 ();
 sg13g2_decap_8 FILLER_0_227 ();
 sg13g2_decap_8 FILLER_0_234 ();
 sg13g2_decap_8 FILLER_0_241 ();
 sg13g2_decap_8 FILLER_0_248 ();
 sg13g2_decap_8 FILLER_0_255 ();
 sg13g2_decap_8 FILLER_0_262 ();
 sg13g2_decap_8 FILLER_0_269 ();
 sg13g2_decap_8 FILLER_0_276 ();
 sg13g2_decap_8 FILLER_0_283 ();
 sg13g2_decap_8 FILLER_0_290 ();
 sg13g2_decap_8 FILLER_0_297 ();
 sg13g2_decap_8 FILLER_0_304 ();
 sg13g2_decap_8 FILLER_0_311 ();
 sg13g2_decap_8 FILLER_0_318 ();
 sg13g2_decap_8 FILLER_0_325 ();
 sg13g2_decap_8 FILLER_0_332 ();
 sg13g2_decap_8 FILLER_0_339 ();
 sg13g2_decap_8 FILLER_0_346 ();
 sg13g2_decap_8 FILLER_0_353 ();
 sg13g2_decap_8 FILLER_0_360 ();
 sg13g2_decap_8 FILLER_0_367 ();
 sg13g2_decap_8 FILLER_0_374 ();
 sg13g2_decap_8 FILLER_0_381 ();
 sg13g2_decap_8 FILLER_0_388 ();
 sg13g2_decap_8 FILLER_0_395 ();
 sg13g2_decap_8 FILLER_0_402 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_fill_2 FILLER_1_98 ();
 sg13g2_fill_1 FILLER_1_100 ();
 sg13g2_fill_1 FILLER_1_125 ();
 sg13g2_fill_2 FILLER_1_142 ();
 sg13g2_fill_2 FILLER_1_184 ();
 sg13g2_decap_8 FILLER_1_207 ();
 sg13g2_decap_8 FILLER_1_214 ();
 sg13g2_decap_8 FILLER_1_221 ();
 sg13g2_decap_8 FILLER_1_228 ();
 sg13g2_decap_8 FILLER_1_235 ();
 sg13g2_decap_8 FILLER_1_242 ();
 sg13g2_decap_8 FILLER_1_249 ();
 sg13g2_decap_8 FILLER_1_256 ();
 sg13g2_decap_8 FILLER_1_263 ();
 sg13g2_decap_8 FILLER_1_270 ();
 sg13g2_decap_8 FILLER_1_277 ();
 sg13g2_fill_1 FILLER_1_284 ();
 sg13g2_decap_8 FILLER_1_290 ();
 sg13g2_decap_8 FILLER_1_297 ();
 sg13g2_decap_8 FILLER_1_304 ();
 sg13g2_decap_8 FILLER_1_311 ();
 sg13g2_decap_8 FILLER_1_318 ();
 sg13g2_decap_8 FILLER_1_325 ();
 sg13g2_decap_8 FILLER_1_332 ();
 sg13g2_decap_8 FILLER_1_339 ();
 sg13g2_decap_8 FILLER_1_346 ();
 sg13g2_decap_8 FILLER_1_353 ();
 sg13g2_decap_8 FILLER_1_360 ();
 sg13g2_decap_8 FILLER_1_367 ();
 sg13g2_decap_8 FILLER_1_374 ();
 sg13g2_decap_8 FILLER_1_381 ();
 sg13g2_decap_8 FILLER_1_388 ();
 sg13g2_decap_8 FILLER_1_395 ();
 sg13g2_decap_8 FILLER_1_402 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_4 FILLER_2_49 ();
 sg13g2_fill_1 FILLER_2_53 ();
 sg13g2_fill_2 FILLER_2_59 ();
 sg13g2_decap_8 FILLER_2_69 ();
 sg13g2_decap_8 FILLER_2_76 ();
 sg13g2_decap_8 FILLER_2_83 ();
 sg13g2_decap_8 FILLER_2_90 ();
 sg13g2_decap_8 FILLER_2_97 ();
 sg13g2_decap_4 FILLER_2_104 ();
 sg13g2_fill_2 FILLER_2_108 ();
 sg13g2_decap_4 FILLER_2_115 ();
 sg13g2_fill_1 FILLER_2_119 ();
 sg13g2_fill_2 FILLER_2_125 ();
 sg13g2_fill_1 FILLER_2_127 ();
 sg13g2_fill_2 FILLER_2_132 ();
 sg13g2_fill_1 FILLER_2_138 ();
 sg13g2_decap_4 FILLER_2_143 ();
 sg13g2_fill_1 FILLER_2_156 ();
 sg13g2_decap_4 FILLER_2_162 ();
 sg13g2_fill_2 FILLER_2_166 ();
 sg13g2_decap_8 FILLER_2_173 ();
 sg13g2_decap_4 FILLER_2_180 ();
 sg13g2_fill_2 FILLER_2_184 ();
 sg13g2_decap_4 FILLER_2_190 ();
 sg13g2_decap_4 FILLER_2_198 ();
 sg13g2_fill_1 FILLER_2_202 ();
 sg13g2_fill_2 FILLER_2_225 ();
 sg13g2_fill_1 FILLER_2_227 ();
 sg13g2_decap_8 FILLER_2_233 ();
 sg13g2_decap_4 FILLER_2_240 ();
 sg13g2_decap_8 FILLER_2_248 ();
 sg13g2_decap_8 FILLER_2_255 ();
 sg13g2_decap_8 FILLER_2_262 ();
 sg13g2_fill_2 FILLER_2_274 ();
 sg13g2_fill_1 FILLER_2_276 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_81 ();
 sg13g2_decap_8 FILLER_3_88 ();
 sg13g2_decap_8 FILLER_3_95 ();
 sg13g2_fill_2 FILLER_3_102 ();
 sg13g2_fill_2 FILLER_3_108 ();
 sg13g2_fill_1 FILLER_3_110 ();
 sg13g2_decap_4 FILLER_3_116 ();
 sg13g2_fill_1 FILLER_3_148 ();
 sg13g2_fill_2 FILLER_3_154 ();
 sg13g2_fill_1 FILLER_3_176 ();
 sg13g2_fill_2 FILLER_3_193 ();
 sg13g2_fill_2 FILLER_3_215 ();
 sg13g2_fill_1 FILLER_3_230 ();
 sg13g2_fill_2 FILLER_3_249 ();
 sg13g2_fill_1 FILLER_3_251 ();
 sg13g2_fill_2 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_286 ();
 sg13g2_fill_2 FILLER_3_293 ();
 sg13g2_decap_8 FILLER_3_316 ();
 sg13g2_decap_8 FILLER_3_323 ();
 sg13g2_decap_8 FILLER_3_330 ();
 sg13g2_decap_8 FILLER_3_337 ();
 sg13g2_decap_8 FILLER_3_344 ();
 sg13g2_decap_8 FILLER_3_351 ();
 sg13g2_decap_8 FILLER_3_358 ();
 sg13g2_decap_8 FILLER_3_365 ();
 sg13g2_decap_8 FILLER_3_372 ();
 sg13g2_decap_8 FILLER_3_379 ();
 sg13g2_decap_8 FILLER_3_386 ();
 sg13g2_decap_8 FILLER_3_393 ();
 sg13g2_decap_8 FILLER_3_400 ();
 sg13g2_fill_2 FILLER_3_407 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_fill_2 FILLER_4_42 ();
 sg13g2_fill_1 FILLER_4_44 ();
 sg13g2_decap_4 FILLER_4_51 ();
 sg13g2_decap_4 FILLER_4_58 ();
 sg13g2_fill_1 FILLER_4_62 ();
 sg13g2_decap_8 FILLER_4_83 ();
 sg13g2_decap_8 FILLER_4_90 ();
 sg13g2_fill_2 FILLER_4_97 ();
 sg13g2_fill_1 FILLER_4_99 ();
 sg13g2_fill_1 FILLER_4_118 ();
 sg13g2_fill_1 FILLER_4_131 ();
 sg13g2_decap_4 FILLER_4_136 ();
 sg13g2_fill_1 FILLER_4_140 ();
 sg13g2_fill_1 FILLER_4_154 ();
 sg13g2_fill_2 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_178 ();
 sg13g2_decap_8 FILLER_4_185 ();
 sg13g2_decap_8 FILLER_4_192 ();
 sg13g2_fill_1 FILLER_4_199 ();
 sg13g2_fill_1 FILLER_4_205 ();
 sg13g2_fill_2 FILLER_4_216 ();
 sg13g2_fill_1 FILLER_4_218 ();
 sg13g2_decap_8 FILLER_4_228 ();
 sg13g2_decap_4 FILLER_4_235 ();
 sg13g2_fill_2 FILLER_4_239 ();
 sg13g2_fill_2 FILLER_4_265 ();
 sg13g2_fill_1 FILLER_4_275 ();
 sg13g2_fill_2 FILLER_4_302 ();
 sg13g2_decap_8 FILLER_4_317 ();
 sg13g2_decap_8 FILLER_4_324 ();
 sg13g2_decap_8 FILLER_4_331 ();
 sg13g2_decap_8 FILLER_4_338 ();
 sg13g2_decap_8 FILLER_4_345 ();
 sg13g2_decap_8 FILLER_4_352 ();
 sg13g2_decap_8 FILLER_4_359 ();
 sg13g2_decap_8 FILLER_4_366 ();
 sg13g2_decap_8 FILLER_4_373 ();
 sg13g2_decap_8 FILLER_4_380 ();
 sg13g2_decap_8 FILLER_4_387 ();
 sg13g2_decap_8 FILLER_4_394 ();
 sg13g2_decap_8 FILLER_4_401 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_fill_1 FILLER_5_42 ();
 sg13g2_fill_2 FILLER_5_51 ();
 sg13g2_fill_1 FILLER_5_53 ();
 sg13g2_decap_8 FILLER_5_78 ();
 sg13g2_decap_8 FILLER_5_85 ();
 sg13g2_decap_8 FILLER_5_92 ();
 sg13g2_decap_8 FILLER_5_99 ();
 sg13g2_fill_2 FILLER_5_106 ();
 sg13g2_decap_8 FILLER_5_120 ();
 sg13g2_fill_1 FILLER_5_137 ();
 sg13g2_decap_4 FILLER_5_142 ();
 sg13g2_fill_2 FILLER_5_153 ();
 sg13g2_fill_1 FILLER_5_155 ();
 sg13g2_fill_2 FILLER_5_161 ();
 sg13g2_fill_2 FILLER_5_173 ();
 sg13g2_fill_2 FILLER_5_201 ();
 sg13g2_fill_1 FILLER_5_223 ();
 sg13g2_decap_8 FILLER_5_232 ();
 sg13g2_fill_1 FILLER_5_239 ();
 sg13g2_fill_2 FILLER_5_254 ();
 sg13g2_fill_2 FILLER_5_260 ();
 sg13g2_fill_1 FILLER_5_262 ();
 sg13g2_fill_1 FILLER_5_288 ();
 sg13g2_decap_8 FILLER_5_307 ();
 sg13g2_decap_8 FILLER_5_314 ();
 sg13g2_decap_8 FILLER_5_321 ();
 sg13g2_decap_8 FILLER_5_328 ();
 sg13g2_decap_8 FILLER_5_335 ();
 sg13g2_decap_8 FILLER_5_342 ();
 sg13g2_decap_8 FILLER_5_349 ();
 sg13g2_decap_8 FILLER_5_356 ();
 sg13g2_decap_8 FILLER_5_363 ();
 sg13g2_decap_8 FILLER_5_370 ();
 sg13g2_decap_8 FILLER_5_377 ();
 sg13g2_decap_8 FILLER_5_384 ();
 sg13g2_decap_8 FILLER_5_391 ();
 sg13g2_decap_8 FILLER_5_398 ();
 sg13g2_decap_4 FILLER_5_405 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_50 ();
 sg13g2_fill_2 FILLER_6_57 ();
 sg13g2_fill_1 FILLER_6_59 ();
 sg13g2_fill_1 FILLER_6_65 ();
 sg13g2_fill_1 FILLER_6_70 ();
 sg13g2_decap_4 FILLER_6_84 ();
 sg13g2_fill_1 FILLER_6_100 ();
 sg13g2_decap_4 FILLER_6_109 ();
 sg13g2_fill_1 FILLER_6_113 ();
 sg13g2_fill_2 FILLER_6_127 ();
 sg13g2_fill_1 FILLER_6_145 ();
 sg13g2_decap_4 FILLER_6_154 ();
 sg13g2_decap_4 FILLER_6_166 ();
 sg13g2_decap_4 FILLER_6_185 ();
 sg13g2_fill_1 FILLER_6_194 ();
 sg13g2_decap_4 FILLER_6_200 ();
 sg13g2_fill_2 FILLER_6_204 ();
 sg13g2_decap_8 FILLER_6_211 ();
 sg13g2_decap_8 FILLER_6_218 ();
 sg13g2_fill_1 FILLER_6_225 ();
 sg13g2_fill_1 FILLER_6_264 ();
 sg13g2_fill_1 FILLER_6_270 ();
 sg13g2_fill_2 FILLER_6_275 ();
 sg13g2_fill_1 FILLER_6_277 ();
 sg13g2_decap_4 FILLER_6_291 ();
 sg13g2_fill_1 FILLER_6_295 ();
 sg13g2_decap_8 FILLER_6_304 ();
 sg13g2_decap_8 FILLER_6_311 ();
 sg13g2_decap_8 FILLER_6_318 ();
 sg13g2_decap_8 FILLER_6_325 ();
 sg13g2_decap_8 FILLER_6_332 ();
 sg13g2_decap_8 FILLER_6_339 ();
 sg13g2_decap_8 FILLER_6_346 ();
 sg13g2_decap_8 FILLER_6_353 ();
 sg13g2_decap_8 FILLER_6_360 ();
 sg13g2_decap_8 FILLER_6_367 ();
 sg13g2_decap_8 FILLER_6_374 ();
 sg13g2_decap_8 FILLER_6_381 ();
 sg13g2_decap_8 FILLER_6_388 ();
 sg13g2_decap_8 FILLER_6_395 ();
 sg13g2_decap_8 FILLER_6_402 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_fill_2 FILLER_7_65 ();
 sg13g2_fill_1 FILLER_7_79 ();
 sg13g2_decap_4 FILLER_7_88 ();
 sg13g2_fill_2 FILLER_7_92 ();
 sg13g2_fill_1 FILLER_7_102 ();
 sg13g2_decap_4 FILLER_7_121 ();
 sg13g2_fill_2 FILLER_7_125 ();
 sg13g2_fill_2 FILLER_7_132 ();
 sg13g2_fill_1 FILLER_7_134 ();
 sg13g2_fill_2 FILLER_7_141 ();
 sg13g2_fill_1 FILLER_7_143 ();
 sg13g2_decap_4 FILLER_7_149 ();
 sg13g2_decap_4 FILLER_7_161 ();
 sg13g2_decap_4 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_184 ();
 sg13g2_fill_2 FILLER_7_199 ();
 sg13g2_fill_1 FILLER_7_201 ();
 sg13g2_decap_4 FILLER_7_210 ();
 sg13g2_fill_1 FILLER_7_214 ();
 sg13g2_fill_1 FILLER_7_227 ();
 sg13g2_decap_8 FILLER_7_232 ();
 sg13g2_fill_2 FILLER_7_239 ();
 sg13g2_fill_1 FILLER_7_241 ();
 sg13g2_fill_2 FILLER_7_254 ();
 sg13g2_fill_1 FILLER_7_266 ();
 sg13g2_fill_1 FILLER_7_275 ();
 sg13g2_fill_1 FILLER_7_281 ();
 sg13g2_fill_1 FILLER_7_290 ();
 sg13g2_fill_1 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_310 ();
 sg13g2_decap_8 FILLER_7_317 ();
 sg13g2_decap_8 FILLER_7_324 ();
 sg13g2_decap_8 FILLER_7_331 ();
 sg13g2_decap_8 FILLER_7_338 ();
 sg13g2_decap_8 FILLER_7_345 ();
 sg13g2_decap_8 FILLER_7_352 ();
 sg13g2_decap_8 FILLER_7_359 ();
 sg13g2_decap_8 FILLER_7_366 ();
 sg13g2_decap_8 FILLER_7_373 ();
 sg13g2_decap_8 FILLER_7_380 ();
 sg13g2_decap_8 FILLER_7_387 ();
 sg13g2_decap_8 FILLER_7_394 ();
 sg13g2_decap_8 FILLER_7_401 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_4 FILLER_8_35 ();
 sg13g2_fill_1 FILLER_8_39 ();
 sg13g2_fill_1 FILLER_8_56 ();
 sg13g2_decap_4 FILLER_8_62 ();
 sg13g2_fill_2 FILLER_8_74 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_fill_2 FILLER_8_110 ();
 sg13g2_fill_1 FILLER_8_112 ();
 sg13g2_fill_2 FILLER_8_132 ();
 sg13g2_fill_2 FILLER_8_150 ();
 sg13g2_fill_1 FILLER_8_152 ();
 sg13g2_fill_2 FILLER_8_161 ();
 sg13g2_decap_4 FILLER_8_179 ();
 sg13g2_fill_1 FILLER_8_191 ();
 sg13g2_fill_2 FILLER_8_200 ();
 sg13g2_fill_1 FILLER_8_210 ();
 sg13g2_fill_1 FILLER_8_225 ();
 sg13g2_fill_2 FILLER_8_258 ();
 sg13g2_fill_1 FILLER_8_260 ();
 sg13g2_fill_2 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_274 ();
 sg13g2_decap_8 FILLER_8_286 ();
 sg13g2_decap_8 FILLER_8_293 ();
 sg13g2_fill_2 FILLER_8_300 ();
 sg13g2_fill_1 FILLER_8_302 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_4 FILLER_9_49 ();
 sg13g2_fill_2 FILLER_9_53 ();
 sg13g2_decap_4 FILLER_9_60 ();
 sg13g2_fill_2 FILLER_9_72 ();
 sg13g2_fill_1 FILLER_9_78 ();
 sg13g2_fill_2 FILLER_9_100 ();
 sg13g2_fill_1 FILLER_9_102 ();
 sg13g2_decap_8 FILLER_9_108 ();
 sg13g2_fill_2 FILLER_9_120 ();
 sg13g2_decap_4 FILLER_9_131 ();
 sg13g2_fill_2 FILLER_9_135 ();
 sg13g2_decap_8 FILLER_9_141 ();
 sg13g2_fill_2 FILLER_9_155 ();
 sg13g2_fill_1 FILLER_9_157 ();
 sg13g2_decap_4 FILLER_9_182 ();
 sg13g2_fill_1 FILLER_9_186 ();
 sg13g2_fill_2 FILLER_9_204 ();
 sg13g2_fill_1 FILLER_9_210 ();
 sg13g2_fill_2 FILLER_9_226 ();
 sg13g2_decap_8 FILLER_9_232 ();
 sg13g2_fill_2 FILLER_9_244 ();
 sg13g2_fill_2 FILLER_9_250 ();
 sg13g2_fill_1 FILLER_9_252 ();
 sg13g2_fill_1 FILLER_9_271 ();
 sg13g2_fill_1 FILLER_9_284 ();
 sg13g2_fill_1 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_4 FILLER_10_35 ();
 sg13g2_fill_2 FILLER_10_71 ();
 sg13g2_fill_2 FILLER_10_78 ();
 sg13g2_fill_1 FILLER_10_80 ();
 sg13g2_fill_2 FILLER_10_94 ();
 sg13g2_fill_1 FILLER_10_96 ();
 sg13g2_fill_1 FILLER_10_113 ();
 sg13g2_fill_2 FILLER_10_122 ();
 sg13g2_fill_2 FILLER_10_132 ();
 sg13g2_fill_1 FILLER_10_134 ();
 sg13g2_fill_2 FILLER_10_148 ();
 sg13g2_fill_2 FILLER_10_163 ();
 sg13g2_fill_1 FILLER_10_165 ();
 sg13g2_decap_4 FILLER_10_169 ();
 sg13g2_fill_1 FILLER_10_173 ();
 sg13g2_fill_2 FILLER_10_178 ();
 sg13g2_fill_2 FILLER_10_188 ();
 sg13g2_fill_2 FILLER_10_213 ();
 sg13g2_decap_4 FILLER_10_244 ();
 sg13g2_fill_2 FILLER_10_248 ();
 sg13g2_decap_8 FILLER_10_262 ();
 sg13g2_decap_8 FILLER_10_269 ();
 sg13g2_fill_1 FILLER_10_276 ();
 sg13g2_decap_8 FILLER_10_309 ();
 sg13g2_decap_8 FILLER_10_316 ();
 sg13g2_decap_8 FILLER_10_323 ();
 sg13g2_decap_8 FILLER_10_330 ();
 sg13g2_decap_8 FILLER_10_337 ();
 sg13g2_decap_8 FILLER_10_344 ();
 sg13g2_decap_8 FILLER_10_351 ();
 sg13g2_decap_8 FILLER_10_358 ();
 sg13g2_decap_8 FILLER_10_365 ();
 sg13g2_decap_8 FILLER_10_372 ();
 sg13g2_decap_8 FILLER_10_379 ();
 sg13g2_decap_8 FILLER_10_386 ();
 sg13g2_decap_8 FILLER_10_393 ();
 sg13g2_decap_8 FILLER_10_400 ();
 sg13g2_fill_2 FILLER_10_407 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_fill_2 FILLER_11_53 ();
 sg13g2_fill_1 FILLER_11_71 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_fill_1 FILLER_11_100 ();
 sg13g2_fill_2 FILLER_11_119 ();
 sg13g2_fill_2 FILLER_11_131 ();
 sg13g2_fill_1 FILLER_11_133 ();
 sg13g2_fill_1 FILLER_11_140 ();
 sg13g2_fill_1 FILLER_11_149 ();
 sg13g2_fill_2 FILLER_11_162 ();
 sg13g2_fill_2 FILLER_11_180 ();
 sg13g2_fill_1 FILLER_11_182 ();
 sg13g2_fill_1 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_201 ();
 sg13g2_decap_4 FILLER_11_208 ();
 sg13g2_fill_2 FILLER_11_212 ();
 sg13g2_decap_4 FILLER_11_222 ();
 sg13g2_fill_2 FILLER_11_226 ();
 sg13g2_fill_2 FILLER_11_236 ();
 sg13g2_fill_2 FILLER_11_252 ();
 sg13g2_fill_2 FILLER_11_261 ();
 sg13g2_fill_1 FILLER_11_263 ();
 sg13g2_fill_1 FILLER_11_268 ();
 sg13g2_decap_8 FILLER_11_281 ();
 sg13g2_fill_1 FILLER_11_288 ();
 sg13g2_fill_2 FILLER_11_298 ();
 sg13g2_fill_1 FILLER_11_300 ();
 sg13g2_decap_8 FILLER_11_309 ();
 sg13g2_decap_4 FILLER_11_316 ();
 sg13g2_fill_2 FILLER_11_320 ();
 sg13g2_fill_1 FILLER_11_327 ();
 sg13g2_decap_8 FILLER_11_333 ();
 sg13g2_decap_8 FILLER_11_340 ();
 sg13g2_decap_8 FILLER_11_347 ();
 sg13g2_decap_8 FILLER_11_354 ();
 sg13g2_decap_8 FILLER_11_361 ();
 sg13g2_decap_8 FILLER_11_368 ();
 sg13g2_decap_8 FILLER_11_375 ();
 sg13g2_decap_8 FILLER_11_382 ();
 sg13g2_decap_8 FILLER_11_389 ();
 sg13g2_decap_8 FILLER_11_396 ();
 sg13g2_decap_4 FILLER_11_403 ();
 sg13g2_fill_2 FILLER_11_407 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_4 FILLER_12_35 ();
 sg13g2_fill_1 FILLER_12_39 ();
 sg13g2_fill_1 FILLER_12_45 ();
 sg13g2_fill_1 FILLER_12_70 ();
 sg13g2_fill_1 FILLER_12_79 ();
 sg13g2_fill_2 FILLER_12_93 ();
 sg13g2_decap_4 FILLER_12_111 ();
 sg13g2_fill_1 FILLER_12_121 ();
 sg13g2_fill_2 FILLER_12_128 ();
 sg13g2_fill_2 FILLER_12_135 ();
 sg13g2_decap_8 FILLER_12_145 ();
 sg13g2_decap_4 FILLER_12_152 ();
 sg13g2_fill_1 FILLER_12_156 ();
 sg13g2_decap_8 FILLER_12_162 ();
 sg13g2_decap_4 FILLER_12_169 ();
 sg13g2_decap_8 FILLER_12_177 ();
 sg13g2_decap_4 FILLER_12_194 ();
 sg13g2_decap_8 FILLER_12_211 ();
 sg13g2_decap_8 FILLER_12_218 ();
 sg13g2_fill_2 FILLER_12_225 ();
 sg13g2_fill_1 FILLER_12_227 ();
 sg13g2_fill_1 FILLER_12_237 ();
 sg13g2_fill_1 FILLER_12_252 ();
 sg13g2_fill_2 FILLER_12_257 ();
 sg13g2_fill_1 FILLER_12_259 ();
 sg13g2_fill_2 FILLER_12_265 ();
 sg13g2_fill_1 FILLER_12_276 ();
 sg13g2_fill_1 FILLER_12_282 ();
 sg13g2_fill_2 FILLER_12_289 ();
 sg13g2_fill_1 FILLER_12_299 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_fill_2 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_fill_2 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_54 ();
 sg13g2_decap_4 FILLER_13_61 ();
 sg13g2_fill_2 FILLER_13_65 ();
 sg13g2_decap_8 FILLER_13_76 ();
 sg13g2_fill_1 FILLER_13_83 ();
 sg13g2_fill_2 FILLER_13_88 ();
 sg13g2_fill_1 FILLER_13_90 ();
 sg13g2_fill_2 FILLER_13_103 ();
 sg13g2_fill_1 FILLER_13_135 ();
 sg13g2_fill_2 FILLER_13_140 ();
 sg13g2_fill_1 FILLER_13_155 ();
 sg13g2_fill_1 FILLER_13_164 ();
 sg13g2_fill_2 FILLER_13_170 ();
 sg13g2_fill_1 FILLER_13_188 ();
 sg13g2_fill_2 FILLER_13_197 ();
 sg13g2_fill_2 FILLER_13_206 ();
 sg13g2_fill_2 FILLER_13_221 ();
 sg13g2_fill_2 FILLER_13_254 ();
 sg13g2_decap_4 FILLER_13_274 ();
 sg13g2_fill_2 FILLER_13_278 ();
 sg13g2_fill_2 FILLER_13_293 ();
 sg13g2_decap_8 FILLER_13_303 ();
 sg13g2_fill_2 FILLER_13_318 ();
 sg13g2_decap_4 FILLER_13_324 ();
 sg13g2_fill_1 FILLER_13_328 ();
 sg13g2_decap_8 FILLER_13_342 ();
 sg13g2_decap_8 FILLER_13_349 ();
 sg13g2_decap_8 FILLER_13_356 ();
 sg13g2_decap_8 FILLER_13_363 ();
 sg13g2_decap_8 FILLER_13_370 ();
 sg13g2_decap_8 FILLER_13_377 ();
 sg13g2_decap_8 FILLER_13_384 ();
 sg13g2_decap_8 FILLER_13_391 ();
 sg13g2_decap_8 FILLER_13_398 ();
 sg13g2_decap_4 FILLER_13_405 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_4 FILLER_14_28 ();
 sg13g2_fill_2 FILLER_14_32 ();
 sg13g2_decap_8 FILLER_14_39 ();
 sg13g2_fill_1 FILLER_14_46 ();
 sg13g2_decap_4 FILLER_14_52 ();
 sg13g2_fill_1 FILLER_14_56 ();
 sg13g2_fill_1 FILLER_14_62 ();
 sg13g2_decap_4 FILLER_14_73 ();
 sg13g2_fill_1 FILLER_14_82 ();
 sg13g2_fill_2 FILLER_14_88 ();
 sg13g2_fill_2 FILLER_14_95 ();
 sg13g2_decap_8 FILLER_14_113 ();
 sg13g2_fill_2 FILLER_14_120 ();
 sg13g2_fill_1 FILLER_14_122 ();
 sg13g2_fill_2 FILLER_14_126 ();
 sg13g2_fill_1 FILLER_14_128 ();
 sg13g2_decap_8 FILLER_14_139 ();
 sg13g2_decap_4 FILLER_14_150 ();
 sg13g2_fill_1 FILLER_14_160 ();
 sg13g2_fill_1 FILLER_14_171 ();
 sg13g2_fill_2 FILLER_14_177 ();
 sg13g2_fill_2 FILLER_14_189 ();
 sg13g2_fill_1 FILLER_14_214 ();
 sg13g2_decap_8 FILLER_14_234 ();
 sg13g2_decap_4 FILLER_14_241 ();
 sg13g2_fill_1 FILLER_14_245 ();
 sg13g2_decap_4 FILLER_14_251 ();
 sg13g2_decap_4 FILLER_14_259 ();
 sg13g2_fill_1 FILLER_14_263 ();
 sg13g2_decap_4 FILLER_14_282 ();
 sg13g2_fill_1 FILLER_14_304 ();
 sg13g2_fill_1 FILLER_14_313 ();
 sg13g2_fill_2 FILLER_14_333 ();
 sg13g2_decap_8 FILLER_14_361 ();
 sg13g2_decap_8 FILLER_14_368 ();
 sg13g2_decap_8 FILLER_14_375 ();
 sg13g2_decap_8 FILLER_14_382 ();
 sg13g2_decap_8 FILLER_14_389 ();
 sg13g2_decap_8 FILLER_14_396 ();
 sg13g2_decap_4 FILLER_14_403 ();
 sg13g2_fill_2 FILLER_14_407 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_4 FILLER_15_21 ();
 sg13g2_fill_1 FILLER_15_25 ();
 sg13g2_fill_2 FILLER_15_39 ();
 sg13g2_fill_2 FILLER_15_53 ();
 sg13g2_decap_4 FILLER_15_62 ();
 sg13g2_fill_1 FILLER_15_73 ();
 sg13g2_fill_1 FILLER_15_86 ();
 sg13g2_decap_8 FILLER_15_95 ();
 sg13g2_fill_1 FILLER_15_102 ();
 sg13g2_decap_8 FILLER_15_107 ();
 sg13g2_fill_2 FILLER_15_114 ();
 sg13g2_fill_1 FILLER_15_128 ();
 sg13g2_fill_2 FILLER_15_142 ();
 sg13g2_fill_1 FILLER_15_144 ();
 sg13g2_decap_8 FILLER_15_157 ();
 sg13g2_decap_4 FILLER_15_164 ();
 sg13g2_fill_1 FILLER_15_181 ();
 sg13g2_decap_8 FILLER_15_204 ();
 sg13g2_decap_8 FILLER_15_211 ();
 sg13g2_fill_2 FILLER_15_218 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_4 FILLER_15_231 ();
 sg13g2_fill_2 FILLER_15_235 ();
 sg13g2_fill_2 FILLER_15_266 ();
 sg13g2_fill_1 FILLER_15_268 ();
 sg13g2_decap_4 FILLER_15_277 ();
 sg13g2_fill_2 FILLER_15_292 ();
 sg13g2_fill_1 FILLER_15_302 ();
 sg13g2_decap_8 FILLER_15_307 ();
 sg13g2_fill_2 FILLER_15_314 ();
 sg13g2_fill_1 FILLER_15_316 ();
 sg13g2_decap_8 FILLER_15_322 ();
 sg13g2_fill_1 FILLER_15_329 ();
 sg13g2_decap_8 FILLER_15_344 ();
 sg13g2_decap_8 FILLER_15_351 ();
 sg13g2_decap_8 FILLER_15_358 ();
 sg13g2_decap_8 FILLER_15_365 ();
 sg13g2_decap_8 FILLER_15_372 ();
 sg13g2_decap_8 FILLER_15_379 ();
 sg13g2_decap_8 FILLER_15_386 ();
 sg13g2_decap_8 FILLER_15_393 ();
 sg13g2_decap_8 FILLER_15_400 ();
 sg13g2_fill_2 FILLER_15_407 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_4 FILLER_16_35 ();
 sg13g2_fill_1 FILLER_16_39 ();
 sg13g2_fill_2 FILLER_16_52 ();
 sg13g2_fill_2 FILLER_16_59 ();
 sg13g2_fill_1 FILLER_16_61 ();
 sg13g2_fill_1 FILLER_16_68 ();
 sg13g2_decap_4 FILLER_16_75 ();
 sg13g2_fill_2 FILLER_16_89 ();
 sg13g2_fill_2 FILLER_16_102 ();
 sg13g2_fill_1 FILLER_16_104 ();
 sg13g2_fill_2 FILLER_16_128 ();
 sg13g2_fill_1 FILLER_16_130 ();
 sg13g2_decap_4 FILLER_16_167 ();
 sg13g2_fill_1 FILLER_16_171 ();
 sg13g2_decap_8 FILLER_16_178 ();
 sg13g2_decap_8 FILLER_16_185 ();
 sg13g2_decap_4 FILLER_16_197 ();
 sg13g2_fill_1 FILLER_16_201 ();
 sg13g2_fill_1 FILLER_16_214 ();
 sg13g2_fill_2 FILLER_16_265 ();
 sg13g2_fill_2 FILLER_16_284 ();
 sg13g2_fill_1 FILLER_16_286 ();
 sg13g2_fill_2 FILLER_16_301 ();
 sg13g2_decap_4 FILLER_16_323 ();
 sg13g2_fill_1 FILLER_16_327 ();
 sg13g2_fill_2 FILLER_16_343 ();
 sg13g2_fill_1 FILLER_16_345 ();
 sg13g2_decap_8 FILLER_16_354 ();
 sg13g2_decap_8 FILLER_16_361 ();
 sg13g2_decap_8 FILLER_16_368 ();
 sg13g2_decap_8 FILLER_16_375 ();
 sg13g2_decap_8 FILLER_16_382 ();
 sg13g2_decap_8 FILLER_16_389 ();
 sg13g2_decap_8 FILLER_16_396 ();
 sg13g2_decap_4 FILLER_16_403 ();
 sg13g2_fill_2 FILLER_16_407 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_fill_2 FILLER_17_28 ();
 sg13g2_fill_1 FILLER_17_30 ();
 sg13g2_fill_2 FILLER_17_44 ();
 sg13g2_fill_2 FILLER_17_65 ();
 sg13g2_decap_4 FILLER_17_75 ();
 sg13g2_decap_4 FILLER_17_88 ();
 sg13g2_decap_8 FILLER_17_107 ();
 sg13g2_fill_2 FILLER_17_120 ();
 sg13g2_fill_1 FILLER_17_122 ();
 sg13g2_fill_1 FILLER_17_128 ();
 sg13g2_fill_1 FILLER_17_134 ();
 sg13g2_fill_2 FILLER_17_140 ();
 sg13g2_fill_1 FILLER_17_142 ();
 sg13g2_fill_2 FILLER_17_151 ();
 sg13g2_fill_1 FILLER_17_153 ();
 sg13g2_decap_8 FILLER_17_167 ();
 sg13g2_decap_4 FILLER_17_178 ();
 sg13g2_fill_2 FILLER_17_203 ();
 sg13g2_decap_4 FILLER_17_210 ();
 sg13g2_decap_4 FILLER_17_222 ();
 sg13g2_fill_1 FILLER_17_226 ();
 sg13g2_fill_1 FILLER_17_231 ();
 sg13g2_fill_1 FILLER_17_237 ();
 sg13g2_decap_4 FILLER_17_242 ();
 sg13g2_decap_4 FILLER_17_251 ();
 sg13g2_fill_1 FILLER_17_255 ();
 sg13g2_fill_2 FILLER_17_261 ();
 sg13g2_fill_1 FILLER_17_267 ();
 sg13g2_fill_2 FILLER_17_276 ();
 sg13g2_fill_2 FILLER_17_287 ();
 sg13g2_fill_1 FILLER_17_297 ();
 sg13g2_fill_2 FILLER_17_302 ();
 sg13g2_fill_1 FILLER_17_304 ();
 sg13g2_fill_2 FILLER_17_310 ();
 sg13g2_fill_1 FILLER_17_312 ();
 sg13g2_fill_2 FILLER_17_334 ();
 sg13g2_decap_8 FILLER_17_355 ();
 sg13g2_decap_8 FILLER_17_362 ();
 sg13g2_decap_8 FILLER_17_369 ();
 sg13g2_decap_8 FILLER_17_376 ();
 sg13g2_decap_8 FILLER_17_383 ();
 sg13g2_decap_8 FILLER_17_390 ();
 sg13g2_decap_8 FILLER_17_397 ();
 sg13g2_decap_4 FILLER_17_404 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_fill_2 FILLER_18_28 ();
 sg13g2_decap_4 FILLER_18_38 ();
 sg13g2_decap_4 FILLER_18_57 ();
 sg13g2_fill_2 FILLER_18_61 ();
 sg13g2_fill_2 FILLER_18_72 ();
 sg13g2_fill_1 FILLER_18_74 ();
 sg13g2_fill_2 FILLER_18_85 ();
 sg13g2_decap_8 FILLER_18_92 ();
 sg13g2_fill_1 FILLER_18_99 ();
 sg13g2_fill_1 FILLER_18_115 ();
 sg13g2_fill_1 FILLER_18_125 ();
 sg13g2_fill_2 FILLER_18_134 ();
 sg13g2_fill_1 FILLER_18_136 ();
 sg13g2_decap_4 FILLER_18_145 ();
 sg13g2_fill_2 FILLER_18_157 ();
 sg13g2_fill_1 FILLER_18_159 ();
 sg13g2_fill_2 FILLER_18_172 ();
 sg13g2_fill_1 FILLER_18_188 ();
 sg13g2_fill_2 FILLER_18_201 ();
 sg13g2_decap_4 FILLER_18_211 ();
 sg13g2_fill_2 FILLER_18_223 ();
 sg13g2_fill_1 FILLER_18_258 ();
 sg13g2_fill_1 FILLER_18_279 ();
 sg13g2_decap_8 FILLER_18_285 ();
 sg13g2_fill_1 FILLER_18_292 ();
 sg13g2_fill_2 FILLER_18_303 ();
 sg13g2_fill_2 FILLER_18_310 ();
 sg13g2_fill_2 FILLER_18_324 ();
 sg13g2_fill_1 FILLER_18_326 ();
 sg13g2_fill_1 FILLER_18_330 ();
 sg13g2_fill_1 FILLER_18_335 ();
 sg13g2_decap_4 FILLER_18_340 ();
 sg13g2_fill_1 FILLER_18_344 ();
 sg13g2_decap_8 FILLER_18_363 ();
 sg13g2_decap_8 FILLER_18_370 ();
 sg13g2_decap_8 FILLER_18_377 ();
 sg13g2_decap_8 FILLER_18_384 ();
 sg13g2_decap_8 FILLER_18_391 ();
 sg13g2_decap_8 FILLER_18_398 ();
 sg13g2_decap_4 FILLER_18_405 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_4 FILLER_19_35 ();
 sg13g2_fill_2 FILLER_19_39 ();
 sg13g2_fill_1 FILLER_19_48 ();
 sg13g2_fill_2 FILLER_19_87 ();
 sg13g2_fill_1 FILLER_19_89 ();
 sg13g2_decap_4 FILLER_19_111 ();
 sg13g2_fill_1 FILLER_19_115 ();
 sg13g2_decap_4 FILLER_19_120 ();
 sg13g2_fill_1 FILLER_19_124 ();
 sg13g2_fill_2 FILLER_19_135 ();
 sg13g2_fill_2 FILLER_19_152 ();
 sg13g2_decap_4 FILLER_19_164 ();
 sg13g2_fill_1 FILLER_19_168 ();
 sg13g2_decap_4 FILLER_19_173 ();
 sg13g2_fill_2 FILLER_19_177 ();
 sg13g2_fill_2 FILLER_19_191 ();
 sg13g2_fill_2 FILLER_19_198 ();
 sg13g2_fill_1 FILLER_19_200 ();
 sg13g2_fill_2 FILLER_19_209 ();
 sg13g2_decap_8 FILLER_19_227 ();
 sg13g2_decap_8 FILLER_19_234 ();
 sg13g2_decap_4 FILLER_19_241 ();
 sg13g2_fill_1 FILLER_19_245 ();
 sg13g2_decap_8 FILLER_19_266 ();
 sg13g2_decap_8 FILLER_19_273 ();
 sg13g2_fill_1 FILLER_19_280 ();
 sg13g2_decap_4 FILLER_19_285 ();
 sg13g2_fill_2 FILLER_19_319 ();
 sg13g2_decap_8 FILLER_19_359 ();
 sg13g2_decap_8 FILLER_19_366 ();
 sg13g2_decap_8 FILLER_19_373 ();
 sg13g2_decap_8 FILLER_19_380 ();
 sg13g2_decap_8 FILLER_19_387 ();
 sg13g2_decap_8 FILLER_19_394 ();
 sg13g2_decap_8 FILLER_19_401 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_fill_1 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_55 ();
 sg13g2_decap_4 FILLER_20_76 ();
 sg13g2_fill_1 FILLER_20_80 ();
 sg13g2_decap_4 FILLER_20_86 ();
 sg13g2_fill_1 FILLER_20_90 ();
 sg13g2_fill_1 FILLER_20_110 ();
 sg13g2_decap_8 FILLER_20_129 ();
 sg13g2_fill_2 FILLER_20_136 ();
 sg13g2_fill_1 FILLER_20_138 ();
 sg13g2_fill_1 FILLER_20_155 ();
 sg13g2_fill_1 FILLER_20_160 ();
 sg13g2_fill_1 FILLER_20_174 ();
 sg13g2_fill_1 FILLER_20_180 ();
 sg13g2_fill_2 FILLER_20_202 ();
 sg13g2_fill_2 FILLER_20_213 ();
 sg13g2_fill_1 FILLER_20_215 ();
 sg13g2_decap_4 FILLER_20_221 ();
 sg13g2_fill_2 FILLER_20_233 ();
 sg13g2_decap_8 FILLER_20_249 ();
 sg13g2_decap_4 FILLER_20_256 ();
 sg13g2_fill_1 FILLER_20_270 ();
 sg13g2_fill_2 FILLER_20_287 ();
 sg13g2_fill_1 FILLER_20_289 ();
 sg13g2_decap_8 FILLER_20_300 ();
 sg13g2_fill_2 FILLER_20_307 ();
 sg13g2_fill_2 FILLER_20_318 ();
 sg13g2_fill_1 FILLER_20_320 ();
 sg13g2_decap_4 FILLER_20_326 ();
 sg13g2_decap_8 FILLER_20_334 ();
 sg13g2_decap_8 FILLER_20_341 ();
 sg13g2_decap_8 FILLER_20_348 ();
 sg13g2_decap_8 FILLER_20_355 ();
 sg13g2_decap_8 FILLER_20_362 ();
 sg13g2_decap_8 FILLER_20_369 ();
 sg13g2_decap_8 FILLER_20_376 ();
 sg13g2_decap_8 FILLER_20_383 ();
 sg13g2_decap_8 FILLER_20_390 ();
 sg13g2_decap_8 FILLER_20_397 ();
 sg13g2_decap_4 FILLER_20_404 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_fill_2 FILLER_21_49 ();
 sg13g2_fill_1 FILLER_21_51 ();
 sg13g2_decap_4 FILLER_21_66 ();
 sg13g2_fill_1 FILLER_21_70 ();
 sg13g2_fill_2 FILLER_21_89 ();
 sg13g2_fill_1 FILLER_21_91 ();
 sg13g2_fill_2 FILLER_21_103 ();
 sg13g2_fill_2 FILLER_21_110 ();
 sg13g2_decap_4 FILLER_21_120 ();
 sg13g2_fill_2 FILLER_21_124 ();
 sg13g2_decap_8 FILLER_21_141 ();
 sg13g2_fill_1 FILLER_21_148 ();
 sg13g2_fill_2 FILLER_21_189 ();
 sg13g2_decap_4 FILLER_21_194 ();
 sg13g2_fill_2 FILLER_21_198 ();
 sg13g2_fill_2 FILLER_21_210 ();
 sg13g2_fill_2 FILLER_21_227 ();
 sg13g2_fill_2 FILLER_21_233 ();
 sg13g2_decap_8 FILLER_21_249 ();
 sg13g2_decap_4 FILLER_21_256 ();
 sg13g2_fill_2 FILLER_21_268 ();
 sg13g2_fill_2 FILLER_21_287 ();
 sg13g2_fill_2 FILLER_21_295 ();
 sg13g2_decap_4 FILLER_21_307 ();
 sg13g2_fill_2 FILLER_21_311 ();
 sg13g2_fill_1 FILLER_21_318 ();
 sg13g2_fill_1 FILLER_21_343 ();
 sg13g2_decap_8 FILLER_21_357 ();
 sg13g2_decap_8 FILLER_21_364 ();
 sg13g2_decap_8 FILLER_21_371 ();
 sg13g2_decap_8 FILLER_21_378 ();
 sg13g2_decap_8 FILLER_21_385 ();
 sg13g2_decap_8 FILLER_21_392 ();
 sg13g2_decap_8 FILLER_21_399 ();
 sg13g2_fill_2 FILLER_21_406 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_fill_1 FILLER_22_42 ();
 sg13g2_fill_2 FILLER_22_56 ();
 sg13g2_fill_1 FILLER_22_58 ();
 sg13g2_fill_1 FILLER_22_69 ();
 sg13g2_decap_8 FILLER_22_75 ();
 sg13g2_decap_4 FILLER_22_87 ();
 sg13g2_fill_2 FILLER_22_91 ();
 sg13g2_fill_2 FILLER_22_113 ();
 sg13g2_decap_8 FILLER_22_133 ();
 sg13g2_decap_8 FILLER_22_140 ();
 sg13g2_fill_1 FILLER_22_147 ();
 sg13g2_decap_8 FILLER_22_152 ();
 sg13g2_fill_1 FILLER_22_159 ();
 sg13g2_decap_8 FILLER_22_176 ();
 sg13g2_fill_2 FILLER_22_183 ();
 sg13g2_fill_1 FILLER_22_185 ();
 sg13g2_fill_1 FILLER_22_202 ();
 sg13g2_decap_4 FILLER_22_208 ();
 sg13g2_fill_1 FILLER_22_212 ();
 sg13g2_decap_4 FILLER_22_226 ();
 sg13g2_fill_1 FILLER_22_234 ();
 sg13g2_decap_4 FILLER_22_242 ();
 sg13g2_decap_4 FILLER_22_270 ();
 sg13g2_fill_1 FILLER_22_274 ();
 sg13g2_fill_2 FILLER_22_285 ();
 sg13g2_fill_1 FILLER_22_320 ();
 sg13g2_decap_4 FILLER_22_325 ();
 sg13g2_fill_1 FILLER_22_329 ();
 sg13g2_decap_8 FILLER_22_356 ();
 sg13g2_decap_8 FILLER_22_363 ();
 sg13g2_decap_8 FILLER_22_370 ();
 sg13g2_decap_8 FILLER_22_377 ();
 sg13g2_decap_8 FILLER_22_384 ();
 sg13g2_decap_8 FILLER_22_391 ();
 sg13g2_decap_8 FILLER_22_398 ();
 sg13g2_decap_4 FILLER_22_405 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_4 FILLER_23_49 ();
 sg13g2_fill_1 FILLER_23_58 ();
 sg13g2_decap_8 FILLER_23_64 ();
 sg13g2_fill_2 FILLER_23_71 ();
 sg13g2_fill_1 FILLER_23_73 ();
 sg13g2_fill_2 FILLER_23_80 ();
 sg13g2_decap_4 FILLER_23_90 ();
 sg13g2_fill_1 FILLER_23_111 ();
 sg13g2_fill_1 FILLER_23_122 ();
 sg13g2_decap_8 FILLER_23_166 ();
 sg13g2_decap_4 FILLER_23_173 ();
 sg13g2_fill_2 FILLER_23_177 ();
 sg13g2_fill_1 FILLER_23_187 ();
 sg13g2_fill_2 FILLER_23_208 ();
 sg13g2_fill_1 FILLER_23_210 ();
 sg13g2_fill_2 FILLER_23_219 ();
 sg13g2_fill_1 FILLER_23_221 ();
 sg13g2_fill_1 FILLER_23_243 ();
 sg13g2_decap_4 FILLER_23_249 ();
 sg13g2_fill_2 FILLER_23_253 ();
 sg13g2_decap_4 FILLER_23_288 ();
 sg13g2_fill_2 FILLER_23_292 ();
 sg13g2_decap_4 FILLER_23_299 ();
 sg13g2_fill_1 FILLER_23_303 ();
 sg13g2_fill_2 FILLER_23_319 ();
 sg13g2_fill_2 FILLER_23_327 ();
 sg13g2_fill_1 FILLER_23_329 ();
 sg13g2_decap_8 FILLER_23_341 ();
 sg13g2_decap_8 FILLER_23_348 ();
 sg13g2_decap_8 FILLER_23_355 ();
 sg13g2_decap_4 FILLER_23_362 ();
 sg13g2_fill_1 FILLER_23_366 ();
 sg13g2_decap_8 FILLER_23_375 ();
 sg13g2_decap_8 FILLER_23_387 ();
 sg13g2_decap_8 FILLER_23_394 ();
 sg13g2_decap_8 FILLER_23_401 ();
 sg13g2_fill_1 FILLER_23_408 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_4 FILLER_24_42 ();
 sg13g2_fill_1 FILLER_24_60 ();
 sg13g2_fill_1 FILLER_24_76 ();
 sg13g2_decap_8 FILLER_24_83 ();
 sg13g2_fill_2 FILLER_24_90 ();
 sg13g2_fill_2 FILLER_24_102 ();
 sg13g2_fill_1 FILLER_24_104 ();
 sg13g2_fill_1 FILLER_24_111 ();
 sg13g2_fill_1 FILLER_24_135 ();
 sg13g2_decap_4 FILLER_24_141 ();
 sg13g2_fill_1 FILLER_24_145 ();
 sg13g2_decap_4 FILLER_24_163 ();
 sg13g2_fill_1 FILLER_24_167 ();
 sg13g2_decap_8 FILLER_24_181 ();
 sg13g2_decap_4 FILLER_24_188 ();
 sg13g2_fill_1 FILLER_24_192 ();
 sg13g2_decap_4 FILLER_24_211 ();
 sg13g2_decap_8 FILLER_24_223 ();
 sg13g2_decap_4 FILLER_24_230 ();
 sg13g2_decap_4 FILLER_24_260 ();
 sg13g2_decap_4 FILLER_24_274 ();
 sg13g2_fill_1 FILLER_24_291 ();
 sg13g2_decap_4 FILLER_24_296 ();
 sg13g2_decap_8 FILLER_24_322 ();
 sg13g2_fill_2 FILLER_24_329 ();
 sg13g2_fill_1 FILLER_24_331 ();
 sg13g2_decap_8 FILLER_24_336 ();
 sg13g2_decap_8 FILLER_24_343 ();
 sg13g2_decap_8 FILLER_24_350 ();
 sg13g2_decap_8 FILLER_24_357 ();
 sg13g2_fill_2 FILLER_24_364 ();
 sg13g2_fill_1 FILLER_24_366 ();
 sg13g2_fill_1 FILLER_24_380 ();
 sg13g2_decap_8 FILLER_24_397 ();
 sg13g2_decap_4 FILLER_24_404 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_4 FILLER_25_42 ();
 sg13g2_fill_1 FILLER_25_46 ();
 sg13g2_fill_1 FILLER_25_57 ();
 sg13g2_fill_1 FILLER_25_63 ();
 sg13g2_decap_4 FILLER_25_74 ();
 sg13g2_fill_2 FILLER_25_78 ();
 sg13g2_decap_8 FILLER_25_89 ();
 sg13g2_decap_4 FILLER_25_100 ();
 sg13g2_decap_8 FILLER_25_116 ();
 sg13g2_decap_4 FILLER_25_123 ();
 sg13g2_fill_2 FILLER_25_135 ();
 sg13g2_fill_1 FILLER_25_137 ();
 sg13g2_fill_1 FILLER_25_143 ();
 sg13g2_decap_4 FILLER_25_149 ();
 sg13g2_fill_2 FILLER_25_165 ();
 sg13g2_fill_2 FILLER_25_195 ();
 sg13g2_fill_1 FILLER_25_197 ();
 sg13g2_fill_1 FILLER_25_203 ();
 sg13g2_decap_8 FILLER_25_213 ();
 sg13g2_decap_4 FILLER_25_220 ();
 sg13g2_fill_2 FILLER_25_224 ();
 sg13g2_fill_1 FILLER_25_231 ();
 sg13g2_fill_2 FILLER_25_251 ();
 sg13g2_fill_1 FILLER_25_261 ();
 sg13g2_fill_2 FILLER_25_276 ();
 sg13g2_fill_1 FILLER_25_278 ();
 sg13g2_fill_1 FILLER_25_300 ();
 sg13g2_fill_1 FILLER_25_305 ();
 sg13g2_fill_2 FILLER_25_326 ();
 sg13g2_decap_8 FILLER_25_344 ();
 sg13g2_decap_8 FILLER_25_351 ();
 sg13g2_decap_8 FILLER_25_358 ();
 sg13g2_decap_4 FILLER_25_365 ();
 sg13g2_fill_1 FILLER_25_369 ();
 sg13g2_fill_1 FILLER_25_379 ();
 sg13g2_fill_2 FILLER_25_394 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_4 FILLER_26_56 ();
 sg13g2_fill_1 FILLER_26_60 ();
 sg13g2_fill_1 FILLER_26_86 ();
 sg13g2_fill_2 FILLER_26_112 ();
 sg13g2_fill_1 FILLER_26_114 ();
 sg13g2_decap_8 FILLER_26_125 ();
 sg13g2_fill_1 FILLER_26_132 ();
 sg13g2_fill_1 FILLER_26_138 ();
 sg13g2_decap_4 FILLER_26_152 ();
 sg13g2_fill_1 FILLER_26_164 ();
 sg13g2_fill_1 FILLER_26_177 ();
 sg13g2_decap_8 FILLER_26_243 ();
 sg13g2_decap_4 FILLER_26_250 ();
 sg13g2_decap_4 FILLER_26_271 ();
 sg13g2_decap_8 FILLER_26_287 ();
 sg13g2_fill_1 FILLER_26_294 ();
 sg13g2_fill_1 FILLER_26_298 ();
 sg13g2_decap_8 FILLER_26_304 ();
 sg13g2_fill_2 FILLER_26_311 ();
 sg13g2_fill_1 FILLER_26_313 ();
 sg13g2_fill_1 FILLER_26_319 ();
 sg13g2_fill_2 FILLER_26_324 ();
 sg13g2_fill_1 FILLER_26_331 ();
 sg13g2_decap_8 FILLER_26_337 ();
 sg13g2_decap_8 FILLER_26_344 ();
 sg13g2_decap_8 FILLER_26_351 ();
 sg13g2_fill_1 FILLER_26_358 ();
 sg13g2_fill_2 FILLER_26_407 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_fill_1 FILLER_27_42 ();
 sg13g2_decap_4 FILLER_27_85 ();
 sg13g2_fill_1 FILLER_27_89 ();
 sg13g2_fill_2 FILLER_27_98 ();
 sg13g2_fill_1 FILLER_27_127 ();
 sg13g2_decap_8 FILLER_27_144 ();
 sg13g2_fill_1 FILLER_27_151 ();
 sg13g2_fill_2 FILLER_27_162 ();
 sg13g2_fill_2 FILLER_27_180 ();
 sg13g2_fill_2 FILLER_27_187 ();
 sg13g2_fill_1 FILLER_27_189 ();
 sg13g2_fill_2 FILLER_27_198 ();
 sg13g2_decap_4 FILLER_27_208 ();
 sg13g2_decap_8 FILLER_27_233 ();
 sg13g2_decap_4 FILLER_27_273 ();
 sg13g2_decap_4 FILLER_27_281 ();
 sg13g2_fill_1 FILLER_27_285 ();
 sg13g2_decap_8 FILLER_27_342 ();
 sg13g2_decap_8 FILLER_27_349 ();
 sg13g2_fill_2 FILLER_27_356 ();
 sg13g2_fill_1 FILLER_27_358 ();
 sg13g2_decap_8 FILLER_27_363 ();
 sg13g2_fill_1 FILLER_27_370 ();
 sg13g2_fill_1 FILLER_27_386 ();
 sg13g2_decap_4 FILLER_27_391 ();
 sg13g2_fill_1 FILLER_27_395 ();
 sg13g2_fill_1 FILLER_27_408 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_4 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_57 ();
 sg13g2_decap_4 FILLER_28_64 ();
 sg13g2_fill_1 FILLER_28_68 ();
 sg13g2_decap_4 FILLER_28_74 ();
 sg13g2_fill_1 FILLER_28_78 ();
 sg13g2_fill_2 FILLER_28_84 ();
 sg13g2_decap_8 FILLER_28_105 ();
 sg13g2_fill_2 FILLER_28_112 ();
 sg13g2_fill_2 FILLER_28_132 ();
 sg13g2_fill_2 FILLER_28_157 ();
 sg13g2_fill_2 FILLER_28_170 ();
 sg13g2_fill_1 FILLER_28_172 ();
 sg13g2_fill_2 FILLER_28_185 ();
 sg13g2_fill_2 FILLER_28_192 ();
 sg13g2_fill_1 FILLER_28_194 ();
 sg13g2_decap_4 FILLER_28_215 ();
 sg13g2_fill_2 FILLER_28_227 ();
 sg13g2_fill_1 FILLER_28_229 ();
 sg13g2_fill_2 FILLER_28_258 ();
 sg13g2_fill_1 FILLER_28_260 ();
 sg13g2_fill_2 FILLER_28_272 ();
 sg13g2_fill_1 FILLER_28_282 ();
 sg13g2_decap_8 FILLER_28_295 ();
 sg13g2_decap_4 FILLER_28_302 ();
 sg13g2_fill_1 FILLER_28_306 ();
 sg13g2_decap_8 FILLER_28_321 ();
 sg13g2_fill_2 FILLER_28_328 ();
 sg13g2_fill_1 FILLER_28_330 ();
 sg13g2_decap_8 FILLER_28_335 ();
 sg13g2_decap_8 FILLER_28_342 ();
 sg13g2_decap_4 FILLER_28_349 ();
 sg13g2_fill_2 FILLER_28_366 ();
 sg13g2_fill_1 FILLER_28_381 ();
 sg13g2_fill_2 FILLER_28_387 ();
 sg13g2_fill_1 FILLER_28_408 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_fill_1 FILLER_29_65 ();
 sg13g2_fill_2 FILLER_29_87 ();
 sg13g2_decap_4 FILLER_29_101 ();
 sg13g2_decap_4 FILLER_29_119 ();
 sg13g2_fill_1 FILLER_29_123 ();
 sg13g2_fill_2 FILLER_29_129 ();
 sg13g2_fill_1 FILLER_29_131 ();
 sg13g2_fill_2 FILLER_29_140 ();
 sg13g2_decap_8 FILLER_29_148 ();
 sg13g2_fill_2 FILLER_29_179 ();
 sg13g2_decap_8 FILLER_29_189 ();
 sg13g2_decap_4 FILLER_29_200 ();
 sg13g2_fill_2 FILLER_29_204 ();
 sg13g2_decap_8 FILLER_29_214 ();
 sg13g2_decap_8 FILLER_29_229 ();
 sg13g2_decap_4 FILLER_29_236 ();
 sg13g2_decap_8 FILLER_29_252 ();
 sg13g2_fill_2 FILLER_29_259 ();
 sg13g2_fill_2 FILLER_29_269 ();
 sg13g2_fill_1 FILLER_29_271 ();
 sg13g2_fill_2 FILLER_29_283 ();
 sg13g2_decap_8 FILLER_29_308 ();
 sg13g2_fill_1 FILLER_29_315 ();
 sg13g2_decap_8 FILLER_29_333 ();
 sg13g2_decap_8 FILLER_29_340 ();
 sg13g2_decap_8 FILLER_29_347 ();
 sg13g2_decap_4 FILLER_29_354 ();
 sg13g2_fill_1 FILLER_29_358 ();
 sg13g2_decap_8 FILLER_29_365 ();
 sg13g2_decap_4 FILLER_29_372 ();
 sg13g2_fill_1 FILLER_29_376 ();
 sg13g2_fill_1 FILLER_29_394 ();
 sg13g2_fill_2 FILLER_29_399 ();
 sg13g2_fill_2 FILLER_29_406 ();
 sg13g2_fill_1 FILLER_29_408 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_4 FILLER_30_42 ();
 sg13g2_fill_1 FILLER_30_46 ();
 sg13g2_decap_8 FILLER_30_55 ();
 sg13g2_decap_8 FILLER_30_62 ();
 sg13g2_decap_8 FILLER_30_69 ();
 sg13g2_fill_2 FILLER_30_81 ();
 sg13g2_fill_1 FILLER_30_91 ();
 sg13g2_fill_2 FILLER_30_131 ();
 sg13g2_fill_1 FILLER_30_133 ();
 sg13g2_fill_1 FILLER_30_146 ();
 sg13g2_fill_2 FILLER_30_156 ();
 sg13g2_fill_1 FILLER_30_158 ();
 sg13g2_decap_8 FILLER_30_167 ();
 sg13g2_decap_8 FILLER_30_174 ();
 sg13g2_fill_2 FILLER_30_181 ();
 sg13g2_fill_1 FILLER_30_194 ();
 sg13g2_decap_8 FILLER_30_211 ();
 sg13g2_fill_2 FILLER_30_218 ();
 sg13g2_fill_1 FILLER_30_220 ();
 sg13g2_decap_4 FILLER_30_227 ();
 sg13g2_fill_2 FILLER_30_231 ();
 sg13g2_fill_1 FILLER_30_256 ();
 sg13g2_fill_2 FILLER_30_271 ();
 sg13g2_fill_2 FILLER_30_279 ();
 sg13g2_fill_1 FILLER_30_281 ();
 sg13g2_fill_2 FILLER_30_295 ();
 sg13g2_fill_1 FILLER_30_297 ();
 sg13g2_fill_2 FILLER_30_312 ();
 sg13g2_decap_4 FILLER_30_321 ();
 sg13g2_fill_2 FILLER_30_325 ();
 sg13g2_fill_2 FILLER_30_339 ();
 sg13g2_fill_1 FILLER_30_349 ();
 sg13g2_decap_4 FILLER_30_380 ();
 sg13g2_fill_1 FILLER_30_384 ();
 sg13g2_fill_1 FILLER_30_399 ();
 sg13g2_fill_1 FILLER_30_408 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_4 FILLER_31_42 ();
 sg13g2_fill_2 FILLER_31_71 ();
 sg13g2_decap_4 FILLER_31_82 ();
 sg13g2_fill_1 FILLER_31_96 ();
 sg13g2_decap_8 FILLER_31_104 ();
 sg13g2_decap_4 FILLER_31_111 ();
 sg13g2_fill_2 FILLER_31_120 ();
 sg13g2_fill_1 FILLER_31_127 ();
 sg13g2_decap_8 FILLER_31_137 ();
 sg13g2_fill_2 FILLER_31_144 ();
 sg13g2_fill_1 FILLER_31_146 ();
 sg13g2_decap_8 FILLER_31_158 ();
 sg13g2_decap_4 FILLER_31_165 ();
 sg13g2_fill_2 FILLER_31_185 ();
 sg13g2_fill_1 FILLER_31_187 ();
 sg13g2_decap_8 FILLER_31_192 ();
 sg13g2_fill_1 FILLER_31_244 ();
 sg13g2_decap_4 FILLER_31_253 ();
 sg13g2_decap_4 FILLER_31_265 ();
 sg13g2_decap_8 FILLER_31_279 ();
 sg13g2_fill_1 FILLER_31_286 ();
 sg13g2_fill_1 FILLER_31_305 ();
 sg13g2_fill_1 FILLER_31_325 ();
 sg13g2_decap_4 FILLER_31_339 ();
 sg13g2_fill_1 FILLER_31_343 ();
 sg13g2_fill_2 FILLER_31_353 ();
 sg13g2_fill_2 FILLER_31_364 ();
 sg13g2_fill_2 FILLER_31_376 ();
 sg13g2_fill_1 FILLER_31_378 ();
 sg13g2_fill_1 FILLER_31_399 ();
 sg13g2_fill_1 FILLER_31_408 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_4 FILLER_32_49 ();
 sg13g2_fill_1 FILLER_32_53 ();
 sg13g2_fill_2 FILLER_32_79 ();
 sg13g2_fill_1 FILLER_32_93 ();
 sg13g2_fill_1 FILLER_32_102 ();
 sg13g2_fill_2 FILLER_32_108 ();
 sg13g2_fill_1 FILLER_32_110 ();
 sg13g2_fill_1 FILLER_32_119 ();
 sg13g2_fill_2 FILLER_32_125 ();
 sg13g2_fill_1 FILLER_32_127 ();
 sg13g2_fill_2 FILLER_32_144 ();
 sg13g2_fill_1 FILLER_32_146 ();
 sg13g2_fill_2 FILLER_32_151 ();
 sg13g2_fill_1 FILLER_32_153 ();
 sg13g2_fill_2 FILLER_32_164 ();
 sg13g2_fill_1 FILLER_32_166 ();
 sg13g2_fill_2 FILLER_32_175 ();
 sg13g2_fill_2 FILLER_32_185 ();
 sg13g2_fill_1 FILLER_32_187 ();
 sg13g2_decap_8 FILLER_32_214 ();
 sg13g2_decap_4 FILLER_32_221 ();
 sg13g2_fill_2 FILLER_32_225 ();
 sg13g2_decap_8 FILLER_32_257 ();
 sg13g2_decap_4 FILLER_32_264 ();
 sg13g2_fill_1 FILLER_32_268 ();
 sg13g2_fill_2 FILLER_32_278 ();
 sg13g2_decap_4 FILLER_32_295 ();
 sg13g2_fill_2 FILLER_32_306 ();
 sg13g2_fill_2 FILLER_32_328 ();
 sg13g2_fill_2 FILLER_32_338 ();
 sg13g2_fill_1 FILLER_32_340 ();
 sg13g2_fill_2 FILLER_32_356 ();
 sg13g2_fill_2 FILLER_32_368 ();
 sg13g2_fill_1 FILLER_32_370 ();
 sg13g2_fill_2 FILLER_32_383 ();
 sg13g2_fill_1 FILLER_32_385 ();
 sg13g2_fill_2 FILLER_32_407 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_fill_1 FILLER_33_56 ();
 sg13g2_fill_2 FILLER_33_61 ();
 sg13g2_fill_1 FILLER_33_63 ();
 sg13g2_decap_4 FILLER_33_69 ();
 sg13g2_fill_1 FILLER_33_73 ();
 sg13g2_decap_4 FILLER_33_94 ();
 sg13g2_fill_1 FILLER_33_98 ();
 sg13g2_fill_2 FILLER_33_115 ();
 sg13g2_fill_1 FILLER_33_117 ();
 sg13g2_fill_2 FILLER_33_130 ();
 sg13g2_fill_1 FILLER_33_136 ();
 sg13g2_fill_1 FILLER_33_152 ();
 sg13g2_fill_1 FILLER_33_158 ();
 sg13g2_fill_1 FILLER_33_164 ();
 sg13g2_fill_2 FILLER_33_173 ();
 sg13g2_fill_1 FILLER_33_175 ();
 sg13g2_fill_2 FILLER_33_212 ();
 sg13g2_fill_1 FILLER_33_223 ();
 sg13g2_decap_4 FILLER_33_274 ();
 sg13g2_fill_2 FILLER_33_278 ();
 sg13g2_fill_2 FILLER_33_286 ();
 sg13g2_decap_8 FILLER_33_301 ();
 sg13g2_decap_8 FILLER_33_308 ();
 sg13g2_fill_2 FILLER_33_324 ();
 sg13g2_fill_1 FILLER_33_326 ();
 sg13g2_decap_4 FILLER_33_340 ();
 sg13g2_decap_4 FILLER_33_349 ();
 sg13g2_fill_2 FILLER_33_374 ();
 sg13g2_fill_1 FILLER_33_376 ();
 sg13g2_decap_4 FILLER_33_384 ();
 sg13g2_decap_4 FILLER_33_396 ();
 sg13g2_fill_1 FILLER_33_408 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_4 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_72 ();
 sg13g2_decap_8 FILLER_34_79 ();
 sg13g2_decap_4 FILLER_34_86 ();
 sg13g2_fill_2 FILLER_34_90 ();
 sg13g2_fill_2 FILLER_34_100 ();
 sg13g2_fill_1 FILLER_34_102 ();
 sg13g2_fill_2 FILLER_34_115 ();
 sg13g2_fill_1 FILLER_34_117 ();
 sg13g2_decap_4 FILLER_34_123 ();
 sg13g2_fill_1 FILLER_34_127 ();
 sg13g2_fill_1 FILLER_34_140 ();
 sg13g2_decap_8 FILLER_34_147 ();
 sg13g2_decap_4 FILLER_34_154 ();
 sg13g2_fill_1 FILLER_34_158 ();
 sg13g2_fill_1 FILLER_34_167 ();
 sg13g2_fill_2 FILLER_34_188 ();
 sg13g2_fill_1 FILLER_34_190 ();
 sg13g2_fill_1 FILLER_34_196 ();
 sg13g2_fill_2 FILLER_34_204 ();
 sg13g2_fill_1 FILLER_34_206 ();
 sg13g2_fill_2 FILLER_34_215 ();
 sg13g2_decap_8 FILLER_34_229 ();
 sg13g2_decap_8 FILLER_34_236 ();
 sg13g2_decap_8 FILLER_34_248 ();
 sg13g2_fill_1 FILLER_34_255 ();
 sg13g2_decap_4 FILLER_34_274 ();
 sg13g2_fill_1 FILLER_34_286 ();
 sg13g2_decap_8 FILLER_34_297 ();
 sg13g2_decap_4 FILLER_34_304 ();
 sg13g2_fill_2 FILLER_34_330 ();
 sg13g2_decap_4 FILLER_34_337 ();
 sg13g2_fill_2 FILLER_34_363 ();
 sg13g2_decap_8 FILLER_34_377 ();
 sg13g2_fill_2 FILLER_34_384 ();
 sg13g2_fill_2 FILLER_34_394 ();
 sg13g2_fill_1 FILLER_34_401 ();
 sg13g2_fill_2 FILLER_34_407 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_fill_2 FILLER_35_42 ();
 sg13g2_fill_2 FILLER_35_76 ();
 sg13g2_fill_1 FILLER_35_105 ();
 sg13g2_fill_2 FILLER_35_130 ();
 sg13g2_decap_8 FILLER_35_142 ();
 sg13g2_fill_2 FILLER_35_160 ();
 sg13g2_fill_2 FILLER_35_183 ();
 sg13g2_fill_1 FILLER_35_185 ();
 sg13g2_fill_1 FILLER_35_205 ();
 sg13g2_decap_8 FILLER_35_214 ();
 sg13g2_decap_8 FILLER_35_221 ();
 sg13g2_decap_4 FILLER_35_228 ();
 sg13g2_fill_2 FILLER_35_232 ();
 sg13g2_fill_1 FILLER_35_243 ();
 sg13g2_decap_8 FILLER_35_266 ();
 sg13g2_fill_1 FILLER_35_273 ();
 sg13g2_decap_4 FILLER_35_284 ();
 sg13g2_fill_1 FILLER_35_314 ();
 sg13g2_fill_2 FILLER_35_340 ();
 sg13g2_decap_8 FILLER_35_347 ();
 sg13g2_decap_8 FILLER_35_365 ();
 sg13g2_fill_2 FILLER_35_378 ();
 sg13g2_fill_2 FILLER_35_388 ();
 sg13g2_fill_1 FILLER_35_390 ();
 sg13g2_fill_1 FILLER_35_399 ();
 sg13g2_fill_1 FILLER_35_408 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_fill_1 FILLER_36_14 ();
 sg13g2_decap_4 FILLER_36_48 ();
 sg13g2_decap_4 FILLER_36_62 ();
 sg13g2_fill_2 FILLER_36_76 ();
 sg13g2_fill_1 FILLER_36_78 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_fill_2 FILLER_36_98 ();
 sg13g2_fill_2 FILLER_36_114 ();
 sg13g2_decap_4 FILLER_36_120 ();
 sg13g2_fill_1 FILLER_36_124 ();
 sg13g2_fill_1 FILLER_36_137 ();
 sg13g2_fill_1 FILLER_36_156 ();
 sg13g2_fill_2 FILLER_36_167 ();
 sg13g2_fill_1 FILLER_36_169 ();
 sg13g2_decap_4 FILLER_36_186 ();
 sg13g2_fill_2 FILLER_36_195 ();
 sg13g2_fill_1 FILLER_36_197 ();
 sg13g2_decap_8 FILLER_36_252 ();
 sg13g2_fill_2 FILLER_36_259 ();
 sg13g2_fill_1 FILLER_36_281 ();
 sg13g2_decap_8 FILLER_36_295 ();
 sg13g2_fill_2 FILLER_36_311 ();
 sg13g2_fill_1 FILLER_36_313 ();
 sg13g2_fill_1 FILLER_36_327 ();
 sg13g2_fill_2 FILLER_36_337 ();
 sg13g2_fill_1 FILLER_36_339 ();
 sg13g2_decap_4 FILLER_36_348 ();
 sg13g2_fill_1 FILLER_36_352 ();
 sg13g2_decap_4 FILLER_36_364 ();
 sg13g2_decap_4 FILLER_36_376 ();
 sg13g2_fill_1 FILLER_36_380 ();
 sg13g2_decap_4 FILLER_36_390 ();
 sg13g2_fill_1 FILLER_36_394 ();
 sg13g2_fill_1 FILLER_36_408 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_4 FILLER_37_7 ();
 sg13g2_fill_2 FILLER_37_19 ();
 sg13g2_fill_2 FILLER_37_36 ();
 sg13g2_fill_1 FILLER_37_51 ();
 sg13g2_fill_1 FILLER_37_75 ();
 sg13g2_decap_4 FILLER_37_81 ();
 sg13g2_fill_2 FILLER_37_85 ();
 sg13g2_decap_4 FILLER_37_113 ();
 sg13g2_decap_8 FILLER_37_135 ();
 sg13g2_fill_1 FILLER_37_142 ();
 sg13g2_fill_1 FILLER_37_148 ();
 sg13g2_fill_1 FILLER_37_165 ();
 sg13g2_decap_4 FILLER_37_175 ();
 sg13g2_decap_4 FILLER_37_184 ();
 sg13g2_decap_4 FILLER_37_203 ();
 sg13g2_fill_1 FILLER_37_207 ();
 sg13g2_fill_1 FILLER_37_212 ();
 sg13g2_fill_2 FILLER_37_217 ();
 sg13g2_fill_1 FILLER_37_219 ();
 sg13g2_fill_2 FILLER_37_228 ();
 sg13g2_decap_4 FILLER_37_248 ();
 sg13g2_fill_1 FILLER_37_252 ();
 sg13g2_fill_1 FILLER_37_273 ();
 sg13g2_fill_1 FILLER_37_284 ();
 sg13g2_decap_4 FILLER_37_301 ();
 sg13g2_fill_2 FILLER_37_313 ();
 sg13g2_fill_2 FILLER_37_335 ();
 sg13g2_fill_1 FILLER_37_337 ();
 sg13g2_decap_8 FILLER_37_348 ();
 sg13g2_decap_4 FILLER_37_355 ();
 sg13g2_fill_2 FILLER_37_379 ();
 sg13g2_fill_1 FILLER_37_381 ();
 sg13g2_decap_4 FILLER_37_387 ();
 sg13g2_fill_2 FILLER_37_407 ();
 sg13g2_decap_4 FILLER_38_0 ();
 sg13g2_fill_2 FILLER_38_4 ();
 sg13g2_decap_8 FILLER_38_24 ();
 sg13g2_decap_4 FILLER_38_41 ();
 sg13g2_fill_2 FILLER_38_45 ();
 sg13g2_decap_8 FILLER_38_51 ();
 sg13g2_decap_4 FILLER_38_63 ();
 sg13g2_decap_4 FILLER_38_78 ();
 sg13g2_decap_4 FILLER_38_94 ();
 sg13g2_fill_2 FILLER_38_102 ();
 sg13g2_fill_2 FILLER_38_117 ();
 sg13g2_fill_2 FILLER_38_127 ();
 sg13g2_fill_2 FILLER_38_136 ();
 sg13g2_decap_8 FILLER_38_157 ();
 sg13g2_fill_2 FILLER_38_168 ();
 sg13g2_decap_4 FILLER_38_175 ();
 sg13g2_fill_1 FILLER_38_179 ();
 sg13g2_decap_8 FILLER_38_223 ();
 sg13g2_decap_8 FILLER_38_230 ();
 sg13g2_fill_1 FILLER_38_237 ();
 sg13g2_fill_1 FILLER_38_258 ();
 sg13g2_fill_1 FILLER_38_279 ();
 sg13g2_fill_2 FILLER_38_285 ();
 sg13g2_fill_1 FILLER_38_287 ();
 sg13g2_decap_8 FILLER_38_292 ();
 sg13g2_fill_2 FILLER_38_299 ();
 sg13g2_decap_8 FILLER_38_308 ();
 sg13g2_fill_1 FILLER_38_315 ();
 sg13g2_fill_2 FILLER_38_336 ();
 sg13g2_decap_4 FILLER_38_362 ();
 sg13g2_fill_2 FILLER_38_366 ();
 sg13g2_decap_4 FILLER_38_381 ();
 sg13g2_fill_1 FILLER_38_385 ();
 sg13g2_fill_2 FILLER_38_398 ();
 sg13g2_fill_1 FILLER_38_408 ();
 sg13g2_fill_2 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_10 ();
 sg13g2_fill_1 FILLER_39_62 ();
 sg13g2_decap_4 FILLER_39_69 ();
 sg13g2_fill_1 FILLER_39_73 ();
 sg13g2_decap_4 FILLER_39_79 ();
 sg13g2_fill_1 FILLER_39_83 ();
 sg13g2_decap_4 FILLER_39_92 ();
 sg13g2_fill_1 FILLER_39_96 ();
 sg13g2_fill_2 FILLER_39_109 ();
 sg13g2_fill_1 FILLER_39_111 ();
 sg13g2_decap_8 FILLER_39_118 ();
 sg13g2_fill_2 FILLER_39_125 ();
 sg13g2_fill_1 FILLER_39_127 ();
 sg13g2_fill_1 FILLER_39_132 ();
 sg13g2_fill_1 FILLER_39_143 ();
 sg13g2_decap_4 FILLER_39_151 ();
 sg13g2_fill_2 FILLER_39_155 ();
 sg13g2_decap_4 FILLER_39_204 ();
 sg13g2_fill_2 FILLER_39_208 ();
 sg13g2_decap_4 FILLER_39_215 ();
 sg13g2_fill_1 FILLER_39_219 ();
 sg13g2_fill_1 FILLER_39_237 ();
 sg13g2_decap_4 FILLER_39_249 ();
 sg13g2_fill_1 FILLER_39_253 ();
 sg13g2_decap_4 FILLER_39_276 ();
 sg13g2_fill_1 FILLER_39_325 ();
 sg13g2_fill_1 FILLER_39_331 ();
 sg13g2_decap_8 FILLER_39_348 ();
 sg13g2_fill_1 FILLER_39_355 ();
 sg13g2_fill_1 FILLER_39_384 ();
 sg13g2_fill_2 FILLER_39_393 ();
 sg13g2_decap_4 FILLER_39_405 ();
 sg13g2_decap_4 FILLER_40_0 ();
 sg13g2_fill_2 FILLER_40_4 ();
 sg13g2_decap_4 FILLER_40_22 ();
 sg13g2_fill_1 FILLER_40_26 ();
 sg13g2_fill_1 FILLER_40_33 ();
 sg13g2_decap_4 FILLER_40_44 ();
 sg13g2_fill_1 FILLER_40_48 ();
 sg13g2_decap_4 FILLER_40_54 ();
 sg13g2_fill_1 FILLER_40_58 ();
 sg13g2_decap_4 FILLER_40_69 ();
 sg13g2_fill_1 FILLER_40_73 ();
 sg13g2_fill_2 FILLER_40_106 ();
 sg13g2_fill_1 FILLER_40_108 ();
 sg13g2_fill_1 FILLER_40_134 ();
 sg13g2_fill_1 FILLER_40_141 ();
 sg13g2_decap_4 FILLER_40_147 ();
 sg13g2_fill_2 FILLER_40_151 ();
 sg13g2_fill_2 FILLER_40_158 ();
 sg13g2_decap_8 FILLER_40_174 ();
 sg13g2_fill_1 FILLER_40_181 ();
 sg13g2_decap_4 FILLER_40_190 ();
 sg13g2_fill_2 FILLER_40_208 ();
 sg13g2_fill_2 FILLER_40_223 ();
 sg13g2_fill_1 FILLER_40_225 ();
 sg13g2_decap_4 FILLER_40_266 ();
 sg13g2_decap_4 FILLER_40_296 ();
 sg13g2_fill_1 FILLER_40_300 ();
 sg13g2_decap_4 FILLER_40_314 ();
 sg13g2_fill_2 FILLER_40_318 ();
 sg13g2_fill_2 FILLER_40_324 ();
 sg13g2_fill_1 FILLER_40_326 ();
 sg13g2_decap_4 FILLER_40_344 ();
 sg13g2_fill_1 FILLER_40_366 ();
 sg13g2_fill_2 FILLER_40_372 ();
 sg13g2_fill_1 FILLER_40_374 ();
 sg13g2_fill_2 FILLER_40_380 ();
 sg13g2_fill_1 FILLER_40_382 ();
 sg13g2_fill_2 FILLER_40_407 ();
 sg13g2_fill_1 FILLER_41_0 ();
 sg13g2_fill_1 FILLER_41_30 ();
 sg13g2_fill_2 FILLER_41_57 ();
 sg13g2_fill_1 FILLER_41_59 ();
 sg13g2_fill_2 FILLER_41_65 ();
 sg13g2_fill_1 FILLER_41_67 ();
 sg13g2_decap_4 FILLER_41_96 ();
 sg13g2_decap_8 FILLER_41_105 ();
 sg13g2_fill_2 FILLER_41_122 ();
 sg13g2_decap_8 FILLER_41_129 ();
 sg13g2_decap_4 FILLER_41_144 ();
 sg13g2_fill_2 FILLER_41_160 ();
 sg13g2_fill_2 FILLER_41_180 ();
 sg13g2_decap_4 FILLER_41_213 ();
 sg13g2_fill_2 FILLER_41_222 ();
 sg13g2_fill_1 FILLER_41_224 ();
 sg13g2_fill_1 FILLER_41_242 ();
 sg13g2_decap_4 FILLER_41_257 ();
 sg13g2_fill_2 FILLER_41_261 ();
 sg13g2_fill_2 FILLER_41_286 ();
 sg13g2_fill_2 FILLER_41_293 ();
 sg13g2_fill_1 FILLER_41_332 ();
 sg13g2_fill_2 FILLER_41_338 ();
 sg13g2_decap_8 FILLER_41_344 ();
 sg13g2_fill_2 FILLER_41_351 ();
 sg13g2_decap_4 FILLER_41_363 ();
 sg13g2_fill_2 FILLER_41_373 ();
 sg13g2_fill_2 FILLER_41_395 ();
 sg13g2_fill_1 FILLER_41_397 ();
 sg13g2_fill_2 FILLER_41_406 ();
 sg13g2_fill_1 FILLER_41_408 ();
 sg13g2_fill_1 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_13 ();
 sg13g2_fill_1 FILLER_42_20 ();
 sg13g2_fill_1 FILLER_42_26 ();
 sg13g2_fill_1 FILLER_42_35 ();
 sg13g2_decap_4 FILLER_42_41 ();
 sg13g2_fill_2 FILLER_42_45 ();
 sg13g2_decap_8 FILLER_42_78 ();
 sg13g2_fill_2 FILLER_42_85 ();
 sg13g2_fill_1 FILLER_42_87 ();
 sg13g2_fill_1 FILLER_42_111 ();
 sg13g2_fill_2 FILLER_42_119 ();
 sg13g2_fill_1 FILLER_42_121 ();
 sg13g2_decap_8 FILLER_42_134 ();
 sg13g2_fill_2 FILLER_42_141 ();
 sg13g2_fill_1 FILLER_42_143 ();
 sg13g2_decap_8 FILLER_42_149 ();
 sg13g2_decap_4 FILLER_42_202 ();
 sg13g2_fill_1 FILLER_42_206 ();
 sg13g2_fill_2 FILLER_42_236 ();
 sg13g2_fill_1 FILLER_42_251 ();
 sg13g2_fill_2 FILLER_42_275 ();
 sg13g2_fill_1 FILLER_42_277 ();
 sg13g2_fill_1 FILLER_42_288 ();
 sg13g2_fill_1 FILLER_42_304 ();
 sg13g2_decap_8 FILLER_42_309 ();
 sg13g2_decap_4 FILLER_42_373 ();
 sg13g2_fill_1 FILLER_42_377 ();
 sg13g2_fill_2 FILLER_42_395 ();
 sg13g2_fill_1 FILLER_42_397 ();
 sg13g2_decap_4 FILLER_43_0 ();
 sg13g2_fill_1 FILLER_43_4 ();
 sg13g2_decap_4 FILLER_43_24 ();
 sg13g2_fill_2 FILLER_43_28 ();
 sg13g2_decap_4 FILLER_43_42 ();
 sg13g2_decap_8 FILLER_43_53 ();
 sg13g2_fill_2 FILLER_43_60 ();
 sg13g2_decap_8 FILLER_43_66 ();
 sg13g2_fill_2 FILLER_43_94 ();
 sg13g2_fill_1 FILLER_43_114 ();
 sg13g2_fill_2 FILLER_43_140 ();
 sg13g2_fill_2 FILLER_43_174 ();
 sg13g2_fill_1 FILLER_43_176 ();
 sg13g2_fill_1 FILLER_43_214 ();
 sg13g2_decap_4 FILLER_43_221 ();
 sg13g2_fill_1 FILLER_43_225 ();
 sg13g2_decap_4 FILLER_43_231 ();
 sg13g2_decap_4 FILLER_43_247 ();
 sg13g2_fill_2 FILLER_43_251 ();
 sg13g2_decap_4 FILLER_43_259 ();
 sg13g2_decap_8 FILLER_43_275 ();
 sg13g2_decap_8 FILLER_43_282 ();
 sg13g2_fill_2 FILLER_43_289 ();
 sg13g2_fill_1 FILLER_43_291 ();
 sg13g2_fill_1 FILLER_43_301 ();
 sg13g2_fill_1 FILLER_43_311 ();
 sg13g2_decap_8 FILLER_43_325 ();
 sg13g2_fill_1 FILLER_43_332 ();
 sg13g2_decap_8 FILLER_43_338 ();
 sg13g2_fill_1 FILLER_43_361 ();
 sg13g2_decap_4 FILLER_43_365 ();
 sg13g2_fill_2 FILLER_43_369 ();
 sg13g2_decap_8 FILLER_43_381 ();
 sg13g2_fill_1 FILLER_43_388 ();
 sg13g2_fill_2 FILLER_43_393 ();
 sg13g2_fill_1 FILLER_43_400 ();
 sg13g2_decap_4 FILLER_44_0 ();
 sg13g2_fill_2 FILLER_44_4 ();
 sg13g2_fill_1 FILLER_44_19 ();
 sg13g2_decap_4 FILLER_44_38 ();
 sg13g2_fill_1 FILLER_44_42 ();
 sg13g2_fill_1 FILLER_44_56 ();
 sg13g2_fill_2 FILLER_44_81 ();
 sg13g2_fill_2 FILLER_44_92 ();
 sg13g2_fill_1 FILLER_44_94 ();
 sg13g2_decap_4 FILLER_44_101 ();
 sg13g2_fill_2 FILLER_44_105 ();
 sg13g2_decap_8 FILLER_44_119 ();
 sg13g2_decap_8 FILLER_44_126 ();
 sg13g2_decap_8 FILLER_44_133 ();
 sg13g2_decap_4 FILLER_44_140 ();
 sg13g2_fill_2 FILLER_44_150 ();
 sg13g2_fill_1 FILLER_44_152 ();
 sg13g2_fill_2 FILLER_44_163 ();
 sg13g2_decap_4 FILLER_44_174 ();
 sg13g2_decap_4 FILLER_44_184 ();
 sg13g2_decap_8 FILLER_44_196 ();
 sg13g2_fill_1 FILLER_44_203 ();
 sg13g2_fill_1 FILLER_44_208 ();
 sg13g2_fill_1 FILLER_44_214 ();
 sg13g2_fill_1 FILLER_44_220 ();
 sg13g2_fill_1 FILLER_44_229 ();
 sg13g2_decap_8 FILLER_44_243 ();
 sg13g2_fill_2 FILLER_44_250 ();
 sg13g2_decap_4 FILLER_44_256 ();
 sg13g2_fill_1 FILLER_44_260 ();
 sg13g2_fill_2 FILLER_44_267 ();
 sg13g2_fill_1 FILLER_44_273 ();
 sg13g2_fill_1 FILLER_44_323 ();
 sg13g2_decap_4 FILLER_44_343 ();
 sg13g2_fill_2 FILLER_44_398 ();
 sg13g2_fill_1 FILLER_44_408 ();
 sg13g2_fill_1 FILLER_45_0 ();
 sg13g2_fill_2 FILLER_45_17 ();
 sg13g2_fill_1 FILLER_45_19 ();
 sg13g2_fill_1 FILLER_45_42 ();
 sg13g2_decap_4 FILLER_45_47 ();
 sg13g2_fill_1 FILLER_45_51 ();
 sg13g2_decap_4 FILLER_45_57 ();
 sg13g2_decap_4 FILLER_45_66 ();
 sg13g2_fill_1 FILLER_45_70 ();
 sg13g2_fill_2 FILLER_45_77 ();
 sg13g2_fill_2 FILLER_45_102 ();
 sg13g2_fill_1 FILLER_45_104 ();
 sg13g2_fill_1 FILLER_45_153 ();
 sg13g2_decap_4 FILLER_45_178 ();
 sg13g2_fill_1 FILLER_45_182 ();
 sg13g2_fill_2 FILLER_45_188 ();
 sg13g2_fill_1 FILLER_45_190 ();
 sg13g2_fill_1 FILLER_45_196 ();
 sg13g2_decap_8 FILLER_45_216 ();
 sg13g2_decap_4 FILLER_45_231 ();
 sg13g2_fill_2 FILLER_45_235 ();
 sg13g2_fill_2 FILLER_45_298 ();
 sg13g2_fill_1 FILLER_45_300 ();
 sg13g2_fill_1 FILLER_45_307 ();
 sg13g2_fill_2 FILLER_45_312 ();
 sg13g2_decap_8 FILLER_45_320 ();
 sg13g2_decap_4 FILLER_45_327 ();
 sg13g2_fill_2 FILLER_45_352 ();
 sg13g2_fill_1 FILLER_45_354 ();
 sg13g2_fill_1 FILLER_45_358 ();
 sg13g2_fill_2 FILLER_45_368 ();
 sg13g2_fill_1 FILLER_45_370 ();
 sg13g2_fill_1 FILLER_45_381 ();
 sg13g2_fill_1 FILLER_45_391 ();
 sg13g2_fill_1 FILLER_45_395 ();
 sg13g2_fill_1 FILLER_46_0 ();
 sg13g2_fill_2 FILLER_46_14 ();
 sg13g2_fill_2 FILLER_46_32 ();
 sg13g2_fill_2 FILLER_46_38 ();
 sg13g2_fill_2 FILLER_46_49 ();
 sg13g2_fill_2 FILLER_46_58 ();
 sg13g2_fill_1 FILLER_46_60 ();
 sg13g2_fill_2 FILLER_46_72 ();
 sg13g2_fill_1 FILLER_46_74 ();
 sg13g2_fill_1 FILLER_46_80 ();
 sg13g2_decap_4 FILLER_46_91 ();
 sg13g2_fill_1 FILLER_46_95 ();
 sg13g2_decap_8 FILLER_46_106 ();
 sg13g2_decap_4 FILLER_46_113 ();
 sg13g2_decap_8 FILLER_46_129 ();
 sg13g2_fill_1 FILLER_46_136 ();
 sg13g2_fill_1 FILLER_46_140 ();
 sg13g2_fill_1 FILLER_46_150 ();
 sg13g2_fill_2 FILLER_46_179 ();
 sg13g2_fill_2 FILLER_46_200 ();
 sg13g2_fill_1 FILLER_46_224 ();
 sg13g2_fill_1 FILLER_46_234 ();
 sg13g2_fill_2 FILLER_46_245 ();
 sg13g2_fill_1 FILLER_46_247 ();
 sg13g2_fill_2 FILLER_46_256 ();
 sg13g2_fill_1 FILLER_46_258 ();
 sg13g2_decap_4 FILLER_46_281 ();
 sg13g2_decap_4 FILLER_46_316 ();
 sg13g2_fill_1 FILLER_46_320 ();
 sg13g2_decap_4 FILLER_46_329 ();
 sg13g2_decap_8 FILLER_46_362 ();
 sg13g2_fill_2 FILLER_46_387 ();
 sg13g2_fill_1 FILLER_46_389 ();
 sg13g2_fill_2 FILLER_46_398 ();
 sg13g2_fill_1 FILLER_46_400 ();
 sg13g2_fill_2 FILLER_46_406 ();
 sg13g2_fill_1 FILLER_46_408 ();
 sg13g2_decap_4 FILLER_47_0 ();
 sg13g2_fill_2 FILLER_47_25 ();
 sg13g2_fill_1 FILLER_47_27 ();
 sg13g2_fill_1 FILLER_47_41 ();
 sg13g2_fill_2 FILLER_47_50 ();
 sg13g2_fill_1 FILLER_47_52 ();
 sg13g2_fill_2 FILLER_47_58 ();
 sg13g2_fill_1 FILLER_47_60 ();
 sg13g2_fill_2 FILLER_47_65 ();
 sg13g2_decap_8 FILLER_47_81 ();
 sg13g2_decap_4 FILLER_47_88 ();
 sg13g2_fill_1 FILLER_47_92 ();
 sg13g2_fill_2 FILLER_47_102 ();
 sg13g2_decap_4 FILLER_47_126 ();
 sg13g2_fill_1 FILLER_47_130 ();
 sg13g2_fill_1 FILLER_47_144 ();
 sg13g2_decap_8 FILLER_47_154 ();
 sg13g2_decap_8 FILLER_47_161 ();
 sg13g2_decap_8 FILLER_47_168 ();
 sg13g2_decap_4 FILLER_47_175 ();
 sg13g2_decap_8 FILLER_47_184 ();
 sg13g2_fill_2 FILLER_47_199 ();
 sg13g2_decap_4 FILLER_47_223 ();
 sg13g2_fill_2 FILLER_47_227 ();
 sg13g2_decap_4 FILLER_47_237 ();
 sg13g2_decap_4 FILLER_47_246 ();
 sg13g2_fill_2 FILLER_47_261 ();
 sg13g2_fill_2 FILLER_47_277 ();
 sg13g2_fill_1 FILLER_47_279 ();
 sg13g2_fill_2 FILLER_47_293 ();
 sg13g2_fill_2 FILLER_47_321 ();
 sg13g2_decap_4 FILLER_47_331 ();
 sg13g2_fill_1 FILLER_47_343 ();
 sg13g2_fill_2 FILLER_47_376 ();
 sg13g2_fill_1 FILLER_47_378 ();
 sg13g2_fill_1 FILLER_47_387 ();
 sg13g2_fill_1 FILLER_47_408 ();
 sg13g2_decap_4 FILLER_48_0 ();
 sg13g2_fill_1 FILLER_48_4 ();
 sg13g2_fill_2 FILLER_48_10 ();
 sg13g2_fill_1 FILLER_48_12 ();
 sg13g2_decap_4 FILLER_48_17 ();
 sg13g2_fill_1 FILLER_48_21 ();
 sg13g2_decap_4 FILLER_48_30 ();
 sg13g2_fill_1 FILLER_48_34 ();
 sg13g2_fill_2 FILLER_48_65 ();
 sg13g2_fill_2 FILLER_48_109 ();
 sg13g2_fill_1 FILLER_48_119 ();
 sg13g2_fill_2 FILLER_48_125 ();
 sg13g2_fill_1 FILLER_48_153 ();
 sg13g2_decap_8 FILLER_48_162 ();
 sg13g2_fill_1 FILLER_48_177 ();
 sg13g2_decap_8 FILLER_48_188 ();
 sg13g2_decap_4 FILLER_48_199 ();
 sg13g2_decap_8 FILLER_48_211 ();
 sg13g2_fill_2 FILLER_48_218 ();
 sg13g2_fill_1 FILLER_48_220 ();
 sg13g2_fill_2 FILLER_48_239 ();
 sg13g2_fill_2 FILLER_48_249 ();
 sg13g2_fill_1 FILLER_48_251 ();
 sg13g2_fill_2 FILLER_48_286 ();
 sg13g2_fill_1 FILLER_48_288 ();
 sg13g2_fill_1 FILLER_48_297 ();
 sg13g2_fill_2 FILLER_48_302 ();
 sg13g2_fill_1 FILLER_48_304 ();
 sg13g2_fill_2 FILLER_48_309 ();
 sg13g2_fill_1 FILLER_48_316 ();
 sg13g2_fill_2 FILLER_48_321 ();
 sg13g2_decap_4 FILLER_48_332 ();
 sg13g2_decap_8 FILLER_48_341 ();
 sg13g2_decap_4 FILLER_48_348 ();
 sg13g2_fill_2 FILLER_48_352 ();
 sg13g2_decap_8 FILLER_48_377 ();
 sg13g2_decap_8 FILLER_48_388 ();
 sg13g2_decap_4 FILLER_48_403 ();
 sg13g2_fill_2 FILLER_48_407 ();
 sg13g2_decap_4 FILLER_49_0 ();
 sg13g2_decap_4 FILLER_49_12 ();
 sg13g2_fill_1 FILLER_49_16 ();
 sg13g2_fill_1 FILLER_49_25 ();
 sg13g2_fill_1 FILLER_49_34 ();
 sg13g2_decap_8 FILLER_49_40 ();
 sg13g2_decap_8 FILLER_49_47 ();
 sg13g2_decap_8 FILLER_49_54 ();
 sg13g2_decap_8 FILLER_49_78 ();
 sg13g2_fill_2 FILLER_49_85 ();
 sg13g2_fill_1 FILLER_49_93 ();
 sg13g2_decap_4 FILLER_49_103 ();
 sg13g2_decap_8 FILLER_49_112 ();
 sg13g2_fill_2 FILLER_49_124 ();
 sg13g2_fill_1 FILLER_49_139 ();
 sg13g2_fill_2 FILLER_49_148 ();
 sg13g2_fill_1 FILLER_49_150 ();
 sg13g2_fill_2 FILLER_49_181 ();
 sg13g2_fill_1 FILLER_49_183 ();
 sg13g2_fill_2 FILLER_49_248 ();
 sg13g2_fill_2 FILLER_49_259 ();
 sg13g2_fill_1 FILLER_49_261 ();
 sg13g2_fill_2 FILLER_49_266 ();
 sg13g2_decap_4 FILLER_49_273 ();
 sg13g2_fill_2 FILLER_49_277 ();
 sg13g2_fill_2 FILLER_49_300 ();
 sg13g2_fill_1 FILLER_49_310 ();
 sg13g2_decap_8 FILLER_49_316 ();
 sg13g2_fill_2 FILLER_49_334 ();
 sg13g2_decap_4 FILLER_49_344 ();
 sg13g2_fill_1 FILLER_49_360 ();
 sg13g2_fill_1 FILLER_49_365 ();
 sg13g2_decap_8 FILLER_49_370 ();
 sg13g2_fill_2 FILLER_49_377 ();
 sg13g2_fill_1 FILLER_49_379 ();
 sg13g2_decap_4 FILLER_49_404 ();
 sg13g2_fill_1 FILLER_49_408 ();
 sg13g2_fill_1 FILLER_50_0 ();
 sg13g2_fill_1 FILLER_50_22 ();
 sg13g2_fill_2 FILLER_50_27 ();
 sg13g2_fill_1 FILLER_50_33 ();
 sg13g2_decap_8 FILLER_50_50 ();
 sg13g2_decap_8 FILLER_50_57 ();
 sg13g2_decap_4 FILLER_50_64 ();
 sg13g2_fill_2 FILLER_50_68 ();
 sg13g2_fill_2 FILLER_50_80 ();
 sg13g2_decap_4 FILLER_50_102 ();
 sg13g2_fill_2 FILLER_50_112 ();
 sg13g2_fill_1 FILLER_50_114 ();
 sg13g2_decap_4 FILLER_50_129 ();
 sg13g2_fill_2 FILLER_50_147 ();
 sg13g2_fill_1 FILLER_50_158 ();
 sg13g2_fill_2 FILLER_50_194 ();
 sg13g2_fill_1 FILLER_50_196 ();
 sg13g2_fill_2 FILLER_50_210 ();
 sg13g2_decap_4 FILLER_50_217 ();
 sg13g2_fill_2 FILLER_50_221 ();
 sg13g2_fill_2 FILLER_50_278 ();
 sg13g2_decap_4 FILLER_50_298 ();
 sg13g2_fill_2 FILLER_50_312 ();
 sg13g2_fill_1 FILLER_50_334 ();
 sg13g2_decap_8 FILLER_50_342 ();
 sg13g2_decap_4 FILLER_50_349 ();
 sg13g2_decap_4 FILLER_50_382 ();
 sg13g2_fill_1 FILLER_50_399 ();
 sg13g2_fill_1 FILLER_50_408 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_decap_8 FILLER_51_7 ();
 sg13g2_decap_4 FILLER_51_14 ();
 sg13g2_fill_2 FILLER_51_21 ();
 sg13g2_fill_1 FILLER_51_33 ();
 sg13g2_fill_1 FILLER_51_61 ();
 sg13g2_fill_2 FILLER_51_66 ();
 sg13g2_fill_1 FILLER_51_68 ();
 sg13g2_fill_1 FILLER_51_83 ();
 sg13g2_decap_4 FILLER_51_89 ();
 sg13g2_fill_2 FILLER_51_93 ();
 sg13g2_fill_2 FILLER_51_103 ();
 sg13g2_decap_4 FILLER_51_115 ();
 sg13g2_decap_8 FILLER_51_124 ();
 sg13g2_fill_2 FILLER_51_136 ();
 sg13g2_fill_1 FILLER_51_138 ();
 sg13g2_fill_1 FILLER_51_253 ();
 sg13g2_fill_2 FILLER_51_260 ();
 sg13g2_decap_8 FILLER_51_271 ();
 sg13g2_fill_2 FILLER_51_288 ();
 sg13g2_fill_1 FILLER_51_290 ();
 sg13g2_decap_4 FILLER_51_298 ();
 sg13g2_fill_2 FILLER_51_302 ();
 sg13g2_fill_2 FILLER_51_312 ();
 sg13g2_fill_1 FILLER_51_314 ();
 sg13g2_fill_2 FILLER_51_322 ();
 sg13g2_fill_1 FILLER_51_324 ();
 sg13g2_fill_1 FILLER_51_333 ();
 sg13g2_fill_2 FILLER_51_342 ();
 sg13g2_fill_1 FILLER_51_344 ();
 sg13g2_fill_1 FILLER_51_357 ();
 sg13g2_fill_2 FILLER_51_363 ();
 sg13g2_fill_1 FILLER_51_365 ();
 sg13g2_decap_4 FILLER_51_395 ();
 sg13g2_fill_1 FILLER_51_399 ();
 sg13g2_fill_2 FILLER_51_407 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_decap_4 FILLER_52_7 ();
 sg13g2_fill_2 FILLER_52_11 ();
 sg13g2_decap_4 FILLER_52_17 ();
 sg13g2_fill_2 FILLER_52_25 ();
 sg13g2_fill_2 FILLER_52_45 ();
 sg13g2_fill_1 FILLER_52_47 ();
 sg13g2_fill_2 FILLER_52_63 ();
 sg13g2_fill_1 FILLER_52_65 ();
 sg13g2_decap_4 FILLER_52_75 ();
 sg13g2_fill_1 FILLER_52_79 ();
 sg13g2_fill_2 FILLER_52_88 ();
 sg13g2_fill_1 FILLER_52_90 ();
 sg13g2_fill_1 FILLER_52_103 ();
 sg13g2_decap_8 FILLER_52_112 ();
 sg13g2_fill_1 FILLER_52_127 ();
 sg13g2_decap_8 FILLER_52_142 ();
 sg13g2_fill_2 FILLER_52_165 ();
 sg13g2_decap_4 FILLER_52_207 ();
 sg13g2_fill_1 FILLER_52_216 ();
 sg13g2_decap_4 FILLER_52_230 ();
 sg13g2_fill_2 FILLER_52_234 ();
 sg13g2_fill_1 FILLER_52_252 ();
 sg13g2_decap_4 FILLER_52_273 ();
 sg13g2_fill_2 FILLER_52_277 ();
 sg13g2_fill_2 FILLER_52_284 ();
 sg13g2_fill_2 FILLER_52_296 ();
 sg13g2_fill_2 FILLER_52_329 ();
 sg13g2_fill_1 FILLER_52_331 ();
 sg13g2_fill_1 FILLER_52_340 ();
 sg13g2_fill_1 FILLER_52_355 ();
 sg13g2_fill_2 FILLER_52_365 ();
 sg13g2_fill_2 FILLER_52_372 ();
 sg13g2_fill_1 FILLER_52_374 ();
 sg13g2_decap_8 FILLER_52_383 ();
 sg13g2_fill_1 FILLER_52_390 ();
 sg13g2_fill_2 FILLER_52_407 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_decap_4 FILLER_53_7 ();
 sg13g2_decap_4 FILLER_53_23 ();
 sg13g2_fill_1 FILLER_53_27 ();
 sg13g2_fill_1 FILLER_53_53 ();
 sg13g2_fill_2 FILLER_53_92 ();
 sg13g2_fill_1 FILLER_53_94 ();
 sg13g2_decap_4 FILLER_53_99 ();
 sg13g2_fill_2 FILLER_53_103 ();
 sg13g2_fill_1 FILLER_53_129 ();
 sg13g2_fill_1 FILLER_53_134 ();
 sg13g2_fill_2 FILLER_53_151 ();
 sg13g2_fill_2 FILLER_53_179 ();
 sg13g2_fill_2 FILLER_53_189 ();
 sg13g2_fill_1 FILLER_53_191 ();
 sg13g2_decap_8 FILLER_53_196 ();
 sg13g2_decap_4 FILLER_53_203 ();
 sg13g2_fill_2 FILLER_53_207 ();
 sg13g2_fill_2 FILLER_53_221 ();
 sg13g2_fill_1 FILLER_53_223 ();
 sg13g2_decap_8 FILLER_53_242 ();
 sg13g2_decap_4 FILLER_53_249 ();
 sg13g2_fill_1 FILLER_53_253 ();
 sg13g2_decap_4 FILLER_53_294 ();
 sg13g2_fill_2 FILLER_53_298 ();
 sg13g2_fill_2 FILLER_53_305 ();
 sg13g2_fill_1 FILLER_53_307 ();
 sg13g2_decap_8 FILLER_53_312 ();
 sg13g2_fill_2 FILLER_53_319 ();
 sg13g2_fill_1 FILLER_53_321 ();
 sg13g2_fill_2 FILLER_53_350 ();
 sg13g2_fill_1 FILLER_53_352 ();
 sg13g2_fill_1 FILLER_53_391 ();
 sg13g2_fill_1 FILLER_53_396 ();
 sg13g2_fill_2 FILLER_53_406 ();
 sg13g2_fill_1 FILLER_53_408 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_fill_1 FILLER_54_7 ();
 sg13g2_fill_2 FILLER_54_28 ();
 sg13g2_decap_8 FILLER_54_34 ();
 sg13g2_decap_4 FILLER_54_41 ();
 sg13g2_fill_1 FILLER_54_45 ();
 sg13g2_decap_8 FILLER_54_66 ();
 sg13g2_decap_8 FILLER_54_73 ();
 sg13g2_decap_8 FILLER_54_80 ();
 sg13g2_fill_1 FILLER_54_99 ();
 sg13g2_fill_1 FILLER_54_116 ();
 sg13g2_fill_2 FILLER_54_125 ();
 sg13g2_decap_8 FILLER_54_148 ();
 sg13g2_decap_8 FILLER_54_155 ();
 sg13g2_fill_2 FILLER_54_162 ();
 sg13g2_fill_1 FILLER_54_164 ();
 sg13g2_decap_4 FILLER_54_182 ();
 sg13g2_fill_2 FILLER_54_198 ();
 sg13g2_fill_1 FILLER_54_212 ();
 sg13g2_decap_4 FILLER_54_226 ();
 sg13g2_fill_2 FILLER_54_230 ();
 sg13g2_decap_4 FILLER_54_240 ();
 sg13g2_fill_1 FILLER_54_250 ();
 sg13g2_fill_2 FILLER_54_278 ();
 sg13g2_fill_1 FILLER_54_285 ();
 sg13g2_decap_4 FILLER_54_309 ();
 sg13g2_decap_4 FILLER_54_330 ();
 sg13g2_fill_2 FILLER_54_334 ();
 sg13g2_fill_2 FILLER_54_342 ();
 sg13g2_fill_1 FILLER_54_349 ();
 sg13g2_fill_2 FILLER_54_364 ();
 sg13g2_decap_8 FILLER_54_370 ();
 sg13g2_decap_4 FILLER_54_377 ();
 sg13g2_fill_1 FILLER_54_381 ();
 sg13g2_fill_2 FILLER_54_397 ();
 sg13g2_fill_2 FILLER_54_407 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_decap_8 FILLER_55_7 ();
 sg13g2_decap_8 FILLER_55_14 ();
 sg13g2_fill_2 FILLER_55_46 ();
 sg13g2_fill_1 FILLER_55_48 ();
 sg13g2_decap_4 FILLER_55_58 ();
 sg13g2_decap_4 FILLER_55_77 ();
 sg13g2_decap_8 FILLER_55_93 ();
 sg13g2_fill_1 FILLER_55_100 ();
 sg13g2_decap_4 FILLER_55_111 ();
 sg13g2_decap_4 FILLER_55_126 ();
 sg13g2_fill_1 FILLER_55_130 ();
 sg13g2_decap_4 FILLER_55_141 ();
 sg13g2_fill_1 FILLER_55_145 ();
 sg13g2_decap_4 FILLER_55_165 ();
 sg13g2_fill_2 FILLER_55_191 ();
 sg13g2_decap_4 FILLER_55_198 ();
 sg13g2_fill_2 FILLER_55_202 ();
 sg13g2_decap_8 FILLER_55_217 ();
 sg13g2_decap_8 FILLER_55_224 ();
 sg13g2_decap_8 FILLER_55_236 ();
 sg13g2_fill_1 FILLER_55_243 ();
 sg13g2_decap_8 FILLER_55_249 ();
 sg13g2_fill_1 FILLER_55_256 ();
 sg13g2_fill_2 FILLER_55_263 ();
 sg13g2_fill_1 FILLER_55_265 ();
 sg13g2_decap_8 FILLER_55_270 ();
 sg13g2_decap_8 FILLER_55_291 ();
 sg13g2_decap_4 FILLER_55_298 ();
 sg13g2_fill_2 FILLER_55_307 ();
 sg13g2_fill_1 FILLER_55_318 ();
 sg13g2_fill_2 FILLER_55_327 ();
 sg13g2_fill_1 FILLER_55_329 ();
 sg13g2_fill_2 FILLER_55_350 ();
 sg13g2_fill_2 FILLER_55_368 ();
 sg13g2_fill_1 FILLER_55_380 ();
 sg13g2_decap_8 FILLER_55_386 ();
 sg13g2_fill_1 FILLER_55_399 ();
 sg13g2_fill_1 FILLER_55_408 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_decap_8 FILLER_56_7 ();
 sg13g2_decap_8 FILLER_56_14 ();
 sg13g2_decap_8 FILLER_56_21 ();
 sg13g2_decap_8 FILLER_56_28 ();
 sg13g2_decap_8 FILLER_56_35 ();
 sg13g2_fill_2 FILLER_56_84 ();
 sg13g2_fill_1 FILLER_56_86 ();
 sg13g2_decap_4 FILLER_56_99 ();
 sg13g2_fill_2 FILLER_56_115 ();
 sg13g2_fill_1 FILLER_56_117 ();
 sg13g2_decap_4 FILLER_56_137 ();
 sg13g2_fill_2 FILLER_56_157 ();
 sg13g2_fill_1 FILLER_56_159 ();
 sg13g2_fill_2 FILLER_56_225 ();
 sg13g2_fill_1 FILLER_56_227 ();
 sg13g2_fill_1 FILLER_56_236 ();
 sg13g2_fill_2 FILLER_56_263 ();
 sg13g2_fill_1 FILLER_56_265 ();
 sg13g2_fill_1 FILLER_56_281 ();
 sg13g2_fill_2 FILLER_56_288 ();
 sg13g2_fill_2 FILLER_56_304 ();
 sg13g2_fill_1 FILLER_56_306 ();
 sg13g2_decap_4 FILLER_56_317 ();
 sg13g2_fill_2 FILLER_56_329 ();
 sg13g2_decap_8 FILLER_56_339 ();
 sg13g2_decap_8 FILLER_56_346 ();
 sg13g2_decap_4 FILLER_56_353 ();
 sg13g2_fill_1 FILLER_56_362 ();
 sg13g2_fill_1 FILLER_56_382 ();
 sg13g2_fill_1 FILLER_56_399 ();
 sg13g2_fill_2 FILLER_56_407 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_decap_8 FILLER_57_7 ();
 sg13g2_decap_8 FILLER_57_14 ();
 sg13g2_decap_8 FILLER_57_21 ();
 sg13g2_decap_8 FILLER_57_28 ();
 sg13g2_decap_8 FILLER_57_35 ();
 sg13g2_decap_8 FILLER_57_42 ();
 sg13g2_fill_2 FILLER_57_49 ();
 sg13g2_fill_1 FILLER_57_51 ();
 sg13g2_fill_2 FILLER_57_65 ();
 sg13g2_decap_8 FILLER_57_71 ();
 sg13g2_decap_4 FILLER_57_78 ();
 sg13g2_fill_1 FILLER_57_82 ();
 sg13g2_fill_2 FILLER_57_105 ();
 sg13g2_fill_1 FILLER_57_107 ();
 sg13g2_fill_1 FILLER_57_118 ();
 sg13g2_decap_8 FILLER_57_124 ();
 sg13g2_fill_2 FILLER_57_131 ();
 sg13g2_fill_1 FILLER_57_133 ();
 sg13g2_decap_8 FILLER_57_140 ();
 sg13g2_decap_4 FILLER_57_155 ();
 sg13g2_fill_1 FILLER_57_159 ();
 sg13g2_decap_8 FILLER_57_170 ();
 sg13g2_fill_2 FILLER_57_177 ();
 sg13g2_decap_4 FILLER_57_192 ();
 sg13g2_fill_1 FILLER_57_196 ();
 sg13g2_decap_8 FILLER_57_207 ();
 sg13g2_fill_1 FILLER_57_214 ();
 sg13g2_fill_2 FILLER_57_220 ();
 sg13g2_fill_1 FILLER_57_222 ();
 sg13g2_fill_2 FILLER_57_241 ();
 sg13g2_fill_1 FILLER_57_243 ();
 sg13g2_fill_2 FILLER_57_253 ();
 sg13g2_fill_1 FILLER_57_255 ();
 sg13g2_decap_8 FILLER_57_265 ();
 sg13g2_decap_8 FILLER_57_272 ();
 sg13g2_fill_2 FILLER_57_289 ();
 sg13g2_fill_1 FILLER_57_300 ();
 sg13g2_fill_1 FILLER_57_330 ();
 sg13g2_fill_2 FILLER_57_339 ();
 sg13g2_fill_1 FILLER_57_341 ();
 sg13g2_decap_8 FILLER_57_356 ();
 sg13g2_decap_4 FILLER_57_363 ();
 sg13g2_fill_1 FILLER_57_367 ();
 sg13g2_fill_1 FILLER_57_372 ();
 sg13g2_decap_8 FILLER_57_380 ();
 sg13g2_decap_4 FILLER_57_387 ();
 sg13g2_fill_1 FILLER_57_408 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_decap_8 FILLER_58_7 ();
 sg13g2_decap_8 FILLER_58_14 ();
 sg13g2_decap_8 FILLER_58_21 ();
 sg13g2_decap_8 FILLER_58_28 ();
 sg13g2_decap_8 FILLER_58_35 ();
 sg13g2_decap_8 FILLER_58_42 ();
 sg13g2_decap_8 FILLER_58_49 ();
 sg13g2_decap_4 FILLER_58_56 ();
 sg13g2_fill_1 FILLER_58_70 ();
 sg13g2_decap_4 FILLER_58_98 ();
 sg13g2_fill_1 FILLER_58_102 ();
 sg13g2_decap_4 FILLER_58_110 ();
 sg13g2_decap_8 FILLER_58_119 ();
 sg13g2_fill_1 FILLER_58_126 ();
 sg13g2_fill_1 FILLER_58_149 ();
 sg13g2_decap_4 FILLER_58_158 ();
 sg13g2_fill_2 FILLER_58_169 ();
 sg13g2_fill_2 FILLER_58_179 ();
 sg13g2_fill_1 FILLER_58_181 ();
 sg13g2_fill_2 FILLER_58_195 ();
 sg13g2_fill_2 FILLER_58_227 ();
 sg13g2_fill_1 FILLER_58_229 ();
 sg13g2_fill_2 FILLER_58_238 ();
 sg13g2_fill_1 FILLER_58_240 ();
 sg13g2_fill_2 FILLER_58_249 ();
 sg13g2_fill_1 FILLER_58_251 ();
 sg13g2_fill_2 FILLER_58_261 ();
 sg13g2_fill_1 FILLER_58_268 ();
 sg13g2_fill_1 FILLER_58_274 ();
 sg13g2_fill_2 FILLER_58_289 ();
 sg13g2_fill_2 FILLER_58_318 ();
 sg13g2_fill_1 FILLER_58_320 ();
 sg13g2_fill_2 FILLER_58_335 ();
 sg13g2_fill_1 FILLER_58_337 ();
 sg13g2_fill_2 FILLER_58_352 ();
 sg13g2_fill_1 FILLER_58_354 ();
 sg13g2_fill_1 FILLER_58_408 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_decap_8 FILLER_59_7 ();
 sg13g2_decap_8 FILLER_59_14 ();
 sg13g2_decap_8 FILLER_59_21 ();
 sg13g2_decap_8 FILLER_59_28 ();
 sg13g2_decap_8 FILLER_59_35 ();
 sg13g2_decap_8 FILLER_59_42 ();
 sg13g2_fill_1 FILLER_59_49 ();
 sg13g2_fill_1 FILLER_59_66 ();
 sg13g2_fill_2 FILLER_59_80 ();
 sg13g2_fill_1 FILLER_59_82 ();
 sg13g2_decap_4 FILLER_59_91 ();
 sg13g2_fill_1 FILLER_59_109 ();
 sg13g2_fill_2 FILLER_59_122 ();
 sg13g2_fill_2 FILLER_59_140 ();
 sg13g2_fill_1 FILLER_59_142 ();
 sg13g2_fill_1 FILLER_59_158 ();
 sg13g2_fill_2 FILLER_59_167 ();
 sg13g2_decap_4 FILLER_59_186 ();
 sg13g2_fill_2 FILLER_59_206 ();
 sg13g2_fill_1 FILLER_59_208 ();
 sg13g2_decap_4 FILLER_59_217 ();
 sg13g2_fill_2 FILLER_59_234 ();
 sg13g2_fill_2 FILLER_59_244 ();
 sg13g2_fill_1 FILLER_59_246 ();
 sg13g2_decap_8 FILLER_59_280 ();
 sg13g2_fill_1 FILLER_59_287 ();
 sg13g2_decap_4 FILLER_59_318 ();
 sg13g2_fill_1 FILLER_59_338 ();
 sg13g2_fill_2 FILLER_59_364 ();
 sg13g2_decap_8 FILLER_59_379 ();
 sg13g2_fill_2 FILLER_59_386 ();
 sg13g2_fill_1 FILLER_59_392 ();
 sg13g2_fill_2 FILLER_59_406 ();
 sg13g2_fill_1 FILLER_59_408 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_decap_8 FILLER_60_7 ();
 sg13g2_decap_8 FILLER_60_14 ();
 sg13g2_decap_8 FILLER_60_21 ();
 sg13g2_decap_8 FILLER_60_28 ();
 sg13g2_decap_4 FILLER_60_35 ();
 sg13g2_fill_2 FILLER_60_39 ();
 sg13g2_fill_2 FILLER_60_49 ();
 sg13g2_fill_1 FILLER_60_51 ();
 sg13g2_fill_1 FILLER_60_57 ();
 sg13g2_decap_8 FILLER_60_113 ();
 sg13g2_decap_4 FILLER_60_120 ();
 sg13g2_fill_2 FILLER_60_133 ();
 sg13g2_fill_1 FILLER_60_135 ();
 sg13g2_fill_2 FILLER_60_141 ();
 sg13g2_decap_8 FILLER_60_147 ();
 sg13g2_fill_2 FILLER_60_169 ();
 sg13g2_decap_8 FILLER_60_176 ();
 sg13g2_fill_1 FILLER_60_183 ();
 sg13g2_decap_8 FILLER_60_188 ();
 sg13g2_fill_2 FILLER_60_206 ();
 sg13g2_decap_8 FILLER_60_211 ();
 sg13g2_decap_4 FILLER_60_231 ();
 sg13g2_decap_8 FILLER_60_243 ();
 sg13g2_decap_8 FILLER_60_250 ();
 sg13g2_decap_8 FILLER_60_257 ();
 sg13g2_fill_1 FILLER_60_264 ();
 sg13g2_fill_2 FILLER_60_275 ();
 sg13g2_fill_1 FILLER_60_277 ();
 sg13g2_decap_8 FILLER_60_286 ();
 sg13g2_decap_4 FILLER_60_293 ();
 sg13g2_fill_2 FILLER_60_309 ();
 sg13g2_fill_1 FILLER_60_311 ();
 sg13g2_decap_4 FILLER_60_339 ();
 sg13g2_decap_4 FILLER_60_347 ();
 sg13g2_fill_2 FILLER_60_351 ();
 sg13g2_decap_4 FILLER_60_379 ();
 sg13g2_fill_1 FILLER_60_408 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_decap_8 FILLER_61_7 ();
 sg13g2_decap_8 FILLER_61_14 ();
 sg13g2_decap_8 FILLER_61_21 ();
 sg13g2_decap_8 FILLER_61_28 ();
 sg13g2_fill_2 FILLER_61_35 ();
 sg13g2_decap_4 FILLER_61_53 ();
 sg13g2_decap_8 FILLER_61_63 ();
 sg13g2_decap_8 FILLER_61_74 ();
 sg13g2_decap_8 FILLER_61_81 ();
 sg13g2_fill_1 FILLER_61_88 ();
 sg13g2_fill_2 FILLER_61_94 ();
 sg13g2_fill_1 FILLER_61_96 ();
 sg13g2_decap_4 FILLER_61_103 ();
 sg13g2_fill_1 FILLER_61_107 ();
 sg13g2_fill_1 FILLER_61_126 ();
 sg13g2_fill_2 FILLER_61_135 ();
 sg13g2_fill_1 FILLER_61_137 ();
 sg13g2_decap_4 FILLER_61_154 ();
 sg13g2_fill_2 FILLER_61_195 ();
 sg13g2_fill_2 FILLER_61_201 ();
 sg13g2_fill_1 FILLER_61_203 ();
 sg13g2_fill_2 FILLER_61_220 ();
 sg13g2_fill_2 FILLER_61_239 ();
 sg13g2_fill_1 FILLER_61_267 ();
 sg13g2_decap_4 FILLER_61_277 ();
 sg13g2_fill_1 FILLER_61_281 ();
 sg13g2_fill_2 FILLER_61_298 ();
 sg13g2_fill_1 FILLER_61_300 ();
 sg13g2_fill_1 FILLER_61_321 ();
 sg13g2_decap_4 FILLER_61_326 ();
 sg13g2_fill_1 FILLER_61_330 ();
 sg13g2_decap_8 FILLER_61_336 ();
 sg13g2_fill_2 FILLER_61_343 ();
 sg13g2_decap_4 FILLER_61_350 ();
 sg13g2_decap_4 FILLER_61_366 ();
 sg13g2_fill_1 FILLER_61_379 ();
 sg13g2_decap_8 FILLER_61_391 ();
 sg13g2_fill_2 FILLER_61_398 ();
 sg13g2_decap_4 FILLER_61_405 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_decap_8 FILLER_62_7 ();
 sg13g2_decap_8 FILLER_62_14 ();
 sg13g2_decap_8 FILLER_62_21 ();
 sg13g2_decap_8 FILLER_62_28 ();
 sg13g2_fill_1 FILLER_62_35 ();
 sg13g2_decap_8 FILLER_62_41 ();
 sg13g2_fill_2 FILLER_62_48 ();
 sg13g2_decap_4 FILLER_62_56 ();
 sg13g2_fill_1 FILLER_62_60 ();
 sg13g2_fill_2 FILLER_62_65 ();
 sg13g2_fill_1 FILLER_62_67 ();
 sg13g2_fill_2 FILLER_62_74 ();
 sg13g2_fill_1 FILLER_62_76 ();
 sg13g2_fill_2 FILLER_62_87 ();
 sg13g2_fill_1 FILLER_62_89 ();
 sg13g2_decap_4 FILLER_62_99 ();
 sg13g2_fill_1 FILLER_62_103 ();
 sg13g2_fill_2 FILLER_62_117 ();
 sg13g2_fill_2 FILLER_62_123 ();
 sg13g2_decap_4 FILLER_62_128 ();
 sg13g2_decap_8 FILLER_62_138 ();
 sg13g2_fill_2 FILLER_62_145 ();
 sg13g2_fill_1 FILLER_62_147 ();
 sg13g2_decap_4 FILLER_62_168 ();
 sg13g2_fill_1 FILLER_62_172 ();
 sg13g2_fill_2 FILLER_62_184 ();
 sg13g2_fill_1 FILLER_62_186 ();
 sg13g2_decap_4 FILLER_62_191 ();
 sg13g2_decap_4 FILLER_62_203 ();
 sg13g2_fill_2 FILLER_62_207 ();
 sg13g2_decap_4 FILLER_62_214 ();
 sg13g2_fill_1 FILLER_62_218 ();
 sg13g2_decap_4 FILLER_62_224 ();
 sg13g2_fill_1 FILLER_62_228 ();
 sg13g2_fill_1 FILLER_62_247 ();
 sg13g2_fill_2 FILLER_62_252 ();
 sg13g2_fill_1 FILLER_62_254 ();
 sg13g2_fill_2 FILLER_62_281 ();
 sg13g2_fill_1 FILLER_62_283 ();
 sg13g2_decap_8 FILLER_62_290 ();
 sg13g2_fill_1 FILLER_62_297 ();
 sg13g2_fill_2 FILLER_62_334 ();
 sg13g2_fill_2 FILLER_62_381 ();
 sg13g2_fill_1 FILLER_62_388 ();
 sg13g2_fill_2 FILLER_62_406 ();
 sg13g2_fill_1 FILLER_62_408 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_decap_8 FILLER_63_7 ();
 sg13g2_decap_8 FILLER_63_14 ();
 sg13g2_fill_1 FILLER_63_21 ();
 sg13g2_fill_2 FILLER_63_73 ();
 sg13g2_decap_8 FILLER_63_87 ();
 sg13g2_decap_8 FILLER_63_110 ();
 sg13g2_fill_2 FILLER_63_117 ();
 sg13g2_decap_4 FILLER_63_151 ();
 sg13g2_fill_1 FILLER_63_155 ();
 sg13g2_fill_2 FILLER_63_172 ();
 sg13g2_fill_1 FILLER_63_174 ();
 sg13g2_fill_2 FILLER_63_208 ();
 sg13g2_fill_2 FILLER_63_214 ();
 sg13g2_decap_8 FILLER_63_222 ();
 sg13g2_fill_2 FILLER_63_261 ();
 sg13g2_fill_1 FILLER_63_263 ();
 sg13g2_fill_1 FILLER_63_307 ();
 sg13g2_decap_8 FILLER_63_312 ();
 sg13g2_fill_2 FILLER_63_327 ();
 sg13g2_fill_1 FILLER_63_329 ();
 sg13g2_decap_8 FILLER_63_338 ();
 sg13g2_decap_4 FILLER_63_345 ();
 sg13g2_decap_8 FILLER_63_354 ();
 sg13g2_decap_4 FILLER_63_361 ();
 sg13g2_fill_2 FILLER_63_376 ();
 sg13g2_fill_1 FILLER_63_383 ();
 sg13g2_fill_2 FILLER_63_406 ();
 sg13g2_fill_1 FILLER_63_408 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_8 FILLER_64_7 ();
 sg13g2_decap_8 FILLER_64_14 ();
 sg13g2_decap_8 FILLER_64_21 ();
 sg13g2_decap_8 FILLER_64_28 ();
 sg13g2_decap_8 FILLER_64_35 ();
 sg13g2_fill_1 FILLER_64_42 ();
 sg13g2_decap_8 FILLER_64_60 ();
 sg13g2_fill_1 FILLER_64_67 ();
 sg13g2_fill_2 FILLER_64_73 ();
 sg13g2_fill_1 FILLER_64_75 ();
 sg13g2_fill_2 FILLER_64_92 ();
 sg13g2_fill_1 FILLER_64_112 ();
 sg13g2_fill_2 FILLER_64_124 ();
 sg13g2_decap_4 FILLER_64_139 ();
 sg13g2_decap_4 FILLER_64_146 ();
 sg13g2_fill_2 FILLER_64_171 ();
 sg13g2_fill_1 FILLER_64_173 ();
 sg13g2_decap_8 FILLER_64_180 ();
 sg13g2_decap_8 FILLER_64_187 ();
 sg13g2_fill_1 FILLER_64_194 ();
 sg13g2_fill_2 FILLER_64_204 ();
 sg13g2_fill_1 FILLER_64_215 ();
 sg13g2_decap_8 FILLER_64_237 ();
 sg13g2_decap_4 FILLER_64_244 ();
 sg13g2_decap_4 FILLER_64_252 ();
 sg13g2_fill_1 FILLER_64_256 ();
 sg13g2_decap_8 FILLER_64_265 ();
 sg13g2_fill_1 FILLER_64_272 ();
 sg13g2_fill_1 FILLER_64_281 ();
 sg13g2_fill_1 FILLER_64_318 ();
 sg13g2_decap_8 FILLER_64_339 ();
 sg13g2_decap_4 FILLER_64_350 ();
 sg13g2_fill_2 FILLER_64_354 ();
 sg13g2_fill_1 FILLER_64_361 ();
 sg13g2_fill_2 FILLER_64_377 ();
 sg13g2_fill_2 FILLER_64_391 ();
 sg13g2_fill_2 FILLER_64_398 ();
 sg13g2_fill_1 FILLER_64_400 ();
 sg13g2_fill_2 FILLER_64_406 ();
 sg13g2_fill_1 FILLER_64_408 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_8 FILLER_65_7 ();
 sg13g2_decap_8 FILLER_65_14 ();
 sg13g2_decap_8 FILLER_65_21 ();
 sg13g2_fill_1 FILLER_65_28 ();
 sg13g2_fill_1 FILLER_65_44 ();
 sg13g2_decap_4 FILLER_65_88 ();
 sg13g2_decap_8 FILLER_65_110 ();
 sg13g2_fill_2 FILLER_65_117 ();
 sg13g2_fill_1 FILLER_65_124 ();
 sg13g2_fill_2 FILLER_65_130 ();
 sg13g2_fill_1 FILLER_65_138 ();
 sg13g2_fill_1 FILLER_65_173 ();
 sg13g2_fill_1 FILLER_65_186 ();
 sg13g2_fill_1 FILLER_65_193 ();
 sg13g2_fill_2 FILLER_65_202 ();
 sg13g2_decap_4 FILLER_65_213 ();
 sg13g2_fill_1 FILLER_65_217 ();
 sg13g2_fill_1 FILLER_65_221 ();
 sg13g2_fill_2 FILLER_65_232 ();
 sg13g2_fill_1 FILLER_65_258 ();
 sg13g2_fill_2 FILLER_65_278 ();
 sg13g2_decap_8 FILLER_65_295 ();
 sg13g2_fill_2 FILLER_65_302 ();
 sg13g2_fill_1 FILLER_65_304 ();
 sg13g2_decap_4 FILLER_65_316 ();
 sg13g2_decap_8 FILLER_65_329 ();
 sg13g2_fill_2 FILLER_65_367 ();
 sg13g2_fill_2 FILLER_65_388 ();
 sg13g2_fill_1 FILLER_65_390 ();
 sg13g2_fill_1 FILLER_65_401 ();
 sg13g2_fill_2 FILLER_65_407 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_8 FILLER_66_7 ();
 sg13g2_decap_8 FILLER_66_14 ();
 sg13g2_decap_8 FILLER_66_21 ();
 sg13g2_fill_1 FILLER_66_28 ();
 sg13g2_fill_1 FILLER_66_37 ();
 sg13g2_fill_1 FILLER_66_49 ();
 sg13g2_fill_1 FILLER_66_56 ();
 sg13g2_decap_4 FILLER_66_67 ();
 sg13g2_fill_1 FILLER_66_71 ();
 sg13g2_fill_1 FILLER_66_92 ();
 sg13g2_fill_1 FILLER_66_97 ();
 sg13g2_fill_2 FILLER_66_103 ();
 sg13g2_fill_1 FILLER_66_120 ();
 sg13g2_decap_4 FILLER_66_136 ();
 sg13g2_fill_1 FILLER_66_152 ();
 sg13g2_fill_2 FILLER_66_161 ();
 sg13g2_fill_2 FILLER_66_173 ();
 sg13g2_fill_1 FILLER_66_179 ();
 sg13g2_fill_2 FILLER_66_188 ();
 sg13g2_fill_1 FILLER_66_190 ();
 sg13g2_fill_1 FILLER_66_205 ();
 sg13g2_decap_4 FILLER_66_225 ();
 sg13g2_fill_1 FILLER_66_229 ();
 sg13g2_fill_2 FILLER_66_235 ();
 sg13g2_fill_1 FILLER_66_237 ();
 sg13g2_fill_1 FILLER_66_242 ();
 sg13g2_decap_4 FILLER_66_248 ();
 sg13g2_fill_2 FILLER_66_275 ();
 sg13g2_fill_2 FILLER_66_285 ();
 sg13g2_fill_1 FILLER_66_300 ();
 sg13g2_fill_2 FILLER_66_311 ();
 sg13g2_fill_1 FILLER_66_325 ();
 sg13g2_fill_1 FILLER_66_347 ();
 sg13g2_fill_1 FILLER_66_364 ();
 sg13g2_decap_8 FILLER_66_371 ();
 sg13g2_fill_1 FILLER_66_378 ();
 sg13g2_fill_1 FILLER_66_387 ();
 sg13g2_fill_1 FILLER_66_408 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_8 FILLER_67_7 ();
 sg13g2_decap_8 FILLER_67_14 ();
 sg13g2_decap_8 FILLER_67_21 ();
 sg13g2_decap_8 FILLER_67_28 ();
 sg13g2_decap_4 FILLER_67_35 ();
 sg13g2_decap_4 FILLER_67_44 ();
 sg13g2_decap_4 FILLER_67_53 ();
 sg13g2_fill_2 FILLER_67_57 ();
 sg13g2_fill_2 FILLER_67_71 ();
 sg13g2_fill_1 FILLER_67_73 ();
 sg13g2_decap_8 FILLER_67_79 ();
 sg13g2_fill_2 FILLER_67_94 ();
 sg13g2_fill_2 FILLER_67_102 ();
 sg13g2_fill_2 FILLER_67_115 ();
 sg13g2_decap_8 FILLER_67_120 ();
 sg13g2_fill_1 FILLER_67_127 ();
 sg13g2_fill_1 FILLER_67_133 ();
 sg13g2_decap_8 FILLER_67_139 ();
 sg13g2_fill_2 FILLER_67_146 ();
 sg13g2_fill_1 FILLER_67_148 ();
 sg13g2_decap_4 FILLER_67_154 ();
 sg13g2_fill_2 FILLER_67_158 ();
 sg13g2_fill_2 FILLER_67_168 ();
 sg13g2_fill_1 FILLER_67_170 ();
 sg13g2_decap_8 FILLER_67_180 ();
 sg13g2_fill_1 FILLER_67_187 ();
 sg13g2_decap_4 FILLER_67_199 ();
 sg13g2_decap_4 FILLER_67_212 ();
 sg13g2_fill_2 FILLER_67_220 ();
 sg13g2_fill_1 FILLER_67_222 ();
 sg13g2_fill_2 FILLER_67_227 ();
 sg13g2_fill_2 FILLER_67_232 ();
 sg13g2_fill_2 FILLER_67_247 ();
 sg13g2_fill_1 FILLER_67_249 ();
 sg13g2_fill_2 FILLER_67_263 ();
 sg13g2_fill_1 FILLER_67_265 ();
 sg13g2_decap_4 FILLER_67_271 ();
 sg13g2_fill_1 FILLER_67_275 ();
 sg13g2_fill_2 FILLER_67_288 ();
 sg13g2_decap_4 FILLER_67_298 ();
 sg13g2_fill_1 FILLER_67_302 ();
 sg13g2_fill_1 FILLER_67_312 ();
 sg13g2_decap_8 FILLER_67_328 ();
 sg13g2_decap_8 FILLER_67_335 ();
 sg13g2_fill_1 FILLER_67_342 ();
 sg13g2_decap_8 FILLER_67_356 ();
 sg13g2_decap_4 FILLER_67_371 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_8 FILLER_68_7 ();
 sg13g2_decap_8 FILLER_68_14 ();
 sg13g2_decap_8 FILLER_68_21 ();
 sg13g2_decap_8 FILLER_68_28 ();
 sg13g2_decap_4 FILLER_68_35 ();
 sg13g2_fill_1 FILLER_68_39 ();
 sg13g2_fill_1 FILLER_68_48 ();
 sg13g2_decap_8 FILLER_68_67 ();
 sg13g2_decap_8 FILLER_68_74 ();
 sg13g2_fill_1 FILLER_68_91 ();
 sg13g2_decap_8 FILLER_68_96 ();
 sg13g2_decap_4 FILLER_68_103 ();
 sg13g2_fill_2 FILLER_68_107 ();
 sg13g2_fill_2 FILLER_68_119 ();
 sg13g2_fill_2 FILLER_68_133 ();
 sg13g2_fill_1 FILLER_68_135 ();
 sg13g2_fill_2 FILLER_68_147 ();
 sg13g2_fill_2 FILLER_68_157 ();
 sg13g2_fill_1 FILLER_68_159 ();
 sg13g2_fill_1 FILLER_68_168 ();
 sg13g2_fill_2 FILLER_68_194 ();
 sg13g2_fill_1 FILLER_68_205 ();
 sg13g2_decap_4 FILLER_68_217 ();
 sg13g2_fill_2 FILLER_68_239 ();
 sg13g2_fill_1 FILLER_68_241 ();
 sg13g2_decap_4 FILLER_68_275 ();
 sg13g2_fill_2 FILLER_68_285 ();
 sg13g2_fill_1 FILLER_68_287 ();
 sg13g2_decap_8 FILLER_68_293 ();
 sg13g2_decap_8 FILLER_68_300 ();
 sg13g2_fill_2 FILLER_68_307 ();
 sg13g2_decap_8 FILLER_68_319 ();
 sg13g2_fill_1 FILLER_68_326 ();
 sg13g2_fill_1 FILLER_68_338 ();
 sg13g2_fill_2 FILLER_68_348 ();
 sg13g2_fill_2 FILLER_68_371 ();
 sg13g2_decap_4 FILLER_68_378 ();
 sg13g2_fill_2 FILLER_68_398 ();
 sg13g2_fill_1 FILLER_68_408 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_8 FILLER_69_7 ();
 sg13g2_decap_8 FILLER_69_14 ();
 sg13g2_decap_8 FILLER_69_21 ();
 sg13g2_decap_8 FILLER_69_28 ();
 sg13g2_decap_8 FILLER_69_35 ();
 sg13g2_fill_1 FILLER_69_42 ();
 sg13g2_decap_4 FILLER_69_53 ();
 sg13g2_fill_1 FILLER_69_57 ();
 sg13g2_fill_2 FILLER_69_79 ();
 sg13g2_fill_2 FILLER_69_91 ();
 sg13g2_fill_2 FILLER_69_106 ();
 sg13g2_fill_2 FILLER_69_127 ();
 sg13g2_decap_4 FILLER_69_142 ();
 sg13g2_fill_2 FILLER_69_146 ();
 sg13g2_decap_8 FILLER_69_155 ();
 sg13g2_fill_2 FILLER_69_162 ();
 sg13g2_fill_1 FILLER_69_164 ();
 sg13g2_fill_2 FILLER_69_174 ();
 sg13g2_fill_1 FILLER_69_176 ();
 sg13g2_fill_1 FILLER_69_181 ();
 sg13g2_decap_4 FILLER_69_187 ();
 sg13g2_fill_1 FILLER_69_191 ();
 sg13g2_decap_4 FILLER_69_200 ();
 sg13g2_fill_2 FILLER_69_204 ();
 sg13g2_decap_4 FILLER_69_211 ();
 sg13g2_decap_8 FILLER_69_228 ();
 sg13g2_fill_2 FILLER_69_235 ();
 sg13g2_fill_2 FILLER_69_250 ();
 sg13g2_fill_1 FILLER_69_252 ();
 sg13g2_decap_4 FILLER_69_258 ();
 sg13g2_fill_1 FILLER_69_262 ();
 sg13g2_fill_2 FILLER_69_271 ();
 sg13g2_fill_1 FILLER_69_277 ();
 sg13g2_fill_2 FILLER_69_286 ();
 sg13g2_fill_1 FILLER_69_288 ();
 sg13g2_fill_2 FILLER_69_316 ();
 sg13g2_fill_2 FILLER_69_357 ();
 sg13g2_fill_1 FILLER_69_359 ();
 sg13g2_fill_1 FILLER_69_384 ();
 sg13g2_fill_1 FILLER_69_394 ();
 sg13g2_fill_2 FILLER_69_407 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_decap_8 FILLER_70_14 ();
 sg13g2_decap_8 FILLER_70_21 ();
 sg13g2_decap_8 FILLER_70_28 ();
 sg13g2_decap_8 FILLER_70_35 ();
 sg13g2_decap_4 FILLER_70_42 ();
 sg13g2_fill_1 FILLER_70_46 ();
 sg13g2_decap_4 FILLER_70_57 ();
 sg13g2_fill_1 FILLER_70_61 ();
 sg13g2_decap_4 FILLER_70_70 ();
 sg13g2_fill_2 FILLER_70_74 ();
 sg13g2_decap_4 FILLER_70_93 ();
 sg13g2_fill_1 FILLER_70_97 ();
 sg13g2_fill_2 FILLER_70_103 ();
 sg13g2_decap_4 FILLER_70_114 ();
 sg13g2_fill_2 FILLER_70_126 ();
 sg13g2_fill_2 FILLER_70_133 ();
 sg13g2_fill_1 FILLER_70_135 ();
 sg13g2_fill_1 FILLER_70_140 ();
 sg13g2_decap_4 FILLER_70_146 ();
 sg13g2_fill_2 FILLER_70_176 ();
 sg13g2_fill_2 FILLER_70_186 ();
 sg13g2_fill_1 FILLER_70_188 ();
 sg13g2_decap_4 FILLER_70_207 ();
 sg13g2_fill_1 FILLER_70_224 ();
 sg13g2_fill_2 FILLER_70_246 ();
 sg13g2_fill_2 FILLER_70_292 ();
 sg13g2_fill_1 FILLER_70_294 ();
 sg13g2_decap_8 FILLER_70_301 ();
 sg13g2_fill_1 FILLER_70_308 ();
 sg13g2_fill_1 FILLER_70_313 ();
 sg13g2_fill_1 FILLER_70_318 ();
 sg13g2_decap_8 FILLER_70_323 ();
 sg13g2_decap_4 FILLER_70_330 ();
 sg13g2_fill_2 FILLER_70_334 ();
 sg13g2_fill_2 FILLER_70_346 ();
 sg13g2_decap_4 FILLER_70_361 ();
 sg13g2_fill_2 FILLER_70_365 ();
 sg13g2_fill_2 FILLER_70_371 ();
 sg13g2_fill_2 FILLER_70_377 ();
 sg13g2_decap_4 FILLER_70_395 ();
 sg13g2_fill_2 FILLER_70_399 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_decap_8 FILLER_71_7 ();
 sg13g2_decap_8 FILLER_71_14 ();
 sg13g2_decap_8 FILLER_71_21 ();
 sg13g2_decap_8 FILLER_71_28 ();
 sg13g2_decap_8 FILLER_71_35 ();
 sg13g2_fill_2 FILLER_71_42 ();
 sg13g2_fill_1 FILLER_71_52 ();
 sg13g2_fill_1 FILLER_71_61 ();
 sg13g2_decap_4 FILLER_71_82 ();
 sg13g2_fill_2 FILLER_71_86 ();
 sg13g2_fill_1 FILLER_71_96 ();
 sg13g2_fill_2 FILLER_71_103 ();
 sg13g2_fill_1 FILLER_71_115 ();
 sg13g2_fill_2 FILLER_71_122 ();
 sg13g2_fill_1 FILLER_71_153 ();
 sg13g2_decap_8 FILLER_71_157 ();
 sg13g2_fill_1 FILLER_71_164 ();
 sg13g2_fill_2 FILLER_71_169 ();
 sg13g2_fill_1 FILLER_71_171 ();
 sg13g2_fill_2 FILLER_71_184 ();
 sg13g2_decap_8 FILLER_71_190 ();
 sg13g2_decap_4 FILLER_71_197 ();
 sg13g2_decap_8 FILLER_71_209 ();
 sg13g2_decap_8 FILLER_71_221 ();
 sg13g2_decap_8 FILLER_71_228 ();
 sg13g2_decap_4 FILLER_71_235 ();
 sg13g2_fill_1 FILLER_71_239 ();
 sg13g2_decap_8 FILLER_71_249 ();
 sg13g2_fill_2 FILLER_71_261 ();
 sg13g2_fill_1 FILLER_71_263 ();
 sg13g2_decap_4 FILLER_71_272 ();
 sg13g2_fill_2 FILLER_71_276 ();
 sg13g2_fill_2 FILLER_71_300 ();
 sg13g2_fill_2 FILLER_71_325 ();
 sg13g2_fill_1 FILLER_71_327 ();
 sg13g2_fill_2 FILLER_71_336 ();
 sg13g2_decap_8 FILLER_71_365 ();
 sg13g2_decap_8 FILLER_71_372 ();
 sg13g2_decap_8 FILLER_71_379 ();
 sg13g2_decap_8 FILLER_71_386 ();
 sg13g2_decap_8 FILLER_71_393 ();
 sg13g2_decap_8 FILLER_71_400 ();
 sg13g2_fill_2 FILLER_71_407 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_decap_8 FILLER_72_14 ();
 sg13g2_decap_8 FILLER_72_21 ();
 sg13g2_decap_8 FILLER_72_28 ();
 sg13g2_decap_8 FILLER_72_35 ();
 sg13g2_decap_4 FILLER_72_42 ();
 sg13g2_fill_1 FILLER_72_46 ();
 sg13g2_decap_8 FILLER_72_52 ();
 sg13g2_decap_4 FILLER_72_59 ();
 sg13g2_decap_8 FILLER_72_71 ();
 sg13g2_fill_2 FILLER_72_78 ();
 sg13g2_fill_1 FILLER_72_80 ();
 sg13g2_decap_8 FILLER_72_101 ();
 sg13g2_decap_8 FILLER_72_113 ();
 sg13g2_fill_1 FILLER_72_132 ();
 sg13g2_fill_1 FILLER_72_138 ();
 sg13g2_fill_2 FILLER_72_143 ();
 sg13g2_fill_2 FILLER_72_150 ();
 sg13g2_decap_4 FILLER_72_165 ();
 sg13g2_fill_1 FILLER_72_169 ();
 sg13g2_fill_2 FILLER_72_175 ();
 sg13g2_fill_1 FILLER_72_181 ();
 sg13g2_fill_2 FILLER_72_204 ();
 sg13g2_fill_1 FILLER_72_206 ();
 sg13g2_decap_4 FILLER_72_220 ();
 sg13g2_decap_8 FILLER_72_251 ();
 sg13g2_decap_8 FILLER_72_258 ();
 sg13g2_decap_8 FILLER_72_265 ();
 sg13g2_decap_8 FILLER_72_280 ();
 sg13g2_fill_2 FILLER_72_287 ();
 sg13g2_fill_1 FILLER_72_299 ();
 sg13g2_decap_4 FILLER_72_304 ();
 sg13g2_decap_4 FILLER_72_311 ();
 sg13g2_fill_2 FILLER_72_315 ();
 sg13g2_fill_1 FILLER_72_324 ();
 sg13g2_fill_2 FILLER_72_333 ();
 sg13g2_fill_1 FILLER_72_335 ();
 sg13g2_decap_8 FILLER_72_342 ();
 sg13g2_decap_8 FILLER_72_370 ();
 sg13g2_decap_8 FILLER_72_377 ();
 sg13g2_decap_8 FILLER_72_384 ();
 sg13g2_decap_8 FILLER_72_391 ();
 sg13g2_decap_8 FILLER_72_398 ();
 sg13g2_decap_4 FILLER_72_405 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_decap_8 FILLER_73_14 ();
 sg13g2_decap_8 FILLER_73_21 ();
 sg13g2_decap_8 FILLER_73_28 ();
 sg13g2_decap_8 FILLER_73_35 ();
 sg13g2_decap_8 FILLER_73_42 ();
 sg13g2_decap_8 FILLER_73_49 ();
 sg13g2_decap_8 FILLER_73_56 ();
 sg13g2_decap_8 FILLER_73_63 ();
 sg13g2_decap_8 FILLER_73_70 ();
 sg13g2_decap_8 FILLER_73_77 ();
 sg13g2_decap_8 FILLER_73_84 ();
 sg13g2_fill_2 FILLER_73_127 ();
 sg13g2_fill_1 FILLER_73_129 ();
 sg13g2_fill_2 FILLER_73_137 ();
 sg13g2_fill_2 FILLER_73_147 ();
 sg13g2_fill_1 FILLER_73_149 ();
 sg13g2_fill_2 FILLER_73_193 ();
 sg13g2_fill_1 FILLER_73_206 ();
 sg13g2_fill_2 FILLER_73_212 ();
 sg13g2_fill_1 FILLER_73_214 ();
 sg13g2_decap_8 FILLER_73_231 ();
 sg13g2_fill_2 FILLER_73_238 ();
 sg13g2_fill_1 FILLER_73_240 ();
 sg13g2_fill_2 FILLER_73_246 ();
 sg13g2_fill_1 FILLER_73_271 ();
 sg13g2_decap_8 FILLER_73_280 ();
 sg13g2_fill_1 FILLER_73_300 ();
 sg13g2_fill_1 FILLER_73_320 ();
 sg13g2_decap_4 FILLER_73_338 ();
 sg13g2_fill_2 FILLER_73_351 ();
 sg13g2_fill_1 FILLER_73_353 ();
 sg13g2_fill_2 FILLER_73_357 ();
 sg13g2_fill_1 FILLER_73_359 ();
 sg13g2_decap_8 FILLER_73_365 ();
 sg13g2_decap_8 FILLER_73_372 ();
 sg13g2_decap_8 FILLER_73_379 ();
 sg13g2_decap_8 FILLER_73_386 ();
 sg13g2_decap_8 FILLER_73_393 ();
 sg13g2_decap_8 FILLER_73_400 ();
 sg13g2_fill_2 FILLER_73_407 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_decap_8 FILLER_74_14 ();
 sg13g2_decap_8 FILLER_74_21 ();
 sg13g2_decap_8 FILLER_74_28 ();
 sg13g2_decap_8 FILLER_74_35 ();
 sg13g2_decap_8 FILLER_74_42 ();
 sg13g2_decap_8 FILLER_74_49 ();
 sg13g2_decap_8 FILLER_74_56 ();
 sg13g2_decap_8 FILLER_74_63 ();
 sg13g2_decap_8 FILLER_74_70 ();
 sg13g2_decap_8 FILLER_74_77 ();
 sg13g2_decap_4 FILLER_74_84 ();
 sg13g2_fill_1 FILLER_74_88 ();
 sg13g2_decap_8 FILLER_74_94 ();
 sg13g2_fill_1 FILLER_74_101 ();
 sg13g2_fill_1 FILLER_74_107 ();
 sg13g2_fill_2 FILLER_74_113 ();
 sg13g2_fill_1 FILLER_74_115 ();
 sg13g2_decap_4 FILLER_74_121 ();
 sg13g2_fill_1 FILLER_74_125 ();
 sg13g2_decap_4 FILLER_74_138 ();
 sg13g2_decap_4 FILLER_74_146 ();
 sg13g2_fill_1 FILLER_74_150 ();
 sg13g2_fill_2 FILLER_74_163 ();
 sg13g2_fill_1 FILLER_74_165 ();
 sg13g2_decap_8 FILLER_74_171 ();
 sg13g2_decap_8 FILLER_74_192 ();
 sg13g2_fill_2 FILLER_74_213 ();
 sg13g2_fill_2 FILLER_74_222 ();
 sg13g2_fill_1 FILLER_74_224 ();
 sg13g2_fill_2 FILLER_74_238 ();
 sg13g2_fill_1 FILLER_74_240 ();
 sg13g2_fill_1 FILLER_74_249 ();
 sg13g2_fill_1 FILLER_74_255 ();
 sg13g2_fill_2 FILLER_74_279 ();
 sg13g2_decap_4 FILLER_74_308 ();
 sg13g2_fill_1 FILLER_74_312 ();
 sg13g2_fill_2 FILLER_74_325 ();
 sg13g2_fill_1 FILLER_74_327 ();
 sg13g2_fill_2 FILLER_74_343 ();
 sg13g2_fill_1 FILLER_74_353 ();
 sg13g2_decap_8 FILLER_74_367 ();
 sg13g2_decap_8 FILLER_74_374 ();
 sg13g2_decap_8 FILLER_74_381 ();
 sg13g2_decap_8 FILLER_74_388 ();
 sg13g2_decap_8 FILLER_74_395 ();
 sg13g2_decap_8 FILLER_74_402 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_14 ();
 sg13g2_decap_8 FILLER_75_21 ();
 sg13g2_decap_8 FILLER_75_28 ();
 sg13g2_decap_8 FILLER_75_35 ();
 sg13g2_decap_8 FILLER_75_42 ();
 sg13g2_decap_8 FILLER_75_49 ();
 sg13g2_decap_8 FILLER_75_56 ();
 sg13g2_decap_8 FILLER_75_63 ();
 sg13g2_decap_8 FILLER_75_70 ();
 sg13g2_decap_4 FILLER_75_77 ();
 sg13g2_fill_2 FILLER_75_81 ();
 sg13g2_fill_2 FILLER_75_99 ();
 sg13g2_decap_4 FILLER_75_105 ();
 sg13g2_decap_8 FILLER_75_130 ();
 sg13g2_fill_2 FILLER_75_137 ();
 sg13g2_fill_1 FILLER_75_139 ();
 sg13g2_decap_8 FILLER_75_154 ();
 sg13g2_fill_2 FILLER_75_161 ();
 sg13g2_fill_2 FILLER_75_175 ();
 sg13g2_fill_1 FILLER_75_177 ();
 sg13g2_decap_4 FILLER_75_199 ();
 sg13g2_fill_1 FILLER_75_203 ();
 sg13g2_fill_1 FILLER_75_228 ();
 sg13g2_fill_2 FILLER_75_234 ();
 sg13g2_fill_1 FILLER_75_236 ();
 sg13g2_decap_8 FILLER_75_263 ();
 sg13g2_decap_4 FILLER_75_270 ();
 sg13g2_decap_8 FILLER_75_284 ();
 sg13g2_decap_8 FILLER_75_291 ();
 sg13g2_fill_2 FILLER_75_298 ();
 sg13g2_fill_2 FILLER_75_315 ();
 sg13g2_decap_4 FILLER_75_324 ();
 sg13g2_fill_1 FILLER_75_333 ();
 sg13g2_fill_2 FILLER_75_344 ();
 sg13g2_decap_4 FILLER_75_356 ();
 sg13g2_fill_2 FILLER_75_360 ();
 sg13g2_decap_8 FILLER_75_367 ();
 sg13g2_decap_8 FILLER_75_374 ();
 sg13g2_decap_8 FILLER_75_381 ();
 sg13g2_decap_8 FILLER_75_388 ();
 sg13g2_decap_8 FILLER_75_395 ();
 sg13g2_decap_8 FILLER_75_402 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_8 FILLER_76_21 ();
 sg13g2_decap_8 FILLER_76_28 ();
 sg13g2_decap_8 FILLER_76_35 ();
 sg13g2_decap_8 FILLER_76_42 ();
 sg13g2_decap_8 FILLER_76_49 ();
 sg13g2_decap_8 FILLER_76_56 ();
 sg13g2_decap_8 FILLER_76_63 ();
 sg13g2_decap_8 FILLER_76_70 ();
 sg13g2_decap_8 FILLER_76_77 ();
 sg13g2_decap_4 FILLER_76_84 ();
 sg13g2_fill_2 FILLER_76_113 ();
 sg13g2_fill_1 FILLER_76_140 ();
 sg13g2_fill_2 FILLER_76_176 ();
 sg13g2_fill_1 FILLER_76_178 ();
 sg13g2_decap_4 FILLER_76_191 ();
 sg13g2_fill_2 FILLER_76_195 ();
 sg13g2_fill_1 FILLER_76_201 ();
 sg13g2_fill_2 FILLER_76_207 ();
 sg13g2_decap_4 FILLER_76_212 ();
 sg13g2_fill_1 FILLER_76_216 ();
 sg13g2_decap_4 FILLER_76_225 ();
 sg13g2_fill_2 FILLER_76_238 ();
 sg13g2_fill_1 FILLER_76_240 ();
 sg13g2_fill_2 FILLER_76_245 ();
 sg13g2_fill_1 FILLER_76_247 ();
 sg13g2_fill_2 FILLER_76_253 ();
 sg13g2_fill_2 FILLER_76_263 ();
 sg13g2_fill_1 FILLER_76_265 ();
 sg13g2_decap_8 FILLER_76_279 ();
 sg13g2_fill_1 FILLER_76_303 ();
 sg13g2_fill_2 FILLER_76_312 ();
 sg13g2_fill_2 FILLER_76_322 ();
 sg13g2_fill_2 FILLER_76_345 ();
 sg13g2_fill_1 FILLER_76_360 ();
 sg13g2_decap_8 FILLER_76_374 ();
 sg13g2_decap_8 FILLER_76_381 ();
 sg13g2_decap_8 FILLER_76_388 ();
 sg13g2_decap_8 FILLER_76_395 ();
 sg13g2_decap_8 FILLER_76_402 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_decap_8 FILLER_77_28 ();
 sg13g2_decap_8 FILLER_77_35 ();
 sg13g2_decap_8 FILLER_77_42 ();
 sg13g2_decap_8 FILLER_77_49 ();
 sg13g2_decap_8 FILLER_77_56 ();
 sg13g2_decap_8 FILLER_77_63 ();
 sg13g2_decap_8 FILLER_77_70 ();
 sg13g2_decap_8 FILLER_77_77 ();
 sg13g2_decap_4 FILLER_77_84 ();
 sg13g2_fill_1 FILLER_77_88 ();
 sg13g2_fill_2 FILLER_77_98 ();
 sg13g2_fill_2 FILLER_77_107 ();
 sg13g2_fill_1 FILLER_77_122 ();
 sg13g2_decap_4 FILLER_77_128 ();
 sg13g2_fill_1 FILLER_77_137 ();
 sg13g2_decap_8 FILLER_77_143 ();
 sg13g2_decap_8 FILLER_77_150 ();
 sg13g2_decap_4 FILLER_77_157 ();
 sg13g2_fill_1 FILLER_77_161 ();
 sg13g2_decap_8 FILLER_77_167 ();
 sg13g2_fill_2 FILLER_77_174 ();
 sg13g2_fill_2 FILLER_77_205 ();
 sg13g2_fill_1 FILLER_77_207 ();
 sg13g2_fill_2 FILLER_77_221 ();
 sg13g2_fill_2 FILLER_77_239 ();
 sg13g2_fill_1 FILLER_77_255 ();
 sg13g2_fill_1 FILLER_77_272 ();
 sg13g2_fill_1 FILLER_77_299 ();
 sg13g2_fill_1 FILLER_77_305 ();
 sg13g2_decap_4 FILLER_77_311 ();
 sg13g2_fill_1 FILLER_77_315 ();
 sg13g2_decap_4 FILLER_77_323 ();
 sg13g2_decap_4 FILLER_77_332 ();
 sg13g2_fill_1 FILLER_77_336 ();
 sg13g2_decap_4 FILLER_77_345 ();
 sg13g2_fill_2 FILLER_77_349 ();
 sg13g2_fill_1 FILLER_77_359 ();
 sg13g2_decap_8 FILLER_77_368 ();
 sg13g2_decap_8 FILLER_77_375 ();
 sg13g2_decap_8 FILLER_77_382 ();
 sg13g2_decap_8 FILLER_77_389 ();
 sg13g2_decap_8 FILLER_77_396 ();
 sg13g2_decap_4 FILLER_77_403 ();
 sg13g2_fill_2 FILLER_77_407 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_decap_8 FILLER_78_28 ();
 sg13g2_decap_8 FILLER_78_35 ();
 sg13g2_decap_8 FILLER_78_42 ();
 sg13g2_decap_8 FILLER_78_49 ();
 sg13g2_decap_8 FILLER_78_56 ();
 sg13g2_decap_8 FILLER_78_63 ();
 sg13g2_decap_8 FILLER_78_70 ();
 sg13g2_decap_8 FILLER_78_77 ();
 sg13g2_decap_4 FILLER_78_84 ();
 sg13g2_fill_2 FILLER_78_88 ();
 sg13g2_decap_4 FILLER_78_98 ();
 sg13g2_fill_1 FILLER_78_102 ();
 sg13g2_decap_4 FILLER_78_120 ();
 sg13g2_fill_1 FILLER_78_124 ();
 sg13g2_fill_2 FILLER_78_130 ();
 sg13g2_fill_1 FILLER_78_132 ();
 sg13g2_fill_1 FILLER_78_144 ();
 sg13g2_fill_1 FILLER_78_155 ();
 sg13g2_fill_2 FILLER_78_170 ();
 sg13g2_fill_1 FILLER_78_172 ();
 sg13g2_fill_2 FILLER_78_182 ();
 sg13g2_decap_4 FILLER_78_202 ();
 sg13g2_fill_2 FILLER_78_206 ();
 sg13g2_fill_1 FILLER_78_230 ();
 sg13g2_decap_8 FILLER_78_241 ();
 sg13g2_fill_1 FILLER_78_248 ();
 sg13g2_fill_1 FILLER_78_259 ();
 sg13g2_fill_1 FILLER_78_270 ();
 sg13g2_fill_1 FILLER_78_279 ();
 sg13g2_fill_2 FILLER_78_285 ();
 sg13g2_fill_2 FILLER_78_296 ();
 sg13g2_fill_2 FILLER_78_307 ();
 sg13g2_decap_4 FILLER_78_320 ();
 sg13g2_fill_2 FILLER_78_324 ();
 sg13g2_fill_2 FILLER_78_331 ();
 sg13g2_fill_1 FILLER_78_333 ();
 sg13g2_decap_8 FILLER_78_348 ();
 sg13g2_decap_4 FILLER_78_355 ();
 sg13g2_fill_1 FILLER_78_359 ();
 sg13g2_decap_8 FILLER_78_369 ();
 sg13g2_decap_8 FILLER_78_376 ();
 sg13g2_decap_8 FILLER_78_383 ();
 sg13g2_decap_8 FILLER_78_390 ();
 sg13g2_decap_8 FILLER_78_397 ();
 sg13g2_decap_4 FILLER_78_404 ();
 sg13g2_fill_1 FILLER_78_408 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_decap_8 FILLER_79_35 ();
 sg13g2_decap_8 FILLER_79_42 ();
 sg13g2_decap_8 FILLER_79_49 ();
 sg13g2_decap_8 FILLER_79_56 ();
 sg13g2_decap_8 FILLER_79_63 ();
 sg13g2_decap_8 FILLER_79_70 ();
 sg13g2_decap_8 FILLER_79_77 ();
 sg13g2_decap_8 FILLER_79_84 ();
 sg13g2_fill_2 FILLER_79_91 ();
 sg13g2_fill_1 FILLER_79_93 ();
 sg13g2_fill_1 FILLER_79_110 ();
 sg13g2_fill_1 FILLER_79_123 ();
 sg13g2_decap_4 FILLER_79_137 ();
 sg13g2_decap_8 FILLER_79_145 ();
 sg13g2_decap_8 FILLER_79_152 ();
 sg13g2_fill_1 FILLER_79_159 ();
 sg13g2_fill_2 FILLER_79_173 ();
 sg13g2_fill_1 FILLER_79_175 ();
 sg13g2_fill_1 FILLER_79_191 ();
 sg13g2_fill_1 FILLER_79_222 ();
 sg13g2_fill_1 FILLER_79_231 ();
 sg13g2_fill_1 FILLER_79_239 ();
 sg13g2_fill_1 FILLER_79_306 ();
 sg13g2_decap_8 FILLER_79_374 ();
 sg13g2_decap_8 FILLER_79_381 ();
 sg13g2_decap_8 FILLER_79_388 ();
 sg13g2_decap_8 FILLER_79_395 ();
 sg13g2_decap_8 FILLER_79_402 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_42 ();
 sg13g2_decap_8 FILLER_80_49 ();
 sg13g2_decap_4 FILLER_80_60 ();
 sg13g2_decap_4 FILLER_80_68 ();
 sg13g2_decap_4 FILLER_80_76 ();
 sg13g2_decap_4 FILLER_80_84 ();
 sg13g2_decap_4 FILLER_80_92 ();
 sg13g2_decap_4 FILLER_80_100 ();
 sg13g2_fill_2 FILLER_80_108 ();
 sg13g2_fill_2 FILLER_80_142 ();
 sg13g2_decap_4 FILLER_80_148 ();
 sg13g2_decap_4 FILLER_80_156 ();
 sg13g2_fill_2 FILLER_80_164 ();
 sg13g2_decap_4 FILLER_80_182 ();
 sg13g2_fill_1 FILLER_80_186 ();
 sg13g2_decap_4 FILLER_80_190 ();
 sg13g2_fill_1 FILLER_80_194 ();
 sg13g2_decap_8 FILLER_80_200 ();
 sg13g2_decap_8 FILLER_80_207 ();
 sg13g2_decap_4 FILLER_80_228 ();
 sg13g2_fill_1 FILLER_80_232 ();
 sg13g2_decap_8 FILLER_80_238 ();
 sg13g2_decap_8 FILLER_80_245 ();
 sg13g2_decap_4 FILLER_80_256 ();
 sg13g2_decap_8 FILLER_80_265 ();
 sg13g2_decap_8 FILLER_80_272 ();
 sg13g2_decap_4 FILLER_80_279 ();
 sg13g2_fill_2 FILLER_80_283 ();
 sg13g2_decap_8 FILLER_80_295 ();
 sg13g2_fill_2 FILLER_80_310 ();
 sg13g2_fill_1 FILLER_80_312 ();
 sg13g2_decap_8 FILLER_80_318 ();
 sg13g2_decap_8 FILLER_80_329 ();
 sg13g2_decap_8 FILLER_80_340 ();
 sg13g2_decap_8 FILLER_80_347 ();
 sg13g2_fill_2 FILLER_80_354 ();
 sg13g2_fill_1 FILLER_80_356 ();
 sg13g2_decap_8 FILLER_80_366 ();
 sg13g2_fill_2 FILLER_80_373 ();
 sg13g2_fill_1 FILLER_80_375 ();
 sg13g2_decap_8 FILLER_80_384 ();
 sg13g2_decap_8 FILLER_80_391 ();
 sg13g2_decap_8 FILLER_80_398 ();
 sg13g2_decap_4 FILLER_80_405 ();
 assign uio_oe[0] = net2;
 assign uio_oe[1] = net3;
 assign uio_oe[2] = net4;
 assign uio_oe[3] = net5;
 assign uio_oe[4] = net6;
 assign uio_oe[5] = net7;
 assign uio_oe[6] = net8;
 assign uio_oe[7] = net9;
 assign uio_out[0] = net10;
 assign uio_out[1] = net11;
 assign uio_out[2] = net12;
 assign uio_out[3] = net13;
 assign uio_out[4] = net14;
 assign uio_out[5] = net15;
 assign uio_out[6] = net16;
 assign uio_out[7] = net17;
endmodule

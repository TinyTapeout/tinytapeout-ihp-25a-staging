module tt_um_wokwi_group_2 (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire \proj_10.net10 ;
 wire \proj_10.net11 ;
 wire \proj_10.net12 ;
 wire \proj_10.net13 ;
 wire \proj_10.net14 ;
 wire \proj_10.net15 ;
 wire \proj_10.net16 ;
 wire \proj_10.net17 ;
 wire \proj_10.net23 ;
 wire \proj_10.net24 ;
 wire \proj_10.net25 ;
 wire \proj_10.net26 ;
 wire \proj_10.net27 ;
 wire \proj_10.net28 ;
 wire \proj_10.net29 ;
 wire \proj_10.net30 ;
 wire \proj_10.net31 ;
 wire \proj_10.net32 ;
 wire \proj_10.net33 ;
 wire \proj_10.net34 ;
 wire \proj_10.net35 ;
 wire \proj_10.net36 ;
 wire \proj_10.net37 ;
 wire \proj_10.net38 ;
 wire \proj_10.net39 ;
 wire \proj_10.net40 ;
 wire \proj_10.net41 ;
 wire \proj_10.net42 ;
 wire \proj_10.net43 ;
 wire \proj_10.net44 ;
 wire \proj_10.net45 ;
 wire \proj_10.net46 ;
 wire \proj_11.net10 ;
 wire \proj_11.net11 ;
 wire \proj_11.net12 ;
 wire \proj_11.net13 ;
 wire \proj_11.net19 ;
 wire \proj_11.net20 ;
 wire \proj_11.net21 ;
 wire \proj_11.net22 ;
 wire \proj_11.net23 ;
 wire \proj_11.net24 ;
 wire \proj_11.net25 ;
 wire \proj_11.net26 ;
 wire \proj_11.net27 ;
 wire \proj_11.net28 ;
 wire \proj_11.net29 ;
 wire \proj_11.net30 ;
 wire \proj_11.net9 ;
 wire clk_regs;
 wire \proj_12.net12 ;
 wire \proj_12.net13 ;
 wire \proj_12.net14 ;
 wire \proj_12.net20 ;
 wire \proj_12.net21 ;
 wire \proj_12.net22 ;
 wire \proj_13.net10 ;
 wire \proj_13.net11 ;
 wire \proj_13.net12 ;
 wire \proj_13.net13 ;
 wire \proj_13.net14 ;
 wire \proj_13.net20 ;
 wire \proj_13.net21 ;
 wire \proj_13.net22 ;
 wire \proj_13.net23 ;
 wire \proj_13.net24 ;
 wire \proj_13.net9 ;
 wire \proj_14.net100 ;
 wire \proj_14.net102 ;
 wire \proj_14.net103 ;
 wire \proj_14.net105 ;
 wire \proj_14.net106 ;
 wire \proj_14.net108 ;
 wire \proj_14.net109 ;
 wire \proj_14.net11 ;
 wire \proj_14.net111 ;
 wire \proj_14.net112 ;
 wire \proj_14.net114 ;
 wire \proj_14.net116 ;
 wire \proj_14.net118 ;
 wire \proj_14.net119 ;
 wire \proj_14.net12 ;
 wire \proj_14.net121 ;
 wire \proj_14.net122 ;
 wire \proj_14.net124 ;
 wire \proj_14.net125 ;
 wire \proj_14.net127 ;
 wire \proj_14.net128 ;
 wire \proj_14.net130 ;
 wire \proj_14.net131 ;
 wire \proj_14.net133 ;
 wire \proj_14.net134 ;
 wire \proj_14.net136 ;
 wire \proj_14.net137 ;
 wire \proj_14.net139 ;
 wire \proj_14.net14 ;
 wire \proj_14.net140 ;
 wire \proj_14.net142 ;
 wire \proj_14.net143 ;
 wire \proj_14.net145 ;
 wire \proj_14.net146 ;
 wire \proj_14.net148 ;
 wire \proj_14.net149 ;
 wire \proj_14.net15 ;
 wire \proj_14.net151 ;
 wire \proj_14.net152 ;
 wire \proj_14.net154 ;
 wire \proj_14.net155 ;
 wire \proj_14.net157 ;
 wire \proj_14.net158 ;
 wire \proj_14.net160 ;
 wire \proj_14.net161 ;
 wire \proj_14.net163 ;
 wire \proj_14.net164 ;
 wire \proj_14.net166 ;
 wire \proj_14.net167 ;
 wire \proj_14.net169 ;
 wire \proj_14.net17 ;
 wire \proj_14.net170 ;
 wire \proj_14.net172 ;
 wire \proj_14.net173 ;
 wire \proj_14.net175 ;
 wire \proj_14.net176 ;
 wire \proj_14.net178 ;
 wire \proj_14.net179 ;
 wire \proj_14.net18 ;
 wire \proj_14.net181 ;
 wire \proj_14.net182 ;
 wire \proj_14.net184 ;
 wire \proj_14.net185 ;
 wire \proj_14.net187 ;
 wire \proj_14.net188 ;
 wire \proj_14.net190 ;
 wire \proj_14.net192 ;
 wire \proj_14.net194 ;
 wire \proj_14.net195 ;
 wire \proj_14.net197 ;
 wire \proj_14.net198 ;
 wire \proj_14.net20 ;
 wire \proj_14.net200 ;
 wire \proj_14.net201 ;
 wire \proj_14.net203 ;
 wire \proj_14.net204 ;
 wire \proj_14.net206 ;
 wire \proj_14.net207 ;
 wire \proj_14.net209 ;
 wire \proj_14.net21 ;
 wire \proj_14.net210 ;
 wire \proj_14.net212 ;
 wire \proj_14.net213 ;
 wire \proj_14.net215 ;
 wire \proj_14.net216 ;
 wire \proj_14.net218 ;
 wire \proj_14.net219 ;
 wire \proj_14.net221 ;
 wire \proj_14.net222 ;
 wire \proj_14.net224 ;
 wire \proj_14.net225 ;
 wire \proj_14.net227 ;
 wire \proj_14.net228 ;
 wire \proj_14.net23 ;
 wire \proj_14.net230 ;
 wire \proj_14.net231 ;
 wire \proj_14.net233 ;
 wire \proj_14.net234 ;
 wire \proj_14.net236 ;
 wire \proj_14.net237 ;
 wire \proj_14.net239 ;
 wire \proj_14.net24 ;
 wire \proj_14.net240 ;
 wire \proj_14.net242 ;
 wire \proj_14.net243 ;
 wire \proj_14.net245 ;
 wire \proj_14.net246 ;
 wire \proj_14.net248 ;
 wire \proj_14.net249 ;
 wire \proj_14.net251 ;
 wire \proj_14.net252 ;
 wire \proj_14.net254 ;
 wire \proj_14.net256 ;
 wire \proj_14.net258 ;
 wire \proj_14.net259 ;
 wire \proj_14.net26 ;
 wire \proj_14.net261 ;
 wire \proj_14.net262 ;
 wire \proj_14.net264 ;
 wire \proj_14.net265 ;
 wire \proj_14.net267 ;
 wire \proj_14.net268 ;
 wire \proj_14.net27 ;
 wire \proj_14.net270 ;
 wire \proj_14.net271 ;
 wire \proj_14.net273 ;
 wire \proj_14.net274 ;
 wire \proj_14.net276 ;
 wire \proj_14.net277 ;
 wire \proj_14.net279 ;
 wire \proj_14.net280 ;
 wire \proj_14.net282 ;
 wire \proj_14.net283 ;
 wire \proj_14.net285 ;
 wire \proj_14.net286 ;
 wire \proj_14.net288 ;
 wire \proj_14.net289 ;
 wire \proj_14.net29 ;
 wire \proj_14.net291 ;
 wire \proj_14.net292 ;
 wire \proj_14.net294 ;
 wire \proj_14.net295 ;
 wire \proj_14.net297 ;
 wire \proj_14.net298 ;
 wire \proj_14.net30 ;
 wire \proj_14.net300 ;
 wire \proj_14.net301 ;
 wire \proj_14.net303 ;
 wire \proj_14.net304 ;
 wire \proj_14.net306 ;
 wire \proj_14.net307 ;
 wire \proj_14.net309 ;
 wire \proj_14.net310 ;
 wire \proj_14.net312 ;
 wire \proj_14.net313 ;
 wire \proj_14.net315 ;
 wire \proj_14.net316 ;
 wire \proj_14.net318 ;
 wire \proj_14.net32 ;
 wire \proj_14.net320 ;
 wire \proj_14.net322 ;
 wire \proj_14.net323 ;
 wire \proj_14.net325 ;
 wire \proj_14.net326 ;
 wire \proj_14.net328 ;
 wire \proj_14.net329 ;
 wire \proj_14.net33 ;
 wire \proj_14.net332 ;
 wire \proj_14.net333 ;
 wire \proj_14.net335 ;
 wire \proj_14.net336 ;
 wire \proj_14.net338 ;
 wire \proj_14.net339 ;
 wire \proj_14.net341 ;
 wire \proj_14.net342 ;
 wire \proj_14.net344 ;
 wire \proj_14.net345 ;
 wire \proj_14.net347 ;
 wire \proj_14.net348 ;
 wire \proj_14.net35 ;
 wire \proj_14.net350 ;
 wire \proj_14.net351 ;
 wire \proj_14.net353 ;
 wire \proj_14.net354 ;
 wire \proj_14.net356 ;
 wire \proj_14.net357 ;
 wire \proj_14.net359 ;
 wire \proj_14.net36 ;
 wire \proj_14.net360 ;
 wire \proj_14.net362 ;
 wire \proj_14.net363 ;
 wire \proj_14.net365 ;
 wire \proj_14.net366 ;
 wire \proj_14.net368 ;
 wire \proj_14.net369 ;
 wire \proj_14.net371 ;
 wire \proj_14.net372 ;
 wire \proj_14.net374 ;
 wire \proj_14.net375 ;
 wire \proj_14.net377 ;
 wire \proj_14.net378 ;
 wire \proj_14.net38 ;
 wire \proj_14.net380 ;
 wire \proj_14.net381 ;
 wire \proj_14.net383 ;
 wire \proj_14.net385 ;
 wire \proj_14.net387 ;
 wire \proj_14.net388 ;
 wire \proj_14.net39 ;
 wire \proj_14.net390 ;
 wire \proj_14.net391 ;
 wire \proj_14.net393 ;
 wire \proj_14.net394 ;
 wire \proj_14.net396 ;
 wire \proj_14.net397 ;
 wire \proj_14.net399 ;
 wire \proj_14.net4 ;
 wire \proj_14.net400 ;
 wire \proj_14.net402 ;
 wire \proj_14.net403 ;
 wire \proj_14.net405 ;
 wire \proj_14.net406 ;
 wire \proj_14.net408 ;
 wire \proj_14.net409 ;
 wire \proj_14.net41 ;
 wire \proj_14.net411 ;
 wire \proj_14.net412 ;
 wire \proj_14.net414 ;
 wire \proj_14.net415 ;
 wire \proj_14.net417 ;
 wire \proj_14.net418 ;
 wire \proj_14.net42 ;
 wire \proj_14.net420 ;
 wire \proj_14.net421 ;
 wire \proj_14.net423 ;
 wire \proj_14.net424 ;
 wire \proj_14.net426 ;
 wire \proj_14.net427 ;
 wire \proj_14.net429 ;
 wire \proj_14.net430 ;
 wire \proj_14.net432 ;
 wire \proj_14.net433 ;
 wire \proj_14.net435 ;
 wire \proj_14.net436 ;
 wire \proj_14.net438 ;
 wire \proj_14.net439 ;
 wire \proj_14.net44 ;
 wire \proj_14.net441 ;
 wire \proj_14.net442 ;
 wire \proj_14.net444 ;
 wire \proj_14.net445 ;
 wire \proj_14.net447 ;
 wire \proj_14.net449 ;
 wire \proj_14.net45 ;
 wire \proj_14.net451 ;
 wire \proj_14.net452 ;
 wire \proj_14.net454 ;
 wire \proj_14.net455 ;
 wire \proj_14.net457 ;
 wire \proj_14.net458 ;
 wire \proj_14.net460 ;
 wire \proj_14.net461 ;
 wire \proj_14.net463 ;
 wire \proj_14.net464 ;
 wire \proj_14.net466 ;
 wire \proj_14.net467 ;
 wire \proj_14.net469 ;
 wire \proj_14.net47 ;
 wire \proj_14.net470 ;
 wire \proj_14.net472 ;
 wire \proj_14.net473 ;
 wire \proj_14.net475 ;
 wire \proj_14.net476 ;
 wire \proj_14.net478 ;
 wire \proj_14.net479 ;
 wire \proj_14.net48 ;
 wire \proj_14.net481 ;
 wire \proj_14.net482 ;
 wire \proj_14.net484 ;
 wire \proj_14.net485 ;
 wire \proj_14.net487 ;
 wire \proj_14.net488 ;
 wire \proj_14.net490 ;
 wire \proj_14.net491 ;
 wire \proj_14.net493 ;
 wire \proj_14.net494 ;
 wire \proj_14.net496 ;
 wire \proj_14.net497 ;
 wire \proj_14.net499 ;
 wire \proj_14.net50 ;
 wire \proj_14.net500 ;
 wire \proj_14.net502 ;
 wire \proj_14.net503 ;
 wire \proj_14.net505 ;
 wire \proj_14.net506 ;
 wire \proj_14.net508 ;
 wire \proj_14.net509 ;
 wire \proj_14.net51 ;
 wire \proj_14.net512 ;
 wire \proj_14.net514 ;
 wire \proj_14.net515 ;
 wire \proj_14.net517 ;
 wire \proj_14.net518 ;
 wire \proj_14.net520 ;
 wire \proj_14.net521 ;
 wire \proj_14.net53 ;
 wire \proj_14.net54 ;
 wire \proj_14.net56 ;
 wire \proj_14.net57 ;
 wire \proj_14.net59 ;
 wire \proj_14.net63 ;
 wire \proj_14.net64 ;
 wire \proj_14.net66 ;
 wire \proj_14.net67 ;
 wire \proj_14.net69 ;
 wire \proj_14.net70 ;
 wire \proj_14.net72 ;
 wire \proj_14.net73 ;
 wire \proj_14.net75 ;
 wire \proj_14.net76 ;
 wire \proj_14.net78 ;
 wire \proj_14.net79 ;
 wire \proj_14.net8 ;
 wire \proj_14.net81 ;
 wire \proj_14.net82 ;
 wire \proj_14.net84 ;
 wire \proj_14.net85 ;
 wire \proj_14.net87 ;
 wire \proj_14.net88 ;
 wire \proj_14.net9 ;
 wire \proj_14.net90 ;
 wire \proj_14.net91 ;
 wire \proj_14.net93 ;
 wire \proj_14.net94 ;
 wire \proj_14.net96 ;
 wire \proj_14.net97 ;
 wire \proj_14.net99 ;
 wire \proj_15.net10 ;
 wire \proj_15.net11 ;
 wire \proj_15.net12 ;
 wire \proj_15.net13 ;
 wire \proj_15.net14 ;
 wire \proj_15.net15 ;
 wire \proj_15.net16 ;
 wire \proj_15.net9 ;
 wire \proj__0.net10 ;
 wire \proj__0.net11 ;
 wire \proj__0.net3 ;
 wire \proj__0.net4 ;
 wire \proj__1.net10 ;
 wire \proj__1.net11 ;
 wire \proj__1.net9 ;
 wire \proj__2.net14 ;
 wire \proj__2.net3 ;
 wire \proj__2.net5 ;
 wire \proj__2.net6 ;
 wire \proj__2.net7 ;
 wire \proj__3.net10 ;
 wire \proj__3.net11 ;
 wire \proj__3.net12 ;
 wire \proj__3.net13 ;
 wire \proj__3.net3 ;
 wire \proj__3.net4 ;
 wire \proj__4.net10 ;
 wire \proj__4.net11 ;
 wire \proj__4.net12 ;
 wire \proj__4.net9 ;
 wire \proj__5.net8 ;
 wire \proj__5.net9 ;
 wire \proj__6.net3 ;
 wire \proj__6.net4 ;
 wire \proj__7.net3 ;
 wire \proj__8.net10 ;
 wire \proj__8.net11 ;
 wire \proj__8.net12 ;
 wire \proj__8.net18 ;
 wire \proj__8.net19 ;
 wire \proj__8.net20 ;
 wire \proj__8.net7 ;
 wire \proj__8.net8 ;
 wire \proj__8.net9 ;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net245;
 wire \proj_10.flop1/notq ;
 wire net246;
 wire \proj_10.flop10/notq ;
 wire net247;
 wire \proj_10.flop11/notq ;
 wire net248;
 wire \proj_10.flop12/notq ;
 wire net249;
 wire \proj_10.flop13/notq ;
 wire net250;
 wire \proj_10.flop14/notq ;
 wire net251;
 wire \proj_10.flop2/notq ;
 wire net252;
 wire \proj_10.flop3/notq ;
 wire net253;
 wire \proj_10.flop4/notq ;
 wire net254;
 wire \proj_10.flop5/notq ;
 wire net255;
 wire \proj_10.flop6/notq ;
 wire net256;
 wire \proj_10.flop7/notq ;
 wire net257;
 wire \proj_10.flop8/notq ;
 wire net258;
 wire \proj_10.flop9/notq ;
 wire net259;
 wire \proj_14.flop1/notq ;
 wire net260;
 wire \proj_14.flop10/notq ;
 wire net261;
 wire \proj_14.flop100/notq ;
 wire net262;
 wire \proj_14.flop101/notq ;
 wire net263;
 wire \proj_14.flop102/notq ;
 wire net264;
 wire \proj_14.flop103/notq ;
 wire net265;
 wire \proj_14.flop104/notq ;
 wire net266;
 wire \proj_14.flop105/notq ;
 wire net267;
 wire \proj_14.flop106/notq ;
 wire net268;
 wire \proj_14.flop107/notq ;
 wire net269;
 wire \proj_14.flop108/notq ;
 wire net270;
 wire \proj_14.flop109/notq ;
 wire net271;
 wire \proj_14.flop11/notq ;
 wire net272;
 wire \proj_14.flop110/notq ;
 wire net273;
 wire \proj_14.flop111/notq ;
 wire net274;
 wire \proj_14.flop112/notq ;
 wire net275;
 wire \proj_14.flop113/notq ;
 wire net276;
 wire \proj_14.flop114/notq ;
 wire net277;
 wire \proj_14.flop115/notq ;
 wire net278;
 wire \proj_14.flop116/notq ;
 wire net279;
 wire \proj_14.flop117/notq ;
 wire net280;
 wire \proj_14.flop118/notq ;
 wire net281;
 wire \proj_14.flop119/notq ;
 wire net282;
 wire \proj_14.flop12/notq ;
 wire net283;
 wire \proj_14.flop120/notq ;
 wire net284;
 wire \proj_14.flop121/notq ;
 wire net285;
 wire \proj_14.flop122/notq ;
 wire net286;
 wire \proj_14.flop123/notq ;
 wire net287;
 wire \proj_14.flop124/notq ;
 wire net288;
 wire \proj_14.flop125/notq ;
 wire net289;
 wire \proj_14.flop126/notq ;
 wire net290;
 wire \proj_14.flop127/notq ;
 wire net291;
 wire \proj_14.flop128/notq ;
 wire net292;
 wire \proj_14.flop129/notq ;
 wire net293;
 wire \proj_14.flop13/notq ;
 wire net294;
 wire \proj_14.flop130/notq ;
 wire net295;
 wire \proj_14.flop131/notq ;
 wire net296;
 wire \proj_14.flop132/notq ;
 wire net297;
 wire \proj_14.flop133/notq ;
 wire net298;
 wire \proj_14.flop134/notq ;
 wire net299;
 wire \proj_14.flop135/notq ;
 wire net300;
 wire \proj_14.flop136/notq ;
 wire net301;
 wire \proj_14.flop137/notq ;
 wire net302;
 wire \proj_14.flop138/notq ;
 wire net303;
 wire \proj_14.flop139/notq ;
 wire net304;
 wire \proj_14.flop14/notq ;
 wire net305;
 wire \proj_14.flop140/notq ;
 wire net306;
 wire \proj_14.flop141/notq ;
 wire net307;
 wire \proj_14.flop142/notq ;
 wire net308;
 wire \proj_14.flop143/notq ;
 wire net309;
 wire \proj_14.flop144/notq ;
 wire net310;
 wire \proj_14.flop145/notq ;
 wire net311;
 wire \proj_14.flop146/notq ;
 wire net312;
 wire \proj_14.flop147/notq ;
 wire net313;
 wire \proj_14.flop148/notq ;
 wire net314;
 wire \proj_14.flop149/notq ;
 wire net315;
 wire \proj_14.flop15/notq ;
 wire net316;
 wire \proj_14.flop150/notq ;
 wire net317;
 wire \proj_14.flop151/notq ;
 wire net318;
 wire \proj_14.flop152/notq ;
 wire net319;
 wire \proj_14.flop153/notq ;
 wire net320;
 wire \proj_14.flop154/notq ;
 wire net321;
 wire \proj_14.flop155/notq ;
 wire net322;
 wire \proj_14.flop156/notq ;
 wire net323;
 wire \proj_14.flop157/notq ;
 wire net324;
 wire \proj_14.flop158/notq ;
 wire net325;
 wire \proj_14.flop159/notq ;
 wire net326;
 wire \proj_14.flop16/notq ;
 wire net327;
 wire \proj_14.flop160/notq ;
 wire net328;
 wire \proj_14.flop161/notq ;
 wire net329;
 wire \proj_14.flop162/notq ;
 wire net330;
 wire \proj_14.flop163/notq ;
 wire net331;
 wire \proj_14.flop164/notq ;
 wire net332;
 wire \proj_14.flop165/notq ;
 wire net333;
 wire \proj_14.flop166/notq ;
 wire net334;
 wire \proj_14.flop167/notq ;
 wire net335;
 wire \proj_14.flop168/notq ;
 wire net336;
 wire \proj_14.flop17/notq ;
 wire net337;
 wire \proj_14.flop18/notq ;
 wire net338;
 wire \proj_14.flop19/notq ;
 wire net339;
 wire \proj_14.flop2/notq ;
 wire net340;
 wire \proj_14.flop20/notq ;
 wire net341;
 wire \proj_14.flop21/notq ;
 wire net342;
 wire \proj_14.flop22/notq ;
 wire net343;
 wire \proj_14.flop23/notq ;
 wire net344;
 wire \proj_14.flop24/notq ;
 wire net345;
 wire \proj_14.flop25/notq ;
 wire net346;
 wire \proj_14.flop26/notq ;
 wire net347;
 wire \proj_14.flop27/notq ;
 wire net348;
 wire \proj_14.flop28/notq ;
 wire net349;
 wire \proj_14.flop29/notq ;
 wire net350;
 wire \proj_14.flop3/notq ;
 wire net351;
 wire \proj_14.flop30/notq ;
 wire net352;
 wire \proj_14.flop31/notq ;
 wire net353;
 wire \proj_14.flop32/notq ;
 wire net354;
 wire \proj_14.flop33/notq ;
 wire net355;
 wire \proj_14.flop34/notq ;
 wire net356;
 wire \proj_14.flop35/notq ;
 wire net357;
 wire \proj_14.flop36/notq ;
 wire net358;
 wire \proj_14.flop37/notq ;
 wire net359;
 wire \proj_14.flop38/notq ;
 wire net360;
 wire \proj_14.flop39/notq ;
 wire net361;
 wire \proj_14.flop4/notq ;
 wire net362;
 wire \proj_14.flop40/notq ;
 wire net363;
 wire \proj_14.flop41/notq ;
 wire net364;
 wire \proj_14.flop42/notq ;
 wire net365;
 wire \proj_14.flop43/notq ;
 wire net366;
 wire \proj_14.flop44/notq ;
 wire net367;
 wire \proj_14.flop45/notq ;
 wire net368;
 wire \proj_14.flop46/notq ;
 wire net369;
 wire \proj_14.flop47/notq ;
 wire net370;
 wire \proj_14.flop48/notq ;
 wire net371;
 wire \proj_14.flop49/notq ;
 wire net372;
 wire \proj_14.flop5/notq ;
 wire net373;
 wire \proj_14.flop50/notq ;
 wire net374;
 wire \proj_14.flop51/notq ;
 wire net375;
 wire \proj_14.flop52/notq ;
 wire net376;
 wire \proj_14.flop53/notq ;
 wire net377;
 wire \proj_14.flop54/notq ;
 wire net378;
 wire \proj_14.flop55/notq ;
 wire net379;
 wire \proj_14.flop56/notq ;
 wire net380;
 wire \proj_14.flop57/notq ;
 wire net381;
 wire \proj_14.flop58/notq ;
 wire net382;
 wire \proj_14.flop59/notq ;
 wire net383;
 wire \proj_14.flop6/notq ;
 wire net384;
 wire \proj_14.flop60/notq ;
 wire net385;
 wire \proj_14.flop61/notq ;
 wire net386;
 wire \proj_14.flop62/notq ;
 wire net387;
 wire \proj_14.flop63/notq ;
 wire net388;
 wire \proj_14.flop64/notq ;
 wire net389;
 wire \proj_14.flop65/notq ;
 wire net390;
 wire \proj_14.flop66/notq ;
 wire net391;
 wire \proj_14.flop67/notq ;
 wire net392;
 wire \proj_14.flop68/notq ;
 wire net393;
 wire \proj_14.flop69/notq ;
 wire net394;
 wire \proj_14.flop7/notq ;
 wire net395;
 wire \proj_14.flop70/notq ;
 wire net396;
 wire \proj_14.flop71/notq ;
 wire net397;
 wire \proj_14.flop72/notq ;
 wire net398;
 wire \proj_14.flop73/notq ;
 wire net399;
 wire \proj_14.flop74/notq ;
 wire net400;
 wire \proj_14.flop75/notq ;
 wire net401;
 wire \proj_14.flop76/notq ;
 wire net402;
 wire \proj_14.flop77/notq ;
 wire net403;
 wire \proj_14.flop78/notq ;
 wire net404;
 wire \proj_14.flop79/notq ;
 wire net405;
 wire \proj_14.flop8/notq ;
 wire net406;
 wire \proj_14.flop80/notq ;
 wire net407;
 wire \proj_14.flop81/notq ;
 wire net408;
 wire \proj_14.flop82/notq ;
 wire net409;
 wire \proj_14.flop83/notq ;
 wire net410;
 wire \proj_14.flop84/notq ;
 wire net411;
 wire \proj_14.flop85/notq ;
 wire net412;
 wire \proj_14.flop86/notq ;
 wire net413;
 wire \proj_14.flop87/notq ;
 wire net414;
 wire \proj_14.flop88/notq ;
 wire net415;
 wire \proj_14.flop89/notq ;
 wire net416;
 wire \proj_14.flop9/notq ;
 wire net417;
 wire \proj_14.flop90/notq ;
 wire net418;
 wire \proj_14.flop91/notq ;
 wire net419;
 wire \proj_14.flop92/notq ;
 wire net420;
 wire \proj_14.flop93/notq ;
 wire net421;
 wire \proj_14.flop94/notq ;
 wire net422;
 wire \proj_14.flop95/notq ;
 wire net423;
 wire \proj_14.flop96/notq ;
 wire net424;
 wire \proj_14.flop97/notq ;
 wire net425;
 wire \proj_14.flop98/notq ;
 wire net426;
 wire \proj_14.flop99/notq ;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;
 wire clknet_0_clk_regs;
 wire clknet_4_0_0_clk_regs;
 wire clknet_4_1_0_clk_regs;
 wire clknet_4_2_0_clk_regs;
 wire clknet_4_3_0_clk_regs;
 wire clknet_4_4_0_clk_regs;
 wire clknet_4_5_0_clk_regs;
 wire clknet_4_6_0_clk_regs;
 wire clknet_4_7_0_clk_regs;
 wire clknet_4_8_0_clk_regs;
 wire clknet_4_9_0_clk_regs;
 wire clknet_4_10_0_clk_regs;
 wire clknet_4_11_0_clk_regs;
 wire clknet_4_12_0_clk_regs;
 wire clknet_4_13_0_clk_regs;
 wire clknet_4_14_0_clk_regs;
 wire clknet_4_15_0_clk_regs;
 wire clknet_5_0__leaf_clk_regs;
 wire clknet_5_1__leaf_clk_regs;
 wire clknet_5_2__leaf_clk_regs;
 wire clknet_5_3__leaf_clk_regs;
 wire clknet_5_4__leaf_clk_regs;
 wire clknet_5_5__leaf_clk_regs;
 wire clknet_5_6__leaf_clk_regs;
 wire clknet_5_7__leaf_clk_regs;
 wire clknet_5_8__leaf_clk_regs;
 wire clknet_5_9__leaf_clk_regs;
 wire clknet_5_10__leaf_clk_regs;
 wire clknet_5_11__leaf_clk_regs;
 wire clknet_5_12__leaf_clk_regs;
 wire clknet_5_13__leaf_clk_regs;
 wire clknet_5_14__leaf_clk_regs;
 wire clknet_5_15__leaf_clk_regs;
 wire clknet_5_16__leaf_clk_regs;
 wire clknet_5_17__leaf_clk_regs;
 wire clknet_5_18__leaf_clk_regs;
 wire clknet_5_19__leaf_clk_regs;
 wire clknet_5_20__leaf_clk_regs;
 wire clknet_5_21__leaf_clk_regs;
 wire clknet_5_22__leaf_clk_regs;
 wire clknet_5_23__leaf_clk_regs;
 wire clknet_5_24__leaf_clk_regs;
 wire clknet_5_25__leaf_clk_regs;
 wire clknet_5_26__leaf_clk_regs;
 wire clknet_5_27__leaf_clk_regs;
 wire clknet_5_28__leaf_clk_regs;
 wire clknet_5_29__leaf_clk_regs;
 wire clknet_5_30__leaf_clk_regs;
 wire clknet_5_31__leaf_clk_regs;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;

 sg13g2_inv_1 _239_ (.Y(_048_),
    .A(\proj__0.net3 ));
 sg13g2_inv_1 _240_ (.Y(_049_),
    .A(\proj__0.net4 ));
 sg13g2_nor2_2 _241_ (.A(net11),
    .B(net12),
    .Y(_050_));
 sg13g2_nand2b_1 _242_ (.Y(_051_),
    .B(_050_),
    .A_N(net135));
 sg13g2_nor2_1 _243_ (.A(net135),
    .B(net10),
    .Y(_052_));
 sg13g2_and2_1 _244_ (.A(_050_),
    .B(_052_),
    .X(_053_));
 sg13g2_nor2b_2 _245_ (.A(net12),
    .B_N(net11),
    .Y(_054_));
 sg13g2_nand3_1 _246_ (.B(net179),
    .C(_054_),
    .A(net9),
    .Y(_055_));
 sg13g2_and2_1 _247_ (.A(net11),
    .B(net12),
    .X(_056_));
 sg13g2_and2_2 _248_ (.A(_052_),
    .B(_056_),
    .X(_057_));
 sg13g2_nor2b_1 _249_ (.A(net10),
    .B_N(net135),
    .Y(_058_));
 sg13g2_and2_2 _250_ (.A(_050_),
    .B(_058_),
    .X(_059_));
 sg13g2_nand2_1 _251_ (.Y(_060_),
    .A(\proj__1.net9 ),
    .B(_059_));
 sg13g2_nor2b_1 _252_ (.A(net135),
    .B_N(net10),
    .Y(_061_));
 sg13g2_and2_1 _253_ (.A(_054_),
    .B(_061_),
    .X(_062_));
 sg13g2_nand2_1 _254_ (.Y(_063_),
    .A(\proj__6.net3 ),
    .B(_062_));
 sg13g2_nor2b_1 _255_ (.A(net11),
    .B_N(net12),
    .Y(_064_));
 sg13g2_and2_2 _256_ (.A(_061_),
    .B(_064_),
    .X(_065_));
 sg13g2_and2_2 _257_ (.A(_050_),
    .B(_061_),
    .X(_066_));
 sg13g2_nand2_1 _258_ (.Y(_067_),
    .A(\proj__2.net3 ),
    .B(_066_));
 sg13g2_and2_2 _259_ (.A(_052_),
    .B(_054_),
    .X(_068_));
 sg13g2_and2_1 _260_ (.A(_056_),
    .B(_061_),
    .X(_069_));
 sg13g2_and3_2 _261_ (.X(_000_),
    .A(net135),
    .B(net10),
    .C(_064_));
 sg13g2_and2_2 _262_ (.A(_056_),
    .B(_058_),
    .X(_001_));
 sg13g2_and3_2 _263_ (.X(_002_),
    .A(net135),
    .B(net10),
    .C(_056_));
 sg13g2_and2_2 _264_ (.A(_052_),
    .B(_064_),
    .X(_003_));
 sg13g2_a22oi_1 _265_ (.Y(_004_),
    .B1(_000_),
    .B2(\proj_11.net9 ),
    .A2(_057_),
    .A1(net426));
 sg13g2_a22oi_1 _266_ (.Y(_005_),
    .B1(_002_),
    .B2(\proj_15.net9 ),
    .A2(_068_),
    .A1(\proj__4.net9 ));
 sg13g2_and4_1 _267_ (.A(_055_),
    .B(_063_),
    .C(_004_),
    .D(_005_),
    .X(_006_));
 sg13g2_a221oi_1 _268_ (.B2(\proj__8.net7 ),
    .C1(_053_),
    .B1(_003_),
    .A1(\proj_10.net10 ),
    .Y(_007_),
    .A2(_065_));
 sg13g2_a22oi_1 _269_ (.Y(_008_),
    .B1(_001_),
    .B2(\proj_13.net9 ),
    .A2(_069_),
    .A1(net8));
 sg13g2_and4_1 _270_ (.A(_060_),
    .B(_067_),
    .C(_007_),
    .D(_008_),
    .X(_009_));
 sg13g2_a22oi_1 _271_ (.Y(uo_out[0]),
    .B1(_006_),
    .B2(_009_),
    .A2(_053_),
    .A1(_048_));
 sg13g2_a22oi_1 _272_ (.Y(_010_),
    .B1(_000_),
    .B2(\proj_11.net10 ),
    .A2(_062_),
    .A1(\proj__6.net4 ));
 sg13g2_a22oi_1 _273_ (.Y(_011_),
    .B1(_002_),
    .B2(\proj_15.net10 ),
    .A2(_065_),
    .A1(\proj_10.net11 ));
 sg13g2_and4_1 _274_ (.A(_051_),
    .B(_060_),
    .C(_010_),
    .D(_011_),
    .X(_012_));
 sg13g2_and3_1 _275_ (.X(_013_),
    .A(net135),
    .B(net10),
    .C(_050_));
 sg13g2_a22oi_1 _276_ (.Y(_014_),
    .B1(_013_),
    .B2(\proj__3.net3 ),
    .A2(_057_),
    .A1(\proj_12.net12 ));
 sg13g2_a22oi_1 _277_ (.Y(_015_),
    .B1(_003_),
    .B2(\proj__8.net8 ),
    .A2(_001_),
    .A1(\proj_13.net10 ));
 sg13g2_a22oi_1 _278_ (.Y(_016_),
    .B1(_069_),
    .B2(net167),
    .A2(_068_),
    .A1(\proj__4.net10 ));
 sg13g2_and3_1 _279_ (.X(_017_),
    .A(net135),
    .B(net10),
    .C(\proj__7.net3 ));
 sg13g2_and2_2 _280_ (.A(_054_),
    .B(_058_),
    .X(_018_));
 sg13g2_a22oi_1 _281_ (.Y(_019_),
    .B1(_018_),
    .B2(net3),
    .A2(_017_),
    .A1(_054_));
 sg13g2_and4_1 _282_ (.A(_014_),
    .B(_015_),
    .C(_016_),
    .D(_019_),
    .X(_020_));
 sg13g2_a22oi_1 _283_ (.Y(uo_out[1]),
    .B1(_012_),
    .B2(_020_),
    .A2(_053_),
    .A1(_049_));
 sg13g2_a22oi_1 _284_ (.Y(_021_),
    .B1(_059_),
    .B2(\proj__1.net10 ),
    .A2(_057_),
    .A1(\proj_12.net13 ));
 sg13g2_a22oi_1 _285_ (.Y(_022_),
    .B1(_000_),
    .B2(\proj_11.net11 ),
    .A2(_066_),
    .A1(\proj__2.net5 ));
 sg13g2_a22oi_1 _286_ (.Y(_023_),
    .B1(_003_),
    .B2(\proj__8.net8 ),
    .A2(_065_),
    .A1(\proj_10.net12 ));
 sg13g2_a22oi_1 _287_ (.Y(_024_),
    .B1(_002_),
    .B2(\proj_15.net11 ),
    .A2(_068_),
    .A1(\proj__4.net11 ));
 sg13g2_a22oi_1 _288_ (.Y(_025_),
    .B1(_018_),
    .B2(net174),
    .A2(_001_),
    .A1(\proj_13.net11 ));
 sg13g2_and3_1 _289_ (.X(_026_),
    .A(_023_),
    .B(_024_),
    .C(_025_));
 sg13g2_nand3_1 _290_ (.B(_022_),
    .C(_026_),
    .A(_021_),
    .Y(uo_out[2]));
 sg13g2_a22oi_1 _291_ (.Y(_027_),
    .B1(_003_),
    .B2(\proj__8.net9 ),
    .A2(_068_),
    .A1(\proj__4.net12 ));
 sg13g2_a22oi_1 _292_ (.Y(_028_),
    .B1(_001_),
    .B2(\proj_13.net12 ),
    .A2(_000_),
    .A1(\proj_11.net12 ));
 sg13g2_and2_1 _293_ (.A(_027_),
    .B(_028_),
    .X(_029_));
 sg13g2_a22oi_1 _294_ (.Y(_030_),
    .B1(_018_),
    .B2(\proj__5.net8 ),
    .A2(_066_),
    .A1(\proj__2.net3 ));
 sg13g2_a22oi_1 _295_ (.Y(_031_),
    .B1(_065_),
    .B2(\proj_10.net13 ),
    .A2(_057_),
    .A1(\proj_12.net14 ));
 sg13g2_a22oi_1 _296_ (.Y(_032_),
    .B1(_002_),
    .B2(\proj_15.net12 ),
    .A2(_059_),
    .A1(\proj__1.net11 ));
 sg13g2_nand4_1 _297_ (.B(_030_),
    .C(_031_),
    .A(_029_),
    .Y(uo_out[3]),
    .D(_032_));
 sg13g2_a22oi_1 _298_ (.Y(_033_),
    .B1(_002_),
    .B2(\proj_15.net13 ),
    .A2(_000_),
    .A1(\proj_11.net13 ));
 sg13g2_a22oi_1 _299_ (.Y(_034_),
    .B1(_003_),
    .B2(\proj__8.net10 ),
    .A2(_065_),
    .A1(\proj_10.net14 ));
 sg13g2_or2_1 _300_ (.X(_035_),
    .B(_068_),
    .A(_059_));
 sg13g2_nand2_1 _301_ (.Y(_036_),
    .A(net172),
    .B(_035_));
 sg13g2_nand4_1 _302_ (.B(_033_),
    .C(_034_),
    .A(_030_),
    .Y(uo_out[4]),
    .D(_036_));
 sg13g2_o21ai_1 _303_ (.B1(net171),
    .Y(_037_),
    .A1(_018_),
    .A2(_035_));
 sg13g2_a22oi_1 _304_ (.Y(_038_),
    .B1(_002_),
    .B2(\proj_15.net14 ),
    .A2(_065_),
    .A1(\proj_10.net15 ));
 sg13g2_a22oi_1 _305_ (.Y(_039_),
    .B1(_013_),
    .B2(\proj__3.net4 ),
    .A2(_001_),
    .A1(\proj_13.net13 ));
 sg13g2_a22oi_1 _306_ (.Y(_040_),
    .B1(_003_),
    .B2(\proj__8.net11 ),
    .A2(_066_),
    .A1(\proj__2.net6 ));
 sg13g2_nand4_1 _307_ (.B(_038_),
    .C(_039_),
    .A(_037_),
    .Y(uo_out[5]),
    .D(_040_));
 sg13g2_a22oi_1 _308_ (.Y(_041_),
    .B1(_018_),
    .B2(\proj__5.net9 ),
    .A2(_066_),
    .A1(\proj__2.net7 ));
 sg13g2_a22oi_1 _309_ (.Y(_042_),
    .B1(_003_),
    .B2(\proj__8.net12 ),
    .A2(_065_),
    .A1(\proj_10.net16 ));
 sg13g2_nand2_1 _310_ (.Y(_043_),
    .A(net164),
    .B(_035_));
 sg13g2_a22oi_1 _311_ (.Y(_044_),
    .B1(_002_),
    .B2(\proj_15.net15 ),
    .A2(_001_),
    .A1(\proj_13.net12 ));
 sg13g2_nand4_1 _312_ (.B(_042_),
    .C(_043_),
    .A(_041_),
    .Y(uo_out[6]),
    .D(_044_));
 sg13g2_nand2_1 _313_ (.Y(_045_),
    .A(net136),
    .B(_035_));
 sg13g2_a22oi_1 _314_ (.Y(_046_),
    .B1(_002_),
    .B2(\proj_15.net16 ),
    .A2(_065_),
    .A1(\proj_10.net17 ));
 sg13g2_a22oi_1 _315_ (.Y(_047_),
    .B1(_001_),
    .B2(\proj_13.net14 ),
    .A2(_069_),
    .A1(\proj_14.net4 ));
 sg13g2_nand3_1 _316_ (.B(_046_),
    .C(_047_),
    .A(_045_),
    .Y(uo_out[7]));
 sg13g2_tiehi \proj_14.mux100/_0__78  (.L_HI(net78));
 sg13g2_tiehi \proj_14.mux101/_0__79  (.L_HI(net79));
 sg13g2_tiehi \proj_14.mux102/_0__80  (.L_HI(net80));
 sg13g2_tiehi \proj_14.mux103/_0__81  (.L_HI(net81));
 sg13g2_tiehi \proj_14.mux104/_0__82  (.L_HI(net82));
 sg13g2_tiehi \proj_14.mux105/_0__83  (.L_HI(net83));
 sg13g2_tiehi \proj_14.mux106/_0__84  (.L_HI(net84));
 sg13g2_tiehi \proj_14.mux107/_0__85  (.L_HI(net85));
 sg13g2_tiehi \proj_14.mux108/_0__86  (.L_HI(net86));
 sg13g2_tiehi \proj_14.mux109/_0__87  (.L_HI(net87));
 sg13g2_tiehi \proj_14.mux11/_0__88  (.L_HI(net88));
 sg13g2_tiehi \proj_14.mux110/_0__89  (.L_HI(net89));
 sg13g2_tiehi \proj_14.mux112/_0__90  (.L_HI(net90));
 sg13g2_tiehi \proj_14.mux118/_0__91  (.L_HI(net91));
 sg13g2_tiehi \proj_14.mux120/_0__92  (.L_HI(net92));
 sg13g2_tiehi \proj_14.mux121/_0__93  (.L_HI(net93));
 sg13g2_tiehi \proj_14.mux122/_0__94  (.L_HI(net94));
 sg13g2_tiehi \proj_14.mux123/_0__95  (.L_HI(net95));
 sg13g2_tiehi \proj_14.mux124/_0__96  (.L_HI(net96));
 sg13g2_tiehi \proj_14.mux125/_0__97  (.L_HI(net97));
 sg13g2_tiehi \proj_14.mux126/_0__98  (.L_HI(net98));
 sg13g2_tiehi \proj_14.mux127/_0__99  (.L_HI(net99));
 sg13g2_tiehi \proj_14.mux128/_0__100  (.L_HI(net100));
 sg13g2_tiehi \proj_14.mux129/_0__101  (.L_HI(net101));
 sg13g2_tiehi \proj_14.mux13/_0__102  (.L_HI(net102));
 sg13g2_tiehi \proj_14.mux130/_0__103  (.L_HI(net103));
 sg13g2_tiehi \proj_14.mux131/_0__104  (.L_HI(net104));
 sg13g2_tiehi \proj_14.mux133/_0__105  (.L_HI(net105));
 sg13g2_tiehi \proj_14.mux136/_0__106  (.L_HI(net106));
 sg13g2_tiehi \proj_14.mux139/_0__107  (.L_HI(net107));
 sg13g2_tiehi \proj_14.mux141/_0__108  (.L_HI(net108));
 sg13g2_tiehi \proj_14.mux142/_0__109  (.L_HI(net109));
 sg13g2_tiehi \proj_14.mux143/_0__110  (.L_HI(net110));
 sg13g2_tiehi \proj_14.mux144/_0__111  (.L_HI(net111));
 sg13g2_tiehi \proj_14.mux145/_0__112  (.L_HI(net112));
 sg13g2_tiehi \proj_14.mux146/_0__113  (.L_HI(net113));
 sg13g2_tiehi \proj_14.mux147/_0__114  (.L_HI(net114));
 sg13g2_tiehi \proj_14.mux148/_0__115  (.L_HI(net115));
 sg13g2_tiehi \proj_14.mux149/_0__116  (.L_HI(net116));
 sg13g2_tiehi \proj_14.mux15/_0__117  (.L_HI(net117));
 sg13g2_tiehi \proj_14.mux150/_0__118  (.L_HI(net118));
 sg13g2_tiehi \proj_14.mux151/_0__119  (.L_HI(net119));
 sg13g2_tiehi \proj_14.mux152/_0__120  (.L_HI(net120));
 sg13g2_tiehi \proj_14.mux155/_0__121  (.L_HI(net121));
 sg13g2_tiehi \proj_14.mux157/_0__122  (.L_HI(net122));
 sg13g2_tiehi \proj_14.mux16/_0__123  (.L_HI(net123));
 sg13g2_tiehi \proj_14.mux162/_0__124  (.L_HI(net124));
 sg13g2_tiehi \proj_14.mux163/_0__125  (.L_HI(net125));
 sg13g2_tiehi \proj_14.mux164/_0__126  (.L_HI(net126));
 sg13g2_tiehi \proj_14.mux165/_0__127  (.L_HI(net127));
 sg13g2_tiehi \proj_14.mux166/_0__128  (.L_HI(net128));
 sg13g2_tiehi \proj_14.mux167/_0__129  (.L_HI(net129));
 sg13g2_tiehi \proj_14.mux168/_0__130  (.L_HI(net130));
 sg13g2_tiehi \proj_14.mux169/_0__131  (.L_HI(net131));
 sg13g2_tiehi \proj_14.mux17/_0__132  (.L_HI(net132));
 sg13g2_tiehi \proj_14.mux18/_0__133  (.L_HI(net133));
 sg13g2_tiehi \proj_14.mux19/_0__134  (.L_HI(net134));
 sg13g2_tiehi \proj_14.mux2/_0__135  (.L_HI(net181));
 sg13g2_tiehi \proj_14.mux20/_0__136  (.L_HI(net182));
 sg13g2_tiehi \proj_14.mux21/_0__137  (.L_HI(net183));
 sg13g2_tiehi \proj_14.mux22/_0__138  (.L_HI(net184));
 sg13g2_tiehi \proj_14.mux27/_0__139  (.L_HI(net185));
 sg13g2_tiehi \proj_14.mux3/_0__140  (.L_HI(net186));
 sg13g2_tiehi \proj_14.mux30/_0__141  (.L_HI(net187));
 sg13g2_tiehi \proj_14.mux32/_0__142  (.L_HI(net188));
 sg13g2_tiehi \proj_14.mux33/_0__143  (.L_HI(net189));
 sg13g2_tiehi \proj_14.mux34/_0__144  (.L_HI(net190));
 sg13g2_tiehi \proj_14.mux35/_0__145  (.L_HI(net191));
 sg13g2_tiehi \proj_14.mux36/_0__146  (.L_HI(net192));
 sg13g2_tiehi \proj_14.mux37/_0__147  (.L_HI(net193));
 sg13g2_tiehi \proj_14.mux38/_0__148  (.L_HI(net194));
 sg13g2_tiehi \proj_14.mux39/_0__149  (.L_HI(net195));
 sg13g2_tiehi \proj_14.mux4/_0__150  (.L_HI(net196));
 sg13g2_tiehi \proj_14.mux40/_0__151  (.L_HI(net197));
 sg13g2_tiehi \proj_14.mux41/_0__152  (.L_HI(net198));
 sg13g2_tiehi \proj_14.mux42/_0__153  (.L_HI(net199));
 sg13g2_tiehi \proj_14.mux43/_0__154  (.L_HI(net200));
 sg13g2_tiehi \proj_14.mux44/_0__155  (.L_HI(net201));
 sg13g2_tiehi \proj_14.mux45/_0__156  (.L_HI(net202));
 sg13g2_tiehi \proj_14.mux46/_0__157  (.L_HI(net203));
 sg13g2_tiehi \proj_14.mux47/_0__158  (.L_HI(net204));
 sg13g2_tiehi \proj_14.mux49/_0__159  (.L_HI(net205));
 sg13g2_tiehi \proj_14.mux5/_0__160  (.L_HI(net206));
 sg13g2_tiehi \proj_14.mux55/_0__161  (.L_HI(net207));
 sg13g2_tiehi \proj_14.mux57/_0__162  (.L_HI(net208));
 sg13g2_tiehi \proj_14.mux58/_0__163  (.L_HI(net209));
 sg13g2_tiehi \proj_14.mux59/_0__164  (.L_HI(net210));
 sg13g2_tiehi \proj_14.mux60/_0__165  (.L_HI(net211));
 sg13g2_tiehi \proj_14.mux61/_0__166  (.L_HI(net212));
 sg13g2_tiehi \proj_14.mux62/_0__167  (.L_HI(net213));
 sg13g2_tiehi \proj_14.mux63/_0__168  (.L_HI(net214));
 sg13g2_tiehi \proj_14.mux64/_0__169  (.L_HI(net215));
 sg13g2_tiehi \proj_14.mux65/_0__170  (.L_HI(net216));
 sg13g2_tiehi \proj_14.mux66/_0__171  (.L_HI(net217));
 sg13g2_tiehi \proj_14.mux67/_0__172  (.L_HI(net218));
 sg13g2_tiehi \proj_14.mux68/_0__173  (.L_HI(net219));
 sg13g2_tiehi \proj_14.mux7/_0__174  (.L_HI(net220));
 sg13g2_tiehi \proj_14.mux70/_0__175  (.L_HI(net221));
 sg13g2_tiehi \proj_14.mux71/_0__176  (.L_HI(net222));
 sg13g2_tiehi \proj_14.mux72/_0__177  (.L_HI(net223));
 sg13g2_tiehi \proj_14.mux73/_0__178  (.L_HI(net224));
 sg13g2_tiehi \proj_14.mux76/_0__179  (.L_HI(net225));
 sg13g2_tiehi \proj_14.mux78/_0__180  (.L_HI(net226));
 sg13g2_tiehi \proj_14.mux79/_0__181  (.L_HI(net227));
 sg13g2_tiehi \proj_14.mux8/_0__182  (.L_HI(net228));
 sg13g2_tiehi \proj_14.mux80/_0__183  (.L_HI(net229));
 sg13g2_tiehi \proj_14.mux81/_0__184  (.L_HI(net230));
 sg13g2_tiehi \proj_14.mux82/_0__185  (.L_HI(net231));
 sg13g2_tiehi \proj_14.mux83/_0__186  (.L_HI(net232));
 sg13g2_tiehi \proj_14.mux84/_0__187  (.L_HI(net233));
 sg13g2_tiehi \proj_14.mux85/_0__188  (.L_HI(net234));
 sg13g2_tiehi \proj_14.mux86/_0__189  (.L_HI(net235));
 sg13g2_tiehi \proj_14.mux87/_0__190  (.L_HI(net236));
 sg13g2_tiehi \proj_14.mux88/_0__191  (.L_HI(net237));
 sg13g2_tiehi \proj_14.mux89/_0__192  (.L_HI(net238));
 sg13g2_tiehi \proj_14.mux91/_0__193  (.L_HI(net239));
 sg13g2_tiehi \proj_14.mux92/_0__194  (.L_HI(net240));
 sg13g2_tiehi \proj_14.mux94/_0__195  (.L_HI(net241));
 sg13g2_tiehi \proj_14.mux97/_0__196  (.L_HI(net242));
 sg13g2_tiehi \proj_14.mux99/_0__197  (.L_HI(net243));
 sg13g2_tiehi \proj_10.flop1/_1__198  (.L_HI(net244));
 sg13g2_tielo \proj_14.mux111/_0__14  (.L_LO(net14));
 sg13g2_tielo \proj_14.mux113/_0__15  (.L_LO(net15));
 sg13g2_tielo \proj_14.mux114/_0__16  (.L_LO(net16));
 sg13g2_tielo \proj_14.mux115/_0__17  (.L_LO(net17));
 sg13g2_tielo \proj_14.mux116/_0__18  (.L_LO(net18));
 sg13g2_tielo \proj_14.mux117/_0__19  (.L_LO(net19));
 sg13g2_tielo \proj_14.mux119/_0__20  (.L_LO(net20));
 sg13g2_tielo \proj_14.mux12/_0__21  (.L_LO(net21));
 sg13g2_tielo \proj_14.mux132/_0__22  (.L_LO(net22));
 sg13g2_tielo \proj_14.mux134/_0__23  (.L_LO(net23));
 sg13g2_tielo \proj_14.mux135/_0__24  (.L_LO(net24));
 sg13g2_tielo \proj_14.mux137/_0__25  (.L_LO(net25));
 sg13g2_tielo \proj_14.mux138/_0__26  (.L_LO(net26));
 sg13g2_tielo \proj_14.mux14/_0__27  (.L_LO(net27));
 sg13g2_tielo \proj_14.mux140/_0__28  (.L_LO(net28));
 sg13g2_tielo \proj_14.mux153/_0__29  (.L_LO(net29));
 sg13g2_tielo \proj_14.mux154/_0__30  (.L_LO(net30));
 sg13g2_tielo \proj_14.mux156/_0__31  (.L_LO(net31));
 sg13g2_tielo \proj_14.mux158/_0__32  (.L_LO(net32));
 sg13g2_tielo \proj_14.mux159/_0__33  (.L_LO(net33));
 sg13g2_tielo \proj_14.mux160/_0__34  (.L_LO(net34));
 sg13g2_tielo \proj_14.mux161/_0__35  (.L_LO(net35));
 sg13g2_tielo \proj_14.mux23/_0__36  (.L_LO(net36));
 sg13g2_tielo \proj_14.mux24/_0__37  (.L_LO(net37));
 sg13g2_tielo \proj_14.mux25/_0__38  (.L_LO(net38));
 sg13g2_tielo \proj_14.mux26/_0__39  (.L_LO(net39));
 sg13g2_tielo \proj_14.mux28/_0__40  (.L_LO(net40));
 sg13g2_tielo \proj_14.mux29/_0__41  (.L_LO(net41));
 sg13g2_tielo \proj_14.mux31/_0__42  (.L_LO(net42));
 sg13g2_tielo \proj_14.mux48/_0__43  (.L_LO(net43));
 sg13g2_tielo \proj_14.mux50/_0__44  (.L_LO(net44));
 sg13g2_tielo \proj_14.mux51/_0__45  (.L_LO(net45));
 sg13g2_tielo \proj_14.mux52/_0__46  (.L_LO(net46));
 sg13g2_tielo \proj_14.mux53/_0__47  (.L_LO(net47));
 sg13g2_tielo \proj_14.mux54/_0__48  (.L_LO(net48));
 sg13g2_tielo \proj_14.mux56/_0__49  (.L_LO(net49));
 sg13g2_tielo \proj_14.mux6/_0__50  (.L_LO(net50));
 sg13g2_tielo \proj_14.mux69/_0__51  (.L_LO(net51));
 sg13g2_tielo \proj_14.mux74/_0__52  (.L_LO(net52));
 sg13g2_tielo \proj_14.mux75/_0__53  (.L_LO(net53));
 sg13g2_tielo \proj_14.mux77/_0__54  (.L_LO(net54));
 sg13g2_tielo \proj_14.mux9/_0__55  (.L_LO(net55));
 sg13g2_tielo \proj_14.mux90/_0__56  (.L_LO(net56));
 sg13g2_tielo \proj_14.mux93/_0__57  (.L_LO(net57));
 sg13g2_tielo \proj_14.mux95/_0__58  (.L_LO(net58));
 sg13g2_tielo \proj_14.mux96/_0__59  (.L_LO(net59));
 sg13g2_tielo \proj_14.mux98/_0__60  (.L_LO(net60));
 sg13g2_tielo tt_um_wokwi_group_2_61 (.L_LO(net61));
 sg13g2_tielo tt_um_wokwi_group_2_62 (.L_LO(net62));
 sg13g2_tielo tt_um_wokwi_group_2_63 (.L_LO(net63));
 sg13g2_tielo tt_um_wokwi_group_2_64 (.L_LO(net64));
 sg13g2_tielo tt_um_wokwi_group_2_65 (.L_LO(net65));
 sg13g2_tielo tt_um_wokwi_group_2_66 (.L_LO(net66));
 sg13g2_tielo tt_um_wokwi_group_2_67 (.L_LO(net67));
 sg13g2_tielo tt_um_wokwi_group_2_68 (.L_LO(net68));
 sg13g2_tielo tt_um_wokwi_group_2_69 (.L_LO(net69));
 sg13g2_tielo tt_um_wokwi_group_2_70 (.L_LO(net70));
 sg13g2_tielo tt_um_wokwi_group_2_71 (.L_LO(net71));
 sg13g2_tielo tt_um_wokwi_group_2_72 (.L_LO(net72));
 sg13g2_tielo tt_um_wokwi_group_2_73 (.L_LO(net73));
 sg13g2_tielo tt_um_wokwi_group_2_74 (.L_LO(net74));
 sg13g2_tielo tt_um_wokwi_group_2_75 (.L_LO(net75));
 sg13g2_tielo tt_um_wokwi_group_2_76 (.L_LO(net76));
 sg13g2_tiehi \proj_14.mux1/_0__77  (.L_HI(net77));
 sg13g2_and2_1 \proj_10.and1/_0_  (.A(\proj_10.net37 ),
    .B(\proj_10.net28 ),
    .X(\proj_10.net41 ));
 sg13g2_and2_1 \proj_10.and10/_0_  (.A(\proj_10.net41 ),
    .B(net435),
    .X(\proj_10.net44 ));
 sg13g2_and2_1 \proj_10.and11/_0_  (.A(net428),
    .B(\proj_10.net43 ),
    .X(\proj_10.net46 ));
 sg13g2_and2_1 \proj_10.and2/_0_  (.A(\proj_10.net24 ),
    .B(\proj_10.net23 ),
    .X(\proj_10.net25 ));
 sg13g2_and2_1 \proj_10.and3/_0_  (.A(\proj_10.net27 ),
    .B(\proj_10.net26 ),
    .X(\proj_10.net28 ));
 sg13g2_and2_1 \proj_10.and4/_0_  (.A(\proj_10.net26 ),
    .B(net434),
    .X(\proj_10.net30 ));
 sg13g2_and2_1 \proj_10.and5/_0_  (.A(net436),
    .B(\proj_10.net23 ),
    .X(\proj_10.net32 ));
 sg13g2_and2_1 \proj_10.and6/_0_  (.A(\proj_10.net33 ),
    .B(\proj_10.net25 ),
    .X(\proj_10.net26 ));
 sg13g2_and2_1 \proj_10.and7/_0_  (.A(net432),
    .B(\proj_10.net25 ),
    .X(\proj_10.net35 ));
 sg13g2_and2_1 \proj_10.and8/_0_  (.A(\proj_10.net28 ),
    .B(net430),
    .X(\proj_10.net42 ));
 sg13g2_and2_1 \proj_10.and9/_0_  (.A(\proj_10.net41 ),
    .B(\proj_10.net39 ),
    .X(\proj_10.net43 ));
 sg13g2_dfrbp_1 \proj_10.flop1/_1_  (.CLK(clknet_5_27__leaf_clk_regs),
    .RESET_B(net244),
    .D(net180),
    .Q_N(\proj_10.flop1/notq ),
    .Q(\proj_10.net40 ));
 sg13g2_tiehi \proj_10.flop10/_1__199  (.L_HI(net245));
 sg13g2_dfrbp_1 \proj_10.flop10/_1_  (.CLK(clknet_5_12__leaf_clk_regs),
    .RESET_B(net245),
    .D(net171),
    .Q_N(\proj_10.flop10/notq ),
    .Q(\proj_10.net38 ));
 sg13g2_tiehi \proj_10.flop11/_1__200  (.L_HI(net246));
 sg13g2_dfrbp_1 \proj_10.flop11/_1_  (.CLK(clknet_5_12__leaf_clk_regs),
    .RESET_B(net246),
    .D(net172),
    .Q_N(\proj_10.flop11/notq ),
    .Q(\proj_10.net36 ));
 sg13g2_tiehi \proj_10.flop12/_1__201  (.L_HI(net247));
 sg13g2_dfrbp_1 \proj_10.flop12/_1_  (.CLK(clknet_5_13__leaf_clk_regs),
    .RESET_B(net247),
    .D(net429),
    .Q_N(\proj_10.flop12/notq ),
    .Q(\proj_10.net16 ));
 sg13g2_tiehi \proj_10.flop13/_1__202  (.L_HI(net248));
 sg13g2_dfrbp_1 \proj_10.flop13/_1_  (.CLK(clknet_5_13__leaf_clk_regs),
    .RESET_B(net248),
    .D(\proj_10.net44 ),
    .Q_N(\proj_10.flop13/notq ),
    .Q(\proj_10.net15 ));
 sg13g2_tiehi \proj_10.flop14/_1__203  (.L_HI(net249));
 sg13g2_dfrbp_1 \proj_10.flop14/_1_  (.CLK(clknet_5_14__leaf_clk_regs),
    .RESET_B(net249),
    .D(net431),
    .Q_N(\proj_10.flop14/notq ),
    .Q(\proj_10.net14 ));
 sg13g2_tiehi \proj_10.flop2/_1__204  (.L_HI(net250));
 sg13g2_dfrbp_1 \proj_10.flop2/_1_  (.CLK(clknet_5_15__leaf_clk_regs),
    .RESET_B(net250),
    .D(net173),
    .Q_N(\proj_10.flop2/notq ),
    .Q(\proj_10.net29 ));
 sg13g2_tiehi \proj_10.flop3/_1__205  (.L_HI(net251));
 sg13g2_dfrbp_1 \proj_10.flop3/_1_  (.CLK(clknet_5_26__leaf_clk_regs),
    .RESET_B(net251),
    .D(net174),
    .Q_N(\proj_10.flop3/notq ),
    .Q(\proj_10.net34 ));
 sg13g2_tiehi \proj_10.flop4/_1__206  (.L_HI(net252));
 sg13g2_dfrbp_1 \proj_10.flop4/_1_  (.CLK(clknet_5_26__leaf_clk_regs),
    .RESET_B(net252),
    .D(net176),
    .Q_N(\proj_10.flop4/notq ),
    .Q(\proj_10.net31 ));
 sg13g2_tiehi \proj_10.flop5/_1__207  (.L_HI(net253));
 sg13g2_dfrbp_1 \proj_10.flop5/_1_  (.CLK(clknet_5_15__leaf_clk_regs),
    .RESET_B(net253),
    .D(\proj_10.net30 ),
    .Q_N(\proj_10.flop5/notq ),
    .Q(\proj_10.net13 ));
 sg13g2_tiehi \proj_10.flop6/_1__208  (.L_HI(net254));
 sg13g2_dfrbp_1 \proj_10.flop6/_1_  (.CLK(clknet_5_26__leaf_clk_regs),
    .RESET_B(net254),
    .D(net433),
    .Q_N(\proj_10.flop6/notq ),
    .Q(\proj_10.net12 ));
 sg13g2_tiehi \proj_10.flop7/_1__209  (.L_HI(net255));
 sg13g2_dfrbp_1 \proj_10.flop7/_1_  (.CLK(clknet_5_27__leaf_clk_regs),
    .RESET_B(net255),
    .D(\proj_10.net32 ),
    .Q_N(\proj_10.flop7/notq ),
    .Q(\proj_10.net11 ));
 sg13g2_tiehi \proj_10.flop8/_1__210  (.L_HI(net256));
 sg13g2_dfrbp_1 \proj_10.flop8/_1_  (.CLK(clknet_5_27__leaf_clk_regs),
    .RESET_B(net256),
    .D(net427),
    .Q_N(\proj_10.flop8/notq ),
    .Q(\proj_10.net10 ));
 sg13g2_tiehi \proj_10.flop9/_1__211  (.L_HI(net257));
 sg13g2_dfrbp_1 \proj_10.flop9/_1_  (.CLK(clknet_5_12__leaf_clk_regs),
    .RESET_B(net257),
    .D(net150),
    .Q_N(\proj_10.flop9/notq ),
    .Q(\proj_10.net45 ));
 sg13g2_tiehi \proj_14.flop1/_1__212  (.L_HI(net258));
 sg13g2_inv_1 \proj_10.not1/_0_  (.Y(\proj_10.net24 ),
    .A(\proj_10.net31 ));
 sg13g2_inv_1 \proj_10.not2/_0_  (.Y(\proj_10.net27 ),
    .A(net434));
 sg13g2_inv_1 \proj_10.not3/_0_  (.Y(\proj_10.net37 ),
    .A(net430));
 sg13g2_inv_1 \proj_10.not5/_0_  (.Y(\proj_10.net39 ),
    .A(\proj_10.net38 ));
 sg13g2_inv_1 \proj_10.not6/_0_  (.Y(\proj_10.net23 ),
    .A(net427));
 sg13g2_inv_1 \proj_10.not7/_0_  (.Y(\proj_10.net33 ),
    .A(net432));
 sg13g2_xor2_1 \proj_10.xor1/_0_  (.B(clknet_1_1__leaf_clk),
    .A(net1),
    .X(\proj_10.net17 ));
 sg13g2_and2_1 \proj_11.and1/_0_  (.A(net6),
    .B(net180),
    .X(\proj_11.net19 ));
 sg13g2_and2_1 \proj_11.and2/_0_  (.A(\proj_11.net20 ),
    .B(\proj_11.net19 ),
    .X(\proj_11.net21 ));
 sg13g2_and2_1 \proj_11.and3/_0_  (.A(net171),
    .B(net176),
    .X(\proj_11.net22 ));
 sg13g2_and2_1 \proj_11.and4/_0_  (.A(net164),
    .B(net174),
    .X(\proj_11.net24 ));
 sg13g2_and2_1 \proj_11.and5/_0_  (.A(\proj_11.net25 ),
    .B(\proj_11.net23 ),
    .X(\proj_11.net26 ));
 sg13g2_and2_1 \proj_11.and6/_0_  (.A(net136),
    .B(net173),
    .X(\proj_11.net28 ));
 sg13g2_and2_1 \proj_11.and7/_0_  (.A(\proj_11.net29 ),
    .B(\proj_11.net27 ),
    .X(\proj_11.net30 ));
 sg13g2_or2_1 \proj_11.or1/_0_  (.X(\proj_11.net23 ),
    .B(\proj_11.net21 ),
    .A(\proj_11.net22 ));
 sg13g2_or2_1 \proj_11.or2/_0_  (.X(\proj_11.net27 ),
    .B(\proj_11.net26 ),
    .A(\proj_11.net24 ));
 sg13g2_or2_1 \proj_11.or3/_0_  (.X(\proj_11.net13 ),
    .B(\proj_11.net30 ),
    .A(\proj_11.net28 ));
 sg13g2_xor2_1 \proj_11.xor1/_0_  (.B(net179),
    .A(net6),
    .X(\proj_11.net9 ));
 sg13g2_xor2_1 \proj_11.xor2/_0_  (.B(net176),
    .A(net7),
    .X(\proj_11.net20 ));
 sg13g2_xor2_1 \proj_11.xor3/_0_  (.B(\proj_11.net20 ),
    .A(\proj_11.net19 ),
    .X(\proj_11.net10 ));
 sg13g2_xor2_1 \proj_11.xor4/_0_  (.B(\proj_11.net25 ),
    .A(\proj_11.net23 ),
    .X(\proj_11.net11 ));
 sg13g2_xor2_1 \proj_11.xor5/_0_  (.B(net174),
    .A(net163),
    .X(\proj_11.net25 ));
 sg13g2_xor2_1 \proj_11.xor6/_0_  (.B(net173),
    .A(net136),
    .X(\proj_11.net29 ));
 sg13g2_xor2_1 \proj_11.xor7/_0_  (.B(\proj_11.net29 ),
    .A(\proj_11.net27 ),
    .X(\proj_11.net12 ));
 sg13g2_and2_1 \proj_12.and1/_0_  (.A(net179),
    .B(net178),
    .X(\proj_12.net21 ));
 sg13g2_and2_1 \proj_12.and2/_0_  (.A(net172),
    .B(net5),
    .X(\proj_12.net12 ));
 sg13g2_mux2_1 \proj_12.mux1/_0_  (.A0(\proj_12.net21 ),
    .A1(\proj_12.net20 ),
    .S(net4),
    .X(\proj_12.net22 ));
 sg13g2_nand2_1 \proj_12.nand1/_0_  (.Y(\proj_12.net20 ),
    .A(net1),
    .B(clknet_1_0__leaf_clk));
 sg13g2_nand2_1 \proj_12.nand2/_0_  (.Y(\proj_12.net13 ),
    .A(net164),
    .B(net171));
 sg13g2_buf_2 clkbuf_regs_0_clk (.A(clk),
    .X(clk_regs));
 sg13g2_xor2_1 \proj_12.xor1/_0_  (.B(net136),
    .A(net152),
    .X(\proj_12.net14 ));
 sg13g2_and2_1 \proj_13.and1/_0_  (.A(net175),
    .B(net136),
    .X(\proj_13.net13 ));
 sg13g2_and2_1 \proj_13.and2/_0_  (.A(\proj_13.net14 ),
    .B(\proj_13.net23 ),
    .X(\proj_13.net10 ));
 sg13g2_and2_1 \proj_13.and3/_0_  (.A(\proj_13.net24 ),
    .B(\proj_13.net22 ),
    .X(\proj_13.net11 ));
 sg13g2_and2_1 \proj_13.and4/_0_  (.A(net164),
    .B(net172),
    .X(\proj_13.net14 ));
 sg13g2_nand2_1 \proj_13.nand1/_0_  (.Y(\proj_13.net9 ),
    .A(net177),
    .B(\proj_13.net21 ));
 sg13g2_nand2_1 \proj_13.nand2/_0_  (.Y(\proj_13.net21 ),
    .A(\proj_13.net13 ),
    .B(\proj_13.net20 ));
 sg13g2_inv_1 \proj_13.not1/_0_  (.Y(\proj_13.net20 ),
    .A(net180));
 sg13g2_inv_1 \proj_13.not2/_0_  (.Y(\proj_13.net24 ),
    .A(net175));
 sg13g2_or2_1 \proj_13.or1/_0_  (.X(\proj_13.net22 ),
    .B(\proj_13.net14 ),
    .A(\proj_13.net12 ));
 sg13g2_or2_1 \proj_13.or2/_0_  (.X(\proj_13.net23 ),
    .B(net173),
    .A(net171));
 sg13g2_xor2_1 \proj_13.xor1/_0_  (.B(net177),
    .A(net174),
    .X(\proj_13.net12 ));
 sg13g2_dfrbp_1 \proj_14.flop1/_1_  (.CLK(clknet_5_14__leaf_clk_regs),
    .RESET_B(net258),
    .D(\proj_14.net8 ),
    .Q_N(\proj_14.flop1/notq ),
    .Q(\proj_14.net9 ));
 sg13g2_tiehi \proj_14.flop10/_1__213  (.L_HI(net259));
 sg13g2_dfrbp_1 \proj_14.flop10/_1_  (.CLK(clknet_5_14__leaf_clk_regs),
    .RESET_B(net259),
    .D(\proj_14.net33 ),
    .Q_N(\proj_14.flop10/notq ),
    .Q(\proj_14.net32 ));
 sg13g2_tiehi \proj_14.flop100/_1__214  (.L_HI(net260));
 sg13g2_dfrbp_1 \proj_14.flop100/_1_  (.CLK(clknet_5_23__leaf_clk_regs),
    .RESET_B(net260),
    .D(\proj_14.net313 ),
    .Q_N(\proj_14.flop100/notq ),
    .Q(\proj_14.net312 ));
 sg13g2_tiehi \proj_14.flop101/_1__215  (.L_HI(net261));
 sg13g2_dfrbp_1 \proj_14.flop101/_1_  (.CLK(clknet_5_22__leaf_clk_regs),
    .RESET_B(net261),
    .D(\proj_14.net316 ),
    .Q_N(\proj_14.flop101/notq ),
    .Q(\proj_14.net315 ));
 sg13g2_tiehi \proj_14.flop102/_1__216  (.L_HI(net262));
 sg13g2_dfrbp_1 \proj_14.flop102/_1_  (.CLK(clknet_5_5__leaf_clk_regs),
    .RESET_B(net262),
    .D(\proj_14.net320 ),
    .Q_N(\proj_14.flop102/notq ),
    .Q(\proj_14.net254 ));
 sg13g2_tiehi \proj_14.flop103/_1__217  (.L_HI(net263));
 sg13g2_dfrbp_1 \proj_14.flop103/_1_  (.CLK(clknet_5_5__leaf_clk_regs),
    .RESET_B(net263),
    .D(\proj_14.net323 ),
    .Q_N(\proj_14.flop103/notq ),
    .Q(\proj_14.net322 ));
 sg13g2_tiehi \proj_14.flop104/_1__218  (.L_HI(net264));
 sg13g2_dfrbp_1 \proj_14.flop104/_1_  (.CLK(clknet_5_17__leaf_clk_regs),
    .RESET_B(net264),
    .D(\proj_14.net326 ),
    .Q_N(\proj_14.flop104/notq ),
    .Q(\proj_14.net325 ));
 sg13g2_tiehi \proj_14.flop105/_1__219  (.L_HI(net265));
 sg13g2_dfrbp_1 \proj_14.flop105/_1_  (.CLK(clknet_5_17__leaf_clk_regs),
    .RESET_B(net265),
    .D(\proj_14.net329 ),
    .Q_N(\proj_14.flop105/notq ),
    .Q(\proj_14.net328 ));
 sg13g2_tiehi \proj_14.flop106/_1__220  (.L_HI(net266));
 sg13g2_dfrbp_1 \proj_14.flop106/_1_  (.CLK(clknet_5_22__leaf_clk_regs),
    .RESET_B(net266),
    .D(\proj_14.net332 ),
    .Q_N(\proj_14.flop106/notq ),
    .Q(\proj_14.net333 ));
 sg13g2_tiehi \proj_14.flop107/_1__221  (.L_HI(net267));
 sg13g2_dfrbp_1 \proj_14.flop107/_1_  (.CLK(clknet_5_25__leaf_clk_regs),
    .RESET_B(net267),
    .D(\proj_14.net336 ),
    .Q_N(\proj_14.flop107/notq ),
    .Q(\proj_14.net335 ));
 sg13g2_tiehi \proj_14.flop108/_1__222  (.L_HI(net268));
 sg13g2_dfrbp_1 \proj_14.flop108/_1_  (.CLK(clknet_5_19__leaf_clk_regs),
    .RESET_B(net268),
    .D(\proj_14.net339 ),
    .Q_N(\proj_14.flop108/notq ),
    .Q(\proj_14.net338 ));
 sg13g2_tiehi \proj_14.flop109/_1__223  (.L_HI(net269));
 sg13g2_dfrbp_1 \proj_14.flop109/_1_  (.CLK(clknet_5_19__leaf_clk_regs),
    .RESET_B(net269),
    .D(\proj_14.net342 ),
    .Q_N(\proj_14.flop109/notq ),
    .Q(\proj_14.net341 ));
 sg13g2_tiehi \proj_14.flop11/_1__224  (.L_HI(net270));
 sg13g2_dfrbp_1 \proj_14.flop11/_1_  (.CLK(clknet_5_11__leaf_clk_regs),
    .RESET_B(net270),
    .D(\proj_14.net36 ),
    .Q_N(\proj_14.flop11/notq ),
    .Q(\proj_14.net35 ));
 sg13g2_tiehi \proj_14.flop110/_1__225  (.L_HI(net271));
 sg13g2_dfrbp_1 \proj_14.flop110/_1_  (.CLK(clknet_5_18__leaf_clk_regs),
    .RESET_B(net271),
    .D(\proj_14.net345 ),
    .Q_N(\proj_14.flop110/notq ),
    .Q(\proj_14.net344 ));
 sg13g2_tiehi \proj_14.flop111/_1__226  (.L_HI(net272));
 sg13g2_dfrbp_1 \proj_14.flop111/_1_  (.CLK(clknet_5_24__leaf_clk_regs),
    .RESET_B(net272),
    .D(\proj_14.net348 ),
    .Q_N(\proj_14.flop111/notq ),
    .Q(\proj_14.net347 ));
 sg13g2_tiehi \proj_14.flop112/_1__227  (.L_HI(net273));
 sg13g2_dfrbp_1 \proj_14.flop112/_1_  (.CLK(clknet_5_24__leaf_clk_regs),
    .RESET_B(net273),
    .D(\proj_14.net351 ),
    .Q_N(\proj_14.flop112/notq ),
    .Q(\proj_14.net350 ));
 sg13g2_tiehi \proj_14.flop113/_1__228  (.L_HI(net274));
 sg13g2_dfrbp_1 \proj_14.flop113/_1_  (.CLK(clknet_5_24__leaf_clk_regs),
    .RESET_B(net274),
    .D(\proj_14.net354 ),
    .Q_N(\proj_14.flop113/notq ),
    .Q(\proj_14.net353 ));
 sg13g2_tiehi \proj_14.flop114/_1__229  (.L_HI(net275));
 sg13g2_dfrbp_1 \proj_14.flop114/_1_  (.CLK(clknet_5_25__leaf_clk_regs),
    .RESET_B(net275),
    .D(\proj_14.net357 ),
    .Q_N(\proj_14.flop114/notq ),
    .Q(\proj_14.net356 ));
 sg13g2_tiehi \proj_14.flop115/_1__230  (.L_HI(net276));
 sg13g2_dfrbp_1 \proj_14.flop115/_1_  (.CLK(clknet_5_25__leaf_clk_regs),
    .RESET_B(net276),
    .D(\proj_14.net360 ),
    .Q_N(\proj_14.flop115/notq ),
    .Q(\proj_14.net359 ));
 sg13g2_tiehi \proj_14.flop116/_1__231  (.L_HI(net277));
 sg13g2_dfrbp_1 \proj_14.flop116/_1_  (.CLK(clknet_5_28__leaf_clk_regs),
    .RESET_B(net277),
    .D(\proj_14.net363 ),
    .Q_N(\proj_14.flop116/notq ),
    .Q(\proj_14.net362 ));
 sg13g2_tiehi \proj_14.flop117/_1__232  (.L_HI(net278));
 sg13g2_dfrbp_1 \proj_14.flop117/_1_  (.CLK(clknet_5_29__leaf_clk_regs),
    .RESET_B(net278),
    .D(\proj_14.net366 ),
    .Q_N(\proj_14.flop117/notq ),
    .Q(\proj_14.net365 ));
 sg13g2_tiehi \proj_14.flop118/_1__233  (.L_HI(net279));
 sg13g2_dfrbp_1 \proj_14.flop118/_1_  (.CLK(clknet_5_28__leaf_clk_regs),
    .RESET_B(net279),
    .D(\proj_14.net369 ),
    .Q_N(\proj_14.flop118/notq ),
    .Q(\proj_14.net368 ));
 sg13g2_tiehi \proj_14.flop119/_1__234  (.L_HI(net280));
 sg13g2_dfrbp_1 \proj_14.flop119/_1_  (.CLK(clknet_5_25__leaf_clk_regs),
    .RESET_B(net280),
    .D(\proj_14.net372 ),
    .Q_N(\proj_14.flop119/notq ),
    .Q(\proj_14.net371 ));
 sg13g2_tiehi \proj_14.flop12/_1__235  (.L_HI(net281));
 sg13g2_dfrbp_1 \proj_14.flop12/_1_  (.CLK(clknet_5_10__leaf_clk_regs),
    .RESET_B(net281),
    .D(\proj_14.net39 ),
    .Q_N(\proj_14.flop12/notq ),
    .Q(\proj_14.net38 ));
 sg13g2_tiehi \proj_14.flop120/_1__236  (.L_HI(net282));
 sg13g2_dfrbp_1 \proj_14.flop120/_1_  (.CLK(clknet_5_24__leaf_clk_regs),
    .RESET_B(net282),
    .D(\proj_14.net375 ),
    .Q_N(\proj_14.flop120/notq ),
    .Q(\proj_14.net374 ));
 sg13g2_tiehi \proj_14.flop121/_1__237  (.L_HI(net283));
 sg13g2_dfrbp_1 \proj_14.flop121/_1_  (.CLK(clknet_5_25__leaf_clk_regs),
    .RESET_B(net283),
    .D(\proj_14.net378 ),
    .Q_N(\proj_14.flop121/notq ),
    .Q(\proj_14.net377 ));
 sg13g2_tiehi \proj_14.flop122/_1__238  (.L_HI(net284));
 sg13g2_dfrbp_1 \proj_14.flop122/_1_  (.CLK(clknet_5_19__leaf_clk_regs),
    .RESET_B(net284),
    .D(\proj_14.net381 ),
    .Q_N(\proj_14.flop122/notq ),
    .Q(\proj_14.net380 ));
 sg13g2_tiehi \proj_14.flop123/_1__239  (.L_HI(net285));
 sg13g2_dfrbp_1 \proj_14.flop123/_1_  (.CLK(clknet_5_22__leaf_clk_regs),
    .RESET_B(net285),
    .D(\proj_14.net385 ),
    .Q_N(\proj_14.flop123/notq ),
    .Q(\proj_14.net318 ));
 sg13g2_tiehi \proj_14.flop124/_1__240  (.L_HI(net286));
 sg13g2_dfrbp_1 \proj_14.flop124/_1_  (.CLK(clknet_5_22__leaf_clk_regs),
    .RESET_B(net286),
    .D(\proj_14.net388 ),
    .Q_N(\proj_14.flop124/notq ),
    .Q(\proj_14.net387 ));
 sg13g2_tiehi \proj_14.flop125/_1__241  (.L_HI(net287));
 sg13g2_dfrbp_1 \proj_14.flop125/_1_  (.CLK(clknet_5_28__leaf_clk_regs),
    .RESET_B(net287),
    .D(\proj_14.net391 ),
    .Q_N(\proj_14.flop125/notq ),
    .Q(\proj_14.net390 ));
 sg13g2_tiehi \proj_14.flop126/_1__242  (.L_HI(net288));
 sg13g2_dfrbp_1 \proj_14.flop126/_1_  (.CLK(clknet_5_28__leaf_clk_regs),
    .RESET_B(net288),
    .D(\proj_14.net394 ),
    .Q_N(\proj_14.flop126/notq ),
    .Q(\proj_14.net393 ));
 sg13g2_tiehi \proj_14.flop127/_1__243  (.L_HI(net289));
 sg13g2_dfrbp_1 \proj_14.flop127/_1_  (.CLK(clknet_5_6__leaf_clk_regs),
    .RESET_B(net289),
    .D(\proj_14.net396 ),
    .Q_N(\proj_14.flop127/notq ),
    .Q(\proj_14.net397 ));
 sg13g2_tiehi \proj_14.flop128/_1__244  (.L_HI(net290));
 sg13g2_dfrbp_1 \proj_14.flop128/_1_  (.CLK(clknet_5_18__leaf_clk_regs),
    .RESET_B(net290),
    .D(\proj_14.net400 ),
    .Q_N(\proj_14.flop128/notq ),
    .Q(\proj_14.net399 ));
 sg13g2_tiehi \proj_14.flop129/_1__245  (.L_HI(net291));
 sg13g2_dfrbp_1 \proj_14.flop129/_1_  (.CLK(clknet_5_6__leaf_clk_regs),
    .RESET_B(net291),
    .D(\proj_14.net403 ),
    .Q_N(\proj_14.flop129/notq ),
    .Q(\proj_14.net402 ));
 sg13g2_tiehi \proj_14.flop13/_1__246  (.L_HI(net292));
 sg13g2_dfrbp_1 \proj_14.flop13/_1_  (.CLK(clknet_5_10__leaf_clk_regs),
    .RESET_B(net292),
    .D(\proj_14.net42 ),
    .Q_N(\proj_14.flop13/notq ),
    .Q(\proj_14.net41 ));
 sg13g2_tiehi \proj_14.flop130/_1__247  (.L_HI(net293));
 sg13g2_dfrbp_1 \proj_14.flop130/_1_  (.CLK(clknet_5_6__leaf_clk_regs),
    .RESET_B(net293),
    .D(\proj_14.net406 ),
    .Q_N(\proj_14.flop130/notq ),
    .Q(\proj_14.net405 ));
 sg13g2_tiehi \proj_14.flop131/_1__248  (.L_HI(net294));
 sg13g2_dfrbp_1 \proj_14.flop131/_1_  (.CLK(clknet_5_6__leaf_clk_regs),
    .RESET_B(net294),
    .D(\proj_14.net409 ),
    .Q_N(\proj_14.flop131/notq ),
    .Q(\proj_14.net408 ));
 sg13g2_tiehi \proj_14.flop132/_1__249  (.L_HI(net295));
 sg13g2_dfrbp_1 \proj_14.flop132/_1_  (.CLK(clknet_5_3__leaf_clk_regs),
    .RESET_B(net295),
    .D(\proj_14.net412 ),
    .Q_N(\proj_14.flop132/notq ),
    .Q(\proj_14.net411 ));
 sg13g2_tiehi \proj_14.flop133/_1__250  (.L_HI(net296));
 sg13g2_dfrbp_1 \proj_14.flop133/_1_  (.CLK(clknet_5_2__leaf_clk_regs),
    .RESET_B(net296),
    .D(\proj_14.net415 ),
    .Q_N(\proj_14.flop133/notq ),
    .Q(\proj_14.net414 ));
 sg13g2_tiehi \proj_14.flop134/_1__251  (.L_HI(net297));
 sg13g2_dfrbp_1 \proj_14.flop134/_1_  (.CLK(clknet_5_5__leaf_clk_regs),
    .RESET_B(net297),
    .D(\proj_14.net418 ),
    .Q_N(\proj_14.flop134/notq ),
    .Q(\proj_14.net417 ));
 sg13g2_tiehi \proj_14.flop135/_1__252  (.L_HI(net298));
 sg13g2_dfrbp_1 \proj_14.flop135/_1_  (.CLK(clknet_5_4__leaf_clk_regs),
    .RESET_B(net298),
    .D(\proj_14.net421 ),
    .Q_N(\proj_14.flop135/notq ),
    .Q(\proj_14.net420 ));
 sg13g2_tiehi \proj_14.flop136/_1__253  (.L_HI(net299));
 sg13g2_dfrbp_1 \proj_14.flop136/_1_  (.CLK(clknet_5_1__leaf_clk_regs),
    .RESET_B(net299),
    .D(\proj_14.net424 ),
    .Q_N(\proj_14.flop136/notq ),
    .Q(\proj_14.net423 ));
 sg13g2_tiehi \proj_14.flop137/_1__254  (.L_HI(net300));
 sg13g2_dfrbp_1 \proj_14.flop137/_1_  (.CLK(clknet_5_4__leaf_clk_regs),
    .RESET_B(net300),
    .D(\proj_14.net427 ),
    .Q_N(\proj_14.flop137/notq ),
    .Q(\proj_14.net426 ));
 sg13g2_tiehi \proj_14.flop138/_1__255  (.L_HI(net301));
 sg13g2_dfrbp_1 \proj_14.flop138/_1_  (.CLK(clknet_5_1__leaf_clk_regs),
    .RESET_B(net301),
    .D(\proj_14.net430 ),
    .Q_N(\proj_14.flop138/notq ),
    .Q(\proj_14.net429 ));
 sg13g2_tiehi \proj_14.flop139/_1__256  (.L_HI(net302));
 sg13g2_dfrbp_1 \proj_14.flop139/_1_  (.CLK(clknet_5_1__leaf_clk_regs),
    .RESET_B(net302),
    .D(\proj_14.net433 ),
    .Q_N(\proj_14.flop139/notq ),
    .Q(\proj_14.net432 ));
 sg13g2_tiehi \proj_14.flop14/_1__257  (.L_HI(net303));
 sg13g2_dfrbp_1 \proj_14.flop14/_1_  (.CLK(clknet_5_10__leaf_clk_regs),
    .RESET_B(net303),
    .D(\proj_14.net45 ),
    .Q_N(\proj_14.flop14/notq ),
    .Q(\proj_14.net44 ));
 sg13g2_tiehi \proj_14.flop140/_1__258  (.L_HI(net304));
 sg13g2_dfrbp_1 \proj_14.flop140/_1_  (.CLK(clknet_5_0__leaf_clk_regs),
    .RESET_B(net304),
    .D(\proj_14.net436 ),
    .Q_N(\proj_14.flop140/notq ),
    .Q(\proj_14.net435 ));
 sg13g2_tiehi \proj_14.flop141/_1__259  (.L_HI(net305));
 sg13g2_dfrbp_1 \proj_14.flop141/_1_  (.CLK(clknet_5_0__leaf_clk_regs),
    .RESET_B(net305),
    .D(\proj_14.net439 ),
    .Q_N(\proj_14.flop141/notq ),
    .Q(\proj_14.net438 ));
 sg13g2_tiehi \proj_14.flop142/_1__260  (.L_HI(net306));
 sg13g2_dfrbp_1 \proj_14.flop142/_1_  (.CLK(clknet_5_0__leaf_clk_regs),
    .RESET_B(net306),
    .D(\proj_14.net442 ),
    .Q_N(\proj_14.flop142/notq ),
    .Q(\proj_14.net441 ));
 sg13g2_tiehi \proj_14.flop143/_1__261  (.L_HI(net307));
 sg13g2_dfrbp_1 \proj_14.flop143/_1_  (.CLK(clknet_5_1__leaf_clk_regs),
    .RESET_B(net307),
    .D(\proj_14.net445 ),
    .Q_N(\proj_14.flop143/notq ),
    .Q(\proj_14.net444 ));
 sg13g2_tiehi \proj_14.flop144/_1__262  (.L_HI(net308));
 sg13g2_dfrbp_1 \proj_14.flop144/_1_  (.CLK(clknet_5_19__leaf_clk_regs),
    .RESET_B(net308),
    .D(\proj_14.net449 ),
    .Q_N(\proj_14.flop144/notq ),
    .Q(\proj_14.net383 ));
 sg13g2_tiehi \proj_14.flop145/_1__263  (.L_HI(net309));
 sg13g2_dfrbp_1 \proj_14.flop145/_1_  (.CLK(clknet_5_18__leaf_clk_regs),
    .RESET_B(net309),
    .D(\proj_14.net452 ),
    .Q_N(\proj_14.flop145/notq ),
    .Q(\proj_14.net451 ));
 sg13g2_tiehi \proj_14.flop146/_1__264  (.L_HI(net310));
 sg13g2_dfrbp_1 \proj_14.flop146/_1_  (.CLK(clknet_5_18__leaf_clk_regs),
    .RESET_B(net310),
    .D(\proj_14.net455 ),
    .Q_N(\proj_14.flop146/notq ),
    .Q(\proj_14.net454 ));
 sg13g2_tiehi \proj_14.flop147/_1__265  (.L_HI(net311));
 sg13g2_dfrbp_1 \proj_14.flop147/_1_  (.CLK(clknet_5_7__leaf_clk_regs),
    .RESET_B(net311),
    .D(\proj_14.net458 ),
    .Q_N(\proj_14.flop147/notq ),
    .Q(\proj_14.net457 ));
 sg13g2_tiehi \proj_14.flop148/_1__266  (.L_HI(net312));
 sg13g2_dfrbp_1 \proj_14.flop148/_1_  (.CLK(clknet_5_2__leaf_clk_regs),
    .RESET_B(net312),
    .D(\proj_14.net460 ),
    .Q_N(\proj_14.flop148/notq ),
    .Q(\proj_14.net461 ));
 sg13g2_tiehi \proj_14.flop149/_1__267  (.L_HI(net313));
 sg13g2_dfrbp_1 \proj_14.flop149/_1_  (.CLK(clknet_5_2__leaf_clk_regs),
    .RESET_B(net313),
    .D(\proj_14.net464 ),
    .Q_N(\proj_14.flop149/notq ),
    .Q(\proj_14.net463 ));
 sg13g2_tiehi \proj_14.flop15/_1__268  (.L_HI(net314));
 sg13g2_dfrbp_1 \proj_14.flop15/_1_  (.CLK(clknet_5_10__leaf_clk_regs),
    .RESET_B(net314),
    .D(\proj_14.net48 ),
    .Q_N(\proj_14.flop15/notq ),
    .Q(\proj_14.net47 ));
 sg13g2_tiehi \proj_14.flop150/_1__269  (.L_HI(net315));
 sg13g2_dfrbp_1 \proj_14.flop150/_1_  (.CLK(clknet_5_2__leaf_clk_regs),
    .RESET_B(net315),
    .D(\proj_14.net467 ),
    .Q_N(\proj_14.flop150/notq ),
    .Q(\proj_14.net466 ));
 sg13g2_tiehi \proj_14.flop151/_1__270  (.L_HI(net316));
 sg13g2_dfrbp_1 \proj_14.flop151/_1_  (.CLK(clknet_5_3__leaf_clk_regs),
    .RESET_B(net316),
    .D(\proj_14.net470 ),
    .Q_N(\proj_14.flop151/notq ),
    .Q(\proj_14.net469 ));
 sg13g2_tiehi \proj_14.flop152/_1__271  (.L_HI(net317));
 sg13g2_dfrbp_1 \proj_14.flop152/_1_  (.CLK(clknet_5_3__leaf_clk_regs),
    .RESET_B(net317),
    .D(\proj_14.net473 ),
    .Q_N(\proj_14.flop152/notq ),
    .Q(\proj_14.net472 ));
 sg13g2_tiehi \proj_14.flop153/_1__272  (.L_HI(net318));
 sg13g2_dfrbp_1 \proj_14.flop153/_1_  (.CLK(clknet_5_3__leaf_clk_regs),
    .RESET_B(net318),
    .D(\proj_14.net476 ),
    .Q_N(\proj_14.flop153/notq ),
    .Q(\proj_14.net475 ));
 sg13g2_tiehi \proj_14.flop154/_1__273  (.L_HI(net319));
 sg13g2_dfrbp_1 \proj_14.flop154/_1_  (.CLK(clknet_5_7__leaf_clk_regs),
    .RESET_B(net319),
    .D(\proj_14.net479 ),
    .Q_N(\proj_14.flop154/notq ),
    .Q(\proj_14.net478 ));
 sg13g2_tiehi \proj_14.flop155/_1__274  (.L_HI(net320));
 sg13g2_dfrbp_1 \proj_14.flop155/_1_  (.CLK(clknet_5_9__leaf_clk_regs),
    .RESET_B(net320),
    .D(\proj_14.net482 ),
    .Q_N(\proj_14.flop155/notq ),
    .Q(\proj_14.net481 ));
 sg13g2_tiehi \proj_14.flop156/_1__275  (.L_HI(net321));
 sg13g2_dfrbp_1 \proj_14.flop156/_1_  (.CLK(clknet_5_9__leaf_clk_regs),
    .RESET_B(net321),
    .D(\proj_14.net485 ),
    .Q_N(\proj_14.flop156/notq ),
    .Q(\proj_14.net484 ));
 sg13g2_tiehi \proj_14.flop157/_1__276  (.L_HI(net322));
 sg13g2_dfrbp_1 \proj_14.flop157/_1_  (.CLK(clknet_5_9__leaf_clk_regs),
    .RESET_B(net322),
    .D(\proj_14.net488 ),
    .Q_N(\proj_14.flop157/notq ),
    .Q(\proj_14.net487 ));
 sg13g2_tiehi \proj_14.flop158/_1__277  (.L_HI(net323));
 sg13g2_dfrbp_1 \proj_14.flop158/_1_  (.CLK(clknet_5_8__leaf_clk_regs),
    .RESET_B(net323),
    .D(\proj_14.net491 ),
    .Q_N(\proj_14.flop158/notq ),
    .Q(\proj_14.net490 ));
 sg13g2_tiehi \proj_14.flop159/_1__278  (.L_HI(net324));
 sg13g2_dfrbp_1 \proj_14.flop159/_1_  (.CLK(clknet_5_14__leaf_clk_regs),
    .RESET_B(net324),
    .D(\proj_14.net494 ),
    .Q_N(\proj_14.flop159/notq ),
    .Q(\proj_14.net493 ));
 sg13g2_tiehi \proj_14.flop16/_1__279  (.L_HI(net325));
 sg13g2_dfrbp_1 \proj_14.flop16/_1_  (.CLK(clknet_5_8__leaf_clk_regs),
    .RESET_B(net325),
    .D(\proj_14.net51 ),
    .Q_N(\proj_14.flop16/notq ),
    .Q(\proj_14.net50 ));
 sg13g2_tiehi \proj_14.flop160/_1__280  (.L_HI(net326));
 sg13g2_dfrbp_1 \proj_14.flop160/_1_  (.CLK(clknet_5_14__leaf_clk_regs),
    .RESET_B(net326),
    .D(\proj_14.net497 ),
    .Q_N(\proj_14.flop160/notq ),
    .Q(\proj_14.net496 ));
 sg13g2_tiehi \proj_14.flop161/_1__281  (.L_HI(net327));
 sg13g2_dfrbp_1 \proj_14.flop161/_1_  (.CLK(clknet_5_11__leaf_clk_regs),
    .RESET_B(net327),
    .D(\proj_14.net500 ),
    .Q_N(\proj_14.flop161/notq ),
    .Q(\proj_14.net499 ));
 sg13g2_tiehi \proj_14.flop162/_1__282  (.L_HI(net328));
 sg13g2_dfrbp_1 \proj_14.flop162/_1_  (.CLK(clknet_5_11__leaf_clk_regs),
    .RESET_B(net328),
    .D(\proj_14.net503 ),
    .Q_N(\proj_14.flop162/notq ),
    .Q(\proj_14.net502 ));
 sg13g2_tiehi \proj_14.flop163/_1__283  (.L_HI(net329));
 sg13g2_dfrbp_1 \proj_14.flop163/_1_  (.CLK(clknet_5_11__leaf_clk_regs),
    .RESET_B(net329),
    .D(\proj_14.net506 ),
    .Q_N(\proj_14.flop163/notq ),
    .Q(\proj_14.net505 ));
 sg13g2_tiehi \proj_14.flop164/_1__284  (.L_HI(net330));
 sg13g2_dfrbp_1 \proj_14.flop164/_1_  (.CLK(clknet_5_15__leaf_clk_regs),
    .RESET_B(net330),
    .D(\proj_14.net509 ),
    .Q_N(\proj_14.flop164/notq ),
    .Q(\proj_14.net508 ));
 sg13g2_tiehi \proj_14.flop165/_1__285  (.L_HI(net331));
 sg13g2_dfrbp_1 \proj_14.flop165/_1_  (.CLK(clknet_5_0__leaf_clk_regs),
    .RESET_B(net331),
    .D(\proj_14.net512 ),
    .Q_N(\proj_14.flop165/notq ),
    .Q(\proj_14.net447 ));
 sg13g2_tiehi \proj_14.flop166/_1__286  (.L_HI(net332));
 sg13g2_dfrbp_1 \proj_14.flop166/_1_  (.CLK(clknet_5_0__leaf_clk_regs),
    .RESET_B(net332),
    .D(\proj_14.net515 ),
    .Q_N(\proj_14.flop166/notq ),
    .Q(\proj_14.net514 ));
 sg13g2_tiehi \proj_14.flop167/_1__287  (.L_HI(net333));
 sg13g2_dfrbp_1 \proj_14.flop167/_1_  (.CLK(clknet_5_0__leaf_clk_regs),
    .RESET_B(net333),
    .D(\proj_14.net518 ),
    .Q_N(\proj_14.flop167/notq ),
    .Q(\proj_14.net517 ));
 sg13g2_tiehi \proj_14.flop168/_1__288  (.L_HI(net334));
 sg13g2_dfrbp_1 \proj_14.flop168/_1_  (.CLK(clknet_5_2__leaf_clk_regs),
    .RESET_B(net334),
    .D(\proj_14.net521 ),
    .Q_N(\proj_14.flop168/notq ),
    .Q(\proj_14.net520 ));
 sg13g2_tiehi \proj_14.flop17/_1__289  (.L_HI(net335));
 sg13g2_dfrbp_1 \proj_14.flop17/_1_  (.CLK(clknet_5_8__leaf_clk_regs),
    .RESET_B(net335),
    .D(\proj_14.net54 ),
    .Q_N(\proj_14.flop17/notq ),
    .Q(\proj_14.net53 ));
 sg13g2_tiehi \proj_14.flop18/_1__290  (.L_HI(net336));
 sg13g2_dfrbp_1 \proj_14.flop18/_1_  (.CLK(clknet_5_8__leaf_clk_regs),
    .RESET_B(net336),
    .D(\proj_14.net57 ),
    .Q_N(\proj_14.flop18/notq ),
    .Q(\proj_14.net56 ));
 sg13g2_tiehi \proj_14.flop19/_1__291  (.L_HI(net337));
 sg13g2_dfrbp_1 \proj_14.flop19/_1_  (.CLK(clknet_5_6__leaf_clk_regs),
    .RESET_B(net337),
    .D(\proj_14.net67 ),
    .Q_N(\proj_14.flop19/notq ),
    .Q(\proj_14.net66 ));
 sg13g2_tiehi \proj_14.flop2/_1__292  (.L_HI(net338));
 sg13g2_dfrbp_1 \proj_14.flop2/_1_  (.CLK(clknet_5_3__leaf_clk_regs),
    .RESET_B(net338),
    .D(\proj_14.net63 ),
    .Q_N(\proj_14.flop2/notq ),
    .Q(\proj_14.net64 ));
 sg13g2_tiehi \proj_14.flop20/_1__293  (.L_HI(net339));
 sg13g2_dfrbp_1 \proj_14.flop20/_1_  (.CLK(clknet_5_6__leaf_clk_regs),
    .RESET_B(net339),
    .D(\proj_14.net70 ),
    .Q_N(\proj_14.flop20/notq ),
    .Q(\proj_14.net69 ));
 sg13g2_tiehi \proj_14.flop21/_1__294  (.L_HI(net340));
 sg13g2_dfrbp_1 \proj_14.flop21/_1_  (.CLK(clknet_5_7__leaf_clk_regs),
    .RESET_B(net340),
    .D(\proj_14.net73 ),
    .Q_N(\proj_14.flop21/notq ),
    .Q(\proj_14.net72 ));
 sg13g2_tiehi \proj_14.flop22/_1__295  (.L_HI(net341));
 sg13g2_dfrbp_1 \proj_14.flop22/_1_  (.CLK(clknet_5_24__leaf_clk_regs),
    .RESET_B(net341),
    .D(\proj_14.net76 ),
    .Q_N(\proj_14.flop22/notq ),
    .Q(\proj_14.net75 ));
 sg13g2_tiehi \proj_14.flop23/_1__296  (.L_HI(net342));
 sg13g2_dfrbp_1 \proj_14.flop23/_1_  (.CLK(clknet_5_7__leaf_clk_regs),
    .RESET_B(net342),
    .D(\proj_14.net79 ),
    .Q_N(\proj_14.flop23/notq ),
    .Q(\proj_14.net78 ));
 sg13g2_tiehi \proj_14.flop24/_1__297  (.L_HI(net343));
 sg13g2_dfrbp_1 \proj_14.flop24/_1_  (.CLK(clknet_5_7__leaf_clk_regs),
    .RESET_B(net343),
    .D(\proj_14.net82 ),
    .Q_N(\proj_14.flop24/notq ),
    .Q(\proj_14.net81 ));
 sg13g2_tiehi \proj_14.flop25/_1__298  (.L_HI(net344));
 sg13g2_dfrbp_1 \proj_14.flop25/_1_  (.CLK(clknet_5_13__leaf_clk_regs),
    .RESET_B(net344),
    .D(\proj_14.net85 ),
    .Q_N(\proj_14.flop25/notq ),
    .Q(\proj_14.net84 ));
 sg13g2_tiehi \proj_14.flop26/_1__299  (.L_HI(net345));
 sg13g2_dfrbp_1 \proj_14.flop26/_1_  (.CLK(clknet_5_13__leaf_clk_regs),
    .RESET_B(net345),
    .D(\proj_14.net88 ),
    .Q_N(\proj_14.flop26/notq ),
    .Q(\proj_14.net87 ));
 sg13g2_tiehi \proj_14.flop27/_1__300  (.L_HI(net346));
 sg13g2_dfrbp_1 \proj_14.flop27/_1_  (.CLK(clknet_5_12__leaf_clk_regs),
    .RESET_B(net346),
    .D(\proj_14.net91 ),
    .Q_N(\proj_14.flop27/notq ),
    .Q(\proj_14.net90 ));
 sg13g2_tiehi \proj_14.flop28/_1__301  (.L_HI(net347));
 sg13g2_dfrbp_1 \proj_14.flop28/_1_  (.CLK(clknet_5_12__leaf_clk_regs),
    .RESET_B(net347),
    .D(\proj_14.net94 ),
    .Q_N(\proj_14.flop28/notq ),
    .Q(\proj_14.net93 ));
 sg13g2_tiehi \proj_14.flop29/_1__302  (.L_HI(net348));
 sg13g2_dfrbp_1 \proj_14.flop29/_1_  (.CLK(clknet_5_13__leaf_clk_regs),
    .RESET_B(net348),
    .D(\proj_14.net97 ),
    .Q_N(\proj_14.flop29/notq ),
    .Q(\proj_14.net96 ));
 sg13g2_tiehi \proj_14.flop3/_1__303  (.L_HI(net349));
 sg13g2_dfrbp_1 \proj_14.flop3/_1_  (.CLK(clknet_5_14__leaf_clk_regs),
    .RESET_B(net349),
    .D(\proj_14.net12 ),
    .Q_N(\proj_14.flop3/notq ),
    .Q(\proj_14.net11 ));
 sg13g2_tiehi \proj_14.flop30/_1__304  (.L_HI(net350));
 sg13g2_dfrbp_1 \proj_14.flop30/_1_  (.CLK(clknet_5_26__leaf_clk_regs),
    .RESET_B(net350),
    .D(\proj_14.net100 ),
    .Q_N(\proj_14.flop30/notq ),
    .Q(\proj_14.net99 ));
 sg13g2_tiehi \proj_14.flop31/_1__305  (.L_HI(net351));
 sg13g2_dfrbp_1 \proj_14.flop31/_1_  (.CLK(clknet_5_24__leaf_clk_regs),
    .RESET_B(net351),
    .D(\proj_14.net103 ),
    .Q_N(\proj_14.flop31/notq ),
    .Q(\proj_14.net102 ));
 sg13g2_tiehi \proj_14.flop32/_1__306  (.L_HI(net352));
 sg13g2_dfrbp_1 \proj_14.flop32/_1_  (.CLK(clknet_5_25__leaf_clk_regs),
    .RESET_B(net352),
    .D(\proj_14.net106 ),
    .Q_N(\proj_14.flop32/notq ),
    .Q(\proj_14.net105 ));
 sg13g2_tiehi \proj_14.flop33/_1__307  (.L_HI(net353));
 sg13g2_dfrbp_1 \proj_14.flop33/_1_  (.CLK(clknet_5_27__leaf_clk_regs),
    .RESET_B(net353),
    .D(\proj_14.net109 ),
    .Q_N(\proj_14.flop33/notq ),
    .Q(\proj_14.net108 ));
 sg13g2_tiehi \proj_14.flop34/_1__308  (.L_HI(net354));
 sg13g2_dfrbp_1 \proj_14.flop34/_1_  (.CLK(clknet_5_27__leaf_clk_regs),
    .RESET_B(net354),
    .D(\proj_14.net112 ),
    .Q_N(\proj_14.flop34/notq ),
    .Q(\proj_14.net111 ));
 sg13g2_tiehi \proj_14.flop35/_1__309  (.L_HI(net355));
 sg13g2_dfrbp_1 \proj_14.flop35/_1_  (.CLK(clknet_5_8__leaf_clk_regs),
    .RESET_B(net355),
    .D(\proj_14.net116 ),
    .Q_N(\proj_14.flop35/notq ),
    .Q(\proj_14.net59 ));
 sg13g2_tiehi \proj_14.flop36/_1__310  (.L_HI(net356));
 sg13g2_dfrbp_1 \proj_14.flop36/_1_  (.CLK(clknet_5_9__leaf_clk_regs),
    .RESET_B(net356),
    .D(\proj_14.net119 ),
    .Q_N(\proj_14.flop36/notq ),
    .Q(\proj_14.net118 ));
 sg13g2_tiehi \proj_14.flop37/_1__311  (.L_HI(net357));
 sg13g2_dfrbp_1 \proj_14.flop37/_1_  (.CLK(clknet_5_8__leaf_clk_regs),
    .RESET_B(net357),
    .D(\proj_14.net122 ),
    .Q_N(\proj_14.flop37/notq ),
    .Q(\proj_14.net121 ));
 sg13g2_tiehi \proj_14.flop38/_1__312  (.L_HI(net358));
 sg13g2_dfrbp_1 \proj_14.flop38/_1_  (.CLK(clknet_5_2__leaf_clk_regs),
    .RESET_B(net358),
    .D(\proj_14.net125 ),
    .Q_N(\proj_14.flop38/notq ),
    .Q(\proj_14.net124 ));
 sg13g2_tiehi \proj_14.flop39/_1__313  (.L_HI(net359));
 sg13g2_dfrbp_1 \proj_14.flop39/_1_  (.CLK(clknet_5_26__leaf_clk_regs),
    .RESET_B(net359),
    .D(\proj_14.net127 ),
    .Q_N(\proj_14.flop39/notq ),
    .Q(\proj_14.net128 ));
 sg13g2_tiehi \proj_14.flop4/_1__314  (.L_HI(net360));
 sg13g2_dfrbp_1 \proj_14.flop4/_1_  (.CLK(clknet_5_12__leaf_clk_regs),
    .RESET_B(net360),
    .D(\proj_14.net15 ),
    .Q_N(\proj_14.flop4/notq ),
    .Q(\proj_14.net14 ));
 sg13g2_tiehi \proj_14.flop40/_1__315  (.L_HI(net361));
 sg13g2_dfrbp_1 \proj_14.flop40/_1_  (.CLK(clknet_5_26__leaf_clk_regs),
    .RESET_B(net361),
    .D(\proj_14.net131 ),
    .Q_N(\proj_14.flop40/notq ),
    .Q(\proj_14.net130 ));
 sg13g2_tiehi \proj_14.flop41/_1__316  (.L_HI(net362));
 sg13g2_dfrbp_1 \proj_14.flop41/_1_  (.CLK(clknet_5_15__leaf_clk_regs),
    .RESET_B(net362),
    .D(\proj_14.net134 ),
    .Q_N(\proj_14.flop41/notq ),
    .Q(\proj_14.net133 ));
 sg13g2_tiehi \proj_14.flop42/_1__317  (.L_HI(net363));
 sg13g2_dfrbp_1 \proj_14.flop42/_1_  (.CLK(clknet_5_15__leaf_clk_regs),
    .RESET_B(net363),
    .D(\proj_14.net137 ),
    .Q_N(\proj_14.flop42/notq ),
    .Q(\proj_14.net136 ));
 sg13g2_tiehi \proj_14.flop43/_1__318  (.L_HI(net364));
 sg13g2_dfrbp_1 \proj_14.flop43/_1_  (.CLK(clknet_5_30__leaf_clk_regs),
    .RESET_B(net364),
    .D(\proj_14.net139 ),
    .Q_N(\proj_14.flop43/notq ),
    .Q(\proj_14.net140 ));
 sg13g2_tiehi \proj_14.flop44/_1__319  (.L_HI(net365));
 sg13g2_dfrbp_1 \proj_14.flop44/_1_  (.CLK(clknet_5_30__leaf_clk_regs),
    .RESET_B(net365),
    .D(\proj_14.net143 ),
    .Q_N(\proj_14.flop44/notq ),
    .Q(\proj_14.net142 ));
 sg13g2_tiehi \proj_14.flop45/_1__320  (.L_HI(net366));
 sg13g2_dfrbp_1 \proj_14.flop45/_1_  (.CLK(clknet_5_31__leaf_clk_regs),
    .RESET_B(net366),
    .D(\proj_14.net146 ),
    .Q_N(\proj_14.flop45/notq ),
    .Q(\proj_14.net145 ));
 sg13g2_tiehi \proj_14.flop46/_1__321  (.L_HI(net367));
 sg13g2_dfrbp_1 \proj_14.flop46/_1_  (.CLK(clknet_5_30__leaf_clk_regs),
    .RESET_B(net367),
    .D(\proj_14.net149 ),
    .Q_N(\proj_14.flop46/notq ),
    .Q(\proj_14.net148 ));
 sg13g2_tiehi \proj_14.flop47/_1__322  (.L_HI(net368));
 sg13g2_dfrbp_1 \proj_14.flop47/_1_  (.CLK(clknet_5_31__leaf_clk_regs),
    .RESET_B(net368),
    .D(\proj_14.net152 ),
    .Q_N(\proj_14.flop47/notq ),
    .Q(\proj_14.net151 ));
 sg13g2_tiehi \proj_14.flop48/_1__323  (.L_HI(net369));
 sg13g2_dfrbp_1 \proj_14.flop48/_1_  (.CLK(clknet_5_30__leaf_clk_regs),
    .RESET_B(net369),
    .D(\proj_14.net155 ),
    .Q_N(\proj_14.flop48/notq ),
    .Q(\proj_14.net154 ));
 sg13g2_tiehi \proj_14.flop49/_1__324  (.L_HI(net370));
 sg13g2_dfrbp_1 \proj_14.flop49/_1_  (.CLK(clknet_5_31__leaf_clk_regs),
    .RESET_B(net370),
    .D(\proj_14.net158 ),
    .Q_N(\proj_14.flop49/notq ),
    .Q(\proj_14.net157 ));
 sg13g2_tiehi \proj_14.flop5/_1__325  (.L_HI(net371));
 sg13g2_dfrbp_1 \proj_14.flop5/_1_  (.CLK(clknet_5_11__leaf_clk_regs),
    .RESET_B(net371),
    .D(\proj_14.net18 ),
    .Q_N(\proj_14.flop5/notq ),
    .Q(\proj_14.net17 ));
 sg13g2_tiehi \proj_14.flop50/_1__326  (.L_HI(net372));
 sg13g2_dfrbp_1 \proj_14.flop50/_1_  (.CLK(clknet_5_30__leaf_clk_regs),
    .RESET_B(net372),
    .D(\proj_14.net161 ),
    .Q_N(\proj_14.flop50/notq ),
    .Q(\proj_14.net160 ));
 sg13g2_tiehi \proj_14.flop51/_1__327  (.L_HI(net373));
 sg13g2_dfrbp_1 \proj_14.flop51/_1_  (.CLK(clknet_5_29__leaf_clk_regs),
    .RESET_B(net373),
    .D(\proj_14.net164 ),
    .Q_N(\proj_14.flop51/notq ),
    .Q(\proj_14.net163 ));
 sg13g2_tiehi \proj_14.flop52/_1__328  (.L_HI(net374));
 sg13g2_dfrbp_1 \proj_14.flop52/_1_  (.CLK(clknet_5_29__leaf_clk_regs),
    .RESET_B(net374),
    .D(\proj_14.net167 ),
    .Q_N(\proj_14.flop52/notq ),
    .Q(\proj_14.net166 ));
 sg13g2_tiehi \proj_14.flop53/_1__329  (.L_HI(net375));
 sg13g2_dfrbp_1 \proj_14.flop53/_1_  (.CLK(clknet_5_29__leaf_clk_regs),
    .RESET_B(net375),
    .D(\proj_14.net170 ),
    .Q_N(\proj_14.flop53/notq ),
    .Q(\proj_14.net169 ));
 sg13g2_tiehi \proj_14.flop54/_1__330  (.L_HI(net376));
 sg13g2_dfrbp_1 \proj_14.flop54/_1_  (.CLK(clknet_5_29__leaf_clk_regs),
    .RESET_B(net376),
    .D(\proj_14.net173 ),
    .Q_N(\proj_14.flop54/notq ),
    .Q(\proj_14.net172 ));
 sg13g2_tiehi \proj_14.flop55/_1__331  (.L_HI(net377));
 sg13g2_dfrbp_1 \proj_14.flop55/_1_  (.CLK(clknet_5_28__leaf_clk_regs),
    .RESET_B(net377),
    .D(\proj_14.net176 ),
    .Q_N(\proj_14.flop55/notq ),
    .Q(\proj_14.net175 ));
 sg13g2_tiehi \proj_14.flop56/_1__332  (.L_HI(net378));
 sg13g2_dfrbp_1 \proj_14.flop56/_1_  (.CLK(clknet_5_22__leaf_clk_regs),
    .RESET_B(net378),
    .D(\proj_14.net179 ),
    .Q_N(\proj_14.flop56/notq ),
    .Q(\proj_14.net178 ));
 sg13g2_tiehi \proj_14.flop57/_1__333  (.L_HI(net379));
 sg13g2_dfrbp_1 \proj_14.flop57/_1_  (.CLK(clknet_5_22__leaf_clk_regs),
    .RESET_B(net379),
    .D(\proj_14.net182 ),
    .Q_N(\proj_14.flop57/notq ),
    .Q(\proj_14.net181 ));
 sg13g2_tiehi \proj_14.flop58/_1__334  (.L_HI(net380));
 sg13g2_dfrbp_1 \proj_14.flop58/_1_  (.CLK(clknet_5_23__leaf_clk_regs),
    .RESET_B(net380),
    .D(\proj_14.net185 ),
    .Q_N(\proj_14.flop58/notq ),
    .Q(\proj_14.net184 ));
 sg13g2_tiehi \proj_14.flop59/_1__335  (.L_HI(net381));
 sg13g2_dfrbp_1 \proj_14.flop59/_1_  (.CLK(clknet_5_20__leaf_clk_regs),
    .RESET_B(net381),
    .D(\proj_14.net188 ),
    .Q_N(\proj_14.flop59/notq ),
    .Q(\proj_14.net187 ));
 sg13g2_tiehi \proj_14.flop6/_1__336  (.L_HI(net382));
 sg13g2_dfrbp_1 \proj_14.flop6/_1_  (.CLK(clknet_5_9__leaf_clk_regs),
    .RESET_B(net382),
    .D(\proj_14.net21 ),
    .Q_N(\proj_14.flop6/notq ),
    .Q(\proj_14.net20 ));
 sg13g2_tiehi \proj_14.flop60/_1__337  (.L_HI(net383));
 sg13g2_dfrbp_1 \proj_14.flop60/_1_  (.CLK(clknet_5_28__leaf_clk_regs),
    .RESET_B(net383),
    .D(\proj_14.net192 ),
    .Q_N(\proj_14.flop60/notq ),
    .Q(\proj_14.net114 ));
 sg13g2_tiehi \proj_14.flop61/_1__338  (.L_HI(net384));
 sg13g2_dfrbp_1 \proj_14.flop61/_1_  (.CLK(clknet_5_30__leaf_clk_regs),
    .RESET_B(net384),
    .D(\proj_14.net195 ),
    .Q_N(\proj_14.flop61/notq ),
    .Q(\proj_14.net194 ));
 sg13g2_tiehi \proj_14.flop62/_1__339  (.L_HI(net385));
 sg13g2_dfrbp_1 \proj_14.flop62/_1_  (.CLK(clknet_5_31__leaf_clk_regs),
    .RESET_B(net385),
    .D(\proj_14.net198 ),
    .Q_N(\proj_14.flop62/notq ),
    .Q(\proj_14.net197 ));
 sg13g2_tiehi \proj_14.flop63/_1__340  (.L_HI(net386));
 sg13g2_dfrbp_1 \proj_14.flop63/_1_  (.CLK(clknet_5_31__leaf_clk_regs),
    .RESET_B(net386),
    .D(\proj_14.net201 ),
    .Q_N(\proj_14.flop63/notq ),
    .Q(\proj_14.net200 ));
 sg13g2_tiehi \proj_14.flop64/_1__341  (.L_HI(net387));
 sg13g2_dfrbp_1 \proj_14.flop64/_1_  (.CLK(clknet_5_16__leaf_clk_regs),
    .RESET_B(net387),
    .D(\proj_14.net203 ),
    .Q_N(\proj_14.flop64/notq ),
    .Q(\proj_14.net204 ));
 sg13g2_tiehi \proj_14.flop65/_1__342  (.L_HI(net388));
 sg13g2_dfrbp_1 \proj_14.flop65/_1_  (.CLK(clknet_5_19__leaf_clk_regs),
    .RESET_B(net388),
    .D(\proj_14.net207 ),
    .Q_N(\proj_14.flop65/notq ),
    .Q(\proj_14.net206 ));
 sg13g2_tiehi \proj_14.flop66/_1__343  (.L_HI(net389));
 sg13g2_dfrbp_1 \proj_14.flop66/_1_  (.CLK(clknet_5_18__leaf_clk_regs),
    .RESET_B(net389),
    .D(\proj_14.net210 ),
    .Q_N(\proj_14.flop66/notq ),
    .Q(\proj_14.net209 ));
 sg13g2_tiehi \proj_14.flop67/_1__344  (.L_HI(net390));
 sg13g2_dfrbp_1 \proj_14.flop67/_1_  (.CLK(clknet_5_18__leaf_clk_regs),
    .RESET_B(net390),
    .D(\proj_14.net213 ),
    .Q_N(\proj_14.flop67/notq ),
    .Q(\proj_14.net212 ));
 sg13g2_tiehi \proj_14.flop68/_1__345  (.L_HI(net391));
 sg13g2_dfrbp_1 \proj_14.flop68/_1_  (.CLK(clknet_5_5__leaf_clk_regs),
    .RESET_B(net391),
    .D(\proj_14.net216 ),
    .Q_N(\proj_14.flop68/notq ),
    .Q(\proj_14.net215 ));
 sg13g2_tiehi \proj_14.flop69/_1__346  (.L_HI(net392));
 sg13g2_dfrbp_1 \proj_14.flop69/_1_  (.CLK(clknet_5_16__leaf_clk_regs),
    .RESET_B(net392),
    .D(\proj_14.net219 ),
    .Q_N(\proj_14.flop69/notq ),
    .Q(\proj_14.net218 ));
 sg13g2_tiehi \proj_14.flop7/_1__347  (.L_HI(net393));
 sg13g2_dfrbp_1 \proj_14.flop7/_1_  (.CLK(clknet_5_9__leaf_clk_regs),
    .RESET_B(net393),
    .D(\proj_14.net24 ),
    .Q_N(\proj_14.flop7/notq ),
    .Q(\proj_14.net23 ));
 sg13g2_tiehi \proj_14.flop70/_1__348  (.L_HI(net394));
 sg13g2_dfrbp_1 \proj_14.flop70/_1_  (.CLK(clknet_5_16__leaf_clk_regs),
    .RESET_B(net394),
    .D(\proj_14.net222 ),
    .Q_N(\proj_14.flop70/notq ),
    .Q(\proj_14.net221 ));
 sg13g2_tiehi \proj_14.flop71/_1__349  (.L_HI(net395));
 sg13g2_dfrbp_1 \proj_14.flop71/_1_  (.CLK(clknet_5_5__leaf_clk_regs),
    .RESET_B(net395),
    .D(\proj_14.net225 ),
    .Q_N(\proj_14.flop71/notq ),
    .Q(\proj_14.net224 ));
 sg13g2_tiehi \proj_14.flop72/_1__350  (.L_HI(net396));
 sg13g2_dfrbp_1 \proj_14.flop72/_1_  (.CLK(clknet_5_4__leaf_clk_regs),
    .RESET_B(net396),
    .D(\proj_14.net228 ),
    .Q_N(\proj_14.flop72/notq ),
    .Q(\proj_14.net227 ));
 sg13g2_tiehi \proj_14.flop73/_1__351  (.L_HI(net397));
 sg13g2_dfrbp_1 \proj_14.flop73/_1_  (.CLK(clknet_5_4__leaf_clk_regs),
    .RESET_B(net397),
    .D(\proj_14.net231 ),
    .Q_N(\proj_14.flop73/notq ),
    .Q(\proj_14.net230 ));
 sg13g2_tiehi \proj_14.flop74/_1__352  (.L_HI(net398));
 sg13g2_dfrbp_1 \proj_14.flop74/_1_  (.CLK(clknet_5_1__leaf_clk_regs),
    .RESET_B(net398),
    .D(\proj_14.net234 ),
    .Q_N(\proj_14.flop74/notq ),
    .Q(\proj_14.net233 ));
 sg13g2_tiehi \proj_14.flop75/_1__353  (.L_HI(net399));
 sg13g2_dfrbp_1 \proj_14.flop75/_1_  (.CLK(clknet_5_1__leaf_clk_regs),
    .RESET_B(net399),
    .D(\proj_14.net237 ),
    .Q_N(\proj_14.flop75/notq ),
    .Q(\proj_14.net236 ));
 sg13g2_tiehi \proj_14.flop76/_1__354  (.L_HI(net400));
 sg13g2_dfrbp_1 \proj_14.flop76/_1_  (.CLK(clknet_5_4__leaf_clk_regs),
    .RESET_B(net400),
    .D(\proj_14.net240 ),
    .Q_N(\proj_14.flop76/notq ),
    .Q(\proj_14.net239 ));
 sg13g2_tiehi \proj_14.flop77/_1__355  (.L_HI(net401));
 sg13g2_dfrbp_1 \proj_14.flop77/_1_  (.CLK(clknet_5_5__leaf_clk_regs),
    .RESET_B(net401),
    .D(\proj_14.net243 ),
    .Q_N(\proj_14.flop77/notq ),
    .Q(\proj_14.net242 ));
 sg13g2_tiehi \proj_14.flop78/_1__356  (.L_HI(net402));
 sg13g2_dfrbp_1 \proj_14.flop78/_1_  (.CLK(clknet_5_4__leaf_clk_regs),
    .RESET_B(net402),
    .D(\proj_14.net246 ),
    .Q_N(\proj_14.flop78/notq ),
    .Q(\proj_14.net245 ));
 sg13g2_tiehi \proj_14.flop79/_1__357  (.L_HI(net403));
 sg13g2_dfrbp_1 \proj_14.flop79/_1_  (.CLK(clknet_5_16__leaf_clk_regs),
    .RESET_B(net403),
    .D(\proj_14.net249 ),
    .Q_N(\proj_14.flop79/notq ),
    .Q(\proj_14.net248 ));
 sg13g2_tiehi \proj_14.flop8/_1__358  (.L_HI(net404));
 sg13g2_dfrbp_1 \proj_14.flop8/_1_  (.CLK(clknet_5_10__leaf_clk_regs),
    .RESET_B(net404),
    .D(\proj_14.net27 ),
    .Q_N(\proj_14.flop8/notq ),
    .Q(\proj_14.net26 ));
 sg13g2_tiehi \proj_14.flop80/_1__359  (.L_HI(net405));
 sg13g2_dfrbp_1 \proj_14.flop80/_1_  (.CLK(clknet_5_16__leaf_clk_regs),
    .RESET_B(net405),
    .D(\proj_14.net252 ),
    .Q_N(\proj_14.flop80/notq ),
    .Q(\proj_14.net251 ));
 sg13g2_tiehi \proj_14.flop81/_1__360  (.L_HI(net406));
 sg13g2_dfrbp_1 \proj_14.flop81/_1_  (.CLK(clknet_5_17__leaf_clk_regs),
    .RESET_B(net406),
    .D(\proj_14.net256 ),
    .Q_N(\proj_14.flop81/notq ),
    .Q(\proj_14.net190 ));
 sg13g2_tiehi \proj_14.flop82/_1__361  (.L_HI(net407));
 sg13g2_dfrbp_1 \proj_14.flop82/_1_  (.CLK(clknet_5_20__leaf_clk_regs),
    .RESET_B(net407),
    .D(\proj_14.net259 ),
    .Q_N(\proj_14.flop82/notq ),
    .Q(\proj_14.net258 ));
 sg13g2_tiehi \proj_14.flop83/_1__362  (.L_HI(net408));
 sg13g2_dfrbp_1 \proj_14.flop83/_1_  (.CLK(clknet_5_17__leaf_clk_regs),
    .RESET_B(net408),
    .D(\proj_14.net262 ),
    .Q_N(\proj_14.flop83/notq ),
    .Q(\proj_14.net261 ));
 sg13g2_tiehi \proj_14.flop84/_1__363  (.L_HI(net409));
 sg13g2_dfrbp_1 \proj_14.flop84/_1_  (.CLK(clknet_5_17__leaf_clk_regs),
    .RESET_B(net409),
    .D(\proj_14.net265 ),
    .Q_N(\proj_14.flop84/notq ),
    .Q(\proj_14.net264 ));
 sg13g2_tiehi \proj_14.flop85/_1__364  (.L_HI(net410));
 sg13g2_dfrbp_1 \proj_14.flop85/_1_  (.CLK(clknet_5_17__leaf_clk_regs),
    .RESET_B(net410),
    .D(\proj_14.net267 ),
    .Q_N(\proj_14.flop85/notq ),
    .Q(\proj_14.net268 ));
 sg13g2_tiehi \proj_14.flop86/_1__365  (.L_HI(net411));
 sg13g2_dfrbp_1 \proj_14.flop86/_1_  (.CLK(clknet_5_16__leaf_clk_regs),
    .RESET_B(net411),
    .D(\proj_14.net271 ),
    .Q_N(\proj_14.flop86/notq ),
    .Q(\proj_14.net270 ));
 sg13g2_tiehi \proj_14.flop87/_1__366  (.L_HI(net412));
 sg13g2_dfrbp_1 \proj_14.flop87/_1_  (.CLK(clknet_5_20__leaf_clk_regs),
    .RESET_B(net412),
    .D(\proj_14.net274 ),
    .Q_N(\proj_14.flop87/notq ),
    .Q(\proj_14.net273 ));
 sg13g2_tiehi \proj_14.flop88/_1__367  (.L_HI(net413));
 sg13g2_dfrbp_1 \proj_14.flop88/_1_  (.CLK(clknet_5_20__leaf_clk_regs),
    .RESET_B(net413),
    .D(\proj_14.net277 ),
    .Q_N(\proj_14.flop88/notq ),
    .Q(\proj_14.net276 ));
 sg13g2_tiehi \proj_14.flop89/_1__368  (.L_HI(net414));
 sg13g2_dfrbp_1 \proj_14.flop89/_1_  (.CLK(clknet_5_20__leaf_clk_regs),
    .RESET_B(net414),
    .D(\proj_14.net280 ),
    .Q_N(\proj_14.flop89/notq ),
    .Q(\proj_14.net279 ));
 sg13g2_tiehi \proj_14.flop9/_1__369  (.L_HI(net415));
 sg13g2_dfrbp_1 \proj_14.flop9/_1_  (.CLK(clknet_5_10__leaf_clk_regs),
    .RESET_B(net415),
    .D(\proj_14.net30 ),
    .Q_N(\proj_14.flop9/notq ),
    .Q(\proj_14.net29 ));
 sg13g2_tiehi \proj_14.flop90/_1__370  (.L_HI(net416));
 sg13g2_dfrbp_1 \proj_14.flop90/_1_  (.CLK(clknet_5_20__leaf_clk_regs),
    .RESET_B(net416),
    .D(\proj_14.net283 ),
    .Q_N(\proj_14.flop90/notq ),
    .Q(\proj_14.net282 ));
 sg13g2_tiehi \proj_14.flop91/_1__371  (.L_HI(net417));
 sg13g2_dfrbp_1 \proj_14.flop91/_1_  (.CLK(clknet_5_21__leaf_clk_regs),
    .RESET_B(net417),
    .D(\proj_14.net286 ),
    .Q_N(\proj_14.flop91/notq ),
    .Q(\proj_14.net285 ));
 sg13g2_tiehi \proj_14.flop92/_1__372  (.L_HI(net418));
 sg13g2_dfrbp_1 \proj_14.flop92/_1_  (.CLK(clknet_5_21__leaf_clk_regs),
    .RESET_B(net418),
    .D(\proj_14.net289 ),
    .Q_N(\proj_14.flop92/notq ),
    .Q(\proj_14.net288 ));
 sg13g2_tiehi \proj_14.flop93/_1__373  (.L_HI(net419));
 sg13g2_dfrbp_1 \proj_14.flop93/_1_  (.CLK(clknet_5_21__leaf_clk_regs),
    .RESET_B(net419),
    .D(\proj_14.net292 ),
    .Q_N(\proj_14.flop93/notq ),
    .Q(\proj_14.net291 ));
 sg13g2_tiehi \proj_14.flop94/_1__374  (.L_HI(net420));
 sg13g2_dfrbp_1 \proj_14.flop94/_1_  (.CLK(clknet_5_23__leaf_clk_regs),
    .RESET_B(net420),
    .D(\proj_14.net295 ),
    .Q_N(\proj_14.flop94/notq ),
    .Q(\proj_14.net294 ));
 sg13g2_tiehi \proj_14.flop95/_1__375  (.L_HI(net421));
 sg13g2_dfrbp_1 \proj_14.flop95/_1_  (.CLK(clknet_5_21__leaf_clk_regs),
    .RESET_B(net421),
    .D(\proj_14.net298 ),
    .Q_N(\proj_14.flop95/notq ),
    .Q(\proj_14.net297 ));
 sg13g2_tiehi \proj_14.flop96/_1__376  (.L_HI(net422));
 sg13g2_dfrbp_1 \proj_14.flop96/_1_  (.CLK(clknet_5_23__leaf_clk_regs),
    .RESET_B(net422),
    .D(\proj_14.net301 ),
    .Q_N(\proj_14.flop96/notq ),
    .Q(\proj_14.net300 ));
 sg13g2_tiehi \proj_14.flop97/_1__377  (.L_HI(net423));
 sg13g2_dfrbp_1 \proj_14.flop97/_1_  (.CLK(clknet_5_21__leaf_clk_regs),
    .RESET_B(net423),
    .D(\proj_14.net304 ),
    .Q_N(\proj_14.flop97/notq ),
    .Q(\proj_14.net303 ));
 sg13g2_tiehi \proj_14.flop98/_1__378  (.L_HI(net424));
 sg13g2_dfrbp_1 \proj_14.flop98/_1_  (.CLK(clknet_5_21__leaf_clk_regs),
    .RESET_B(net424),
    .D(\proj_14.net307 ),
    .Q_N(\proj_14.flop98/notq ),
    .Q(\proj_14.net306 ));
 sg13g2_tiehi \proj_14.flop99/_1__379  (.L_HI(net425));
 sg13g2_dfrbp_1 \proj_14.flop99/_1_  (.CLK(clknet_5_23__leaf_clk_regs),
    .RESET_B(net425),
    .D(\proj_14.net310 ),
    .Q_N(\proj_14.flop99/notq ),
    .Q(\proj_14.net309 ));
 sg13g2_inv_1 \proj_12.not1/_0__1  (.Y(net426),
    .A(\proj_12.net22 ));
 sg13g2_mux2_1 \proj_14.mux1/_0_  (.A0(net77),
    .A1(net589),
    .S(net150),
    .X(\proj_14.net8 ));
 sg13g2_mux2_1 \proj_14.mux10/_0_  (.A0(net13),
    .A1(net554),
    .S(net149),
    .X(\proj_14.net33 ));
 sg13g2_mux2_1 \proj_14.mux100/_0_  (.A0(net78),
    .A1(net548),
    .S(net161),
    .X(\proj_14.net310 ));
 sg13g2_mux2_1 \proj_14.mux101/_0_  (.A0(net79),
    .A1(net486),
    .S(net161),
    .X(\proj_14.net313 ));
 sg13g2_mux2_1 \proj_14.mux102/_0_  (.A0(net80),
    .A1(net522),
    .S(net161),
    .X(\proj_14.net316 ));
 sg13g2_mux2_1 \proj_14.mux103/_0_  (.A0(net81),
    .A1(net562),
    .S(net142),
    .X(\proj_14.net320 ));
 sg13g2_mux2_1 \proj_14.mux104/_0_  (.A0(net82),
    .A1(net600),
    .S(net154),
    .X(\proj_14.net323 ));
 sg13g2_mux2_1 \proj_14.mux105/_0_  (.A0(net83),
    .A1(net549),
    .S(net154),
    .X(\proj_14.net326 ));
 sg13g2_mux2_1 \proj_14.mux106/_0_  (.A0(net84),
    .A1(net505),
    .S(net154),
    .X(\proj_14.net329 ));
 sg13g2_mux2_1 \proj_14.mux107/_0_  (.A0(net85),
    .A1(net547),
    .S(net156),
    .X(\proj_14.net332 ));
 sg13g2_mux2_1 \proj_14.mux108/_0_  (.A0(net86),
    .A1(net469),
    .S(net156),
    .X(\proj_14.net336 ));
 sg13g2_mux2_1 \proj_14.mux109/_0_  (.A0(net87),
    .A1(net489),
    .S(net155),
    .X(\proj_14.net339 ));
 sg13g2_mux2_1 \proj_14.mux11/_0_  (.A0(net88),
    .A1(net454),
    .S(net148),
    .X(\proj_14.net36 ));
 sg13g2_mux2_1 \proj_14.mux110/_0_  (.A0(net89),
    .A1(net509),
    .S(net155),
    .X(\proj_14.net342 ));
 sg13g2_mux2_1 \proj_14.mux111/_0_  (.A0(net14),
    .A1(net526),
    .S(net155),
    .X(\proj_14.net345 ));
 sg13g2_mux2_1 \proj_14.mux112/_0_  (.A0(net90),
    .A1(net525),
    .S(net163),
    .X(\proj_14.net348 ));
 sg13g2_mux2_1 \proj_14.mux113/_0_  (.A0(net15),
    .A1(net559),
    .S(net163),
    .X(\proj_14.net351 ));
 sg13g2_mux2_1 \proj_14.mux114/_0_  (.A0(net16),
    .A1(net560),
    .S(net163),
    .X(\proj_14.net354 ));
 sg13g2_mux2_1 \proj_14.mux115/_0_  (.A0(net17),
    .A1(net521),
    .S(net165),
    .X(\proj_14.net357 ));
 sg13g2_mux2_1 \proj_14.mux116/_0_  (.A0(net18),
    .A1(net602),
    .S(net165),
    .X(\proj_14.net360 ));
 sg13g2_mux2_1 \proj_14.mux117/_0_  (.A0(net19),
    .A1(net442),
    .S(net165),
    .X(\proj_14.net363 ));
 sg13g2_mux2_1 \proj_14.mux118/_0_  (.A0(net91),
    .A1(net594),
    .S(net160),
    .X(\proj_14.net366 ));
 sg13g2_mux2_1 \proj_14.mux119/_0_  (.A0(net20),
    .A1(net440),
    .S(net160),
    .X(\proj_14.net369 ));
 sg13g2_mux2_1 \proj_14.mux12/_0_  (.A0(net21),
    .A1(net496),
    .S(net148),
    .X(\proj_14.net39 ));
 sg13g2_mux2_1 \proj_14.mux120/_0_  (.A0(net92),
    .A1(net479),
    .S(net155),
    .X(\proj_14.net372 ));
 sg13g2_mux2_1 \proj_14.mux121/_0_  (.A0(net93),
    .A1(net561),
    .S(net155),
    .X(\proj_14.net375 ));
 sg13g2_mux2_1 \proj_14.mux122/_0_  (.A0(net94),
    .A1(net537),
    .S(net156),
    .X(\proj_14.net378 ));
 sg13g2_mux2_1 \proj_14.mux123/_0_  (.A0(net95),
    .A1(net482),
    .S(net155),
    .X(\proj_14.net381 ));
 sg13g2_mux2_1 \proj_14.mux124/_0_  (.A0(net96),
    .A1(net467),
    .S(net161),
    .X(\proj_14.net385 ));
 sg13g2_mux2_1 \proj_14.mux125/_0_  (.A0(net97),
    .A1(net593),
    .S(net160),
    .X(\proj_14.net388 ));
 sg13g2_mux2_1 \proj_14.mux126/_0_  (.A0(net98),
    .A1(net520),
    .S(net160),
    .X(\proj_14.net391 ));
 sg13g2_mux2_1 \proj_14.mux127/_0_  (.A0(net99),
    .A1(net439),
    .S(net156),
    .X(\proj_14.net394 ));
 sg13g2_mux2_1 \proj_14.mux128/_0_  (.A0(net100),
    .A1(net514),
    .S(net143),
    .X(\proj_14.net396 ));
 sg13g2_mux2_1 \proj_14.mux129/_0_  (.A0(net101),
    .A1(net563),
    .S(net143),
    .X(\proj_14.net400 ));
 sg13g2_mux2_1 \proj_14.mux13/_0_  (.A0(net102),
    .A1(net550),
    .S(net148),
    .X(\proj_14.net42 ));
 sg13g2_mux2_1 \proj_14.mux130/_0_  (.A0(net103),
    .A1(net462),
    .S(net143),
    .X(\proj_14.net403 ));
 sg13g2_mux2_1 \proj_14.mux131/_0_  (.A0(net104),
    .A1(net506),
    .S(net143),
    .X(\proj_14.net406 ));
 sg13g2_mux2_1 \proj_14.mux132/_0_  (.A0(net22),
    .A1(net478),
    .S(net139),
    .X(\proj_14.net409 ));
 sg13g2_mux2_1 \proj_14.mux133/_0_  (.A0(net105),
    .A1(net452),
    .S(net140),
    .X(\proj_14.net412 ));
 sg13g2_mux2_1 \proj_14.mux134/_0_  (.A0(net23),
    .A1(net599),
    .S(net140),
    .X(\proj_14.net415 ));
 sg13g2_mux2_1 \proj_14.mux135/_0_  (.A0(net24),
    .A1(net508),
    .S(net138),
    .X(\proj_14.net418 ));
 sg13g2_mux2_1 \proj_14.mux136/_0_  (.A0(net106),
    .A1(net524),
    .S(net138),
    .X(\proj_14.net421 ));
 sg13g2_mux2_1 \proj_14.mux137/_0_  (.A0(net25),
    .A1(net455),
    .S(net138),
    .X(\proj_14.net424 ));
 sg13g2_mux2_1 \proj_14.mux138/_0_  (.A0(net26),
    .A1(net557),
    .S(net138),
    .X(\proj_14.net427 ));
 sg13g2_mux2_1 \proj_14.mux139/_0_  (.A0(net107),
    .A1(net461),
    .S(net137),
    .X(\proj_14.net430 ));
 sg13g2_mux2_1 \proj_14.mux14/_0_  (.A0(net27),
    .A1(net533),
    .S(net148),
    .X(\proj_14.net45 ));
 sg13g2_mux2_1 \proj_14.mux140/_0_  (.A0(net28),
    .A1(net495),
    .S(net137),
    .X(\proj_14.net433 ));
 sg13g2_mux2_1 \proj_14.mux141/_0_  (.A0(net108),
    .A1(net498),
    .S(net137),
    .X(\proj_14.net436 ));
 sg13g2_mux2_1 \proj_14.mux142/_0_  (.A0(net109),
    .A1(net564),
    .S(net137),
    .X(\proj_14.net439 ));
 sg13g2_mux2_1 \proj_14.mux143/_0_  (.A0(net110),
    .A1(net515),
    .S(net137),
    .X(\proj_14.net442 ));
 sg13g2_mux2_1 \proj_14.mux144/_0_  (.A0(net111),
    .A1(net538),
    .S(net137),
    .X(\proj_14.net445 ));
 sg13g2_mux2_1 \proj_14.mux145/_0_  (.A0(net112),
    .A1(net484),
    .S(net155),
    .X(\proj_14.net449 ));
 sg13g2_mux2_1 \proj_14.mux146/_0_  (.A0(net113),
    .A1(net499),
    .S(net144),
    .X(\proj_14.net452 ));
 sg13g2_mux2_1 \proj_14.mux147/_0_  (.A0(net114),
    .A1(net453),
    .S(net144),
    .X(\proj_14.net455 ));
 sg13g2_mux2_1 \proj_14.mux148/_0_  (.A0(net115),
    .A1(net543),
    .S(net143),
    .X(\proj_14.net458 ));
 sg13g2_mux2_1 \proj_14.mux149/_0_  (.A0(net116),
    .A1(net490),
    .S(net139),
    .X(\proj_14.net460 ));
 sg13g2_mux2_1 \proj_14.mux15/_0_  (.A0(net117),
    .A1(net457),
    .S(net148),
    .X(\proj_14.net48 ));
 sg13g2_mux2_1 \proj_14.mux150/_0_  (.A0(net118),
    .A1(net471),
    .S(net139),
    .X(\proj_14.net464 ));
 sg13g2_mux2_1 \proj_14.mux151/_0_  (.A0(net119),
    .A1(net541),
    .S(net139),
    .X(\proj_14.net467 ));
 sg13g2_mux2_1 \proj_14.mux152/_0_  (.A0(net120),
    .A1(net518),
    .S(net140),
    .X(\proj_14.net470 ));
 sg13g2_mux2_1 \proj_14.mux153/_0_  (.A0(net29),
    .A1(net544),
    .S(net147),
    .X(\proj_14.net473 ));
 sg13g2_mux2_1 \proj_14.mux154/_0_  (.A0(net30),
    .A1(net443),
    .S(net147),
    .X(\proj_14.net476 ));
 sg13g2_mux2_1 \proj_14.mux155/_0_  (.A0(net121),
    .A1(net582),
    .S(net147),
    .X(\proj_14.net479 ));
 sg13g2_mux2_1 \proj_14.mux156/_0_  (.A0(net31),
    .A1(net458),
    .S(net147),
    .X(\proj_14.net482 ));
 sg13g2_mux2_1 \proj_14.mux157/_0_  (.A0(net122),
    .A1(net535),
    .S(net146),
    .X(\proj_14.net485 ));
 sg13g2_mux2_1 \proj_14.mux158/_0_  (.A0(net32),
    .A1(net466),
    .S(net146),
    .X(\proj_14.net488 ));
 sg13g2_mux2_1 \proj_14.mux159/_0_  (.A0(net33),
    .A1(net603),
    .S(net148),
    .X(\proj_14.net491 ));
 sg13g2_mux2_1 \proj_14.mux16/_0_  (.A0(net123),
    .A1(net512),
    .S(net146),
    .X(\proj_14.net51 ));
 sg13g2_mux2_1 \proj_14.mux160/_0_  (.A0(net34),
    .A1(net531),
    .S(net151),
    .X(\proj_14.net494 ));
 sg13g2_mux2_1 \proj_14.mux161/_0_  (.A0(net35),
    .A1(net468),
    .S(net151),
    .X(\proj_14.net497 ));
 sg13g2_mux2_1 \proj_14.mux162/_0_  (.A0(net124),
    .A1(net497),
    .S(net149),
    .X(\proj_14.net500 ));
 sg13g2_mux2_1 \proj_14.mux163/_0_  (.A0(net125),
    .A1(net507),
    .S(net151),
    .X(\proj_14.net503 ));
 sg13g2_mux2_1 \proj_14.mux164/_0_  (.A0(net126),
    .A1(net459),
    .S(net151),
    .X(\proj_14.net506 ));
 sg13g2_mux2_1 \proj_14.mux165/_0_  (.A0(net127),
    .A1(\proj_14.net4 ),
    .S(net151),
    .X(\proj_14.net509 ));
 sg13g2_mux2_1 \proj_14.mux166/_0_  (.A0(net128),
    .A1(net536),
    .S(net137),
    .X(\proj_14.net512 ));
 sg13g2_mux2_1 \proj_14.mux167/_0_  (.A0(net129),
    .A1(net480),
    .S(net137),
    .X(\proj_14.net515 ));
 sg13g2_mux2_1 \proj_14.mux168/_0_  (.A0(net130),
    .A1(net465),
    .S(net139),
    .X(\proj_14.net518 ));
 sg13g2_mux2_1 \proj_14.mux169/_0_  (.A0(net131),
    .A1(net523),
    .S(net139),
    .X(\proj_14.net521 ));
 sg13g2_mux2_1 \proj_14.mux17/_0_  (.A0(net132),
    .A1(net553),
    .S(net146),
    .X(\proj_14.net54 ));
 sg13g2_mux2_1 \proj_14.mux18/_0_  (.A0(net133),
    .A1(net551),
    .S(net146),
    .X(\proj_14.net57 ));
 sg13g2_mux2_1 \proj_14.mux19/_0_  (.A0(net134),
    .A1(net552),
    .S(net140),
    .X(\proj_14.net63 ));
 sg13g2_mux2_1 \proj_14.mux2/_0_  (.A0(net181),
    .A1(net604),
    .S(net136),
    .X(\proj_14.net4 ));
 sg13g2_mux2_1 \proj_14.mux20/_0_  (.A0(net182),
    .A1(net568),
    .S(net140),
    .X(\proj_14.net67 ));
 sg13g2_mux2_1 \proj_14.mux21/_0_  (.A0(net183),
    .A1(net492),
    .S(net143),
    .X(\proj_14.net70 ));
 sg13g2_mux2_1 \proj_14.mux22/_0_  (.A0(net184),
    .A1(net556),
    .S(net143),
    .X(\proj_14.net73 ));
 sg13g2_mux2_1 \proj_14.mux23/_0_  (.A0(net36),
    .A1(net519),
    .S(net143),
    .X(\proj_14.net76 ));
 sg13g2_mux2_1 \proj_14.mux24/_0_  (.A0(net37),
    .A1(net513),
    .S(net150),
    .X(\proj_14.net79 ));
 sg13g2_mux2_1 \proj_14.mux25/_0_  (.A0(net38),
    .A1(net572),
    .S(net150),
    .X(\proj_14.net82 ));
 sg13g2_mux2_1 \proj_14.mux26/_0_  (.A0(net39),
    .A1(net579),
    .S(net150),
    .X(\proj_14.net85 ));
 sg13g2_mux2_1 \proj_14.mux27/_0_  (.A0(net185),
    .A1(net555),
    .S(net152),
    .X(\proj_14.net88 ));
 sg13g2_mux2_1 \proj_14.mux28/_0_  (.A0(net40),
    .A1(net470),
    .S(net152),
    .X(\proj_14.net91 ));
 sg13g2_mux2_1 \proj_14.mux29/_0_  (.A0(net41),
    .A1(net542),
    .S(net150),
    .X(\proj_14.net94 ));
 sg13g2_mux2_1 \proj_14.mux3/_0_  (.A0(net186),
    .A1(net451),
    .S(net150),
    .X(\proj_14.net12 ));
 sg13g2_mux2_1 \proj_14.mux30/_0_  (.A0(net187),
    .A1(net601),
    .S(net163),
    .X(\proj_14.net97 ));
 sg13g2_mux2_1 \proj_14.mux31/_0_  (.A0(net42),
    .A1(net437),
    .S(net163),
    .X(\proj_14.net100 ));
 sg13g2_mux2_1 \proj_14.mux32/_0_  (.A0(net188),
    .A1(net583),
    .S(net163),
    .X(\proj_14.net103 ));
 sg13g2_mux2_1 \proj_14.mux33/_0_  (.A0(net189),
    .A1(net591),
    .S(net163),
    .X(\proj_14.net106 ));
 sg13g2_mux2_1 \proj_14.mux34/_0_  (.A0(net190),
    .A1(net539),
    .S(net165),
    .X(\proj_14.net109 ));
 sg13g2_mux2_1 \proj_14.mux35/_0_  (.A0(net191),
    .A1(net595),
    .S(net165),
    .X(\proj_14.net112 ));
 sg13g2_mux2_1 \proj_14.mux36/_0_  (.A0(net192),
    .A1(net573),
    .S(net146),
    .X(\proj_14.net116 ));
 sg13g2_mux2_1 \proj_14.mux37/_0_  (.A0(net193),
    .A1(net472),
    .S(net146),
    .X(\proj_14.net119 ));
 sg13g2_mux2_1 \proj_14.mux38/_0_  (.A0(net194),
    .A1(net540),
    .S(net139),
    .X(\proj_14.net122 ));
 sg13g2_mux2_1 \proj_14.mux39/_0_  (.A0(net195),
    .A1(net596),
    .S(net139),
    .X(\proj_14.net125 ));
 sg13g2_mux2_1 \proj_14.mux4/_0_  (.A0(net196),
    .A1(net529),
    .S(net150),
    .X(\proj_14.net15 ));
 sg13g2_mux2_1 \proj_14.mux40/_0_  (.A0(net197),
    .A1(net511),
    .S(net151),
    .X(\proj_14.net127 ));
 sg13g2_mux2_1 \proj_14.mux41/_0_  (.A0(net198),
    .A1(net438),
    .S(net151),
    .X(\proj_14.net131 ));
 sg13g2_mux2_1 \proj_14.mux42/_0_  (.A0(net199),
    .A1(net474),
    .S(net151),
    .X(\proj_14.net134 ));
 sg13g2_mux2_1 \proj_14.mux43/_0_  (.A0(net200),
    .A1(net590),
    .S(net152),
    .X(\proj_14.net137 ));
 sg13g2_mux2_1 \proj_14.mux44/_0_  (.A0(net201),
    .A1(net491),
    .S(net167),
    .X(\proj_14.net139 ));
 sg13g2_mux2_1 \proj_14.mux45/_0_  (.A0(net202),
    .A1(net516),
    .S(net167),
    .X(\proj_14.net143 ));
 sg13g2_mux2_1 \proj_14.mux46/_0_  (.A0(net203),
    .A1(net597),
    .S(net167),
    .X(\proj_14.net146 ));
 sg13g2_mux2_1 \proj_14.mux47/_0_  (.A0(net204),
    .A1(net464),
    .S(net167),
    .X(\proj_14.net149 ));
 sg13g2_mux2_1 \proj_14.mux48/_0_  (.A0(net43),
    .A1(net587),
    .S(net167),
    .X(\proj_14.net152 ));
 sg13g2_mux2_1 \proj_14.mux49/_0_  (.A0(net205),
    .A1(net475),
    .S(net166),
    .X(\proj_14.net155 ));
 sg13g2_mux2_1 \proj_14.mux5/_0_  (.A0(net206),
    .A1(net446),
    .S(net146),
    .X(\proj_14.net18 ));
 sg13g2_mux2_1 \proj_14.mux50/_0_  (.A0(net44),
    .A1(net577),
    .S(net166),
    .X(\proj_14.net158 ));
 sg13g2_mux2_1 \proj_14.mux51/_0_  (.A0(net45),
    .A1(net448),
    .S(net165),
    .X(\proj_14.net161 ));
 sg13g2_mux2_1 \proj_14.mux52/_0_  (.A0(net46),
    .A1(net501),
    .S(net166),
    .X(\proj_14.net164 ));
 sg13g2_mux2_1 \proj_14.mux53/_0_  (.A0(net47),
    .A1(net487),
    .S(net166),
    .X(\proj_14.net167 ));
 sg13g2_mux2_1 \proj_14.mux54/_0_  (.A0(net48),
    .A1(net567),
    .S(net160),
    .X(\proj_14.net170 ));
 sg13g2_mux2_1 \proj_14.mux55/_0_  (.A0(net207),
    .A1(net578),
    .S(net160),
    .X(\proj_14.net173 ));
 sg13g2_mux2_1 \proj_14.mux56/_0_  (.A0(net49),
    .A1(net441),
    .S(net160),
    .X(\proj_14.net176 ));
 sg13g2_mux2_1 \proj_14.mux57/_0_  (.A0(net208),
    .A1(net483),
    .S(net160),
    .X(\proj_14.net179 ));
 sg13g2_mux2_1 \proj_14.mux58/_0_  (.A0(net209),
    .A1(net545),
    .S(net158),
    .X(\proj_14.net182 ));
 sg13g2_mux2_1 \proj_14.mux59/_0_  (.A0(net210),
    .A1(net481),
    .S(net158),
    .X(\proj_14.net185 ));
 sg13g2_mux2_1 \proj_14.mux6/_0_  (.A0(net50),
    .A1(net488),
    .S(net149),
    .X(\proj_14.net21 ));
 sg13g2_mux2_1 \proj_14.mux60/_0_  (.A0(net211),
    .A1(net528),
    .S(net158),
    .X(\proj_14.net188 ));
 sg13g2_mux2_1 \proj_14.mux61/_0_  (.A0(net212),
    .A1(net503),
    .S(net165),
    .X(\proj_14.net192 ));
 sg13g2_mux2_1 \proj_14.mux62/_0_  (.A0(net213),
    .A1(net477),
    .S(net165),
    .X(\proj_14.net195 ));
 sg13g2_mux2_1 \proj_14.mux63/_0_  (.A0(net214),
    .A1(net588),
    .S(net168),
    .X(\proj_14.net198 ));
 sg13g2_mux2_1 \proj_14.mux64/_0_  (.A0(net215),
    .A1(net592),
    .S(net167),
    .X(\proj_14.net201 ));
 sg13g2_mux2_1 \proj_14.mux65/_0_  (.A0(net216),
    .A1(net546),
    .S(net154),
    .X(\proj_14.net203 ));
 sg13g2_mux2_1 \proj_14.mux66/_0_  (.A0(net217),
    .A1(net485),
    .S(net155),
    .X(\proj_14.net207 ));
 sg13g2_mux2_1 \proj_14.mux67/_0_  (.A0(net218),
    .A1(net530),
    .S(net144),
    .X(\proj_14.net210 ));
 sg13g2_mux2_1 \proj_14.mux68/_0_  (.A0(net219),
    .A1(net502),
    .S(net144),
    .X(\proj_14.net213 ));
 sg13g2_mux2_1 \proj_14.mux69/_0_  (.A0(net51),
    .A1(net532),
    .S(net145),
    .X(\proj_14.net216 ));
 sg13g2_mux2_1 \proj_14.mux7/_0_  (.A0(net220),
    .A1(net534),
    .S(net149),
    .X(\proj_14.net24 ));
 sg13g2_mux2_1 \proj_14.mux70/_0_  (.A0(net221),
    .A1(net565),
    .S(net142),
    .X(\proj_14.net219 ));
 sg13g2_mux2_1 \proj_14.mux71/_0_  (.A0(net222),
    .A1(net456),
    .S(net142),
    .X(\proj_14.net222 ));
 sg13g2_mux2_1 \proj_14.mux72/_0_  (.A0(net223),
    .A1(net450),
    .S(net142),
    .X(\proj_14.net225 ));
 sg13g2_mux2_1 \proj_14.mux73/_0_  (.A0(net224),
    .A1(net494),
    .S(net138),
    .X(\proj_14.net228 ));
 sg13g2_mux2_1 \proj_14.mux74/_0_  (.A0(net52),
    .A1(net570),
    .S(net138),
    .X(\proj_14.net231 ));
 sg13g2_mux2_1 \proj_14.mux75/_0_  (.A0(net53),
    .A1(net493),
    .S(net138),
    .X(\proj_14.net234 ));
 sg13g2_mux2_1 \proj_14.mux76/_0_  (.A0(net225),
    .A1(net586),
    .S(net142),
    .X(\proj_14.net237 ));
 sg13g2_mux2_1 \proj_14.mux77/_0_  (.A0(net54),
    .A1(net574),
    .S(net142),
    .X(\proj_14.net240 ));
 sg13g2_mux2_1 \proj_14.mux78/_0_  (.A0(net226),
    .A1(net463),
    .S(net145),
    .X(\proj_14.net243 ));
 sg13g2_mux2_1 \proj_14.mux79/_0_  (.A0(net227),
    .A1(net585),
    .S(net145),
    .X(\proj_14.net246 ));
 sg13g2_mux2_1 \proj_14.mux8/_0_  (.A0(net228),
    .A1(net476),
    .S(net148),
    .X(\proj_14.net27 ));
 sg13g2_mux2_1 \proj_14.mux80/_0_  (.A0(net229),
    .A1(net571),
    .S(net142),
    .X(\proj_14.net249 ));
 sg13g2_mux2_1 \proj_14.mux81/_0_  (.A0(net230),
    .A1(net460),
    .S(net142),
    .X(\proj_14.net252 ));
 sg13g2_mux2_1 \proj_14.mux82/_0_  (.A0(net231),
    .A1(net517),
    .S(net154),
    .X(\proj_14.net256 ));
 sg13g2_mux2_1 \proj_14.mux83/_0_  (.A0(net232),
    .A1(net566),
    .S(net157),
    .X(\proj_14.net259 ));
 sg13g2_mux2_1 \proj_14.mux84/_0_  (.A0(net233),
    .A1(net473),
    .S(net154),
    .X(\proj_14.net262 ));
 sg13g2_mux2_1 \proj_14.mux85/_0_  (.A0(net234),
    .A1(net444),
    .S(net154),
    .X(\proj_14.net265 ));
 sg13g2_mux2_1 \proj_14.mux86/_0_  (.A0(net235),
    .A1(net447),
    .S(net154),
    .X(\proj_14.net267 ));
 sg13g2_mux2_1 \proj_14.mux87/_0_  (.A0(net236),
    .A1(net598),
    .S(net158),
    .X(\proj_14.net271 ));
 sg13g2_mux2_1 \proj_14.mux88/_0_  (.A0(net237),
    .A1(net569),
    .S(net158),
    .X(\proj_14.net274 ));
 sg13g2_mux2_1 \proj_14.mux89/_0_  (.A0(net238),
    .A1(net500),
    .S(net158),
    .X(\proj_14.net277 ));
 sg13g2_mux2_1 \proj_14.mux9/_0_  (.A0(net55),
    .A1(net581),
    .S(net148),
    .X(\proj_14.net30 ));
 sg13g2_mux2_1 \proj_14.mux90/_0_  (.A0(net56),
    .A1(net510),
    .S(net158),
    .X(\proj_14.net280 ));
 sg13g2_mux2_1 \proj_14.mux91/_0_  (.A0(net239),
    .A1(net584),
    .S(net158),
    .X(\proj_14.net283 ));
 sg13g2_mux2_1 \proj_14.mux92/_0_  (.A0(net240),
    .A1(net527),
    .S(net159),
    .X(\proj_14.net286 ));
 sg13g2_mux2_1 \proj_14.mux93/_0_  (.A0(net57),
    .A1(net580),
    .S(net159),
    .X(\proj_14.net289 ));
 sg13g2_mux2_1 \proj_14.mux94/_0_  (.A0(net241),
    .A1(net445),
    .S(net159),
    .X(\proj_14.net292 ));
 sg13g2_mux2_1 \proj_14.mux95/_0_  (.A0(net58),
    .A1(net576),
    .S(net159),
    .X(\proj_14.net295 ));
 sg13g2_mux2_1 \proj_14.mux96/_0_  (.A0(net59),
    .A1(net449),
    .S(net159),
    .X(\proj_14.net298 ));
 sg13g2_mux2_1 \proj_14.mux97/_0_  (.A0(net242),
    .A1(net558),
    .S(net159),
    .X(\proj_14.net301 ));
 sg13g2_mux2_1 \proj_14.mux98/_0_  (.A0(net60),
    .A1(net575),
    .S(net159),
    .X(\proj_14.net304 ));
 sg13g2_mux2_1 \proj_14.mux99/_0_  (.A0(net243),
    .A1(net504),
    .S(net159),
    .X(\proj_14.net307 ));
 sg13g2_and2_1 \proj_15.and1/_0_  (.A(net4),
    .B(net178),
    .X(\proj_15.net10 ));
 sg13g2_and2_1 \proj_15.and2/_0_  (.A(net174),
    .B(net176),
    .X(\proj_15.net14 ));
 sg13g2_nand2_1 \proj_15.nand1/_0_  (.Y(\proj_15.net11 ),
    .A(net172),
    .B(net173));
 sg13g2_inv_1 \proj_15.not1/_0_  (.Y(\proj_15.net9 ),
    .A(net179));
 sg13g2_or2_1 \proj_15.or1/_0_  (.X(\proj_15.net13 ),
    .B(net136),
    .A(net180));
 sg13g2_or2_1 \proj_15.or2/_0_  (.X(\proj_15.net15 ),
    .B(net173),
    .A(net172));
 sg13g2_xor2_1 \proj_15.xor1/_0_  (.B(net171),
    .A(net164),
    .X(\proj_15.net12 ));
 sg13g2_xor2_1 \proj_15.xor2/_0_  (.B(net7),
    .A(net167),
    .X(\proj_15.net16 ));
 sg13g2_inv_1 \proj__0.not1/_0_  (.Y(\proj__0.net4 ),
    .A(\proj__0.net11 ));
 sg13g2_inv_1 \proj__0.not2/_0_  (.Y(\proj__0.net3 ),
    .A(\proj__0.net10 ));
 sg13g2_or2_1 \proj__0.or1/_0_  (.X(\proj__0.net10 ),
    .B(net2),
    .A(\proj__0.net4 ));
 sg13g2_or2_1 \proj__0.or2/_0_  (.X(\proj__0.net11 ),
    .B(\proj__0.net3 ),
    .A(net3));
 sg13g2_nand2_1 \proj__1.nand1/_0_  (.Y(\proj__1.net9 ),
    .A(net176),
    .B(net180));
 sg13g2_inv_1 \proj__1.not3/_0_  (.Y(\proj__1.net10 ),
    .A(net174));
 sg13g2_inv_1 \proj__1.not4/_0_  (.Y(\proj__1.net11 ),
    .A(net173));
 sg13g2_and2_1 \proj__2.and1/_0_  (.A(net177),
    .B(net180),
    .X(\proj__2.net7 ));
 sg13g2_and2_1 \proj__2.and2/_0_  (.A(\proj__2.net3 ),
    .B(\proj__2.net5 ),
    .X(\proj__2.net6 ));
 sg13g2_inv_1 \proj__2.not1/_0_  (.Y(\proj__2.net3 ),
    .A(\proj__2.net14 ));
 sg13g2_inv_1 \proj__2.not2/_0_  (.Y(\proj__2.net5 ),
    .A(\proj__2.net7 ));
 sg13g2_xor2_1 \proj__2.xor1/_0_  (.B(net180),
    .A(net176),
    .X(\proj__2.net14 ));
 sg13g2_and2_1 \proj__3.and1/_0_  (.A(net178),
    .B(\proj__3.net10 ),
    .X(\proj__3.net11 ));
 sg13g2_and2_1 \proj__3.and2/_0_  (.A(net177),
    .B(net7),
    .X(\proj__3.net4 ));
 sg13g2_and2_1 \proj__3.and3/_0_  (.A(\proj__3.net12 ),
    .B(net171),
    .X(\proj__3.net13 ));
 sg13g2_and2_1 \proj__3.and4/_0_  (.A(\proj__3.net13 ),
    .B(\proj__3.net11 ),
    .X(\proj__3.net3 ));
 sg13g2_inv_1 \proj__3.not1/_0_  (.Y(\proj__3.net10 ),
    .A(net171));
 sg13g2_inv_1 \proj__3.not2/_0_  (.Y(\proj__3.net12 ),
    .A(net178));
 sg13g2_inv_1 \proj__4.not1/_0_  (.Y(\proj__4.net9 ),
    .A(net179));
 sg13g2_inv_1 \proj__4.not2/_0_  (.Y(\proj__4.net10 ),
    .A(net177));
 sg13g2_inv_1 \proj__4.not3/_0_  (.Y(\proj__4.net11 ),
    .A(net174));
 sg13g2_inv_1 \proj__4.not4/_0_  (.Y(\proj__4.net12 ),
    .A(net173));
 sg13g2_inv_1 \proj__5.not1/_0_  (.Y(\proj__5.net9 ),
    .A(net164));
 sg13g2_or2_1 \proj__5.or1/_0_  (.X(\proj__5.net8 ),
    .B(net5),
    .A(net172));
 sg13g2_and2_1 \proj__6.and2/_0_  (.A(net176),
    .B(net179),
    .X(\proj__6.net4 ));
 sg13g2_xor2_1 \proj__6.xor1/_0_  (.B(net179),
    .A(net178),
    .X(\proj__6.net3 ));
 sg13g2_xor2_1 \proj__7.xor1/_0_  (.B(net179),
    .A(net178),
    .X(\proj__7.net3 ));
 sg13g2_and2_1 \proj__8.and1/_0_  (.A(net175),
    .B(net176),
    .X(\proj__8.net18 ));
 sg13g2_and2_1 \proj__8.and2/_0_  (.A(net180),
    .B(\proj__8.net19 ),
    .X(\proj__8.net20 ));
 sg13g2_inv_1 \proj__8.not1/_0_  (.Y(\proj__8.net8 ),
    .A(\proj__8.net18 ));
 sg13g2_inv_1 \proj__8.not2/_0_  (.Y(\proj__8.net19 ),
    .A(\proj__8.net18 ));
 sg13g2_or2_1 \proj__8.or1/_0_  (.X(\proj__8.net12 ),
    .B(\proj__8.net18 ),
    .A(net172));
 sg13g2_or2_1 \proj__8.or2/_0_  (.X(\proj__8.net11 ),
    .B(\proj__8.net20 ),
    .A(\proj__8.net12 ));
 sg13g2_or2_1 \proj__8.or3/_0_  (.X(\proj__8.net7 ),
    .B(\proj__8.net20 ),
    .A(net136));
 sg13g2_or2_1 \proj__8.or4/_0_  (.X(\proj__8.net10 ),
    .B(net164),
    .A(\proj__8.net20 ));
 sg13g2_or2_1 \proj__8.or5/_0_  (.X(\proj__8.net9 ),
    .B(\proj__8.net10 ),
    .A(\proj__8.net20 ));
 sg13g2_buf_2 fanout135 (.A(net9),
    .X(net135));
 sg13g2_buf_2 fanout136 (.A(net8),
    .X(net136));
 sg13g2_buf_4 fanout137 (.X(net137),
    .A(net141));
 sg13g2_buf_4 fanout138 (.X(net138),
    .A(net141));
 sg13g2_buf_4 fanout139 (.X(net139),
    .A(net141));
 sg13g2_buf_2 fanout140 (.A(net141),
    .X(net140));
 sg13g2_buf_2 fanout141 (.A(net170),
    .X(net141));
 sg13g2_buf_4 fanout142 (.X(net142),
    .A(net145));
 sg13g2_buf_4 fanout143 (.X(net143),
    .A(net145));
 sg13g2_buf_2 fanout144 (.A(net145),
    .X(net144));
 sg13g2_buf_2 fanout145 (.A(net170),
    .X(net145));
 sg13g2_buf_4 fanout146 (.X(net146),
    .A(net153));
 sg13g2_buf_2 fanout147 (.A(net153),
    .X(net147));
 sg13g2_buf_4 fanout148 (.X(net148),
    .A(net149));
 sg13g2_buf_2 fanout149 (.A(net153),
    .X(net149));
 sg13g2_buf_4 fanout150 (.X(net150),
    .A(net152));
 sg13g2_buf_4 fanout151 (.X(net151),
    .A(net152));
 sg13g2_buf_2 fanout152 (.A(net153),
    .X(net152));
 sg13g2_buf_2 fanout153 (.A(net170),
    .X(net153));
 sg13g2_buf_4 fanout154 (.X(net154),
    .A(net157));
 sg13g2_buf_4 fanout155 (.X(net155),
    .A(net157));
 sg13g2_buf_2 fanout156 (.A(net157),
    .X(net156));
 sg13g2_buf_2 fanout157 (.A(net169),
    .X(net157));
 sg13g2_buf_4 fanout158 (.X(net158),
    .A(net162));
 sg13g2_buf_4 fanout159 (.X(net159),
    .A(net162));
 sg13g2_buf_4 fanout160 (.X(net160),
    .A(net162));
 sg13g2_buf_2 fanout161 (.A(net162),
    .X(net161));
 sg13g2_buf_2 fanout162 (.A(net169),
    .X(net162));
 sg13g2_buf_4 fanout163 (.X(net163),
    .A(net169));
 sg13g2_buf_2 fanout164 (.A(net169),
    .X(net164));
 sg13g2_buf_4 fanout165 (.X(net165),
    .A(net168));
 sg13g2_buf_2 fanout166 (.A(net168),
    .X(net166));
 sg13g2_buf_4 fanout167 (.X(net167),
    .A(net168));
 sg13g2_buf_2 fanout168 (.A(net169),
    .X(net168));
 sg13g2_buf_2 fanout169 (.A(net170),
    .X(net169));
 sg13g2_buf_2 fanout170 (.A(ui_in[6]),
    .X(net170));
 sg13g2_buf_2 fanout171 (.A(net7),
    .X(net171));
 sg13g2_buf_2 fanout172 (.A(net6),
    .X(net172));
 sg13g2_buf_2 fanout173 (.A(net5),
    .X(net173));
 sg13g2_buf_2 fanout174 (.A(net175),
    .X(net174));
 sg13g2_buf_1 fanout175 (.A(net4),
    .X(net175));
 sg13g2_buf_2 fanout176 (.A(net178),
    .X(net176));
 sg13g2_buf_1 fanout177 (.A(net178),
    .X(net177));
 sg13g2_buf_2 fanout178 (.A(net3),
    .X(net178));
 sg13g2_buf_2 fanout179 (.A(net2),
    .X(net179));
 sg13g2_buf_2 fanout180 (.A(net2),
    .X(net180));
 sg13g2_buf_1 input1 (.A(rst_n),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[0]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[1]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[2]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[3]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[4]),
    .X(net6));
 sg13g2_buf_2 input7 (.A(ui_in[5]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(ui_in[7]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(uio_in[0]),
    .X(net9));
 sg13g2_buf_2 input10 (.A(uio_in[1]),
    .X(net10));
 sg13g2_buf_1 input11 (.A(uio_in[2]),
    .X(net11));
 sg13g2_buf_1 input12 (.A(uio_in[3]),
    .X(net12));
 sg13g2_tielo \proj_14.mux10/_0__13  (.L_LO(net13));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_2 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .X(clknet_1_0__leaf_clk));
 sg13g2_buf_2 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .X(clknet_1_1__leaf_clk));
 sg13g2_buf_1 clkload0 (.A(clknet_1_0__leaf_clk));
 sg13g2_buf_2 clkbuf_0_clk_regs (.A(clk_regs),
    .X(clknet_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_0_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_0_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_1_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_1_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_2_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_2_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_3_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_3_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_4_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_4_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_5_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_5_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_6_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_6_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_7_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_7_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_8_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_8_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_9_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_9_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_10_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_10_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_11_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_11_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_12_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_12_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_13_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_13_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_14_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_14_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_15_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_15_0_clk_regs));
 sg13g2_buf_2 clkbuf_5_0__f_clk_regs (.A(clknet_4_0_0_clk_regs),
    .X(clknet_5_0__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_1__f_clk_regs (.A(clknet_4_0_0_clk_regs),
    .X(clknet_5_1__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_2__f_clk_regs (.A(clknet_4_1_0_clk_regs),
    .X(clknet_5_2__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_3__f_clk_regs (.A(clknet_4_1_0_clk_regs),
    .X(clknet_5_3__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_4__f_clk_regs (.A(clknet_4_2_0_clk_regs),
    .X(clknet_5_4__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_5__f_clk_regs (.A(clknet_4_2_0_clk_regs),
    .X(clknet_5_5__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_6__f_clk_regs (.A(clknet_4_3_0_clk_regs),
    .X(clknet_5_6__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_7__f_clk_regs (.A(clknet_4_3_0_clk_regs),
    .X(clknet_5_7__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_8__f_clk_regs (.A(clknet_4_4_0_clk_regs),
    .X(clknet_5_8__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_9__f_clk_regs (.A(clknet_4_4_0_clk_regs),
    .X(clknet_5_9__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_10__f_clk_regs (.A(clknet_4_5_0_clk_regs),
    .X(clknet_5_10__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_11__f_clk_regs (.A(clknet_4_5_0_clk_regs),
    .X(clknet_5_11__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_12__f_clk_regs (.A(clknet_4_6_0_clk_regs),
    .X(clknet_5_12__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_13__f_clk_regs (.A(clknet_4_6_0_clk_regs),
    .X(clknet_5_13__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_14__f_clk_regs (.A(clknet_4_7_0_clk_regs),
    .X(clknet_5_14__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_15__f_clk_regs (.A(clknet_4_7_0_clk_regs),
    .X(clknet_5_15__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_16__f_clk_regs (.A(clknet_4_8_0_clk_regs),
    .X(clknet_5_16__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_17__f_clk_regs (.A(clknet_4_8_0_clk_regs),
    .X(clknet_5_17__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_18__f_clk_regs (.A(clknet_4_9_0_clk_regs),
    .X(clknet_5_18__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_19__f_clk_regs (.A(clknet_4_9_0_clk_regs),
    .X(clknet_5_19__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_20__f_clk_regs (.A(clknet_4_10_0_clk_regs),
    .X(clknet_5_20__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_21__f_clk_regs (.A(clknet_4_10_0_clk_regs),
    .X(clknet_5_21__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_22__f_clk_regs (.A(clknet_4_11_0_clk_regs),
    .X(clknet_5_22__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_23__f_clk_regs (.A(clknet_4_11_0_clk_regs),
    .X(clknet_5_23__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_24__f_clk_regs (.A(clknet_4_12_0_clk_regs),
    .X(clknet_5_24__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_25__f_clk_regs (.A(clknet_4_12_0_clk_regs),
    .X(clknet_5_25__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_26__f_clk_regs (.A(clknet_4_13_0_clk_regs),
    .X(clknet_5_26__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_27__f_clk_regs (.A(clknet_4_13_0_clk_regs),
    .X(clknet_5_27__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_28__f_clk_regs (.A(clknet_4_14_0_clk_regs),
    .X(clknet_5_28__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_29__f_clk_regs (.A(clknet_4_14_0_clk_regs),
    .X(clknet_5_29__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_30__f_clk_regs (.A(clknet_4_15_0_clk_regs),
    .X(clknet_5_30__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_31__f_clk_regs (.A(clknet_4_15_0_clk_regs),
    .X(clknet_5_31__leaf_clk_regs));
 sg13g2_inv_1 clkload1 (.A(clknet_5_3__leaf_clk_regs));
 sg13g2_inv_1 clkload2 (.A(clknet_5_7__leaf_clk_regs));
 sg13g2_inv_1 clkload3 (.A(clknet_5_11__leaf_clk_regs));
 sg13g2_inv_1 clkload4 (.A(clknet_5_13__leaf_clk_regs));
 sg13g2_inv_1 clkload5 (.A(clknet_5_15__leaf_clk_regs));
 sg13g2_inv_1 clkload6 (.A(clknet_5_19__leaf_clk_regs));
 sg13g2_inv_1 clkload7 (.A(clknet_5_23__leaf_clk_regs));
 sg13g2_inv_1 clkload8 (.A(clknet_5_27__leaf_clk_regs));
 sg13g2_inv_1 clkload9 (.A(clknet_5_29__leaf_clk_regs));
 sg13g2_inv_1 clkload10 (.A(clknet_5_31__leaf_clk_regs));
 sg13g2_dlygate4sd3_1 hold1 (.A(\proj_10.net40 ),
    .X(net427));
 sg13g2_dlygate4sd3_1 hold2 (.A(\proj_10.net45 ),
    .X(net428));
 sg13g2_dlygate4sd3_1 hold3 (.A(\proj_10.net46 ),
    .X(net429));
 sg13g2_dlygate4sd3_1 hold4 (.A(\proj_10.net36 ),
    .X(net430));
 sg13g2_dlygate4sd3_1 hold5 (.A(\proj_10.net42 ),
    .X(net431));
 sg13g2_dlygate4sd3_1 hold6 (.A(\proj_10.net34 ),
    .X(net432));
 sg13g2_dlygate4sd3_1 hold7 (.A(\proj_10.net35 ),
    .X(net433));
 sg13g2_dlygate4sd3_1 hold8 (.A(\proj_10.net29 ),
    .X(net434));
 sg13g2_dlygate4sd3_1 hold9 (.A(\proj_10.net38 ),
    .X(net435));
 sg13g2_dlygate4sd3_1 hold10 (.A(\proj_10.net31 ),
    .X(net436));
 sg13g2_dlygate4sd3_1 hold11 (.A(\proj_14.net102 ),
    .X(net437));
 sg13g2_dlygate4sd3_1 hold12 (.A(\proj_14.net133 ),
    .X(net438));
 sg13g2_dlygate4sd3_1 hold13 (.A(\proj_14.net333 ),
    .X(net439));
 sg13g2_dlygate4sd3_1 hold14 (.A(\proj_14.net371 ),
    .X(net440));
 sg13g2_dlygate4sd3_1 hold15 (.A(\proj_14.net178 ),
    .X(net441));
 sg13g2_dlygate4sd3_1 hold16 (.A(\proj_14.net365 ),
    .X(net442));
 sg13g2_dlygate4sd3_1 hold17 (.A(\proj_14.net478 ),
    .X(net443));
 sg13g2_dlygate4sd3_1 hold18 (.A(\proj_14.net204 ),
    .X(net444));
 sg13g2_dlygate4sd3_1 hold19 (.A(\proj_14.net294 ),
    .X(net445));
 sg13g2_dlygate4sd3_1 hold20 (.A(\proj_14.net20 ),
    .X(net446));
 sg13g2_dlygate4sd3_1 hold21 (.A(\proj_14.net270 ),
    .X(net447));
 sg13g2_dlygate4sd3_1 hold22 (.A(\proj_14.net163 ),
    .X(net448));
 sg13g2_dlygate4sd3_1 hold23 (.A(\proj_14.net300 ),
    .X(net449));
 sg13g2_dlygate4sd3_1 hold24 (.A(\proj_14.net227 ),
    .X(net450));
 sg13g2_dlygate4sd3_1 hold25 (.A(\proj_14.net14 ),
    .X(net451));
 sg13g2_dlygate4sd3_1 hold26 (.A(\proj_14.net414 ),
    .X(net452));
 sg13g2_dlygate4sd3_1 hold27 (.A(\proj_14.net457 ),
    .X(net453));
 sg13g2_dlygate4sd3_1 hold28 (.A(\proj_14.net38 ),
    .X(net454));
 sg13g2_dlygate4sd3_1 hold29 (.A(\proj_14.net426 ),
    .X(net455));
 sg13g2_dlygate4sd3_1 hold30 (.A(\proj_14.net224 ),
    .X(net456));
 sg13g2_dlygate4sd3_1 hold31 (.A(\proj_14.net50 ),
    .X(net457));
 sg13g2_dlygate4sd3_1 hold32 (.A(\proj_14.net484 ),
    .X(net458));
 sg13g2_dlygate4sd3_1 hold33 (.A(\proj_14.net508 ),
    .X(net459));
 sg13g2_dlygate4sd3_1 hold34 (.A(\proj_14.net254 ),
    .X(net460));
 sg13g2_dlygate4sd3_1 hold35 (.A(\proj_14.net432 ),
    .X(net461));
 sg13g2_dlygate4sd3_1 hold36 (.A(\proj_14.net405 ),
    .X(net462));
 sg13g2_dlygate4sd3_1 hold37 (.A(\proj_14.net245 ),
    .X(net463));
 sg13g2_dlygate4sd3_1 hold38 (.A(\proj_14.net151 ),
    .X(net464));
 sg13g2_dlygate4sd3_1 hold39 (.A(\proj_14.net520 ),
    .X(net465));
 sg13g2_dlygate4sd3_1 hold40 (.A(\proj_14.net490 ),
    .X(net466));
 sg13g2_dlygate4sd3_1 hold41 (.A(\proj_14.net387 ),
    .X(net467));
 sg13g2_dlygate4sd3_1 hold42 (.A(\proj_14.net499 ),
    .X(net468));
 sg13g2_dlygate4sd3_1 hold43 (.A(\proj_14.net338 ),
    .X(net469));
 sg13g2_dlygate4sd3_1 hold44 (.A(\proj_14.net93 ),
    .X(net470));
 sg13g2_dlygate4sd3_1 hold45 (.A(\proj_14.net466 ),
    .X(net471));
 sg13g2_dlygate4sd3_1 hold46 (.A(\proj_14.net121 ),
    .X(net472));
 sg13g2_dlygate4sd3_1 hold47 (.A(\proj_14.net264 ),
    .X(net473));
 sg13g2_dlygate4sd3_1 hold48 (.A(\proj_14.net136 ),
    .X(net474));
 sg13g2_dlygate4sd3_1 hold49 (.A(\proj_14.net157 ),
    .X(net475));
 sg13g2_dlygate4sd3_1 hold50 (.A(\proj_14.net29 ),
    .X(net476));
 sg13g2_dlygate4sd3_1 hold51 (.A(\proj_14.net197 ),
    .X(net477));
 sg13g2_dlygate4sd3_1 hold52 (.A(\proj_14.net411 ),
    .X(net478));
 sg13g2_dlygate4sd3_1 hold53 (.A(\proj_14.net374 ),
    .X(net479));
 sg13g2_dlygate4sd3_1 hold54 (.A(\proj_14.net517 ),
    .X(net480));
 sg13g2_dlygate4sd3_1 hold55 (.A(\proj_14.net187 ),
    .X(net481));
 sg13g2_dlygate4sd3_1 hold56 (.A(\proj_14.net383 ),
    .X(net482));
 sg13g2_dlygate4sd3_1 hold57 (.A(\proj_14.net181 ),
    .X(net483));
 sg13g2_dlygate4sd3_1 hold58 (.A(\proj_14.net451 ),
    .X(net484));
 sg13g2_dlygate4sd3_1 hold59 (.A(\proj_14.net209 ),
    .X(net485));
 sg13g2_dlygate4sd3_1 hold60 (.A(\proj_14.net315 ),
    .X(net486));
 sg13g2_dlygate4sd3_1 hold61 (.A(\proj_14.net169 ),
    .X(net487));
 sg13g2_dlygate4sd3_1 hold62 (.A(\proj_14.net23 ),
    .X(net488));
 sg13g2_dlygate4sd3_1 hold63 (.A(\proj_14.net341 ),
    .X(net489));
 sg13g2_dlygate4sd3_1 hold64 (.A(\proj_14.net463 ),
    .X(net490));
 sg13g2_dlygate4sd3_1 hold65 (.A(\proj_14.net142 ),
    .X(net491));
 sg13g2_dlygate4sd3_1 hold66 (.A(\proj_14.net72 ),
    .X(net492));
 sg13g2_dlygate4sd3_1 hold67 (.A(\proj_14.net236 ),
    .X(net493));
 sg13g2_dlygate4sd3_1 hold68 (.A(\proj_14.net230 ),
    .X(net494));
 sg13g2_dlygate4sd3_1 hold69 (.A(\proj_14.net435 ),
    .X(net495));
 sg13g2_dlygate4sd3_1 hold70 (.A(\proj_14.net41 ),
    .X(net496));
 sg13g2_dlygate4sd3_1 hold71 (.A(\proj_14.net502 ),
    .X(net497));
 sg13g2_dlygate4sd3_1 hold72 (.A(\proj_14.net438 ),
    .X(net498));
 sg13g2_dlygate4sd3_1 hold73 (.A(\proj_14.net454 ),
    .X(net499));
 sg13g2_dlygate4sd3_1 hold74 (.A(\proj_14.net279 ),
    .X(net500));
 sg13g2_dlygate4sd3_1 hold75 (.A(\proj_14.net166 ),
    .X(net501));
 sg13g2_dlygate4sd3_1 hold76 (.A(\proj_14.net215 ),
    .X(net502));
 sg13g2_dlygate4sd3_1 hold77 (.A(\proj_14.net194 ),
    .X(net503));
 sg13g2_dlygate4sd3_1 hold78 (.A(\proj_14.net309 ),
    .X(net504));
 sg13g2_dlygate4sd3_1 hold79 (.A(\proj_14.net268 ),
    .X(net505));
 sg13g2_dlygate4sd3_1 hold80 (.A(\proj_14.net408 ),
    .X(net506));
 sg13g2_dlygate4sd3_1 hold81 (.A(\proj_14.net505 ),
    .X(net507));
 sg13g2_dlygate4sd3_1 hold82 (.A(\proj_14.net420 ),
    .X(net508));
 sg13g2_dlygate4sd3_1 hold83 (.A(\proj_14.net344 ),
    .X(net509));
 sg13g2_dlygate4sd3_1 hold84 (.A(\proj_14.net282 ),
    .X(net510));
 sg13g2_dlygate4sd3_1 hold85 (.A(\proj_14.net130 ),
    .X(net511));
 sg13g2_dlygate4sd3_1 hold86 (.A(\proj_14.net53 ),
    .X(net512));
 sg13g2_dlygate4sd3_1 hold87 (.A(\proj_14.net81 ),
    .X(net513));
 sg13g2_dlygate4sd3_1 hold88 (.A(\proj_14.net399 ),
    .X(net514));
 sg13g2_dlygate4sd3_1 hold89 (.A(\proj_14.net444 ),
    .X(net515));
 sg13g2_dlygate4sd3_1 hold90 (.A(\proj_14.net145 ),
    .X(net516));
 sg13g2_dlygate4sd3_1 hold91 (.A(\proj_14.net258 ),
    .X(net517));
 sg13g2_dlygate4sd3_1 hold92 (.A(\proj_14.net472 ),
    .X(net518));
 sg13g2_dlygate4sd3_1 hold93 (.A(\proj_14.net78 ),
    .X(net519));
 sg13g2_dlygate4sd3_1 hold94 (.A(\proj_14.net393 ),
    .X(net520));
 sg13g2_dlygate4sd3_1 hold95 (.A(\proj_14.net359 ),
    .X(net521));
 sg13g2_dlygate4sd3_1 hold96 (.A(\proj_14.net318 ),
    .X(net522));
 sg13g2_dlygate4sd3_1 hold97 (.A(\proj_14.net461 ),
    .X(net523));
 sg13g2_dlygate4sd3_1 hold98 (.A(\proj_14.net423 ),
    .X(net524));
 sg13g2_dlygate4sd3_1 hold99 (.A(\proj_14.net350 ),
    .X(net525));
 sg13g2_dlygate4sd3_1 hold100 (.A(\proj_14.net347 ),
    .X(net526));
 sg13g2_dlygate4sd3_1 hold101 (.A(\proj_14.net288 ),
    .X(net527));
 sg13g2_dlygate4sd3_1 hold102 (.A(\proj_14.net190 ),
    .X(net528));
 sg13g2_dlygate4sd3_1 hold103 (.A(\proj_14.net17 ),
    .X(net529));
 sg13g2_dlygate4sd3_1 hold104 (.A(\proj_14.net212 ),
    .X(net530));
 sg13g2_dlygate4sd3_1 hold105 (.A(\proj_14.net496 ),
    .X(net531));
 sg13g2_dlygate4sd3_1 hold106 (.A(\proj_14.net218 ),
    .X(net532));
 sg13g2_dlygate4sd3_1 hold107 (.A(\proj_14.net47 ),
    .X(net533));
 sg13g2_dlygate4sd3_1 hold108 (.A(\proj_14.net26 ),
    .X(net534));
 sg13g2_dlygate4sd3_1 hold109 (.A(\proj_14.net487 ),
    .X(net535));
 sg13g2_dlygate4sd3_1 hold110 (.A(\proj_14.net514 ),
    .X(net536));
 sg13g2_dlygate4sd3_1 hold111 (.A(\proj_14.net380 ),
    .X(net537));
 sg13g2_dlygate4sd3_1 hold112 (.A(\proj_14.net447 ),
    .X(net538));
 sg13g2_dlygate4sd3_1 hold113 (.A(\proj_14.net111 ),
    .X(net539));
 sg13g2_dlygate4sd3_1 hold114 (.A(\proj_14.net124 ),
    .X(net540));
 sg13g2_dlygate4sd3_1 hold115 (.A(\proj_14.net469 ),
    .X(net541));
 sg13g2_dlygate4sd3_1 hold116 (.A(\proj_14.net96 ),
    .X(net542));
 sg13g2_dlygate4sd3_1 hold117 (.A(\proj_14.net397 ),
    .X(net543));
 sg13g2_dlygate4sd3_1 hold118 (.A(\proj_14.net475 ),
    .X(net544));
 sg13g2_dlygate4sd3_1 hold119 (.A(\proj_14.net184 ),
    .X(net545));
 sg13g2_dlygate4sd3_1 hold120 (.A(\proj_14.net206 ),
    .X(net546));
 sg13g2_dlygate4sd3_1 hold121 (.A(\proj_14.net335 ),
    .X(net547));
 sg13g2_dlygate4sd3_1 hold122 (.A(\proj_14.net312 ),
    .X(net548));
 sg13g2_dlygate4sd3_1 hold123 (.A(\proj_14.net328 ),
    .X(net549));
 sg13g2_dlygate4sd3_1 hold124 (.A(\proj_14.net44 ),
    .X(net550));
 sg13g2_dlygate4sd3_1 hold125 (.A(\proj_14.net59 ),
    .X(net551));
 sg13g2_dlygate4sd3_1 hold126 (.A(\proj_14.net66 ),
    .X(net552));
 sg13g2_dlygate4sd3_1 hold127 (.A(\proj_14.net56 ),
    .X(net553));
 sg13g2_dlygate4sd3_1 hold128 (.A(\proj_14.net35 ),
    .X(net554));
 sg13g2_dlygate4sd3_1 hold129 (.A(\proj_14.net90 ),
    .X(net555));
 sg13g2_dlygate4sd3_1 hold130 (.A(\proj_14.net75 ),
    .X(net556));
 sg13g2_dlygate4sd3_1 hold131 (.A(\proj_14.net429 ),
    .X(net557));
 sg13g2_dlygate4sd3_1 hold132 (.A(\proj_14.net303 ),
    .X(net558));
 sg13g2_dlygate4sd3_1 hold133 (.A(\proj_14.net353 ),
    .X(net559));
 sg13g2_dlygate4sd3_1 hold134 (.A(\proj_14.net356 ),
    .X(net560));
 sg13g2_dlygate4sd3_1 hold135 (.A(\proj_14.net377 ),
    .X(net561));
 sg13g2_dlygate4sd3_1 hold136 (.A(\proj_14.net322 ),
    .X(net562));
 sg13g2_dlygate4sd3_1 hold137 (.A(\proj_14.net402 ),
    .X(net563));
 sg13g2_dlygate4sd3_1 hold138 (.A(\proj_14.net441 ),
    .X(net564));
 sg13g2_dlygate4sd3_1 hold139 (.A(\proj_14.net221 ),
    .X(net565));
 sg13g2_dlygate4sd3_1 hold140 (.A(\proj_14.net261 ),
    .X(net566));
 sg13g2_dlygate4sd3_1 hold141 (.A(\proj_14.net172 ),
    .X(net567));
 sg13g2_dlygate4sd3_1 hold142 (.A(\proj_14.net69 ),
    .X(net568));
 sg13g2_dlygate4sd3_1 hold143 (.A(\proj_14.net276 ),
    .X(net569));
 sg13g2_dlygate4sd3_1 hold144 (.A(\proj_14.net233 ),
    .X(net570));
 sg13g2_dlygate4sd3_1 hold145 (.A(\proj_14.net251 ),
    .X(net571));
 sg13g2_dlygate4sd3_1 hold146 (.A(\proj_14.net84 ),
    .X(net572));
 sg13g2_dlygate4sd3_1 hold147 (.A(\proj_14.net118 ),
    .X(net573));
 sg13g2_dlygate4sd3_1 hold148 (.A(\proj_14.net242 ),
    .X(net574));
 sg13g2_dlygate4sd3_1 hold149 (.A(\proj_14.net306 ),
    .X(net575));
 sg13g2_dlygate4sd3_1 hold150 (.A(\proj_14.net297 ),
    .X(net576));
 sg13g2_dlygate4sd3_1 hold151 (.A(\proj_14.net160 ),
    .X(net577));
 sg13g2_dlygate4sd3_1 hold152 (.A(\proj_14.net175 ),
    .X(net578));
 sg13g2_dlygate4sd3_1 hold153 (.A(\proj_14.net87 ),
    .X(net579));
 sg13g2_dlygate4sd3_1 hold154 (.A(\proj_14.net291 ),
    .X(net580));
 sg13g2_dlygate4sd3_1 hold155 (.A(\proj_14.net32 ),
    .X(net581));
 sg13g2_dlygate4sd3_1 hold156 (.A(\proj_14.net481 ),
    .X(net582));
 sg13g2_dlygate4sd3_1 hold157 (.A(\proj_14.net105 ),
    .X(net583));
 sg13g2_dlygate4sd3_1 hold158 (.A(\proj_14.net285 ),
    .X(net584));
 sg13g2_dlygate4sd3_1 hold159 (.A(\proj_14.net248 ),
    .X(net585));
 sg13g2_dlygate4sd3_1 hold160 (.A(\proj_14.net239 ),
    .X(net586));
 sg13g2_dlygate4sd3_1 hold161 (.A(\proj_14.net154 ),
    .X(net587));
 sg13g2_dlygate4sd3_1 hold162 (.A(\proj_14.net200 ),
    .X(net588));
 sg13g2_dlygate4sd3_1 hold163 (.A(\proj_14.net11 ),
    .X(net589));
 sg13g2_dlygate4sd3_1 hold164 (.A(\proj_14.net9 ),
    .X(net590));
 sg13g2_dlygate4sd3_1 hold165 (.A(\proj_14.net108 ),
    .X(net591));
 sg13g2_dlygate4sd3_1 hold166 (.A(\proj_14.net140 ),
    .X(net592));
 sg13g2_dlygate4sd3_1 hold167 (.A(\proj_14.net390 ),
    .X(net593));
 sg13g2_dlygate4sd3_1 hold168 (.A(\proj_14.net368 ),
    .X(net594));
 sg13g2_dlygate4sd3_1 hold169 (.A(\proj_14.net114 ),
    .X(net595));
 sg13g2_dlygate4sd3_1 hold170 (.A(\proj_14.net64 ),
    .X(net596));
 sg13g2_dlygate4sd3_1 hold171 (.A(\proj_14.net148 ),
    .X(net597));
 sg13g2_dlygate4sd3_1 hold172 (.A(\proj_14.net273 ),
    .X(net598));
 sg13g2_dlygate4sd3_1 hold173 (.A(\proj_14.net417 ),
    .X(net599));
 sg13g2_dlygate4sd3_1 hold174 (.A(\proj_14.net325 ),
    .X(net600));
 sg13g2_dlygate4sd3_1 hold175 (.A(\proj_14.net99 ),
    .X(net601));
 sg13g2_dlygate4sd3_1 hold176 (.A(\proj_14.net362 ),
    .X(net602));
 sg13g2_dlygate4sd3_1 hold177 (.A(\proj_14.net493 ),
    .X(net603));
 sg13g2_dlygate4sd3_1 hold178 (.A(\proj_14.net128 ),
    .X(net604));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_fill_2 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_307 ();
 sg13g2_decap_8 FILLER_5_314 ();
 sg13g2_decap_8 FILLER_5_321 ();
 sg13g2_decap_8 FILLER_5_328 ();
 sg13g2_decap_8 FILLER_5_335 ();
 sg13g2_decap_8 FILLER_5_342 ();
 sg13g2_decap_8 FILLER_5_349 ();
 sg13g2_decap_8 FILLER_5_356 ();
 sg13g2_decap_8 FILLER_5_363 ();
 sg13g2_decap_8 FILLER_5_370 ();
 sg13g2_decap_8 FILLER_5_377 ();
 sg13g2_decap_8 FILLER_5_384 ();
 sg13g2_fill_2 FILLER_5_391 ();
 sg13g2_fill_1 FILLER_5_393 ();
 sg13g2_decap_8 FILLER_5_398 ();
 sg13g2_decap_4 FILLER_5_405 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_4 FILLER_6_133 ();
 sg13g2_fill_2 FILLER_6_137 ();
 sg13g2_fill_2 FILLER_6_143 ();
 sg13g2_fill_1 FILLER_6_145 ();
 sg13g2_decap_8 FILLER_6_156 ();
 sg13g2_fill_1 FILLER_6_163 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_fill_2 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_220 ();
 sg13g2_decap_8 FILLER_6_227 ();
 sg13g2_decap_8 FILLER_6_234 ();
 sg13g2_decap_8 FILLER_6_241 ();
 sg13g2_decap_8 FILLER_6_248 ();
 sg13g2_decap_8 FILLER_6_255 ();
 sg13g2_decap_8 FILLER_6_262 ();
 sg13g2_decap_8 FILLER_6_269 ();
 sg13g2_decap_8 FILLER_6_276 ();
 sg13g2_decap_8 FILLER_6_283 ();
 sg13g2_fill_2 FILLER_6_290 ();
 sg13g2_fill_1 FILLER_6_292 ();
 sg13g2_fill_1 FILLER_6_307 ();
 sg13g2_fill_2 FILLER_6_317 ();
 sg13g2_fill_1 FILLER_6_319 ();
 sg13g2_fill_2 FILLER_6_324 ();
 sg13g2_fill_1 FILLER_6_326 ();
 sg13g2_decap_8 FILLER_6_331 ();
 sg13g2_decap_4 FILLER_6_338 ();
 sg13g2_fill_2 FILLER_6_342 ();
 sg13g2_decap_8 FILLER_6_383 ();
 sg13g2_fill_2 FILLER_6_394 ();
 sg13g2_fill_1 FILLER_6_396 ();
 sg13g2_decap_4 FILLER_6_405 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_4 FILLER_7_63 ();
 sg13g2_fill_1 FILLER_7_67 ();
 sg13g2_decap_8 FILLER_7_94 ();
 sg13g2_decap_4 FILLER_7_101 ();
 sg13g2_fill_2 FILLER_7_109 ();
 sg13g2_decap_4 FILLER_7_121 ();
 sg13g2_fill_2 FILLER_7_125 ();
 sg13g2_fill_2 FILLER_7_179 ();
 sg13g2_fill_1 FILLER_7_181 ();
 sg13g2_fill_2 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_234 ();
 sg13g2_fill_1 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_256 ();
 sg13g2_decap_8 FILLER_7_263 ();
 sg13g2_fill_2 FILLER_7_270 ();
 sg13g2_decap_8 FILLER_7_282 ();
 sg13g2_fill_1 FILLER_7_289 ();
 sg13g2_fill_2 FILLER_7_360 ();
 sg13g2_fill_1 FILLER_7_372 ();
 sg13g2_decap_8 FILLER_8_26 ();
 sg13g2_decap_8 FILLER_8_33 ();
 sg13g2_decap_8 FILLER_8_40 ();
 sg13g2_decap_8 FILLER_8_47 ();
 sg13g2_decap_8 FILLER_8_54 ();
 sg13g2_decap_8 FILLER_8_65 ();
 sg13g2_decap_8 FILLER_8_130 ();
 sg13g2_fill_2 FILLER_8_137 ();
 sg13g2_fill_1 FILLER_8_139 ();
 sg13g2_fill_2 FILLER_8_149 ();
 sg13g2_fill_1 FILLER_8_155 ();
 sg13g2_fill_1 FILLER_8_185 ();
 sg13g2_fill_1 FILLER_8_213 ();
 sg13g2_fill_2 FILLER_8_227 ();
 sg13g2_fill_1 FILLER_8_229 ();
 sg13g2_fill_2 FILLER_8_260 ();
 sg13g2_fill_2 FILLER_8_301 ();
 sg13g2_fill_1 FILLER_8_303 ();
 sg13g2_decap_8 FILLER_8_346 ();
 sg13g2_fill_2 FILLER_8_353 ();
 sg13g2_fill_1 FILLER_8_355 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_4 FILLER_9_0 ();
 sg13g2_fill_2 FILLER_9_4 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_fill_2 FILLER_9_84 ();
 sg13g2_fill_1 FILLER_9_86 ();
 sg13g2_fill_2 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_97 ();
 sg13g2_fill_2 FILLER_9_104 ();
 sg13g2_fill_1 FILLER_9_106 ();
 sg13g2_fill_1 FILLER_9_167 ();
 sg13g2_fill_2 FILLER_9_198 ();
 sg13g2_fill_1 FILLER_9_200 ();
 sg13g2_decap_8 FILLER_9_227 ();
 sg13g2_fill_1 FILLER_9_234 ();
 sg13g2_fill_1 FILLER_9_258 ();
 sg13g2_fill_2 FILLER_9_287 ();
 sg13g2_fill_2 FILLER_9_306 ();
 sg13g2_fill_1 FILLER_9_308 ();
 sg13g2_fill_2 FILLER_9_371 ();
 sg13g2_fill_1 FILLER_9_373 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_4 FILLER_10_7 ();
 sg13g2_fill_2 FILLER_10_15 ();
 sg13g2_decap_4 FILLER_10_31 ();
 sg13g2_fill_2 FILLER_10_35 ();
 sg13g2_fill_2 FILLER_10_64 ();
 sg13g2_fill_2 FILLER_10_157 ();
 sg13g2_fill_2 FILLER_10_182 ();
 sg13g2_fill_2 FILLER_10_241 ();
 sg13g2_decap_8 FILLER_10_323 ();
 sg13g2_fill_1 FILLER_10_330 ();
 sg13g2_fill_2 FILLER_10_335 ();
 sg13g2_fill_2 FILLER_10_346 ();
 sg13g2_fill_1 FILLER_10_348 ();
 sg13g2_fill_2 FILLER_10_358 ();
 sg13g2_fill_1 FILLER_10_360 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_fill_1 FILLER_11_30 ();
 sg13g2_fill_1 FILLER_11_35 ();
 sg13g2_fill_1 FILLER_11_46 ();
 sg13g2_fill_2 FILLER_11_56 ();
 sg13g2_fill_1 FILLER_11_58 ();
 sg13g2_fill_1 FILLER_11_82 ();
 sg13g2_fill_2 FILLER_11_98 ();
 sg13g2_decap_4 FILLER_11_156 ();
 sg13g2_fill_2 FILLER_11_173 ();
 sg13g2_fill_1 FILLER_11_225 ();
 sg13g2_decap_4 FILLER_11_230 ();
 sg13g2_fill_2 FILLER_11_234 ();
 sg13g2_decap_8 FILLER_11_253 ();
 sg13g2_fill_1 FILLER_11_264 ();
 sg13g2_fill_1 FILLER_11_274 ();
 sg13g2_decap_8 FILLER_11_285 ();
 sg13g2_decap_4 FILLER_11_296 ();
 sg13g2_fill_1 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_320 ();
 sg13g2_fill_2 FILLER_11_327 ();
 sg13g2_fill_1 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_4 FILLER_12_7 ();
 sg13g2_fill_2 FILLER_12_24 ();
 sg13g2_decap_8 FILLER_12_127 ();
 sg13g2_decap_4 FILLER_12_134 ();
 sg13g2_fill_2 FILLER_12_138 ();
 sg13g2_fill_1 FILLER_12_193 ();
 sg13g2_decap_8 FILLER_12_220 ();
 sg13g2_fill_1 FILLER_12_333 ();
 sg13g2_fill_2 FILLER_12_338 ();
 sg13g2_decap_4 FILLER_12_344 ();
 sg13g2_fill_1 FILLER_12_348 ();
 sg13g2_fill_2 FILLER_12_381 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_4 FILLER_13_25 ();
 sg13g2_fill_1 FILLER_13_29 ();
 sg13g2_decap_4 FILLER_13_34 ();
 sg13g2_fill_1 FILLER_13_38 ();
 sg13g2_fill_1 FILLER_13_57 ();
 sg13g2_decap_8 FILLER_13_79 ();
 sg13g2_fill_2 FILLER_13_86 ();
 sg13g2_fill_1 FILLER_13_88 ();
 sg13g2_fill_2 FILLER_13_147 ();
 sg13g2_fill_1 FILLER_13_149 ();
 sg13g2_fill_1 FILLER_13_163 ();
 sg13g2_fill_2 FILLER_13_178 ();
 sg13g2_decap_8 FILLER_13_197 ();
 sg13g2_fill_1 FILLER_13_252 ();
 sg13g2_fill_2 FILLER_13_298 ();
 sg13g2_fill_1 FILLER_13_300 ();
 sg13g2_decap_4 FILLER_13_350 ();
 sg13g2_fill_1 FILLER_13_362 ();
 sg13g2_fill_2 FILLER_13_407 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_fill_2 FILLER_14_7 ();
 sg13g2_fill_1 FILLER_14_9 ();
 sg13g2_fill_2 FILLER_14_46 ();
 sg13g2_fill_1 FILLER_14_48 ();
 sg13g2_fill_1 FILLER_14_57 ();
 sg13g2_fill_1 FILLER_14_85 ();
 sg13g2_fill_2 FILLER_14_165 ();
 sg13g2_decap_8 FILLER_14_197 ();
 sg13g2_decap_8 FILLER_14_204 ();
 sg13g2_decap_8 FILLER_14_211 ();
 sg13g2_decap_4 FILLER_14_218 ();
 sg13g2_decap_8 FILLER_14_226 ();
 sg13g2_fill_1 FILLER_14_233 ();
 sg13g2_fill_1 FILLER_14_277 ();
 sg13g2_fill_1 FILLER_14_341 ();
 sg13g2_decap_4 FILLER_14_378 ();
 sg13g2_fill_1 FILLER_14_382 ();
 sg13g2_fill_1 FILLER_15_26 ();
 sg13g2_fill_1 FILLER_15_36 ();
 sg13g2_decap_4 FILLER_15_103 ();
 sg13g2_fill_1 FILLER_15_107 ();
 sg13g2_fill_1 FILLER_15_143 ();
 sg13g2_decap_4 FILLER_15_153 ();
 sg13g2_fill_2 FILLER_15_157 ();
 sg13g2_fill_2 FILLER_15_181 ();
 sg13g2_fill_1 FILLER_15_183 ();
 sg13g2_decap_4 FILLER_15_207 ();
 sg13g2_fill_1 FILLER_15_211 ();
 sg13g2_decap_8 FILLER_15_256 ();
 sg13g2_fill_2 FILLER_15_263 ();
 sg13g2_fill_1 FILLER_15_265 ();
 sg13g2_fill_2 FILLER_15_282 ();
 sg13g2_fill_1 FILLER_15_284 ();
 sg13g2_fill_1 FILLER_15_298 ();
 sg13g2_decap_8 FILLER_15_303 ();
 sg13g2_fill_1 FILLER_15_310 ();
 sg13g2_decap_8 FILLER_15_350 ();
 sg13g2_fill_2 FILLER_15_357 ();
 sg13g2_fill_1 FILLER_15_369 ();
 sg13g2_fill_1 FILLER_15_374 ();
 sg13g2_fill_1 FILLER_15_389 ();
 sg13g2_fill_2 FILLER_15_407 ();
 sg13g2_fill_2 FILLER_16_0 ();
 sg13g2_decap_4 FILLER_16_51 ();
 sg13g2_fill_2 FILLER_16_55 ();
 sg13g2_fill_1 FILLER_16_84 ();
 sg13g2_fill_2 FILLER_16_102 ();
 sg13g2_fill_1 FILLER_16_104 ();
 sg13g2_fill_2 FILLER_16_120 ();
 sg13g2_fill_1 FILLER_16_122 ();
 sg13g2_fill_2 FILLER_16_168 ();
 sg13g2_fill_1 FILLER_16_170 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_fill_1 FILLER_16_182 ();
 sg13g2_fill_2 FILLER_16_230 ();
 sg13g2_fill_1 FILLER_16_232 ();
 sg13g2_fill_2 FILLER_16_284 ();
 sg13g2_decap_8 FILLER_16_373 ();
 sg13g2_fill_2 FILLER_16_380 ();
 sg13g2_fill_1 FILLER_16_382 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_11 ();
 sg13g2_decap_4 FILLER_17_18 ();
 sg13g2_decap_8 FILLER_17_26 ();
 sg13g2_fill_2 FILLER_17_33 ();
 sg13g2_fill_1 FILLER_17_71 ();
 sg13g2_fill_2 FILLER_17_131 ();
 sg13g2_fill_1 FILLER_17_133 ();
 sg13g2_fill_2 FILLER_17_147 ();
 sg13g2_fill_1 FILLER_17_149 ();
 sg13g2_decap_8 FILLER_17_186 ();
 sg13g2_fill_1 FILLER_17_193 ();
 sg13g2_decap_4 FILLER_17_199 ();
 sg13g2_decap_4 FILLER_17_213 ();
 sg13g2_fill_1 FILLER_17_217 ();
 sg13g2_fill_2 FILLER_17_294 ();
 sg13g2_fill_1 FILLER_17_296 ();
 sg13g2_fill_2 FILLER_17_301 ();
 sg13g2_fill_1 FILLER_17_303 ();
 sg13g2_decap_4 FILLER_17_344 ();
 sg13g2_fill_2 FILLER_17_348 ();
 sg13g2_fill_1 FILLER_17_354 ();
 sg13g2_fill_2 FILLER_17_369 ();
 sg13g2_fill_1 FILLER_17_371 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_4 FILLER_18_21 ();
 sg13g2_fill_1 FILLER_18_25 ();
 sg13g2_decap_4 FILLER_18_31 ();
 sg13g2_fill_1 FILLER_18_39 ();
 sg13g2_fill_2 FILLER_18_53 ();
 sg13g2_fill_1 FILLER_18_55 ();
 sg13g2_decap_8 FILLER_18_60 ();
 sg13g2_fill_2 FILLER_18_67 ();
 sg13g2_fill_1 FILLER_18_79 ();
 sg13g2_fill_1 FILLER_18_94 ();
 sg13g2_fill_2 FILLER_18_107 ();
 sg13g2_fill_1 FILLER_18_109 ();
 sg13g2_decap_8 FILLER_18_169 ();
 sg13g2_decap_8 FILLER_18_232 ();
 sg13g2_fill_1 FILLER_18_243 ();
 sg13g2_fill_2 FILLER_18_272 ();
 sg13g2_fill_2 FILLER_18_296 ();
 sg13g2_fill_1 FILLER_18_308 ();
 sg13g2_fill_2 FILLER_18_341 ();
 sg13g2_fill_2 FILLER_18_407 ();
 sg13g2_decap_4 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_111 ();
 sg13g2_fill_2 FILLER_19_118 ();
 sg13g2_decap_8 FILLER_19_124 ();
 sg13g2_decap_8 FILLER_19_135 ();
 sg13g2_fill_2 FILLER_19_142 ();
 sg13g2_fill_1 FILLER_19_184 ();
 sg13g2_fill_1 FILLER_19_222 ();
 sg13g2_decap_8 FILLER_19_382 ();
 sg13g2_decap_8 FILLER_19_397 ();
 sg13g2_decap_4 FILLER_19_404 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_fill_1 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_45 ();
 sg13g2_fill_1 FILLER_20_133 ();
 sg13g2_fill_2 FILLER_20_138 ();
 sg13g2_fill_1 FILLER_20_140 ();
 sg13g2_decap_8 FILLER_20_151 ();
 sg13g2_decap_4 FILLER_20_162 ();
 sg13g2_fill_2 FILLER_20_166 ();
 sg13g2_decap_8 FILLER_20_189 ();
 sg13g2_fill_1 FILLER_20_245 ();
 sg13g2_fill_2 FILLER_20_260 ();
 sg13g2_decap_4 FILLER_20_298 ();
 sg13g2_fill_2 FILLER_20_302 ();
 sg13g2_fill_2 FILLER_20_318 ();
 sg13g2_fill_1 FILLER_20_320 ();
 sg13g2_fill_1 FILLER_20_330 ();
 sg13g2_fill_1 FILLER_20_350 ();
 sg13g2_fill_2 FILLER_20_391 ();
 sg13g2_fill_1 FILLER_20_393 ();
 sg13g2_decap_8 FILLER_20_398 ();
 sg13g2_decap_4 FILLER_20_405 ();
 sg13g2_fill_2 FILLER_21_0 ();
 sg13g2_fill_2 FILLER_21_38 ();
 sg13g2_fill_2 FILLER_21_66 ();
 sg13g2_fill_1 FILLER_21_68 ();
 sg13g2_fill_1 FILLER_21_122 ();
 sg13g2_decap_8 FILLER_21_198 ();
 sg13g2_fill_2 FILLER_21_205 ();
 sg13g2_fill_1 FILLER_21_211 ();
 sg13g2_fill_2 FILLER_21_220 ();
 sg13g2_fill_1 FILLER_21_226 ();
 sg13g2_decap_4 FILLER_21_241 ();
 sg13g2_fill_2 FILLER_21_245 ();
 sg13g2_decap_4 FILLER_21_307 ();
 sg13g2_fill_2 FILLER_21_337 ();
 sg13g2_decap_8 FILLER_21_365 ();
 sg13g2_decap_4 FILLER_21_404 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_4 FILLER_22_7 ();
 sg13g2_fill_1 FILLER_22_11 ();
 sg13g2_fill_2 FILLER_22_16 ();
 sg13g2_fill_2 FILLER_22_31 ();
 sg13g2_fill_1 FILLER_22_50 ();
 sg13g2_decap_8 FILLER_22_55 ();
 sg13g2_decap_4 FILLER_22_62 ();
 sg13g2_decap_4 FILLER_22_70 ();
 sg13g2_fill_2 FILLER_22_74 ();
 sg13g2_decap_4 FILLER_22_106 ();
 sg13g2_decap_8 FILLER_22_114 ();
 sg13g2_decap_8 FILLER_22_183 ();
 sg13g2_decap_4 FILLER_22_190 ();
 sg13g2_fill_2 FILLER_22_198 ();
 sg13g2_fill_1 FILLER_22_209 ();
 sg13g2_fill_2 FILLER_22_255 ();
 sg13g2_fill_1 FILLER_22_257 ();
 sg13g2_fill_2 FILLER_22_289 ();
 sg13g2_fill_1 FILLER_22_291 ();
 sg13g2_decap_4 FILLER_22_301 ();
 sg13g2_fill_2 FILLER_22_305 ();
 sg13g2_fill_2 FILLER_22_320 ();
 sg13g2_decap_8 FILLER_22_326 ();
 sg13g2_decap_8 FILLER_22_360 ();
 sg13g2_decap_4 FILLER_22_367 ();
 sg13g2_fill_2 FILLER_22_371 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_4 FILLER_23_21 ();
 sg13g2_decap_4 FILLER_23_51 ();
 sg13g2_fill_2 FILLER_23_95 ();
 sg13g2_fill_1 FILLER_23_231 ();
 sg13g2_fill_1 FILLER_23_247 ();
 sg13g2_fill_2 FILLER_23_336 ();
 sg13g2_fill_1 FILLER_23_338 ();
 sg13g2_fill_2 FILLER_23_375 ();
 sg13g2_fill_1 FILLER_23_377 ();
 sg13g2_decap_4 FILLER_23_404 ();
 sg13g2_fill_1 FILLER_23_408 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_fill_1 FILLER_24_28 ();
 sg13g2_fill_1 FILLER_24_82 ();
 sg13g2_fill_2 FILLER_24_119 ();
 sg13g2_fill_1 FILLER_24_121 ();
 sg13g2_decap_4 FILLER_24_136 ();
 sg13g2_fill_2 FILLER_24_140 ();
 sg13g2_fill_1 FILLER_24_152 ();
 sg13g2_decap_4 FILLER_24_167 ();
 sg13g2_fill_1 FILLER_24_171 ();
 sg13g2_decap_8 FILLER_24_185 ();
 sg13g2_fill_1 FILLER_24_192 ();
 sg13g2_decap_4 FILLER_24_217 ();
 sg13g2_decap_4 FILLER_24_231 ();
 sg13g2_fill_2 FILLER_24_239 ();
 sg13g2_fill_1 FILLER_24_241 ();
 sg13g2_decap_4 FILLER_24_246 ();
 sg13g2_fill_1 FILLER_24_269 ();
 sg13g2_decap_8 FILLER_24_291 ();
 sg13g2_decap_8 FILLER_24_298 ();
 sg13g2_decap_4 FILLER_24_305 ();
 sg13g2_decap_4 FILLER_24_313 ();
 sg13g2_fill_2 FILLER_24_317 ();
 sg13g2_fill_2 FILLER_24_333 ();
 sg13g2_fill_1 FILLER_24_366 ();
 sg13g2_fill_1 FILLER_24_376 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_4 FILLER_25_14 ();
 sg13g2_fill_1 FILLER_25_18 ();
 sg13g2_fill_1 FILLER_25_57 ();
 sg13g2_decap_8 FILLER_25_66 ();
 sg13g2_decap_4 FILLER_25_73 ();
 sg13g2_fill_2 FILLER_25_122 ();
 sg13g2_fill_1 FILLER_25_159 ();
 sg13g2_fill_2 FILLER_25_212 ();
 sg13g2_decap_4 FILLER_25_250 ();
 sg13g2_fill_1 FILLER_25_341 ();
 sg13g2_fill_1 FILLER_25_368 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_4 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_15 ();
 sg13g2_decap_4 FILLER_26_57 ();
 sg13g2_fill_2 FILLER_26_61 ();
 sg13g2_fill_2 FILLER_26_120 ();
 sg13g2_fill_2 FILLER_26_180 ();
 sg13g2_fill_2 FILLER_26_186 ();
 sg13g2_fill_1 FILLER_26_206 ();
 sg13g2_fill_1 FILLER_26_216 ();
 sg13g2_fill_2 FILLER_26_239 ();
 sg13g2_fill_1 FILLER_26_241 ();
 sg13g2_decap_4 FILLER_26_251 ();
 sg13g2_fill_1 FILLER_26_255 ();
 sg13g2_decap_8 FILLER_26_265 ();
 sg13g2_fill_2 FILLER_26_280 ();
 sg13g2_fill_1 FILLER_26_282 ();
 sg13g2_decap_8 FILLER_26_291 ();
 sg13g2_fill_2 FILLER_26_298 ();
 sg13g2_decap_4 FILLER_26_304 ();
 sg13g2_fill_1 FILLER_26_308 ();
 sg13g2_fill_1 FILLER_26_317 ();
 sg13g2_fill_2 FILLER_26_332 ();
 sg13g2_fill_1 FILLER_26_334 ();
 sg13g2_fill_2 FILLER_26_340 ();
 sg13g2_fill_1 FILLER_26_342 ();
 sg13g2_fill_2 FILLER_26_377 ();
 sg13g2_decap_4 FILLER_26_404 ();
 sg13g2_fill_1 FILLER_26_408 ();
 sg13g2_decap_8 FILLER_27_26 ();
 sg13g2_decap_8 FILLER_27_33 ();
 sg13g2_fill_2 FILLER_27_40 ();
 sg13g2_fill_1 FILLER_27_72 ();
 sg13g2_fill_2 FILLER_27_82 ();
 sg13g2_decap_8 FILLER_27_102 ();
 sg13g2_decap_8 FILLER_27_109 ();
 sg13g2_fill_1 FILLER_27_116 ();
 sg13g2_fill_1 FILLER_27_153 ();
 sg13g2_fill_2 FILLER_27_272 ();
 sg13g2_fill_2 FILLER_27_288 ();
 sg13g2_fill_1 FILLER_27_316 ();
 sg13g2_fill_2 FILLER_27_347 ();
 sg13g2_fill_1 FILLER_27_349 ();
 sg13g2_decap_4 FILLER_27_404 ();
 sg13g2_fill_1 FILLER_27_408 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_fill_2 FILLER_28_42 ();
 sg13g2_fill_1 FILLER_28_54 ();
 sg13g2_fill_1 FILLER_28_205 ();
 sg13g2_fill_2 FILLER_28_214 ();
 sg13g2_fill_1 FILLER_28_221 ();
 sg13g2_fill_2 FILLER_28_231 ();
 sg13g2_decap_8 FILLER_28_246 ();
 sg13g2_fill_2 FILLER_28_279 ();
 sg13g2_fill_1 FILLER_28_320 ();
 sg13g2_fill_2 FILLER_28_331 ();
 sg13g2_fill_1 FILLER_28_333 ();
 sg13g2_decap_4 FILLER_28_365 ();
 sg13g2_fill_1 FILLER_28_369 ();
 sg13g2_fill_2 FILLER_29_0 ();
 sg13g2_fill_1 FILLER_29_2 ();
 sg13g2_fill_1 FILLER_29_26 ();
 sg13g2_fill_1 FILLER_29_31 ();
 sg13g2_fill_2 FILLER_29_63 ();
 sg13g2_fill_1 FILLER_29_65 ();
 sg13g2_fill_1 FILLER_29_111 ();
 sg13g2_decap_8 FILLER_29_116 ();
 sg13g2_fill_2 FILLER_29_123 ();
 sg13g2_fill_1 FILLER_29_125 ();
 sg13g2_decap_4 FILLER_29_210 ();
 sg13g2_fill_1 FILLER_29_214 ();
 sg13g2_fill_1 FILLER_29_220 ();
 sg13g2_decap_4 FILLER_29_224 ();
 sg13g2_fill_1 FILLER_29_228 ();
 sg13g2_decap_4 FILLER_29_233 ();
 sg13g2_fill_1 FILLER_29_237 ();
 sg13g2_decap_4 FILLER_29_251 ();
 sg13g2_fill_1 FILLER_29_255 ();
 sg13g2_decap_8 FILLER_29_268 ();
 sg13g2_fill_2 FILLER_29_275 ();
 sg13g2_fill_2 FILLER_29_303 ();
 sg13g2_fill_1 FILLER_29_305 ();
 sg13g2_fill_1 FILLER_29_324 ();
 sg13g2_fill_2 FILLER_29_329 ();
 sg13g2_decap_4 FILLER_29_340 ();
 sg13g2_fill_1 FILLER_29_344 ();
 sg13g2_decap_4 FILLER_29_349 ();
 sg13g2_fill_1 FILLER_29_353 ();
 sg13g2_fill_2 FILLER_29_386 ();
 sg13g2_fill_2 FILLER_29_406 ();
 sg13g2_fill_1 FILLER_29_408 ();
 sg13g2_fill_2 FILLER_30_91 ();
 sg13g2_fill_1 FILLER_30_93 ();
 sg13g2_fill_1 FILLER_30_108 ();
 sg13g2_fill_1 FILLER_30_180 ();
 sg13g2_decap_8 FILLER_30_207 ();
 sg13g2_fill_2 FILLER_30_229 ();
 sg13g2_fill_1 FILLER_30_231 ();
 sg13g2_decap_8 FILLER_30_252 ();
 sg13g2_fill_2 FILLER_30_259 ();
 sg13g2_decap_4 FILLER_30_269 ();
 sg13g2_fill_1 FILLER_30_273 ();
 sg13g2_fill_2 FILLER_30_305 ();
 sg13g2_fill_2 FILLER_30_318 ();
 sg13g2_fill_1 FILLER_30_320 ();
 sg13g2_decap_4 FILLER_30_334 ();
 sg13g2_decap_4 FILLER_30_346 ();
 sg13g2_fill_2 FILLER_30_350 ();
 sg13g2_fill_1 FILLER_30_357 ();
 sg13g2_fill_1 FILLER_30_363 ();
 sg13g2_decap_4 FILLER_31_0 ();
 sg13g2_fill_1 FILLER_31_4 ();
 sg13g2_decap_8 FILLER_31_32 ();
 sg13g2_decap_8 FILLER_31_52 ();
 sg13g2_fill_2 FILLER_31_67 ();
 sg13g2_fill_1 FILLER_31_130 ();
 sg13g2_fill_2 FILLER_31_139 ();
 sg13g2_decap_8 FILLER_31_146 ();
 sg13g2_decap_8 FILLER_31_153 ();
 sg13g2_fill_2 FILLER_31_168 ();
 sg13g2_fill_1 FILLER_31_170 ();
 sg13g2_decap_8 FILLER_31_188 ();
 sg13g2_decap_8 FILLER_31_203 ();
 sg13g2_fill_2 FILLER_31_210 ();
 sg13g2_fill_1 FILLER_31_212 ();
 sg13g2_fill_1 FILLER_31_233 ();
 sg13g2_decap_8 FILLER_31_278 ();
 sg13g2_fill_2 FILLER_31_285 ();
 sg13g2_fill_1 FILLER_31_287 ();
 sg13g2_decap_4 FILLER_31_321 ();
 sg13g2_fill_2 FILLER_31_352 ();
 sg13g2_fill_1 FILLER_31_354 ();
 sg13g2_decap_4 FILLER_31_361 ();
 sg13g2_fill_2 FILLER_31_406 ();
 sg13g2_fill_1 FILLER_31_408 ();
 sg13g2_fill_2 FILLER_32_26 ();
 sg13g2_fill_1 FILLER_32_28 ();
 sg13g2_fill_2 FILLER_32_94 ();
 sg13g2_fill_1 FILLER_32_96 ();
 sg13g2_fill_2 FILLER_32_106 ();
 sg13g2_fill_1 FILLER_32_108 ();
 sg13g2_decap_4 FILLER_32_135 ();
 sg13g2_fill_2 FILLER_32_139 ();
 sg13g2_fill_2 FILLER_32_145 ();
 sg13g2_fill_2 FILLER_32_181 ();
 sg13g2_fill_1 FILLER_32_183 ();
 sg13g2_decap_8 FILLER_32_188 ();
 sg13g2_fill_1 FILLER_32_195 ();
 sg13g2_decap_4 FILLER_32_236 ();
 sg13g2_fill_1 FILLER_32_243 ();
 sg13g2_fill_2 FILLER_32_280 ();
 sg13g2_fill_1 FILLER_32_282 ();
 sg13g2_decap_4 FILLER_32_300 ();
 sg13g2_fill_2 FILLER_32_334 ();
 sg13g2_fill_2 FILLER_32_344 ();
 sg13g2_decap_8 FILLER_32_367 ();
 sg13g2_fill_2 FILLER_32_374 ();
 sg13g2_fill_1 FILLER_32_408 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_fill_2 FILLER_33_7 ();
 sg13g2_fill_1 FILLER_33_9 ();
 sg13g2_decap_4 FILLER_33_33 ();
 sg13g2_fill_2 FILLER_33_37 ();
 sg13g2_fill_2 FILLER_33_43 ();
 sg13g2_fill_1 FILLER_33_45 ();
 sg13g2_fill_2 FILLER_33_55 ();
 sg13g2_fill_1 FILLER_33_57 ();
 sg13g2_fill_1 FILLER_33_98 ();
 sg13g2_fill_2 FILLER_33_103 ();
 sg13g2_fill_1 FILLER_33_105 ();
 sg13g2_fill_1 FILLER_33_110 ();
 sg13g2_decap_8 FILLER_33_124 ();
 sg13g2_fill_2 FILLER_33_157 ();
 sg13g2_fill_1 FILLER_33_159 ();
 sg13g2_decap_4 FILLER_33_200 ();
 sg13g2_fill_2 FILLER_33_204 ();
 sg13g2_decap_8 FILLER_33_234 ();
 sg13g2_fill_2 FILLER_33_241 ();
 sg13g2_decap_8 FILLER_33_252 ();
 sg13g2_decap_4 FILLER_33_259 ();
 sg13g2_decap_8 FILLER_33_273 ();
 sg13g2_fill_1 FILLER_33_280 ();
 sg13g2_fill_2 FILLER_33_298 ();
 sg13g2_decap_8 FILLER_33_309 ();
 sg13g2_fill_2 FILLER_33_316 ();
 sg13g2_decap_4 FILLER_33_342 ();
 sg13g2_decap_8 FILLER_33_364 ();
 sg13g2_decap_8 FILLER_33_371 ();
 sg13g2_fill_1 FILLER_33_378 ();
 sg13g2_decap_8 FILLER_34_26 ();
 sg13g2_decap_4 FILLER_34_33 ();
 sg13g2_fill_2 FILLER_34_37 ();
 sg13g2_decap_4 FILLER_34_49 ();
 sg13g2_fill_1 FILLER_34_53 ();
 sg13g2_decap_8 FILLER_34_121 ();
 sg13g2_fill_2 FILLER_34_132 ();
 sg13g2_fill_2 FILLER_34_148 ();
 sg13g2_fill_2 FILLER_34_169 ();
 sg13g2_fill_1 FILLER_34_171 ();
 sg13g2_decap_8 FILLER_34_198 ();
 sg13g2_fill_2 FILLER_34_205 ();
 sg13g2_fill_1 FILLER_34_207 ();
 sg13g2_fill_2 FILLER_34_230 ();
 sg13g2_decap_8 FILLER_34_277 ();
 sg13g2_fill_2 FILLER_34_311 ();
 sg13g2_decap_8 FILLER_34_331 ();
 sg13g2_fill_2 FILLER_34_338 ();
 sg13g2_fill_1 FILLER_34_340 ();
 sg13g2_fill_1 FILLER_34_345 ();
 sg13g2_decap_4 FILLER_34_359 ();
 sg13g2_fill_1 FILLER_34_363 ();
 sg13g2_decap_4 FILLER_35_0 ();
 sg13g2_fill_1 FILLER_35_4 ();
 sg13g2_fill_2 FILLER_35_79 ();
 sg13g2_fill_1 FILLER_35_81 ();
 sg13g2_fill_1 FILLER_35_231 ();
 sg13g2_decap_4 FILLER_35_253 ();
 sg13g2_decap_4 FILLER_35_283 ();
 sg13g2_fill_2 FILLER_35_293 ();
 sg13g2_fill_2 FILLER_35_312 ();
 sg13g2_fill_1 FILLER_35_314 ();
 sg13g2_fill_1 FILLER_35_340 ();
 sg13g2_decap_8 FILLER_35_353 ();
 sg13g2_decap_4 FILLER_35_360 ();
 sg13g2_fill_2 FILLER_35_364 ();
 sg13g2_decap_4 FILLER_35_370 ();
 sg13g2_fill_1 FILLER_35_374 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_fill_2 FILLER_36_7 ();
 sg13g2_fill_1 FILLER_36_9 ();
 sg13g2_fill_2 FILLER_36_14 ();
 sg13g2_fill_1 FILLER_36_16 ();
 sg13g2_decap_4 FILLER_36_27 ();
 sg13g2_fill_1 FILLER_36_31 ();
 sg13g2_fill_2 FILLER_36_36 ();
 sg13g2_fill_1 FILLER_36_38 ();
 sg13g2_fill_2 FILLER_36_52 ();
 sg13g2_fill_1 FILLER_36_54 ();
 sg13g2_decap_4 FILLER_36_59 ();
 sg13g2_decap_4 FILLER_36_97 ();
 sg13g2_fill_2 FILLER_36_101 ();
 sg13g2_decap_4 FILLER_36_130 ();
 sg13g2_fill_1 FILLER_36_144 ();
 sg13g2_fill_2 FILLER_36_153 ();
 sg13g2_fill_1 FILLER_36_177 ();
 sg13g2_fill_2 FILLER_36_188 ();
 sg13g2_decap_8 FILLER_36_197 ();
 sg13g2_decap_8 FILLER_36_227 ();
 sg13g2_decap_4 FILLER_36_234 ();
 sg13g2_fill_2 FILLER_36_238 ();
 sg13g2_decap_8 FILLER_36_244 ();
 sg13g2_decap_4 FILLER_36_251 ();
 sg13g2_fill_2 FILLER_36_255 ();
 sg13g2_decap_4 FILLER_36_267 ();
 sg13g2_fill_2 FILLER_36_275 ();
 sg13g2_fill_1 FILLER_36_277 ();
 sg13g2_decap_8 FILLER_36_299 ();
 sg13g2_decap_8 FILLER_36_306 ();
 sg13g2_fill_2 FILLER_36_313 ();
 sg13g2_fill_1 FILLER_36_315 ();
 sg13g2_decap_8 FILLER_36_335 ();
 sg13g2_fill_1 FILLER_36_342 ();
 sg13g2_fill_2 FILLER_36_348 ();
 sg13g2_decap_4 FILLER_36_382 ();
 sg13g2_fill_2 FILLER_36_386 ();
 sg13g2_decap_4 FILLER_36_405 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_fill_2 FILLER_37_70 ();
 sg13g2_fill_1 FILLER_37_72 ();
 sg13g2_fill_2 FILLER_37_86 ();
 sg13g2_decap_4 FILLER_37_114 ();
 sg13g2_fill_1 FILLER_37_132 ();
 sg13g2_fill_1 FILLER_37_211 ();
 sg13g2_decap_4 FILLER_37_248 ();
 sg13g2_decap_4 FILLER_37_256 ();
 sg13g2_fill_1 FILLER_37_260 ();
 sg13g2_decap_8 FILLER_37_271 ();
 sg13g2_decap_8 FILLER_37_278 ();
 sg13g2_decap_8 FILLER_37_285 ();
 sg13g2_decap_8 FILLER_37_292 ();
 sg13g2_decap_8 FILLER_37_299 ();
 sg13g2_decap_8 FILLER_37_306 ();
 sg13g2_decap_4 FILLER_37_313 ();
 sg13g2_fill_2 FILLER_37_336 ();
 sg13g2_fill_1 FILLER_37_338 ();
 sg13g2_decap_4 FILLER_37_405 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_4 FILLER_38_60 ();
 sg13g2_decap_4 FILLER_38_68 ();
 sg13g2_decap_4 FILLER_38_76 ();
 sg13g2_fill_1 FILLER_38_84 ();
 sg13g2_fill_1 FILLER_38_122 ();
 sg13g2_fill_2 FILLER_38_140 ();
 sg13g2_fill_1 FILLER_38_142 ();
 sg13g2_fill_1 FILLER_38_151 ();
 sg13g2_decap_4 FILLER_38_164 ();
 sg13g2_decap_4 FILLER_38_172 ();
 sg13g2_fill_2 FILLER_38_180 ();
 sg13g2_fill_1 FILLER_38_182 ();
 sg13g2_decap_8 FILLER_38_200 ();
 sg13g2_fill_2 FILLER_38_207 ();
 sg13g2_fill_1 FILLER_38_222 ();
 sg13g2_fill_1 FILLER_38_227 ();
 sg13g2_decap_4 FILLER_38_284 ();
 sg13g2_decap_4 FILLER_38_292 ();
 sg13g2_fill_2 FILLER_38_301 ();
 sg13g2_fill_1 FILLER_38_303 ();
 sg13g2_fill_2 FILLER_38_308 ();
 sg13g2_fill_2 FILLER_38_368 ();
 sg13g2_fill_1 FILLER_38_370 ();
 sg13g2_fill_1 FILLER_38_408 ();
 assign uio_oe[0] = net61;
 assign uio_oe[1] = net62;
 assign uio_oe[2] = net63;
 assign uio_oe[3] = net64;
 assign uio_oe[4] = net65;
 assign uio_oe[5] = net66;
 assign uio_oe[6] = net67;
 assign uio_oe[7] = net68;
 assign uio_out[0] = net69;
 assign uio_out[1] = net70;
 assign uio_out[2] = net71;
 assign uio_out[3] = net72;
 assign uio_out[4] = net73;
 assign uio_out[5] = net74;
 assign uio_out[6] = net75;
 assign uio_out[7] = net76;
endmodule

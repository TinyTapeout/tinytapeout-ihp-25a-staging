module tt_um_wokwi_group_13 (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire \proj_10.net11 ;
 wire \proj_10.net12 ;
 wire \proj_10.net13 ;
 wire \proj_10.net14 ;
 wire \proj_10.net15 ;
 wire \proj_10.net16 ;
 wire \proj_10.net17 ;
 wire \proj_10.net18 ;
 wire \proj_10.net24 ;
 wire \proj_10.net25 ;
 wire \proj_10.net26 ;
 wire \proj_10.net27 ;
 wire \proj_10.net28 ;
 wire \proj_10.net29 ;
 wire \proj_10.net30 ;
 wire \proj_10.net31 ;
 wire \proj_10.net32 ;
 wire \proj_10.net33 ;
 wire \proj_10.net34 ;
 wire \proj_10.net35 ;
 wire \proj_10.net36 ;
 wire \proj_10.net37 ;
 wire \proj_10.net38 ;
 wire \proj_10.net39 ;
 wire \proj_10.net40 ;
 wire \proj_10.net41 ;
 wire \proj_10.net42 ;
 wire \proj_10.net43 ;
 wire \proj_10.net44 ;
 wire \proj_10.net45 ;
 wire \proj_10.net46 ;
 wire \proj_10.net47 ;
 wire \proj_10.net48 ;
 wire \proj_10.net49 ;
 wire \proj_10.net50 ;
 wire \proj_10.net51 ;
 wire \proj_10.net52 ;
 wire \proj_10.net53 ;
 wire \proj_10.net54 ;
 wire \proj_10.net55 ;
 wire \proj_10.net56 ;
 wire \proj_10.net57 ;
 wire \proj_10.net59 ;
 wire \proj_10.net60 ;
 wire \proj_10.net61 ;
 wire \proj_10.net62 ;
 wire \proj_10.net63 ;
 wire \proj_10.net64 ;
 wire \proj_10.net66 ;
 wire \proj_10.net69 ;
 wire \proj_10.net71 ;
 wire \proj_10.net72 ;
 wire \proj_10.net73 ;
 wire \proj_10.net74 ;
 wire \proj_10.net75 ;
 wire \proj_10.net76 ;
 wire \proj_10.net77 ;
 wire \proj_10.net78 ;
 wire \proj_10.net79 ;
 wire \proj_10.net80 ;
 wire \proj_10.net82 ;
 wire \proj_10.net83 ;
 wire \proj_10.net85 ;
 wire \proj_10.net87 ;
 wire \proj_10.net89 ;
 wire \proj_10.net92 ;
 wire \proj_10.net93 ;
 wire \proj_10.net94 ;
 wire \proj_10.net95 ;
 wire \proj_10.net96 ;
 wire \proj_11.net10 ;
 wire \proj_11.net11 ;
 wire \proj_11.net12 ;
 wire \proj_11.net9 ;
 wire \proj_12.net10 ;
 wire \proj_12.net11 ;
 wire \proj_12.net17 ;
 wire \proj_12.net19 ;
 wire \proj_12.net20 ;
 wire \proj_12.net7 ;
 wire \proj_12.net8 ;
 wire \proj_12.net9 ;
 wire \proj_13.net10 ;
 wire \proj_13.net11 ;
 wire \proj_13.net12 ;
 wire \proj_13.net13 ;
 wire \proj_13.net14 ;
 wire \proj_13.net15 ;
 wire \proj_13.net16 ;
 wire \proj_13.net22 ;
 wire \proj_13.net23 ;
 wire \proj_13.net24 ;
 wire \proj_13.net25 ;
 wire \proj_13.net26 ;
 wire \proj_13.net27 ;
 wire \proj_13.net28 ;
 wire \proj_13.net29 ;
 wire \proj_13.net30 ;
 wire \proj_13.net31 ;
 wire \proj_13.net32 ;
 wire \proj_13.net33 ;
 wire \proj_13.net34 ;
 wire \proj_13.net35 ;
 wire \proj_13.net36 ;
 wire \proj_13.net37 ;
 wire \proj_13.net38 ;
 wire \proj_13.net39 ;
 wire \proj_13.net40 ;
 wire \proj_13.net41 ;
 wire \proj_13.net42 ;
 wire \proj_13.net43 ;
 wire \proj_13.net44 ;
 wire \proj_14.net3 ;
 wire \proj_15.net10 ;
 wire \proj_15.net11 ;
 wire \proj_15.net12 ;
 wire \proj_15.net9 ;
 wire \proj__0.net10 ;
 wire \proj__0.net11 ;
 wire \proj__1.net10 ;
 wire \proj__1.net11 ;
 wire \proj__1.net12 ;
 wire \proj__1.net13 ;
 wire \proj__2.net12 ;
 wire \proj__2.net13 ;
 wire \proj__2.net14 ;
 wire \proj__2.net6 ;
 wire \proj__3.net14 ;
 wire \proj__3.net15 ;
 wire \proj__3.net16 ;
 wire \proj__3.net17 ;
 wire \proj__3.net18 ;
 wire \proj__3.net19 ;
 wire \proj__3.net2 ;
 wire \proj__3.net20 ;
 wire \proj__3.net21 ;
 wire \proj__3.net22 ;
 wire \proj__3.net23 ;
 wire \proj__3.net24 ;
 wire \proj__3.net25 ;
 wire \proj__3.net26 ;
 wire \proj__3.net27 ;
 wire \proj__3.net28 ;
 wire \proj__3.net29 ;
 wire \proj__3.net3 ;
 wire \proj__3.net4 ;
 wire \proj__3.net5 ;
 wire \proj__3.net6 ;
 wire \proj__3.net7 ;
 wire \proj__3.net8 ;
 wire \proj__4.net100 ;
 wire \proj__4.net101 ;
 wire \proj__4.net102 ;
 wire \proj__4.net103 ;
 wire \proj__4.net104 ;
 wire \proj__4.net105 ;
 wire \proj__4.net106 ;
 wire \proj__4.net109 ;
 wire \proj__4.net110 ;
 wire \proj__4.net111 ;
 wire \proj__4.net112 ;
 wire \proj__4.net113 ;
 wire \proj__4.net114 ;
 wire \proj__4.net115 ;
 wire \proj__4.net116 ;
 wire \proj__4.net117 ;
 wire \proj__4.net118 ;
 wire \proj__4.net119 ;
 wire \proj__4.net120 ;
 wire \proj__4.net121 ;
 wire \proj__4.net122 ;
 wire \proj__4.net125 ;
 wire \proj__4.net126 ;
 wire \proj__4.net127 ;
 wire \proj__4.net128 ;
 wire \proj__4.net129 ;
 wire \proj__4.net130 ;
 wire \proj__4.net131 ;
 wire \proj__4.net132 ;
 wire \proj__4.net133 ;
 wire \proj__4.net134 ;
 wire \proj__4.net135 ;
 wire \proj__4.net136 ;
 wire \proj__4.net137 ;
 wire \proj__4.net138 ;
 wire \proj__4.net139 ;
 wire \proj__4.net140 ;
 wire \proj__4.net16 ;
 wire \proj__4.net17 ;
 wire \proj__4.net18 ;
 wire \proj__4.net2 ;
 wire \proj__4.net20 ;
 wire \proj__4.net21 ;
 wire \proj__4.net22 ;
 wire \proj__4.net23 ;
 wire \proj__4.net24 ;
 wire \proj__4.net25 ;
 wire \proj__4.net26 ;
 wire \proj__4.net27 ;
 wire \proj__4.net28 ;
 wire \proj__4.net29 ;
 wire \proj__4.net3 ;
 wire \proj__4.net30 ;
 wire \proj__4.net31 ;
 wire \proj__4.net32 ;
 wire \proj__4.net33 ;
 wire \proj__4.net34 ;
 wire \proj__4.net35 ;
 wire \proj__4.net36 ;
 wire \proj__4.net37 ;
 wire \proj__4.net38 ;
 wire \proj__4.net4 ;
 wire \proj__4.net40 ;
 wire \proj__4.net41 ;
 wire \proj__4.net42 ;
 wire \proj__4.net44 ;
 wire \proj__4.net46 ;
 wire \proj__4.net47 ;
 wire \proj__4.net48 ;
 wire \proj__4.net49 ;
 wire \proj__4.net5 ;
 wire \proj__4.net50 ;
 wire \proj__4.net51 ;
 wire \proj__4.net52 ;
 wire \proj__4.net53 ;
 wire \proj__4.net54 ;
 wire \proj__4.net55 ;
 wire \proj__4.net56 ;
 wire \proj__4.net57 ;
 wire \proj__4.net58 ;
 wire \proj__4.net6 ;
 wire \proj__4.net60 ;
 wire \proj__4.net62 ;
 wire \proj__4.net63 ;
 wire \proj__4.net64 ;
 wire \proj__4.net65 ;
 wire \proj__4.net66 ;
 wire \proj__4.net67 ;
 wire \proj__4.net68 ;
 wire \proj__4.net69 ;
 wire \proj__4.net7 ;
 wire \proj__4.net70 ;
 wire \proj__4.net71 ;
 wire \proj__4.net72 ;
 wire \proj__4.net73 ;
 wire \proj__4.net74 ;
 wire \proj__4.net77 ;
 wire \proj__4.net78 ;
 wire \proj__4.net79 ;
 wire \proj__4.net8 ;
 wire \proj__4.net80 ;
 wire \proj__4.net81 ;
 wire \proj__4.net82 ;
 wire \proj__4.net83 ;
 wire \proj__4.net84 ;
 wire \proj__4.net85 ;
 wire \proj__4.net86 ;
 wire \proj__4.net87 ;
 wire \proj__4.net88 ;
 wire \proj__4.net89 ;
 wire \proj__4.net9 ;
 wire \proj__4.net90 ;
 wire \proj__4.net92 ;
 wire \proj__4.net94 ;
 wire \proj__4.net95 ;
 wire \proj__4.net96 ;
 wire \proj__4.net97 ;
 wire \proj__4.net98 ;
 wire \proj__4.net99 ;
 wire \proj__5.net12 ;
 wire \proj__5.net13 ;
 wire \proj__5.net14 ;
 wire \proj__5.net6 ;
 wire \proj__6.net10 ;
 wire \proj__6.net100 ;
 wire \proj__6.net101 ;
 wire \proj__6.net102 ;
 wire \proj__6.net103 ;
 wire \proj__6.net104 ;
 wire \proj__6.net105 ;
 wire \proj__6.net106 ;
 wire \proj__6.net107 ;
 wire \proj__6.net11 ;
 wire \proj__6.net12 ;
 wire \proj__6.net13 ;
 wire \proj__6.net14 ;
 wire \proj__6.net15 ;
 wire \proj__6.net16 ;
 wire \proj__6.net17 ;
 wire \proj__6.net20 ;
 wire \proj__6.net21 ;
 wire \proj__6.net23 ;
 wire \proj__6.net24 ;
 wire \proj__6.net25 ;
 wire \proj__6.net26 ;
 wire \proj__6.net27 ;
 wire \proj__6.net28 ;
 wire \proj__6.net29 ;
 wire \proj__6.net30 ;
 wire \proj__6.net31 ;
 wire \proj__6.net32 ;
 wire \proj__6.net33 ;
 wire \proj__6.net34 ;
 wire \proj__6.net35 ;
 wire \proj__6.net36 ;
 wire \proj__6.net37 ;
 wire \proj__6.net38 ;
 wire \proj__6.net39 ;
 wire \proj__6.net40 ;
 wire \proj__6.net41 ;
 wire \proj__6.net42 ;
 wire \proj__6.net43 ;
 wire \proj__6.net44 ;
 wire \proj__6.net45 ;
 wire \proj__6.net46 ;
 wire \proj__6.net47 ;
 wire \proj__6.net48 ;
 wire \proj__6.net49 ;
 wire \proj__6.net50 ;
 wire \proj__6.net51 ;
 wire \proj__6.net52 ;
 wire \proj__6.net53 ;
 wire \proj__6.net54 ;
 wire \proj__6.net55 ;
 wire \proj__6.net56 ;
 wire \proj__6.net57 ;
 wire \proj__6.net58 ;
 wire \proj__6.net59 ;
 wire \proj__6.net60 ;
 wire \proj__6.net61 ;
 wire \proj__6.net62 ;
 wire \proj__6.net63 ;
 wire \proj__6.net64 ;
 wire \proj__6.net65 ;
 wire \proj__6.net66 ;
 wire \proj__6.net72 ;
 wire \proj__6.net74 ;
 wire \proj__6.net75 ;
 wire \proj__6.net76 ;
 wire \proj__6.net77 ;
 wire \proj__6.net78 ;
 wire \proj__6.net79 ;
 wire \proj__6.net80 ;
 wire \proj__6.net81 ;
 wire \proj__6.net82 ;
 wire \proj__6.net83 ;
 wire \proj__6.net84 ;
 wire \proj__6.net85 ;
 wire \proj__6.net86 ;
 wire \proj__6.net87 ;
 wire \proj__6.net88 ;
 wire \proj__6.net90 ;
 wire \proj__6.net91 ;
 wire \proj__6.net92 ;
 wire \proj__6.net93 ;
 wire \proj__6.net94 ;
 wire \proj__6.net95 ;
 wire \proj__6.net96 ;
 wire \proj__6.net97 ;
 wire \proj__6.net98 ;
 wire \proj__6.net99 ;
 wire \proj__7.net11 ;
 wire \proj__7.net12 ;
 wire \proj__7.net4 ;
 wire \proj__7.net5 ;
 wire \proj__9.net15 ;
 wire \proj__9.net16 ;
 wire \proj__9.net18 ;
 wire \proj__9.net19 ;
 wire \proj__9.net20 ;
 wire \proj__9.net5 ;
 wire \proj__9.net6 ;
 wire \proj__9.net7 ;
 wire \proj__9.net8 ;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire \proj_10.flop1/_0_ ;
 wire \proj_10.flop1/_1_ ;
 wire net151;
 wire net152;
 wire \proj_10.flop1/notq ;
 wire \proj_10.flop10/_0_ ;
 wire \proj_10.flop10/_1_ ;
 wire net153;
 wire net154;
 wire \proj_10.flop10/notq ;
 wire \proj_10.flop11/_0_ ;
 wire \proj_10.flop11/_1_ ;
 wire net155;
 wire net156;
 wire \proj_10.flop11/notq ;
 wire \proj_10.flop12/_0_ ;
 wire \proj_10.flop12/_1_ ;
 wire net157;
 wire net158;
 wire \proj_10.flop12/notq ;
 wire \proj_10.flop13/_0_ ;
 wire \proj_10.flop13/_1_ ;
 wire net159;
 wire net213;
 wire \proj_10.flop13/notq ;
 wire \proj_10.flop14/_0_ ;
 wire \proj_10.flop14/_1_ ;
 wire net214;
 wire net215;
 wire \proj_10.flop14/notq ;
 wire \proj_10.flop2/_0_ ;
 wire \proj_10.flop2/_1_ ;
 wire net216;
 wire net217;
 wire \proj_10.flop2/notq ;
 wire \proj_10.flop3/_0_ ;
 wire \proj_10.flop3/_1_ ;
 wire net218;
 wire net219;
 wire \proj_10.flop3/notq ;
 wire \proj_10.flop4/_0_ ;
 wire \proj_10.flop4/_1_ ;
 wire net220;
 wire net221;
 wire \proj_10.flop4/notq ;
 wire \proj_10.flop5/_0_ ;
 wire \proj_10.flop5/_1_ ;
 wire net222;
 wire net223;
 wire \proj_10.flop5/notq ;
 wire \proj_10.flop6/_0_ ;
 wire \proj_10.flop6/_1_ ;
 wire net224;
 wire net225;
 wire \proj_10.flop6/notq ;
 wire \proj_10.flop7/_0_ ;
 wire \proj_10.flop7/_1_ ;
 wire net226;
 wire net227;
 wire \proj_10.flop7/notq ;
 wire \proj_10.flop8/_0_ ;
 wire \proj_10.flop8/_1_ ;
 wire net228;
 wire net229;
 wire \proj_10.flop8/notq ;
 wire \proj_10.flop9/_0_ ;
 wire \proj_10.flop9/_1_ ;
 wire net230;
 wire net231;
 wire \proj_10.flop9/notq ;
 wire \proj_12.flop1/_0_ ;
 wire \proj_12.flop1/_1_ ;
 wire net232;
 wire net233;
 wire \proj_12.flop2/_0_ ;
 wire \proj_12.flop2/_1_ ;
 wire net234;
 wire net235;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire \proj__4.flop1/notq ;
 wire net396;
 wire \proj__4.flop2/notq ;
 wire net397;
 wire \proj__4.flop3/notq ;
 wire clk_regs;
 wire \proj__4.flop4/notq ;
 wire \proj__6.flop0/_0_ ;
 wire \proj__6.flop0/_1_ ;
 wire net236;
 wire net237;
 wire \proj__6.flop0/notq ;
 wire \proj__6.flop1/_0_ ;
 wire \proj__6.flop1/_1_ ;
 wire net238;
 wire net239;
 wire \proj__6.flop1/notq ;
 wire \proj__6.flop10/_0_ ;
 wire \proj__6.flop10/_1_ ;
 wire net240;
 wire net241;
 wire \proj__6.flop10/notq ;
 wire \proj__6.flop11/_0_ ;
 wire \proj__6.flop11/_1_ ;
 wire net242;
 wire net243;
 wire \proj__6.flop11/notq ;
 wire \proj__6.flop12/_0_ ;
 wire \proj__6.flop12/_1_ ;
 wire net244;
 wire net245;
 wire \proj__6.flop12/notq ;
 wire \proj__6.flop13/_0_ ;
 wire \proj__6.flop13/_1_ ;
 wire net246;
 wire net247;
 wire \proj__6.flop13/notq ;
 wire \proj__6.flop14/_0_ ;
 wire \proj__6.flop14/_1_ ;
 wire net248;
 wire net249;
 wire \proj__6.flop14/notq ;
 wire \proj__6.flop15/_0_ ;
 wire \proj__6.flop15/_1_ ;
 wire net250;
 wire net251;
 wire \proj__6.flop15/notq ;
 wire \proj__6.flop16/_0_ ;
 wire \proj__6.flop16/_1_ ;
 wire net252;
 wire net253;
 wire \proj__6.flop16/notq ;
 wire \proj__6.flop17/_0_ ;
 wire \proj__6.flop17/_1_ ;
 wire net254;
 wire net255;
 wire \proj__6.flop17/notq ;
 wire \proj__6.flop18/_0_ ;
 wire \proj__6.flop18/_1_ ;
 wire net256;
 wire net257;
 wire \proj__6.flop18/notq ;
 wire \proj__6.flop19/_0_ ;
 wire \proj__6.flop19/_1_ ;
 wire net258;
 wire net259;
 wire \proj__6.flop19/notq ;
 wire \proj__6.flop2/_0_ ;
 wire \proj__6.flop2/_1_ ;
 wire net260;
 wire net261;
 wire \proj__6.flop2/notq ;
 wire \proj__6.flop20/_0_ ;
 wire \proj__6.flop20/_1_ ;
 wire net262;
 wire net263;
 wire \proj__6.flop20/notq ;
 wire \proj__6.flop21/_0_ ;
 wire \proj__6.flop21/_1_ ;
 wire net264;
 wire net265;
 wire \proj__6.flop21/notq ;
 wire \proj__6.flop22/_0_ ;
 wire \proj__6.flop22/_1_ ;
 wire net266;
 wire net267;
 wire \proj__6.flop22/notq ;
 wire \proj__6.flop23/_0_ ;
 wire \proj__6.flop23/_1_ ;
 wire net268;
 wire net269;
 wire \proj__6.flop23/notq ;
 wire \proj__6.flop24/_0_ ;
 wire \proj__6.flop24/_1_ ;
 wire net270;
 wire net271;
 wire \proj__6.flop24/notq ;
 wire \proj__6.flop25/_0_ ;
 wire \proj__6.flop25/_1_ ;
 wire net272;
 wire net273;
 wire \proj__6.flop25/notq ;
 wire \proj__6.flop26/_0_ ;
 wire \proj__6.flop26/_1_ ;
 wire net274;
 wire net275;
 wire \proj__6.flop26/notq ;
 wire \proj__6.flop27/_0_ ;
 wire \proj__6.flop27/_1_ ;
 wire net276;
 wire net277;
 wire \proj__6.flop27/notq ;
 wire \proj__6.flop28/_0_ ;
 wire \proj__6.flop28/_1_ ;
 wire net278;
 wire net279;
 wire \proj__6.flop28/notq ;
 wire \proj__6.flop29/_0_ ;
 wire \proj__6.flop29/_1_ ;
 wire net280;
 wire net281;
 wire \proj__6.flop29/notq ;
 wire \proj__6.flop3/_0_ ;
 wire \proj__6.flop3/_1_ ;
 wire net282;
 wire net283;
 wire \proj__6.flop3/notq ;
 wire \proj__6.flop30/_0_ ;
 wire \proj__6.flop30/_1_ ;
 wire net284;
 wire net285;
 wire \proj__6.flop30/notq ;
 wire \proj__6.flop31/_0_ ;
 wire \proj__6.flop31/_1_ ;
 wire net286;
 wire net287;
 wire \proj__6.flop31/notq ;
 wire \proj__6.flop33/_0_ ;
 wire \proj__6.flop33/_1_ ;
 wire net288;
 wire net289;
 wire \proj__6.flop33/notq ;
 wire \proj__6.flop34/_0_ ;
 wire \proj__6.flop34/_1_ ;
 wire net290;
 wire net291;
 wire \proj__6.flop34/notq ;
 wire \proj__6.flop35/_0_ ;
 wire \proj__6.flop35/_1_ ;
 wire net292;
 wire net293;
 wire \proj__6.flop35/notq ;
 wire \proj__6.flop36/_0_ ;
 wire \proj__6.flop36/_1_ ;
 wire net294;
 wire net295;
 wire \proj__6.flop36/notq ;
 wire \proj__6.flop37/_0_ ;
 wire \proj__6.flop37/_1_ ;
 wire net296;
 wire net297;
 wire \proj__6.flop37/notq ;
 wire \proj__6.flop38/_0_ ;
 wire \proj__6.flop38/_1_ ;
 wire net298;
 wire net299;
 wire \proj__6.flop38/notq ;
 wire \proj__6.flop39/_0_ ;
 wire \proj__6.flop39/_1_ ;
 wire net300;
 wire net301;
 wire \proj__6.flop39/notq ;
 wire \proj__6.flop4/_0_ ;
 wire \proj__6.flop4/_1_ ;
 wire net302;
 wire net303;
 wire \proj__6.flop4/notq ;
 wire \proj__6.flop40/_0_ ;
 wire \proj__6.flop40/_1_ ;
 wire net304;
 wire net305;
 wire \proj__6.flop40/notq ;
 wire \proj__6.flop5/_0_ ;
 wire \proj__6.flop5/_1_ ;
 wire net306;
 wire net307;
 wire \proj__6.flop5/notq ;
 wire \proj__6.flop6/_0_ ;
 wire \proj__6.flop6/_1_ ;
 wire net308;
 wire net309;
 wire \proj__6.flop6/notq ;
 wire \proj__6.flop7/_0_ ;
 wire \proj__6.flop7/_1_ ;
 wire net310;
 wire net311;
 wire \proj__6.flop7/notq ;
 wire \proj__6.flop8/_0_ ;
 wire \proj__6.flop8/_1_ ;
 wire net312;
 wire net313;
 wire \proj__6.flop8/notq ;
 wire \proj__6.flop9/_0_ ;
 wire \proj__6.flop9/_1_ ;
 wire net314;
 wire net315;
 wire \proj__6.flop9/notq ;
 wire \proj__9.flop1/_0_ ;
 wire \proj__9.flop1/_1_ ;
 wire net316;
 wire net317;
 wire \proj__9.flop1/notq ;
 wire \proj__9.flop2/_0_ ;
 wire \proj__9.flop2/_1_ ;
 wire net318;
 wire net319;
 wire \proj__9.flop2/notq ;
 wire \proj__9.flop3/_0_ ;
 wire \proj__9.flop3/_1_ ;
 wire net320;
 wire net321;
 wire \proj__9.flop3/notq ;
 wire \proj__9.flop4/_0_ ;
 wire \proj__9.flop4/_1_ ;
 wire net322;
 wire net323;
 wire \proj__9.flop4/notq ;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;
 wire clknet_0_clk_regs;
 wire clknet_2_0__leaf_clk_regs;
 wire clknet_2_1__leaf_clk_regs;
 wire clknet_2_2__leaf_clk_regs;
 wire clknet_2_3__leaf_clk_regs;
 wire clknet_0__015_;
 wire clknet_1_0__leaf__015_;
 wire clknet_1_1__leaf__015_;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;

 sg13g2_inv_1 _268_ (.Y(_061_),
    .A(net6));
 sg13g2_inv_1 _269_ (.Y(_062_),
    .A(net209));
 sg13g2_inv_1 _270_ (.Y(_063_),
    .A(net199));
 sg13g2_inv_1 _271_ (.Y(_064_),
    .A(\proj__0.net10 ));
 sg13g2_inv_1 _272_ (.Y(_065_),
    .A(\proj__0.net11 ));
 sg13g2_nor2b_1 _273_ (.A(net4),
    .B_N(net3),
    .Y(_066_));
 sg13g2_nor2_1 _274_ (.A(net6),
    .B(net5),
    .Y(_067_));
 sg13g2_or2_1 _275_ (.X(_068_),
    .B(net5),
    .A(net6));
 sg13g2_and2_2 _276_ (.A(_066_),
    .B(_067_),
    .X(_069_));
 sg13g2_nand2_2 _277_ (.Y(_070_),
    .A(net4),
    .B(net3));
 sg13g2_a22oi_1 _278_ (.Y(_071_),
    .B1(_068_),
    .B2(_070_),
    .A2(net3),
    .A1(_061_));
 sg13g2_or2_1 _279_ (.X(_072_),
    .B(_071_),
    .A(_069_));
 sg13g2_nand2_1 _280_ (.Y(_073_),
    .A(net185),
    .B(_072_));
 sg13g2_nor2b_1 _281_ (.A(net6),
    .B_N(net5),
    .Y(_074_));
 sg13g2_nand2b_1 _282_ (.Y(_000_),
    .B(net5),
    .A_N(net6));
 sg13g2_nor3_2 _283_ (.A(net4),
    .B(net3),
    .C(_000_),
    .Y(_001_));
 sg13g2_nand2_2 _284_ (.Y(_002_),
    .A(net6),
    .B(net5));
 sg13g2_and3_2 _285_ (.X(_003_),
    .A(net6),
    .B(net5),
    .C(_066_));
 sg13g2_nor3_2 _286_ (.A(net4),
    .B(net3),
    .C(_002_),
    .Y(_004_));
 sg13g2_nor2b_1 _287_ (.A(net3),
    .B_N(net4),
    .Y(_005_));
 sg13g2_and2_2 _288_ (.A(_074_),
    .B(_005_),
    .X(_006_));
 sg13g2_a22oi_1 _289_ (.Y(_007_),
    .B1(_006_),
    .B2(\proj__6.net17 ),
    .A2(_004_),
    .A1(\proj_12.net11 ));
 sg13g2_nor2_1 _290_ (.A(_070_),
    .B(_000_),
    .Y(_008_));
 sg13g2_nor2b_1 _291_ (.A(net5),
    .B_N(net6),
    .Y(_009_));
 sg13g2_and2_2 _292_ (.A(_005_),
    .B(_009_),
    .X(_010_));
 sg13g2_a22oi_1 _293_ (.Y(_011_),
    .B1(_008_),
    .B2(\proj__7.net5 ),
    .A2(_003_),
    .A1(clknet_1_1__leaf_clk));
 sg13g2_a22oi_1 _294_ (.Y(_012_),
    .B1(_010_),
    .B2(\proj_10.net18 ),
    .A2(_001_),
    .A1(\proj__4.net9 ));
 sg13g2_nand4_1 _295_ (.B(_007_),
    .C(_011_),
    .A(_073_),
    .Y(uo_out[7]),
    .D(_012_));
 sg13g2_nor3_2 _296_ (.A(net4),
    .B(net3),
    .C(_068_),
    .Y(_013_));
 sg13g2_nor2b_1 _297_ (.A(_002_),
    .B_N(_005_),
    .Y(_014_));
 sg13g2_a21oi_1 _298_ (.A1(\proj_14.net3 ),
    .A2(_014_),
    .Y(_015_),
    .B1(_013_));
 sg13g2_a22oi_1 _299_ (.Y(_016_),
    .B1(_008_),
    .B2(\proj__7.net4 ),
    .A2(_004_),
    .A1(\proj_12.net7 ));
 sg13g2_nor2b_2 _300_ (.A(_070_),
    .B_N(_009_),
    .Y(_017_));
 sg13g2_a22oi_1 _301_ (.Y(_018_),
    .B1(_017_),
    .B2(\proj_11.net9 ),
    .A2(_001_),
    .A1(\proj__4.net2 ));
 sg13g2_and2_1 _302_ (.A(_066_),
    .B(_009_),
    .X(_019_));
 sg13g2_nand3_1 _303_ (.B(_067_),
    .C(_005_),
    .A(\proj__2.net6 ),
    .Y(_020_));
 sg13g2_and2_1 _304_ (.A(_066_),
    .B(_074_),
    .X(_021_));
 sg13g2_nor2_2 _305_ (.A(_070_),
    .B(_002_),
    .Y(_022_));
 sg13g2_nor2_2 _306_ (.A(_068_),
    .B(_070_),
    .Y(_023_));
 sg13g2_a22oi_1 _307_ (.Y(_024_),
    .B1(_023_),
    .B2(\proj__3.net2 ),
    .A2(_003_),
    .A1(\proj_13.net10 ));
 sg13g2_a22oi_1 _308_ (.Y(_025_),
    .B1(_006_),
    .B2(\proj__6.net10 ),
    .A2(_069_),
    .A1(\proj__1.net10 ));
 sg13g2_a22oi_1 _309_ (.Y(_026_),
    .B1(_022_),
    .B2(\proj_15.net9 ),
    .A2(_021_),
    .A1(\proj__5.net6 ));
 sg13g2_a22oi_1 _310_ (.Y(_027_),
    .B1(_019_),
    .B2(\proj__9.net5 ),
    .A2(_010_),
    .A1(\proj_10.net11 ));
 sg13g2_and4_1 _311_ (.A(clknet_1_1__leaf__015_),
    .B(_016_),
    .C(_025_),
    .D(_026_),
    .X(_028_));
 sg13g2_and4_1 _312_ (.A(_018_),
    .B(_020_),
    .C(_024_),
    .D(_027_),
    .X(_029_));
 sg13g2_a22oi_1 _313_ (.Y(uo_out[0]),
    .B1(_028_),
    .B2(_029_),
    .A2(_013_),
    .A1(_062_));
 sg13g2_a22oi_1 _314_ (.Y(_030_),
    .B1(_023_),
    .B2(\proj__3.net3 ),
    .A2(_001_),
    .A1(\proj__4.net3 ));
 sg13g2_a22oi_1 _315_ (.Y(_031_),
    .B1(_022_),
    .B2(\proj_15.net10 ),
    .A2(_017_),
    .A1(\proj_11.net10 ));
 sg13g2_a22oi_1 _316_ (.Y(_032_),
    .B1(_019_),
    .B2(\proj__9.net6 ),
    .A2(_010_),
    .A1(\proj_10.net12 ));
 sg13g2_a22oi_1 _317_ (.Y(_033_),
    .B1(_006_),
    .B2(\proj__6.net11 ),
    .A2(_069_),
    .A1(\proj__1.net11 ));
 sg13g2_and2_1 _318_ (.A(_032_),
    .B(_033_),
    .X(_034_));
 sg13g2_a22oi_1 _319_ (.Y(_035_),
    .B1(_004_),
    .B2(\proj_12.net8 ),
    .A2(_003_),
    .A1(\proj_13.net11 ));
 sg13g2_and4_1 _320_ (.A(clknet_1_0__leaf__015_),
    .B(_030_),
    .C(_031_),
    .D(_035_),
    .X(_036_));
 sg13g2_a22oi_1 _321_ (.Y(uo_out[1]),
    .B1(_034_),
    .B2(_036_),
    .A2(_013_),
    .A1(_063_));
 sg13g2_and2_1 _322_ (.A(\proj__9.net7 ),
    .B(_019_),
    .X(_037_));
 sg13g2_a221oi_1 _323_ (.B2(\proj__3.net4 ),
    .C1(_037_),
    .B1(_023_),
    .A1(\proj_12.net9 ),
    .Y(_038_),
    .A2(_004_));
 sg13g2_a22oi_1 _324_ (.Y(_039_),
    .B1(_017_),
    .B2(\proj_11.net11 ),
    .A2(_010_),
    .A1(\proj_10.net13 ));
 sg13g2_a22oi_1 _325_ (.Y(_040_),
    .B1(_003_),
    .B2(\proj_13.net12 ),
    .A2(_001_),
    .A1(\proj__4.net4 ));
 sg13g2_a22oi_1 _326_ (.Y(_041_),
    .B1(_022_),
    .B2(\proj_15.net11 ),
    .A2(_006_),
    .A1(\proj__6.net12 ));
 sg13g2_and4_1 _327_ (.A(clknet_1_0__leaf__015_),
    .B(_039_),
    .C(_040_),
    .D(_041_),
    .X(_042_));
 sg13g2_a22oi_1 _328_ (.Y(uo_out[2]),
    .B1(_038_),
    .B2(_042_),
    .A2(_013_),
    .A1(_064_));
 sg13g2_and2_1 _329_ (.A(\proj__9.net8 ),
    .B(_019_),
    .X(_043_));
 sg13g2_a22oi_1 _330_ (.Y(_044_),
    .B1(_010_),
    .B2(\proj_10.net14 ),
    .A2(_004_),
    .A1(\proj_12.net10 ));
 sg13g2_a221oi_1 _331_ (.B2(\proj_11.net12 ),
    .C1(_043_),
    .B1(_017_),
    .A1(\proj_13.net13 ),
    .Y(_045_),
    .A2(_003_));
 sg13g2_a21oi_1 _332_ (.A1(\proj__6.net13 ),
    .A2(_006_),
    .Y(_046_),
    .B1(_013_));
 sg13g2_a22oi_1 _333_ (.Y(_047_),
    .B1(_023_),
    .B2(\proj__3.net5 ),
    .A2(_069_),
    .A1(\proj__1.net12 ));
 sg13g2_a22oi_1 _334_ (.Y(_048_),
    .B1(_022_),
    .B2(\proj_15.net12 ),
    .A2(_001_),
    .A1(\proj__4.net5 ));
 sg13g2_and4_1 _335_ (.A(_044_),
    .B(_046_),
    .C(_047_),
    .D(_048_),
    .X(_049_));
 sg13g2_a22oi_1 _336_ (.Y(uo_out[3]),
    .B1(_045_),
    .B2(_049_),
    .A2(_013_),
    .A1(_065_));
 sg13g2_o21ai_1 _337_ (.B1(net192),
    .Y(_050_),
    .A1(_071_),
    .A2(_004_));
 sg13g2_a22oi_1 _338_ (.Y(_051_),
    .B1(_023_),
    .B2(\proj__3.net6 ),
    .A2(_069_),
    .A1(\proj__1.net13 ));
 sg13g2_a22oi_1 _339_ (.Y(_052_),
    .B1(_003_),
    .B2(\proj_13.net14 ),
    .A2(_001_),
    .A1(\proj__4.net6 ));
 sg13g2_a22oi_1 _340_ (.Y(_053_),
    .B1(_010_),
    .B2(\proj_10.net15 ),
    .A2(_006_),
    .A1(\proj__6.net14 ));
 sg13g2_nand4_1 _341_ (.B(_051_),
    .C(_052_),
    .A(_050_),
    .Y(uo_out[4]),
    .D(_053_));
 sg13g2_a22oi_1 _342_ (.Y(_054_),
    .B1(_023_),
    .B2(\proj__3.net7 ),
    .A2(_001_),
    .A1(\proj__4.net7 ));
 sg13g2_a22oi_1 _343_ (.Y(_055_),
    .B1(_006_),
    .B2(\proj__6.net15 ),
    .A2(_071_),
    .A1(net190));
 sg13g2_a22oi_1 _344_ (.Y(_056_),
    .B1(_010_),
    .B2(\proj_10.net16 ),
    .A2(_003_),
    .A1(\proj_13.net15 ));
 sg13g2_nand3_1 _345_ (.B(_055_),
    .C(_056_),
    .A(_054_),
    .Y(uo_out[5]));
 sg13g2_nand2_1 _346_ (.Y(_057_),
    .A(net187),
    .B(_072_));
 sg13g2_nand2_1 _347_ (.Y(_058_),
    .A(\proj__4.net8 ),
    .B(_001_));
 sg13g2_a22oi_1 _348_ (.Y(_059_),
    .B1(_010_),
    .B2(\proj_10.net17 ),
    .A2(_003_),
    .A1(\proj_13.net16 ));
 sg13g2_a22oi_1 _349_ (.Y(_060_),
    .B1(_023_),
    .B2(\proj__3.net8 ),
    .A2(_006_),
    .A1(\proj__6.net16 ));
 sg13g2_nand4_1 _350_ (.B(_058_),
    .C(_059_),
    .A(_057_),
    .Y(uo_out[6]),
    .D(_060_));
 sg13g2_tiehi \proj__4.mux106/_0__271  (.L_HI(net324));
 sg13g2_tiehi \proj__4.mux107/_0__272  (.L_HI(net325));
 sg13g2_tiehi \proj__4.mux107/_0__273  (.L_HI(net326));
 sg13g2_tiehi \proj__4.mux108/_0__274  (.L_HI(net327));
 sg13g2_tiehi \proj__4.mux108/_0__275  (.L_HI(net328));
 sg13g2_tiehi \proj__4.mux109/_0__276  (.L_HI(net329));
 sg13g2_tiehi \proj__4.mux109/_0__277  (.L_HI(net330));
 sg13g2_tiehi \proj__4.mux110/_0__278  (.L_HI(net331));
 sg13g2_tiehi \proj__4.mux111/_0__279  (.L_HI(net332));
 sg13g2_tiehi \proj__4.mux111/_0__280  (.L_HI(net333));
 sg13g2_tiehi \proj__4.mux112/_0__281  (.L_HI(net334));
 sg13g2_tiehi \proj__4.mux112/_0__282  (.L_HI(net335));
 sg13g2_tiehi \proj__4.mux113/_0__283  (.L_HI(net336));
 sg13g2_tiehi \proj__4.mux113/_0__284  (.L_HI(net337));
 sg13g2_tiehi \proj__4.mux3/_0__285  (.L_HI(net338));
 sg13g2_tiehi \proj__4.mux32/_0__286  (.L_HI(net339));
 sg13g2_tiehi \proj__4.mux33/_0__287  (.L_HI(net340));
 sg13g2_tiehi \proj__4.mux34/_0__288  (.L_HI(net341));
 sg13g2_tiehi \proj__4.mux34/_0__289  (.L_HI(net342));
 sg13g2_tiehi \proj__4.mux38/_0__290  (.L_HI(net343));
 sg13g2_tiehi \proj__4.mux4/_0__291  (.L_HI(net344));
 sg13g2_tiehi \proj__4.mux4/_0__292  (.L_HI(net345));
 sg13g2_tiehi \proj__4.mux47/_0__293  (.L_HI(net346));
 sg13g2_tiehi \proj__4.mux47/_0__294  (.L_HI(net347));
 sg13g2_tiehi \proj__4.mux48/_0__295  (.L_HI(net348));
 sg13g2_tiehi \proj__4.mux50/_0__296  (.L_HI(net349));
 sg13g2_tiehi \proj__4.mux50/_0__297  (.L_HI(net350));
 sg13g2_tiehi \proj__4.mux52/_0__298  (.L_HI(net351));
 sg13g2_tiehi \proj__4.mux53/_0__299  (.L_HI(net352));
 sg13g2_tiehi \proj__4.mux53/_0__300  (.L_HI(net353));
 sg13g2_tiehi \proj__4.mux61/_0__301  (.L_HI(net354));
 sg13g2_tiehi \proj__4.mux62/_0__302  (.L_HI(net355));
 sg13g2_tiehi \proj__4.mux63/_0__303  (.L_HI(net356));
 sg13g2_tiehi \proj__4.mux63/_0__304  (.L_HI(net357));
 sg13g2_tiehi \proj__4.mux64/_0__305  (.L_HI(net358));
 sg13g2_tiehi \proj__4.mux65/_0__306  (.L_HI(net359));
 sg13g2_tiehi \proj__4.mux65/_0__307  (.L_HI(net360));
 sg13g2_tiehi \proj__4.mux66/_0__308  (.L_HI(net361));
 sg13g2_tiehi \proj__4.mux67/_0__309  (.L_HI(net362));
 sg13g2_tiehi \proj__4.mux67/_0__310  (.L_HI(net363));
 sg13g2_tiehi \proj__4.mux68/_0__311  (.L_HI(net364));
 sg13g2_tiehi \proj__4.mux76/_0__312  (.L_HI(net365));
 sg13g2_tiehi \proj__4.mux76/_0__313  (.L_HI(net366));
 sg13g2_tiehi \proj__4.mux77/_0__314  (.L_HI(net367));
 sg13g2_tiehi \proj__4.mux78/_0__315  (.L_HI(net368));
 sg13g2_tiehi \proj__4.mux78/_0__316  (.L_HI(net369));
 sg13g2_tiehi \proj__4.mux79/_0__317  (.L_HI(net370));
 sg13g2_tiehi \proj__4.mux79/_0__318  (.L_HI(net371));
 sg13g2_tiehi \proj__4.mux8/_0__319  (.L_HI(net372));
 sg13g2_tiehi \proj__4.mux80/_0__320  (.L_HI(net373));
 sg13g2_tiehi \proj__4.mux80/_0__321  (.L_HI(net374));
 sg13g2_tiehi \proj__4.mux81/_0__322  (.L_HI(net375));
 sg13g2_tiehi \proj__4.mux81/_0__323  (.L_HI(net376));
 sg13g2_tiehi \proj__4.mux82/_0__324  (.L_HI(net377));
 sg13g2_tiehi \proj__4.mux82/_0__325  (.L_HI(net378));
 sg13g2_tiehi \proj__4.mux83/_0__326  (.L_HI(net379));
 sg13g2_tiehi \proj__4.mux91/_0__327  (.L_HI(net380));
 sg13g2_tiehi \proj__4.mux92/_0__328  (.L_HI(net381));
 sg13g2_tiehi \proj__4.mux93/_0__329  (.L_HI(net382));
 sg13g2_tiehi \proj__4.mux94/_0__330  (.L_HI(net383));
 sg13g2_tiehi \proj__4.mux94/_0__331  (.L_HI(net384));
 sg13g2_tiehi \proj__4.mux96/_0__332  (.L_HI(net385));
 sg13g2_tiehi \proj__4.mux98/_0__333  (.L_HI(net386));
 sg13g2_tiehi \proj__4.mux98/_0__334  (.L_HI(net387));
 sg13g2_tiehi \proj__4.xor1/_0__335  (.L_HI(net388));
 sg13g2_tiehi \proj__2.flop1/_1__336  (.L_HI(net389));
 sg13g2_tielo \proj_10.flop11/_5__8  (.L_LO(net8));
 sg13g2_tielo \proj_10.flop12/_5__9  (.L_LO(net9));
 sg13g2_tielo \proj_10.flop13/_5__10  (.L_LO(net10));
 sg13g2_tielo \proj_10.flop14/_5__11  (.L_LO(net11));
 sg13g2_tielo \proj_10.mux11/_0__12  (.L_LO(net12));
 sg13g2_tielo \proj_10.mux12/_0__13  (.L_LO(net13));
 sg13g2_tielo \proj_10.mux13/_0__14  (.L_LO(net14));
 sg13g2_tielo \proj_10.mux14/_0__15  (.L_LO(net15));
 sg13g2_tielo \proj_10.mux15/_0__16  (.L_LO(net16));
 sg13g2_tielo \proj_10.mux16/_0__17  (.L_LO(net17));
 sg13g2_tielo \proj_10.mux17/_0__18  (.L_LO(net18));
 sg13g2_tielo \proj_10.mux18/_0__19  (.L_LO(net19));
 sg13g2_tielo \proj_10.mux19/_0__20  (.L_LO(net20));
 sg13g2_tielo \proj_10.mux20/_0__21  (.L_LO(net21));
 sg13g2_tielo \proj_10.mux21/_0__22  (.L_LO(net22));
 sg13g2_tielo \proj_10.mux21/_0__23  (.L_LO(net23));
 sg13g2_tielo \proj_10.mux22/_0__24  (.L_LO(net24));
 sg13g2_tielo \proj_10.mux23/_0__25  (.L_LO(net25));
 sg13g2_tielo \proj_10.mux25/_0__26  (.L_LO(net26));
 sg13g2_tielo \proj_10.mux26/_0__27  (.L_LO(net27));
 sg13g2_tielo \proj_10.mux27/_0__28  (.L_LO(net28));
 sg13g2_tielo \proj_10.mux29/_0__29  (.L_LO(net29));
 sg13g2_tielo \proj_10.mux30/_0__30  (.L_LO(net30));
 sg13g2_tielo \proj_10.mux31/_0__31  (.L_LO(net31));
 sg13g2_tielo \proj_10.mux32/_0__32  (.L_LO(net32));
 sg13g2_tielo \proj_10.mux33/_0__33  (.L_LO(net33));
 sg13g2_tielo \proj_10.mux34/_0__34  (.L_LO(net34));
 sg13g2_tielo \proj_10.mux35/_0__35  (.L_LO(net35));
 sg13g2_tielo \proj_10.mux36/_0__36  (.L_LO(net36));
 sg13g2_tielo \proj_10.not6/_0__37  (.L_LO(net37));
 sg13g2_tielo \proj_12.flop1/_4__38  (.L_LO(net38));
 sg13g2_tielo \proj_12.flop1/_5__39  (.L_LO(net39));
 sg13g2_tielo \proj_12.flop2/_4__40  (.L_LO(net40));
 sg13g2_tielo \proj_12.flop2/_5__41  (.L_LO(net41));
 sg13g2_tielo \proj__4.mux1/_0__42  (.L_LO(net42));
 sg13g2_tielo \proj__4.mux1/_0__43  (.L_LO(net43));
 sg13g2_tielo \proj__4.mux106/_0__44  (.L_LO(net44));
 sg13g2_tielo \proj__4.mux110/_0__45  (.L_LO(net45));
 sg13g2_tielo \proj__4.mux2/_0__46  (.L_LO(net46));
 sg13g2_tielo \proj__4.mux2/_0__47  (.L_LO(net47));
 sg13g2_tielo \proj__4.mux3/_0__48  (.L_LO(net48));
 sg13g2_tielo \proj__4.mux31/_0__49  (.L_LO(net49));
 sg13g2_tielo \proj__4.mux31/_0__50  (.L_LO(net50));
 sg13g2_tielo \proj__4.mux32/_0__51  (.L_LO(net51));
 sg13g2_tielo \proj__4.mux33/_0__52  (.L_LO(net52));
 sg13g2_tielo \proj__4.mux35/_0__53  (.L_LO(net53));
 sg13g2_tielo \proj__4.mux35/_0__54  (.L_LO(net54));
 sg13g2_tielo \proj__4.mux36/_0__55  (.L_LO(net55));
 sg13g2_tielo \proj__4.mux36/_0__56  (.L_LO(net56));
 sg13g2_tielo \proj__4.mux37/_0__57  (.L_LO(net57));
 sg13g2_tielo \proj__4.mux37/_0__58  (.L_LO(net58));
 sg13g2_tielo \proj__4.mux38/_0__59  (.L_LO(net59));
 sg13g2_tielo \proj__4.mux46/_0__60  (.L_LO(net60));
 sg13g2_tielo \proj__4.mux46/_0__61  (.L_LO(net61));
 sg13g2_tielo \proj__4.mux48/_0__62  (.L_LO(net62));
 sg13g2_tielo \proj__4.mux49/_0__63  (.L_LO(net63));
 sg13g2_tielo \proj__4.mux49/_0__64  (.L_LO(net64));
 sg13g2_tielo \proj__4.mux5/_0__65  (.L_LO(net65));
 sg13g2_tielo \proj__4.mux5/_0__66  (.L_LO(net66));
 sg13g2_tielo \proj__4.mux51/_0__67  (.L_LO(net67));
 sg13g2_tielo \proj__4.mux51/_0__68  (.L_LO(net68));
 sg13g2_tielo \proj__4.mux52/_0__69  (.L_LO(net69));
 sg13g2_tielo \proj__4.mux6/_0__70  (.L_LO(net70));
 sg13g2_tielo \proj__4.mux6/_0__71  (.L_LO(net71));
 sg13g2_tielo \proj__4.mux61/_0__72  (.L_LO(net72));
 sg13g2_tielo \proj__4.mux62/_0__73  (.L_LO(net73));
 sg13g2_tielo \proj__4.mux64/_0__74  (.L_LO(net74));
 sg13g2_tielo \proj__4.mux66/_0__75  (.L_LO(net75));
 sg13g2_tielo \proj__4.mux68/_0__76  (.L_LO(net76));
 sg13g2_tielo \proj__4.mux7/_0__77  (.L_LO(net77));
 sg13g2_tielo \proj__4.mux7/_0__78  (.L_LO(net78));
 sg13g2_tielo \proj__4.mux77/_0__79  (.L_LO(net79));
 sg13g2_tielo \proj__4.mux8/_0__80  (.L_LO(net80));
 sg13g2_tielo \proj__4.mux83/_0__81  (.L_LO(net81));
 sg13g2_tielo \proj__4.mux91/_0__82  (.L_LO(net82));
 sg13g2_tielo \proj__4.mux92/_0__83  (.L_LO(net83));
 sg13g2_tielo \proj__4.mux93/_0__84  (.L_LO(net84));
 sg13g2_tielo \proj__4.mux95/_0__85  (.L_LO(net85));
 sg13g2_tielo \proj__4.mux95/_0__86  (.L_LO(net86));
 sg13g2_tielo \proj__4.mux96/_0__87  (.L_LO(net87));
 sg13g2_tielo \proj__4.mux97/_0__88  (.L_LO(net88));
 sg13g2_tielo \proj__4.mux97/_0__89  (.L_LO(net89));
 sg13g2_tielo \proj__6.flop0/_5__90  (.L_LO(net90));
 sg13g2_tielo \proj__6.flop1/_5__91  (.L_LO(net91));
 sg13g2_tielo \proj__6.flop10/_5__92  (.L_LO(net92));
 sg13g2_tielo \proj__6.flop11/_5__93  (.L_LO(net93));
 sg13g2_tielo \proj__6.flop12/_5__94  (.L_LO(net94));
 sg13g2_tielo \proj__6.flop13/_5__95  (.L_LO(net95));
 sg13g2_tielo \proj__6.flop14/_5__96  (.L_LO(net96));
 sg13g2_tielo \proj__6.flop15/_5__97  (.L_LO(net97));
 sg13g2_tielo \proj__6.flop16/_5__98  (.L_LO(net98));
 sg13g2_tielo \proj__6.flop17/_5__99  (.L_LO(net99));
 sg13g2_tielo \proj__6.flop18/_5__100  (.L_LO(net100));
 sg13g2_tielo \proj__6.flop19/_5__101  (.L_LO(net101));
 sg13g2_tielo \proj__6.flop2/_5__102  (.L_LO(net102));
 sg13g2_tielo \proj__6.flop20/_5__103  (.L_LO(net103));
 sg13g2_tielo \proj__6.flop21/_5__104  (.L_LO(net104));
 sg13g2_tielo \proj__6.flop22/_5__105  (.L_LO(net105));
 sg13g2_tielo \proj__6.flop23/_5__106  (.L_LO(net106));
 sg13g2_tielo \proj__6.flop24/_5__107  (.L_LO(net107));
 sg13g2_tielo \proj__6.flop25/_5__108  (.L_LO(net108));
 sg13g2_tielo \proj__6.flop26/_5__109  (.L_LO(net109));
 sg13g2_tielo \proj__6.flop27/_5__110  (.L_LO(net110));
 sg13g2_tielo \proj__6.flop28/_5__111  (.L_LO(net111));
 sg13g2_tielo \proj__6.flop29/_5__112  (.L_LO(net112));
 sg13g2_tielo \proj__6.flop3/_5__113  (.L_LO(net113));
 sg13g2_tielo \proj__6.flop30/_5__114  (.L_LO(net114));
 sg13g2_tielo \proj__6.flop31/_5__115  (.L_LO(net115));
 sg13g2_tielo \proj__6.flop33/_5__116  (.L_LO(net116));
 sg13g2_tielo \proj__6.flop34/_5__117  (.L_LO(net117));
 sg13g2_tielo \proj__6.flop35/_5__118  (.L_LO(net118));
 sg13g2_tielo \proj__6.flop36/_5__119  (.L_LO(net119));
 sg13g2_tielo \proj__6.flop37/_5__120  (.L_LO(net120));
 sg13g2_tielo \proj__6.flop38/_5__121  (.L_LO(net121));
 sg13g2_tielo \proj__6.flop39/_5__122  (.L_LO(net122));
 sg13g2_tielo \proj__6.flop4/_5__123  (.L_LO(net123));
 sg13g2_tielo \proj__6.flop40/_5__124  (.L_LO(net124));
 sg13g2_tielo \proj__6.flop5/_5__125  (.L_LO(net125));
 sg13g2_tielo \proj__6.flop6/_5__126  (.L_LO(net126));
 sg13g2_tielo \proj__6.flop7/_5__127  (.L_LO(net127));
 sg13g2_tielo \proj__6.flop8/_5__128  (.L_LO(net128));
 sg13g2_tielo \proj__6.flop9/_5__129  (.L_LO(net129));
 sg13g2_tielo \proj__9.flop1/_5__130  (.L_LO(net130));
 sg13g2_tielo \proj__9.flop2/_5__131  (.L_LO(net131));
 sg13g2_tielo \proj__9.flop3/_5__132  (.L_LO(net132));
 sg13g2_tielo \proj__9.flop4/_5__133  (.L_LO(net133));
 sg13g2_tielo tt_um_wokwi_group_13_134 (.L_LO(net134));
 sg13g2_tielo tt_um_wokwi_group_13_135 (.L_LO(net135));
 sg13g2_tielo tt_um_wokwi_group_13_136 (.L_LO(net136));
 sg13g2_tielo tt_um_wokwi_group_13_137 (.L_LO(net137));
 sg13g2_tielo tt_um_wokwi_group_13_138 (.L_LO(net138));
 sg13g2_tielo tt_um_wokwi_group_13_139 (.L_LO(net139));
 sg13g2_tielo tt_um_wokwi_group_13_140 (.L_LO(net140));
 sg13g2_tielo tt_um_wokwi_group_13_141 (.L_LO(net141));
 sg13g2_tielo tt_um_wokwi_group_13_142 (.L_LO(net142));
 sg13g2_tielo tt_um_wokwi_group_13_143 (.L_LO(net143));
 sg13g2_tielo tt_um_wokwi_group_13_144 (.L_LO(net144));
 sg13g2_tielo tt_um_wokwi_group_13_145 (.L_LO(net145));
 sg13g2_tielo tt_um_wokwi_group_13_146 (.L_LO(net146));
 sg13g2_tielo tt_um_wokwi_group_13_147 (.L_LO(net147));
 sg13g2_tielo tt_um_wokwi_group_13_148 (.L_LO(net148));
 sg13g2_tielo tt_um_wokwi_group_13_149 (.L_LO(net149));
 sg13g2_tielo \proj_10.flop1/dffsr_150  (.L_LO(net150));
 sg13g2_and2_2 \proj_10.and1/_0_  (.A(net189),
    .B(net195),
    .X(\proj_10.net96 ));
 sg13g2_inv_1 \proj_10.flop1/_4_  (.Y(\proj_10.flop1/_0_ ),
    .A(\proj_10.net43 ));
 sg13g2_inv_1 \proj_10.flop1/_5_  (.Y(\proj_10.flop1/_1_ ),
    .A(\proj_10.net42 ));
 sg13g2_tielo \proj_10.flop1/dffsr_151  (.L_LO(net151));
 sg13g2_tielo \proj_10.flop10/dffsr_152  (.L_LO(net152));
 sg13g2_sdfbbp_1 \proj_10.flop1/dffsr  (.Q(\proj_10.net28 ),
    .Q_N(\proj_10.flop1/notq ),
    .RESET_B(\proj_10.flop1/_0_ ),
    .SET_B(\proj_10.flop1/_1_ ),
    .D(\proj_10.net41 ),
    .SCE(net151),
    .SCD(net150),
    .CLK(clknet_2_2__leaf_clk_regs));
 sg13g2_inv_1 \proj_10.flop10/_4_  (.Y(\proj_10.flop10/_0_ ),
    .A(net183));
 sg13g2_inv_1 \proj_10.flop10/_5_  (.Y(\proj_10.flop10/_1_ ),
    .A(net7));
 sg13g2_tielo \proj_10.flop10/dffsr_153  (.L_LO(net153));
 sg13g2_tielo \proj_10.flop11/dffsr_154  (.L_LO(net154));
 sg13g2_sdfbbp_1 \proj_10.flop10/dffsr  (.Q(\proj_10.net83 ),
    .Q_N(\proj_10.flop10/notq ),
    .RESET_B(\proj_10.flop10/_0_ ),
    .SET_B(\proj_10.flop10/_1_ ),
    .D(net403),
    .SCE(net153),
    .SCD(net152),
    .CLK(clknet_2_1__leaf_clk_regs));
 sg13g2_inv_1 \proj_10.flop11/_4_  (.Y(\proj_10.flop11/_0_ ),
    .A(net183));
 sg13g2_inv_1 \proj_10.flop11/_5_  (.Y(\proj_10.flop11/_1_ ),
    .A(net8));
 sg13g2_tielo \proj_10.flop11/dffsr_155  (.L_LO(net155));
 sg13g2_tielo \proj_10.flop12/dffsr_156  (.L_LO(net156));
 sg13g2_sdfbbp_1 \proj_10.flop11/dffsr  (.Q(\proj_10.net85 ),
    .Q_N(\proj_10.flop11/notq ),
    .RESET_B(\proj_10.flop11/_0_ ),
    .SET_B(\proj_10.flop11/_1_ ),
    .D(net408),
    .SCE(net155),
    .SCD(net154),
    .CLK(clknet_2_3__leaf_clk_regs));
 sg13g2_inv_1 \proj_10.flop12/_4_  (.Y(\proj_10.flop12/_0_ ),
    .A(net183));
 sg13g2_inv_1 \proj_10.flop12/_5_  (.Y(\proj_10.flop12/_1_ ),
    .A(net9));
 sg13g2_tielo \proj_10.flop12/dffsr_157  (.L_LO(net157));
 sg13g2_tielo \proj_10.flop13/dffsr_158  (.L_LO(net158));
 sg13g2_sdfbbp_1 \proj_10.flop12/dffsr  (.Q(\proj_10.net87 ),
    .Q_N(\proj_10.flop12/notq ),
    .RESET_B(\proj_10.flop12/_0_ ),
    .SET_B(\proj_10.flop12/_1_ ),
    .D(net406),
    .SCE(net157),
    .SCD(net156),
    .CLK(clknet_2_3__leaf_clk_regs));
 sg13g2_inv_1 \proj_10.flop13/_4_  (.Y(\proj_10.flop13/_0_ ),
    .A(net183));
 sg13g2_inv_1 \proj_10.flop13/_5_  (.Y(\proj_10.flop13/_1_ ),
    .A(net10));
 sg13g2_tielo \proj_10.flop13/dffsr_159  (.L_LO(net159));
 sg13g2_tielo \proj_10.flop14/dffsr_160  (.L_LO(net213));
 sg13g2_sdfbbp_1 \proj_10.flop13/dffsr  (.Q(\proj_10.net89 ),
    .Q_N(\proj_10.flop13/notq ),
    .RESET_B(\proj_10.flop13/_0_ ),
    .SET_B(\proj_10.flop13/_1_ ),
    .D(net413),
    .SCE(net159),
    .SCD(net158),
    .CLK(clknet_2_3__leaf_clk_regs));
 sg13g2_inv_1 \proj_10.flop14/_4_  (.Y(\proj_10.flop14/_0_ ),
    .A(net183));
 sg13g2_inv_1 \proj_10.flop14/_5_  (.Y(\proj_10.flop14/_1_ ),
    .A(net11));
 sg13g2_tielo \proj_10.flop14/dffsr_161  (.L_LO(net214));
 sg13g2_tielo \proj_10.flop2/dffsr_162  (.L_LO(net215));
 sg13g2_sdfbbp_1 \proj_10.flop14/dffsr  (.Q(\proj_10.net71 ),
    .Q_N(\proj_10.flop14/notq ),
    .RESET_B(\proj_10.flop14/_0_ ),
    .SET_B(\proj_10.flop14/_1_ ),
    .D(net412),
    .SCE(net214),
    .SCD(net213),
    .CLK(clknet_2_3__leaf_clk_regs));
 sg13g2_inv_1 \proj_10.flop2/_4_  (.Y(\proj_10.flop2/_0_ ),
    .A(\proj_10.net45 ));
 sg13g2_inv_1 \proj_10.flop2/_5_  (.Y(\proj_10.flop2/_1_ ),
    .A(\proj_10.net44 ));
 sg13g2_tielo \proj_10.flop2/dffsr_163  (.L_LO(net216));
 sg13g2_tielo \proj_10.flop3/dffsr_164  (.L_LO(net217));
 sg13g2_sdfbbp_1 \proj_10.flop2/dffsr  (.Q(\proj_10.net33 ),
    .Q_N(\proj_10.flop2/notq ),
    .RESET_B(\proj_10.flop2/_0_ ),
    .SET_B(\proj_10.flop2/_1_ ),
    .D(net411),
    .SCE(net216),
    .SCD(net215),
    .CLK(clknet_2_2__leaf_clk_regs));
 sg13g2_inv_1 \proj_10.flop3/_4_  (.Y(\proj_10.flop3/_0_ ),
    .A(\proj_10.net47 ));
 sg13g2_inv_1 \proj_10.flop3/_5_  (.Y(\proj_10.flop3/_1_ ),
    .A(\proj_10.net46 ));
 sg13g2_tielo \proj_10.flop3/dffsr_165  (.L_LO(net218));
 sg13g2_tielo \proj_10.flop4/dffsr_166  (.L_LO(net219));
 sg13g2_sdfbbp_1 \proj_10.flop3/dffsr  (.Q(\proj_10.net48 ),
    .Q_N(\proj_10.flop3/notq ),
    .RESET_B(\proj_10.flop3/_0_ ),
    .SET_B(\proj_10.flop3/_1_ ),
    .D(net417),
    .SCE(net218),
    .SCD(net217),
    .CLK(clknet_2_2__leaf_clk_regs));
 sg13g2_inv_1 \proj_10.flop4/_4_  (.Y(\proj_10.flop4/_0_ ),
    .A(\proj_10.net50 ));
 sg13g2_inv_1 \proj_10.flop4/_5_  (.Y(\proj_10.flop4/_1_ ),
    .A(\proj_10.net49 ));
 sg13g2_tielo \proj_10.flop4/dffsr_167  (.L_LO(net220));
 sg13g2_tielo \proj_10.flop5/dffsr_168  (.L_LO(net221));
 sg13g2_sdfbbp_1 \proj_10.flop4/dffsr  (.Q(\proj_10.net51 ),
    .Q_N(\proj_10.flop4/notq ),
    .RESET_B(\proj_10.flop4/_0_ ),
    .SET_B(\proj_10.flop4/_1_ ),
    .D(net414),
    .SCE(net220),
    .SCD(net219),
    .CLK(clknet_2_2__leaf_clk_regs));
 sg13g2_inv_1 \proj_10.flop5/_4_  (.Y(\proj_10.flop5/_0_ ),
    .A(\proj_10.net53 ));
 sg13g2_inv_1 \proj_10.flop5/_5_  (.Y(\proj_10.flop5/_1_ ),
    .A(\proj_10.net52 ));
 sg13g2_tielo \proj_10.flop5/dffsr_169  (.L_LO(net222));
 sg13g2_tielo \proj_10.flop6/dffsr_170  (.L_LO(net223));
 sg13g2_sdfbbp_1 \proj_10.flop5/dffsr  (.Q(\proj_10.net54 ),
    .Q_N(\proj_10.flop5/notq ),
    .RESET_B(\proj_10.flop5/_0_ ),
    .SET_B(\proj_10.flop5/_1_ ),
    .D(net415),
    .SCE(net222),
    .SCD(net221),
    .CLK(clknet_2_2__leaf_clk_regs));
 sg13g2_inv_1 \proj_10.flop6/_4_  (.Y(\proj_10.flop6/_0_ ),
    .A(\proj_10.net56 ));
 sg13g2_inv_1 \proj_10.flop6/_5_  (.Y(\proj_10.flop6/_1_ ),
    .A(\proj_10.net55 ));
 sg13g2_tielo \proj_10.flop6/dffsr_171  (.L_LO(net224));
 sg13g2_tielo \proj_10.flop7/dffsr_172  (.L_LO(net225));
 sg13g2_sdfbbp_1 \proj_10.flop6/dffsr  (.Q(\proj_10.net57 ),
    .Q_N(\proj_10.flop6/notq ),
    .RESET_B(\proj_10.flop6/_0_ ),
    .SET_B(\proj_10.flop6/_1_ ),
    .D(net402),
    .SCE(net224),
    .SCD(net223),
    .CLK(clknet_2_2__leaf_clk_regs));
 sg13g2_inv_1 \proj_10.flop7/_4_  (.Y(\proj_10.flop7/_0_ ),
    .A(\proj_10.net73 ));
 sg13g2_inv_1 \proj_10.flop7/_5_  (.Y(\proj_10.flop7/_1_ ),
    .A(\proj_10.net72 ));
 sg13g2_tielo \proj_10.flop7/dffsr_173  (.L_LO(net226));
 sg13g2_tielo \proj_10.flop8/dffsr_174  (.L_LO(net227));
 sg13g2_sdfbbp_1 \proj_10.flop7/dffsr  (.Q(\proj_10.net74 ),
    .Q_N(\proj_10.flop7/notq ),
    .RESET_B(\proj_10.flop7/_0_ ),
    .SET_B(\proj_10.flop7/_1_ ),
    .D(net409),
    .SCE(net226),
    .SCD(net225),
    .CLK(clknet_2_3__leaf_clk_regs));
 sg13g2_inv_1 \proj_10.flop8/_4_  (.Y(\proj_10.flop8/_0_ ),
    .A(\proj_10.net76 ));
 sg13g2_inv_1 \proj_10.flop8/_5_  (.Y(\proj_10.flop8/_1_ ),
    .A(\proj_10.net75 ));
 sg13g2_tielo \proj_10.flop8/dffsr_175  (.L_LO(net228));
 sg13g2_tielo \proj_10.flop9/dffsr_176  (.L_LO(net229));
 sg13g2_sdfbbp_1 \proj_10.flop8/dffsr  (.Q(\proj_10.net77 ),
    .Q_N(\proj_10.flop8/notq ),
    .RESET_B(\proj_10.flop8/_0_ ),
    .SET_B(\proj_10.flop8/_1_ ),
    .D(net410),
    .SCE(net228),
    .SCD(net227),
    .CLK(clknet_2_3__leaf_clk_regs));
 sg13g2_inv_1 \proj_10.flop9/_4_  (.Y(\proj_10.flop9/_0_ ),
    .A(\proj_10.net79 ));
 sg13g2_inv_1 \proj_10.flop9/_5_  (.Y(\proj_10.flop9/_1_ ),
    .A(\proj_10.net78 ));
 sg13g2_tielo \proj_10.flop9/dffsr_177  (.L_LO(net230));
 sg13g2_tielo \proj_12.flop1/dffsr_178  (.L_LO(net231));
 sg13g2_sdfbbp_1 \proj_10.flop9/dffsr  (.Q(\proj_10.net80 ),
    .Q_N(\proj_10.flop9/notq ),
    .RESET_B(\proj_10.flop9/_0_ ),
    .SET_B(\proj_10.flop9/_1_ ),
    .D(net416),
    .SCE(net230),
    .SCD(net229),
    .CLK(clknet_2_1__leaf_clk_regs));
 sg13g2_mux2_1 \proj_10.mux1/_0_  (.A0(\proj_10.net24 ),
    .A1(\proj_10.net25 ),
    .S(net187),
    .X(\proj_10.net12 ));
 sg13g2_mux2_1 \proj_10.mux10/_0_  (.A0(\proj_10.net38 ),
    .A1(\proj_10.net37 ),
    .S(\proj_10.net30 ),
    .X(\proj_10.net40 ));
 sg13g2_mux2_1 \proj_10.mux11/_0_  (.A0(net12),
    .A1(net205),
    .S(net181),
    .X(\proj_10.net42 ));
 sg13g2_mux2_1 \proj_10.mux12/_0_  (.A0(net13),
    .A1(\proj_10.net60 ),
    .S(net181),
    .X(\proj_10.net43 ));
 sg13g2_mux2_1 \proj_10.mux13/_0_  (.A0(net14),
    .A1(net202),
    .S(net182),
    .X(\proj_10.net44 ));
 sg13g2_mux2_1 \proj_10.mux14/_0_  (.A0(net15),
    .A1(\proj_10.net61 ),
    .S(net182),
    .X(\proj_10.net45 ));
 sg13g2_mux2_1 \proj_10.mux15/_0_  (.A0(net16),
    .A1(net198),
    .S(net181),
    .X(\proj_10.net46 ));
 sg13g2_mux2_1 \proj_10.mux16/_0_  (.A0(net17),
    .A1(\proj_10.net62 ),
    .S(net181),
    .X(\proj_10.net47 ));
 sg13g2_mux2_1 \proj_10.mux17/_0_  (.A0(net18),
    .A1(net194),
    .S(net181),
    .X(\proj_10.net49 ));
 sg13g2_mux2_1 \proj_10.mux18/_0_  (.A0(net19),
    .A1(\proj_10.net63 ),
    .S(net181),
    .X(\proj_10.net50 ));
 sg13g2_mux2_1 \proj_10.mux19/_0_  (.A0(net20),
    .A1(net193),
    .S(net181),
    .X(\proj_10.net52 ));
 sg13g2_mux2_1 \proj_10.mux2/_0_  (.A0(\proj_10.net25 ),
    .A1(\proj_10.net24 ),
    .S(net187),
    .X(\proj_10.net16 ));
 sg13g2_mux2_1 \proj_10.mux20/_0_  (.A0(net21),
    .A1(\proj_10.net64 ),
    .S(net181),
    .X(\proj_10.net53 ));
 sg13g2_mux2_1 \proj_10.mux21/_0_  (.A0(net22),
    .A1(net23),
    .S(net182),
    .X(\proj_10.net55 ));
 sg13g2_mux2_1 \proj_10.mux22/_0_  (.A0(net24),
    .A1(\proj_10.net66 ),
    .S(net182),
    .X(\proj_10.net56 ));
 sg13g2_mux2_1 \proj_10.mux23/_0_  (.A0(net25),
    .A1(clknet_1_0__leaf_clk),
    .S(net185),
    .X(\proj_10.net18 ));
 sg13g2_mux2_1 \proj_10.mux24/_0_  (.A0(net418),
    .A1(net415),
    .S(net188),
    .X(\proj_10.net41 ));
 sg13g2_mux2_1 \proj_10.mux25/_0_  (.A0(\proj_10.net48 ),
    .A1(net26),
    .S(net188),
    .X(\proj_10.net34 ));
 sg13g2_mux2_1 \proj_10.mux26/_0_  (.A0(\proj_10.net51 ),
    .A1(net27),
    .S(net188),
    .X(\proj_10.net29 ));
 sg13g2_mux2_1 \proj_10.mux27/_0_  (.A0(\proj_10.net54 ),
    .A1(net28),
    .S(net188),
    .X(\proj_10.net37 ));
 sg13g2_mux2_1 \proj_10.mux28/_0_  (.A0(\proj_10.net57 ),
    .A1(\proj_10.net51 ),
    .S(net188),
    .X(\proj_10.net38 ));
 sg13g2_mux2_1 \proj_10.mux29/_0_  (.A0(net29),
    .A1(\proj_10.net48 ),
    .S(net188),
    .X(\proj_10.net69 ));
 sg13g2_mux2_1 \proj_10.mux3/_0_  (.A0(\proj_10.net26 ),
    .A1(\proj_10.net27 ),
    .S(net2),
    .X(\proj_10.net13 ));
 sg13g2_mux2_2 \proj_10.mux30/_0_  (.A0(net30),
    .A1(net193),
    .S(net188),
    .X(\proj_10.net30 ));
 sg13g2_mux2_1 \proj_10.mux31/_0_  (.A0(net31),
    .A1(net205),
    .S(\proj_10.net82 ),
    .X(\proj_10.net72 ));
 sg13g2_mux2_1 \proj_10.mux32/_0_  (.A0(net32),
    .A1(\proj_10.net92 ),
    .S(\proj_10.net82 ),
    .X(\proj_10.net73 ));
 sg13g2_mux2_1 \proj_10.mux33/_0_  (.A0(net33),
    .A1(net202),
    .S(net183),
    .X(\proj_10.net75 ));
 sg13g2_mux2_1 \proj_10.mux34/_0_  (.A0(net34),
    .A1(\proj_10.net93 ),
    .S(\proj_10.net82 ),
    .X(\proj_10.net76 ));
 sg13g2_mux2_1 \proj_10.mux35/_0_  (.A0(net35),
    .A1(net198),
    .S(net183),
    .X(\proj_10.net78 ));
 sg13g2_mux2_1 \proj_10.mux36/_0_  (.A0(net36),
    .A1(\proj_10.net94 ),
    .S(net183),
    .X(\proj_10.net79 ));
 sg13g2_mux2_1 \proj_10.mux37/_0_  (.A0(\proj_10.net31 ),
    .A1(\proj_10.net74 ),
    .S(\proj_10.net96 ),
    .X(\proj_10.net11 ));
 sg13g2_mux2_1 \proj_10.mux38/_0_  (.A0(\proj_10.net35 ),
    .A1(\proj_10.net77 ),
    .S(\proj_10.net96 ),
    .X(\proj_10.net24 ));
 sg13g2_mux2_1 \proj_10.mux39/_0_  (.A0(\proj_10.net36 ),
    .A1(\proj_10.net87 ),
    .S(\proj_10.net96 ),
    .X(\proj_10.net26 ));
 sg13g2_mux2_1 \proj_10.mux4/_0_  (.A0(\proj_10.net27 ),
    .A1(\proj_10.net26 ),
    .S(net2),
    .X(\proj_10.net15 ));
 sg13g2_mux2_1 \proj_10.mux40/_0_  (.A0(\proj_10.net32 ),
    .A1(\proj_10.net85 ),
    .S(\proj_10.net96 ),
    .X(\proj_10.net14 ));
 sg13g2_mux2_1 \proj_10.mux41/_0_  (.A0(\proj_10.net39 ),
    .A1(\proj_10.net83 ),
    .S(\proj_10.net96 ),
    .X(\proj_10.net27 ));
 sg13g2_mux2_1 \proj_10.mux42/_0_  (.A0(\proj_10.net40 ),
    .A1(\proj_10.net71 ),
    .S(\proj_10.net96 ),
    .X(\proj_10.net25 ));
 sg13g2_mux2_1 \proj_10.mux43/_0_  (.A0(\proj_10.net69 ),
    .A1(\proj_10.net95 ),
    .S(\proj_10.net96 ),
    .X(\proj_10.net17 ));
 sg13g2_mux2_1 \proj_10.mux5/_0_  (.A0(\proj_10.net28 ),
    .A1(\proj_10.net29 ),
    .S(\proj_10.net30 ),
    .X(\proj_10.net31 ));
 sg13g2_mux2_1 \proj_10.mux6/_0_  (.A0(\proj_10.net29 ),
    .A1(\proj_10.net28 ),
    .S(\proj_10.net30 ),
    .X(\proj_10.net32 ));
 sg13g2_mux2_1 \proj_10.mux7/_0_  (.A0(\proj_10.net33 ),
    .A1(\proj_10.net34 ),
    .S(\proj_10.net30 ),
    .X(\proj_10.net35 ));
 sg13g2_mux2_1 \proj_10.mux8/_0_  (.A0(\proj_10.net34 ),
    .A1(\proj_10.net33 ),
    .S(\proj_10.net30 ),
    .X(\proj_10.net36 ));
 sg13g2_mux2_1 \proj_10.mux9/_0_  (.A0(\proj_10.net37 ),
    .A1(\proj_10.net38 ),
    .S(\proj_10.net30 ),
    .X(\proj_10.net39 ));
 sg13g2_inv_1 \proj_10.not1/_0_  (.Y(\proj_10.net60 ),
    .A(net205));
 sg13g2_inv_1 \proj_10.not10/_0_  (.Y(\proj_10.net94 ),
    .A(net198));
 sg13g2_inv_2 \proj_10.not16/_0_  (.Y(\proj_10.net82 ),
    .A(net212));
 sg13g2_inv_1 \proj_10.not2/_0_  (.Y(\proj_10.net61 ),
    .A(net202));
 sg13g2_inv_1 \proj_10.not3/_0_  (.Y(\proj_10.net62 ),
    .A(net198));
 sg13g2_inv_1 \proj_10.not4/_0_  (.Y(\proj_10.net63 ),
    .A(net195));
 sg13g2_inv_1 \proj_10.not5/_0_  (.Y(\proj_10.net64 ),
    .A(net193));
 sg13g2_inv_1 \proj_10.not6/_0_  (.Y(\proj_10.net66 ),
    .A(net37));
 sg13g2_inv_1 \proj_10.not7/_0_  (.Y(\proj_10.net59 ),
    .A(net210));
 sg13g2_inv_1 \proj_10.not8/_0_  (.Y(\proj_10.net92 ),
    .A(net205));
 sg13g2_inv_1 \proj_10.not9/_0_  (.Y(\proj_10.net93 ),
    .A(net202));
 sg13g2_or2_1 \proj_10.or1/_0_  (.X(\proj_10.net95 ),
    .B(\proj_10.net80 ),
    .A(\proj_10.net89 ));
 sg13g2_inv_1 \proj_11.not1/_0_  (.Y(\proj_11.net9 ),
    .A(net204));
 sg13g2_inv_1 \proj_11.not2/_0_  (.Y(\proj_11.net10 ),
    .A(net199));
 sg13g2_inv_1 \proj_11.not3/_0_  (.Y(\proj_11.net11 ),
    .A(net197));
 sg13g2_inv_1 \proj_11.not4/_0_  (.Y(\proj_11.net12 ),
    .A(net195));
 sg13g2_inv_1 \proj_12.flop1/_4_  (.Y(\proj_12.flop1/_0_ ),
    .A(net38));
 sg13g2_inv_1 \proj_12.flop1/_5_  (.Y(\proj_12.flop1/_1_ ),
    .A(net39));
 sg13g2_tielo \proj_12.flop1/dffsr_179  (.L_LO(net232));
 sg13g2_tielo \proj_12.flop2/dffsr_180  (.L_LO(net233));
 sg13g2_sdfbbp_1 \proj_12.flop1/dffsr  (.Q(\proj_12.net19 ),
    .Q_N(\proj_12.net17 ),
    .RESET_B(\proj_12.flop1/_0_ ),
    .SET_B(\proj_12.flop1/_1_ ),
    .D(net401),
    .SCE(net232),
    .SCD(net231),
    .CLK(clknet_2_0__leaf_clk_regs));
 sg13g2_inv_1 \proj_12.flop2/_4_  (.Y(\proj_12.flop2/_0_ ),
    .A(net40));
 sg13g2_inv_1 \proj_12.flop2/_5_  (.Y(\proj_12.flop2/_1_ ),
    .A(net41));
 sg13g2_tielo \proj_12.flop2/dffsr_181  (.L_LO(net234));
 sg13g2_tielo \proj__6.flop0/dffsr_182  (.L_LO(net235));
 sg13g2_sdfbbp_1 \proj_12.flop2/dffsr  (.Q(\proj_12.net11 ),
    .Q_N(\proj_12.net20 ),
    .RESET_B(\proj_12.flop2/_0_ ),
    .SET_B(\proj_12.flop2/_1_ ),
    .D(\proj_12.net20 ),
    .SCE(net234),
    .SCD(net233),
    .CLK(\proj_12.net19 ));
 sg13g2_inv_1 \proj_12.not1/_0_  (.Y(\proj_12.net7 ),
    .A(net204));
 sg13g2_inv_1 \proj_12.not2/_0_  (.Y(\proj_12.net8 ),
    .A(net199));
 sg13g2_inv_1 \proj_12.not3/_0_  (.Y(\proj_12.net9 ),
    .A(net197));
 sg13g2_inv_1 \proj_12.not4/_0_  (.Y(\proj_12.net10 ),
    .A(net195));
 sg13g2_or2_1 \proj_13.or1/_0_  (.X(\proj_13.net22 ),
    .B(net187),
    .A(net184));
 sg13g2_or2_1 \proj_13.or10/_0_  (.X(\proj_13.net30 ),
    .B(net203),
    .A(net196));
 sg13g2_or2_1 \proj_13.or11/_0_  (.X(\proj_13.net31 ),
    .B(\proj_13.net30 ),
    .A(net191));
 sg13g2_or2_1 \proj_13.or12/_0_  (.X(\proj_13.net32 ),
    .B(\proj_13.net31 ),
    .A(net194));
 sg13g2_or2_1 \proj_13.or13/_0_  (.X(\proj_13.net33 ),
    .B(\proj_13.net32 ),
    .A(net190));
 sg13g2_or2_1 \proj_13.or14/_0_  (.X(\proj_13.net34 ),
    .B(\proj_13.net33 ),
    .A(net187));
 sg13g2_or2_1 \proj_13.or15/_0_  (.X(\proj_13.net12 ),
    .B(\proj_13.net34 ),
    .A(net184));
 sg13g2_or2_1 \proj_13.or16/_0_  (.X(\proj_13.net35 ),
    .B(net199),
    .A(net196));
 sg13g2_or2_1 \proj_13.or17/_0_  (.X(\proj_13.net27 ),
    .B(\proj_13.net26 ),
    .A(net203));
 sg13g2_or2_1 \proj_13.or18/_0_  (.X(\proj_13.net36 ),
    .B(net192),
    .A(\proj_13.net35 ));
 sg13g2_or2_1 \proj_13.or19/_0_  (.X(\proj_13.net37 ),
    .B(net190),
    .A(\proj_13.net36 ));
 sg13g2_or2_1 \proj_13.or2/_0_  (.X(\proj_13.net23 ),
    .B(net190),
    .A(\proj_13.net22 ));
 sg13g2_or2_1 \proj_13.or20/_0_  (.X(\proj_13.net13 ),
    .B(net186),
    .A(\proj_13.net37 ));
 sg13g2_or2_1 \proj_13.or21/_0_  (.X(\proj_13.net38 ),
    .B(net201),
    .A(net190));
 sg13g2_or2_1 \proj_13.or22/_0_  (.X(\proj_13.net14 ),
    .B(net184),
    .A(\proj_13.net38 ));
 sg13g2_or2_1 \proj_13.or23/_0_  (.X(\proj_13.net39 ),
    .B(net189),
    .A(net193));
 sg13g2_or2_1 \proj_13.or24/_0_  (.X(\proj_13.net40 ),
    .B(net195),
    .A(\proj_13.net39 ));
 sg13g2_or2_1 \proj_13.or25/_0_  (.X(\proj_13.net15 ),
    .B(net186),
    .A(\proj_13.net40 ));
 sg13g2_or2_1 \proj_13.or26/_0_  (.X(\proj_13.net41 ),
    .B(net196),
    .A(net201));
 sg13g2_or2_1 \proj_13.or27/_0_  (.X(\proj_13.net42 ),
    .B(net195),
    .A(\proj_13.net41 ));
 sg13g2_or2_1 \proj_13.or28/_0_  (.X(\proj_13.net43 ),
    .B(net193),
    .A(\proj_13.net42 ));
 sg13g2_or2_1 \proj_13.or29/_0_  (.X(\proj_13.net44 ),
    .B(net188),
    .A(\proj_13.net43 ));
 sg13g2_or2_1 \proj_13.or3/_0_  (.X(\proj_13.net24 ),
    .B(net192),
    .A(\proj_13.net23 ));
 sg13g2_or2_1 \proj_13.or30/_0_  (.X(\proj_13.net16 ),
    .B(net186),
    .A(\proj_13.net44 ));
 sg13g2_or2_1 \proj_13.or4/_0_  (.X(\proj_13.net25 ),
    .B(net197),
    .A(\proj_13.net24 ));
 sg13g2_or2_1 \proj_13.or5/_0_  (.X(\proj_13.net10 ),
    .B(net199),
    .A(\proj_13.net25 ));
 sg13g2_or2_1 \proj_13.or6/_0_  (.X(\proj_13.net26 ),
    .B(net201),
    .A(net196));
 sg13g2_or2_1 \proj_13.or7/_0_  (.X(\proj_13.net28 ),
    .B(\proj_13.net27 ),
    .A(net194));
 sg13g2_or2_1 \proj_13.or8/_0_  (.X(\proj_13.net29 ),
    .B(\proj_13.net28 ),
    .A(net187));
 sg13g2_or2_1 \proj_13.or9/_0_  (.X(\proj_13.net11 ),
    .B(\proj_13.net29 ),
    .A(net184));
 sg13g2_and2_1 \proj_14.and1/_0_  (.A(net187),
    .B(clknet_1_1__leaf_clk),
    .X(\proj_14.net3 ));
 sg13g2_inv_1 \proj_15.not2/_0_  (.Y(\proj_15.net10 ),
    .A(net199));
 sg13g2_inv_1 \proj_15.not3/_0_  (.Y(\proj_15.net11 ),
    .A(net197));
 sg13g2_inv_1 \proj_15.not4/_0_  (.Y(\proj_15.net12 ),
    .A(net1));
 sg13g2_xor2_1 \proj_15.xor1/_0_  (.B(net204),
    .A(net199),
    .X(\proj_15.net9 ));
 sg13g2_inv_1 \proj__0.not1/_0_  (.Y(\proj__0.net10 ),
    .A(net204));
 sg13g2_or2_1 \proj__0.or1/_0_  (.X(\proj__0.net11 ),
    .B(net197),
    .A(net1));
 sg13g2_nand2_1 \proj__1.nand1/_0_  (.Y(\proj__1.net10 ),
    .A(net199),
    .B(net204));
 sg13g2_inv_1 \proj__1.not1/_0_  (.Y(\proj__1.net12 ),
    .A(net192));
 sg13g2_or2_1 \proj__1.or1/_0_  (.X(\proj__1.net11 ),
    .B(net197),
    .A(net195));
 sg13g2_xor2_1 \proj__1.xor1/_0_  (.B(clknet_1_0__leaf_clk),
    .A(net190),
    .X(\proj__1.net13 ));
 sg13g2_dfrbp_1 \proj__2.flop1/_1_  (.CLK(clknet_2_0__leaf_clk_regs),
    .RESET_B(net389),
    .D(net398),
    .Q_N(\proj__2.net12 ),
    .Q(\proj__2.net13 ));
 sg13g2_tiehi \proj__2.flop2/_1__337  (.L_HI(net390));
 sg13g2_dfrbp_1 \proj__2.flop2/_1_  (.CLK(\proj__2.net13 ),
    .RESET_B(net390),
    .D(\proj__2.net14 ),
    .Q_N(\proj__2.net14 ),
    .Q(\proj__2.net6 ));
 sg13g2_tiehi \proj__3.flop1/_1__338  (.L_HI(net391));
 sg13g2_and2_1 \proj__3.and10/_0_  (.A(\proj__3.net14 ),
    .B(\proj__3.net24 ),
    .X(\proj__3.net6 ));
 sg13g2_and2_1 \proj__3.and11/_0_  (.A(\proj__3.net17 ),
    .B(\proj__3.net18 ),
    .X(\proj__3.net25 ));
 sg13g2_and2_1 \proj__3.and12/_0_  (.A(\proj__3.net15 ),
    .B(\proj__3.net25 ),
    .X(\proj__3.net5 ));
 sg13g2_and2_1 \proj__3.and13/_0_  (.A(\proj__3.net17 ),
    .B(\proj__3.net18 ),
    .X(\proj__3.net26 ));
 sg13g2_and2_1 \proj__3.and14/_0_  (.A(\proj__3.net14 ),
    .B(\proj__3.net26 ),
    .X(\proj__3.net4 ));
 sg13g2_and2_1 \proj__3.and15/_0_  (.A(\proj__3.net16 ),
    .B(\proj__3.net18 ),
    .X(\proj__3.net27 ));
 sg13g2_and2_1 \proj__3.and16/_0_  (.A(\proj__3.net15 ),
    .B(\proj__3.net27 ),
    .X(\proj__3.net28 ));
 sg13g2_and2_1 \proj__3.and17/_0_  (.A(\proj__3.net16 ),
    .B(\proj__3.net18 ),
    .X(\proj__3.net29 ));
 sg13g2_and2_1 \proj__3.and18/_0_  (.A(\proj__3.net14 ),
    .B(\proj__3.net29 ),
    .X(\proj__3.net7 ));
 sg13g2_and2_1 \proj__3.and3/_0_  (.A(\proj__3.net17 ),
    .B(\proj__3.net15 ),
    .X(\proj__3.net20 ));
 sg13g2_and2_1 \proj__3.and4/_0_  (.A(\proj__3.net19 ),
    .B(\proj__3.net20 ),
    .X(\proj__3.net2 ));
 sg13g2_and2_1 \proj__3.and5/_0_  (.A(\proj__3.net17 ),
    .B(\proj__3.net19 ),
    .X(\proj__3.net21 ));
 sg13g2_and2_1 \proj__3.and6/_0_  (.A(\proj__3.net14 ),
    .B(\proj__3.net21 ),
    .X(\proj__3.net3 ));
 sg13g2_and2_1 \proj__3.and7/_0_  (.A(\proj__3.net16 ),
    .B(\proj__3.net19 ),
    .X(\proj__3.net22 ));
 sg13g2_and2_1 \proj__3.and8/_0_  (.A(\proj__3.net15 ),
    .B(\proj__3.net22 ),
    .X(\proj__3.net23 ));
 sg13g2_and2_1 \proj__3.and9/_0_  (.A(\proj__3.net16 ),
    .B(\proj__3.net19 ),
    .X(\proj__3.net24 ));
 sg13g2_dfrbp_1 \proj__3.flop1/_1_  (.CLK(clknet_2_0__leaf_clk_regs),
    .RESET_B(net391),
    .D(net399),
    .Q_N(\proj__3.net14 ),
    .Q(\proj__3.net15 ));
 sg13g2_tiehi \proj__3.flop2/_1__339  (.L_HI(net392));
 sg13g2_dfrbp_1 \proj__3.flop2/_1_  (.CLK(\proj__3.net15 ),
    .RESET_B(net392),
    .D(\proj__3.net16 ),
    .Q_N(\proj__3.net16 ),
    .Q(\proj__3.net17 ));
 sg13g2_tiehi \proj__3.flop3/_1__340  (.L_HI(net393));
 sg13g2_dfrbp_1 \proj__3.flop3/_1_  (.CLK(\proj__3.net17 ),
    .RESET_B(net393),
    .D(\proj__3.net18 ),
    .Q_N(\proj__3.net18 ),
    .Q(\proj__3.net19 ));
 sg13g2_tiehi \proj__4.flop1/_1__341  (.L_HI(net394));
 sg13g2_or2_1 \proj__3.or1/_0_  (.X(\proj__3.net8 ),
    .B(\proj__3.net23 ),
    .A(\proj__3.net28 ));
 sg13g2_and2_1 \proj__4.and1/_0_  (.A(net323),
    .B(net175),
    .X(\proj__4.net40 ));
 sg13g2_and2_1 \proj__4.and2/_0_  (.A(\proj__4.net40 ),
    .B(net167),
    .X(\proj__4.net41 ));
 sg13g2_and2_1 \proj__4.and3/_0_  (.A(\proj__4.net41 ),
    .B(net164),
    .X(\proj__4.net42 ));
 sg13g2_and2_1 \proj__4.and5/_0_  (.A(net168),
    .B(net178),
    .X(\proj__4.net139 ));
 sg13g2_and2_1 \proj__4.and6/_0_  (.A(net162),
    .B(net164),
    .X(\proj__4.net140 ));
 sg13g2_and2_1 \proj__4.and7/_0_  (.A(\proj__4.net140 ),
    .B(\proj__4.net139 ),
    .X(\proj__4.net9 ));
 sg13g2_dfrbp_1 \proj__4.flop1/_1_  (.CLK(clknet_2_0__leaf_clk_regs),
    .RESET_B(net394),
    .D(\proj__4.net35 ),
    .Q_N(\proj__4.flop1/notq ),
    .Q(\proj__4.net16 ));
 sg13g2_tiehi \proj__4.flop2/_1__342  (.L_HI(net395));
 sg13g2_dfrbp_1 \proj__4.flop2/_1_  (.CLK(clknet_2_0__leaf_clk_regs),
    .RESET_B(net395),
    .D(\proj__4.net36 ),
    .Q_N(\proj__4.flop2/notq ),
    .Q(\proj__4.net26 ));
 sg13g2_tiehi \proj__4.flop3/_1__343  (.L_HI(net396));
 sg13g2_dfrbp_1 \proj__4.flop3/_1_  (.CLK(clknet_2_0__leaf_clk_regs),
    .RESET_B(net396),
    .D(\proj__4.net37 ),
    .Q_N(\proj__4.flop3/notq ),
    .Q(\proj__4.net31 ));
 sg13g2_tiehi \proj__4.flop4/_1__344  (.L_HI(net397));
 sg13g2_dfrbp_1 \proj__4.flop4/_1_  (.CLK(clknet_2_0__leaf_clk_regs),
    .RESET_B(net397),
    .D(\proj__4.net38 ),
    .Q_N(\proj__4.flop4/notq ),
    .Q(\proj__4.net34 ));
 sg13g2_buf_2 clkbuf_regs_0_clk (.A(clk),
    .X(clk_regs));
 sg13g2_mux2_1 \proj__4.mux1/_0_  (.A0(net42),
    .A1(net43),
    .S(net177),
    .X(\proj__4.net17 ));
 sg13g2_mux2_1 \proj__4.mux10/_0_  (.A0(\proj__4.net20 ),
    .A1(\proj__4.net21 ),
    .S(net168),
    .X(\proj__4.net28 ));
 sg13g2_mux2_1 \proj__4.mux100/_0_  (.A0(\proj__4.net111 ),
    .A1(\proj__4.net112 ),
    .S(net166),
    .X(\proj__4.net118 ));
 sg13g2_mux2_1 \proj__4.mux101/_0_  (.A0(\proj__4.net113 ),
    .A1(\proj__4.net114 ),
    .S(net168),
    .X(\proj__4.net119 ));
 sg13g2_mux2_1 \proj__4.mux102/_0_  (.A0(\proj__4.net115 ),
    .A1(\proj__4.net116 ),
    .S(net168),
    .X(\proj__4.net120 ));
 sg13g2_mux2_1 \proj__4.mux103/_0_  (.A0(\proj__4.net119 ),
    .A1(\proj__4.net120 ),
    .S(\proj__4.net31 ),
    .X(\proj__4.net121 ));
 sg13g2_mux2_1 \proj__4.mux104/_0_  (.A0(\proj__4.net117 ),
    .A1(\proj__4.net118 ),
    .S(net163),
    .X(\proj__4.net122 ));
 sg13g2_mux2_1 \proj__4.mux105/_0_  (.A0(\proj__4.net122 ),
    .A1(\proj__4.net121 ),
    .S(net162),
    .X(\proj__4.net7 ));
 sg13g2_mux2_1 \proj__4.mux106/_0_  (.A0(net324),
    .A1(net44),
    .S(net174),
    .X(\proj__4.net125 ));
 sg13g2_mux2_1 \proj__4.mux107/_0_  (.A0(net325),
    .A1(net326),
    .S(net174),
    .X(\proj__4.net126 ));
 sg13g2_mux2_1 \proj__4.mux108/_0_  (.A0(net327),
    .A1(net328),
    .S(net173),
    .X(\proj__4.net127 ));
 sg13g2_mux2_1 \proj__4.mux109/_0_  (.A0(net329),
    .A1(net330),
    .S(net173),
    .X(\proj__4.net128 ));
 sg13g2_mux2_1 \proj__4.mux11/_0_  (.A0(\proj__4.net22 ),
    .A1(\proj__4.net23 ),
    .S(net168),
    .X(\proj__4.net29 ));
 sg13g2_mux2_1 \proj__4.mux110/_0_  (.A0(net331),
    .A1(net45),
    .S(net171),
    .X(\proj__4.net129 ));
 sg13g2_mux2_1 \proj__4.mux111/_0_  (.A0(net332),
    .A1(net333),
    .S(net171),
    .X(\proj__4.net130 ));
 sg13g2_mux2_1 \proj__4.mux112/_0_  (.A0(net334),
    .A1(net335),
    .S(net171),
    .X(\proj__4.net131 ));
 sg13g2_mux2_1 \proj__4.mux113/_0_  (.A0(net336),
    .A1(net337),
    .S(net171),
    .X(\proj__4.net132 ));
 sg13g2_mux2_1 \proj__4.mux114/_0_  (.A0(\proj__4.net125 ),
    .A1(\proj__4.net126 ),
    .S(net166),
    .X(\proj__4.net133 ));
 sg13g2_mux2_1 \proj__4.mux115/_0_  (.A0(\proj__4.net127 ),
    .A1(\proj__4.net128 ),
    .S(net166),
    .X(\proj__4.net134 ));
 sg13g2_mux2_1 \proj__4.mux116/_0_  (.A0(\proj__4.net129 ),
    .A1(\proj__4.net130 ),
    .S(net165),
    .X(\proj__4.net135 ));
 sg13g2_mux2_1 \proj__4.mux117/_0_  (.A0(\proj__4.net131 ),
    .A1(\proj__4.net132 ),
    .S(net165),
    .X(\proj__4.net136 ));
 sg13g2_mux2_1 \proj__4.mux118/_0_  (.A0(\proj__4.net135 ),
    .A1(\proj__4.net136 ),
    .S(net163),
    .X(\proj__4.net137 ));
 sg13g2_mux2_1 \proj__4.mux119/_0_  (.A0(\proj__4.net133 ),
    .A1(\proj__4.net134 ),
    .S(net164),
    .X(\proj__4.net138 ));
 sg13g2_mux2_1 \proj__4.mux12/_0_  (.A0(\proj__4.net24 ),
    .A1(\proj__4.net25 ),
    .S(net168),
    .X(\proj__4.net30 ));
 sg13g2_mux2_1 \proj__4.mux120/_0_  (.A0(\proj__4.net138 ),
    .A1(\proj__4.net137 ),
    .S(net162),
    .X(\proj__4.net8 ));
 sg13g2_mux2_1 \proj__4.mux13/_0_  (.A0(\proj__4.net29 ),
    .A1(\proj__4.net30 ),
    .S(net164),
    .X(\proj__4.net32 ));
 sg13g2_mux2_1 \proj__4.mux14/_0_  (.A0(\proj__4.net27 ),
    .A1(\proj__4.net28 ),
    .S(net164),
    .X(\proj__4.net33 ));
 sg13g2_mux2_1 \proj__4.mux15/_0_  (.A0(\proj__4.net33 ),
    .A1(\proj__4.net32 ),
    .S(net162),
    .X(\proj__4.net2 ));
 sg13g2_mux2_1 \proj__4.mux2/_0_  (.A0(net46),
    .A1(net47),
    .S(net177),
    .X(\proj__4.net18 ));
 sg13g2_mux2_1 \proj__4.mux3/_0_  (.A0(net48),
    .A1(net338),
    .S(net177),
    .X(\proj__4.net20 ));
 sg13g2_mux2_1 \proj__4.mux31/_0_  (.A0(net49),
    .A1(net50),
    .S(net173),
    .X(\proj__4.net44 ));
 sg13g2_mux2_1 \proj__4.mux32/_0_  (.A0(net51),
    .A1(net339),
    .S(net173),
    .X(\proj__4.net46 ));
 sg13g2_mux2_1 \proj__4.mux33/_0_  (.A0(net52),
    .A1(net340),
    .S(net173),
    .X(\proj__4.net47 ));
 sg13g2_mux2_1 \proj__4.mux34/_0_  (.A0(net341),
    .A1(net342),
    .S(net173),
    .X(\proj__4.net48 ));
 sg13g2_mux2_1 \proj__4.mux35/_0_  (.A0(net53),
    .A1(net54),
    .S(net174),
    .X(\proj__4.net49 ));
 sg13g2_mux2_1 \proj__4.mux36/_0_  (.A0(net55),
    .A1(net56),
    .S(net174),
    .X(\proj__4.net50 ));
 sg13g2_mux2_1 \proj__4.mux37/_0_  (.A0(net57),
    .A1(net58),
    .S(net173),
    .X(\proj__4.net51 ));
 sg13g2_mux2_1 \proj__4.mux38/_0_  (.A0(net343),
    .A1(net59),
    .S(net173),
    .X(\proj__4.net52 ));
 sg13g2_mux2_1 \proj__4.mux39/_0_  (.A0(\proj__4.net44 ),
    .A1(\proj__4.net46 ),
    .S(net166),
    .X(\proj__4.net53 ));
 sg13g2_mux2_1 \proj__4.mux4/_0_  (.A0(net344),
    .A1(net345),
    .S(net177),
    .X(\proj__4.net21 ));
 sg13g2_mux2_1 \proj__4.mux40/_0_  (.A0(\proj__4.net47 ),
    .A1(\proj__4.net48 ),
    .S(net166),
    .X(\proj__4.net54 ));
 sg13g2_mux2_1 \proj__4.mux41/_0_  (.A0(\proj__4.net49 ),
    .A1(\proj__4.net50 ),
    .S(net166),
    .X(\proj__4.net55 ));
 sg13g2_mux2_1 \proj__4.mux42/_0_  (.A0(\proj__4.net51 ),
    .A1(\proj__4.net52 ),
    .S(net166),
    .X(\proj__4.net56 ));
 sg13g2_mux2_1 \proj__4.mux43/_0_  (.A0(\proj__4.net55 ),
    .A1(\proj__4.net56 ),
    .S(net163),
    .X(\proj__4.net57 ));
 sg13g2_mux2_1 \proj__4.mux44/_0_  (.A0(\proj__4.net53 ),
    .A1(\proj__4.net54 ),
    .S(net163),
    .X(\proj__4.net58 ));
 sg13g2_mux2_1 \proj__4.mux45/_0_  (.A0(\proj__4.net58 ),
    .A1(\proj__4.net57 ),
    .S(net162),
    .X(\proj__4.net3 ));
 sg13g2_mux2_1 \proj__4.mux46/_0_  (.A0(net60),
    .A1(net61),
    .S(net175),
    .X(\proj__4.net60 ));
 sg13g2_mux2_1 \proj__4.mux47/_0_  (.A0(net346),
    .A1(net347),
    .S(net176),
    .X(\proj__4.net62 ));
 sg13g2_mux2_1 \proj__4.mux48/_0_  (.A0(net62),
    .A1(net348),
    .S(net175),
    .X(\proj__4.net63 ));
 sg13g2_mux2_1 \proj__4.mux49/_0_  (.A0(net63),
    .A1(net64),
    .S(net176),
    .X(\proj__4.net64 ));
 sg13g2_mux2_1 \proj__4.mux5/_0_  (.A0(net65),
    .A1(net66),
    .S(net178),
    .X(\proj__4.net22 ));
 sg13g2_mux2_1 \proj__4.mux50/_0_  (.A0(net349),
    .A1(net350),
    .S(net176),
    .X(\proj__4.net65 ));
 sg13g2_mux2_1 \proj__4.mux51/_0_  (.A0(net67),
    .A1(net68),
    .S(net176),
    .X(\proj__4.net66 ));
 sg13g2_mux2_1 \proj__4.mux52/_0_  (.A0(net351),
    .A1(net69),
    .S(net176),
    .X(\proj__4.net67 ));
 sg13g2_mux2_1 \proj__4.mux53/_0_  (.A0(net352),
    .A1(net353),
    .S(net176),
    .X(\proj__4.net68 ));
 sg13g2_mux2_1 \proj__4.mux54/_0_  (.A0(\proj__4.net60 ),
    .A1(\proj__4.net62 ),
    .S(net167),
    .X(\proj__4.net69 ));
 sg13g2_mux2_1 \proj__4.mux55/_0_  (.A0(\proj__4.net63 ),
    .A1(\proj__4.net64 ),
    .S(net167),
    .X(\proj__4.net70 ));
 sg13g2_mux2_1 \proj__4.mux56/_0_  (.A0(\proj__4.net65 ),
    .A1(\proj__4.net66 ),
    .S(net167),
    .X(\proj__4.net71 ));
 sg13g2_mux2_1 \proj__4.mux57/_0_  (.A0(\proj__4.net67 ),
    .A1(\proj__4.net68 ),
    .S(net167),
    .X(\proj__4.net72 ));
 sg13g2_mux2_1 \proj__4.mux58/_0_  (.A0(\proj__4.net71 ),
    .A1(\proj__4.net72 ),
    .S(net164),
    .X(\proj__4.net73 ));
 sg13g2_mux2_1 \proj__4.mux59/_0_  (.A0(\proj__4.net69 ),
    .A1(\proj__4.net70 ),
    .S(\proj__4.net31 ),
    .X(\proj__4.net74 ));
 sg13g2_mux2_1 \proj__4.mux6/_0_  (.A0(net70),
    .A1(net71),
    .S(net178),
    .X(\proj__4.net23 ));
 sg13g2_mux2_1 \proj__4.mux60/_0_  (.A0(\proj__4.net74 ),
    .A1(\proj__4.net73 ),
    .S(net162),
    .X(\proj__4.net4 ));
 sg13g2_mux2_1 \proj__4.mux61/_0_  (.A0(net354),
    .A1(net72),
    .S(net172),
    .X(\proj__4.net77 ));
 sg13g2_mux2_1 \proj__4.mux62/_0_  (.A0(net73),
    .A1(net355),
    .S(net172),
    .X(\proj__4.net78 ));
 sg13g2_mux2_1 \proj__4.mux63/_0_  (.A0(net356),
    .A1(net357),
    .S(net172),
    .X(\proj__4.net79 ));
 sg13g2_mux2_1 \proj__4.mux64/_0_  (.A0(net74),
    .A1(net358),
    .S(net172),
    .X(\proj__4.net80 ));
 sg13g2_mux2_1 \proj__4.mux65/_0_  (.A0(net359),
    .A1(net360),
    .S(net175),
    .X(\proj__4.net81 ));
 sg13g2_mux2_1 \proj__4.mux66/_0_  (.A0(net361),
    .A1(net75),
    .S(net175),
    .X(\proj__4.net82 ));
 sg13g2_mux2_1 \proj__4.mux67/_0_  (.A0(net362),
    .A1(net363),
    .S(net175),
    .X(\proj__4.net83 ));
 sg13g2_mux2_1 \proj__4.mux68/_0_  (.A0(net76),
    .A1(net364),
    .S(net175),
    .X(\proj__4.net84 ));
 sg13g2_mux2_1 \proj__4.mux69/_0_  (.A0(\proj__4.net77 ),
    .A1(\proj__4.net78 ),
    .S(net165),
    .X(\proj__4.net85 ));
 sg13g2_mux2_1 \proj__4.mux7/_0_  (.A0(net77),
    .A1(net78),
    .S(net178),
    .X(\proj__4.net24 ));
 sg13g2_mux2_1 \proj__4.mux70/_0_  (.A0(\proj__4.net79 ),
    .A1(\proj__4.net80 ),
    .S(net165),
    .X(\proj__4.net86 ));
 sg13g2_mux2_1 \proj__4.mux71/_0_  (.A0(\proj__4.net81 ),
    .A1(\proj__4.net82 ),
    .S(net167),
    .X(\proj__4.net87 ));
 sg13g2_mux2_1 \proj__4.mux72/_0_  (.A0(\proj__4.net83 ),
    .A1(\proj__4.net84 ),
    .S(net167),
    .X(\proj__4.net88 ));
 sg13g2_mux2_1 \proj__4.mux73/_0_  (.A0(\proj__4.net87 ),
    .A1(\proj__4.net88 ),
    .S(net163),
    .X(\proj__4.net89 ));
 sg13g2_mux2_1 \proj__4.mux74/_0_  (.A0(\proj__4.net85 ),
    .A1(\proj__4.net86 ),
    .S(net163),
    .X(\proj__4.net90 ));
 sg13g2_mux2_1 \proj__4.mux75/_0_  (.A0(\proj__4.net90 ),
    .A1(\proj__4.net89 ),
    .S(net162),
    .X(\proj__4.net5 ));
 sg13g2_mux2_1 \proj__4.mux76/_0_  (.A0(net365),
    .A1(net366),
    .S(net170),
    .X(\proj__4.net92 ));
 sg13g2_mux2_1 \proj__4.mux77/_0_  (.A0(net367),
    .A1(net79),
    .S(net170),
    .X(\proj__4.net94 ));
 sg13g2_mux2_1 \proj__4.mux78/_0_  (.A0(net368),
    .A1(net369),
    .S(net170),
    .X(\proj__4.net95 ));
 sg13g2_mux2_1 \proj__4.mux79/_0_  (.A0(net370),
    .A1(net371),
    .S(net170),
    .X(\proj__4.net96 ));
 sg13g2_mux2_1 \proj__4.mux8/_0_  (.A0(net80),
    .A1(net372),
    .S(net178),
    .X(\proj__4.net25 ));
 sg13g2_mux2_1 \proj__4.mux80/_0_  (.A0(net373),
    .A1(net374),
    .S(net170),
    .X(\proj__4.net97 ));
 sg13g2_mux2_1 \proj__4.mux81/_0_  (.A0(net375),
    .A1(net376),
    .S(net170),
    .X(\proj__4.net98 ));
 sg13g2_mux2_1 \proj__4.mux82/_0_  (.A0(net377),
    .A1(net378),
    .S(net170),
    .X(\proj__4.net99 ));
 sg13g2_mux2_1 \proj__4.mux83/_0_  (.A0(net379),
    .A1(net81),
    .S(net170),
    .X(\proj__4.net100 ));
 sg13g2_mux2_1 \proj__4.mux84/_0_  (.A0(\proj__4.net92 ),
    .A1(\proj__4.net94 ),
    .S(net165),
    .X(\proj__4.net101 ));
 sg13g2_mux2_1 \proj__4.mux85/_0_  (.A0(\proj__4.net95 ),
    .A1(\proj__4.net96 ),
    .S(net165),
    .X(\proj__4.net102 ));
 sg13g2_mux2_1 \proj__4.mux86/_0_  (.A0(\proj__4.net97 ),
    .A1(\proj__4.net98 ),
    .S(net165),
    .X(\proj__4.net103 ));
 sg13g2_mux2_1 \proj__4.mux87/_0_  (.A0(\proj__4.net99 ),
    .A1(\proj__4.net100 ),
    .S(net165),
    .X(\proj__4.net104 ));
 sg13g2_mux2_1 \proj__4.mux88/_0_  (.A0(\proj__4.net103 ),
    .A1(\proj__4.net104 ),
    .S(net163),
    .X(\proj__4.net105 ));
 sg13g2_mux2_1 \proj__4.mux89/_0_  (.A0(\proj__4.net101 ),
    .A1(\proj__4.net102 ),
    .S(net163),
    .X(\proj__4.net106 ));
 sg13g2_mux2_1 \proj__4.mux9/_0_  (.A0(\proj__4.net17 ),
    .A1(\proj__4.net18 ),
    .S(net168),
    .X(\proj__4.net27 ));
 sg13g2_mux2_1 \proj__4.mux90/_0_  (.A0(\proj__4.net106 ),
    .A1(\proj__4.net105 ),
    .S(net162),
    .X(\proj__4.net6 ));
 sg13g2_mux2_1 \proj__4.mux91/_0_  (.A0(net380),
    .A1(net82),
    .S(net180),
    .X(\proj__4.net109 ));
 sg13g2_mux2_1 \proj__4.mux92/_0_  (.A0(net83),
    .A1(net381),
    .S(net174),
    .X(\proj__4.net110 ));
 sg13g2_mux2_1 \proj__4.mux93/_0_  (.A0(net382),
    .A1(net84),
    .S(net174),
    .X(\proj__4.net111 ));
 sg13g2_mux2_1 \proj__4.mux94/_0_  (.A0(net383),
    .A1(net384),
    .S(net174),
    .X(\proj__4.net112 ));
 sg13g2_mux2_1 \proj__4.mux95/_0_  (.A0(net85),
    .A1(net86),
    .S(net177),
    .X(\proj__4.net113 ));
 sg13g2_mux2_1 \proj__4.mux96/_0_  (.A0(net385),
    .A1(net87),
    .S(net177),
    .X(\proj__4.net114 ));
 sg13g2_mux2_1 \proj__4.mux97/_0_  (.A0(net88),
    .A1(net89),
    .S(net177),
    .X(\proj__4.net115 ));
 sg13g2_mux2_1 \proj__4.mux98/_0_  (.A0(net386),
    .A1(net387),
    .S(net177),
    .X(\proj__4.net116 ));
 sg13g2_mux2_1 \proj__4.mux99/_0_  (.A0(\proj__4.net109 ),
    .A1(\proj__4.net110 ),
    .S(net166),
    .X(\proj__4.net117 ));
 sg13g2_xor2_1 \proj__4.xor1/_0_  (.B(net175),
    .A(net388),
    .X(\proj__4.net35 ));
 sg13g2_xor2_1 \proj__4.xor2/_0_  (.B(net167),
    .A(\proj__4.net40 ),
    .X(\proj__4.net36 ));
 sg13g2_xor2_1 \proj__4.xor3/_0_  (.B(net164),
    .A(\proj__4.net41 ),
    .X(\proj__4.net37 ));
 sg13g2_xor2_1 \proj__4.xor4/_0_  (.B(net400),
    .A(\proj__4.net42 ),
    .X(\proj__4.net38 ));
 sg13g2_and2_1 \proj__5.and1/_0_  (.A(net201),
    .B(net203),
    .X(\proj__5.net12 ));
 sg13g2_and2_1 \proj__5.and2/_0_  (.A(net194),
    .B(net196),
    .X(\proj__5.net13 ));
 sg13g2_and2_1 \proj__5.and3/_0_  (.A(net186),
    .B(\proj__5.net13 ),
    .X(\proj__5.net14 ));
 sg13g2_and2_1 \proj__5.and4/_0_  (.A(\proj__5.net14 ),
    .B(\proj__5.net12 ),
    .X(\proj__5.net6 ));
 sg13g2_and2_1 \proj__6.and1/_0_  (.A(\proj__6.net61 ),
    .B(\proj__6.net62 ),
    .X(\proj__6.net63 ));
 sg13g2_and2_2 \proj__6.and10/_0_  (.A(\proj__6.net64 ),
    .B(net194),
    .X(\proj__6.net32 ));
 sg13g2_and2_2 \proj__6.and11/_0_  (.A(\proj__6.net65 ),
    .B(net194),
    .X(\proj__6.net42 ));
 sg13g2_and2_2 \proj__6.and12/_0_  (.A(\proj__6.net66 ),
    .B(net194),
    .X(\proj__6.net52 ));
 sg13g2_and2_1 \proj__6.and13/_0_  (.A(net184),
    .B(\proj__6.net74 ),
    .X(\proj__6.net10 ));
 sg13g2_and2_1 \proj__6.and14/_0_  (.A(net186),
    .B(\proj__6.net76 ),
    .X(\proj__6.net11 ));
 sg13g2_and2_1 \proj__6.and15/_0_  (.A(net184),
    .B(\proj__6.net78 ),
    .X(\proj__6.net12 ));
 sg13g2_and2_1 \proj__6.and16/_0_  (.A(net184),
    .B(\proj__6.net80 ),
    .X(\proj__6.net13 ));
 sg13g2_and2_1 \proj__6.and17/_0_  (.A(net186),
    .B(\proj__6.net82 ),
    .X(\proj__6.net14 ));
 sg13g2_and2_1 \proj__6.and18/_0_  (.A(net185),
    .B(\proj__6.net84 ),
    .X(\proj__6.net15 ));
 sg13g2_and2_1 \proj__6.and19/_0_  (.A(net184),
    .B(\proj__6.net86 ),
    .X(\proj__6.net16 ));
 sg13g2_and2_1 \proj__6.and2/_0_  (.A(net203),
    .B(net201),
    .X(\proj__6.net66 ));
 sg13g2_and2_1 \proj__6.and20/_0_  (.A(net186),
    .B(\proj__6.net88 ),
    .X(\proj__6.net17 ));
 sg13g2_and2_1 \proj__6.and3/_0_  (.A(net196),
    .B(\proj__6.net63 ),
    .X(\proj__6.net20 ));
 sg13g2_and2_1 \proj__6.and4/_0_  (.A(net203),
    .B(\proj__6.net62 ),
    .X(\proj__6.net64 ));
 sg13g2_and2_1 \proj__6.and5/_0_  (.A(net198),
    .B(\proj__6.net66 ),
    .X(\proj__6.net51 ));
 sg13g2_and2_1 \proj__6.and6/_0_  (.A(net196),
    .B(\proj__6.net64 ),
    .X(\proj__6.net31 ));
 sg13g2_and2_1 \proj__6.and7/_0_  (.A(\proj__6.net61 ),
    .B(net201),
    .X(\proj__6.net65 ));
 sg13g2_and2_2 \proj__6.and8/_0_  (.A(\proj__6.net63 ),
    .B(net194),
    .X(\proj__6.net21 ));
 sg13g2_and2_1 \proj__6.and9/_0_  (.A(net196),
    .B(\proj__6.net65 ),
    .X(\proj__6.net41 ));
 sg13g2_inv_1 \proj__6.flop0/_4_  (.Y(\proj__6.flop0/_0_ ),
    .A(net207));
 sg13g2_inv_1 \proj__6.flop0/_5_  (.Y(\proj__6.flop0/_1_ ),
    .A(net90));
 sg13g2_tielo \proj__6.flop0/dffsr_183  (.L_LO(net236));
 sg13g2_tielo \proj__6.flop1/dffsr_184  (.L_LO(net237));
 sg13g2_sdfbbp_1 \proj__6.flop0/dffsr  (.Q(\proj__6.net23 ),
    .Q_N(\proj__6.flop0/notq ),
    .RESET_B(\proj__6.flop0/_0_ ),
    .SET_B(\proj__6.flop0/_1_ ),
    .D(\proj__6.net20 ),
    .SCE(net236),
    .SCD(net235),
    .CLK(\proj__6.net21 ));
 sg13g2_inv_1 \proj__6.flop1/_4_  (.Y(\proj__6.flop1/_0_ ),
    .A(net207));
 sg13g2_inv_1 \proj__6.flop1/_5_  (.Y(\proj__6.flop1/_1_ ),
    .A(net91));
 sg13g2_tielo \proj__6.flop1/dffsr_185  (.L_LO(net238));
 sg13g2_tielo \proj__6.flop10/dffsr_186  (.L_LO(net239));
 sg13g2_sdfbbp_1 \proj__6.flop1/dffsr  (.Q(\proj__6.net24 ),
    .Q_N(\proj__6.flop1/notq ),
    .RESET_B(\proj__6.flop1/_0_ ),
    .SET_B(\proj__6.flop1/_1_ ),
    .D(\proj__6.net23 ),
    .SCE(net238),
    .SCD(net237),
    .CLK(\proj__6.net21 ));
 sg13g2_inv_1 \proj__6.flop10/_4_  (.Y(\proj__6.flop10/_0_ ),
    .A(net209));
 sg13g2_inv_1 \proj__6.flop10/_5_  (.Y(\proj__6.flop10/_1_ ),
    .A(net92));
 sg13g2_tielo \proj__6.flop10/dffsr_187  (.L_LO(net240));
 sg13g2_tielo \proj__6.flop11/dffsr_188  (.L_LO(net241));
 sg13g2_sdfbbp_1 \proj__6.flop10/dffsr  (.Q(\proj__6.net36 ),
    .Q_N(\proj__6.flop10/notq ),
    .RESET_B(\proj__6.flop10/_0_ ),
    .SET_B(\proj__6.flop10/_1_ ),
    .D(\proj__6.net35 ),
    .SCE(net240),
    .SCD(net239),
    .CLK(\proj__6.net32 ));
 sg13g2_inv_1 \proj__6.flop11/_4_  (.Y(\proj__6.flop11/_0_ ),
    .A(net208));
 sg13g2_inv_1 \proj__6.flop11/_5_  (.Y(\proj__6.flop11/_1_ ),
    .A(net93));
 sg13g2_tielo \proj__6.flop11/dffsr_189  (.L_LO(net242));
 sg13g2_tielo \proj__6.flop12/dffsr_190  (.L_LO(net243));
 sg13g2_sdfbbp_1 \proj__6.flop11/dffsr  (.Q(\proj__6.net35 ),
    .Q_N(\proj__6.flop11/notq ),
    .RESET_B(\proj__6.flop11/_0_ ),
    .SET_B(\proj__6.flop11/_1_ ),
    .D(\proj__6.net37 ),
    .SCE(net242),
    .SCD(net241),
    .CLK(\proj__6.net32 ));
 sg13g2_inv_1 \proj__6.flop12/_4_  (.Y(\proj__6.flop12/_0_ ),
    .A(net206));
 sg13g2_inv_1 \proj__6.flop12/_5_  (.Y(\proj__6.flop12/_1_ ),
    .A(net94));
 sg13g2_tielo \proj__6.flop12/dffsr_191  (.L_LO(net244));
 sg13g2_tielo \proj__6.flop13/dffsr_192  (.L_LO(net245));
 sg13g2_sdfbbp_1 \proj__6.flop12/dffsr  (.Q(\proj__6.net38 ),
    .Q_N(\proj__6.flop12/notq ),
    .RESET_B(\proj__6.flop12/_0_ ),
    .SET_B(\proj__6.flop12/_1_ ),
    .D(\proj__6.net34 ),
    .SCE(net244),
    .SCD(net243),
    .CLK(\proj__6.net32 ));
 sg13g2_inv_1 \proj__6.flop13/_4_  (.Y(\proj__6.flop13/_0_ ),
    .A(net206));
 sg13g2_inv_1 \proj__6.flop13/_5_  (.Y(\proj__6.flop13/_1_ ),
    .A(net95));
 sg13g2_tielo \proj__6.flop13/dffsr_193  (.L_LO(net246));
 sg13g2_tielo \proj__6.flop14/dffsr_194  (.L_LO(net247));
 sg13g2_sdfbbp_1 \proj__6.flop13/dffsr  (.Q(\proj__6.net39 ),
    .Q_N(\proj__6.flop13/notq ),
    .RESET_B(\proj__6.flop13/_0_ ),
    .SET_B(\proj__6.flop13/_1_ ),
    .D(\proj__6.net38 ),
    .SCE(net246),
    .SCD(net245),
    .CLK(\proj__6.net32 ));
 sg13g2_inv_1 \proj__6.flop14/_4_  (.Y(\proj__6.flop14/_0_ ),
    .A(net206));
 sg13g2_inv_1 \proj__6.flop14/_5_  (.Y(\proj__6.flop14/_1_ ),
    .A(net96));
 sg13g2_tielo \proj__6.flop14/dffsr_195  (.L_LO(net248));
 sg13g2_tielo \proj__6.flop15/dffsr_196  (.L_LO(net249));
 sg13g2_sdfbbp_1 \proj__6.flop14/dffsr  (.Q(\proj__6.net40 ),
    .Q_N(\proj__6.flop14/notq ),
    .RESET_B(\proj__6.flop14/_0_ ),
    .SET_B(\proj__6.flop14/_1_ ),
    .D(\proj__6.net39 ),
    .SCE(net248),
    .SCD(net247),
    .CLK(\proj__6.net32 ));
 sg13g2_inv_1 \proj__6.flop15/_4_  (.Y(\proj__6.flop15/_0_ ),
    .A(net206));
 sg13g2_inv_1 \proj__6.flop15/_5_  (.Y(\proj__6.flop15/_1_ ),
    .A(net97));
 sg13g2_tielo \proj__6.flop15/dffsr_197  (.L_LO(net250));
 sg13g2_tielo \proj__6.flop16/dffsr_198  (.L_LO(net251));
 sg13g2_sdfbbp_1 \proj__6.flop15/dffsr  (.Q(\proj__6.net37 ),
    .Q_N(\proj__6.flop15/notq ),
    .RESET_B(\proj__6.flop15/_0_ ),
    .SET_B(\proj__6.flop15/_1_ ),
    .D(\proj__6.net40 ),
    .SCE(net250),
    .SCD(net249),
    .CLK(\proj__6.net32 ));
 sg13g2_inv_1 \proj__6.flop16/_4_  (.Y(\proj__6.flop16/_0_ ),
    .A(net208));
 sg13g2_inv_1 \proj__6.flop16/_5_  (.Y(\proj__6.flop16/_1_ ),
    .A(net98));
 sg13g2_tielo \proj__6.flop16/dffsr_199  (.L_LO(net252));
 sg13g2_tielo \proj__6.flop17/dffsr_200  (.L_LO(net253));
 sg13g2_sdfbbp_1 \proj__6.flop16/dffsr  (.Q(\proj__6.net43 ),
    .Q_N(\proj__6.flop16/notq ),
    .RESET_B(\proj__6.flop16/_0_ ),
    .SET_B(\proj__6.flop16/_1_ ),
    .D(\proj__6.net41 ),
    .SCE(net252),
    .SCD(net251),
    .CLK(\proj__6.net42 ));
 sg13g2_inv_1 \proj__6.flop17/_4_  (.Y(\proj__6.flop17/_0_ ),
    .A(net211));
 sg13g2_inv_1 \proj__6.flop17/_5_  (.Y(\proj__6.flop17/_1_ ),
    .A(net99));
 sg13g2_tielo \proj__6.flop17/dffsr_201  (.L_LO(net254));
 sg13g2_tielo \proj__6.flop18/dffsr_202  (.L_LO(net255));
 sg13g2_sdfbbp_1 \proj__6.flop17/dffsr  (.Q(\proj__6.net44 ),
    .Q_N(\proj__6.flop17/notq ),
    .RESET_B(\proj__6.flop17/_0_ ),
    .SET_B(\proj__6.flop17/_1_ ),
    .D(\proj__6.net43 ),
    .SCE(net254),
    .SCD(net253),
    .CLK(\proj__6.net42 ));
 sg13g2_inv_1 \proj__6.flop18/_4_  (.Y(\proj__6.flop18/_0_ ),
    .A(net210));
 sg13g2_inv_1 \proj__6.flop18/_5_  (.Y(\proj__6.flop18/_1_ ),
    .A(net100));
 sg13g2_tielo \proj__6.flop18/dffsr_203  (.L_LO(net256));
 sg13g2_tielo \proj__6.flop19/dffsr_204  (.L_LO(net257));
 sg13g2_sdfbbp_1 \proj__6.flop18/dffsr  (.Q(\proj__6.net46 ),
    .Q_N(\proj__6.flop18/notq ),
    .RESET_B(\proj__6.flop18/_0_ ),
    .SET_B(\proj__6.flop18/_1_ ),
    .D(\proj__6.net45 ),
    .SCE(net256),
    .SCD(net255),
    .CLK(\proj__6.net42 ));
 sg13g2_inv_1 \proj__6.flop19/_4_  (.Y(\proj__6.flop19/_0_ ),
    .A(net210));
 sg13g2_inv_1 \proj__6.flop19/_5_  (.Y(\proj__6.flop19/_1_ ),
    .A(net101));
 sg13g2_tielo \proj__6.flop19/dffsr_205  (.L_LO(net258));
 sg13g2_tielo \proj__6.flop2/dffsr_206  (.L_LO(net259));
 sg13g2_sdfbbp_1 \proj__6.flop19/dffsr  (.Q(\proj__6.net45 ),
    .Q_N(\proj__6.flop19/notq ),
    .RESET_B(\proj__6.flop19/_0_ ),
    .SET_B(\proj__6.flop19/_1_ ),
    .D(\proj__6.net47 ),
    .SCE(net258),
    .SCD(net257),
    .CLK(\proj__6.net42 ));
 sg13g2_inv_1 \proj__6.flop2/_4_  (.Y(\proj__6.flop2/_0_ ),
    .A(net209));
 sg13g2_inv_1 \proj__6.flop2/_5_  (.Y(\proj__6.flop2/_1_ ),
    .A(net102));
 sg13g2_tielo \proj__6.flop2/dffsr_207  (.L_LO(net260));
 sg13g2_tielo \proj__6.flop20/dffsr_208  (.L_LO(net261));
 sg13g2_sdfbbp_1 \proj__6.flop2/dffsr  (.Q(\proj__6.net26 ),
    .Q_N(\proj__6.flop2/notq ),
    .RESET_B(\proj__6.flop2/_0_ ),
    .SET_B(\proj__6.flop2/_1_ ),
    .D(\proj__6.net25 ),
    .SCE(net260),
    .SCD(net259),
    .CLK(\proj__6.net21 ));
 sg13g2_inv_1 \proj__6.flop20/_4_  (.Y(\proj__6.flop20/_0_ ),
    .A(net211));
 sg13g2_inv_1 \proj__6.flop20/_5_  (.Y(\proj__6.flop20/_1_ ),
    .A(net103));
 sg13g2_tielo \proj__6.flop20/dffsr_209  (.L_LO(net262));
 sg13g2_tielo \proj__6.flop21/dffsr_210  (.L_LO(net263));
 sg13g2_sdfbbp_1 \proj__6.flop20/dffsr  (.Q(\proj__6.net48 ),
    .Q_N(\proj__6.flop20/notq ),
    .RESET_B(\proj__6.flop20/_0_ ),
    .SET_B(\proj__6.flop20/_1_ ),
    .D(\proj__6.net44 ),
    .SCE(net262),
    .SCD(net261),
    .CLK(\proj__6.net42 ));
 sg13g2_inv_1 \proj__6.flop21/_4_  (.Y(\proj__6.flop21/_0_ ),
    .A(net211));
 sg13g2_inv_1 \proj__6.flop21/_5_  (.Y(\proj__6.flop21/_1_ ),
    .A(net104));
 sg13g2_tielo \proj__6.flop21/dffsr_211  (.L_LO(net264));
 sg13g2_tielo \proj__6.flop22/dffsr_212  (.L_LO(net265));
 sg13g2_sdfbbp_1 \proj__6.flop21/dffsr  (.Q(\proj__6.net49 ),
    .Q_N(\proj__6.flop21/notq ),
    .RESET_B(\proj__6.flop21/_0_ ),
    .SET_B(\proj__6.flop21/_1_ ),
    .D(\proj__6.net48 ),
    .SCE(net264),
    .SCD(net263),
    .CLK(\proj__6.net42 ));
 sg13g2_inv_1 \proj__6.flop22/_4_  (.Y(\proj__6.flop22/_0_ ),
    .A(net211));
 sg13g2_inv_1 \proj__6.flop22/_5_  (.Y(\proj__6.flop22/_1_ ),
    .A(net105));
 sg13g2_tielo \proj__6.flop22/dffsr_213  (.L_LO(net266));
 sg13g2_tielo \proj__6.flop23/dffsr_214  (.L_LO(net267));
 sg13g2_sdfbbp_1 \proj__6.flop22/dffsr  (.Q(\proj__6.net50 ),
    .Q_N(\proj__6.flop22/notq ),
    .RESET_B(\proj__6.flop22/_0_ ),
    .SET_B(\proj__6.flop22/_1_ ),
    .D(\proj__6.net49 ),
    .SCE(net266),
    .SCD(net265),
    .CLK(\proj__6.net42 ));
 sg13g2_inv_1 \proj__6.flop23/_4_  (.Y(\proj__6.flop23/_0_ ),
    .A(net210));
 sg13g2_inv_1 \proj__6.flop23/_5_  (.Y(\proj__6.flop23/_1_ ),
    .A(net106));
 sg13g2_tielo \proj__6.flop23/dffsr_215  (.L_LO(net268));
 sg13g2_tielo \proj__6.flop24/dffsr_216  (.L_LO(net269));
 sg13g2_sdfbbp_1 \proj__6.flop23/dffsr  (.Q(\proj__6.net47 ),
    .Q_N(\proj__6.flop23/notq ),
    .RESET_B(\proj__6.flop23/_0_ ),
    .SET_B(\proj__6.flop23/_1_ ),
    .D(\proj__6.net50 ),
    .SCE(net268),
    .SCD(net267),
    .CLK(\proj__6.net42 ));
 sg13g2_inv_1 \proj__6.flop24/_4_  (.Y(\proj__6.flop24/_0_ ),
    .A(net211));
 sg13g2_inv_1 \proj__6.flop24/_5_  (.Y(\proj__6.flop24/_1_ ),
    .A(net107));
 sg13g2_tielo \proj__6.flop24/dffsr_217  (.L_LO(net270));
 sg13g2_tielo \proj__6.flop25/dffsr_218  (.L_LO(net271));
 sg13g2_sdfbbp_1 \proj__6.flop24/dffsr  (.Q(\proj__6.net53 ),
    .Q_N(\proj__6.flop24/notq ),
    .RESET_B(\proj__6.flop24/_0_ ),
    .SET_B(\proj__6.flop24/_1_ ),
    .D(\proj__6.net51 ),
    .SCE(net270),
    .SCD(net269),
    .CLK(\proj__6.net52 ));
 sg13g2_inv_1 \proj__6.flop25/_4_  (.Y(\proj__6.flop25/_0_ ),
    .A(net212));
 sg13g2_inv_1 \proj__6.flop25/_5_  (.Y(\proj__6.flop25/_1_ ),
    .A(net108));
 sg13g2_tielo \proj__6.flop25/dffsr_219  (.L_LO(net272));
 sg13g2_tielo \proj__6.flop26/dffsr_220  (.L_LO(net273));
 sg13g2_sdfbbp_1 \proj__6.flop25/dffsr  (.Q(\proj__6.net54 ),
    .Q_N(\proj__6.flop25/notq ),
    .RESET_B(\proj__6.flop25/_0_ ),
    .SET_B(\proj__6.flop25/_1_ ),
    .D(\proj__6.net53 ),
    .SCE(net272),
    .SCD(net271),
    .CLK(\proj__6.net52 ));
 sg13g2_inv_1 \proj__6.flop26/_4_  (.Y(\proj__6.flop26/_0_ ),
    .A(net210));
 sg13g2_inv_1 \proj__6.flop26/_5_  (.Y(\proj__6.flop26/_1_ ),
    .A(net109));
 sg13g2_tielo \proj__6.flop26/dffsr_221  (.L_LO(net274));
 sg13g2_tielo \proj__6.flop27/dffsr_222  (.L_LO(net275));
 sg13g2_sdfbbp_1 \proj__6.flop26/dffsr  (.Q(\proj__6.net56 ),
    .Q_N(\proj__6.flop26/notq ),
    .RESET_B(\proj__6.flop26/_0_ ),
    .SET_B(\proj__6.flop26/_1_ ),
    .D(\proj__6.net55 ),
    .SCE(net274),
    .SCD(net273),
    .CLK(\proj__6.net52 ));
 sg13g2_inv_1 \proj__6.flop27/_4_  (.Y(\proj__6.flop27/_0_ ),
    .A(net210));
 sg13g2_inv_1 \proj__6.flop27/_5_  (.Y(\proj__6.flop27/_1_ ),
    .A(net110));
 sg13g2_tielo \proj__6.flop27/dffsr_223  (.L_LO(net276));
 sg13g2_tielo \proj__6.flop28/dffsr_224  (.L_LO(net277));
 sg13g2_sdfbbp_1 \proj__6.flop27/dffsr  (.Q(\proj__6.net55 ),
    .Q_N(\proj__6.flop27/notq ),
    .RESET_B(\proj__6.flop27/_0_ ),
    .SET_B(\proj__6.flop27/_1_ ),
    .D(\proj__6.net57 ),
    .SCE(net276),
    .SCD(net275),
    .CLK(\proj__6.net52 ));
 sg13g2_inv_1 \proj__6.flop28/_4_  (.Y(\proj__6.flop28/_0_ ),
    .A(net212));
 sg13g2_inv_1 \proj__6.flop28/_5_  (.Y(\proj__6.flop28/_1_ ),
    .A(net111));
 sg13g2_tielo \proj__6.flop28/dffsr_225  (.L_LO(net278));
 sg13g2_tielo \proj__6.flop29/dffsr_226  (.L_LO(net279));
 sg13g2_sdfbbp_1 \proj__6.flop28/dffsr  (.Q(\proj__6.net58 ),
    .Q_N(\proj__6.flop28/notq ),
    .RESET_B(\proj__6.flop28/_0_ ),
    .SET_B(\proj__6.flop28/_1_ ),
    .D(\proj__6.net54 ),
    .SCE(net278),
    .SCD(net277),
    .CLK(\proj__6.net52 ));
 sg13g2_inv_1 \proj__6.flop29/_4_  (.Y(\proj__6.flop29/_0_ ),
    .A(net210));
 sg13g2_inv_1 \proj__6.flop29/_5_  (.Y(\proj__6.flop29/_1_ ),
    .A(net112));
 sg13g2_tielo \proj__6.flop29/dffsr_227  (.L_LO(net280));
 sg13g2_tielo \proj__6.flop3/dffsr_228  (.L_LO(net281));
 sg13g2_sdfbbp_1 \proj__6.flop29/dffsr  (.Q(\proj__6.net59 ),
    .Q_N(\proj__6.flop29/notq ),
    .RESET_B(\proj__6.flop29/_0_ ),
    .SET_B(\proj__6.flop29/_1_ ),
    .D(\proj__6.net58 ),
    .SCE(net280),
    .SCD(net279),
    .CLK(\proj__6.net52 ));
 sg13g2_inv_1 \proj__6.flop3/_4_  (.Y(\proj__6.flop3/_0_ ),
    .A(net208));
 sg13g2_inv_1 \proj__6.flop3/_5_  (.Y(\proj__6.flop3/_1_ ),
    .A(net113));
 sg13g2_tielo \proj__6.flop3/dffsr_229  (.L_LO(net282));
 sg13g2_tielo \proj__6.flop30/dffsr_230  (.L_LO(net283));
 sg13g2_sdfbbp_1 \proj__6.flop3/dffsr  (.Q(\proj__6.net25 ),
    .Q_N(\proj__6.flop3/notq ),
    .RESET_B(\proj__6.flop3/_0_ ),
    .SET_B(\proj__6.flop3/_1_ ),
    .D(\proj__6.net27 ),
    .SCE(net282),
    .SCD(net281),
    .CLK(\proj__6.net21 ));
 sg13g2_inv_1 \proj__6.flop30/_4_  (.Y(\proj__6.flop30/_0_ ),
    .A(net211));
 sg13g2_inv_1 \proj__6.flop30/_5_  (.Y(\proj__6.flop30/_1_ ),
    .A(net114));
 sg13g2_tielo \proj__6.flop30/dffsr_231  (.L_LO(net284));
 sg13g2_tielo \proj__6.flop31/dffsr_232  (.L_LO(net285));
 sg13g2_sdfbbp_1 \proj__6.flop30/dffsr  (.Q(\proj__6.net60 ),
    .Q_N(\proj__6.flop30/notq ),
    .RESET_B(\proj__6.flop30/_0_ ),
    .SET_B(\proj__6.flop30/_1_ ),
    .D(\proj__6.net59 ),
    .SCE(net284),
    .SCD(net283),
    .CLK(\proj__6.net52 ));
 sg13g2_inv_1 \proj__6.flop31/_4_  (.Y(\proj__6.flop31/_0_ ),
    .A(net210));
 sg13g2_inv_1 \proj__6.flop31/_5_  (.Y(\proj__6.flop31/_1_ ),
    .A(net115));
 sg13g2_tielo \proj__6.flop31/dffsr_233  (.L_LO(net286));
 sg13g2_tielo \proj__6.flop33/dffsr_234  (.L_LO(net287));
 sg13g2_sdfbbp_1 \proj__6.flop31/dffsr  (.Q(\proj__6.net57 ),
    .Q_N(\proj__6.flop31/notq ),
    .RESET_B(\proj__6.flop31/_0_ ),
    .SET_B(\proj__6.flop31/_1_ ),
    .D(\proj__6.net60 ),
    .SCE(net286),
    .SCD(net285),
    .CLK(\proj__6.net52 ));
 sg13g2_inv_1 \proj__6.flop33/_4_  (.Y(\proj__6.flop33/_0_ ),
    .A(net209));
 sg13g2_inv_1 \proj__6.flop33/_5_  (.Y(\proj__6.flop33/_1_ ),
    .A(net116));
 sg13g2_tielo \proj__6.flop33/dffsr_235  (.L_LO(net288));
 sg13g2_tielo \proj__6.flop34/dffsr_236  (.L_LO(net289));
 sg13g2_sdfbbp_1 \proj__6.flop33/dffsr  (.Q(\proj__6.net74 ),
    .Q_N(\proj__6.flop33/notq ),
    .RESET_B(\proj__6.flop33/_0_ ),
    .SET_B(\proj__6.flop33/_1_ ),
    .D(\proj__6.net72 ),
    .SCE(net288),
    .SCD(net287),
    .CLK(net191));
 sg13g2_inv_1 \proj__6.flop34/_4_  (.Y(\proj__6.flop34/_0_ ),
    .A(net209));
 sg13g2_inv_1 \proj__6.flop34/_5_  (.Y(\proj__6.flop34/_1_ ),
    .A(net117));
 sg13g2_tielo \proj__6.flop34/dffsr_237  (.L_LO(net290));
 sg13g2_tielo \proj__6.flop35/dffsr_238  (.L_LO(net291));
 sg13g2_sdfbbp_1 \proj__6.flop34/dffsr  (.Q(\proj__6.net76 ),
    .Q_N(\proj__6.flop34/notq ),
    .RESET_B(\proj__6.flop34/_0_ ),
    .SET_B(\proj__6.flop34/_1_ ),
    .D(\proj__6.net75 ),
    .SCE(net290),
    .SCD(net289),
    .CLK(net192));
 sg13g2_inv_1 \proj__6.flop35/_4_  (.Y(\proj__6.flop35/_0_ ),
    .A(net208));
 sg13g2_inv_1 \proj__6.flop35/_5_  (.Y(\proj__6.flop35/_1_ ),
    .A(net118));
 sg13g2_tielo \proj__6.flop35/dffsr_239  (.L_LO(net292));
 sg13g2_tielo \proj__6.flop36/dffsr_240  (.L_LO(net293));
 sg13g2_sdfbbp_1 \proj__6.flop35/dffsr  (.Q(\proj__6.net78 ),
    .Q_N(\proj__6.flop35/notq ),
    .RESET_B(\proj__6.flop35/_0_ ),
    .SET_B(\proj__6.flop35/_1_ ),
    .D(\proj__6.net77 ),
    .SCE(net292),
    .SCD(net291),
    .CLK(net191));
 sg13g2_inv_1 \proj__6.flop36/_4_  (.Y(\proj__6.flop36/_0_ ),
    .A(net208));
 sg13g2_inv_1 \proj__6.flop36/_5_  (.Y(\proj__6.flop36/_1_ ),
    .A(net119));
 sg13g2_tielo \proj__6.flop36/dffsr_241  (.L_LO(net294));
 sg13g2_tielo \proj__6.flop37/dffsr_242  (.L_LO(net295));
 sg13g2_sdfbbp_1 \proj__6.flop36/dffsr  (.Q(\proj__6.net80 ),
    .Q_N(\proj__6.flop36/notq ),
    .RESET_B(\proj__6.flop36/_0_ ),
    .SET_B(\proj__6.flop36/_1_ ),
    .D(\proj__6.net79 ),
    .SCE(net294),
    .SCD(net293),
    .CLK(net191));
 sg13g2_inv_1 \proj__6.flop37/_4_  (.Y(\proj__6.flop37/_0_ ),
    .A(net211));
 sg13g2_inv_1 \proj__6.flop37/_5_  (.Y(\proj__6.flop37/_1_ ),
    .A(net120));
 sg13g2_tielo \proj__6.flop37/dffsr_243  (.L_LO(net296));
 sg13g2_tielo \proj__6.flop38/dffsr_244  (.L_LO(net297));
 sg13g2_sdfbbp_1 \proj__6.flop37/dffsr  (.Q(\proj__6.net82 ),
    .Q_N(\proj__6.flop37/notq ),
    .RESET_B(\proj__6.flop37/_0_ ),
    .SET_B(\proj__6.flop37/_1_ ),
    .D(\proj__6.net81 ),
    .SCE(net296),
    .SCD(net295),
    .CLK(net191));
 sg13g2_inv_1 \proj__6.flop38/_4_  (.Y(\proj__6.flop38/_0_ ),
    .A(net209));
 sg13g2_inv_1 \proj__6.flop38/_5_  (.Y(\proj__6.flop38/_1_ ),
    .A(net121));
 sg13g2_tielo \proj__6.flop38/dffsr_245  (.L_LO(net298));
 sg13g2_tielo \proj__6.flop39/dffsr_246  (.L_LO(net299));
 sg13g2_sdfbbp_1 \proj__6.flop38/dffsr  (.Q(\proj__6.net84 ),
    .Q_N(\proj__6.flop38/notq ),
    .RESET_B(\proj__6.flop38/_0_ ),
    .SET_B(\proj__6.flop38/_1_ ),
    .D(\proj__6.net83 ),
    .SCE(net298),
    .SCD(net297),
    .CLK(net191));
 sg13g2_inv_1 \proj__6.flop39/_4_  (.Y(\proj__6.flop39/_0_ ),
    .A(net208));
 sg13g2_inv_1 \proj__6.flop39/_5_  (.Y(\proj__6.flop39/_1_ ),
    .A(net122));
 sg13g2_tielo \proj__6.flop39/dffsr_247  (.L_LO(net300));
 sg13g2_tielo \proj__6.flop4/dffsr_248  (.L_LO(net301));
 sg13g2_sdfbbp_1 \proj__6.flop39/dffsr  (.Q(\proj__6.net86 ),
    .Q_N(\proj__6.flop39/notq ),
    .RESET_B(\proj__6.flop39/_0_ ),
    .SET_B(\proj__6.flop39/_1_ ),
    .D(\proj__6.net85 ),
    .SCE(net300),
    .SCD(net299),
    .CLK(net191));
 sg13g2_inv_1 \proj__6.flop4/_4_  (.Y(\proj__6.flop4/_0_ ),
    .A(net206));
 sg13g2_inv_1 \proj__6.flop4/_5_  (.Y(\proj__6.flop4/_1_ ),
    .A(net123));
 sg13g2_tielo \proj__6.flop4/dffsr_249  (.L_LO(net302));
 sg13g2_tielo \proj__6.flop40/dffsr_250  (.L_LO(net303));
 sg13g2_sdfbbp_1 \proj__6.flop4/dffsr  (.Q(\proj__6.net28 ),
    .Q_N(\proj__6.flop4/notq ),
    .RESET_B(\proj__6.flop4/_0_ ),
    .SET_B(\proj__6.flop4/_1_ ),
    .D(\proj__6.net24 ),
    .SCE(net302),
    .SCD(net301),
    .CLK(\proj__6.net21 ));
 sg13g2_inv_1 \proj__6.flop40/_4_  (.Y(\proj__6.flop40/_0_ ),
    .A(net212));
 sg13g2_inv_1 \proj__6.flop40/_5_  (.Y(\proj__6.flop40/_1_ ),
    .A(net124));
 sg13g2_tielo \proj__6.flop40/dffsr_251  (.L_LO(net304));
 sg13g2_tielo \proj__6.flop5/dffsr_252  (.L_LO(net305));
 sg13g2_sdfbbp_1 \proj__6.flop40/dffsr  (.Q(\proj__6.net88 ),
    .Q_N(\proj__6.flop40/notq ),
    .RESET_B(\proj__6.flop40/_0_ ),
    .SET_B(\proj__6.flop40/_1_ ),
    .D(\proj__6.net87 ),
    .SCE(net304),
    .SCD(net303),
    .CLK(net191));
 sg13g2_inv_1 \proj__6.flop5/_4_  (.Y(\proj__6.flop5/_0_ ),
    .A(net206));
 sg13g2_inv_1 \proj__6.flop5/_5_  (.Y(\proj__6.flop5/_1_ ),
    .A(net125));
 sg13g2_tielo \proj__6.flop5/dffsr_253  (.L_LO(net306));
 sg13g2_tielo \proj__6.flop6/dffsr_254  (.L_LO(net307));
 sg13g2_sdfbbp_1 \proj__6.flop5/dffsr  (.Q(\proj__6.net29 ),
    .Q_N(\proj__6.flop5/notq ),
    .RESET_B(\proj__6.flop5/_0_ ),
    .SET_B(\proj__6.flop5/_1_ ),
    .D(\proj__6.net28 ),
    .SCE(net306),
    .SCD(net305),
    .CLK(\proj__6.net21 ));
 sg13g2_inv_1 \proj__6.flop6/_4_  (.Y(\proj__6.flop6/_0_ ),
    .A(net206));
 sg13g2_inv_1 \proj__6.flop6/_5_  (.Y(\proj__6.flop6/_1_ ),
    .A(net126));
 sg13g2_tielo \proj__6.flop6/dffsr_255  (.L_LO(net308));
 sg13g2_tielo \proj__6.flop7/dffsr_256  (.L_LO(net309));
 sg13g2_sdfbbp_1 \proj__6.flop6/dffsr  (.Q(\proj__6.net30 ),
    .Q_N(\proj__6.flop6/notq ),
    .RESET_B(\proj__6.flop6/_0_ ),
    .SET_B(\proj__6.flop6/_1_ ),
    .D(\proj__6.net29 ),
    .SCE(net308),
    .SCD(net307),
    .CLK(\proj__6.net21 ));
 sg13g2_inv_1 \proj__6.flop7/_4_  (.Y(\proj__6.flop7/_0_ ),
    .A(net206));
 sg13g2_inv_1 \proj__6.flop7/_5_  (.Y(\proj__6.flop7/_1_ ),
    .A(net127));
 sg13g2_tielo \proj__6.flop7/dffsr_257  (.L_LO(net310));
 sg13g2_tielo \proj__6.flop8/dffsr_258  (.L_LO(net311));
 sg13g2_sdfbbp_1 \proj__6.flop7/dffsr  (.Q(\proj__6.net27 ),
    .Q_N(\proj__6.flop7/notq ),
    .RESET_B(\proj__6.flop7/_0_ ),
    .SET_B(\proj__6.flop7/_1_ ),
    .D(\proj__6.net30 ),
    .SCE(net310),
    .SCD(net309),
    .CLK(\proj__6.net21 ));
 sg13g2_inv_1 \proj__6.flop8/_4_  (.Y(\proj__6.flop8/_0_ ),
    .A(net207));
 sg13g2_inv_1 \proj__6.flop8/_5_  (.Y(\proj__6.flop8/_1_ ),
    .A(net128));
 sg13g2_tielo \proj__6.flop8/dffsr_259  (.L_LO(net312));
 sg13g2_tielo \proj__6.flop9/dffsr_260  (.L_LO(net313));
 sg13g2_sdfbbp_1 \proj__6.flop8/dffsr  (.Q(\proj__6.net33 ),
    .Q_N(\proj__6.flop8/notq ),
    .RESET_B(\proj__6.flop8/_0_ ),
    .SET_B(\proj__6.flop8/_1_ ),
    .D(\proj__6.net31 ),
    .SCE(net312),
    .SCD(net311),
    .CLK(\proj__6.net32 ));
 sg13g2_inv_1 \proj__6.flop9/_4_  (.Y(\proj__6.flop9/_0_ ),
    .A(net207));
 sg13g2_inv_1 \proj__6.flop9/_5_  (.Y(\proj__6.flop9/_1_ ),
    .A(net129));
 sg13g2_tielo \proj__6.flop9/dffsr_261  (.L_LO(net314));
 sg13g2_tielo \proj__9.flop1/dffsr_262  (.L_LO(net315));
 sg13g2_sdfbbp_1 \proj__6.flop9/dffsr  (.Q(\proj__6.net34 ),
    .Q_N(\proj__6.flop9/notq ),
    .RESET_B(\proj__6.flop9/_0_ ),
    .SET_B(\proj__6.flop9/_1_ ),
    .D(\proj__6.net33 ),
    .SCE(net314),
    .SCD(net313),
    .CLK(\proj__6.net32 ));
 sg13g2_mux2_1 \proj__6.mux1/_0_  (.A0(\proj__6.net53 ),
    .A1(\proj__6.net43 ),
    .S(net160),
    .X(\proj__6.net91 ));
 sg13g2_mux2_1 \proj__6.mux10/_0_  (.A0(\proj__6.net59 ),
    .A1(\proj__6.net49 ),
    .S(net161),
    .X(\proj__6.net98 ));
 sg13g2_mux2_1 \proj__6.mux11/_0_  (.A0(\proj__6.net39 ),
    .A1(\proj__6.net29 ),
    .S(net160),
    .X(\proj__6.net99 ));
 sg13g2_mux2_1 \proj__6.mux12/_0_  (.A0(\proj__6.net98 ),
    .A1(\proj__6.net99 ),
    .S(\proj__6.net93 ),
    .X(\proj__6.net79 ));
 sg13g2_mux2_1 \proj__6.mux13/_0_  (.A0(\proj__6.net60 ),
    .A1(\proj__6.net50 ),
    .S(net161),
    .X(\proj__6.net100 ));
 sg13g2_mux2_1 \proj__6.mux14/_0_  (.A0(\proj__6.net40 ),
    .A1(\proj__6.net30 ),
    .S(net160),
    .X(\proj__6.net101 ));
 sg13g2_mux2_1 \proj__6.mux15/_0_  (.A0(\proj__6.net100 ),
    .A1(\proj__6.net101 ),
    .S(\proj__6.net93 ),
    .X(\proj__6.net81 ));
 sg13g2_mux2_1 \proj__6.mux16/_0_  (.A0(\proj__6.net57 ),
    .A1(\proj__6.net47 ),
    .S(net161),
    .X(\proj__6.net102 ));
 sg13g2_mux2_1 \proj__6.mux17/_0_  (.A0(\proj__6.net37 ),
    .A1(\proj__6.net27 ),
    .S(net160),
    .X(\proj__6.net103 ));
 sg13g2_mux2_1 \proj__6.mux18/_0_  (.A0(\proj__6.net102 ),
    .A1(\proj__6.net103 ),
    .S(\proj__6.net93 ),
    .X(\proj__6.net83 ));
 sg13g2_mux2_1 \proj__6.mux19/_0_  (.A0(\proj__6.net55 ),
    .A1(\proj__6.net45 ),
    .S(net161),
    .X(\proj__6.net104 ));
 sg13g2_mux2_1 \proj__6.mux2/_0_  (.A0(\proj__6.net54 ),
    .A1(\proj__6.net44 ),
    .S(\proj__6.net90 ),
    .X(\proj__6.net94 ));
 sg13g2_mux2_1 \proj__6.mux20/_0_  (.A0(\proj__6.net35 ),
    .A1(\proj__6.net25 ),
    .S(net161),
    .X(\proj__6.net105 ));
 sg13g2_mux2_1 \proj__6.mux21/_0_  (.A0(\proj__6.net104 ),
    .A1(\proj__6.net105 ),
    .S(\proj__6.net93 ),
    .X(\proj__6.net85 ));
 sg13g2_mux2_1 \proj__6.mux22/_0_  (.A0(\proj__6.net56 ),
    .A1(\proj__6.net46 ),
    .S(net161),
    .X(\proj__6.net106 ));
 sg13g2_mux2_1 \proj__6.mux23/_0_  (.A0(\proj__6.net36 ),
    .A1(\proj__6.net26 ),
    .S(net160),
    .X(\proj__6.net107 ));
 sg13g2_mux2_1 \proj__6.mux24/_0_  (.A0(\proj__6.net106 ),
    .A1(\proj__6.net107 ),
    .S(\proj__6.net93 ),
    .X(\proj__6.net87 ));
 sg13g2_mux2_1 \proj__6.mux3/_0_  (.A0(\proj__6.net34 ),
    .A1(\proj__6.net24 ),
    .S(net160),
    .X(\proj__6.net95 ));
 sg13g2_mux2_1 \proj__6.mux4/_0_  (.A0(\proj__6.net94 ),
    .A1(\proj__6.net95 ),
    .S(\proj__6.net93 ),
    .X(\proj__6.net75 ));
 sg13g2_mux2_1 \proj__6.mux5/_0_  (.A0(\proj__6.net33 ),
    .A1(\proj__6.net23 ),
    .S(net160),
    .X(\proj__6.net92 ));
 sg13g2_mux2_1 \proj__6.mux6/_0_  (.A0(\proj__6.net58 ),
    .A1(\proj__6.net48 ),
    .S(net161),
    .X(\proj__6.net96 ));
 sg13g2_mux2_1 \proj__6.mux7/_0_  (.A0(\proj__6.net38 ),
    .A1(\proj__6.net28 ),
    .S(net160),
    .X(\proj__6.net97 ));
 sg13g2_mux2_1 \proj__6.mux8/_0_  (.A0(\proj__6.net96 ),
    .A1(\proj__6.net97 ),
    .S(\proj__6.net93 ),
    .X(\proj__6.net77 ));
 sg13g2_mux2_1 \proj__6.mux9/_0_  (.A0(\proj__6.net91 ),
    .A1(\proj__6.net92 ),
    .S(\proj__6.net93 ),
    .X(\proj__6.net72 ));
 sg13g2_inv_1 \proj__6.not1/_0_  (.Y(\proj__6.net61 ),
    .A(net203));
 sg13g2_inv_1 \proj__6.not2/_0_  (.Y(\proj__6.net62 ),
    .A(net201));
 sg13g2_inv_1 \proj__6.not3/_0_  (.Y(\proj__6.net90 ),
    .A(net189));
 sg13g2_inv_4 \proj__6.not4/_0_  (.A(net187),
    .Y(\proj__6.net93 ));
 sg13g2_nand2_1 \proj__7.nand1/_0_  (.Y(\proj__7.net11 ),
    .A(net200),
    .B(net203));
 sg13g2_nand2_1 \proj__7.nand2/_0_  (.Y(\proj__7.net12 ),
    .A(net197),
    .B(net200));
 sg13g2_nand2_1 \proj__7.nand3/_0_  (.Y(\proj__7.net4 ),
    .A(\proj__7.net5 ),
    .B(\proj__7.net11 ));
 sg13g2_nand2_1 \proj__7.nand4/_0_  (.Y(\proj__7.net5 ),
    .A(\proj__7.net12 ),
    .B(\proj__7.net4 ));
 sg13g2_and2_1 \proj__9.and1/_0_  (.A(net200),
    .B(\proj__9.net16 ),
    .X(\proj__9.net5 ));
 sg13g2_and2_1 \proj__9.and2/_0_  (.A(net200),
    .B(\proj__9.net18 ),
    .X(\proj__9.net6 ));
 sg13g2_and2_1 \proj__9.and3/_0_  (.A(net200),
    .B(\proj__9.net19 ),
    .X(\proj__9.net7 ));
 sg13g2_and2_1 \proj__9.and4/_0_  (.A(net202),
    .B(\proj__9.net20 ),
    .X(\proj__9.net8 ));
 sg13g2_inv_1 \proj__9.flop1/_4_  (.Y(\proj__9.flop1/_0_ ),
    .A(\proj__9.net15 ));
 sg13g2_inv_1 \proj__9.flop1/_5_  (.Y(\proj__9.flop1/_1_ ),
    .A(net130));
 sg13g2_tielo \proj__9.flop1/dffsr_263  (.L_LO(net316));
 sg13g2_tielo \proj__9.flop2/dffsr_264  (.L_LO(net317));
 sg13g2_sdfbbp_1 \proj__9.flop1/dffsr  (.Q(\proj__9.net16 ),
    .Q_N(\proj__9.flop1/notq ),
    .RESET_B(\proj__9.flop1/_0_ ),
    .SET_B(\proj__9.flop1/_1_ ),
    .D(net203),
    .SCE(net316),
    .SCD(net315),
    .CLK(clknet_2_1__leaf_clk_regs));
 sg13g2_inv_1 \proj__9.flop2/_4_  (.Y(\proj__9.flop2/_0_ ),
    .A(\proj__9.net15 ));
 sg13g2_inv_1 \proj__9.flop2/_5_  (.Y(\proj__9.flop2/_1_ ),
    .A(net131));
 sg13g2_tielo \proj__9.flop2/dffsr_265  (.L_LO(net318));
 sg13g2_tielo \proj__9.flop3/dffsr_266  (.L_LO(net319));
 sg13g2_sdfbbp_1 \proj__9.flop2/dffsr  (.Q(\proj__9.net18 ),
    .Q_N(\proj__9.flop2/notq ),
    .RESET_B(\proj__9.flop2/_0_ ),
    .SET_B(\proj__9.flop2/_1_ ),
    .D(net404),
    .SCE(net318),
    .SCD(net317),
    .CLK(clknet_2_1__leaf_clk_regs));
 sg13g2_inv_1 \proj__9.flop3/_4_  (.Y(\proj__9.flop3/_0_ ),
    .A(\proj__9.net15 ));
 sg13g2_inv_1 \proj__9.flop3/_5_  (.Y(\proj__9.flop3/_1_ ),
    .A(net132));
 sg13g2_tielo \proj__9.flop3/dffsr_267  (.L_LO(net320));
 sg13g2_tielo \proj__9.flop4/dffsr_268  (.L_LO(net321));
 sg13g2_sdfbbp_1 \proj__9.flop3/dffsr  (.Q(\proj__9.net19 ),
    .Q_N(\proj__9.flop3/notq ),
    .RESET_B(\proj__9.flop3/_0_ ),
    .SET_B(\proj__9.flop3/_1_ ),
    .D(net405),
    .SCE(net320),
    .SCD(net319),
    .CLK(clknet_2_1__leaf_clk_regs));
 sg13g2_inv_1 \proj__9.flop4/_4_  (.Y(\proj__9.flop4/_0_ ),
    .A(\proj__9.net15 ));
 sg13g2_inv_1 \proj__9.flop4/_5_  (.Y(\proj__9.flop4/_1_ ),
    .A(net133));
 sg13g2_tielo \proj__9.flop4/dffsr_269  (.L_LO(net322));
 sg13g2_tiehi \proj__4.and1/_0__270  (.L_HI(net323));
 sg13g2_sdfbbp_1 \proj__9.flop4/dffsr  (.Q(\proj__9.net20 ),
    .Q_N(\proj__9.flop4/notq ),
    .RESET_B(\proj__9.flop4/_0_ ),
    .SET_B(\proj__9.flop4/_1_ ),
    .D(net407),
    .SCE(net322),
    .SCD(net321),
    .CLK(clknet_2_1__leaf_clk_regs));
 sg13g2_inv_1 \proj__9.not1/_0_  (.Y(\proj__9.net15 ),
    .A(net212));
 sg13g2_buf_4 fanout160 (.X(net160),
    .A(net161));
 sg13g2_buf_4 fanout161 (.X(net161),
    .A(\proj__6.net90 ));
 sg13g2_buf_4 fanout162 (.X(net162),
    .A(\proj__4.net34 ));
 sg13g2_buf_4 fanout163 (.X(net163),
    .A(net164));
 sg13g2_buf_4 fanout164 (.X(net164),
    .A(net419));
 sg13g2_buf_4 fanout165 (.X(net165),
    .A(net169));
 sg13g2_buf_4 fanout166 (.X(net166),
    .A(net169));
 sg13g2_buf_4 fanout167 (.X(net167),
    .A(net169));
 sg13g2_buf_4 fanout168 (.X(net168),
    .A(net169));
 sg13g2_buf_2 fanout169 (.A(\proj__4.net26 ),
    .X(net169));
 sg13g2_buf_4 fanout170 (.X(net170),
    .A(net172));
 sg13g2_buf_2 fanout171 (.A(net172),
    .X(net171));
 sg13g2_buf_2 fanout172 (.A(net180),
    .X(net172));
 sg13g2_buf_4 fanout173 (.X(net173),
    .A(net174));
 sg13g2_buf_4 fanout174 (.X(net174),
    .A(net180));
 sg13g2_buf_4 fanout175 (.X(net175),
    .A(net179));
 sg13g2_buf_2 fanout176 (.A(net179),
    .X(net176));
 sg13g2_buf_4 fanout177 (.X(net177),
    .A(net179));
 sg13g2_buf_2 fanout178 (.A(net179),
    .X(net178));
 sg13g2_buf_2 fanout179 (.A(net180),
    .X(net179));
 sg13g2_buf_2 fanout180 (.A(\proj__4.net16 ),
    .X(net180));
 sg13g2_buf_4 fanout181 (.X(net181),
    .A(\proj_10.net59 ));
 sg13g2_buf_2 fanout182 (.A(\proj_10.net59 ),
    .X(net182));
 sg13g2_buf_2 fanout183 (.A(\proj_10.net82 ),
    .X(net183));
 sg13g2_buf_2 fanout184 (.A(net185),
    .X(net184));
 sg13g2_buf_1 fanout185 (.A(net186),
    .X(net185));
 sg13g2_buf_2 fanout186 (.A(ui_in[7]),
    .X(net186));
 sg13g2_buf_4 fanout187 (.X(net187),
    .A(net2));
 sg13g2_buf_4 fanout188 (.X(net188),
    .A(net189));
 sg13g2_buf_1 fanout189 (.A(net190),
    .X(net189));
 sg13g2_buf_2 fanout190 (.A(ui_in[5]),
    .X(net190));
 sg13g2_buf_2 fanout191 (.A(net192),
    .X(net191));
 sg13g2_buf_2 fanout192 (.A(net193),
    .X(net192));
 sg13g2_buf_2 fanout193 (.A(ui_in[4]),
    .X(net193));
 sg13g2_buf_2 fanout194 (.A(net195),
    .X(net194));
 sg13g2_buf_2 fanout195 (.A(net1),
    .X(net195));
 sg13g2_buf_2 fanout196 (.A(net198),
    .X(net196));
 sg13g2_buf_2 fanout197 (.A(net198),
    .X(net197));
 sg13g2_buf_2 fanout198 (.A(ui_in[2]),
    .X(net198));
 sg13g2_buf_2 fanout199 (.A(net200),
    .X(net199));
 sg13g2_buf_2 fanout200 (.A(net201),
    .X(net200));
 sg13g2_buf_2 fanout201 (.A(net202),
    .X(net201));
 sg13g2_buf_2 fanout202 (.A(ui_in[1]),
    .X(net202));
 sg13g2_buf_2 fanout203 (.A(net205),
    .X(net203));
 sg13g2_buf_2 fanout204 (.A(net205),
    .X(net204));
 sg13g2_buf_2 fanout205 (.A(ui_in[0]),
    .X(net205));
 sg13g2_buf_2 fanout206 (.A(net208),
    .X(net206));
 sg13g2_buf_1 fanout207 (.A(net208),
    .X(net207));
 sg13g2_buf_2 fanout208 (.A(net209),
    .X(net208));
 sg13g2_buf_2 fanout209 (.A(rst_n),
    .X(net209));
 sg13g2_buf_2 fanout210 (.A(net211),
    .X(net210));
 sg13g2_buf_2 fanout211 (.A(net212),
    .X(net211));
 sg13g2_buf_4 fanout212 (.X(net212),
    .A(rst_n));
 sg13g2_buf_1 input1 (.A(ui_in[3]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[6]),
    .X(net2));
 sg13g2_buf_4 input3 (.X(net3),
    .A(uio_in[0]));
 sg13g2_buf_2 input4 (.A(uio_in[1]),
    .X(net4));
 sg13g2_buf_2 input5 (.A(uio_in[2]),
    .X(net5));
 sg13g2_buf_2 input6 (.A(uio_in[3]),
    .X(net6));
 sg13g2_tielo \proj_10.flop10/_5__7  (.L_LO(net7));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_2 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .X(clknet_1_0__leaf_clk));
 sg13g2_buf_2 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .X(clknet_1_1__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_1_1__leaf_clk));
 sg13g2_buf_2 clkbuf_0_clk_regs (.A(clk_regs),
    .X(clknet_0_clk_regs));
 sg13g2_buf_2 clkbuf_2_0__f_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_2_0__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_2_1__f_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_2_1__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_2_2__f_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_2_2__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_2_3__f_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_2_3__leaf_clk_regs));
 sg13g2_buf_1 clkload1 (.A(clknet_2_1__leaf_clk_regs));
 sg13g2_buf_1 clkload2 (.A(clknet_2_2__leaf_clk_regs));
 sg13g2_buf_1 clkload3 (.A(clknet_2_3__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_0__015_ (.A(_015_),
    .X(clknet_0__015_));
 sg13g2_buf_2 clkbuf_1_0__f__015_ (.A(clknet_0__015_),
    .X(clknet_1_0__leaf__015_));
 sg13g2_buf_2 clkbuf_1_1__f__015_ (.A(clknet_0__015_),
    .X(clknet_1_1__leaf__015_));
 sg13g2_buf_1 clkload4 (.A(clknet_1_1__leaf__015_));
 sg13g2_dlygate4sd3_1 hold1 (.A(\proj__2.net12 ),
    .X(net398));
 sg13g2_dlygate4sd3_1 hold2 (.A(\proj__3.net14 ),
    .X(net399));
 sg13g2_dlygate4sd3_1 hold3 (.A(\proj__4.net34 ),
    .X(net400));
 sg13g2_dlygate4sd3_1 hold4 (.A(\proj_12.net17 ),
    .X(net401));
 sg13g2_dlygate4sd3_1 hold5 (.A(\proj_10.net54 ),
    .X(net402));
 sg13g2_dlygate4sd3_1 hold6 (.A(\proj_10.net80 ),
    .X(net403));
 sg13g2_dlygate4sd3_1 hold7 (.A(\proj__9.net16 ),
    .X(net404));
 sg13g2_dlygate4sd3_1 hold8 (.A(\proj__9.net18 ),
    .X(net405));
 sg13g2_dlygate4sd3_1 hold9 (.A(\proj_10.net85 ),
    .X(net406));
 sg13g2_dlygate4sd3_1 hold10 (.A(\proj__9.net19 ),
    .X(net407));
 sg13g2_dlygate4sd3_1 hold11 (.A(\proj_10.net83 ),
    .X(net408));
 sg13g2_dlygate4sd3_1 hold12 (.A(\proj_10.net71 ),
    .X(net409));
 sg13g2_dlygate4sd3_1 hold13 (.A(\proj_10.net74 ),
    .X(net410));
 sg13g2_dlygate4sd3_1 hold14 (.A(\proj_10.net28 ),
    .X(net411));
 sg13g2_dlygate4sd3_1 hold15 (.A(\proj_10.net89 ),
    .X(net412));
 sg13g2_dlygate4sd3_1 hold16 (.A(\proj_10.net87 ),
    .X(net413));
 sg13g2_dlygate4sd3_1 hold17 (.A(\proj_10.net48 ),
    .X(net414));
 sg13g2_dlygate4sd3_1 hold18 (.A(\proj_10.net51 ),
    .X(net415));
 sg13g2_dlygate4sd3_1 hold19 (.A(\proj_10.net77 ),
    .X(net416));
 sg13g2_dlygate4sd3_1 hold20 (.A(\proj_10.net33 ),
    .X(net417));
 sg13g2_dlygate4sd3_1 hold21 (.A(\proj_10.net57 ),
    .X(net418));
 sg13g2_dlygate4sd3_1 hold22 (.A(\proj__4.net31 ),
    .X(net419));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_4 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_155 ();
 sg13g2_decap_4 FILLER_12_162 ();
 sg13g2_fill_1 FILLER_12_166 ();
 sg13g2_decap_4 FILLER_12_177 ();
 sg13g2_decap_4 FILLER_12_189 ();
 sg13g2_fill_2 FILLER_12_193 ();
 sg13g2_fill_2 FILLER_12_202 ();
 sg13g2_fill_2 FILLER_12_207 ();
 sg13g2_fill_1 FILLER_12_209 ();
 sg13g2_decap_8 FILLER_12_223 ();
 sg13g2_decap_4 FILLER_12_230 ();
 sg13g2_decap_8 FILLER_12_241 ();
 sg13g2_decap_8 FILLER_12_248 ();
 sg13g2_decap_8 FILLER_12_255 ();
 sg13g2_decap_8 FILLER_12_262 ();
 sg13g2_decap_8 FILLER_12_269 ();
 sg13g2_decap_8 FILLER_12_276 ();
 sg13g2_decap_4 FILLER_12_283 ();
 sg13g2_fill_1 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_291 ();
 sg13g2_decap_8 FILLER_12_298 ();
 sg13g2_decap_8 FILLER_12_305 ();
 sg13g2_decap_8 FILLER_12_312 ();
 sg13g2_decap_8 FILLER_12_319 ();
 sg13g2_decap_8 FILLER_12_326 ();
 sg13g2_decap_8 FILLER_12_333 ();
 sg13g2_decap_8 FILLER_12_340 ();
 sg13g2_decap_8 FILLER_12_347 ();
 sg13g2_decap_8 FILLER_12_354 ();
 sg13g2_decap_8 FILLER_12_361 ();
 sg13g2_decap_8 FILLER_12_368 ();
 sg13g2_decap_8 FILLER_12_375 ();
 sg13g2_decap_8 FILLER_12_382 ();
 sg13g2_decap_8 FILLER_12_389 ();
 sg13g2_decap_8 FILLER_12_396 ();
 sg13g2_decap_4 FILLER_12_403 ();
 sg13g2_fill_2 FILLER_12_407 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_fill_1 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_89 ();
 sg13g2_fill_2 FILLER_13_96 ();
 sg13g2_fill_1 FILLER_13_98 ();
 sg13g2_decap_4 FILLER_13_106 ();
 sg13g2_decap_4 FILLER_13_113 ();
 sg13g2_fill_1 FILLER_13_117 ();
 sg13g2_decap_4 FILLER_13_126 ();
 sg13g2_fill_2 FILLER_13_137 ();
 sg13g2_decap_8 FILLER_13_251 ();
 sg13g2_decap_8 FILLER_13_258 ();
 sg13g2_decap_4 FILLER_13_265 ();
 sg13g2_fill_2 FILLER_13_304 ();
 sg13g2_fill_1 FILLER_13_306 ();
 sg13g2_decap_8 FILLER_13_311 ();
 sg13g2_fill_2 FILLER_13_318 ();
 sg13g2_fill_1 FILLER_13_320 ();
 sg13g2_decap_4 FILLER_13_325 ();
 sg13g2_fill_2 FILLER_13_329 ();
 sg13g2_decap_4 FILLER_13_334 ();
 sg13g2_fill_1 FILLER_13_338 ();
 sg13g2_decap_8 FILLER_13_347 ();
 sg13g2_decap_4 FILLER_13_354 ();
 sg13g2_decap_8 FILLER_13_365 ();
 sg13g2_decap_8 FILLER_13_372 ();
 sg13g2_decap_8 FILLER_13_379 ();
 sg13g2_decap_8 FILLER_13_386 ();
 sg13g2_decap_8 FILLER_13_393 ();
 sg13g2_decap_8 FILLER_13_400 ();
 sg13g2_fill_2 FILLER_13_407 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_fill_2 FILLER_14_77 ();
 sg13g2_fill_1 FILLER_14_79 ();
 sg13g2_decap_4 FILLER_14_119 ();
 sg13g2_fill_2 FILLER_14_123 ();
 sg13g2_decap_8 FILLER_14_128 ();
 sg13g2_decap_4 FILLER_14_138 ();
 sg13g2_fill_1 FILLER_14_145 ();
 sg13g2_decap_8 FILLER_14_156 ();
 sg13g2_fill_2 FILLER_14_166 ();
 sg13g2_decap_8 FILLER_14_171 ();
 sg13g2_decap_8 FILLER_14_188 ();
 sg13g2_fill_2 FILLER_14_195 ();
 sg13g2_decap_4 FILLER_14_200 ();
 sg13g2_fill_2 FILLER_14_204 ();
 sg13g2_decap_8 FILLER_14_209 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_fill_2 FILLER_14_231 ();
 sg13g2_fill_1 FILLER_14_233 ();
 sg13g2_decap_4 FILLER_14_238 ();
 sg13g2_decap_4 FILLER_14_255 ();
 sg13g2_decap_8 FILLER_14_263 ();
 sg13g2_decap_8 FILLER_14_282 ();
 sg13g2_fill_2 FILLER_14_293 ();
 sg13g2_fill_1 FILLER_14_295 ();
 sg13g2_fill_1 FILLER_14_299 ();
 sg13g2_decap_4 FILLER_14_377 ();
 sg13g2_fill_1 FILLER_14_381 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_fill_2 FILLER_14_406 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_fill_2 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_83 ();
 sg13g2_decap_4 FILLER_15_90 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_fill_2 FILLER_15_105 ();
 sg13g2_fill_1 FILLER_15_107 ();
 sg13g2_fill_2 FILLER_15_178 ();
 sg13g2_fill_2 FILLER_15_250 ();
 sg13g2_fill_1 FILLER_15_252 ();
 sg13g2_decap_4 FILLER_15_295 ();
 sg13g2_fill_2 FILLER_15_299 ();
 sg13g2_fill_1 FILLER_15_311 ();
 sg13g2_decap_4 FILLER_15_315 ();
 sg13g2_decap_8 FILLER_15_326 ();
 sg13g2_fill_2 FILLER_15_333 ();
 sg13g2_fill_1 FILLER_15_335 ();
 sg13g2_decap_4 FILLER_15_349 ();
 sg13g2_decap_8 FILLER_15_396 ();
 sg13g2_decap_4 FILLER_15_403 ();
 sg13g2_fill_2 FILLER_15_407 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_4 FILLER_16_70 ();
 sg13g2_fill_2 FILLER_16_117 ();
 sg13g2_fill_1 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_134 ();
 sg13g2_decap_4 FILLER_16_141 ();
 sg13g2_fill_1 FILLER_16_145 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_fill_2 FILLER_16_161 ();
 sg13g2_fill_1 FILLER_16_163 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_4 FILLER_16_193 ();
 sg13g2_fill_1 FILLER_16_197 ();
 sg13g2_decap_8 FILLER_16_202 ();
 sg13g2_decap_4 FILLER_16_209 ();
 sg13g2_decap_8 FILLER_16_223 ();
 sg13g2_fill_2 FILLER_16_230 ();
 sg13g2_fill_1 FILLER_16_232 ();
 sg13g2_fill_2 FILLER_16_236 ();
 sg13g2_fill_1 FILLER_16_238 ();
 sg13g2_decap_8 FILLER_16_259 ();
 sg13g2_fill_1 FILLER_16_266 ();
 sg13g2_decap_4 FILLER_16_280 ();
 sg13g2_decap_4 FILLER_16_357 ();
 sg13g2_decap_8 FILLER_16_375 ();
 sg13g2_fill_2 FILLER_16_382 ();
 sg13g2_fill_2 FILLER_16_388 ();
 sg13g2_decap_8 FILLER_16_400 ();
 sg13g2_fill_2 FILLER_16_407 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_4 FILLER_17_88 ();
 sg13g2_fill_1 FILLER_17_92 ();
 sg13g2_fill_2 FILLER_17_96 ();
 sg13g2_fill_1 FILLER_17_98 ();
 sg13g2_decap_4 FILLER_17_103 ();
 sg13g2_decap_4 FILLER_17_117 ();
 sg13g2_fill_1 FILLER_17_121 ();
 sg13g2_decap_8 FILLER_17_130 ();
 sg13g2_fill_1 FILLER_17_137 ();
 sg13g2_decap_4 FILLER_17_142 ();
 sg13g2_decap_8 FILLER_17_149 ();
 sg13g2_fill_2 FILLER_17_156 ();
 sg13g2_fill_1 FILLER_17_158 ();
 sg13g2_decap_8 FILLER_17_178 ();
 sg13g2_fill_2 FILLER_17_185 ();
 sg13g2_fill_1 FILLER_17_187 ();
 sg13g2_decap_4 FILLER_17_192 ();
 sg13g2_decap_8 FILLER_17_199 ();
 sg13g2_decap_8 FILLER_17_206 ();
 sg13g2_fill_2 FILLER_17_213 ();
 sg13g2_fill_1 FILLER_17_215 ();
 sg13g2_decap_4 FILLER_17_226 ();
 sg13g2_fill_2 FILLER_17_230 ();
 sg13g2_fill_2 FILLER_17_236 ();
 sg13g2_fill_1 FILLER_17_238 ();
 sg13g2_decap_8 FILLER_17_242 ();
 sg13g2_decap_4 FILLER_17_249 ();
 sg13g2_fill_2 FILLER_17_253 ();
 sg13g2_decap_8 FILLER_17_259 ();
 sg13g2_decap_4 FILLER_17_266 ();
 sg13g2_decap_4 FILLER_17_274 ();
 sg13g2_fill_2 FILLER_17_278 ();
 sg13g2_fill_2 FILLER_17_283 ();
 sg13g2_fill_1 FILLER_17_285 ();
 sg13g2_decap_8 FILLER_17_294 ();
 sg13g2_fill_2 FILLER_17_301 ();
 sg13g2_fill_1 FILLER_17_303 ();
 sg13g2_decap_8 FILLER_17_311 ();
 sg13g2_fill_2 FILLER_17_318 ();
 sg13g2_decap_4 FILLER_17_324 ();
 sg13g2_decap_8 FILLER_17_331 ();
 sg13g2_decap_8 FILLER_17_346 ();
 sg13g2_fill_2 FILLER_17_353 ();
 sg13g2_fill_2 FILLER_17_359 ();
 sg13g2_decap_8 FILLER_17_400 ();
 sg13g2_fill_2 FILLER_17_407 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_fill_1 FILLER_18_77 ();
 sg13g2_fill_2 FILLER_18_117 ();
 sg13g2_fill_2 FILLER_18_164 ();
 sg13g2_decap_4 FILLER_18_297 ();
 sg13g2_fill_1 FILLER_18_336 ();
 sg13g2_decap_8 FILLER_18_375 ();
 sg13g2_fill_1 FILLER_18_382 ();
 sg13g2_decap_4 FILLER_18_386 ();
 sg13g2_decap_8 FILLER_18_393 ();
 sg13g2_decap_8 FILLER_18_400 ();
 sg13g2_fill_2 FILLER_18_407 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_4 FILLER_19_84 ();
 sg13g2_fill_1 FILLER_19_88 ();
 sg13g2_decap_4 FILLER_19_93 ();
 sg13g2_fill_1 FILLER_19_97 ();
 sg13g2_decap_4 FILLER_19_101 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_4 FILLER_19_119 ();
 sg13g2_decap_4 FILLER_19_133 ();
 sg13g2_decap_8 FILLER_19_140 ();
 sg13g2_decap_4 FILLER_19_151 ();
 sg13g2_fill_2 FILLER_19_155 ();
 sg13g2_decap_8 FILLER_19_164 ();
 sg13g2_fill_2 FILLER_19_171 ();
 sg13g2_fill_1 FILLER_19_173 ();
 sg13g2_decap_4 FILLER_19_184 ();
 sg13g2_fill_1 FILLER_19_188 ();
 sg13g2_fill_2 FILLER_19_197 ();
 sg13g2_decap_4 FILLER_19_203 ();
 sg13g2_fill_1 FILLER_19_207 ();
 sg13g2_fill_2 FILLER_19_211 ();
 sg13g2_fill_1 FILLER_19_213 ();
 sg13g2_fill_1 FILLER_19_230 ();
 sg13g2_decap_4 FILLER_19_234 ();
 sg13g2_fill_1 FILLER_19_238 ();
 sg13g2_decap_8 FILLER_19_246 ();
 sg13g2_decap_4 FILLER_19_253 ();
 sg13g2_decap_8 FILLER_19_261 ();
 sg13g2_fill_1 FILLER_19_268 ();
 sg13g2_decap_4 FILLER_19_272 ();
 sg13g2_fill_2 FILLER_19_280 ();
 sg13g2_fill_1 FILLER_19_282 ();
 sg13g2_decap_4 FILLER_19_286 ();
 sg13g2_fill_2 FILLER_19_290 ();
 sg13g2_fill_2 FILLER_19_300 ();
 sg13g2_decap_8 FILLER_19_310 ();
 sg13g2_fill_1 FILLER_19_317 ();
 sg13g2_fill_1 FILLER_19_321 ();
 sg13g2_decap_8 FILLER_19_331 ();
 sg13g2_fill_1 FILLER_19_338 ();
 sg13g2_decap_4 FILLER_19_343 ();
 sg13g2_fill_2 FILLER_19_347 ();
 sg13g2_decap_8 FILLER_19_360 ();
 sg13g2_fill_2 FILLER_19_367 ();
 sg13g2_decap_8 FILLER_19_376 ();
 sg13g2_decap_8 FILLER_19_383 ();
 sg13g2_decap_8 FILLER_19_390 ();
 sg13g2_decap_8 FILLER_19_397 ();
 sg13g2_decap_4 FILLER_19_404 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_fill_2 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_27 ();
 sg13g2_decap_8 FILLER_20_34 ();
 sg13g2_decap_4 FILLER_20_41 ();
 sg13g2_decap_8 FILLER_20_59 ();
 sg13g2_decap_8 FILLER_20_66 ();
 sg13g2_decap_8 FILLER_20_73 ();
 sg13g2_fill_2 FILLER_20_80 ();
 sg13g2_fill_1 FILLER_20_82 ();
 sg13g2_decap_4 FILLER_20_125 ();
 sg13g2_fill_2 FILLER_20_129 ();
 sg13g2_fill_2 FILLER_20_176 ();
 sg13g2_fill_2 FILLER_20_217 ();
 sg13g2_fill_1 FILLER_20_219 ();
 sg13g2_fill_1 FILLER_20_255 ();
 sg13g2_fill_1 FILLER_20_291 ();
 sg13g2_fill_2 FILLER_20_302 ();
 sg13g2_decap_8 FILLER_20_307 ();
 sg13g2_fill_2 FILLER_20_317 ();
 sg13g2_decap_8 FILLER_20_328 ();
 sg13g2_decap_8 FILLER_20_335 ();
 sg13g2_fill_2 FILLER_20_346 ();
 sg13g2_decap_4 FILLER_20_383 ();
 sg13g2_fill_1 FILLER_20_387 ();
 sg13g2_decap_8 FILLER_20_391 ();
 sg13g2_decap_8 FILLER_20_398 ();
 sg13g2_decap_4 FILLER_20_405 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_fill_1 FILLER_21_7 ();
 sg13g2_fill_2 FILLER_21_38 ();
 sg13g2_fill_1 FILLER_21_40 ();
 sg13g2_decap_8 FILLER_21_65 ();
 sg13g2_decap_4 FILLER_21_72 ();
 sg13g2_decap_8 FILLER_21_86 ();
 sg13g2_fill_2 FILLER_21_93 ();
 sg13g2_decap_4 FILLER_21_141 ();
 sg13g2_fill_1 FILLER_21_145 ();
 sg13g2_decap_4 FILLER_21_149 ();
 sg13g2_fill_1 FILLER_21_153 ();
 sg13g2_decap_4 FILLER_21_157 ();
 sg13g2_fill_2 FILLER_21_181 ();
 sg13g2_fill_2 FILLER_21_187 ();
 sg13g2_fill_1 FILLER_21_189 ();
 sg13g2_decap_4 FILLER_21_193 ();
 sg13g2_fill_1 FILLER_21_197 ();
 sg13g2_decap_8 FILLER_21_201 ();
 sg13g2_fill_2 FILLER_21_208 ();
 sg13g2_fill_1 FILLER_21_210 ();
 sg13g2_fill_1 FILLER_21_222 ();
 sg13g2_decap_4 FILLER_21_234 ();
 sg13g2_decap_4 FILLER_21_241 ();
 sg13g2_decap_4 FILLER_21_255 ();
 sg13g2_fill_1 FILLER_21_263 ();
 sg13g2_decap_8 FILLER_21_268 ();
 sg13g2_decap_8 FILLER_21_281 ();
 sg13g2_decap_8 FILLER_21_358 ();
 sg13g2_decap_4 FILLER_21_365 ();
 sg13g2_fill_1 FILLER_21_369 ();
 sg13g2_decap_8 FILLER_21_373 ();
 sg13g2_decap_8 FILLER_21_380 ();
 sg13g2_fill_1 FILLER_21_387 ();
 sg13g2_decap_4 FILLER_21_393 ();
 sg13g2_fill_1 FILLER_21_397 ();
 sg13g2_decap_8 FILLER_21_401 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_decap_4 FILLER_22_0 ();
 sg13g2_fill_2 FILLER_22_4 ();
 sg13g2_fill_2 FILLER_22_20 ();
 sg13g2_fill_1 FILLER_22_22 ();
 sg13g2_decap_4 FILLER_22_31 ();
 sg13g2_fill_2 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_59 ();
 sg13g2_decap_8 FILLER_22_66 ();
 sg13g2_decap_4 FILLER_22_73 ();
 sg13g2_decap_8 FILLER_22_87 ();
 sg13g2_decap_4 FILLER_22_94 ();
 sg13g2_decap_4 FILLER_22_106 ();
 sg13g2_fill_2 FILLER_22_110 ();
 sg13g2_decap_8 FILLER_22_119 ();
 sg13g2_decap_8 FILLER_22_126 ();
 sg13g2_fill_2 FILLER_22_168 ();
 sg13g2_fill_2 FILLER_22_209 ();
 sg13g2_decap_4 FILLER_22_235 ();
 sg13g2_fill_1 FILLER_22_239 ();
 sg13g2_decap_4 FILLER_22_279 ();
 sg13g2_fill_1 FILLER_22_283 ();
 sg13g2_fill_2 FILLER_22_303 ();
 sg13g2_decap_8 FILLER_22_309 ();
 sg13g2_fill_2 FILLER_22_316 ();
 sg13g2_fill_1 FILLER_22_318 ();
 sg13g2_fill_1 FILLER_22_322 ();
 sg13g2_decap_4 FILLER_22_327 ();
 sg13g2_fill_2 FILLER_22_331 ();
 sg13g2_fill_2 FILLER_22_346 ();
 sg13g2_decap_8 FILLER_22_351 ();
 sg13g2_decap_8 FILLER_22_358 ();
 sg13g2_decap_8 FILLER_22_365 ();
 sg13g2_decap_8 FILLER_22_372 ();
 sg13g2_decap_4 FILLER_22_379 ();
 sg13g2_fill_1 FILLER_22_383 ();
 sg13g2_fill_2 FILLER_22_406 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_fill_2 FILLER_23_0 ();
 sg13g2_fill_1 FILLER_23_2 ();
 sg13g2_decap_4 FILLER_23_27 ();
 sg13g2_decap_8 FILLER_23_65 ();
 sg13g2_fill_2 FILLER_23_72 ();
 sg13g2_decap_4 FILLER_23_96 ();
 sg13g2_decap_8 FILLER_23_110 ();
 sg13g2_fill_2 FILLER_23_117 ();
 sg13g2_fill_1 FILLER_23_119 ();
 sg13g2_decap_8 FILLER_23_124 ();
 sg13g2_decap_4 FILLER_23_131 ();
 sg13g2_fill_1 FILLER_23_135 ();
 sg13g2_decap_8 FILLER_23_144 ();
 sg13g2_decap_4 FILLER_23_151 ();
 sg13g2_decap_8 FILLER_23_162 ();
 sg13g2_fill_2 FILLER_23_173 ();
 sg13g2_decap_8 FILLER_23_179 ();
 sg13g2_fill_1 FILLER_23_186 ();
 sg13g2_decap_4 FILLER_23_195 ();
 sg13g2_fill_1 FILLER_23_199 ();
 sg13g2_decap_8 FILLER_23_203 ();
 sg13g2_fill_2 FILLER_23_210 ();
 sg13g2_fill_1 FILLER_23_212 ();
 sg13g2_fill_2 FILLER_23_221 ();
 sg13g2_decap_8 FILLER_23_228 ();
 sg13g2_fill_1 FILLER_23_235 ();
 sg13g2_decap_4 FILLER_23_242 ();
 sg13g2_decap_4 FILLER_23_254 ();
 sg13g2_fill_2 FILLER_23_258 ();
 sg13g2_decap_8 FILLER_23_270 ();
 sg13g2_fill_2 FILLER_23_277 ();
 sg13g2_decap_8 FILLER_23_284 ();
 sg13g2_fill_1 FILLER_23_291 ();
 sg13g2_fill_2 FILLER_23_295 ();
 sg13g2_fill_1 FILLER_23_297 ();
 sg13g2_decap_8 FILLER_23_350 ();
 sg13g2_decap_8 FILLER_23_357 ();
 sg13g2_fill_2 FILLER_23_364 ();
 sg13g2_fill_1 FILLER_23_366 ();
 sg13g2_decap_8 FILLER_23_371 ();
 sg13g2_decap_8 FILLER_23_378 ();
 sg13g2_decap_4 FILLER_23_385 ();
 sg13g2_fill_2 FILLER_23_407 ();
 sg13g2_decap_4 FILLER_24_0 ();
 sg13g2_fill_1 FILLER_24_4 ();
 sg13g2_fill_1 FILLER_24_25 ();
 sg13g2_fill_2 FILLER_24_36 ();
 sg13g2_fill_1 FILLER_24_38 ();
 sg13g2_decap_8 FILLER_24_57 ();
 sg13g2_decap_8 FILLER_24_86 ();
 sg13g2_decap_8 FILLER_24_93 ();
 sg13g2_decap_8 FILLER_24_132 ();
 sg13g2_fill_2 FILLER_24_139 ();
 sg13g2_decap_8 FILLER_24_155 ();
 sg13g2_fill_1 FILLER_24_162 ();
 sg13g2_decap_4 FILLER_24_205 ();
 sg13g2_fill_2 FILLER_24_209 ();
 sg13g2_fill_1 FILLER_24_236 ();
 sg13g2_fill_1 FILLER_24_279 ();
 sg13g2_decap_4 FILLER_24_290 ();
 sg13g2_fill_2 FILLER_24_294 ();
 sg13g2_decap_8 FILLER_24_300 ();
 sg13g2_fill_1 FILLER_24_307 ();
 sg13g2_fill_1 FILLER_24_320 ();
 sg13g2_fill_2 FILLER_24_330 ();
 sg13g2_fill_1 FILLER_24_332 ();
 sg13g2_decap_8 FILLER_24_336 ();
 sg13g2_decap_4 FILLER_24_343 ();
 sg13g2_fill_2 FILLER_24_347 ();
 sg13g2_fill_1 FILLER_24_359 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_4 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_29 ();
 sg13g2_decap_4 FILLER_25_36 ();
 sg13g2_decap_8 FILLER_25_54 ();
 sg13g2_decap_4 FILLER_25_61 ();
 sg13g2_decap_4 FILLER_25_95 ();
 sg13g2_fill_1 FILLER_25_99 ();
 sg13g2_decap_4 FILLER_25_110 ();
 sg13g2_fill_2 FILLER_25_114 ();
 sg13g2_decap_8 FILLER_25_130 ();
 sg13g2_fill_2 FILLER_25_165 ();
 sg13g2_fill_1 FILLER_25_167 ();
 sg13g2_decap_8 FILLER_25_172 ();
 sg13g2_decap_4 FILLER_25_179 ();
 sg13g2_fill_1 FILLER_25_183 ();
 sg13g2_decap_4 FILLER_25_191 ();
 sg13g2_decap_8 FILLER_25_198 ();
 sg13g2_decap_4 FILLER_25_210 ();
 sg13g2_fill_2 FILLER_25_214 ();
 sg13g2_decap_8 FILLER_25_221 ();
 sg13g2_decap_4 FILLER_25_238 ();
 sg13g2_fill_1 FILLER_25_247 ();
 sg13g2_decap_4 FILLER_25_253 ();
 sg13g2_fill_1 FILLER_25_257 ();
 sg13g2_fill_2 FILLER_25_263 ();
 sg13g2_fill_2 FILLER_25_273 ();
 sg13g2_fill_2 FILLER_25_284 ();
 sg13g2_fill_2 FILLER_25_331 ();
 sg13g2_fill_1 FILLER_25_333 ();
 sg13g2_fill_2 FILLER_25_366 ();
 sg13g2_decap_4 FILLER_25_380 ();
 sg13g2_fill_1 FILLER_25_384 ();
 sg13g2_decap_4 FILLER_25_405 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_fill_2 FILLER_26_7 ();
 sg13g2_decap_4 FILLER_26_71 ();
 sg13g2_fill_2 FILLER_26_75 ();
 sg13g2_decap_4 FILLER_26_85 ();
 sg13g2_fill_2 FILLER_26_89 ();
 sg13g2_fill_2 FILLER_26_101 ();
 sg13g2_fill_1 FILLER_26_103 ();
 sg13g2_fill_2 FILLER_26_112 ();
 sg13g2_decap_4 FILLER_26_138 ();
 sg13g2_fill_2 FILLER_26_142 ();
 sg13g2_decap_4 FILLER_26_158 ();
 sg13g2_fill_1 FILLER_26_162 ();
 sg13g2_fill_1 FILLER_26_217 ();
 sg13g2_fill_2 FILLER_26_238 ();
 sg13g2_fill_1 FILLER_26_240 ();
 sg13g2_decap_4 FILLER_26_259 ();
 sg13g2_fill_2 FILLER_26_283 ();
 sg13g2_fill_1 FILLER_26_285 ();
 sg13g2_decap_8 FILLER_26_291 ();
 sg13g2_fill_2 FILLER_26_309 ();
 sg13g2_fill_2 FILLER_26_327 ();
 sg13g2_fill_1 FILLER_26_329 ();
 sg13g2_fill_1 FILLER_26_408 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_fill_1 FILLER_27_7 ();
 sg13g2_decap_4 FILLER_27_27 ();
 sg13g2_fill_2 FILLER_27_31 ();
 sg13g2_fill_2 FILLER_27_43 ();
 sg13g2_fill_2 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_4 FILLER_27_63 ();
 sg13g2_fill_1 FILLER_27_67 ();
 sg13g2_fill_1 FILLER_27_76 ();
 sg13g2_decap_8 FILLER_27_108 ();
 sg13g2_fill_2 FILLER_27_115 ();
 sg13g2_fill_2 FILLER_27_137 ();
 sg13g2_fill_1 FILLER_27_139 ();
 sg13g2_decap_8 FILLER_27_176 ();
 sg13g2_decap_8 FILLER_27_186 ();
 sg13g2_fill_2 FILLER_27_204 ();
 sg13g2_decap_8 FILLER_27_211 ();
 sg13g2_decap_8 FILLER_27_218 ();
 sg13g2_decap_4 FILLER_27_225 ();
 sg13g2_fill_1 FILLER_27_245 ();
 sg13g2_decap_8 FILLER_27_255 ();
 sg13g2_fill_2 FILLER_27_262 ();
 sg13g2_fill_2 FILLER_27_279 ();
 sg13g2_decap_8 FILLER_27_301 ();
 sg13g2_fill_2 FILLER_27_308 ();
 sg13g2_fill_1 FILLER_27_310 ();
 sg13g2_decap_4 FILLER_27_315 ();
 sg13g2_fill_1 FILLER_27_319 ();
 sg13g2_decap_8 FILLER_27_333 ();
 sg13g2_fill_2 FILLER_27_354 ();
 sg13g2_fill_1 FILLER_27_356 ();
 sg13g2_fill_2 FILLER_27_367 ();
 sg13g2_fill_2 FILLER_27_377 ();
 sg13g2_fill_1 FILLER_27_379 ();
 sg13g2_fill_1 FILLER_27_389 ();
 sg13g2_fill_2 FILLER_28_0 ();
 sg13g2_fill_1 FILLER_28_2 ();
 sg13g2_fill_1 FILLER_28_27 ();
 sg13g2_fill_2 FILLER_28_85 ();
 sg13g2_fill_1 FILLER_28_87 ();
 sg13g2_decap_8 FILLER_28_92 ();
 sg13g2_fill_2 FILLER_28_99 ();
 sg13g2_decap_4 FILLER_28_109 ();
 sg13g2_fill_2 FILLER_28_113 ();
 sg13g2_fill_2 FILLER_28_138 ();
 sg13g2_fill_1 FILLER_28_140 ();
 sg13g2_fill_1 FILLER_28_145 ();
 sg13g2_decap_4 FILLER_28_150 ();
 sg13g2_fill_2 FILLER_28_154 ();
 sg13g2_fill_1 FILLER_28_175 ();
 sg13g2_fill_1 FILLER_28_186 ();
 sg13g2_decap_8 FILLER_28_204 ();
 sg13g2_fill_2 FILLER_28_211 ();
 sg13g2_fill_1 FILLER_28_213 ();
 sg13g2_fill_2 FILLER_28_219 ();
 sg13g2_fill_2 FILLER_28_237 ();
 sg13g2_decap_4 FILLER_28_244 ();
 sg13g2_fill_1 FILLER_28_248 ();
 sg13g2_fill_1 FILLER_28_252 ();
 sg13g2_decap_8 FILLER_28_263 ();
 sg13g2_decap_4 FILLER_28_275 ();
 sg13g2_fill_2 FILLER_28_294 ();
 sg13g2_fill_1 FILLER_28_296 ();
 sg13g2_fill_1 FILLER_28_305 ();
 sg13g2_fill_2 FILLER_28_356 ();
 sg13g2_decap_4 FILLER_28_368 ();
 sg13g2_fill_1 FILLER_28_372 ();
 sg13g2_fill_1 FILLER_28_408 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_4 FILLER_29_7 ();
 sg13g2_fill_2 FILLER_29_11 ();
 sg13g2_decap_8 FILLER_29_25 ();
 sg13g2_decap_4 FILLER_29_32 ();
 sg13g2_fill_1 FILLER_29_36 ();
 sg13g2_decap_8 FILLER_29_51 ();
 sg13g2_fill_2 FILLER_29_66 ();
 sg13g2_decap_4 FILLER_29_111 ();
 sg13g2_fill_1 FILLER_29_115 ();
 sg13g2_fill_2 FILLER_29_133 ();
 sg13g2_decap_8 FILLER_29_161 ();
 sg13g2_fill_2 FILLER_29_168 ();
 sg13g2_decap_8 FILLER_29_180 ();
 sg13g2_decap_4 FILLER_29_187 ();
 sg13g2_fill_2 FILLER_29_215 ();
 sg13g2_fill_1 FILLER_29_217 ();
 sg13g2_fill_1 FILLER_29_235 ();
 sg13g2_fill_1 FILLER_29_250 ();
 sg13g2_fill_1 FILLER_29_268 ();
 sg13g2_fill_2 FILLER_29_294 ();
 sg13g2_decap_4 FILLER_29_312 ();
 sg13g2_decap_4 FILLER_29_330 ();
 sg13g2_fill_1 FILLER_29_334 ();
 sg13g2_fill_2 FILLER_29_339 ();
 sg13g2_decap_8 FILLER_29_351 ();
 sg13g2_fill_2 FILLER_29_358 ();
 sg13g2_fill_1 FILLER_29_360 ();
 sg13g2_decap_8 FILLER_29_383 ();
 sg13g2_fill_1 FILLER_29_390 ();
 sg13g2_fill_1 FILLER_29_399 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_fill_1 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_22 ();
 sg13g2_decap_8 FILLER_30_29 ();
 sg13g2_fill_2 FILLER_30_36 ();
 sg13g2_fill_1 FILLER_30_38 ();
 sg13g2_decap_8 FILLER_30_59 ();
 sg13g2_decap_8 FILLER_30_66 ();
 sg13g2_fill_2 FILLER_30_73 ();
 sg13g2_decap_4 FILLER_30_80 ();
 sg13g2_fill_2 FILLER_30_89 ();
 sg13g2_fill_2 FILLER_30_95 ();
 sg13g2_fill_2 FILLER_30_139 ();
 sg13g2_fill_2 FILLER_30_150 ();
 sg13g2_fill_1 FILLER_30_172 ();
 sg13g2_fill_2 FILLER_30_183 ();
 sg13g2_fill_1 FILLER_30_210 ();
 sg13g2_decap_8 FILLER_30_215 ();
 sg13g2_fill_1 FILLER_30_222 ();
 sg13g2_decap_4 FILLER_30_226 ();
 sg13g2_fill_2 FILLER_30_230 ();
 sg13g2_fill_1 FILLER_30_237 ();
 sg13g2_fill_1 FILLER_30_252 ();
 sg13g2_decap_4 FILLER_30_265 ();
 sg13g2_decap_8 FILLER_30_275 ();
 sg13g2_decap_4 FILLER_30_282 ();
 sg13g2_fill_2 FILLER_30_286 ();
 sg13g2_decap_4 FILLER_30_306 ();
 sg13g2_fill_1 FILLER_30_310 ();
 sg13g2_decap_8 FILLER_30_331 ();
 sg13g2_decap_4 FILLER_30_338 ();
 sg13g2_fill_2 FILLER_30_382 ();
 sg13g2_fill_2 FILLER_30_407 ();
 sg13g2_fill_2 FILLER_31_0 ();
 sg13g2_fill_1 FILLER_31_26 ();
 sg13g2_decap_4 FILLER_31_51 ();
 sg13g2_fill_1 FILLER_31_55 ();
 sg13g2_decap_8 FILLER_31_72 ();
 sg13g2_decap_4 FILLER_31_95 ();
 sg13g2_fill_1 FILLER_31_99 ();
 sg13g2_decap_8 FILLER_31_105 ();
 sg13g2_decap_4 FILLER_31_112 ();
 sg13g2_decap_4 FILLER_31_120 ();
 sg13g2_fill_1 FILLER_31_124 ();
 sg13g2_fill_1 FILLER_31_156 ();
 sg13g2_decap_8 FILLER_31_177 ();
 sg13g2_decap_4 FILLER_31_184 ();
 sg13g2_fill_1 FILLER_31_188 ();
 sg13g2_fill_2 FILLER_31_199 ();
 sg13g2_fill_1 FILLER_31_201 ();
 sg13g2_fill_2 FILLER_31_217 ();
 sg13g2_fill_1 FILLER_31_238 ();
 sg13g2_fill_1 FILLER_31_259 ();
 sg13g2_fill_1 FILLER_31_275 ();
 sg13g2_fill_1 FILLER_31_281 ();
 sg13g2_fill_2 FILLER_31_288 ();
 sg13g2_decap_8 FILLER_31_300 ();
 sg13g2_decap_4 FILLER_31_307 ();
 sg13g2_fill_2 FILLER_31_331 ();
 sg13g2_decap_4 FILLER_31_336 ();
 sg13g2_fill_2 FILLER_31_340 ();
 sg13g2_decap_8 FILLER_31_352 ();
 sg13g2_decap_8 FILLER_31_359 ();
 sg13g2_decap_8 FILLER_31_366 ();
 sg13g2_fill_2 FILLER_31_373 ();
 sg13g2_fill_2 FILLER_31_379 ();
 sg13g2_fill_1 FILLER_31_381 ();
 sg13g2_decap_4 FILLER_31_385 ();
 sg13g2_fill_2 FILLER_31_389 ();
 sg13g2_decap_4 FILLER_31_405 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_fill_2 FILLER_32_7 ();
 sg13g2_decap_4 FILLER_32_21 ();
 sg13g2_fill_2 FILLER_32_25 ();
 sg13g2_decap_8 FILLER_32_45 ();
 sg13g2_decap_4 FILLER_32_52 ();
 sg13g2_fill_1 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_79 ();
 sg13g2_fill_2 FILLER_32_86 ();
 sg13g2_decap_4 FILLER_32_114 ();
 sg13g2_fill_1 FILLER_32_118 ();
 sg13g2_decap_4 FILLER_32_136 ();
 sg13g2_fill_2 FILLER_32_145 ();
 sg13g2_decap_8 FILLER_32_157 ();
 sg13g2_fill_2 FILLER_32_164 ();
 sg13g2_fill_1 FILLER_32_166 ();
 sg13g2_decap_8 FILLER_32_184 ();
 sg13g2_decap_8 FILLER_32_207 ();
 sg13g2_fill_2 FILLER_32_214 ();
 sg13g2_fill_1 FILLER_32_216 ();
 sg13g2_decap_4 FILLER_32_227 ();
 sg13g2_fill_1 FILLER_32_231 ();
 sg13g2_decap_8 FILLER_32_257 ();
 sg13g2_fill_2 FILLER_32_274 ();
 sg13g2_decap_4 FILLER_32_287 ();
 sg13g2_decap_8 FILLER_32_306 ();
 sg13g2_decap_8 FILLER_32_313 ();
 sg13g2_fill_2 FILLER_32_330 ();
 sg13g2_decap_8 FILLER_32_352 ();
 sg13g2_decap_4 FILLER_32_359 ();
 sg13g2_fill_1 FILLER_32_408 ();
 sg13g2_fill_2 FILLER_33_24 ();
 sg13g2_fill_2 FILLER_33_38 ();
 sg13g2_fill_1 FILLER_33_40 ();
 sg13g2_decap_8 FILLER_33_91 ();
 sg13g2_fill_1 FILLER_33_98 ();
 sg13g2_decap_4 FILLER_33_103 ();
 sg13g2_fill_2 FILLER_33_115 ();
 sg13g2_fill_1 FILLER_33_117 ();
 sg13g2_decap_4 FILLER_33_128 ();
 sg13g2_decap_4 FILLER_33_160 ();
 sg13g2_fill_2 FILLER_33_164 ();
 sg13g2_decap_4 FILLER_33_190 ();
 sg13g2_fill_2 FILLER_33_234 ();
 sg13g2_fill_1 FILLER_33_240 ();
 sg13g2_decap_4 FILLER_33_255 ();
 sg13g2_fill_1 FILLER_33_259 ();
 sg13g2_decap_4 FILLER_33_272 ();
 sg13g2_fill_1 FILLER_33_276 ();
 sg13g2_decap_8 FILLER_33_282 ();
 sg13g2_decap_8 FILLER_33_289 ();
 sg13g2_fill_2 FILLER_33_296 ();
 sg13g2_fill_1 FILLER_33_342 ();
 sg13g2_fill_1 FILLER_33_391 ();
 sg13g2_fill_1 FILLER_34_0 ();
 sg13g2_fill_2 FILLER_34_15 ();
 sg13g2_fill_1 FILLER_34_27 ();
 sg13g2_fill_2 FILLER_34_38 ();
 sg13g2_fill_1 FILLER_34_40 ();
 sg13g2_decap_4 FILLER_34_51 ();
 sg13g2_fill_2 FILLER_34_55 ();
 sg13g2_decap_8 FILLER_34_71 ();
 sg13g2_decap_8 FILLER_34_102 ();
 sg13g2_decap_4 FILLER_34_109 ();
 sg13g2_fill_2 FILLER_34_113 ();
 sg13g2_decap_4 FILLER_34_125 ();
 sg13g2_fill_2 FILLER_34_129 ();
 sg13g2_fill_2 FILLER_34_166 ();
 sg13g2_fill_1 FILLER_34_168 ();
 sg13g2_fill_2 FILLER_34_189 ();
 sg13g2_fill_2 FILLER_34_209 ();
 sg13g2_fill_1 FILLER_34_211 ();
 sg13g2_fill_2 FILLER_34_229 ();
 sg13g2_fill_1 FILLER_34_269 ();
 sg13g2_fill_1 FILLER_34_275 ();
 sg13g2_decap_8 FILLER_34_291 ();
 sg13g2_fill_1 FILLER_34_298 ();
 sg13g2_decap_8 FILLER_34_307 ();
 sg13g2_fill_1 FILLER_34_314 ();
 sg13g2_fill_1 FILLER_34_327 ();
 sg13g2_fill_2 FILLER_34_353 ();
 sg13g2_fill_2 FILLER_34_368 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_fill_2 FILLER_35_7 ();
 sg13g2_fill_2 FILLER_35_17 ();
 sg13g2_fill_1 FILLER_35_19 ();
 sg13g2_fill_1 FILLER_35_52 ();
 sg13g2_fill_2 FILLER_35_73 ();
 sg13g2_fill_1 FILLER_35_75 ();
 sg13g2_fill_2 FILLER_35_98 ();
 sg13g2_decap_8 FILLER_35_124 ();
 sg13g2_decap_8 FILLER_35_149 ();
 sg13g2_decap_8 FILLER_35_156 ();
 sg13g2_decap_8 FILLER_35_163 ();
 sg13g2_decap_8 FILLER_35_170 ();
 sg13g2_decap_8 FILLER_35_177 ();
 sg13g2_fill_1 FILLER_35_184 ();
 sg13g2_fill_2 FILLER_35_189 ();
 sg13g2_fill_1 FILLER_35_191 ();
 sg13g2_decap_8 FILLER_35_197 ();
 sg13g2_fill_2 FILLER_35_204 ();
 sg13g2_fill_2 FILLER_35_211 ();
 sg13g2_fill_1 FILLER_35_213 ();
 sg13g2_fill_2 FILLER_35_239 ();
 sg13g2_fill_1 FILLER_35_249 ();
 sg13g2_fill_2 FILLER_35_271 ();
 sg13g2_fill_1 FILLER_35_364 ();
 sg13g2_fill_2 FILLER_35_375 ();
 sg13g2_fill_1 FILLER_35_384 ();
 sg13g2_fill_2 FILLER_35_407 ();
 sg13g2_decap_8 FILLER_36_24 ();
 sg13g2_decap_8 FILLER_36_45 ();
 sg13g2_decap_4 FILLER_36_52 ();
 sg13g2_fill_1 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_73 ();
 sg13g2_fill_2 FILLER_36_94 ();
 sg13g2_fill_2 FILLER_36_110 ();
 sg13g2_decap_8 FILLER_36_120 ();
 sg13g2_fill_1 FILLER_36_127 ();
 sg13g2_decap_8 FILLER_36_209 ();
 sg13g2_decap_4 FILLER_36_216 ();
 sg13g2_fill_1 FILLER_36_220 ();
 sg13g2_fill_2 FILLER_36_276 ();
 sg13g2_decap_8 FILLER_36_286 ();
 sg13g2_decap_4 FILLER_36_293 ();
 sg13g2_fill_2 FILLER_36_316 ();
 sg13g2_decap_4 FILLER_36_326 ();
 sg13g2_fill_2 FILLER_36_336 ();
 sg13g2_fill_2 FILLER_36_348 ();
 sg13g2_decap_4 FILLER_37_0 ();
 sg13g2_fill_2 FILLER_37_4 ();
 sg13g2_decap_8 FILLER_37_16 ();
 sg13g2_decap_4 FILLER_37_23 ();
 sg13g2_decap_8 FILLER_37_47 ();
 sg13g2_decap_8 FILLER_37_54 ();
 sg13g2_decap_8 FILLER_37_61 ();
 sg13g2_decap_8 FILLER_37_68 ();
 sg13g2_fill_2 FILLER_37_95 ();
 sg13g2_fill_1 FILLER_37_97 ();
 sg13g2_decap_8 FILLER_37_126 ();
 sg13g2_fill_2 FILLER_37_133 ();
 sg13g2_fill_1 FILLER_37_139 ();
 sg13g2_fill_1 FILLER_37_182 ();
 sg13g2_decap_8 FILLER_37_199 ();
 sg13g2_decap_4 FILLER_37_206 ();
 sg13g2_fill_2 FILLER_37_210 ();
 sg13g2_decap_4 FILLER_37_216 ();
 sg13g2_fill_2 FILLER_37_220 ();
 sg13g2_decap_8 FILLER_37_230 ();
 sg13g2_fill_2 FILLER_37_237 ();
 sg13g2_fill_2 FILLER_37_243 ();
 sg13g2_fill_2 FILLER_37_388 ();
 sg13g2_fill_2 FILLER_37_407 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_4 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_19 ();
 sg13g2_decap_4 FILLER_38_26 ();
 sg13g2_fill_2 FILLER_38_30 ();
 sg13g2_decap_4 FILLER_38_48 ();
 sg13g2_fill_1 FILLER_38_52 ();
 sg13g2_fill_2 FILLER_38_115 ();
 sg13g2_fill_1 FILLER_38_166 ();
 sg13g2_decap_8 FILLER_38_227 ();
 sg13g2_decap_8 FILLER_38_234 ();
 sg13g2_fill_1 FILLER_38_241 ();
 sg13g2_fill_2 FILLER_38_250 ();
 sg13g2_fill_2 FILLER_38_261 ();
 sg13g2_fill_1 FILLER_38_267 ();
 sg13g2_fill_1 FILLER_38_295 ();
 sg13g2_fill_1 FILLER_38_328 ();
 sg13g2_decap_4 FILLER_38_333 ();
 sg13g2_fill_2 FILLER_38_337 ();
 sg13g2_fill_1 FILLER_38_380 ();
 sg13g2_fill_1 FILLER_38_397 ();
 sg13g2_decap_8 FILLER_38_401 ();
 sg13g2_fill_1 FILLER_38_408 ();
 assign uio_oe[0] = net134;
 assign uio_oe[1] = net135;
 assign uio_oe[2] = net136;
 assign uio_oe[3] = net137;
 assign uio_oe[4] = net138;
 assign uio_oe[5] = net139;
 assign uio_oe[6] = net140;
 assign uio_oe[7] = net141;
 assign uio_out[0] = net142;
 assign uio_out[1] = net143;
 assign uio_out[2] = net144;
 assign uio_out[3] = net145;
 assign uio_out[4] = net146;
 assign uio_out[5] = net147;
 assign uio_out[6] = net148;
 assign uio_out[7] = net149;
endmodule

module tt_um_warp (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire _3093_;
 wire _3094_;
 wire _3095_;
 wire _3096_;
 wire _3097_;
 wire _3098_;
 wire _3099_;
 wire _3100_;
 wire _3101_;
 wire _3102_;
 wire _3103_;
 wire _3104_;
 wire _3105_;
 wire _3106_;
 wire _3107_;
 wire _3108_;
 wire _3109_;
 wire _3110_;
 wire _3111_;
 wire _3112_;
 wire _3113_;
 wire _3114_;
 wire _3115_;
 wire _3116_;
 wire _3117_;
 wire _3118_;
 wire _3119_;
 wire _3120_;
 wire _3121_;
 wire _3122_;
 wire _3123_;
 wire _3124_;
 wire _3125_;
 wire _3126_;
 wire _3127_;
 wire _3128_;
 wire _3129_;
 wire _3130_;
 wire _3131_;
 wire _3132_;
 wire _3133_;
 wire _3134_;
 wire _3135_;
 wire _3136_;
 wire _3137_;
 wire _3138_;
 wire _3139_;
 wire _3140_;
 wire _3141_;
 wire _3142_;
 wire _3143_;
 wire _3144_;
 wire _3145_;
 wire _3146_;
 wire _3147_;
 wire _3148_;
 wire _3149_;
 wire _3150_;
 wire _3151_;
 wire _3152_;
 wire _3153_;
 wire _3154_;
 wire _3155_;
 wire _3156_;
 wire _3157_;
 wire _3158_;
 wire _3159_;
 wire _3160_;
 wire _3161_;
 wire _3162_;
 wire _3163_;
 wire _3164_;
 wire _3165_;
 wire _3166_;
 wire _3167_;
 wire _3168_;
 wire _3169_;
 wire _3170_;
 wire _3171_;
 wire _3172_;
 wire _3173_;
 wire _3174_;
 wire _3175_;
 wire _3176_;
 wire _3177_;
 wire _3178_;
 wire _3179_;
 wire _3180_;
 wire _3181_;
 wire _3182_;
 wire _3183_;
 wire _3184_;
 wire _3185_;
 wire _3186_;
 wire _3187_;
 wire _3188_;
 wire _3189_;
 wire _3190_;
 wire _3191_;
 wire _3192_;
 wire _3193_;
 wire _3194_;
 wire _3195_;
 wire _3196_;
 wire _3197_;
 wire _3198_;
 wire _3199_;
 wire _3200_;
 wire _3201_;
 wire _3202_;
 wire _3203_;
 wire _3204_;
 wire _3205_;
 wire _3206_;
 wire _3207_;
 wire _3208_;
 wire _3209_;
 wire _3210_;
 wire _3211_;
 wire _3212_;
 wire _3213_;
 wire _3214_;
 wire _3215_;
 wire _3216_;
 wire _3217_;
 wire _3218_;
 wire _3219_;
 wire _3220_;
 wire _3221_;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire \main._w_demo_audio1 ;
 wire \main._w_demo_video_hs ;
 wire \main._w_demo_video_vs ;
 wire \main.demo._d___pip_58_1_1___stage___block_3_a[1] ;
 wire \main.demo._d___pip_58_1_1___stage___block_3_a[2] ;
 wire \main.demo._d___pip_58_1_1___stage___block_3_a[3] ;
 wire \main.demo._d___pip_58_1_1___stage___block_3_a[4] ;
 wire \main.demo._d___pip_58_1_1___stage___block_3_a[6] ;
 wire \main.demo._d___pip_58_1_1___stage___block_3_a[7] ;
 wire \main.demo._d___pip_58_1_1___stage___block_3_cx[0] ;
 wire \main.demo._d___pip_58_1_1___stage___block_3_cx[10] ;
 wire \main.demo._d___pip_58_1_1___stage___block_3_cx[1] ;
 wire \main.demo._d___pip_58_1_1___stage___block_3_cx[2] ;
 wire \main.demo._d___pip_58_1_1___stage___block_3_cx[3] ;
 wire \main.demo._d___pip_58_1_1___stage___block_3_cx[4] ;
 wire \main.demo._d___pip_58_1_1___stage___block_3_cx[5] ;
 wire \main.demo._d___pip_58_1_1___stage___block_3_cx[6] ;
 wire \main.demo._d___pip_58_1_1___stage___block_3_cx[7] ;
 wire \main.demo._d___pip_58_1_1___stage___block_3_cx[8] ;
 wire \main.demo._d___pip_58_1_1___stage___block_3_cx[9] ;
 wire \main.demo._d___pip_58_1_1___stage___block_3_cy[0] ;
 wire \main.demo._d___pip_58_1_1___stage___block_3_cy[10] ;
 wire \main.demo._d___pip_58_1_1___stage___block_3_cy[1] ;
 wire \main.demo._d___pip_58_1_1___stage___block_3_cy[2] ;
 wire \main.demo._d___pip_58_1_1___stage___block_3_cy[3] ;
 wire \main.demo._d___pip_58_1_1___stage___block_3_cy[4] ;
 wire \main.demo._d___pip_58_1_1___stage___block_3_cy[5] ;
 wire \main.demo._d___pip_58_1_1___stage___block_3_cy[6] ;
 wire \main.demo._d___pip_58_1_1___stage___block_3_cy[7] ;
 wire \main.demo._d___pip_58_1_1___stage___block_3_cy[8] ;
 wire \main.demo._d___pip_58_1_1___stage___block_3_cy[9] ;
 wire \main.demo._d___pip_58_1_2___stage___block_3_a[1] ;
 wire \main.demo._d___pip_58_1_2___stage___block_3_a[2] ;
 wire \main.demo._d___pip_58_1_2___stage___block_3_a[3] ;
 wire \main.demo._d___pip_58_1_2___stage___block_3_a[4] ;
 wire \main.demo._d___pip_58_1_2___stage___block_3_a[5] ;
 wire \main.demo._d___pip_58_1_2___stage___block_3_a[6] ;
 wire \main.demo._d___pip_58_1_2___stage___block_3_a[7] ;
 wire \main.demo._d___pip_58_1_2___stage___block_3_cx[0] ;
 wire \main.demo._d___pip_58_1_2___stage___block_3_cx[10] ;
 wire \main.demo._d___pip_58_1_2___stage___block_3_cx[1] ;
 wire \main.demo._d___pip_58_1_2___stage___block_3_cx[2] ;
 wire \main.demo._d___pip_58_1_2___stage___block_3_cx[3] ;
 wire \main.demo._d___pip_58_1_2___stage___block_3_cx[4] ;
 wire \main.demo._d___pip_58_1_2___stage___block_3_cx[5] ;
 wire \main.demo._d___pip_58_1_2___stage___block_3_cx[6] ;
 wire \main.demo._d___pip_58_1_2___stage___block_3_cx[7] ;
 wire \main.demo._d___pip_58_1_2___stage___block_3_cx[8] ;
 wire \main.demo._d___pip_58_1_2___stage___block_3_cx[9] ;
 wire \main.demo._d___pip_58_1_3___stage___block_3_a[1] ;
 wire \main.demo._d___pip_58_1_3___stage___block_3_a[2] ;
 wire \main.demo._d___pip_58_1_3___stage___block_3_a[3] ;
 wire \main.demo._d___pip_58_1_3___stage___block_3_a[4] ;
 wire \main.demo._d___pip_58_1_3___stage___block_3_a[5] ;
 wire \main.demo._d___pip_58_1_3___stage___block_3_a[6] ;
 wire \main.demo._d___pip_58_1_3___stage___block_3_a[7] ;
 wire \main.demo._d___pip_58_1_3___stage___block_3_cx[0] ;
 wire \main.demo._d___pip_58_1_3___stage___block_3_cx[10] ;
 wire \main.demo._d___pip_58_1_3___stage___block_3_cx[1] ;
 wire \main.demo._d___pip_58_1_3___stage___block_3_cx[2] ;
 wire \main.demo._d___pip_58_1_3___stage___block_3_cx[3] ;
 wire \main.demo._d___pip_58_1_3___stage___block_3_cx[4] ;
 wire \main.demo._d___pip_58_1_3___stage___block_3_cx[5] ;
 wire \main.demo._d___pip_58_1_3___stage___block_3_cx[6] ;
 wire \main.demo._d___pip_58_1_3___stage___block_3_cx[7] ;
 wire \main.demo._d___pip_58_1_3___stage___block_3_cx[8] ;
 wire \main.demo._d___pip_58_1_3___stage___block_3_cx[9] ;
 wire \main.demo._d___pip_58_1_4___block_68_frag[0] ;
 wire \main.demo._d___pip_58_1_4___block_68_frag[1] ;
 wire \main.demo._d___pip_58_1_4___block_68_frag[2] ;
 wire \main.demo._d___pip_58_1_4___block_68_frag[3] ;
 wire \main.demo._d___pip_58_1_4___block_68_frag[4] ;
 wire \main.demo._d___pip_58_1_4___block_68_frag[5] ;
 wire \main.demo._d___pip_58_1_4___block_87_atten_h[0] ;
 wire \main.demo._d___pip_58_1_4___block_87_atten_h[1] ;
 wire \main.demo._d___pip_58_1_4___block_87_atten_h[2] ;
 wire \main.demo._d___pip_58_1_4___block_87_atten_l[0] ;
 wire \main.demo._d___pip_58_1_4___block_87_atten_l[1] ;
 wire \main.demo._d___pip_58_1_4___stage___block_3_cx[1] ;
 wire \main.demo._d___pip_58_1_4___stage___block_3_cx[2] ;
 wire \main.demo._d___pip_58_1_4___stage___block_3_cx[3] ;
 wire \main.demo._d___pip_58_1_4___stage___block_3_cx[4] ;
 wire \main.demo._d___pip_58_1_4___stage___block_3_cx[5] ;
 wire \main.demo._d___pip_58_1_4___stage___block_3_cx[6] ;
 wire \main.demo._d___pip_58_1_4___stage___block_3_cx[9] ;
 wire \main.demo._d_prev_b[0] ;
 wire \main.demo._d_prev_b[1] ;
 wire \main.demo._d_prev_b[2] ;
 wire \main.demo._d_prev_b[3] ;
 wire \main.demo._d_prev_b[4] ;
 wire \main.demo._d_prev_b[5] ;
 wire \main.demo._d_prev_b[6] ;
 wire \main.demo._d_prev_b[7] ;
 wire \main.demo._q___pip_58_1_1___stage___block_3_cx[0] ;
 wire \main.demo._q___pip_58_1_1___stage___block_3_cx[10] ;
 wire \main.demo._q___pip_58_1_1___stage___block_3_cx[1] ;
 wire \main.demo._q___pip_58_1_1___stage___block_3_cx[2] ;
 wire \main.demo._q___pip_58_1_1___stage___block_3_cx[3] ;
 wire \main.demo._q___pip_58_1_1___stage___block_3_cx[4] ;
 wire \main.demo._q___pip_58_1_1___stage___block_3_cx[5] ;
 wire \main.demo._q___pip_58_1_1___stage___block_3_cx[6] ;
 wire \main.demo._q___pip_58_1_1___stage___block_3_cx[7] ;
 wire \main.demo._q___pip_58_1_1___stage___block_3_cx[8] ;
 wire \main.demo._q___pip_58_1_1___stage___block_3_cx[9] ;
 wire \main.demo._q___pip_58_1_1___stage___block_3_cy[0] ;
 wire \main.demo._q___pip_58_1_1___stage___block_3_cy[10] ;
 wire \main.demo._q___pip_58_1_1___stage___block_3_cy[1] ;
 wire \main.demo._q___pip_58_1_1___stage___block_3_cy[2] ;
 wire \main.demo._q___pip_58_1_1___stage___block_3_cy[3] ;
 wire \main.demo._q___pip_58_1_1___stage___block_3_cy[4] ;
 wire \main.demo._q___pip_58_1_1___stage___block_3_cy[5] ;
 wire \main.demo._q___pip_58_1_1___stage___block_3_cy[6] ;
 wire \main.demo._q___pip_58_1_1___stage___block_3_cy[7] ;
 wire \main.demo._q___pip_58_1_1___stage___block_3_cy[8] ;
 wire \main.demo._q___pip_58_1_1___stage___block_3_cy[9] ;
 wire \main.demo._q___pip_58_1_2___stage___block_3_a[1] ;
 wire \main.demo._q___pip_58_1_2___stage___block_3_a[2] ;
 wire \main.demo._q___pip_58_1_2___stage___block_3_a[3] ;
 wire \main.demo._q___pip_58_1_2___stage___block_3_a[4] ;
 wire \main.demo._q___pip_58_1_2___stage___block_3_a[6] ;
 wire \main.demo._q___pip_58_1_2___stage___block_3_a[7] ;
 wire \main.demo._q___pip_58_1_2___stage___block_3_cx[0] ;
 wire \main.demo._q___pip_58_1_2___stage___block_3_cx[10] ;
 wire \main.demo._q___pip_58_1_2___stage___block_3_cx[1] ;
 wire \main.demo._q___pip_58_1_2___stage___block_3_cx[2] ;
 wire \main.demo._q___pip_58_1_2___stage___block_3_cx[3] ;
 wire \main.demo._q___pip_58_1_2___stage___block_3_cx[4] ;
 wire \main.demo._q___pip_58_1_2___stage___block_3_cx[5] ;
 wire \main.demo._q___pip_58_1_2___stage___block_3_cx[6] ;
 wire \main.demo._q___pip_58_1_2___stage___block_3_cx[7] ;
 wire \main.demo._q___pip_58_1_2___stage___block_3_cx[8] ;
 wire \main.demo._q___pip_58_1_2___stage___block_3_cx[9] ;
 wire \main.demo._q___pip_58_1_2___stage___block_3_cy[0] ;
 wire \main.demo._q___pip_58_1_2___stage___block_3_cy[10] ;
 wire \main.demo._q___pip_58_1_2___stage___block_3_cy[1] ;
 wire \main.demo._q___pip_58_1_2___stage___block_3_cy[2] ;
 wire \main.demo._q___pip_58_1_2___stage___block_3_cy[3] ;
 wire \main.demo._q___pip_58_1_2___stage___block_3_cy[4] ;
 wire \main.demo._q___pip_58_1_2___stage___block_3_cy[5] ;
 wire \main.demo._q___pip_58_1_2___stage___block_3_cy[6] ;
 wire \main.demo._q___pip_58_1_2___stage___block_3_cy[7] ;
 wire \main.demo._q___pip_58_1_2___stage___block_3_cy[8] ;
 wire \main.demo._q___pip_58_1_2___stage___block_3_cy[9] ;
 wire \main.demo._q_effect[0] ;
 wire \main.demo._q_effect[1] ;
 wire \main.demo._q_frame[0] ;
 wire \main.demo._q_frame[10] ;
 wire \main.demo._q_frame[11] ;
 wire \main.demo._q_frame[12] ;
 wire \main.demo._q_frame[13] ;
 wire \main.demo._q_frame[14] ;
 wire \main.demo._q_frame[1] ;
 wire \main.demo._q_frame[2] ;
 wire \main.demo._q_frame[3] ;
 wire \main.demo._q_frame[4] ;
 wire \main.demo._q_frame[5] ;
 wire \main.demo._q_frame[6] ;
 wire \main.demo._q_frame[7] ;
 wire \main.demo._q_frame[8] ;
 wire \main.demo._q_frame[9] ;
 wire \main.demo._q_go ;
 wire \main.demo._q_prev_b[6] ;
 wire \main.demo._q_prev_b[7] ;
 wire \main.demo._q_prev_vs ;
 wire \main.demo._q_rot_en ;
 wire \main.demo._q_speed[0] ;
 wire \main.demo._q_speed[10] ;
 wire \main.demo._q_speed[11] ;
 wire \main.demo._q_speed[12] ;
 wire \main.demo._q_speed[13] ;
 wire \main.demo._q_speed[14] ;
 wire \main.demo._q_speed[15] ;
 wire \main.demo._q_speed[1] ;
 wire \main.demo._q_speed[2] ;
 wire \main.demo._q_speed[3] ;
 wire \main.demo._q_speed[4] ;
 wire \main.demo._q_speed[5] ;
 wire \main.demo._q_speed[6] ;
 wire \main.demo._q_speed[7] ;
 wire \main.demo._q_speed[8] ;
 wire \main.demo._q_speed[9] ;
 wire \main.demo._q_th[0] ;
 wire \main.demo._q_th[1] ;
 wire \main.demo._q_th[2] ;
 wire \main.demo._q_th[3] ;
 wire \main.demo._q_th[4] ;
 wire \main.demo._q_th[5] ;
 wire \main.demo._q_th[6] ;
 wire \main.demo._q_th[7] ;
 wire \main.demo._q_th[8] ;
 wire \main.demo._t___block_68_frag[0] ;
 wire \main.demo._t___block_68_frag[1] ;
 wire \main.demo._t___block_68_frag[2] ;
 wire \main.demo._t___block_68_frag[3] ;
 wire \main.demo._t___block_68_frag[4] ;
 wire \main.demo._t___block_68_frag[5] ;
 wire \main.demo._t___pip_58_1_0___stage___block_3_a[6] ;
 wire \main.demo._t___pip_58_1_0___stage___block_3_a[7] ;
 wire \main.demo._t___pip_58_1_0___stage___block_3_cx[0] ;
 wire \main.demo._t___pip_58_1_0___stage___block_3_cx[10] ;
 wire \main.demo._t___pip_58_1_0___stage___block_3_cx[1] ;
 wire \main.demo._t___pip_58_1_0___stage___block_3_cx[2] ;
 wire \main.demo._t___pip_58_1_0___stage___block_3_cx[3] ;
 wire \main.demo._t___pip_58_1_0___stage___block_3_cx[4] ;
 wire \main.demo._t___pip_58_1_0___stage___block_3_cx[5] ;
 wire \main.demo._t___pip_58_1_0___stage___block_3_cx[6] ;
 wire \main.demo._t___pip_58_1_0___stage___block_3_cx[7] ;
 wire \main.demo._t___pip_58_1_0___stage___block_3_cx[8] ;
 wire \main.demo._t___pip_58_1_0___stage___block_3_cx[9] ;
 wire \main.demo._t___pip_58_1_0___stage___block_3_cy[0] ;
 wire \main.demo._t___pip_58_1_0___stage___block_3_cy[10] ;
 wire \main.demo._t___pip_58_1_0___stage___block_3_cy[1] ;
 wire \main.demo._t___pip_58_1_0___stage___block_3_cy[2] ;
 wire \main.demo._t___pip_58_1_0___stage___block_3_cy[3] ;
 wire \main.demo._t___pip_58_1_0___stage___block_3_cy[4] ;
 wire \main.demo._t___pip_58_1_0___stage___block_3_cy[5] ;
 wire \main.demo._t___pip_58_1_0___stage___block_3_cy[6] ;
 wire \main.demo._t___pip_58_1_0___stage___block_3_cy[7] ;
 wire \main.demo._t___pip_58_1_0___stage___block_3_cy[8] ;
 wire \main.demo._t___pip_58_1_0___stage___block_3_cy[9] ;
 wire \main.demo._t___pip_58_1_3___block_87_atten_h[0] ;
 wire \main.demo._t___pip_58_1_3___block_87_atten_h[1] ;
 wire \main.demo._t___pip_58_1_3___block_87_atten_h[2] ;
 wire \main.demo._t___pip_58_1_3___block_87_atten_l[0] ;
 wire \main.demo._t___pip_58_1_3___block_87_atten_l[1] ;
 wire \main.demo._t___stage___block_3_x[0] ;
 wire \main.demo._t___stage___block_3_x[1] ;
 wire \main.demo._t___stage___block_3_x[2] ;
 wire \main.demo._t___stage___block_3_y[0] ;
 wire \main.demo._t___stage___block_3_y[1] ;
 wire \main.demo._t___stage___block_3_y[2] ;
 wire \main.demo._w_vga_active ;
 wire \main.demo._w_vga_vga_x[10] ;
 wire \main.demo._w_vga_vga_x[3] ;
 wire \main.demo._w_vga_vga_x[4] ;
 wire \main.demo._w_vga_vga_x[5] ;
 wire \main.demo._w_vga_vga_x[6] ;
 wire \main.demo._w_vga_vga_x[7] ;
 wire \main.demo._w_vga_vga_x[8] ;
 wire \main.demo._w_vga_vga_x[9] ;
 wire \main.demo._w_vga_vga_y[10] ;
 wire \main.demo._w_vga_vga_y[3] ;
 wire \main.demo._w_vga_vga_y[4] ;
 wire \main.demo._w_vga_vga_y[5] ;
 wire \main.demo._w_vga_vga_y[6] ;
 wire \main.demo._w_vga_vga_y[7] ;
 wire \main.demo._w_vga_vga_y[8] ;
 wire \main.demo.vga._d_active ;
 wire \main.demo.vga._d_vblank ;
 wire \main.demo.vga._q_active_h ;
 wire \main.demo.vga._q_active_v ;
 wire \main.demo.vga._q_xcount[0] ;
 wire \main.demo.vga._q_xcount[10] ;
 wire \main.demo.vga._q_xcount[1] ;
 wire \main.demo.vga._q_xcount[2] ;
 wire \main.demo.vga._q_xcount[3] ;
 wire \main.demo.vga._q_xcount[4] ;
 wire \main.demo.vga._q_xcount[5] ;
 wire \main.demo.vga._q_xcount[6] ;
 wire \main.demo.vga._q_xcount[7] ;
 wire \main.demo.vga._q_xcount[8] ;
 wire \main.demo.vga._q_xcount[9] ;
 wire \main.demo.vga._q_ycount[0] ;
 wire \main.demo.vga._q_ycount[1] ;
 wire \main.demo.vga._q_ycount[2] ;
 wire \main.demo.vga._q_ycount[3] ;
 wire \main.demo.vga._q_ycount[4] ;
 wire \main.demo.vga._q_ycount[5] ;
 wire \main.demo.vga._q_ycount[6] ;
 wire \main.demo.vga._q_ycount[7] ;
 wire \main.demo.vga._q_ycount[8] ;
 wire \main.demo.zic._q_clock_count[0] ;
 wire \main.demo.zic._q_clock_count[1] ;
 wire \main.demo.zic._q_clock_count[2] ;
 wire \main.demo.zic._q_clock_count[3] ;
 wire \main.demo.zic._q_clock_count[4] ;
 wire \main.demo.zic._q_clock_count[5] ;
 wire \main.demo.zic._q_clock_count[6] ;
 wire \main.demo.zic._q_clock_count[7] ;
 wire \main.demo.zic._q_clock_count[8] ;
 wire \main.demo.zic._q_drum_inc[0] ;
 wire \main.demo.zic._q_drum_inc[1] ;
 wire \main.demo.zic._q_drum_inc[2] ;
 wire \main.demo.zic._q_drum_inc[3] ;
 wire \main.demo.zic._q_idx[0] ;
 wire \main.demo.zic._q_idx[1] ;
 wire \main.demo.zic._q_idx[2] ;
 wire \main.demo.zic._q_idx[3] ;
 wire \main.demo.zic._q_idx[4] ;
 wire \main.demo.zic._q_idx[5] ;
 wire \main.demo.zic._q_idx[6] ;
 wire \main.demo.zic._q_qpos[0] ;
 wire \main.demo.zic._q_qpos[10] ;
 wire \main.demo.zic._q_qpos[11] ;
 wire \main.demo.zic._q_qpos[12] ;
 wire \main.demo.zic._q_qpos[1] ;
 wire \main.demo.zic._q_qpos[2] ;
 wire \main.demo.zic._q_qpos[3] ;
 wire \main.demo.zic._q_qpos[4] ;
 wire \main.demo.zic._q_qpos[5] ;
 wire \main.demo.zic._q_qpos[6] ;
 wire \main.demo.zic._q_qpos[7] ;
 wire \main.demo.zic._q_qpos[8] ;
 wire \main.demo.zic._q_qpos[9] ;
 wire \main.demo.zic._q_rythm_count[0] ;
 wire \main.demo.zic._q_rythm_count[10] ;
 wire \main.demo.zic._q_rythm_count[11] ;
 wire \main.demo.zic._q_rythm_count[12] ;
 wire \main.demo.zic._q_rythm_count[1] ;
 wire \main.demo.zic._q_rythm_count[2] ;
 wire \main.demo.zic._q_rythm_count[3] ;
 wire \main.demo.zic._q_rythm_count[4] ;
 wire \main.demo.zic._q_rythm_count[5] ;
 wire \main.demo.zic._q_rythm_count[6] ;
 wire \main.demo.zic._q_rythm_count[7] ;
 wire \main.demo.zic._q_rythm_count[8] ;
 wire \main.demo.zic._q_rythm_count[9] ;
 wire \main.demo.zic._q_squ_env[0] ;
 wire \main.demo.zic._q_squ_env[1] ;
 wire \main.demo.zic._q_squ_env[2] ;
 wire \main.demo.zic._q_squ_env[3] ;
 wire \main.demo.zic._q_squ_env[4] ;
 wire \main.demo.zic._q_squ_env[5] ;
 wire \main.demo.zic._q_tpos[0] ;
 wire \main.demo.zic._q_tpos[10] ;
 wire \main.demo.zic._q_tpos[11] ;
 wire \main.demo.zic._q_tpos[1] ;
 wire \main.demo.zic._q_tpos[2] ;
 wire \main.demo.zic._q_tpos[3] ;
 wire \main.demo.zic._q_tpos[4] ;
 wire \main.demo.zic._q_tpos[5] ;
 wire \main.demo.zic._q_tpos[6] ;
 wire \main.demo.zic._q_tpos[7] ;
 wire \main.demo.zic._q_tpos[8] ;
 wire \main.demo.zic._q_tpos[9] ;
 wire rst_n_q;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire clknet_leaf_0_clk;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net1;
 wire net2;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;

 sg13g2_inv_1 _3483_ (.Y(_2604_),
    .A(net529));
 sg13g2_inv_1 _3484_ (.Y(_2605_),
    .A(net543));
 sg13g2_inv_1 _3485_ (.Y(_2606_),
    .A(net566));
 sg13g2_inv_1 _3486_ (.Y(_2607_),
    .A(\main.demo.zic._q_rythm_count[10] ));
 sg13g2_inv_1 _3487_ (.Y(_2608_),
    .A(net319));
 sg13g2_inv_2 _3488_ (.Y(_2609_),
    .A(\main.demo._q_th[7] ));
 sg13g2_inv_1 _3489_ (.Y(_2610_),
    .A(\main.demo._q_th[6] ));
 sg13g2_inv_2 _3490_ (.Y(_2611_),
    .A(\main.demo._q_th[5] ));
 sg13g2_inv_1 _3491_ (.Y(_2612_),
    .A(\main.demo._q_th[4] ));
 sg13g2_inv_1 _3492_ (.Y(_2613_),
    .A(\main.demo._q_th[3] ));
 sg13g2_inv_1 _3493_ (.Y(_2614_),
    .A(net419));
 sg13g2_inv_2 _3494_ (.Y(_2615_),
    .A(net422));
 sg13g2_inv_1 _3495_ (.Y(_2616_),
    .A(\main.demo.zic._q_qpos[12] ));
 sg13g2_inv_1 _3496_ (.Y(_2617_),
    .A(net310));
 sg13g2_inv_1 _3497_ (.Y(_2618_),
    .A(net410));
 sg13g2_inv_1 _3498_ (.Y(_2619_),
    .A(\main.demo.zic._q_idx[4] ));
 sg13g2_inv_2 _3499_ (.Y(_2620_),
    .A(\main.demo._d___pip_58_1_3___stage___block_3_cx[7] ));
 sg13g2_inv_1 _3500_ (.Y(_2621_),
    .A(net450));
 sg13g2_inv_1 _3501_ (.Y(_2622_),
    .A(_0041_));
 sg13g2_inv_1 _3502_ (.Y(_2623_),
    .A(_0047_));
 sg13g2_inv_1 _3503_ (.Y(_2624_),
    .A(_0048_));
 sg13g2_inv_1 _3504_ (.Y(_2625_),
    .A(_0049_));
 sg13g2_inv_1 _3505_ (.Y(_2626_),
    .A(_0050_));
 sg13g2_inv_1 _3506_ (.Y(_2627_),
    .A(_0051_));
 sg13g2_inv_1 _3507_ (.Y(_2628_),
    .A(\main.demo._q___pip_58_1_1___stage___block_3_cx[5] ));
 sg13g2_inv_1 _3508_ (.Y(_2629_),
    .A(\main.demo._q___pip_58_1_1___stage___block_3_cy[5] ));
 sg13g2_inv_1 _3509_ (.Y(_2630_),
    .A(\main.demo._w_vga_vga_x[9] ));
 sg13g2_inv_2 _3510_ (.Y(_2631_),
    .A(\main.demo._w_vga_vga_x[7] ));
 sg13g2_inv_2 _3511_ (.Y(_2632_),
    .A(net414));
 sg13g2_inv_1 _3512_ (.Y(_2633_),
    .A(\main.demo._w_vga_vga_x[5] ));
 sg13g2_inv_1 _3513_ (.Y(_2634_),
    .A(\main.demo._q_frame[2] ));
 sg13g2_inv_1 _3514_ (.Y(_2635_),
    .A(_0060_));
 sg13g2_inv_1 _3515_ (.Y(_2636_),
    .A(\main.demo._w_vga_vga_y[5] ));
 sg13g2_inv_1 _3516_ (.Y(_2637_),
    .A(net437));
 sg13g2_inv_1 _3517_ (.Y(_2638_),
    .A(\main.demo.zic._q_clock_count[2] ));
 sg13g2_inv_1 _3518_ (.Y(_2639_),
    .A(\main.demo.vga._q_active_h ));
 sg13g2_inv_2 _3519_ (.Y(_2640_),
    .A(\main.demo._t___stage___block_3_y[0] ));
 sg13g2_inv_1 _3520_ (.Y(_2641_),
    .A(\main.demo._t___stage___block_3_y[1] ));
 sg13g2_inv_1 _3521_ (.Y(_2642_),
    .A(\main.demo._t___stage___block_3_x[1] ));
 sg13g2_inv_1 _3522_ (.Y(_2643_),
    .A(\main.demo._t___stage___block_3_y[2] ));
 sg13g2_inv_2 _3523_ (.Y(_2644_),
    .A(\main.demo._t___stage___block_3_x[2] ));
 sg13g2_inv_1 _3524_ (.Y(_2645_),
    .A(_0005_));
 sg13g2_inv_2 _3525_ (.Y(_2646_),
    .A(net426));
 sg13g2_inv_1 _3526_ (.Y(_2647_),
    .A(\main.demo._q_frame[13] ));
 sg13g2_inv_2 _3527_ (.Y(_2648_),
    .A(net641));
 sg13g2_inv_1 _3528_ (.Y(_2649_),
    .A(net610));
 sg13g2_inv_1 _3529_ (.Y(_2650_),
    .A(\main.demo._d___pip_58_1_3___stage___block_3_cx[6] ));
 sg13g2_inv_2 _3530_ (.Y(_2651_),
    .A(_0008_));
 sg13g2_inv_2 _3531_ (.Y(_2652_),
    .A(_0009_));
 sg13g2_inv_1 _3532_ (.Y(_2653_),
    .A(_0010_));
 sg13g2_inv_1 _3533_ (.Y(_2654_),
    .A(_0012_));
 sg13g2_inv_1 _3534_ (.Y(_2655_),
    .A(_0015_));
 sg13g2_inv_1 _3535_ (.Y(_2656_),
    .A(\main.demo._d___pip_58_1_3___stage___block_3_a[1] ));
 sg13g2_inv_1 _3536_ (.Y(_2657_),
    .A(_0017_));
 sg13g2_inv_1 _3537_ (.Y(_2658_),
    .A(_0019_));
 sg13g2_inv_1 _3538_ (.Y(_2659_),
    .A(_0020_));
 sg13g2_inv_1 _3539_ (.Y(_2660_),
    .A(_0021_));
 sg13g2_inv_1 _3540_ (.Y(_2661_),
    .A(_0023_));
 sg13g2_inv_1 _3541_ (.Y(_2662_),
    .A(net612));
 sg13g2_inv_1 _3542_ (.Y(_2663_),
    .A(net607));
 sg13g2_inv_1 _3543_ (.Y(_2664_),
    .A(net567));
 sg13g2_inv_1 _3544_ (.Y(_2665_),
    .A(net550));
 sg13g2_inv_1 _3545_ (.Y(_2666_),
    .A(_0028_));
 sg13g2_inv_1 _3546_ (.Y(_2667_),
    .A(_0031_));
 sg13g2_inv_1 _3547_ (.Y(_2668_),
    .A(\main.demo._q___pip_58_1_2___stage___block_3_a[4] ));
 sg13g2_inv_1 _3548_ (.Y(_2669_),
    .A(\main.demo._d___pip_58_1_4___block_68_frag[3] ));
 sg13g2_inv_1 _3549_ (.Y(_2670_),
    .A(\main.demo._d___pip_58_1_4___stage___block_3_cx[6] ));
 sg13g2_inv_1 _3550_ (.Y(_2671_),
    .A(\main.demo._d___pip_58_1_4___stage___block_3_cx[5] ));
 sg13g2_inv_1 _3551_ (.Y(_2672_),
    .A(\main.demo._d___pip_58_1_4___stage___block_3_cx[3] ));
 sg13g2_inv_1 _3552_ (.Y(_2673_),
    .A(net284));
 sg13g2_nor2_1 _3553_ (.A(\main.demo._d___pip_58_1_3___stage___block_3_cx[10] ),
    .B(net425),
    .Y(_2674_));
 sg13g2_or2_1 _3554_ (.X(_2675_),
    .B(net425),
    .A(\main.demo._d___pip_58_1_3___stage___block_3_cx[10] ));
 sg13g2_nand2_2 _3555_ (.Y(\main.demo._t___pip_58_1_3___block_87_atten_l[0] ),
    .A(net556),
    .B(net399));
 sg13g2_inv_1 _3556_ (.Y(\main.demo._t___pip_58_1_3___block_87_atten_h[0] ),
    .A(\main.demo._t___pip_58_1_3___block_87_atten_l[0] ));
 sg13g2_nor2b_1 _3557_ (.A(\main.demo._q___pip_58_1_2___stage___block_3_cx[0] ),
    .B_N(\main.demo._q___pip_58_1_2___stage___block_3_cy[3] ),
    .Y(_2676_));
 sg13g2_xor2_1 _3558_ (.B(\main.demo._q___pip_58_1_2___stage___block_3_cy[3] ),
    .A(\main.demo._q___pip_58_1_2___stage___block_3_cx[0] ),
    .X(_2677_));
 sg13g2_nor3_2 _3559_ (.A(\main.demo._q___pip_58_1_2___stage___block_3_cx[5] ),
    .B(\main.demo._q___pip_58_1_2___stage___block_3_cx[3] ),
    .C(\main.demo._q___pip_58_1_2___stage___block_3_cx[4] ),
    .Y(_2678_));
 sg13g2_nand2b_1 _3560_ (.Y(_2679_),
    .B(\main.demo._q___pip_58_1_2___stage___block_3_cx[6] ),
    .A_N(_2678_));
 sg13g2_nand2b_1 _3561_ (.Y(_2680_),
    .B(_2678_),
    .A_N(\main.demo._q___pip_58_1_2___stage___block_3_cx[6] ));
 sg13g2_nand3_1 _3562_ (.B(_2679_),
    .C(_2680_),
    .A(net404),
    .Y(_2681_));
 sg13g2_o21ai_1 _3563_ (.B1(_2681_),
    .Y(_2682_),
    .A1(net404),
    .A2(_0040_));
 sg13g2_nand2b_1 _3564_ (.Y(_2683_),
    .B(_2682_),
    .A_N(_0039_));
 sg13g2_o21ai_1 _3565_ (.B1(\main.demo._q___pip_58_1_2___stage___block_3_cx[5] ),
    .Y(_2684_),
    .A1(\main.demo._q___pip_58_1_2___stage___block_3_cx[3] ),
    .A2(\main.demo._q___pip_58_1_2___stage___block_3_cx[4] ));
 sg13g2_nor2_1 _3566_ (.A(net448),
    .B(_2678_),
    .Y(_2685_));
 sg13g2_a22oi_1 _3567_ (.Y(_2686_),
    .B1(_2684_),
    .B2(_2685_),
    .A2(_2622_),
    .A1(net448));
 sg13g2_nor2b_1 _3568_ (.A(_2686_),
    .B_N(\main.demo._q___pip_58_1_2___stage___block_3_cy[2] ),
    .Y(_2687_));
 sg13g2_xnor2_1 _3569_ (.Y(_2688_),
    .A(\main.demo._q___pip_58_1_2___stage___block_3_cx[3] ),
    .B(\main.demo._q___pip_58_1_2___stage___block_3_cx[4] ));
 sg13g2_mux2_1 _3570_ (.A0(_0042_),
    .A1(_2688_),
    .S(net404),
    .X(_2689_));
 sg13g2_nand2b_1 _3571_ (.Y(_2690_),
    .B(\main.demo._q___pip_58_1_2___stage___block_3_cy[1] ),
    .A_N(_2689_));
 sg13g2_nand2_1 _3572_ (.Y(_2691_),
    .A(\main.demo._q___pip_58_1_2___stage___block_3_cx[3] ),
    .B(\main.demo._q___pip_58_1_2___stage___block_3_cy[0] ));
 sg13g2_xor2_1 _3573_ (.B(_2689_),
    .A(\main.demo._q___pip_58_1_2___stage___block_3_cy[1] ),
    .X(_2692_));
 sg13g2_nor2_1 _3574_ (.A(_2691_),
    .B(_2692_),
    .Y(_2693_));
 sg13g2_o21ai_1 _3575_ (.B1(_2690_),
    .Y(_2694_),
    .A1(_2691_),
    .A2(_2692_));
 sg13g2_xnor2_1 _3576_ (.Y(_2695_),
    .A(\main.demo._q___pip_58_1_2___stage___block_3_cy[2] ),
    .B(_2686_));
 sg13g2_a21oi_2 _3577_ (.B1(_2687_),
    .Y(_2696_),
    .A2(_2695_),
    .A1(_2694_));
 sg13g2_xor2_1 _3578_ (.B(_2682_),
    .A(_0039_),
    .X(_2697_));
 sg13g2_o21ai_1 _3579_ (.B1(_2683_),
    .Y(_2698_),
    .A1(_2696_),
    .A2(_2697_));
 sg13g2_nand2_1 _3580_ (.Y(_2699_),
    .A(\main.demo._q___pip_58_1_2___stage___block_3_cx[7] ),
    .B(_2680_));
 sg13g2_or2_1 _3581_ (.X(_2700_),
    .B(_2680_),
    .A(\main.demo._q___pip_58_1_2___stage___block_3_cx[7] ));
 sg13g2_a21oi_1 _3582_ (.A1(_2699_),
    .A2(_2700_),
    .Y(_2701_),
    .B1(net447));
 sg13g2_a21oi_1 _3583_ (.A1(_0038_),
    .A2(net447),
    .Y(_2702_),
    .B1(_2701_));
 sg13g2_xor2_1 _3584_ (.B(_2702_),
    .A(\main.demo._q___pip_58_1_2___stage___block_3_cy[4] ),
    .X(_2703_));
 sg13g2_xnor2_1 _3585_ (.Y(_2704_),
    .A(_2698_),
    .B(_2703_));
 sg13g2_nor2_1 _3586_ (.A(_2677_),
    .B(_2704_),
    .Y(_2705_));
 sg13g2_inv_1 _3587_ (.Y(_2706_),
    .A(_2705_));
 sg13g2_xnor2_1 _3588_ (.Y(_2707_),
    .A(_2677_),
    .B(_2704_));
 sg13g2_a22oi_1 _3589_ (.Y(_2708_),
    .B1(_2703_),
    .B2(_2698_),
    .A2(_2702_),
    .A1(_2627_));
 sg13g2_inv_1 _3590_ (.Y(_2709_),
    .A(_2708_));
 sg13g2_a21oi_1 _3591_ (.A1(\main.demo._q___pip_58_1_2___stage___block_3_cx[8] ),
    .A2(_2700_),
    .Y(_2710_),
    .B1(net445));
 sg13g2_o21ai_1 _3592_ (.B1(_2710_),
    .Y(_2711_),
    .A1(\main.demo._q___pip_58_1_2___stage___block_3_cx[8] ),
    .A2(_2700_));
 sg13g2_o21ai_1 _3593_ (.B1(_2711_),
    .Y(_2712_),
    .A1(net404),
    .A2(_0045_));
 sg13g2_xor2_1 _3594_ (.B(_2712_),
    .A(\main.demo._q___pip_58_1_2___stage___block_3_cy[5] ),
    .X(_2713_));
 sg13g2_xor2_1 _3595_ (.B(_2713_),
    .A(_2708_),
    .X(_2714_));
 sg13g2_nor2_1 _3596_ (.A(\main.demo._q___pip_58_1_2___stage___block_3_cy[3] ),
    .B(\main.demo._q___pip_58_1_2___stage___block_3_cy[4] ),
    .Y(_2715_));
 sg13g2_nor3_1 _3597_ (.A(\main.demo._q___pip_58_1_2___stage___block_3_cy[3] ),
    .B(\main.demo._q___pip_58_1_2___stage___block_3_cy[4] ),
    .C(\main.demo._q___pip_58_1_2___stage___block_3_cy[5] ),
    .Y(_2716_));
 sg13g2_nor2b_1 _3598_ (.A(\main.demo._q___pip_58_1_2___stage___block_3_cy[6] ),
    .B_N(_2716_),
    .Y(_2717_));
 sg13g2_nand2b_1 _3599_ (.Y(_2718_),
    .B(_2717_),
    .A_N(\main.demo._q___pip_58_1_2___stage___block_3_cy[7] ));
 sg13g2_nand2_1 _3600_ (.Y(_2719_),
    .A(\main.demo._q___pip_58_1_2___stage___block_3_cy[8] ),
    .B(_2718_));
 sg13g2_nor2_2 _3601_ (.A(\main.demo._q___pip_58_1_2___stage___block_3_cy[8] ),
    .B(_2718_),
    .Y(_2720_));
 sg13g2_nor2_1 _3602_ (.A(net446),
    .B(_2720_),
    .Y(_2721_));
 sg13g2_a22oi_1 _3603_ (.Y(_2722_),
    .B1(_2719_),
    .B2(_2721_),
    .A2(_2623_),
    .A1(net446));
 sg13g2_nand2b_1 _3604_ (.Y(_2723_),
    .B(\main.demo._q___pip_58_1_2___stage___block_3_cy[7] ),
    .A_N(_2717_));
 sg13g2_and2_1 _3605_ (.A(net404),
    .B(_2718_),
    .X(_2724_));
 sg13g2_a22oi_1 _3606_ (.Y(_2725_),
    .B1(_2723_),
    .B2(_2724_),
    .A2(_2624_),
    .A1(net445));
 sg13g2_and2_1 _3607_ (.A(\main.demo._q___pip_58_1_2___stage___block_3_cx[4] ),
    .B(_2725_),
    .X(_2726_));
 sg13g2_nand2b_1 _3608_ (.Y(_2727_),
    .B(\main.demo._q___pip_58_1_2___stage___block_3_cy[6] ),
    .A_N(_2716_));
 sg13g2_nor2_1 _3609_ (.A(net447),
    .B(_2717_),
    .Y(_2728_));
 sg13g2_a22oi_1 _3610_ (.Y(_2729_),
    .B1(_2727_),
    .B2(_2728_),
    .A2(_2625_),
    .A1(net447));
 sg13g2_o21ai_1 _3611_ (.B1(\main.demo._q___pip_58_1_2___stage___block_3_cy[5] ),
    .Y(_2730_),
    .A1(\main.demo._q___pip_58_1_2___stage___block_3_cy[3] ),
    .A2(\main.demo._q___pip_58_1_2___stage___block_3_cy[4] ));
 sg13g2_nor2_1 _3612_ (.A(net447),
    .B(_2716_),
    .Y(_2731_));
 sg13g2_a22oi_1 _3613_ (.Y(_2732_),
    .B1(_2730_),
    .B2(_2731_),
    .A2(_2626_),
    .A1(net447));
 sg13g2_nand2_1 _3614_ (.Y(_2733_),
    .A(\main.demo._q___pip_58_1_2___stage___block_3_cy[3] ),
    .B(\main.demo._q___pip_58_1_2___stage___block_3_cy[4] ));
 sg13g2_nor2_1 _3615_ (.A(net448),
    .B(_2715_),
    .Y(_2734_));
 sg13g2_a22oi_1 _3616_ (.Y(_2735_),
    .B1(_2733_),
    .B2(_2734_),
    .A2(_2627_),
    .A1(net448));
 sg13g2_nand2_1 _3617_ (.Y(_2736_),
    .A(\main.demo._q___pip_58_1_2___stage___block_3_cx[1] ),
    .B(_2735_));
 sg13g2_xnor2_1 _3618_ (.Y(_2737_),
    .A(\main.demo._q___pip_58_1_2___stage___block_3_cx[1] ),
    .B(_2735_));
 sg13g2_o21ai_1 _3619_ (.B1(_2736_),
    .Y(_2738_),
    .A1(_2676_),
    .A2(_2737_));
 sg13g2_xnor2_1 _3620_ (.Y(_2739_),
    .A(\main.demo._q___pip_58_1_2___stage___block_3_cx[2] ),
    .B(_2732_));
 sg13g2_nor2b_1 _3621_ (.A(_2739_),
    .B_N(_2738_),
    .Y(_2740_));
 sg13g2_a21o_1 _3622_ (.A2(_2732_),
    .A1(\main.demo._q___pip_58_1_2___stage___block_3_cx[2] ),
    .B1(_2740_),
    .X(_2741_));
 sg13g2_xnor2_1 _3623_ (.Y(_2742_),
    .A(\main.demo._q___pip_58_1_2___stage___block_3_cx[3] ),
    .B(_2729_));
 sg13g2_nor2b_1 _3624_ (.A(_2742_),
    .B_N(_2741_),
    .Y(_2743_));
 sg13g2_a21o_1 _3625_ (.A2(_2729_),
    .A1(\main.demo._q___pip_58_1_2___stage___block_3_cx[3] ),
    .B1(_2743_),
    .X(_2744_));
 sg13g2_xnor2_1 _3626_ (.Y(_2745_),
    .A(_0042_),
    .B(_2725_));
 sg13g2_a21o_1 _3627_ (.A2(_2745_),
    .A1(_2744_),
    .B1(_2726_),
    .X(_2746_));
 sg13g2_xnor2_1 _3628_ (.Y(_2747_),
    .A(_0041_),
    .B(_2722_));
 sg13g2_a22oi_1 _3629_ (.Y(_2748_),
    .B1(_2746_),
    .B2(_2747_),
    .A2(_2722_),
    .A1(\main.demo._q___pip_58_1_2___stage___block_3_cx[5] ));
 sg13g2_xnor2_1 _3630_ (.Y(_2749_),
    .A(\main.demo._q___pip_58_1_2___stage___block_3_cy[9] ),
    .B(_2720_));
 sg13g2_nand2_1 _3631_ (.Y(_2750_),
    .A(net445),
    .B(_0046_));
 sg13g2_o21ai_1 _3632_ (.B1(_2750_),
    .Y(_2751_),
    .A1(net446),
    .A2(_2749_));
 sg13g2_xnor2_1 _3633_ (.Y(_2752_),
    .A(_0040_),
    .B(_2751_));
 sg13g2_nor2b_1 _3634_ (.A(_2748_),
    .B_N(_2752_),
    .Y(_2753_));
 sg13g2_a21o_1 _3635_ (.A2(_2751_),
    .A1(\main.demo._q___pip_58_1_2___stage___block_3_cx[6] ),
    .B1(_2753_),
    .X(_2754_));
 sg13g2_nand2_1 _3636_ (.Y(_2755_),
    .A(_0044_),
    .B(_2720_));
 sg13g2_nand3_1 _3637_ (.B(_0046_),
    .C(_2720_),
    .A(_0044_),
    .Y(_2756_));
 sg13g2_xor2_1 _3638_ (.B(_2756_),
    .A(_0038_),
    .X(_2757_));
 sg13g2_nand2_1 _3639_ (.Y(_2758_),
    .A(_2754_),
    .B(_2757_));
 sg13g2_nand4_1 _3640_ (.B(_0044_),
    .C(_0046_),
    .A(\main.demo._q___pip_58_1_2___stage___block_3_cx[7] ),
    .Y(_2759_),
    .D(_2720_));
 sg13g2_nor3_2 _3641_ (.A(net445),
    .B(\main.demo._q___pip_58_1_2___stage___block_3_cy[9] ),
    .C(_2755_),
    .Y(_2760_));
 sg13g2_inv_1 _3642_ (.Y(_2761_),
    .A(_2760_));
 sg13g2_xor2_1 _3643_ (.B(_2760_),
    .A(_0045_),
    .X(_2762_));
 sg13g2_a21oi_1 _3644_ (.A1(_2758_),
    .A2(_2759_),
    .Y(_2763_),
    .B1(_2762_));
 sg13g2_a21oi_1 _3645_ (.A1(\main.demo._q___pip_58_1_2___stage___block_3_cx[8] ),
    .A2(_2760_),
    .Y(_2764_),
    .B1(_2763_));
 sg13g2_xor2_1 _3646_ (.B(_2760_),
    .A(_0043_),
    .X(_2765_));
 sg13g2_nor2_1 _3647_ (.A(_2764_),
    .B(_2765_),
    .Y(_2766_));
 sg13g2_xor2_1 _3648_ (.B(_2765_),
    .A(_2764_),
    .X(_2767_));
 sg13g2_xnor2_1 _3649_ (.Y(_2768_),
    .A(_2748_),
    .B(_2752_));
 sg13g2_xor2_1 _3650_ (.B(_2747_),
    .A(_2746_),
    .X(_2769_));
 sg13g2_xnor2_1 _3651_ (.Y(_2770_),
    .A(_2744_),
    .B(_2745_));
 sg13g2_inv_1 _3652_ (.Y(_2771_),
    .A(_2770_));
 sg13g2_nor2_1 _3653_ (.A(_2769_),
    .B(_2771_),
    .Y(_2772_));
 sg13g2_nand2b_1 _3654_ (.Y(_2773_),
    .B(_2772_),
    .A_N(_2768_));
 sg13g2_xor2_1 _3655_ (.B(_2757_),
    .A(_2754_),
    .X(_2774_));
 sg13g2_nor2_1 _3656_ (.A(_2773_),
    .B(_2774_),
    .Y(_2775_));
 sg13g2_nand3_1 _3657_ (.B(_2759_),
    .C(_2762_),
    .A(_2758_),
    .Y(_2776_));
 sg13g2_nand2b_2 _3658_ (.Y(_2777_),
    .B(_2776_),
    .A_N(_2763_));
 sg13g2_nand2_1 _3659_ (.Y(_2778_),
    .A(_2775_),
    .B(_2777_));
 sg13g2_or3_1 _3660_ (.A(\main.demo._q___pip_58_1_2___stage___block_3_cx[9] ),
    .B(\main.demo._q___pip_58_1_2___stage___block_3_cx[8] ),
    .C(_2700_),
    .X(_2779_));
 sg13g2_nor2_1 _3661_ (.A(net445),
    .B(_2779_),
    .Y(_2780_));
 sg13g2_nor2_1 _3662_ (.A(\main.demo._q___pip_58_1_2___stage___block_3_cx[10] ),
    .B(_2780_),
    .Y(_2781_));
 sg13g2_nand2_1 _3663_ (.Y(_2782_),
    .A(net404),
    .B(\main.demo._q___pip_58_1_2___stage___block_3_cx[10] ));
 sg13g2_a21oi_1 _3664_ (.A1(net445),
    .A2(_0052_),
    .Y(_2783_),
    .B1(_2780_));
 sg13g2_nand2_2 _3665_ (.Y(_2784_),
    .A(_2782_),
    .B(_2783_));
 sg13g2_o21ai_1 _3666_ (.B1(_2784_),
    .Y(_2785_),
    .A1(_2779_),
    .A2(_2782_));
 sg13g2_o21ai_1 _3667_ (.B1(\main.demo._q___pip_58_1_2___stage___block_3_cx[9] ),
    .Y(_2786_),
    .A1(\main.demo._q___pip_58_1_2___stage___block_3_cx[8] ),
    .A2(_2700_));
 sg13g2_a21oi_1 _3668_ (.A1(_2779_),
    .A2(_2786_),
    .Y(_2787_),
    .B1(net445));
 sg13g2_a21oi_1 _3669_ (.A1(net445),
    .A2(_0043_),
    .Y(_2788_),
    .B1(_2787_));
 sg13g2_a22oi_1 _3670_ (.Y(_2789_),
    .B1(_2713_),
    .B2(_2709_),
    .A2(_2712_),
    .A1(_2626_));
 sg13g2_inv_1 _3671_ (.Y(_2790_),
    .A(_2789_));
 sg13g2_xor2_1 _3672_ (.B(_2788_),
    .A(\main.demo._q___pip_58_1_2___stage___block_3_cy[6] ),
    .X(_2791_));
 sg13g2_a22oi_1 _3673_ (.Y(_2792_),
    .B1(_2790_),
    .B2(_2791_),
    .A2(_2788_),
    .A1(_2625_));
 sg13g2_inv_1 _3674_ (.Y(_2793_),
    .A(_2792_));
 sg13g2_xor2_1 _3675_ (.B(_2785_),
    .A(\main.demo._q___pip_58_1_2___stage___block_3_cy[7] ),
    .X(_2794_));
 sg13g2_a22oi_1 _3676_ (.Y(_2795_),
    .B1(_2793_),
    .B2(_2794_),
    .A2(_2785_),
    .A1(_2624_));
 sg13g2_xor2_1 _3677_ (.B(_2784_),
    .A(\main.demo._q___pip_58_1_2___stage___block_3_cy[8] ),
    .X(_2796_));
 sg13g2_or2_1 _3678_ (.X(_2797_),
    .B(_2796_),
    .A(_2795_));
 sg13g2_xor2_1 _3679_ (.B(_2784_),
    .A(\main.demo._q___pip_58_1_2___stage___block_3_cy[9] ),
    .X(_2798_));
 sg13g2_o21ai_1 _3680_ (.B1(_0046_),
    .Y(_2799_),
    .A1(\main.demo._q___pip_58_1_2___stage___block_3_cy[9] ),
    .A2(_0047_));
 sg13g2_nand3_1 _3681_ (.B(_2783_),
    .C(_2799_),
    .A(_2782_),
    .Y(_2800_));
 sg13g2_o21ai_1 _3682_ (.B1(_2800_),
    .Y(_2801_),
    .A1(_2797_),
    .A2(_2798_));
 sg13g2_xor2_1 _3683_ (.B(_2801_),
    .A(_2781_),
    .X(_2802_));
 sg13g2_xnor2_1 _3684_ (.Y(_2803_),
    .A(_2781_),
    .B(_2801_));
 sg13g2_nand2_1 _3685_ (.Y(_2804_),
    .A(_2778_),
    .B(net349));
 sg13g2_xor2_1 _3686_ (.B(_2804_),
    .A(_2767_),
    .X(_2805_));
 sg13g2_nor2_1 _3687_ (.A(_2714_),
    .B(_2805_),
    .Y(_2806_));
 sg13g2_nand2_1 _3688_ (.Y(_2807_),
    .A(_2714_),
    .B(_2805_));
 sg13g2_nand2b_1 _3689_ (.Y(_2808_),
    .B(_2807_),
    .A_N(_2806_));
 sg13g2_nor2_1 _3690_ (.A(_2775_),
    .B(net351),
    .Y(_2809_));
 sg13g2_xnor2_1 _3691_ (.Y(_2810_),
    .A(_2777_),
    .B(_2809_));
 sg13g2_inv_1 _3692_ (.Y(_2811_),
    .A(_2810_));
 sg13g2_o21ai_1 _3693_ (.B1(_2771_),
    .Y(_2812_),
    .A1(\main.demo._q___pip_58_1_2___stage___block_3_cx[3] ),
    .A2(\main.demo._q___pip_58_1_2___stage___block_3_cy[0] ));
 sg13g2_nor2_1 _3694_ (.A(_2692_),
    .B(_2812_),
    .Y(_2813_));
 sg13g2_nand2_1 _3695_ (.Y(_2814_),
    .A(_2691_),
    .B(_2813_));
 sg13g2_nor2_1 _3696_ (.A(_2770_),
    .B(net352),
    .Y(_2815_));
 sg13g2_and2_1 _3697_ (.A(_2691_),
    .B(_2692_),
    .X(_2816_));
 sg13g2_a221oi_1 _3698_ (.B2(_2812_),
    .C1(_2693_),
    .B1(_2816_),
    .A1(_2769_),
    .Y(_2817_),
    .A2(_2815_));
 sg13g2_o21ai_1 _3699_ (.B1(_2817_),
    .Y(_2818_),
    .A1(_2769_),
    .A2(_2815_));
 sg13g2_xnor2_1 _3700_ (.Y(_2819_),
    .A(_2694_),
    .B(_2695_));
 sg13g2_nor2_1 _3701_ (.A(_2772_),
    .B(net351),
    .Y(_2820_));
 sg13g2_xnor2_1 _3702_ (.Y(_2821_),
    .A(_2768_),
    .B(_2820_));
 sg13g2_a22oi_1 _3703_ (.Y(_2822_),
    .B1(_2819_),
    .B2(_2821_),
    .A2(_2818_),
    .A1(_2814_));
 sg13g2_xnor2_1 _3704_ (.Y(_2823_),
    .A(_2696_),
    .B(_2697_));
 sg13g2_nand2_1 _3705_ (.Y(_2824_),
    .A(_2773_),
    .B(net349));
 sg13g2_xor2_1 _3706_ (.B(_2824_),
    .A(_2774_),
    .X(_2825_));
 sg13g2_or2_1 _3707_ (.X(_2826_),
    .B(_2825_),
    .A(_2823_));
 sg13g2_o21ai_1 _3708_ (.B1(_2826_),
    .Y(_2827_),
    .A1(_2819_),
    .A2(_2821_));
 sg13g2_a22oi_1 _3709_ (.Y(_2828_),
    .B1(_2823_),
    .B2(_2825_),
    .A2(_2811_),
    .A1(_2704_));
 sg13g2_o21ai_1 _3710_ (.B1(_2828_),
    .Y(_2829_),
    .A1(_2822_),
    .A2(_2827_));
 sg13g2_o21ai_1 _3711_ (.B1(_2829_),
    .Y(_2830_),
    .A1(_2704_),
    .A2(_2811_));
 sg13g2_xnor2_1 _3712_ (.Y(_2831_),
    .A(_2808_),
    .B(_2830_));
 sg13g2_nor2b_1 _3713_ (.A(_2707_),
    .B_N(_2831_),
    .Y(_2832_));
 sg13g2_xor2_1 _3714_ (.B(_2831_),
    .A(_2707_),
    .X(\main.demo._d___pip_58_1_2___stage___block_3_cx[0] ));
 sg13g2_nand2b_1 _3715_ (.Y(_2833_),
    .B(\main.demo._q___pip_58_1_1___stage___block_3_cy[9] ),
    .A_N(\main.demo._q___pip_58_1_1___stage___block_3_cx[9] ));
 sg13g2_nor2b_1 _3716_ (.A(\main.demo._q___pip_58_1_1___stage___block_3_cy[9] ),
    .B_N(\main.demo._q___pip_58_1_1___stage___block_3_cx[9] ),
    .Y(_2834_));
 sg13g2_nor2b_1 _3717_ (.A(\main.demo._q___pip_58_1_1___stage___block_3_cy[8] ),
    .B_N(\main.demo._q___pip_58_1_1___stage___block_3_cx[8] ),
    .Y(_2835_));
 sg13g2_nand2b_1 _3718_ (.Y(_2836_),
    .B(\main.demo._q___pip_58_1_1___stage___block_3_cy[8] ),
    .A_N(\main.demo._q___pip_58_1_1___stage___block_3_cx[8] ));
 sg13g2_nor2b_2 _3719_ (.A(_2835_),
    .B_N(_2836_),
    .Y(_2837_));
 sg13g2_nor2b_1 _3720_ (.A(\main.demo._q___pip_58_1_1___stage___block_3_cx[7] ),
    .B_N(\main.demo._q___pip_58_1_1___stage___block_3_cy[7] ),
    .Y(_2838_));
 sg13g2_nand2b_1 _3721_ (.Y(_2839_),
    .B(\main.demo._q___pip_58_1_1___stage___block_3_cx[7] ),
    .A_N(\main.demo._q___pip_58_1_1___stage___block_3_cy[7] ));
 sg13g2_nor2b_1 _3722_ (.A(\main.demo._q___pip_58_1_1___stage___block_3_cy[6] ),
    .B_N(\main.demo._q___pip_58_1_1___stage___block_3_cx[6] ),
    .Y(_2840_));
 sg13g2_nand2b_2 _3723_ (.Y(_2841_),
    .B(\main.demo._q___pip_58_1_1___stage___block_3_cy[6] ),
    .A_N(\main.demo._q___pip_58_1_1___stage___block_3_cx[6] ));
 sg13g2_nor2b_1 _3724_ (.A(_2840_),
    .B_N(_2841_),
    .Y(_2842_));
 sg13g2_nand2b_2 _3725_ (.Y(_2843_),
    .B(_2841_),
    .A_N(_2840_));
 sg13g2_nor2b_1 _3726_ (.A(\main.demo._q___pip_58_1_1___stage___block_3_cy[4] ),
    .B_N(\main.demo._q___pip_58_1_1___stage___block_3_cx[4] ),
    .Y(_2844_));
 sg13g2_nand2b_2 _3727_ (.Y(_2845_),
    .B(\main.demo._q___pip_58_1_1___stage___block_3_cy[4] ),
    .A_N(\main.demo._q___pip_58_1_1___stage___block_3_cx[4] ));
 sg13g2_nand2b_2 _3728_ (.Y(_2846_),
    .B(_2845_),
    .A_N(_2844_));
 sg13g2_nand2b_1 _3729_ (.Y(_2847_),
    .B(\main.demo._q___pip_58_1_1___stage___block_3_cy[3] ),
    .A_N(\main.demo._q___pip_58_1_1___stage___block_3_cx[3] ));
 sg13g2_nand2b_1 _3730_ (.Y(_2848_),
    .B(\main.demo._q___pip_58_1_1___stage___block_3_cx[3] ),
    .A_N(\main.demo._q___pip_58_1_1___stage___block_3_cy[3] ));
 sg13g2_nor2b_1 _3731_ (.A(\main.demo._q___pip_58_1_1___stage___block_3_cy[2] ),
    .B_N(\main.demo._q___pip_58_1_1___stage___block_3_cx[2] ),
    .Y(_2849_));
 sg13g2_nand2b_2 _3732_ (.Y(_2850_),
    .B(\main.demo._q___pip_58_1_1___stage___block_3_cy[2] ),
    .A_N(\main.demo._q___pip_58_1_1___stage___block_3_cx[2] ));
 sg13g2_nand2b_2 _3733_ (.Y(_2851_),
    .B(_2850_),
    .A_N(_2849_));
 sg13g2_nor2b_1 _3734_ (.A(\main.demo._q___pip_58_1_1___stage___block_3_cx[1] ),
    .B_N(\main.demo._q___pip_58_1_1___stage___block_3_cy[1] ),
    .Y(_2852_));
 sg13g2_nand2b_1 _3735_ (.Y(_2853_),
    .B(\main.demo._q___pip_58_1_1___stage___block_3_cx[1] ),
    .A_N(\main.demo._q___pip_58_1_1___stage___block_3_cy[1] ));
 sg13g2_nor2b_1 _3736_ (.A(\main.demo._q___pip_58_1_1___stage___block_3_cx[0] ),
    .B_N(\main.demo._q___pip_58_1_1___stage___block_3_cy[0] ),
    .Y(_2854_));
 sg13g2_a21oi_1 _3737_ (.A1(_2853_),
    .A2(_2854_),
    .Y(_2855_),
    .B1(_2852_));
 sg13g2_a21o_1 _3738_ (.A2(_2855_),
    .A1(_2850_),
    .B1(_2849_),
    .X(_2856_));
 sg13g2_nand2_1 _3739_ (.Y(_2857_),
    .A(_2847_),
    .B(_2856_));
 sg13g2_nand2_1 _3740_ (.Y(_2858_),
    .A(_2848_),
    .B(_2857_));
 sg13g2_a21o_1 _3741_ (.A2(_2858_),
    .A1(_2845_),
    .B1(_2844_),
    .X(_2859_));
 sg13g2_a21oi_1 _3742_ (.A1(\main.demo._q___pip_58_1_1___stage___block_3_cx[5] ),
    .A2(_2629_),
    .Y(_2860_),
    .B1(_2859_));
 sg13g2_a21oi_2 _3743_ (.B1(_2860_),
    .Y(_2861_),
    .A2(\main.demo._q___pip_58_1_1___stage___block_3_cy[5] ),
    .A1(_2628_));
 sg13g2_a21oi_1 _3744_ (.A1(_2842_),
    .A2(_2861_),
    .Y(_2862_),
    .B1(_2840_));
 sg13g2_o21ai_1 _3745_ (.B1(_2839_),
    .Y(_2863_),
    .A1(_2838_),
    .A2(_2862_));
 sg13g2_a21o_1 _3746_ (.A2(_2863_),
    .A1(_2837_),
    .B1(_2835_),
    .X(_2864_));
 sg13g2_a21oi_1 _3747_ (.A1(_2833_),
    .A2(_2864_),
    .Y(_2865_),
    .B1(_2834_));
 sg13g2_xnor2_1 _3748_ (.Y(_2866_),
    .A(\main.demo._q___pip_58_1_1___stage___block_3_cx[9] ),
    .B(\main.demo._q___pip_58_1_1___stage___block_3_cy[9] ));
 sg13g2_xnor2_1 _3749_ (.Y(_2867_),
    .A(\main.demo._q___pip_58_1_1___stage___block_3_cx[5] ),
    .B(\main.demo._q___pip_58_1_1___stage___block_3_cy[5] ));
 sg13g2_xor2_1 _3750_ (.B(\main.demo._q___pip_58_1_1___stage___block_3_cy[5] ),
    .A(\main.demo._q___pip_58_1_1___stage___block_3_cx[5] ),
    .X(_2868_));
 sg13g2_nand2b_1 _3751_ (.Y(_2869_),
    .B(\main.demo._q___pip_58_1_1___stage___block_3_cx[0] ),
    .A_N(\main.demo._q___pip_58_1_1___stage___block_3_cy[0] ));
 sg13g2_o21ai_1 _3752_ (.B1(_2853_),
    .Y(_2870_),
    .A1(_2852_),
    .A2(_2869_));
 sg13g2_nor2_1 _3753_ (.A(_2851_),
    .B(_2870_),
    .Y(_2871_));
 sg13g2_o21ai_1 _3754_ (.B1(_2848_),
    .Y(_2872_),
    .A1(_2857_),
    .A2(_2871_));
 sg13g2_nor2_1 _3755_ (.A(_2846_),
    .B(_2872_),
    .Y(_2873_));
 sg13g2_nand2_1 _3756_ (.Y(_2874_),
    .A(_2867_),
    .B(_2873_));
 sg13g2_nand2b_2 _3757_ (.Y(_2875_),
    .B(_2839_),
    .A_N(_2838_));
 sg13g2_nor3_1 _3758_ (.A(_2843_),
    .B(_2874_),
    .C(_2875_),
    .Y(_2876_));
 sg13g2_nor2b_1 _3759_ (.A(_2876_),
    .B_N(_2863_),
    .Y(_2877_));
 sg13g2_nor2b_1 _3760_ (.A(_2877_),
    .B_N(_2837_),
    .Y(_2878_));
 sg13g2_a21oi_1 _3761_ (.A1(_2866_),
    .A2(_2878_),
    .Y(_2879_),
    .B1(_2865_));
 sg13g2_and2_1 _3762_ (.A(\main.demo._q___pip_58_1_1___stage___block_3_cx[7] ),
    .B(\main.demo._q___pip_58_1_1___stage___block_3_cy[7] ),
    .X(_2880_));
 sg13g2_nand2_1 _3763_ (.Y(_2881_),
    .A(\main.demo._q___pip_58_1_1___stage___block_3_cx[5] ),
    .B(\main.demo._q___pip_58_1_1___stage___block_3_cy[5] ));
 sg13g2_and2_1 _3764_ (.A(\main.demo._q___pip_58_1_1___stage___block_3_cx[4] ),
    .B(\main.demo._q___pip_58_1_1___stage___block_3_cy[4] ),
    .X(_2882_));
 sg13g2_and2_1 _3765_ (.A(\main.demo._q___pip_58_1_1___stage___block_3_cy[3] ),
    .B(\main.demo._q___pip_58_1_1___stage___block_3_cx[3] ),
    .X(_2883_));
 sg13g2_nand2_2 _3766_ (.Y(_2884_),
    .A(_2847_),
    .B(_2848_));
 sg13g2_and2_1 _3767_ (.A(\main.demo._q___pip_58_1_1___stage___block_3_cx[2] ),
    .B(\main.demo._q___pip_58_1_1___stage___block_3_cy[2] ),
    .X(_2885_));
 sg13g2_nand2_1 _3768_ (.Y(_2886_),
    .A(\main.demo._q___pip_58_1_1___stage___block_3_cx[1] ),
    .B(\main.demo._q___pip_58_1_1___stage___block_3_cy[1] ));
 sg13g2_nor2b_1 _3769_ (.A(_2852_),
    .B_N(_2853_),
    .Y(_2887_));
 sg13g2_nand2_1 _3770_ (.Y(_2888_),
    .A(\main.demo._q___pip_58_1_1___stage___block_3_cx[0] ),
    .B(\main.demo._q___pip_58_1_1___stage___block_3_cy[0] ));
 sg13g2_o21ai_1 _3771_ (.B1(_2886_),
    .Y(_2889_),
    .A1(_2887_),
    .A2(_2888_));
 sg13g2_a21o_1 _3772_ (.A2(_2889_),
    .A1(_2851_),
    .B1(_2885_),
    .X(_2890_));
 sg13g2_a21o_1 _3773_ (.A2(_2890_),
    .A1(_2884_),
    .B1(_2883_),
    .X(_2891_));
 sg13g2_a21o_1 _3774_ (.A2(_2891_),
    .A1(_2846_),
    .B1(_2882_),
    .X(_2892_));
 sg13g2_nand2_1 _3775_ (.Y(_2893_),
    .A(_2868_),
    .B(_2892_));
 sg13g2_a21oi_1 _3776_ (.A1(_2881_),
    .A2(_2893_),
    .Y(_2894_),
    .B1(_2842_));
 sg13g2_a21o_1 _3777_ (.A2(\main.demo._q___pip_58_1_1___stage___block_3_cy[6] ),
    .A1(\main.demo._q___pip_58_1_1___stage___block_3_cx[6] ),
    .B1(_2894_),
    .X(_2895_));
 sg13g2_a21o_1 _3778_ (.A2(_2895_),
    .A1(_2875_),
    .B1(_2880_),
    .X(_2896_));
 sg13g2_nor2b_1 _3779_ (.A(_2837_),
    .B_N(_2896_),
    .Y(_2897_));
 sg13g2_a21o_1 _3780_ (.A2(\main.demo._q___pip_58_1_1___stage___block_3_cy[8] ),
    .A1(\main.demo._q___pip_58_1_1___stage___block_3_cx[8] ),
    .B1(_2897_),
    .X(_2898_));
 sg13g2_nor2b_1 _3781_ (.A(_2866_),
    .B_N(_2898_),
    .Y(_2899_));
 sg13g2_a21oi_1 _3782_ (.A1(\main.demo._q___pip_58_1_1___stage___block_3_cx[9] ),
    .A2(\main.demo._q___pip_58_1_1___stage___block_3_cy[9] ),
    .Y(_2900_),
    .B1(_2899_));
 sg13g2_mux2_1 _3783_ (.A0(_2879_),
    .A1(_2900_),
    .S(net429),
    .X(_2901_));
 sg13g2_xor2_1 _3784_ (.B(_2901_),
    .A(net631),
    .X(\main.demo._d___pip_58_1_1___stage___block_3_a[3] ));
 sg13g2_inv_1 _3785_ (.Y(\main.demo._d___pip_58_1_1___stage___block_3_a[2] ),
    .A(net348));
 sg13g2_xnor2_1 _3786_ (.Y(_2902_),
    .A(\main.demo._q___pip_58_1_1___stage___block_3_cx[0] ),
    .B(\main.demo._q___pip_58_1_1___stage___block_3_cy[0] ));
 sg13g2_xnor2_1 _3787_ (.Y(_2903_),
    .A(_2887_),
    .B(_2888_));
 sg13g2_nand2b_1 _3788_ (.Y(_2904_),
    .B(\main.demo._q___pip_58_1_1___stage___block_3_cx[0] ),
    .A_N(net433));
 sg13g2_xnor2_1 _3789_ (.Y(_2905_),
    .A(_2903_),
    .B(_2904_));
 sg13g2_nand2b_1 _3790_ (.Y(_2906_),
    .B(_2902_),
    .A_N(_2905_));
 sg13g2_xnor2_1 _3791_ (.Y(_2907_),
    .A(_2902_),
    .B(_2905_));
 sg13g2_nand2_1 _3792_ (.Y(_2908_),
    .A(\main.demo._q___pip_58_1_1___stage___block_3_cy[0] ),
    .B(net432));
 sg13g2_xnor2_1 _3793_ (.Y(_2909_),
    .A(_2903_),
    .B(_2908_));
 sg13g2_nor2_1 _3794_ (.A(net347),
    .B(_2909_),
    .Y(_2910_));
 sg13g2_xnor2_1 _3795_ (.Y(_2911_),
    .A(_2851_),
    .B(_2889_));
 sg13g2_inv_1 _3796_ (.Y(_2912_),
    .A(_2911_));
 sg13g2_nor2_1 _3797_ (.A(net433),
    .B(_2911_),
    .Y(_2913_));
 sg13g2_xnor2_1 _3798_ (.Y(_2914_),
    .A(_2851_),
    .B(_2855_));
 sg13g2_a21oi_2 _3799_ (.B1(_2913_),
    .Y(_2915_),
    .A2(_2914_),
    .A1(net433));
 sg13g2_xnor2_1 _3800_ (.Y(_2916_),
    .A(_2910_),
    .B(_2915_));
 sg13g2_nor2b_1 _3801_ (.A(_2905_),
    .B_N(_2916_),
    .Y(_2917_));
 sg13g2_nor2_1 _3802_ (.A(_2902_),
    .B(_2909_),
    .Y(_2918_));
 sg13g2_xnor2_1 _3803_ (.Y(_2919_),
    .A(_2905_),
    .B(_2916_));
 sg13g2_a21oi_1 _3804_ (.A1(_2918_),
    .A2(_2919_),
    .Y(_2920_),
    .B1(_2917_));
 sg13g2_nand2_1 _3805_ (.Y(_2921_),
    .A(_2851_),
    .B(_2870_));
 sg13g2_nor2_1 _3806_ (.A(net432),
    .B(_2871_),
    .Y(_2922_));
 sg13g2_a22oi_1 _3807_ (.Y(_2923_),
    .B1(_2921_),
    .B2(_2922_),
    .A2(_2912_),
    .A1(net433));
 sg13g2_inv_1 _3808_ (.Y(_2924_),
    .A(_2923_));
 sg13g2_nand2_1 _3809_ (.Y(_2925_),
    .A(_2909_),
    .B(_2915_));
 sg13g2_nand2_1 _3810_ (.Y(_2926_),
    .A(\main.demo._d___pip_58_1_1___stage___block_3_a[2] ),
    .B(_2925_));
 sg13g2_nand2_1 _3811_ (.Y(_2927_),
    .A(net432),
    .B(_2856_));
 sg13g2_o21ai_1 _3812_ (.B1(_2927_),
    .Y(_2928_),
    .A1(net432),
    .A2(_2890_));
 sg13g2_xnor2_1 _3813_ (.Y(_2929_),
    .A(_2884_),
    .B(_2928_));
 sg13g2_inv_1 _3814_ (.Y(_2930_),
    .A(_2929_));
 sg13g2_xnor2_1 _3815_ (.Y(_2931_),
    .A(_2926_),
    .B(_2929_));
 sg13g2_xnor2_1 _3816_ (.Y(_2932_),
    .A(_2923_),
    .B(_2931_));
 sg13g2_nor2b_1 _3817_ (.A(_2920_),
    .B_N(_2932_),
    .Y(_2933_));
 sg13g2_xnor2_1 _3818_ (.Y(_2934_),
    .A(_2920_),
    .B(_2932_));
 sg13g2_nand2_1 _3819_ (.Y(_2935_),
    .A(_2907_),
    .B(_2934_));
 sg13g2_xnor2_1 _3820_ (.Y(\main.demo._d___pip_58_1_1___stage___block_3_cx[0] ),
    .A(_2907_),
    .B(_2934_));
 sg13g2_nand2_2 _3821_ (.Y(_2936_),
    .A(net422),
    .B(\main.demo._q_frame[6] ));
 sg13g2_nor2_1 _3822_ (.A(_0060_),
    .B(_2936_),
    .Y(_2937_));
 sg13g2_and2_1 _3823_ (.A(\main.demo._q_frame[6] ),
    .B(\main.demo._q_frame[5] ),
    .X(_2938_));
 sg13g2_xor2_1 _3824_ (.B(\main.demo._q_frame[5] ),
    .A(\main.demo._q_frame[6] ),
    .X(_2939_));
 sg13g2_a21oi_1 _3825_ (.A1(net435),
    .A2(net391),
    .Y(_2940_),
    .B1(_2615_));
 sg13g2_o21ai_1 _3826_ (.B1(_2940_),
    .Y(_2941_),
    .A1(net435),
    .A2(net391));
 sg13g2_nor2_1 _3827_ (.A(_0061_),
    .B(_2941_),
    .Y(_2942_));
 sg13g2_xor2_1 _3828_ (.B(_2936_),
    .A(\main.demo._w_vga_vga_y[8] ),
    .X(_2943_));
 sg13g2_nand2_1 _3829_ (.Y(_2944_),
    .A(_2942_),
    .B(_2943_));
 sg13g2_xnor2_1 _3830_ (.Y(_2945_),
    .A(_2942_),
    .B(_2943_));
 sg13g2_a21oi_1 _3831_ (.A1(net436),
    .A2(net391),
    .Y(_2946_),
    .B1(_2615_));
 sg13g2_o21ai_1 _3832_ (.B1(_2946_),
    .Y(_2947_),
    .A1(net436),
    .A2(net391));
 sg13g2_nor2_1 _3833_ (.A(_0062_),
    .B(_2947_),
    .Y(_2948_));
 sg13g2_xnor2_1 _3834_ (.Y(_2949_),
    .A(_0061_),
    .B(_2941_));
 sg13g2_nand2b_1 _3835_ (.Y(_2950_),
    .B(_2949_),
    .A_N(_2948_));
 sg13g2_xor2_1 _3836_ (.B(_2947_),
    .A(_0062_),
    .X(_2951_));
 sg13g2_a21oi_1 _3837_ (.A1(\main.demo._q_frame[2] ),
    .A2(net391),
    .Y(_2952_),
    .B1(_2615_));
 sg13g2_o21ai_1 _3838_ (.B1(_2952_),
    .Y(_2953_),
    .A1(\main.demo._q_frame[2] ),
    .A2(net391));
 sg13g2_nor2_1 _3839_ (.A(_0063_),
    .B(_2953_),
    .Y(_2954_));
 sg13g2_xnor2_1 _3840_ (.Y(_2955_),
    .A(_2951_),
    .B(_2954_));
 sg13g2_xor2_1 _3841_ (.B(net391),
    .A(\main.demo._q_frame[1] ),
    .X(_2956_));
 sg13g2_a21oi_2 _3842_ (.B1(\main.demo._w_vga_vga_y[4] ),
    .Y(_2957_),
    .A2(_2956_),
    .A1(net422));
 sg13g2_xor2_1 _3843_ (.B(_2953_),
    .A(_0063_),
    .X(_2958_));
 sg13g2_inv_1 _3844_ (.Y(_2959_),
    .A(_2958_));
 sg13g2_a21oi_1 _3845_ (.A1(\main.demo._q_frame[0] ),
    .A2(net392),
    .Y(_2960_),
    .B1(_2615_));
 sg13g2_o21ai_1 _3846_ (.B1(_2960_),
    .Y(_2961_),
    .A1(\main.demo._q_frame[0] ),
    .A2(net391));
 sg13g2_nor2_1 _3847_ (.A(_0001_),
    .B(_2961_),
    .Y(_2962_));
 sg13g2_nand3_1 _3848_ (.B(\main.demo._w_vga_vga_y[4] ),
    .C(_2956_),
    .A(net422),
    .Y(_2963_));
 sg13g2_nand2b_1 _3849_ (.Y(_2964_),
    .B(_2963_),
    .A_N(_2957_));
 sg13g2_nand2_1 _3850_ (.Y(_2965_),
    .A(_2962_),
    .B(_2964_));
 sg13g2_xor2_1 _3851_ (.B(_2964_),
    .A(_2962_),
    .X(_2966_));
 sg13g2_xnor2_1 _3852_ (.Y(_2967_),
    .A(_2957_),
    .B(_2958_));
 sg13g2_xnor2_1 _3853_ (.Y(_2968_),
    .A(_2965_),
    .B(_2967_));
 sg13g2_or2_1 _3854_ (.X(_2969_),
    .B(_2968_),
    .A(_2966_));
 sg13g2_o21ai_1 _3855_ (.B1(_2969_),
    .Y(_2970_),
    .A1(_2957_),
    .A2(_2959_));
 sg13g2_nor2b_1 _3856_ (.A(_2955_),
    .B_N(_2970_),
    .Y(_2971_));
 sg13g2_a21oi_1 _3857_ (.A1(_2951_),
    .A2(_2954_),
    .Y(_2972_),
    .B1(_2948_));
 sg13g2_nor2_1 _3858_ (.A(_2949_),
    .B(_2972_),
    .Y(_2973_));
 sg13g2_o21ai_1 _3859_ (.B1(_2950_),
    .Y(_2974_),
    .A1(_2971_),
    .A2(_2973_));
 sg13g2_xor2_1 _3860_ (.B(_2974_),
    .A(_2945_),
    .X(_2975_));
 sg13g2_o21ai_1 _3861_ (.B1(_2944_),
    .Y(_2976_),
    .A1(_2945_),
    .A2(_2974_));
 sg13g2_a21oi_1 _3862_ (.A1(\main.demo._w_vga_vga_y[8] ),
    .A2(_2936_),
    .Y(_2977_),
    .B1(\main.demo._w_vga_vga_y[10] ));
 sg13g2_nand3_1 _3863_ (.B(\main.demo._w_vga_vga_y[8] ),
    .C(_2936_),
    .A(\main.demo._w_vga_vga_y[10] ),
    .Y(_2978_));
 sg13g2_nand2b_1 _3864_ (.Y(_2979_),
    .B(_2978_),
    .A_N(_2977_));
 sg13g2_xor2_1 _3865_ (.B(_2979_),
    .A(_2976_),
    .X(_2980_));
 sg13g2_nor2_1 _3866_ (.A(_2975_),
    .B(_2980_),
    .Y(_2981_));
 sg13g2_a22oi_1 _3867_ (.Y(_2982_),
    .B1(_2944_),
    .B2(_2977_),
    .A2(_2936_),
    .A1(\main.demo._w_vga_vga_y[10] ));
 sg13g2_nor2_1 _3868_ (.A(_2981_),
    .B(_2982_),
    .Y(_2983_));
 sg13g2_xnor2_1 _3869_ (.Y(\main.demo._t___pip_58_1_0___stage___block_3_a[6] ),
    .A(_2937_),
    .B(_2983_));
 sg13g2_nand2_1 _3870_ (.Y(_2984_),
    .A(\main.demo._q_rot_en ),
    .B(net434));
 sg13g2_nor2_1 _3871_ (.A(_0054_),
    .B(_2984_),
    .Y(_2985_));
 sg13g2_xor2_1 _3872_ (.B(_2984_),
    .A(_0054_),
    .X(_2986_));
 sg13g2_a21oi_1 _3873_ (.A1(net434),
    .A2(net392),
    .Y(_2987_),
    .B1(_2615_));
 sg13g2_o21ai_1 _3874_ (.B1(_2987_),
    .Y(_2988_),
    .A1(net434),
    .A2(net392));
 sg13g2_nand2_1 _3875_ (.Y(_2989_),
    .A(_0055_),
    .B(_2988_));
 sg13g2_and2_1 _3876_ (.A(_2986_),
    .B(_2989_),
    .X(_2990_));
 sg13g2_xor2_1 _3877_ (.B(\main.demo._q_frame[6] ),
    .A(net434),
    .X(_2991_));
 sg13g2_a21oi_1 _3878_ (.A1(net435),
    .A2(_2991_),
    .Y(_2992_),
    .B1(_2615_));
 sg13g2_o21ai_1 _3879_ (.B1(_2992_),
    .Y(_2993_),
    .A1(net435),
    .A2(_2991_));
 sg13g2_nand2_1 _3880_ (.Y(_2994_),
    .A(_0056_),
    .B(_2993_));
 sg13g2_xnor2_1 _3881_ (.Y(_2995_),
    .A(_2631_),
    .B(_2988_));
 sg13g2_nand2_1 _3882_ (.Y(_2996_),
    .A(_2994_),
    .B(_2995_));
 sg13g2_xor2_1 _3883_ (.B(_2995_),
    .A(_2994_),
    .X(_2997_));
 sg13g2_inv_1 _3884_ (.Y(_2998_),
    .A(_2997_));
 sg13g2_a21oi_1 _3885_ (.A1(net436),
    .A2(_2991_),
    .Y(_2999_),
    .B1(_2615_));
 sg13g2_o21ai_1 _3886_ (.B1(_2999_),
    .Y(_3000_),
    .A1(net436),
    .A2(_2991_));
 sg13g2_xnor2_1 _3887_ (.Y(_3001_),
    .A(_0057_),
    .B(_3000_));
 sg13g2_o21ai_1 _3888_ (.B1(net422),
    .Y(_3002_),
    .A1(\main.demo._q_frame[2] ),
    .A2(_2991_));
 sg13g2_a21oi_1 _3889_ (.A1(\main.demo._q_frame[2] ),
    .A2(_2991_),
    .Y(_3003_),
    .B1(_3002_));
 sg13g2_nand2b_1 _3890_ (.Y(_3004_),
    .B(_3003_),
    .A_N(_0058_));
 sg13g2_o21ai_1 _3891_ (.B1(net422),
    .Y(_3005_),
    .A1(\main.demo._q_frame[1] ),
    .A2(_2991_));
 sg13g2_a21oi_1 _3892_ (.A1(\main.demo._q_frame[1] ),
    .A2(_2991_),
    .Y(_3006_),
    .B1(_3005_));
 sg13g2_nor2b_1 _3893_ (.A(_0059_),
    .B_N(_3006_),
    .Y(_3007_));
 sg13g2_xnor2_1 _3894_ (.Y(_3008_),
    .A(_0058_),
    .B(_3003_));
 sg13g2_nand2_1 _3895_ (.Y(_3009_),
    .A(_3007_),
    .B(_3008_));
 sg13g2_a21o_1 _3896_ (.A2(_3009_),
    .A1(_3004_),
    .B1(_3001_),
    .X(_3010_));
 sg13g2_o21ai_1 _3897_ (.B1(_3010_),
    .Y(_3011_),
    .A1(_0057_),
    .A2(_3000_));
 sg13g2_xnor2_1 _3898_ (.Y(_3012_),
    .A(_2632_),
    .B(_2993_));
 sg13g2_nand2_1 _3899_ (.Y(_3013_),
    .A(_3011_),
    .B(_3012_));
 sg13g2_o21ai_1 _3900_ (.B1(_2996_),
    .Y(_3014_),
    .A1(_2998_),
    .A2(_3013_));
 sg13g2_xor2_1 _3901_ (.B(_2989_),
    .A(_2986_),
    .X(_3015_));
 sg13g2_a21o_1 _3902_ (.A2(_3015_),
    .A1(_3014_),
    .B1(_2990_),
    .X(_3016_));
 sg13g2_nand3_1 _3903_ (.B(net434),
    .C(_0054_),
    .A(net422),
    .Y(_3017_));
 sg13g2_xnor2_1 _3904_ (.Y(_3018_),
    .A(_2630_),
    .B(_3017_));
 sg13g2_a22oi_1 _3905_ (.Y(_3019_),
    .B1(_3016_),
    .B2(_3018_),
    .A2(_2985_),
    .A1(\main.demo._w_vga_vga_x[9] ));
 sg13g2_a21oi_1 _3906_ (.A1(net422),
    .A2(net434),
    .Y(_3020_),
    .B1(_0053_));
 sg13g2_xor2_1 _3907_ (.B(_3020_),
    .A(\main.demo._w_vga_vga_x[10] ),
    .X(_3021_));
 sg13g2_xnor2_1 _3908_ (.Y(_3022_),
    .A(_3019_),
    .B(_3021_));
 sg13g2_nor2b_1 _3909_ (.A(net353),
    .B_N(_3022_),
    .Y(_3023_));
 sg13g2_inv_2 _3910_ (.Y(\main.demo._t___pip_58_1_0___stage___block_3_a[7] ),
    .A(net346));
 sg13g2_nor2_1 _3911_ (.A(net452),
    .B(net309),
    .Y(_3024_));
 sg13g2_nor4_2 _3912_ (.A(\main.demo.vga._q_xcount[1] ),
    .B(\main.demo.vga._q_xcount[0] ),
    .C(\main.demo.vga._q_xcount[3] ),
    .Y(_3025_),
    .D(\main.demo.vga._q_xcount[2] ));
 sg13g2_nor2_1 _3913_ (.A(\main.demo.vga._q_xcount[5] ),
    .B(\main.demo.vga._q_xcount[4] ),
    .Y(_3026_));
 sg13g2_and2_1 _3914_ (.A(\main.demo.vga._q_xcount[7] ),
    .B(_3026_),
    .X(_3027_));
 sg13g2_nor2_1 _3915_ (.A(\main.demo.vga._q_xcount[6] ),
    .B(\main.demo.vga._q_xcount[10] ),
    .Y(_3028_));
 sg13g2_nor2b_1 _3916_ (.A(\main.demo.vga._q_xcount[8] ),
    .B_N(\main.demo.vga._q_xcount[9] ),
    .Y(_0230_));
 sg13g2_and4_1 _3917_ (.A(_3025_),
    .B(_3027_),
    .C(_3028_),
    .D(_0230_),
    .X(_0231_));
 sg13g2_nor3_1 _3918_ (.A(\main.demo.vga._q_xcount[7] ),
    .B(\main.demo.vga._q_xcount[9] ),
    .C(\main.demo.vga._q_xcount[8] ),
    .Y(_0232_));
 sg13g2_nand4_1 _3919_ (.B(_3026_),
    .C(_3028_),
    .A(_3025_),
    .Y(_0233_),
    .D(_0232_));
 sg13g2_o21ai_1 _3920_ (.B1(_0233_),
    .Y(_0234_),
    .A1(_2639_),
    .A2(_0231_));
 sg13g2_inv_1 _3921_ (.Y(_0235_),
    .A(net366));
 sg13g2_nand4_1 _3922_ (.B(net620),
    .C(\main.demo.vga._q_ycount[6] ),
    .A(net469),
    .Y(_0236_),
    .D(net319));
 sg13g2_nor4_2 _3923_ (.A(\main.demo.vga._q_ycount[3] ),
    .B(\main.demo.vga._q_ycount[2] ),
    .C(net645),
    .Y(_0237_),
    .D(\main.demo.vga._q_ycount[0] ));
 sg13g2_inv_1 _3924_ (.Y(_0238_),
    .A(_0237_));
 sg13g2_nor4_2 _3925_ (.A(net501),
    .B(net485),
    .C(net621),
    .Y(_0239_),
    .D(_0238_));
 sg13g2_nor2b_2 _3926_ (.A(_0239_),
    .B_N(net553),
    .Y(_0240_));
 sg13g2_or4_1 _3927_ (.A(\main.demo.vga._q_ycount[8] ),
    .B(\main.demo.vga._q_ycount[7] ),
    .C(\main.demo.vga._q_ycount[6] ),
    .D(\main.demo.vga._q_ycount[5] ),
    .X(_0241_));
 sg13g2_nor3_1 _3928_ (.A(\main.demo.vga._q_ycount[4] ),
    .B(\main.demo.vga._d_vblank ),
    .C(_0241_),
    .Y(_0242_));
 sg13g2_a21oi_2 _3929_ (.B1(_0240_),
    .Y(_0243_),
    .A2(_0242_),
    .A1(_0237_));
 sg13g2_nor2_1 _3930_ (.A(_0235_),
    .B(_0243_),
    .Y(\main.demo.vga._d_active ));
 sg13g2_nand2_1 _3931_ (.Y(_0244_),
    .A(net415),
    .B(net356));
 sg13g2_o21ai_1 _3932_ (.B1(_0244_),
    .Y(\main.demo._t___pip_58_1_0___stage___block_3_cy[0] ),
    .A1(_2640_),
    .A2(net356));
 sg13g2_xor2_1 _3933_ (.B(\main.demo._t___stage___block_3_x[1] ),
    .A(net415),
    .X(_0245_));
 sg13g2_nand2_1 _3934_ (.Y(_0246_),
    .A(net355),
    .B(_0245_));
 sg13g2_nor2_1 _3935_ (.A(_2640_),
    .B(_3022_),
    .Y(_0247_));
 sg13g2_xnor2_1 _3936_ (.Y(_0248_),
    .A(net407),
    .B(_0247_));
 sg13g2_o21ai_1 _3937_ (.B1(_0246_),
    .Y(\main.demo._t___pip_58_1_0___stage___block_3_cy[1] ),
    .A1(net356),
    .A2(_0248_));
 sg13g2_nor3_2 _3938_ (.A(net415),
    .B(\main.demo._t___stage___block_3_x[1] ),
    .C(\main.demo._t___stage___block_3_x[2] ),
    .Y(_0249_));
 sg13g2_o21ai_1 _3939_ (.B1(\main.demo._t___stage___block_3_x[2] ),
    .Y(_0250_),
    .A1(net415),
    .A2(\main.demo._t___stage___block_3_x[1] ));
 sg13g2_nor2b_1 _3940_ (.A(_0249_),
    .B_N(_0250_),
    .Y(_0251_));
 sg13g2_nand2_1 _3941_ (.Y(_0252_),
    .A(net355),
    .B(_0251_));
 sg13g2_nor2_1 _3942_ (.A(\main.demo._t___stage___block_3_y[0] ),
    .B(net407),
    .Y(_0253_));
 sg13g2_nor2_1 _3943_ (.A(_3022_),
    .B(_0253_),
    .Y(_0254_));
 sg13g2_xor2_1 _3944_ (.B(_0254_),
    .A(net632),
    .X(_0255_));
 sg13g2_o21ai_1 _3945_ (.B1(_0252_),
    .Y(\main.demo._t___pip_58_1_0___stage___block_3_cy[2] ),
    .A1(net356),
    .A2(_0255_));
 sg13g2_xnor2_1 _3946_ (.Y(_0256_),
    .A(_0059_),
    .B(_3006_));
 sg13g2_nor2b_1 _3947_ (.A(_0256_),
    .B_N(_0249_),
    .Y(_0257_));
 sg13g2_xnor2_1 _3948_ (.Y(_0258_),
    .A(_0249_),
    .B(_0256_));
 sg13g2_xor2_1 _3949_ (.B(_2961_),
    .A(net643),
    .X(_0259_));
 sg13g2_a21oi_1 _3950_ (.A1(_2643_),
    .A2(_0253_),
    .Y(_0260_),
    .B1(_3022_));
 sg13g2_xor2_1 _3951_ (.B(_0260_),
    .A(_0259_),
    .X(_0261_));
 sg13g2_mux2_1 _3952_ (.A0(_0261_),
    .A1(_0258_),
    .S(net355),
    .X(\main.demo._t___pip_58_1_0___stage___block_3_cy[3] ));
 sg13g2_xor2_1 _3953_ (.B(_3008_),
    .A(_3007_),
    .X(_0262_));
 sg13g2_nand2b_1 _3954_ (.Y(_0263_),
    .B(_0257_),
    .A_N(_0262_));
 sg13g2_xnor2_1 _3955_ (.Y(_0264_),
    .A(_0257_),
    .B(_0262_));
 sg13g2_nand2_1 _3956_ (.Y(_0265_),
    .A(net355),
    .B(_0264_));
 sg13g2_nand3b_1 _3957_ (.B(_0253_),
    .C(_0003_),
    .Y(_0266_),
    .A_N(_0259_));
 sg13g2_nor2b_1 _3958_ (.A(_3022_),
    .B_N(_0266_),
    .Y(_0267_));
 sg13g2_xnor2_1 _3959_ (.Y(_0268_),
    .A(_2966_),
    .B(_0267_));
 sg13g2_o21ai_1 _3960_ (.B1(_0265_),
    .Y(\main.demo._t___pip_58_1_0___stage___block_3_cy[4] ),
    .A1(net353),
    .A2(_0268_));
 sg13g2_o21ai_1 _3961_ (.B1(_2968_),
    .Y(_0269_),
    .A1(_2966_),
    .A2(_0266_));
 sg13g2_nor2_1 _3962_ (.A(_2969_),
    .B(_0266_),
    .Y(_0270_));
 sg13g2_nor2_1 _3963_ (.A(_3022_),
    .B(_0270_),
    .Y(_0271_));
 sg13g2_nand2_1 _3964_ (.Y(_0272_),
    .A(_0269_),
    .B(_0271_));
 sg13g2_nand3_1 _3965_ (.B(_3004_),
    .C(_3009_),
    .A(_3001_),
    .Y(_0273_));
 sg13g2_and2_1 _3966_ (.A(_3010_),
    .B(_0273_),
    .X(_0274_));
 sg13g2_nor2_1 _3967_ (.A(_0263_),
    .B(_0274_),
    .Y(_0275_));
 sg13g2_xor2_1 _3968_ (.B(_0274_),
    .A(_0263_),
    .X(_0276_));
 sg13g2_nor2_2 _3969_ (.A(net353),
    .B(_3022_),
    .Y(_0277_));
 sg13g2_inv_1 _3970_ (.Y(_0278_),
    .A(net345));
 sg13g2_a22oi_1 _3971_ (.Y(_0279_),
    .B1(_0276_),
    .B2(net353),
    .A2(_3023_),
    .A1(_2968_));
 sg13g2_o21ai_1 _3972_ (.B1(_0279_),
    .Y(\main.demo._t___pip_58_1_0___stage___block_3_cy[5] ),
    .A1(net353),
    .A2(_0272_));
 sg13g2_xnor2_1 _3973_ (.Y(_0280_),
    .A(_3011_),
    .B(_3012_));
 sg13g2_nand2_1 _3974_ (.Y(_0281_),
    .A(_0275_),
    .B(_0280_));
 sg13g2_xor2_1 _3975_ (.B(_0280_),
    .A(_0275_),
    .X(_0282_));
 sg13g2_xor2_1 _3976_ (.B(_2970_),
    .A(_2955_),
    .X(_0283_));
 sg13g2_inv_1 _3977_ (.Y(_0284_),
    .A(_0283_));
 sg13g2_xnor2_1 _3978_ (.Y(_0285_),
    .A(_0271_),
    .B(_0284_));
 sg13g2_nand2_1 _3979_ (.Y(_0286_),
    .A(net357),
    .B(_0282_));
 sg13g2_o21ai_1 _3980_ (.B1(_0286_),
    .Y(\main.demo._t___pip_58_1_0___stage___block_3_cy[6] ),
    .A1(net354),
    .A2(_0285_));
 sg13g2_a21oi_1 _3981_ (.A1(_2951_),
    .A2(_2954_),
    .Y(_0287_),
    .B1(_2971_));
 sg13g2_xnor2_1 _3982_ (.Y(_0288_),
    .A(_2948_),
    .B(_2949_));
 sg13g2_xnor2_1 _3983_ (.Y(_0289_),
    .A(_0287_),
    .B(_0288_));
 sg13g2_nand2_1 _3984_ (.Y(_0290_),
    .A(_0270_),
    .B(_0283_));
 sg13g2_or2_1 _3985_ (.X(_0291_),
    .B(_0290_),
    .A(_0289_));
 sg13g2_inv_1 _3986_ (.Y(_0292_),
    .A(_0291_));
 sg13g2_xnor2_1 _3987_ (.Y(_0293_),
    .A(_0289_),
    .B(_0290_));
 sg13g2_xnor2_1 _3988_ (.Y(_0294_),
    .A(_2998_),
    .B(_3013_));
 sg13g2_nor2b_1 _3989_ (.A(_0281_),
    .B_N(_0294_),
    .Y(_0295_));
 sg13g2_xnor2_1 _3990_ (.Y(_0296_),
    .A(_0281_),
    .B(_0294_));
 sg13g2_a22oi_1 _3991_ (.Y(_0297_),
    .B1(_0296_),
    .B2(net354),
    .A2(_0289_),
    .A1(net346));
 sg13g2_o21ai_1 _3992_ (.B1(_0297_),
    .Y(\main.demo._t___pip_58_1_0___stage___block_3_cy[7] ),
    .A1(_0278_),
    .A2(_0293_));
 sg13g2_xnor2_1 _3993_ (.Y(_0298_),
    .A(_2975_),
    .B(_0291_));
 sg13g2_xor2_1 _3994_ (.B(_3015_),
    .A(_3014_),
    .X(_0299_));
 sg13g2_nor2b_1 _3995_ (.A(_0299_),
    .B_N(_0295_),
    .Y(_0300_));
 sg13g2_xnor2_1 _3996_ (.Y(_0301_),
    .A(_0295_),
    .B(_0299_));
 sg13g2_a22oi_1 _3997_ (.Y(_0302_),
    .B1(_0301_),
    .B2(net354),
    .A2(net346),
    .A1(_2975_));
 sg13g2_o21ai_1 _3998_ (.B1(_0302_),
    .Y(\main.demo._t___pip_58_1_0___stage___block_3_cy[8] ),
    .A1(_0278_),
    .A2(_0298_));
 sg13g2_o21ai_1 _3999_ (.B1(_2980_),
    .Y(_0303_),
    .A1(_2975_),
    .A2(_0291_));
 sg13g2_a21oi_1 _4000_ (.A1(_2981_),
    .A2(_0292_),
    .Y(_0304_),
    .B1(_0278_));
 sg13g2_xor2_1 _4001_ (.B(_3018_),
    .A(_3016_),
    .X(_0305_));
 sg13g2_nand2b_1 _4002_ (.Y(_0306_),
    .B(_0300_),
    .A_N(_0305_));
 sg13g2_xnor2_1 _4003_ (.Y(_0307_),
    .A(_0300_),
    .B(_0305_));
 sg13g2_nand2_1 _4004_ (.Y(_0308_),
    .A(net354),
    .B(_0307_));
 sg13g2_a22oi_1 _4005_ (.Y(_0309_),
    .B1(_0303_),
    .B2(_0304_),
    .A2(net346),
    .A1(_2980_));
 sg13g2_nand2_1 _4006_ (.Y(\main.demo._t___pip_58_1_0___stage___block_3_cy[9] ),
    .A(_0308_),
    .B(_0309_));
 sg13g2_xor2_1 _4007_ (.B(_0306_),
    .A(_3022_),
    .X(_0310_));
 sg13g2_a21oi_1 _4008_ (.A1(net354),
    .A2(_0310_),
    .Y(\main.demo._t___pip_58_1_0___stage___block_3_cy[10] ),
    .B1(_0304_));
 sg13g2_a22oi_1 _4009_ (.Y(_0311_),
    .B1(_0277_),
    .B2(net415),
    .A2(net355),
    .A1(\main.demo._t___stage___block_3_y[0] ));
 sg13g2_o21ai_1 _4010_ (.B1(_0311_),
    .Y(\main.demo._t___pip_58_1_0___stage___block_3_cx[0] ),
    .A1(net600),
    .A2(\main.demo._t___pip_58_1_0___stage___block_3_a[7] ));
 sg13g2_a22oi_1 _4011_ (.Y(_0312_),
    .B1(_0245_),
    .B2(_0277_),
    .A2(net355),
    .A1(net407));
 sg13g2_o21ai_1 _4012_ (.B1(_0312_),
    .Y(\main.demo._t___pip_58_1_0___stage___block_3_cx[1] ),
    .A1(net517),
    .A2(\main.demo._t___pip_58_1_0___stage___block_3_a[7] ));
 sg13g2_nand2_1 _4013_ (.Y(_0313_),
    .A(net587),
    .B(net355));
 sg13g2_a22oi_1 _4014_ (.Y(_0314_),
    .B1(_0251_),
    .B2(net345),
    .A2(net346),
    .A1(\main.demo._t___stage___block_3_x[2] ));
 sg13g2_nand2_1 _4015_ (.Y(\main.demo._t___pip_58_1_0___stage___block_3_cx[2] ),
    .A(_0313_),
    .B(_0314_));
 sg13g2_nand2_1 _4016_ (.Y(_0315_),
    .A(net355),
    .B(_0259_));
 sg13g2_a22oi_1 _4017_ (.Y(_0316_),
    .B1(_0258_),
    .B2(net345),
    .A2(_0256_),
    .A1(net346));
 sg13g2_nand2_1 _4018_ (.Y(\main.demo._t___pip_58_1_0___stage___block_3_cx[3] ),
    .A(_0315_),
    .B(_0316_));
 sg13g2_nand2_1 _4019_ (.Y(_0317_),
    .A(_2966_),
    .B(net353));
 sg13g2_a22oi_1 _4020_ (.Y(_0318_),
    .B1(_0264_),
    .B2(_0277_),
    .A2(_0262_),
    .A1(_3023_));
 sg13g2_nand2_1 _4021_ (.Y(\main.demo._t___pip_58_1_0___stage___block_3_cx[4] ),
    .A(_0317_),
    .B(_0318_));
 sg13g2_nand2_1 _4022_ (.Y(_0319_),
    .A(_2968_),
    .B(net353));
 sg13g2_a22oi_1 _4023_ (.Y(_0320_),
    .B1(_0276_),
    .B2(net345),
    .A2(_0274_),
    .A1(_3023_));
 sg13g2_nand2_1 _4024_ (.Y(\main.demo._t___pip_58_1_0___stage___block_3_cx[5] ),
    .A(_0319_),
    .B(_0320_));
 sg13g2_a22oi_1 _4025_ (.Y(_0321_),
    .B1(_0284_),
    .B2(net353),
    .A2(_0282_),
    .A1(net345));
 sg13g2_o21ai_1 _4026_ (.B1(_0321_),
    .Y(\main.demo._t___pip_58_1_0___stage___block_3_cx[6] ),
    .A1(\main.demo._t___pip_58_1_0___stage___block_3_a[7] ),
    .A2(_0280_));
 sg13g2_a22oi_1 _4027_ (.Y(_0322_),
    .B1(_0296_),
    .B2(net345),
    .A2(_0289_),
    .A1(net354));
 sg13g2_o21ai_1 _4028_ (.B1(_0322_),
    .Y(\main.demo._t___pip_58_1_0___stage___block_3_cx[7] ),
    .A1(\main.demo._t___pip_58_1_0___stage___block_3_a[7] ),
    .A2(_0294_));
 sg13g2_nand2_1 _4029_ (.Y(_0323_),
    .A(_2975_),
    .B(net354));
 sg13g2_a22oi_1 _4030_ (.Y(_0324_),
    .B1(_0301_),
    .B2(net345),
    .A2(_0299_),
    .A1(net346));
 sg13g2_nand2_1 _4031_ (.Y(\main.demo._t___pip_58_1_0___stage___block_3_cx[8] ),
    .A(_0323_),
    .B(_0324_));
 sg13g2_nand2_1 _4032_ (.Y(_0325_),
    .A(_2980_),
    .B(net354));
 sg13g2_a22oi_1 _4033_ (.Y(_0326_),
    .B1(_0307_),
    .B2(net345),
    .A2(_0305_),
    .A1(net346));
 sg13g2_nand2_1 _4034_ (.Y(\main.demo._t___pip_58_1_0___stage___block_3_cx[9] ),
    .A(_0325_),
    .B(_0326_));
 sg13g2_nor2_1 _4035_ (.A(_0278_),
    .B(_0306_),
    .Y(\main.demo._t___pip_58_1_0___stage___block_3_cx[10] ));
 sg13g2_nor2_1 _4036_ (.A(_2925_),
    .B(_2929_),
    .Y(_0327_));
 sg13g2_xor2_1 _4037_ (.B(_2891_),
    .A(_2846_),
    .X(_0328_));
 sg13g2_nor2b_1 _4038_ (.A(net432),
    .B_N(_0328_),
    .Y(_0329_));
 sg13g2_xnor2_1 _4039_ (.Y(_0330_),
    .A(_2846_),
    .B(_2858_));
 sg13g2_a21oi_2 _4040_ (.B1(_0329_),
    .Y(_0331_),
    .A2(_0330_),
    .A1(net432));
 sg13g2_nand2_1 _4041_ (.Y(_0332_),
    .A(_0327_),
    .B(_0331_));
 sg13g2_nor2_1 _4042_ (.A(net431),
    .B(_2892_),
    .Y(_0333_));
 sg13g2_a21oi_1 _4043_ (.A1(net431),
    .A2(_2859_),
    .Y(_0334_),
    .B1(_0333_));
 sg13g2_xnor2_1 _4044_ (.Y(_0335_),
    .A(_2867_),
    .B(_0334_));
 sg13g2_inv_1 _4045_ (.Y(_0336_),
    .A(_0335_));
 sg13g2_nor2_1 _4046_ (.A(_0332_),
    .B(_0335_),
    .Y(_0337_));
 sg13g2_nand3_1 _4047_ (.B(_2881_),
    .C(_2893_),
    .A(_2842_),
    .Y(_0338_));
 sg13g2_nor2b_1 _4048_ (.A(_2894_),
    .B_N(_0338_),
    .Y(_0339_));
 sg13g2_nor2b_1 _4049_ (.A(net431),
    .B_N(_0339_),
    .Y(_0340_));
 sg13g2_xnor2_1 _4050_ (.Y(_0341_),
    .A(_2843_),
    .B(_2861_));
 sg13g2_a21oi_2 _4051_ (.B1(_0340_),
    .Y(_0342_),
    .A2(_0341_),
    .A1(net431));
 sg13g2_nand2_1 _4052_ (.Y(_0343_),
    .A(_0337_),
    .B(_0342_));
 sg13g2_mux2_1 _4053_ (.A0(_2895_),
    .A1(_2862_),
    .S(net430),
    .X(_0344_));
 sg13g2_xnor2_1 _4054_ (.Y(_0345_),
    .A(_2875_),
    .B(_0344_));
 sg13g2_nor2b_1 _4055_ (.A(_0343_),
    .B_N(_0345_),
    .Y(_0346_));
 sg13g2_xnor2_1 _4056_ (.Y(_0347_),
    .A(_2837_),
    .B(_2896_));
 sg13g2_xor2_1 _4057_ (.B(_2863_),
    .A(_2837_),
    .X(_0348_));
 sg13g2_mux2_1 _4058_ (.A0(_0347_),
    .A1(_0348_),
    .S(net429),
    .X(_0349_));
 sg13g2_inv_1 _4059_ (.Y(_0350_),
    .A(_0349_));
 sg13g2_nand2_1 _4060_ (.Y(_0351_),
    .A(_0346_),
    .B(_0350_));
 sg13g2_nor2_1 _4061_ (.A(net429),
    .B(_2898_),
    .Y(_0352_));
 sg13g2_a21oi_1 _4062_ (.A1(net429),
    .A2(_2864_),
    .Y(_0353_),
    .B1(_0352_));
 sg13g2_xnor2_1 _4063_ (.Y(_0354_),
    .A(_2866_),
    .B(_0353_));
 sg13g2_nor2_1 _4064_ (.A(_0351_),
    .B(_0354_),
    .Y(_0355_));
 sg13g2_mux2_1 _4065_ (.A0(_2900_),
    .A1(_2865_),
    .S(net429),
    .X(_0356_));
 sg13g2_xnor2_1 _4066_ (.Y(_0357_),
    .A(\main.demo._q___pip_58_1_1___stage___block_3_cx[10] ),
    .B(_0356_));
 sg13g2_a21oi_2 _4067_ (.B1(_0357_),
    .Y(_0358_),
    .A2(_0355_),
    .A1(net344));
 sg13g2_nor2_1 _4068_ (.A(net429),
    .B(_2878_),
    .Y(_0359_));
 sg13g2_a22oi_1 _4069_ (.Y(_0360_),
    .B1(_0359_),
    .B2(_2836_),
    .A2(_2898_),
    .A1(net429));
 sg13g2_xnor2_1 _4070_ (.Y(_0361_),
    .A(_2866_),
    .B(_0360_));
 sg13g2_nor2_1 _4071_ (.A(net347),
    .B(_0355_),
    .Y(_0362_));
 sg13g2_xnor2_1 _4072_ (.Y(_0363_),
    .A(_0357_),
    .B(_0362_));
 sg13g2_nand2b_1 _4073_ (.Y(_0364_),
    .B(_2877_),
    .A_N(_2837_));
 sg13g2_a22oi_1 _4074_ (.Y(_0365_),
    .B1(_0359_),
    .B2(_0364_),
    .A2(_0347_),
    .A1(net429));
 sg13g2_nand2_1 _4075_ (.Y(_0366_),
    .A(net344),
    .B(_0351_));
 sg13g2_xor2_1 _4076_ (.B(_0366_),
    .A(_0354_),
    .X(_0367_));
 sg13g2_nor2_1 _4077_ (.A(_0365_),
    .B(_0367_),
    .Y(_0368_));
 sg13g2_a21oi_1 _4078_ (.A1(_2861_),
    .A2(_2874_),
    .Y(_0369_),
    .B1(_2843_));
 sg13g2_nor2_1 _4079_ (.A(net430),
    .B(_0369_),
    .Y(_0370_));
 sg13g2_a22oi_1 _4080_ (.Y(_0371_),
    .B1(_0370_),
    .B2(_2841_),
    .A2(_2895_),
    .A1(net430));
 sg13g2_xnor2_1 _4081_ (.Y(_0372_),
    .A(_2875_),
    .B(_0371_));
 sg13g2_nor2_1 _4082_ (.A(net347),
    .B(_0346_),
    .Y(_0373_));
 sg13g2_xnor2_1 _4083_ (.Y(_0374_),
    .A(_0350_),
    .B(_0373_));
 sg13g2_nand3_1 _4084_ (.B(_2861_),
    .C(_2874_),
    .A(_2843_),
    .Y(_0375_));
 sg13g2_a22oi_1 _4085_ (.Y(_0376_),
    .B1(_0370_),
    .B2(_0375_),
    .A2(_0339_),
    .A1(net431));
 sg13g2_nand2_1 _4086_ (.Y(_0377_),
    .A(net344),
    .B(_0343_));
 sg13g2_xnor2_1 _4087_ (.Y(_0378_),
    .A(_0345_),
    .B(_0377_));
 sg13g2_nor2_1 _4088_ (.A(_0376_),
    .B(_0378_),
    .Y(_0379_));
 sg13g2_nand2_1 _4089_ (.Y(_0380_),
    .A(_0376_),
    .B(_0378_));
 sg13g2_nand2b_1 _4090_ (.Y(_0381_),
    .B(_0380_),
    .A_N(_0379_));
 sg13g2_nor2_1 _4091_ (.A(net431),
    .B(_2873_),
    .Y(_0382_));
 sg13g2_a22oi_1 _4092_ (.Y(_0383_),
    .B1(_0382_),
    .B2(_2845_),
    .A2(_2892_),
    .A1(net431));
 sg13g2_xnor2_1 _4093_ (.Y(_0384_),
    .A(_2868_),
    .B(_0383_));
 sg13g2_nor2_1 _4094_ (.A(net347),
    .B(_0337_),
    .Y(_0385_));
 sg13g2_xnor2_1 _4095_ (.Y(_0386_),
    .A(_0342_),
    .B(_0385_));
 sg13g2_nand2_1 _4096_ (.Y(_0387_),
    .A(_2846_),
    .B(_2872_));
 sg13g2_a22oi_1 _4097_ (.Y(_0388_),
    .B1(_0382_),
    .B2(_0387_),
    .A2(_0328_),
    .A1(net432));
 sg13g2_nand2_1 _4098_ (.Y(_0389_),
    .A(net344),
    .B(_0332_));
 sg13g2_xnor2_1 _4099_ (.Y(_0390_),
    .A(_0336_),
    .B(_0389_));
 sg13g2_nor2_1 _4100_ (.A(_0388_),
    .B(_0390_),
    .Y(_0391_));
 sg13g2_xnor2_1 _4101_ (.Y(_0392_),
    .A(_0388_),
    .B(_0390_));
 sg13g2_inv_1 _4102_ (.Y(_0393_),
    .A(_0392_));
 sg13g2_a22oi_1 _4103_ (.Y(_0394_),
    .B1(_2922_),
    .B2(_2850_),
    .A2(_2890_),
    .A1(net432));
 sg13g2_xnor2_1 _4104_ (.Y(_0395_),
    .A(_2884_),
    .B(_0394_));
 sg13g2_nor2_1 _4105_ (.A(net348),
    .B(_0327_),
    .Y(_0396_));
 sg13g2_xnor2_1 _4106_ (.Y(_0397_),
    .A(_0331_),
    .B(_0396_));
 sg13g2_a21oi_1 _4107_ (.A1(_2924_),
    .A2(_2931_),
    .Y(_0398_),
    .B1(_2933_));
 sg13g2_xor2_1 _4108_ (.B(_0397_),
    .A(_0395_),
    .X(_0399_));
 sg13g2_nor2b_1 _4109_ (.A(_0398_),
    .B_N(_0399_),
    .Y(_0400_));
 sg13g2_a21o_1 _4110_ (.A2(_0397_),
    .A1(_0395_),
    .B1(_0400_),
    .X(_0401_));
 sg13g2_a21oi_1 _4111_ (.A1(_0393_),
    .A2(_0401_),
    .Y(_0402_),
    .B1(_0391_));
 sg13g2_xor2_1 _4112_ (.B(_0386_),
    .A(_0384_),
    .X(_0403_));
 sg13g2_nor2b_1 _4113_ (.A(_0402_),
    .B_N(_0403_),
    .Y(_0404_));
 sg13g2_a21o_1 _4114_ (.A2(_0386_),
    .A1(_0384_),
    .B1(_0404_),
    .X(_0405_));
 sg13g2_a21oi_1 _4115_ (.A1(_0380_),
    .A2(_0405_),
    .Y(_0406_),
    .B1(_0379_));
 sg13g2_xor2_1 _4116_ (.B(_0374_),
    .A(_0372_),
    .X(_0407_));
 sg13g2_nor2b_1 _4117_ (.A(_0406_),
    .B_N(_0407_),
    .Y(_0408_));
 sg13g2_a21o_1 _4118_ (.A2(_0374_),
    .A1(_0372_),
    .B1(_0408_),
    .X(_0409_));
 sg13g2_xor2_1 _4119_ (.B(_0367_),
    .A(_0365_),
    .X(_0410_));
 sg13g2_a21oi_1 _4120_ (.A1(_0409_),
    .A2(_0410_),
    .Y(_0411_),
    .B1(_0368_));
 sg13g2_xor2_1 _4121_ (.B(_0363_),
    .A(_0361_),
    .X(_0412_));
 sg13g2_nand2b_1 _4122_ (.Y(_0413_),
    .B(_0412_),
    .A_N(_0411_));
 sg13g2_o21ai_1 _4123_ (.B1(_0413_),
    .Y(_0414_),
    .A1(_0361_),
    .A2(_0363_));
 sg13g2_xor2_1 _4124_ (.B(_0414_),
    .A(_0358_),
    .X(\main.demo._d___pip_58_1_1___stage___block_3_a[1] ));
 sg13g2_inv_2 _4125_ (.Y(_0415_),
    .A(net339));
 sg13g2_nand2_1 _4126_ (.Y(\main.demo._t___pip_58_1_3___block_87_atten_l[1] ),
    .A(net551),
    .B(net399));
 sg13g2_a21oi_2 _4127_ (.B1(\main.demo._d___pip_58_1_3___stage___block_3_cx[10] ),
    .Y(_0416_),
    .A2(\main.demo._d___pip_58_1_3___stage___block_3_cx[8] ),
    .A1(net425));
 sg13g2_a21o_2 _4128_ (.A2(\main.demo._d___pip_58_1_3___stage___block_3_cx[8] ),
    .A1(net425),
    .B1(\main.demo._d___pip_58_1_3___stage___block_3_cx[10] ),
    .X(_0417_));
 sg13g2_and2_1 _4129_ (.A(\main.demo._d___pip_58_1_3___stage___block_3_cx[6] ),
    .B(net427),
    .X(_0418_));
 sg13g2_nand2_2 _4130_ (.Y(_0419_),
    .A(\main.demo._d___pip_58_1_3___stage___block_3_cx[6] ),
    .B(net427));
 sg13g2_nor2_1 _4131_ (.A(\main.demo._d___pip_58_1_3___stage___block_3_cx[7] ),
    .B(\main.demo._d___pip_58_1_3___stage___block_3_cx[10] ),
    .Y(_0420_));
 sg13g2_or2_1 _4132_ (.X(_0421_),
    .B(\main.demo._d___pip_58_1_3___stage___block_3_cx[10] ),
    .A(\main.demo._d___pip_58_1_3___stage___block_3_cx[7] ));
 sg13g2_a21oi_2 _4133_ (.B1(_0416_),
    .Y(_0422_),
    .A2(_0420_),
    .A1(_0419_));
 sg13g2_o21ai_1 _4134_ (.B1(_0417_),
    .Y(_0423_),
    .A1(_0418_),
    .A2(_0421_));
 sg13g2_nand2_2 _4135_ (.Y(_0424_),
    .A(net426),
    .B(_0423_));
 sg13g2_nand2_2 _4136_ (.Y(_0425_),
    .A(\main.demo._d___pip_58_1_3___stage___block_3_cx[7] ),
    .B(_0416_));
 sg13g2_nand2_1 _4137_ (.Y(_0426_),
    .A(_0416_),
    .B(_0418_));
 sg13g2_nor3_2 _4138_ (.A(_2620_),
    .B(_0417_),
    .C(_0419_),
    .Y(_0427_));
 sg13g2_nand3_1 _4139_ (.B(_0416_),
    .C(_0418_),
    .A(\main.demo._d___pip_58_1_3___stage___block_3_cx[7] ),
    .Y(_0428_));
 sg13g2_a21oi_2 _4140_ (.B1(_0428_),
    .Y(_0429_),
    .A2(_0423_),
    .A1(net426));
 sg13g2_o21ai_1 _4141_ (.B1(_0427_),
    .Y(_0430_),
    .A1(_2646_),
    .A2(_0422_));
 sg13g2_nor3_2 _4142_ (.A(_2646_),
    .B(_0422_),
    .C(_0427_),
    .Y(_0431_));
 sg13g2_nand3_1 _4143_ (.B(_0423_),
    .C(_0428_),
    .A(net426),
    .Y(_0432_));
 sg13g2_nand2_1 _4144_ (.Y(_0433_),
    .A(_0430_),
    .B(_0432_));
 sg13g2_nand2_1 _4145_ (.Y(_0434_),
    .A(_0425_),
    .B(_0426_));
 sg13g2_nand2_1 _4146_ (.Y(_0435_),
    .A(_0428_),
    .B(_0434_));
 sg13g2_a21oi_2 _4147_ (.B1(\main.demo._d___pip_58_1_3___stage___block_3_cx[6] ),
    .Y(_0436_),
    .A2(_0421_),
    .A1(_0417_));
 sg13g2_nor2b_1 _4148_ (.A(\main.demo._d___pip_58_1_3___stage___block_3_cx[5] ),
    .B_N(_0436_),
    .Y(_0437_));
 sg13g2_nand2b_2 _4149_ (.Y(_0438_),
    .B(_0436_),
    .A_N(net427));
 sg13g2_a221oi_1 _4150_ (.B2(_0428_),
    .C1(_0438_),
    .B1(_0434_),
    .A1(_0430_),
    .Y(_0439_),
    .A2(_0432_));
 sg13g2_nand3_1 _4151_ (.B(_0435_),
    .C(_0437_),
    .A(_0433_),
    .Y(_0440_));
 sg13g2_nor2_2 _4152_ (.A(_2650_),
    .B(\main.demo._d___pip_58_1_3___stage___block_3_cx[5] ),
    .Y(_0441_));
 sg13g2_nor2_2 _4153_ (.A(_0422_),
    .B(_0441_),
    .Y(_0442_));
 sg13g2_inv_1 _4154_ (.Y(_0443_),
    .A(_0442_));
 sg13g2_a221oi_1 _4155_ (.B2(_0428_),
    .C1(_0442_),
    .B1(_0434_),
    .A1(_0430_),
    .Y(_0444_),
    .A2(_0432_));
 sg13g2_nand3_1 _4156_ (.B(_0435_),
    .C(_0443_),
    .A(_0433_),
    .Y(_0445_));
 sg13g2_o21ai_1 _4157_ (.B1(_0425_),
    .Y(_0446_),
    .A1(_2646_),
    .A2(_0422_));
 sg13g2_nor2_1 _4158_ (.A(_0426_),
    .B(_0446_),
    .Y(_0447_));
 sg13g2_nor3_1 _4159_ (.A(_0439_),
    .B(_0444_),
    .C(_0447_),
    .Y(_0448_));
 sg13g2_nor2_2 _4160_ (.A(net396),
    .B(_0448_),
    .Y(_0449_));
 sg13g2_nand4_1 _4161_ (.B(net427),
    .C(_0423_),
    .A(_2650_),
    .Y(_0450_),
    .D(_0425_));
 sg13g2_a21oi_2 _4162_ (.B1(_0450_),
    .Y(_0451_),
    .A2(_0432_),
    .A1(_0430_));
 sg13g2_nor2_2 _4163_ (.A(net393),
    .B(_0430_),
    .Y(_0452_));
 sg13g2_xnor2_1 _4164_ (.Y(_0453_),
    .A(net398),
    .B(_0429_));
 sg13g2_nand2_1 _4165_ (.Y(_0454_),
    .A(_0451_),
    .B(_0453_));
 sg13g2_nor4_2 _4166_ (.A(net398),
    .B(_0429_),
    .C(_0431_),
    .Y(_0455_),
    .D(_0450_));
 sg13g2_nor3_1 _4167_ (.A(net398),
    .B(_0424_),
    .C(_0428_),
    .Y(_0456_));
 sg13g2_nand4_1 _4168_ (.B(net393),
    .C(_0423_),
    .A(net426),
    .Y(_0457_),
    .D(_0427_));
 sg13g2_nor2_2 _4169_ (.A(_0438_),
    .B(_0446_),
    .Y(_0458_));
 sg13g2_nor3_1 _4170_ (.A(net398),
    .B(_0438_),
    .C(_0446_),
    .Y(_0459_));
 sg13g2_nand2_1 _4171_ (.Y(_0460_),
    .A(net394),
    .B(_0458_));
 sg13g2_nor3_2 _4172_ (.A(_0455_),
    .B(_0456_),
    .C(_0459_),
    .Y(_0461_));
 sg13g2_nor3_2 _4173_ (.A(_2620_),
    .B(_2646_),
    .C(_0417_),
    .Y(_0462_));
 sg13g2_nand4_1 _4174_ (.B(net393),
    .C(_0436_),
    .A(net427),
    .Y(_0463_),
    .D(_0462_));
 sg13g2_nand4_1 _4175_ (.B(net426),
    .C(_0416_),
    .A(_2620_),
    .Y(_0464_),
    .D(_0418_));
 sg13g2_nor2_1 _4176_ (.A(net395),
    .B(_0464_),
    .Y(_0465_));
 sg13g2_nor4_2 _4177_ (.A(_2620_),
    .B(net398),
    .C(_0424_),
    .Y(_0466_),
    .D(_0438_));
 sg13g2_nand2_2 _4178_ (.Y(_0467_),
    .A(_0441_),
    .B(_0462_));
 sg13g2_nor2_1 _4179_ (.A(net397),
    .B(_0467_),
    .Y(_0468_));
 sg13g2_nor3_2 _4180_ (.A(net397),
    .B(_0442_),
    .C(_0446_),
    .Y(_0469_));
 sg13g2_o21ai_1 _4181_ (.B1(_0463_),
    .Y(_0470_),
    .A1(net395),
    .A2(_0467_));
 sg13g2_nor2_1 _4182_ (.A(_0466_),
    .B(_0470_),
    .Y(_0471_));
 sg13g2_nor4_2 _4183_ (.A(_0465_),
    .B(_0466_),
    .C(_0469_),
    .Y(_0472_),
    .D(_0470_));
 sg13g2_nand3_1 _4184_ (.B(_0461_),
    .C(_0472_),
    .A(_0454_),
    .Y(_0473_));
 sg13g2_nor2_1 _4185_ (.A(_0449_),
    .B(_0473_),
    .Y(_0474_));
 sg13g2_a221oi_1 _4186_ (.B2(_0426_),
    .C1(_0427_),
    .B1(_0425_),
    .A1(net426),
    .Y(_0475_),
    .A2(_0423_));
 sg13g2_and3_1 _4187_ (.X(_0476_),
    .A(net395),
    .B(_0441_),
    .C(_0475_));
 sg13g2_nand3_1 _4188_ (.B(_0441_),
    .C(_0475_),
    .A(net395),
    .Y(_0477_));
 sg13g2_nor2_1 _4189_ (.A(_0452_),
    .B(_0476_),
    .Y(_0478_));
 sg13g2_and3_1 _4190_ (.X(_0479_),
    .A(_2650_),
    .B(net398),
    .C(_0475_));
 sg13g2_nor4_1 _4191_ (.A(_0452_),
    .B(_0462_),
    .C(_0476_),
    .D(_0479_),
    .Y(_0480_));
 sg13g2_nor4_2 _4192_ (.A(net393),
    .B(_0429_),
    .C(_0431_),
    .Y(_0481_),
    .D(_0450_));
 sg13g2_nor3_2 _4193_ (.A(net393),
    .B(_0442_),
    .C(_0446_),
    .Y(_0482_));
 sg13g2_nor2_2 _4194_ (.A(_0481_),
    .B(_0482_),
    .Y(_0483_));
 sg13g2_nor3_2 _4195_ (.A(net393),
    .B(_0419_),
    .C(_0446_),
    .Y(_0484_));
 sg13g2_nand2_1 _4196_ (.Y(_0485_),
    .A(net396),
    .B(_0458_));
 sg13g2_nor2_2 _4197_ (.A(\main.demo._t___pip_58_1_3___block_87_atten_l[1] ),
    .B(_0428_),
    .Y(_0486_));
 sg13g2_a21oi_2 _4198_ (.B1(_0481_),
    .Y(_0487_),
    .A2(_0458_),
    .A1(net396));
 sg13g2_nor2_2 _4199_ (.A(_0482_),
    .B(_0484_),
    .Y(_0488_));
 sg13g2_nand3b_1 _4200_ (.B(_0487_),
    .C(_0488_),
    .Y(_0489_),
    .A_N(_0486_));
 sg13g2_nand3_1 _4201_ (.B(_0487_),
    .C(_0488_),
    .A(_0480_),
    .Y(_0490_));
 sg13g2_nand2_2 _4202_ (.Y(_0491_),
    .A(net396),
    .B(_0451_));
 sg13g2_inv_1 _4203_ (.Y(_0492_),
    .A(_0491_));
 sg13g2_nand2_2 _4204_ (.Y(_0493_),
    .A(net396),
    .B(_0444_));
 sg13g2_o21ai_1 _4205_ (.B1(net396),
    .Y(_0494_),
    .A1(_0444_),
    .A2(_0451_));
 sg13g2_nor2_1 _4206_ (.A(net394),
    .B(_0467_),
    .Y(_0495_));
 sg13g2_nand3_1 _4207_ (.B(_0441_),
    .C(_0462_),
    .A(net395),
    .Y(_0496_));
 sg13g2_nor2_2 _4208_ (.A(net394),
    .B(_0464_),
    .Y(_0497_));
 sg13g2_or2_1 _4209_ (.X(_0498_),
    .B(_0464_),
    .A(net393));
 sg13g2_nand3_1 _4210_ (.B(_0496_),
    .C(_0498_),
    .A(_0494_),
    .Y(_0499_));
 sg13g2_nor4_2 _4211_ (.A(_0449_),
    .B(_0473_),
    .C(_0490_),
    .Y(_0500_),
    .D(_0499_));
 sg13g2_or4_2 _4212_ (.A(_0449_),
    .B(_0473_),
    .C(_0490_),
    .D(_0499_),
    .X(_0501_));
 sg13g2_nand2_2 _4213_ (.Y(_0502_),
    .A(net427),
    .B(_0479_));
 sg13g2_nand2_1 _4214_ (.Y(_0503_),
    .A(_0477_),
    .B(_0502_));
 sg13g2_nand2_2 _4215_ (.Y(_0504_),
    .A(_0478_),
    .B(_0502_));
 sg13g2_nor2_1 _4216_ (.A(_0456_),
    .B(_0469_),
    .Y(_0505_));
 sg13g2_nor4_2 _4217_ (.A(_2620_),
    .B(net393),
    .C(_0424_),
    .Y(_0506_),
    .D(_0438_));
 sg13g2_nor2_1 _4218_ (.A(_0484_),
    .B(_0506_),
    .Y(_0507_));
 sg13g2_nand3_1 _4219_ (.B(_0464_),
    .C(_0507_),
    .A(_0463_),
    .Y(_0508_));
 sg13g2_o21ai_1 _4220_ (.B1(_0505_),
    .Y(_0509_),
    .A1(net395),
    .A2(_0440_));
 sg13g2_nor4_2 _4221_ (.A(_0500_),
    .B(_0504_),
    .C(_0508_),
    .Y(_0510_),
    .D(_0509_));
 sg13g2_a22oi_1 _4222_ (.Y(_0511_),
    .B1(_0451_),
    .B2(_0453_),
    .A2(_0439_),
    .A1(net394));
 sg13g2_nor2_1 _4223_ (.A(net395),
    .B(_0445_),
    .Y(_0512_));
 sg13g2_nand2_1 _4224_ (.Y(_0513_),
    .A(net394),
    .B(_0444_));
 sg13g2_a221oi_1 _4225_ (.B2(_0453_),
    .C1(_0452_),
    .B1(_0451_),
    .A1(net394),
    .Y(_0514_),
    .A2(_0439_));
 sg13g2_nand2_1 _4226_ (.Y(_0515_),
    .A(_0513_),
    .B(_0514_));
 sg13g2_and4_2 _4227_ (.A(_0461_),
    .B(_0472_),
    .C(_0513_),
    .D(_0514_),
    .X(_0516_));
 sg13g2_and2_2 _4228_ (.A(\main.demo._d___pip_58_1_3___stage___block_3_cx[9] ),
    .B(_0516_),
    .X(_0517_));
 sg13g2_nand2_2 _4229_ (.Y(_0518_),
    .A(net425),
    .B(_0516_));
 sg13g2_or2_2 _4230_ (.X(_0519_),
    .B(_0453_),
    .A(_0440_));
 sg13g2_nand2_1 _4231_ (.Y(_0520_),
    .A(_0491_),
    .B(_0519_));
 sg13g2_nand2_1 _4232_ (.Y(_0521_),
    .A(_0437_),
    .B(_0475_));
 sg13g2_nor2_1 _4233_ (.A(net394),
    .B(_0521_),
    .Y(_0522_));
 sg13g2_or4_1 _4234_ (.A(_0455_),
    .B(_0503_),
    .C(_0512_),
    .D(_0522_),
    .X(_0523_));
 sg13g2_nor2_1 _4235_ (.A(_0465_),
    .B(_0466_),
    .Y(_0524_));
 sg13g2_nand2_1 _4236_ (.Y(_0525_),
    .A(_0463_),
    .B(_0524_));
 sg13g2_nand4_1 _4237_ (.B(net398),
    .C(_0436_),
    .A(net427),
    .Y(_0526_),
    .D(_0462_));
 sg13g2_and2_1 _4238_ (.A(_0498_),
    .B(_0526_),
    .X(_0527_));
 sg13g2_nand3_1 _4239_ (.B(_0485_),
    .C(_0527_),
    .A(_0457_),
    .Y(_0528_));
 sg13g2_or2_1 _4240_ (.X(_0529_),
    .B(_0528_),
    .A(_0525_));
 sg13g2_nor4_2 _4241_ (.A(_0517_),
    .B(_0520_),
    .C(_0523_),
    .Y(_0530_),
    .D(_0529_));
 sg13g2_nand2_2 _4242_ (.Y(_0531_),
    .A(_0494_),
    .B(_0501_));
 sg13g2_nor2_1 _4243_ (.A(_0495_),
    .B(_0506_),
    .Y(_0532_));
 sg13g2_nand3_1 _4244_ (.B(_0472_),
    .C(_0532_),
    .A(_0460_),
    .Y(_0533_));
 sg13g2_nor3_2 _4245_ (.A(_0481_),
    .B(_0504_),
    .C(_0533_),
    .Y(_0534_));
 sg13g2_nor2b_1 _4246_ (.A(_0531_),
    .B_N(_0534_),
    .Y(_0535_));
 sg13g2_nand3_1 _4247_ (.B(_0501_),
    .C(_0534_),
    .A(_0494_),
    .Y(_0536_));
 sg13g2_a221oi_1 _4248_ (.B2(_0441_),
    .C1(_0452_),
    .B1(_0462_),
    .A1(_0451_),
    .Y(_0537_),
    .A2(_0453_));
 sg13g2_nor2_1 _4249_ (.A(_0452_),
    .B(_0468_),
    .Y(_0538_));
 sg13g2_nand4_1 _4250_ (.B(_0505_),
    .C(_0527_),
    .A(_0487_),
    .Y(_0539_),
    .D(_0537_));
 sg13g2_a21oi_1 _4251_ (.A1(net425),
    .A2(_0516_),
    .Y(_0540_),
    .B1(_0539_));
 sg13g2_nor2_1 _4252_ (.A(_0486_),
    .B(_0506_),
    .Y(_0541_));
 sg13g2_nand4_1 _4253_ (.B(_0460_),
    .C(_0483_),
    .A(_0457_),
    .Y(_0542_),
    .D(_0541_));
 sg13g2_nor3_1 _4254_ (.A(_0449_),
    .B(_0495_),
    .C(_0542_),
    .Y(_0543_));
 sg13g2_and2_1 _4255_ (.A(_0501_),
    .B(_0543_),
    .X(_0544_));
 sg13g2_nor2b_1 _4256_ (.A(_0540_),
    .B_N(_0544_),
    .Y(_0545_));
 sg13g2_nand3_1 _4257_ (.B(_0540_),
    .C(_0543_),
    .A(_0501_),
    .Y(_0546_));
 sg13g2_a21o_1 _4258_ (.A2(_0543_),
    .A1(_0501_),
    .B1(_0540_),
    .X(_0547_));
 sg13g2_a22oi_1 _4259_ (.Y(_0548_),
    .B1(_0546_),
    .B2(_0547_),
    .A2(_0536_),
    .A1(_0530_));
 sg13g2_nand4_1 _4260_ (.B(_0536_),
    .C(_0546_),
    .A(_0530_),
    .Y(_0549_),
    .D(_0547_));
 sg13g2_nor2b_2 _4261_ (.A(_0548_),
    .B_N(_0549_),
    .Y(_0550_));
 sg13g2_and2_1 _4262_ (.A(_2651_),
    .B(_0550_),
    .X(_0551_));
 sg13g2_xnor2_1 _4263_ (.Y(_0552_),
    .A(_0530_),
    .B(_0536_));
 sg13g2_and2_1 _4264_ (.A(_2652_),
    .B(_0552_),
    .X(_0553_));
 sg13g2_nand2_1 _4265_ (.Y(_0554_),
    .A(_0551_),
    .B(_0553_));
 sg13g2_xnor2_1 _4266_ (.Y(_0555_),
    .A(_0551_),
    .B(_0553_));
 sg13g2_a21oi_1 _4267_ (.A1(net395),
    .A2(_0444_),
    .Y(_0556_),
    .B1(_0497_));
 sg13g2_and3_1 _4268_ (.X(_0557_),
    .A(_0478_),
    .B(_0501_),
    .C(_0556_));
 sg13g2_nand2b_2 _4269_ (.Y(_0558_),
    .B(_0526_),
    .A_N(_0465_));
 sg13g2_inv_1 _4270_ (.Y(_0559_),
    .A(_0558_));
 sg13g2_nor4_1 _4271_ (.A(_0484_),
    .B(_0506_),
    .C(_0522_),
    .D(_0558_),
    .Y(_0560_));
 sg13g2_nand4_1 _4272_ (.B(_0487_),
    .C(_0557_),
    .A(_0471_),
    .Y(_0561_),
    .D(_0560_));
 sg13g2_nor2_1 _4273_ (.A(_0497_),
    .B(_0506_),
    .Y(_0562_));
 sg13g2_and2_1 _4274_ (.A(_0485_),
    .B(_0541_),
    .X(_0563_));
 sg13g2_nand3_1 _4275_ (.B(_0488_),
    .C(_0562_),
    .A(_0445_),
    .Y(_0564_));
 sg13g2_nor3_1 _4276_ (.A(_0503_),
    .B(_0525_),
    .C(_0564_),
    .Y(_0565_));
 sg13g2_nand4_1 _4277_ (.B(_0518_),
    .C(_0563_),
    .A(_0491_),
    .Y(_0566_),
    .D(_0565_));
 sg13g2_nor2b_1 _4278_ (.A(_0561_),
    .B_N(_0566_),
    .Y(_0567_));
 sg13g2_xor2_1 _4279_ (.B(_0566_),
    .A(_0561_),
    .X(_0568_));
 sg13g2_nand4_1 _4280_ (.B(_0502_),
    .C(_0532_),
    .A(_0457_),
    .Y(_0569_),
    .D(_0538_));
 sg13g2_nand2_1 _4281_ (.Y(_0570_),
    .A(_0440_),
    .B(_0483_));
 sg13g2_or4_1 _4282_ (.A(_0458_),
    .B(_0512_),
    .C(_0569_),
    .D(_0570_),
    .X(_0571_));
 sg13g2_nor3_2 _4283_ (.A(_0517_),
    .B(_0558_),
    .C(_0571_),
    .Y(_0572_));
 sg13g2_nor3_1 _4284_ (.A(_0466_),
    .B(_0484_),
    .C(_0486_),
    .Y(_0573_));
 sg13g2_nand4_1 _4285_ (.B(_0477_),
    .C(_0559_),
    .A(_0461_),
    .Y(_0574_),
    .D(_0573_));
 sg13g2_nand3_1 _4286_ (.B(_0496_),
    .C(_0511_),
    .A(_0483_),
    .Y(_0575_));
 sg13g2_nor4_2 _4287_ (.A(_0492_),
    .B(_0500_),
    .C(_0574_),
    .Y(_0576_),
    .D(_0575_));
 sg13g2_inv_1 _4288_ (.Y(_0577_),
    .A(_0576_));
 sg13g2_nor2_1 _4289_ (.A(_0466_),
    .B(_0482_),
    .Y(_0578_));
 sg13g2_nand3_1 _4290_ (.B(_0556_),
    .C(_0578_),
    .A(_0538_),
    .Y(_0579_));
 sg13g2_or3_1 _4291_ (.A(_0517_),
    .B(_0523_),
    .C(_0579_),
    .X(_0580_));
 sg13g2_nand2_1 _4292_ (.Y(_0581_),
    .A(_0510_),
    .B(_0580_));
 sg13g2_xor2_1 _4293_ (.B(_0580_),
    .A(_0510_),
    .X(_0582_));
 sg13g2_o21ai_1 _4294_ (.B1(_0582_),
    .Y(_0583_),
    .A1(_0545_),
    .A2(_0548_));
 sg13g2_nand2b_1 _4295_ (.Y(_0584_),
    .B(_0576_),
    .A_N(_0572_));
 sg13g2_and2_1 _4296_ (.A(_0581_),
    .B(_0584_),
    .X(_0585_));
 sg13g2_a22oi_1 _4297_ (.Y(_0586_),
    .B1(_0583_),
    .B2(_0585_),
    .A2(_0577_),
    .A1(_0572_));
 sg13g2_a221oi_1 _4298_ (.B2(_0585_),
    .C1(_0568_),
    .B1(_0583_),
    .A1(_0572_),
    .Y(_0587_),
    .A2(_0577_));
 sg13g2_xnor2_1 _4299_ (.Y(_0588_),
    .A(_0568_),
    .B(_0586_));
 sg13g2_xor2_1 _4300_ (.B(_0586_),
    .A(_0568_),
    .X(_0589_));
 sg13g2_and2_1 _4301_ (.A(\main.demo._d___pip_58_1_3___stage___block_3_cx[0] ),
    .B(_0588_),
    .X(_0590_));
 sg13g2_xor2_1 _4302_ (.B(_0576_),
    .A(_0572_),
    .X(_0591_));
 sg13g2_nand3_1 _4303_ (.B(_0583_),
    .C(_0591_),
    .A(_0581_),
    .Y(_0592_));
 sg13g2_a21o_1 _4304_ (.A2(_0583_),
    .A1(_0581_),
    .B1(_0591_),
    .X(_0593_));
 sg13g2_nand2_1 _4305_ (.Y(_0594_),
    .A(_0592_),
    .B(_0593_));
 sg13g2_and2_2 _4306_ (.A(_0592_),
    .B(_0593_),
    .X(_0595_));
 sg13g2_or3_1 _4307_ (.A(_0545_),
    .B(_0548_),
    .C(_0582_),
    .X(_0596_));
 sg13g2_and2_2 _4308_ (.A(_0583_),
    .B(_0596_),
    .X(_0597_));
 sg13g2_nand2_1 _4309_ (.Y(_0598_),
    .A(\main.demo._d___pip_58_1_3___stage___block_3_cx[2] ),
    .B(_0597_));
 sg13g2_nand3_1 _4310_ (.B(_0592_),
    .C(_0593_),
    .A(net428),
    .Y(_0599_));
 sg13g2_xor2_1 _4311_ (.B(_0599_),
    .A(_0598_),
    .X(_0600_));
 sg13g2_nand2_1 _4312_ (.Y(_0601_),
    .A(_0590_),
    .B(_0600_));
 sg13g2_xor2_1 _4313_ (.B(_0600_),
    .A(_0590_),
    .X(_0602_));
 sg13g2_nand2b_1 _4314_ (.Y(_0603_),
    .B(_0602_),
    .A_N(_0555_));
 sg13g2_nand4_1 _4315_ (.B(_0483_),
    .C(_0526_),
    .A(_0477_),
    .Y(_0604_),
    .D(_0541_));
 sg13g2_nor3_2 _4316_ (.A(_0515_),
    .B(_0531_),
    .C(_0604_),
    .Y(_0605_));
 sg13g2_nand4_1 _4317_ (.B(_0496_),
    .C(_0511_),
    .A(_0487_),
    .Y(_0606_),
    .D(_0562_));
 sg13g2_nor2_1 _4318_ (.A(_0504_),
    .B(_0606_),
    .Y(_0607_));
 sg13g2_nand4_1 _4319_ (.B(_0518_),
    .C(_0519_),
    .A(_0491_),
    .Y(_0608_),
    .D(_0607_));
 sg13g2_nand2_1 _4320_ (.Y(_0609_),
    .A(_0605_),
    .B(_0608_));
 sg13g2_xor2_1 _4321_ (.B(_0608_),
    .A(_0605_),
    .X(_0610_));
 sg13g2_o21ai_1 _4322_ (.B1(_0610_),
    .Y(_0611_),
    .A1(_0567_),
    .A2(_0587_));
 sg13g2_or3_1 _4323_ (.A(_0567_),
    .B(_0587_),
    .C(_0610_),
    .X(_0612_));
 sg13g2_and2_1 _4324_ (.A(_0611_),
    .B(_0612_),
    .X(_0613_));
 sg13g2_nand3_1 _4325_ (.B(_0611_),
    .C(_0612_),
    .A(_2654_),
    .Y(_0614_));
 sg13g2_and4_1 _4326_ (.A(\main.demo._d___pip_58_1_3___stage___block_3_cx[2] ),
    .B(_2653_),
    .C(_0588_),
    .D(_0595_),
    .X(_0615_));
 sg13g2_a22oi_1 _4327_ (.Y(_0616_),
    .B1(_0595_),
    .B2(\main.demo._d___pip_58_1_3___stage___block_3_cx[2] ),
    .A2(_0588_),
    .A1(_2653_));
 sg13g2_or3_1 _4328_ (.A(_0614_),
    .B(_0615_),
    .C(_0616_),
    .X(_0617_));
 sg13g2_o21ai_1 _4329_ (.B1(_0614_),
    .Y(_0618_),
    .A1(_0615_),
    .A2(_0616_));
 sg13g2_and2_1 _4330_ (.A(_2651_),
    .B(_0597_),
    .X(_0619_));
 sg13g2_nand2_1 _4331_ (.Y(_0620_),
    .A(_2651_),
    .B(_0597_));
 sg13g2_and2_1 _4332_ (.A(_2652_),
    .B(_0550_),
    .X(_0621_));
 sg13g2_nand2_1 _4333_ (.Y(_0622_),
    .A(_0619_),
    .B(_0621_));
 sg13g2_xnor2_1 _4334_ (.Y(_0623_),
    .A(_0620_),
    .B(_0621_));
 sg13g2_nor2b_1 _4335_ (.A(_0554_),
    .B_N(_0623_),
    .Y(_0624_));
 sg13g2_nor2_1 _4336_ (.A(_0009_),
    .B(_0594_),
    .Y(_0625_));
 sg13g2_nand2_1 _4337_ (.Y(_0626_),
    .A(_2652_),
    .B(_0595_));
 sg13g2_nor2_1 _4338_ (.A(_0620_),
    .B(_0626_),
    .Y(_0627_));
 sg13g2_a22oi_1 _4339_ (.Y(_0628_),
    .B1(_0597_),
    .B2(_2652_),
    .A2(_0595_),
    .A1(_2651_));
 sg13g2_a21oi_1 _4340_ (.A1(_0619_),
    .A2(_0625_),
    .Y(_0629_),
    .B1(_0628_));
 sg13g2_xnor2_1 _4341_ (.Y(_0630_),
    .A(_0554_),
    .B(_0623_));
 sg13g2_and3_1 _4342_ (.X(_0631_),
    .A(_0617_),
    .B(_0618_),
    .C(_0630_));
 sg13g2_a21oi_2 _4343_ (.B1(_0630_),
    .Y(_0632_),
    .A2(_0618_),
    .A1(_0617_));
 sg13g2_nor3_1 _4344_ (.A(_0603_),
    .B(_0631_),
    .C(_0632_),
    .Y(_0633_));
 sg13g2_or3_1 _4345_ (.A(_0603_),
    .B(_0631_),
    .C(_0632_),
    .X(_0634_));
 sg13g2_o21ai_1 _4346_ (.B1(_0601_),
    .Y(_0635_),
    .A1(_0598_),
    .A2(_0599_));
 sg13g2_o21ai_1 _4347_ (.B1(_0603_),
    .Y(_0636_),
    .A1(_0631_),
    .A2(_0632_));
 sg13g2_and3_1 _4348_ (.X(_0637_),
    .A(_0634_),
    .B(_0635_),
    .C(_0636_));
 sg13g2_nor2_1 _4349_ (.A(_0633_),
    .B(_0637_),
    .Y(_0638_));
 sg13g2_nor2b_1 _4350_ (.A(_0615_),
    .B_N(_0617_),
    .Y(_0639_));
 sg13g2_nor2_1 _4351_ (.A(_0624_),
    .B(_0631_),
    .Y(_0640_));
 sg13g2_nor2b_1 _4352_ (.A(_0622_),
    .B_N(_0629_),
    .Y(_0641_));
 sg13g2_xor2_1 _4353_ (.B(_0629_),
    .A(_0622_),
    .X(_0642_));
 sg13g2_nand3_1 _4354_ (.B(_0557_),
    .C(_0563_),
    .A(_0474_),
    .Y(_0643_));
 sg13g2_nor4_1 _4355_ (.A(net425),
    .B(_0486_),
    .C(_0499_),
    .D(_0503_),
    .Y(_0644_));
 sg13g2_and2_1 _4356_ (.A(_0516_),
    .B(_0644_),
    .X(_0645_));
 sg13g2_or2_1 _4357_ (.X(_0646_),
    .B(_0645_),
    .A(_0643_));
 sg13g2_xnor2_1 _4358_ (.Y(_0647_),
    .A(_0643_),
    .B(_0645_));
 sg13g2_a21o_1 _4359_ (.A2(_0611_),
    .A1(_0609_),
    .B1(_0647_),
    .X(_0648_));
 sg13g2_and2_1 _4360_ (.A(_0519_),
    .B(_0648_),
    .X(_0649_));
 sg13g2_nand3_1 _4361_ (.B(_0519_),
    .C(_0648_),
    .A(\main.demo._d___pip_58_1_3___stage___block_3_cx[0] ),
    .Y(_0650_));
 sg13g2_nor2_1 _4362_ (.A(_0011_),
    .B(_0589_),
    .Y(_0651_));
 sg13g2_and3_1 _4363_ (.X(_0652_),
    .A(net428),
    .B(_0611_),
    .C(_0612_));
 sg13g2_nand2_1 _4364_ (.Y(_0653_),
    .A(_0651_),
    .B(_0652_));
 sg13g2_xnor2_1 _4365_ (.Y(_0654_),
    .A(_0651_),
    .B(_0652_));
 sg13g2_xnor2_1 _4366_ (.Y(_0655_),
    .A(_0650_),
    .B(_0654_));
 sg13g2_nor2_1 _4367_ (.A(_0642_),
    .B(_0655_),
    .Y(_0656_));
 sg13g2_xnor2_1 _4368_ (.Y(_0657_),
    .A(_0642_),
    .B(_0655_));
 sg13g2_xor2_1 _4369_ (.B(_0657_),
    .A(_0640_),
    .X(_0658_));
 sg13g2_nand2b_1 _4370_ (.Y(_0659_),
    .B(_0658_),
    .A_N(_0639_));
 sg13g2_xnor2_1 _4371_ (.Y(_0660_),
    .A(_0639_),
    .B(_0658_));
 sg13g2_nand2b_1 _4372_ (.Y(_0661_),
    .B(_0660_),
    .A_N(_0638_));
 sg13g2_nor2_1 _4373_ (.A(_0012_),
    .B(_0594_),
    .Y(_0662_));
 sg13g2_and2_1 _4374_ (.A(\main.demo._d___pip_58_1_3___stage___block_3_cx[2] ),
    .B(_0550_),
    .X(_0663_));
 sg13g2_nand3_1 _4375_ (.B(_0597_),
    .C(_0663_),
    .A(\main.demo._d___pip_58_1_3___stage___block_3_cx[1] ),
    .Y(_0664_));
 sg13g2_a21o_1 _4376_ (.A2(_0597_),
    .A1(\main.demo._d___pip_58_1_3___stage___block_3_cx[1] ),
    .B1(_0663_),
    .X(_0665_));
 sg13g2_and2_1 _4377_ (.A(_0664_),
    .B(_0665_),
    .X(_0666_));
 sg13g2_nand2_1 _4378_ (.Y(_0667_),
    .A(_0662_),
    .B(_0666_));
 sg13g2_xnor2_1 _4379_ (.Y(_0668_),
    .A(_0662_),
    .B(_0666_));
 sg13g2_nand2_1 _4380_ (.Y(_0669_),
    .A(\main.demo._d___pip_58_1_3___stage___block_3_cx[3] ),
    .B(_0552_));
 sg13g2_nor2_1 _4381_ (.A(_0668_),
    .B(_0669_),
    .Y(_0670_));
 sg13g2_xnor2_1 _4382_ (.Y(_0671_),
    .A(_0555_),
    .B(_0602_));
 sg13g2_and2_1 _4383_ (.A(_0670_),
    .B(_0671_),
    .X(_0672_));
 sg13g2_nand2_1 _4384_ (.Y(_0673_),
    .A(_0664_),
    .B(_0667_));
 sg13g2_xor2_1 _4385_ (.B(_0671_),
    .A(_0670_),
    .X(_0674_));
 sg13g2_a21oi_1 _4386_ (.A1(_0673_),
    .A2(_0674_),
    .Y(_0675_),
    .B1(_0672_));
 sg13g2_a21oi_1 _4387_ (.A1(_0634_),
    .A2(_0636_),
    .Y(_0676_),
    .B1(_0635_));
 sg13g2_nor3_1 _4388_ (.A(_0637_),
    .B(_0675_),
    .C(_0676_),
    .Y(_0677_));
 sg13g2_nand2_1 _4389_ (.Y(_0678_),
    .A(\main.demo._d___pip_58_1_3___stage___block_3_cx[0] ),
    .B(_0597_));
 sg13g2_nand2_1 _4390_ (.Y(_0679_),
    .A(_2653_),
    .B(_0550_));
 sg13g2_nand2_1 _4391_ (.Y(_0680_),
    .A(_2654_),
    .B(_0552_));
 sg13g2_nor4_1 _4392_ (.A(_0011_),
    .B(_0678_),
    .C(_0679_),
    .D(_0680_),
    .Y(_0681_));
 sg13g2_nand2_1 _4393_ (.Y(_0682_),
    .A(_0668_),
    .B(_0669_));
 sg13g2_nand2b_1 _4394_ (.Y(_0683_),
    .B(_0552_),
    .A_N(_0011_));
 sg13g2_a21o_1 _4395_ (.A2(_0683_),
    .A1(_0680_),
    .B1(_0679_),
    .X(_0684_));
 sg13g2_a221oi_1 _4396_ (.B2(_0678_),
    .C1(_0670_),
    .B1(_0684_),
    .A1(_0679_),
    .Y(_0685_),
    .A2(_0683_));
 sg13g2_a21oi_1 _4397_ (.A1(_0682_),
    .A2(_0685_),
    .Y(_0686_),
    .B1(_0681_));
 sg13g2_xnor2_1 _4398_ (.Y(_0687_),
    .A(_0673_),
    .B(_0674_));
 sg13g2_nor2_1 _4399_ (.A(_0686_),
    .B(_0687_),
    .Y(_0688_));
 sg13g2_o21ai_1 _4400_ (.B1(_0675_),
    .Y(_0689_),
    .A1(_0637_),
    .A2(_0676_));
 sg13g2_nor2b_1 _4401_ (.A(_0677_),
    .B_N(_0689_),
    .Y(_0690_));
 sg13g2_a21oi_1 _4402_ (.A1(_0688_),
    .A2(_0689_),
    .Y(_0691_),
    .B1(_0677_));
 sg13g2_nor2b_1 _4403_ (.A(_0660_),
    .B_N(_0638_),
    .Y(_0692_));
 sg13g2_xnor2_1 _4404_ (.Y(_0693_),
    .A(_0638_),
    .B(_0660_));
 sg13g2_o21ai_1 _4405_ (.B1(_0661_),
    .Y(_0694_),
    .A1(_0691_),
    .A2(_0692_));
 sg13g2_o21ai_1 _4406_ (.B1(_0659_),
    .Y(_0695_),
    .A1(_0640_),
    .A2(_0657_));
 sg13g2_o21ai_1 _4407_ (.B1(_0653_),
    .Y(_0696_),
    .A1(_0650_),
    .A2(_0654_));
 sg13g2_nor2_1 _4408_ (.A(_0641_),
    .B(_0656_),
    .Y(_0697_));
 sg13g2_nor3_2 _4409_ (.A(_0492_),
    .B(_0497_),
    .C(_0500_),
    .Y(_0698_));
 sg13g2_nor2_1 _4410_ (.A(_0479_),
    .B(_0489_),
    .Y(_0699_));
 sg13g2_nand2_2 _4411_ (.Y(_0700_),
    .A(_0698_),
    .B(_0699_));
 sg13g2_nand4_1 _4412_ (.B(_0496_),
    .C(_0519_),
    .A(_0493_),
    .Y(_0701_),
    .D(_0521_));
 sg13g2_nor3_1 _4413_ (.A(_0489_),
    .B(_0517_),
    .C(_0701_),
    .Y(_0702_));
 sg13g2_xnor2_1 _4414_ (.Y(_0703_),
    .A(_0700_),
    .B(_0702_));
 sg13g2_a21o_1 _4415_ (.A2(_0648_),
    .A1(_0646_),
    .B1(_0703_),
    .X(_0704_));
 sg13g2_nand2_1 _4416_ (.Y(_0705_),
    .A(\main.demo._d___pip_58_1_3___stage___block_3_cx[0] ),
    .B(_0704_));
 sg13g2_and2_1 _4417_ (.A(_0493_),
    .B(net358),
    .X(_0706_));
 sg13g2_inv_1 _4418_ (.Y(_0707_),
    .A(_0706_));
 sg13g2_nand3_1 _4419_ (.B(_0493_),
    .C(_0704_),
    .A(\main.demo._d___pip_58_1_3___stage___block_3_cx[0] ),
    .Y(_0708_));
 sg13g2_nand3_1 _4420_ (.B(_0519_),
    .C(_0648_),
    .A(net428),
    .Y(_0709_));
 sg13g2_nor2b_1 _4421_ (.A(_0011_),
    .B_N(_0613_),
    .Y(_0710_));
 sg13g2_nand2b_1 _4422_ (.Y(_0711_),
    .B(_0710_),
    .A_N(_0709_));
 sg13g2_xnor2_1 _4423_ (.Y(_0712_),
    .A(_0709_),
    .B(_0710_));
 sg13g2_nand2b_1 _4424_ (.Y(_0713_),
    .B(_0712_),
    .A_N(_0708_));
 sg13g2_xnor2_1 _4425_ (.Y(_0714_),
    .A(_0708_),
    .B(_0712_));
 sg13g2_nand2_2 _4426_ (.Y(_0715_),
    .A(\main.demo._d___pip_58_1_3___stage___block_3_cx[3] ),
    .B(_0588_));
 sg13g2_nor2_1 _4427_ (.A(_0619_),
    .B(_0626_),
    .Y(_0716_));
 sg13g2_xnor2_1 _4428_ (.Y(_0717_),
    .A(_0715_),
    .B(_0716_));
 sg13g2_xnor2_1 _4429_ (.Y(_0718_),
    .A(_0714_),
    .B(_0717_));
 sg13g2_nor2_1 _4430_ (.A(_0697_),
    .B(_0718_),
    .Y(_0719_));
 sg13g2_xor2_1 _4431_ (.B(_0718_),
    .A(_0697_),
    .X(_0720_));
 sg13g2_xnor2_1 _4432_ (.Y(_0721_),
    .A(_0696_),
    .B(_0720_));
 sg13g2_nor2b_1 _4433_ (.A(_0721_),
    .B_N(_0695_),
    .Y(_0722_));
 sg13g2_nand2b_1 _4434_ (.Y(_0723_),
    .B(_0721_),
    .A_N(_0695_));
 sg13g2_xnor2_1 _4435_ (.Y(_0724_),
    .A(_0695_),
    .B(_0721_));
 sg13g2_xnor2_1 _4436_ (.Y(_0725_),
    .A(_0694_),
    .B(_0724_));
 sg13g2_or2_1 _4437_ (.X(_0726_),
    .B(_0725_),
    .A(_0510_));
 sg13g2_xnor2_1 _4438_ (.Y(_0727_),
    .A(_0691_),
    .B(_0693_));
 sg13g2_nor2b_1 _4439_ (.A(_0544_),
    .B_N(_0727_),
    .Y(_0728_));
 sg13g2_xnor2_1 _4440_ (.Y(_0729_),
    .A(_0688_),
    .B(_0690_));
 sg13g2_nor2_1 _4441_ (.A(_0535_),
    .B(_0729_),
    .Y(_0730_));
 sg13g2_xnor2_1 _4442_ (.Y(_0731_),
    .A(_0544_),
    .B(_0727_));
 sg13g2_a21oi_1 _4443_ (.A1(_0730_),
    .A2(_0731_),
    .Y(_0732_),
    .B1(_0728_));
 sg13g2_and2_1 _4444_ (.A(_0510_),
    .B(_0725_),
    .X(_0733_));
 sg13g2_xor2_1 _4445_ (.B(_0725_),
    .A(_0510_),
    .X(_0734_));
 sg13g2_o21ai_1 _4446_ (.B1(_0726_),
    .Y(_0735_),
    .A1(_0732_),
    .A2(_0733_));
 sg13g2_a21o_1 _4447_ (.A2(_0723_),
    .A1(_0694_),
    .B1(_0722_),
    .X(_0736_));
 sg13g2_a21oi_1 _4448_ (.A1(_0696_),
    .A2(_0720_),
    .Y(_0737_),
    .B1(_0719_));
 sg13g2_nand2_1 _4449_ (.Y(_0738_),
    .A(_0711_),
    .B(_0713_));
 sg13g2_a22oi_1 _4450_ (.Y(_0739_),
    .B1(_0717_),
    .B2(_0714_),
    .A2(_0715_),
    .A1(_0627_));
 sg13g2_or2_1 _4451_ (.X(_0740_),
    .B(_0715_),
    .A(_0626_));
 sg13g2_nand2_1 _4452_ (.Y(_0741_),
    .A(_2651_),
    .B(_0613_));
 sg13g2_nor2_1 _4453_ (.A(_0009_),
    .B(_0589_),
    .Y(_0742_));
 sg13g2_nand3_1 _4454_ (.B(_0613_),
    .C(_0742_),
    .A(_2651_),
    .Y(_0743_));
 sg13g2_xor2_1 _4455_ (.B(_0742_),
    .A(_0741_),
    .X(_0744_));
 sg13g2_nor2_1 _4456_ (.A(_0740_),
    .B(_0744_),
    .Y(_0745_));
 sg13g2_xor2_1 _4457_ (.B(_0744_),
    .A(_0740_),
    .X(_0746_));
 sg13g2_and2_2 _4458_ (.A(_0491_),
    .B(net358),
    .X(_0747_));
 sg13g2_nand2_1 _4459_ (.Y(_0748_),
    .A(\main.demo._d___pip_58_1_3___stage___block_3_cx[0] ),
    .B(_0747_));
 sg13g2_nand2_1 _4460_ (.Y(_0749_),
    .A(\main.demo._d___pip_58_1_3___stage___block_3_cx[2] ),
    .B(net358));
 sg13g2_nand2_1 _4461_ (.Y(_0750_),
    .A(\main.demo._d___pip_58_1_3___stage___block_3_cx[2] ),
    .B(_0706_));
 sg13g2_nand2_1 _4462_ (.Y(_0751_),
    .A(\main.demo._d___pip_58_1_3___stage___block_3_cx[2] ),
    .B(_0649_));
 sg13g2_nand2_1 _4463_ (.Y(_0752_),
    .A(net428),
    .B(net358));
 sg13g2_nand3_1 _4464_ (.B(_0493_),
    .C(net358),
    .A(net428),
    .Y(_0753_));
 sg13g2_xor2_1 _4465_ (.B(_0753_),
    .A(_0751_),
    .X(_0754_));
 sg13g2_nand2b_1 _4466_ (.Y(_0755_),
    .B(_0754_),
    .A_N(_0748_));
 sg13g2_xnor2_1 _4467_ (.Y(_0756_),
    .A(_0748_),
    .B(_0754_));
 sg13g2_xnor2_1 _4468_ (.Y(_0757_),
    .A(_0746_),
    .B(_0756_));
 sg13g2_nor2_1 _4469_ (.A(_0739_),
    .B(_0757_),
    .Y(_0758_));
 sg13g2_xor2_1 _4470_ (.B(_0757_),
    .A(_0739_),
    .X(_0759_));
 sg13g2_xnor2_1 _4471_ (.Y(_0760_),
    .A(_0738_),
    .B(_0759_));
 sg13g2_nor2_1 _4472_ (.A(_0737_),
    .B(_0760_),
    .Y(_0761_));
 sg13g2_xor2_1 _4473_ (.B(_0760_),
    .A(_0737_),
    .X(_0762_));
 sg13g2_xnor2_1 _4474_ (.Y(_0763_),
    .A(_0736_),
    .B(_0762_));
 sg13g2_nor2_1 _4475_ (.A(_0576_),
    .B(_0763_),
    .Y(_0764_));
 sg13g2_xnor2_1 _4476_ (.Y(_0765_),
    .A(_0577_),
    .B(_0763_));
 sg13g2_xor2_1 _4477_ (.B(_0765_),
    .A(_0735_),
    .X(_0766_));
 sg13g2_nand2b_1 _4478_ (.Y(_0767_),
    .B(_0766_),
    .A_N(_0016_));
 sg13g2_xnor2_1 _4479_ (.Y(_0768_),
    .A(_0732_),
    .B(_0734_));
 sg13g2_nand2_1 _4480_ (.Y(_0769_),
    .A(\main.demo._q_speed[0] ),
    .B(_0768_));
 sg13g2_nor2b_1 _4481_ (.A(_0766_),
    .B_N(_0016_),
    .Y(_0770_));
 sg13g2_xnor2_1 _4482_ (.Y(_0771_),
    .A(_0016_),
    .B(_0766_));
 sg13g2_o21ai_1 _4483_ (.B1(_0767_),
    .Y(_0772_),
    .A1(_0769_),
    .A2(_0770_));
 sg13g2_a21oi_1 _4484_ (.A1(_0735_),
    .A2(_0765_),
    .Y(_0773_),
    .B1(_0764_));
 sg13g2_a21oi_1 _4485_ (.A1(_0736_),
    .A2(_0762_),
    .Y(_0774_),
    .B1(_0761_));
 sg13g2_a21oi_1 _4486_ (.A1(_0738_),
    .A2(_0759_),
    .Y(_0775_),
    .B1(_0758_));
 sg13g2_o21ai_1 _4487_ (.B1(_0755_),
    .Y(_0776_),
    .A1(_0751_),
    .A2(_0753_));
 sg13g2_a21oi_1 _4488_ (.A1(_0746_),
    .A2(_0756_),
    .Y(_0777_),
    .B1(_0745_));
 sg13g2_nand2_1 _4489_ (.Y(_0778_),
    .A(net428),
    .B(_0747_));
 sg13g2_nor2_1 _4490_ (.A(_0750_),
    .B(_0778_),
    .Y(_0779_));
 sg13g2_xor2_1 _4491_ (.B(_0778_),
    .A(_0750_),
    .X(_0780_));
 sg13g2_nor2b_1 _4492_ (.A(_0705_),
    .B_N(_0780_),
    .Y(_0781_));
 sg13g2_xnor2_1 _4493_ (.Y(_0782_),
    .A(_0705_),
    .B(_0780_));
 sg13g2_nand2_1 _4494_ (.Y(_0783_),
    .A(_2652_),
    .B(_0649_));
 sg13g2_nor2_1 _4495_ (.A(_0741_),
    .B(_0783_),
    .Y(_0784_));
 sg13g2_a22oi_1 _4496_ (.Y(_0785_),
    .B1(_0649_),
    .B2(_2651_),
    .A2(_0613_),
    .A1(_2652_));
 sg13g2_or2_1 _4497_ (.X(_0786_),
    .B(_0785_),
    .A(_0784_));
 sg13g2_nor2_1 _4498_ (.A(_0743_),
    .B(_0786_),
    .Y(_0787_));
 sg13g2_xor2_1 _4499_ (.B(_0786_),
    .A(_0743_),
    .X(_0788_));
 sg13g2_xnor2_1 _4500_ (.Y(_0789_),
    .A(_0782_),
    .B(_0788_));
 sg13g2_nor2_1 _4501_ (.A(_0777_),
    .B(_0789_),
    .Y(_0790_));
 sg13g2_xor2_1 _4502_ (.B(_0789_),
    .A(_0777_),
    .X(_0791_));
 sg13g2_xnor2_1 _4503_ (.Y(_0792_),
    .A(_0776_),
    .B(_0791_));
 sg13g2_or2_1 _4504_ (.X(_0793_),
    .B(_0792_),
    .A(_0775_));
 sg13g2_and2_1 _4505_ (.A(_0775_),
    .B(_0792_),
    .X(_0794_));
 sg13g2_xor2_1 _4506_ (.B(_0792_),
    .A(_0775_),
    .X(_0795_));
 sg13g2_xnor2_1 _4507_ (.Y(_0796_),
    .A(_0774_),
    .B(_0795_));
 sg13g2_nand2_1 _4508_ (.Y(_0797_),
    .A(_0561_),
    .B(_0796_));
 sg13g2_xnor2_1 _4509_ (.Y(_0798_),
    .A(_0561_),
    .B(_0796_));
 sg13g2_xnor2_1 _4510_ (.Y(_0799_),
    .A(_0773_),
    .B(_0798_));
 sg13g2_xnor2_1 _4511_ (.Y(_0800_),
    .A(\main.demo._q_speed[2] ),
    .B(_0799_));
 sg13g2_xor2_1 _4512_ (.B(_0800_),
    .A(_0772_),
    .X(_0801_));
 sg13g2_inv_2 _4513_ (.Y(_0802_),
    .A(_0801_));
 sg13g2_o21ai_1 _4514_ (.B1(_0793_),
    .Y(_0803_),
    .A1(_0774_),
    .A2(_0794_));
 sg13g2_a21oi_1 _4515_ (.A1(_0776_),
    .A2(_0791_),
    .Y(_0804_),
    .B1(_0790_));
 sg13g2_nor2_1 _4516_ (.A(_0779_),
    .B(_0781_),
    .Y(_0805_));
 sg13g2_a21oi_1 _4517_ (.A1(_0782_),
    .A2(_0788_),
    .Y(_0806_),
    .B1(_0787_));
 sg13g2_nand2_2 _4518_ (.Y(_0807_),
    .A(\main.demo._d___pip_58_1_3___stage___block_3_cx[0] ),
    .B(_0518_));
 sg13g2_inv_1 _4519_ (.Y(_0808_),
    .A(_0807_));
 sg13g2_nor2b_1 _4520_ (.A(_0011_),
    .B_N(_0747_),
    .Y(_0809_));
 sg13g2_xnor2_1 _4521_ (.Y(_0810_),
    .A(_0752_),
    .B(_0809_));
 sg13g2_xnor2_1 _4522_ (.Y(_0811_),
    .A(_0807_),
    .B(_0810_));
 sg13g2_nand2b_1 _4523_ (.Y(_0812_),
    .B(net358),
    .A_N(_0008_));
 sg13g2_nor2_1 _4524_ (.A(_0008_),
    .B(_0707_),
    .Y(_0813_));
 sg13g2_nor2b_1 _4525_ (.A(_0783_),
    .B_N(_0741_),
    .Y(_0814_));
 sg13g2_xnor2_1 _4526_ (.Y(_0815_),
    .A(_0813_),
    .B(_0814_));
 sg13g2_inv_1 _4527_ (.Y(_0816_),
    .A(_0815_));
 sg13g2_xnor2_1 _4528_ (.Y(_0817_),
    .A(_0811_),
    .B(_0815_));
 sg13g2_nor2b_1 _4529_ (.A(_0806_),
    .B_N(_0817_),
    .Y(_0818_));
 sg13g2_xnor2_1 _4530_ (.Y(_0819_),
    .A(_0806_),
    .B(_0817_));
 sg13g2_nor2b_1 _4531_ (.A(_0805_),
    .B_N(_0819_),
    .Y(_0820_));
 sg13g2_xor2_1 _4532_ (.B(_0819_),
    .A(_0805_),
    .X(_0821_));
 sg13g2_nor2_1 _4533_ (.A(_0804_),
    .B(_0821_),
    .Y(_0822_));
 sg13g2_xor2_1 _4534_ (.B(_0821_),
    .A(_0804_),
    .X(_0823_));
 sg13g2_xnor2_1 _4535_ (.Y(_0824_),
    .A(_0803_),
    .B(_0823_));
 sg13g2_nor2_1 _4536_ (.A(_0605_),
    .B(_0824_),
    .Y(_0825_));
 sg13g2_o21ai_1 _4537_ (.B1(_0797_),
    .Y(_0826_),
    .A1(_0773_),
    .A2(_0798_));
 sg13g2_xor2_1 _4538_ (.B(_0824_),
    .A(_0605_),
    .X(_0827_));
 sg13g2_a21oi_1 _4539_ (.A1(_0826_),
    .A2(_0827_),
    .Y(_0828_),
    .B1(_0825_));
 sg13g2_a21oi_1 _4540_ (.A1(_0803_),
    .A2(_0823_),
    .Y(_0829_),
    .B1(_0822_));
 sg13g2_nor2_1 _4541_ (.A(_0818_),
    .B(_0820_),
    .Y(_0830_));
 sg13g2_a22oi_1 _4542_ (.Y(_0831_),
    .B1(_0810_),
    .B2(_0808_),
    .A2(_0809_),
    .A1(net428));
 sg13g2_a22oi_1 _4543_ (.Y(_0832_),
    .B1(_0811_),
    .B2(_0816_),
    .A2(_0784_),
    .A1(_0707_));
 sg13g2_nor3_1 _4544_ (.A(_0008_),
    .B(_0707_),
    .C(_0783_),
    .Y(_0833_));
 sg13g2_and4_1 _4545_ (.A(\main.demo._d___pip_58_1_3___stage___block_3_cx[4] ),
    .B(\main.demo._d___pip_58_1_3___stage___block_3_cx[3] ),
    .C(_0706_),
    .D(_0747_),
    .X(_0834_));
 sg13g2_a22oi_1 _4546_ (.Y(_0835_),
    .B1(_0747_),
    .B2(\main.demo._d___pip_58_1_3___stage___block_3_cx[3] ),
    .A2(_0706_),
    .A1(\main.demo._d___pip_58_1_3___stage___block_3_cx[4] ));
 sg13g2_nor2_1 _4547_ (.A(_0834_),
    .B(_0835_),
    .Y(_0836_));
 sg13g2_xnor2_1 _4548_ (.Y(_0837_),
    .A(_0833_),
    .B(_0836_));
 sg13g2_nor2_1 _4549_ (.A(_0010_),
    .B(_0517_),
    .Y(_0838_));
 sg13g2_inv_1 _4550_ (.Y(_0839_),
    .A(_0838_));
 sg13g2_xnor2_1 _4551_ (.Y(_0840_),
    .A(_0749_),
    .B(_0838_));
 sg13g2_nand2_1 _4552_ (.Y(_0841_),
    .A(_0808_),
    .B(_0840_));
 sg13g2_xnor2_1 _4553_ (.Y(_0842_),
    .A(_0807_),
    .B(_0840_));
 sg13g2_nor2b_1 _4554_ (.A(_0837_),
    .B_N(_0842_),
    .Y(_0843_));
 sg13g2_xnor2_1 _4555_ (.Y(_0844_),
    .A(_0837_),
    .B(_0842_));
 sg13g2_nand2b_1 _4556_ (.Y(_0845_),
    .B(_0844_),
    .A_N(_0832_));
 sg13g2_xnor2_1 _4557_ (.Y(_0846_),
    .A(_0832_),
    .B(_0844_));
 sg13g2_inv_1 _4558_ (.Y(_0847_),
    .A(_0846_));
 sg13g2_xnor2_1 _4559_ (.Y(_0848_),
    .A(_0831_),
    .B(_0846_));
 sg13g2_nand2b_1 _4560_ (.Y(_0849_),
    .B(_0848_),
    .A_N(_0830_));
 sg13g2_xor2_1 _4561_ (.B(_0848_),
    .A(_0830_),
    .X(_0850_));
 sg13g2_xor2_1 _4562_ (.B(_0850_),
    .A(_0829_),
    .X(_0851_));
 sg13g2_nand2_1 _4563_ (.Y(_0852_),
    .A(_0643_),
    .B(_0851_));
 sg13g2_xnor2_1 _4564_ (.Y(_0853_),
    .A(_0643_),
    .B(_0851_));
 sg13g2_xor2_1 _4565_ (.B(_0853_),
    .A(_0828_),
    .X(_0854_));
 sg13g2_nor2b_1 _4566_ (.A(_0013_),
    .B_N(_0854_),
    .Y(_0855_));
 sg13g2_xnor2_1 _4567_ (.Y(_0856_),
    .A(_0826_),
    .B(_0827_));
 sg13g2_or2_1 _4568_ (.X(_0857_),
    .B(_0856_),
    .A(_0014_));
 sg13g2_nor2_1 _4569_ (.A(_0015_),
    .B(_0799_),
    .Y(_0858_));
 sg13g2_a21oi_1 _4570_ (.A1(_0772_),
    .A2(_0800_),
    .Y(_0859_),
    .B1(_0858_));
 sg13g2_xnor2_1 _4571_ (.Y(_0860_),
    .A(_0014_),
    .B(_0856_));
 sg13g2_o21ai_1 _4572_ (.B1(_0857_),
    .Y(_0861_),
    .A1(_0859_),
    .A2(_0860_));
 sg13g2_xnor2_1 _4573_ (.Y(_0862_),
    .A(_0013_),
    .B(_0854_));
 sg13g2_a21oi_2 _4574_ (.B1(_0855_),
    .Y(_0863_),
    .A2(_0862_),
    .A1(_0861_));
 sg13g2_o21ai_1 _4575_ (.B1(_0852_),
    .Y(_0864_),
    .A1(_0828_),
    .A2(_0853_));
 sg13g2_o21ai_1 _4576_ (.B1(_0849_),
    .Y(_0865_),
    .A1(_0829_),
    .A2(_0850_));
 sg13g2_o21ai_1 _4577_ (.B1(_0845_),
    .Y(_0866_),
    .A1(_0831_),
    .A2(_0847_));
 sg13g2_inv_1 _4578_ (.Y(_0867_),
    .A(_0866_));
 sg13g2_o21ai_1 _4579_ (.B1(_0841_),
    .Y(_0868_),
    .A1(_0749_),
    .A2(_0839_));
 sg13g2_a21o_1 _4580_ (.A2(_0836_),
    .A1(_0833_),
    .B1(_0843_),
    .X(_0869_));
 sg13g2_nor2_1 _4581_ (.A(_0011_),
    .B(_0839_),
    .Y(_0870_));
 sg13g2_a21oi_1 _4582_ (.A1(_0010_),
    .A2(_0011_),
    .Y(_0871_),
    .B1(_0517_));
 sg13g2_nor2b_1 _4583_ (.A(_0870_),
    .B_N(_0871_),
    .Y(_0872_));
 sg13g2_xnor2_1 _4584_ (.Y(_0873_),
    .A(_0807_),
    .B(_0872_));
 sg13g2_nor2b_1 _4585_ (.A(_0009_),
    .B_N(_0747_),
    .Y(_0874_));
 sg13g2_nor2b_1 _4586_ (.A(_0008_),
    .B_N(_0874_),
    .Y(_0875_));
 sg13g2_xnor2_1 _4587_ (.Y(_0876_),
    .A(_0812_),
    .B(_0874_));
 sg13g2_nand2_1 _4588_ (.Y(_0877_),
    .A(_0834_),
    .B(_0876_));
 sg13g2_xnor2_1 _4589_ (.Y(_0878_),
    .A(_0834_),
    .B(_0876_));
 sg13g2_inv_1 _4590_ (.Y(_0879_),
    .A(_0878_));
 sg13g2_nand2_1 _4591_ (.Y(_0880_),
    .A(_0873_),
    .B(_0879_));
 sg13g2_xor2_1 _4592_ (.B(_0878_),
    .A(_0873_),
    .X(_0881_));
 sg13g2_nor2b_1 _4593_ (.A(_0881_),
    .B_N(_0869_),
    .Y(_0882_));
 sg13g2_xnor2_1 _4594_ (.Y(_0883_),
    .A(_0869_),
    .B(_0881_));
 sg13g2_xnor2_1 _4595_ (.Y(_0884_),
    .A(_0868_),
    .B(_0883_));
 sg13g2_xor2_1 _4596_ (.B(_0884_),
    .A(_0866_),
    .X(_0885_));
 sg13g2_nand2b_1 _4597_ (.Y(_0886_),
    .B(_0865_),
    .A_N(_0885_));
 sg13g2_xor2_1 _4598_ (.B(_0885_),
    .A(_0865_),
    .X(_0887_));
 sg13g2_nor2b_1 _4599_ (.A(_0887_),
    .B_N(_0700_),
    .Y(_0888_));
 sg13g2_xor2_1 _4600_ (.B(_0887_),
    .A(_0700_),
    .X(_0889_));
 sg13g2_nor2b_1 _4601_ (.A(_0889_),
    .B_N(_0864_),
    .Y(_0890_));
 sg13g2_xor2_1 _4602_ (.B(_0889_),
    .A(_0864_),
    .X(_0891_));
 sg13g2_nor2_1 _4603_ (.A(_0007_),
    .B(_0891_),
    .Y(_0892_));
 sg13g2_xor2_1 _4604_ (.B(_0891_),
    .A(_0007_),
    .X(_0893_));
 sg13g2_nand2b_1 _4605_ (.Y(_0894_),
    .B(_0893_),
    .A_N(_0863_));
 sg13g2_xnor2_1 _4606_ (.Y(_0895_),
    .A(_0863_),
    .B(_0893_));
 sg13g2_xor2_1 _4607_ (.B(_0893_),
    .A(_0863_),
    .X(_0896_));
 sg13g2_nor2_1 _4608_ (.A(net416),
    .B(net421),
    .Y(_0897_));
 sg13g2_or2_1 _4609_ (.X(_0898_),
    .B(net420),
    .A(net416));
 sg13g2_nand2_2 _4610_ (.Y(_0899_),
    .A(\main.demo._q_speed[1] ),
    .B(net389));
 sg13g2_inv_1 _4611_ (.Y(_0900_),
    .A(_0899_));
 sg13g2_nor2_1 _4612_ (.A(_2648_),
    .B(net387),
    .Y(_0901_));
 sg13g2_nand2_2 _4613_ (.Y(_0902_),
    .A(\main.demo._q_speed[2] ),
    .B(net388));
 sg13g2_nor3_1 _4614_ (.A(\main.demo._q_speed[2] ),
    .B(_0896_),
    .C(_0899_),
    .Y(_0903_));
 sg13g2_a21oi_1 _4615_ (.A1(_0895_),
    .A2(_0900_),
    .Y(_0904_),
    .B1(_0902_));
 sg13g2_nor2_1 _4616_ (.A(_0903_),
    .B(_0904_),
    .Y(_0905_));
 sg13g2_o21ai_1 _4617_ (.B1(\main.demo._d___pip_58_1_3___stage___block_3_a[1] ),
    .Y(_0906_),
    .A1(_0903_),
    .A2(_0904_));
 sg13g2_nor3_1 _4618_ (.A(\main.demo._d___pip_58_1_3___stage___block_3_a[1] ),
    .B(_0903_),
    .C(_0904_),
    .Y(_0907_));
 sg13g2_xnor2_1 _4619_ (.Y(_0908_),
    .A(_2656_),
    .B(_0905_));
 sg13g2_inv_2 _4620_ (.Y(_0909_),
    .A(_0908_));
 sg13g2_o21ai_1 _4621_ (.B1(_0906_),
    .Y(_0910_),
    .A1(_0899_),
    .A2(_0907_));
 sg13g2_a21oi_1 _4622_ (.A1(_0899_),
    .A2(_0902_),
    .Y(_0911_),
    .B1(_0896_));
 sg13g2_nand2_1 _4623_ (.Y(_0912_),
    .A(\main.demo._q_speed[3] ),
    .B(net388));
 sg13g2_xor2_1 _4624_ (.B(_0912_),
    .A(_0911_),
    .X(_0913_));
 sg13g2_xnor2_1 _4625_ (.Y(_0914_),
    .A(\main.demo._d___pip_58_1_3___stage___block_3_a[2] ),
    .B(_0913_));
 sg13g2_xor2_1 _4626_ (.B(_0914_),
    .A(_0910_),
    .X(_0915_));
 sg13g2_and2_1 _4627_ (.A(net421),
    .B(_0915_),
    .X(_0916_));
 sg13g2_and2_2 _4628_ (.A(net416),
    .B(net421),
    .X(_0917_));
 sg13g2_nand2_1 _4629_ (.Y(_0918_),
    .A(net417),
    .B(net420));
 sg13g2_nor2_1 _4630_ (.A(_0916_),
    .B(_0917_),
    .Y(_0919_));
 sg13g2_nor2_1 _4631_ (.A(_0802_),
    .B(_0919_),
    .Y(_0920_));
 sg13g2_xnor2_1 _4632_ (.Y(_0921_),
    .A(_0802_),
    .B(_0919_));
 sg13g2_nor2b_1 _4633_ (.A(net416),
    .B_N(net420),
    .Y(_0922_));
 sg13g2_nand2_2 _4634_ (.Y(_0923_),
    .A(net405),
    .B(net420));
 sg13g2_nor2_2 _4635_ (.A(_0908_),
    .B(_0923_),
    .Y(_0924_));
 sg13g2_xnor2_1 _4636_ (.Y(_0925_),
    .A(_0769_),
    .B(_0771_));
 sg13g2_and2_1 _4637_ (.A(_0924_),
    .B(_0925_),
    .X(_0926_));
 sg13g2_xnor2_1 _4638_ (.Y(_0927_),
    .A(_0924_),
    .B(_0925_));
 sg13g2_or2_1 _4639_ (.X(_0928_),
    .B(_0768_),
    .A(\main.demo._q_speed[0] ));
 sg13g2_and3_1 _4640_ (.X(_0929_),
    .A(_0769_),
    .B(net385),
    .C(_0928_));
 sg13g2_nor2b_2 _4641_ (.A(_0927_),
    .B_N(_0929_),
    .Y(_0930_));
 sg13g2_nor2_1 _4642_ (.A(_0926_),
    .B(_0930_),
    .Y(_0931_));
 sg13g2_xnor2_1 _4643_ (.Y(_0932_),
    .A(_0921_),
    .B(_0931_));
 sg13g2_nand2_1 _4644_ (.Y(_0933_),
    .A(net418),
    .B(_0932_));
 sg13g2_nor2_1 _4645_ (.A(_0019_),
    .B(_0913_),
    .Y(_0934_));
 sg13g2_a21oi_2 _4646_ (.B1(_0934_),
    .Y(_0935_),
    .A2(_0914_),
    .A1(_0910_));
 sg13g2_nand2_2 _4647_ (.Y(_0936_),
    .A(\main.demo._q_speed[4] ),
    .B(net389));
 sg13g2_o21ai_1 _4648_ (.B1(net388),
    .Y(_0937_),
    .A1(\main.demo._q_speed[2] ),
    .A2(\main.demo._q_speed[3] ));
 sg13g2_a21oi_1 _4649_ (.A1(_0899_),
    .A2(_0937_),
    .Y(_0938_),
    .B1(_0896_));
 sg13g2_xnor2_1 _4650_ (.Y(_0939_),
    .A(_0936_),
    .B(_0938_));
 sg13g2_nand2b_1 _4651_ (.Y(_0940_),
    .B(_0939_),
    .A_N(_0018_));
 sg13g2_nor2b_1 _4652_ (.A(_0939_),
    .B_N(_0018_),
    .Y(_0941_));
 sg13g2_xnor2_1 _4653_ (.Y(_0942_),
    .A(_0018_),
    .B(_0939_));
 sg13g2_xnor2_1 _4654_ (.Y(_0943_),
    .A(_0935_),
    .B(_0942_));
 sg13g2_nand2_2 _4655_ (.Y(_0944_),
    .A(net385),
    .B(_0943_));
 sg13g2_xnor2_1 _4656_ (.Y(_0945_),
    .A(_0859_),
    .B(_0860_));
 sg13g2_inv_1 _4657_ (.Y(_0946_),
    .A(_0945_));
 sg13g2_nand3_1 _4658_ (.B(_0943_),
    .C(_0946_),
    .A(net386),
    .Y(_0947_));
 sg13g2_xnor2_1 _4659_ (.Y(_0948_),
    .A(_0944_),
    .B(_0945_));
 sg13g2_nand4_1 _4660_ (.B(net420),
    .C(_0909_),
    .A(net416),
    .Y(_0949_),
    .D(_0946_));
 sg13g2_and2_1 _4661_ (.A(_0947_),
    .B(_0949_),
    .X(_0950_));
 sg13g2_nand2_1 _4662_ (.Y(_0951_),
    .A(_0947_),
    .B(_0949_));
 sg13g2_and2_1 _4663_ (.A(_0915_),
    .B(_0917_),
    .X(_0952_));
 sg13g2_o21ai_1 _4664_ (.B1(_0940_),
    .Y(_0953_),
    .A1(_0935_),
    .A2(_0941_));
 sg13g2_nand2_2 _4665_ (.Y(_0954_),
    .A(\main.demo._q_speed[5] ),
    .B(net388));
 sg13g2_nand2_1 _4666_ (.Y(_0955_),
    .A(_0936_),
    .B(_0937_));
 sg13g2_nand4_1 _4667_ (.B(_0902_),
    .C(_0912_),
    .A(_0899_),
    .Y(_0956_),
    .D(_0936_));
 sg13g2_nand2_1 _4668_ (.Y(_0957_),
    .A(_0895_),
    .B(_0956_));
 sg13g2_xor2_1 _4669_ (.B(_0957_),
    .A(_0954_),
    .X(_0958_));
 sg13g2_xor2_1 _4670_ (.B(_0958_),
    .A(\main.demo._d___pip_58_1_3___stage___block_3_a[4] ),
    .X(_0959_));
 sg13g2_xor2_1 _4671_ (.B(_0959_),
    .A(_0953_),
    .X(_0960_));
 sg13g2_xor2_1 _4672_ (.B(_0862_),
    .A(_0861_),
    .X(_0961_));
 sg13g2_nand3_1 _4673_ (.B(_0960_),
    .C(_0961_),
    .A(_0922_),
    .Y(_0962_));
 sg13g2_a21o_1 _4674_ (.A2(_0960_),
    .A1(net386),
    .B1(_0961_),
    .X(_0963_));
 sg13g2_nand3_1 _4675_ (.B(_0916_),
    .C(_0961_),
    .A(net417),
    .Y(_0964_));
 sg13g2_inv_1 _4676_ (.Y(_0965_),
    .A(_0964_));
 sg13g2_a21oi_1 _4677_ (.A1(_0962_),
    .A2(_0963_),
    .Y(_0966_),
    .B1(_0952_));
 sg13g2_a21o_1 _4678_ (.A2(_0963_),
    .A1(_0962_),
    .B1(_0952_),
    .X(_0967_));
 sg13g2_nor3_1 _4679_ (.A(_0950_),
    .B(_0965_),
    .C(_0966_),
    .Y(_0968_));
 sg13g2_nor2_2 _4680_ (.A(net405),
    .B(net420),
    .Y(_0969_));
 sg13g2_nand2b_1 _4681_ (.Y(_0970_),
    .B(net416),
    .A_N(net421));
 sg13g2_a21oi_1 _4682_ (.A1(_0964_),
    .A2(_0967_),
    .Y(_0971_),
    .B1(_0951_));
 sg13g2_nor3_1 _4683_ (.A(_0951_),
    .B(_0965_),
    .C(_0966_),
    .Y(_0972_));
 sg13g2_a21oi_1 _4684_ (.A1(_0964_),
    .A2(_0967_),
    .Y(_0973_),
    .B1(_0950_));
 sg13g2_nor3_1 _4685_ (.A(_0968_),
    .B(_0970_),
    .C(_0971_),
    .Y(_0974_));
 sg13g2_or2_1 _4686_ (.X(_0975_),
    .B(_0974_),
    .A(_0968_));
 sg13g2_nor2_1 _4687_ (.A(_0908_),
    .B(_0970_),
    .Y(_0976_));
 sg13g2_nand2_2 _4688_ (.Y(_0977_),
    .A(_0909_),
    .B(_0969_));
 sg13g2_nand2_1 _4689_ (.Y(_0978_),
    .A(_0962_),
    .B(_0964_));
 sg13g2_inv_1 _4690_ (.Y(_0979_),
    .A(_0978_));
 sg13g2_a22oi_1 _4691_ (.Y(_0980_),
    .B1(_0959_),
    .B2(_0953_),
    .A2(_0958_),
    .A1(_2657_));
 sg13g2_nand2_2 _4692_ (.Y(_0981_),
    .A(\main.demo._q_speed[6] ),
    .B(net388));
 sg13g2_nand3_1 _4693_ (.B(_0937_),
    .C(_0954_),
    .A(_0936_),
    .Y(_0982_));
 sg13g2_nor2b_1 _4694_ (.A(_0956_),
    .B_N(_0954_),
    .Y(_0983_));
 sg13g2_nor2_1 _4695_ (.A(_0896_),
    .B(_0983_),
    .Y(_0984_));
 sg13g2_xnor2_1 _4696_ (.Y(_0985_),
    .A(_0981_),
    .B(_0984_));
 sg13g2_xor2_1 _4697_ (.B(_0985_),
    .A(\main.demo._d___pip_58_1_3___stage___block_3_a[5] ),
    .X(_0986_));
 sg13g2_inv_1 _4698_ (.Y(_0987_),
    .A(_0986_));
 sg13g2_xnor2_1 _4699_ (.Y(_0988_),
    .A(_0980_),
    .B(_0986_));
 sg13g2_nand3_1 _4700_ (.B(net386),
    .C(_0988_),
    .A(_0895_),
    .Y(_0989_));
 sg13g2_a21o_1 _4701_ (.A2(_0988_),
    .A1(net386),
    .B1(_0895_),
    .X(_0990_));
 sg13g2_nand4_1 _4702_ (.B(net420),
    .C(_0895_),
    .A(net416),
    .Y(_0991_),
    .D(_0943_));
 sg13g2_inv_1 _4703_ (.Y(_0992_),
    .A(_0991_));
 sg13g2_a22oi_1 _4704_ (.Y(_0993_),
    .B1(_0989_),
    .B2(_0990_),
    .A2(_0943_),
    .A1(_0917_));
 sg13g2_nor3_1 _4705_ (.A(_0979_),
    .B(_0992_),
    .C(_0993_),
    .Y(_0994_));
 sg13g2_o21ai_1 _4706_ (.B1(_0979_),
    .Y(_0995_),
    .A1(_0992_),
    .A2(_0993_));
 sg13g2_nor2b_1 _4707_ (.A(_0994_),
    .B_N(_0995_),
    .Y(_0996_));
 sg13g2_xnor2_1 _4708_ (.Y(_0997_),
    .A(_0977_),
    .B(_0996_));
 sg13g2_nand2_1 _4709_ (.Y(_0998_),
    .A(_0975_),
    .B(_0997_));
 sg13g2_o21ai_1 _4710_ (.B1(_0948_),
    .Y(_0999_),
    .A1(_0908_),
    .A2(_0918_));
 sg13g2_nand2_2 _4711_ (.Y(_1000_),
    .A(_0949_),
    .B(_0999_));
 sg13g2_or3_1 _4712_ (.A(_0802_),
    .B(_0919_),
    .C(_1000_),
    .X(_1001_));
 sg13g2_nor3_1 _4713_ (.A(_0969_),
    .B(_0972_),
    .C(_0973_),
    .Y(_1002_));
 sg13g2_nor3_1 _4714_ (.A(_0974_),
    .B(_1001_),
    .C(_1002_),
    .Y(_1003_));
 sg13g2_nor2b_1 _4715_ (.A(_0921_),
    .B_N(_0926_),
    .Y(_1004_));
 sg13g2_nor2b_1 _4716_ (.A(_1000_),
    .B_N(_1004_),
    .Y(_1005_));
 sg13g2_nor2b_1 _4717_ (.A(_0921_),
    .B_N(_0930_),
    .Y(_1006_));
 sg13g2_nor2_1 _4718_ (.A(_0920_),
    .B(_1004_),
    .Y(_1007_));
 sg13g2_xor2_1 _4719_ (.B(_1007_),
    .A(_1000_),
    .X(_1008_));
 sg13g2_a21o_1 _4720_ (.A2(_1008_),
    .A1(_1006_),
    .B1(_1005_),
    .X(_1009_));
 sg13g2_o21ai_1 _4721_ (.B1(_1001_),
    .Y(_1010_),
    .A1(_0974_),
    .A2(_1002_));
 sg13g2_nor2b_1 _4722_ (.A(_1003_),
    .B_N(_1010_),
    .Y(_1011_));
 sg13g2_a21oi_1 _4723_ (.A1(_1009_),
    .A2(_1010_),
    .Y(_1012_),
    .B1(_1003_));
 sg13g2_xnor2_1 _4724_ (.Y(_1013_),
    .A(_0975_),
    .B(_0997_));
 sg13g2_o21ai_1 _4725_ (.B1(_0998_),
    .Y(_1014_),
    .A1(_1012_),
    .A2(_1013_));
 sg13g2_a21oi_1 _4726_ (.A1(_0976_),
    .A2(_0995_),
    .Y(_1015_),
    .B1(_0994_));
 sg13g2_xor2_1 _4727_ (.B(net415),
    .A(\main.demo._t___stage___block_3_y[0] ),
    .X(_1016_));
 sg13g2_xnor2_1 _4728_ (.Y(_1017_),
    .A(\main.demo._t___stage___block_3_y[0] ),
    .B(net415));
 sg13g2_mux2_1 _4729_ (.A0(_0799_),
    .A1(_0856_),
    .S(net381),
    .X(_1018_));
 sg13g2_nor2_1 _4730_ (.A(_0013_),
    .B(_1018_),
    .Y(_1019_));
 sg13g2_nand2_1 _4731_ (.Y(_1020_),
    .A(_0766_),
    .B(net383));
 sg13g2_o21ai_1 _4732_ (.B1(_1020_),
    .Y(_1021_),
    .A1(_0799_),
    .A2(net382));
 sg13g2_nand2b_1 _4733_ (.Y(_1022_),
    .B(_1021_),
    .A_N(_0014_));
 sg13g2_xnor2_1 _4734_ (.Y(_1023_),
    .A(_0730_),
    .B(_0731_));
 sg13g2_nor2_1 _4735_ (.A(net381),
    .B(_1023_),
    .Y(_1024_));
 sg13g2_a21oi_1 _4736_ (.A1(_0768_),
    .A2(net381),
    .Y(_1025_),
    .B1(_1024_));
 sg13g2_or2_1 _4737_ (.X(_1026_),
    .B(_1025_),
    .A(_0016_));
 sg13g2_nand2_1 _4738_ (.Y(_1027_),
    .A(_0535_),
    .B(_0729_));
 sg13g2_nand3b_1 _4739_ (.B(net382),
    .C(_1027_),
    .Y(_1028_),
    .A_N(_0730_));
 sg13g2_o21ai_1 _4740_ (.B1(_1028_),
    .Y(_1029_),
    .A1(net382),
    .A2(_1023_));
 sg13g2_nand2_1 _4741_ (.Y(_1030_),
    .A(\main.demo._q_speed[0] ),
    .B(_1029_));
 sg13g2_xnor2_1 _4742_ (.Y(_1031_),
    .A(_0016_),
    .B(_1025_));
 sg13g2_o21ai_1 _4743_ (.B1(_1026_),
    .Y(_1032_),
    .A1(_1030_),
    .A2(_1031_));
 sg13g2_mux2_1 _4744_ (.A0(_0766_),
    .A1(_0768_),
    .S(net382),
    .X(_1033_));
 sg13g2_xnor2_1 _4745_ (.Y(_1034_),
    .A(_2648_),
    .B(_1033_));
 sg13g2_a22oi_1 _4746_ (.Y(_1035_),
    .B1(_1034_),
    .B2(_1032_),
    .A2(_1033_),
    .A1(_2655_));
 sg13g2_xor2_1 _4747_ (.B(_1021_),
    .A(_0014_),
    .X(_1036_));
 sg13g2_o21ai_1 _4748_ (.B1(_1022_),
    .Y(_1037_),
    .A1(_1035_),
    .A2(_1036_));
 sg13g2_xor2_1 _4749_ (.B(_1018_),
    .A(_0013_),
    .X(_1038_));
 sg13g2_a21oi_1 _4750_ (.A1(_1037_),
    .A2(_1038_),
    .Y(_1039_),
    .B1(_1019_));
 sg13g2_nor2_1 _4751_ (.A(_0856_),
    .B(net381),
    .Y(_1040_));
 sg13g2_a21oi_1 _4752_ (.A1(_0854_),
    .A2(net381),
    .Y(_1041_),
    .B1(_1040_));
 sg13g2_or2_1 _4753_ (.X(_1042_),
    .B(_1041_),
    .A(_0007_));
 sg13g2_xnor2_1 _4754_ (.Y(_1043_),
    .A(_0007_),
    .B(_1041_));
 sg13g2_xor2_1 _4755_ (.B(_1043_),
    .A(_1039_),
    .X(_1044_));
 sg13g2_nand3_1 _4756_ (.B(_0901_),
    .C(_1044_),
    .A(_2649_),
    .Y(_1045_));
 sg13g2_a21o_1 _4757_ (.A2(_1044_),
    .A1(_0901_),
    .B1(_0912_),
    .X(_1046_));
 sg13g2_a21o_1 _4758_ (.A2(_1046_),
    .A1(_1045_),
    .B1(_2656_),
    .X(_1047_));
 sg13g2_and3_1 _4759_ (.X(_1048_),
    .A(_2656_),
    .B(_1045_),
    .C(_1046_));
 sg13g2_nand3_1 _4760_ (.B(_1045_),
    .C(_1046_),
    .A(_2656_),
    .Y(_1049_));
 sg13g2_nand2_1 _4761_ (.Y(_1050_),
    .A(_1047_),
    .B(_1049_));
 sg13g2_o21ai_1 _4762_ (.B1(_1047_),
    .Y(_1051_),
    .A1(_0902_),
    .A2(_1048_));
 sg13g2_nor2b_1 _4763_ (.A(_0937_),
    .B_N(net342),
    .Y(_1052_));
 sg13g2_xnor2_1 _4764_ (.Y(_1053_),
    .A(_0936_),
    .B(_1052_));
 sg13g2_xor2_1 _4765_ (.B(_1053_),
    .A(\main.demo._d___pip_58_1_3___stage___block_3_a[2] ),
    .X(_1054_));
 sg13g2_xor2_1 _4766_ (.B(_1054_),
    .A(_1051_),
    .X(_1055_));
 sg13g2_nand2_1 _4767_ (.Y(_1056_),
    .A(_0969_),
    .B(_1055_));
 sg13g2_inv_1 _4768_ (.Y(_1057_),
    .A(_1056_));
 sg13g2_nand2_1 _4769_ (.Y(_1058_),
    .A(_0989_),
    .B(_0991_));
 sg13g2_inv_1 _4770_ (.Y(_1059_),
    .A(_1058_));
 sg13g2_nand2b_1 _4771_ (.Y(_1060_),
    .B(_0985_),
    .A_N(_0022_));
 sg13g2_o21ai_1 _4772_ (.B1(_1060_),
    .Y(_1061_),
    .A1(_0980_),
    .A2(_0987_));
 sg13g2_nand2_2 _4773_ (.Y(_1062_),
    .A(\main.demo._q_speed[7] ),
    .B(net388));
 sg13g2_nand2b_1 _4774_ (.Y(_1063_),
    .B(_0981_),
    .A_N(_0982_));
 sg13g2_nor2_1 _4775_ (.A(_0956_),
    .B(_1063_),
    .Y(_1064_));
 sg13g2_nor2_1 _4776_ (.A(_0896_),
    .B(_1064_),
    .Y(_1065_));
 sg13g2_xnor2_1 _4777_ (.Y(_1066_),
    .A(_1062_),
    .B(_1065_));
 sg13g2_xor2_1 _4778_ (.B(_1066_),
    .A(\main.demo._d___pip_58_1_3___stage___block_3_a[6] ),
    .X(_1067_));
 sg13g2_xor2_1 _4779_ (.B(_1067_),
    .A(_1061_),
    .X(_1068_));
 sg13g2_xnor2_1 _4780_ (.Y(_1069_),
    .A(_1061_),
    .B(_1067_));
 sg13g2_nor2b_1 _4781_ (.A(_0892_),
    .B_N(_0894_),
    .Y(_1070_));
 sg13g2_nor2_1 _4782_ (.A(_0888_),
    .B(_0890_),
    .Y(_1071_));
 sg13g2_nand3_1 _4783_ (.B(_0532_),
    .C(_0698_),
    .A(_0526_),
    .Y(_1072_));
 sg13g2_o21ai_1 _4784_ (.B1(_0886_),
    .Y(_1073_),
    .A1(_0867_),
    .A2(_0884_));
 sg13g2_a21oi_1 _4785_ (.A1(_0868_),
    .A2(_0883_),
    .Y(_1074_),
    .B1(_0882_));
 sg13g2_a21o_1 _4786_ (.A2(_0872_),
    .A1(_0808_),
    .B1(_0870_),
    .X(_1075_));
 sg13g2_nand2_1 _4787_ (.Y(_1076_),
    .A(\main.demo._d___pip_58_1_3___stage___block_3_cx[3] ),
    .B(_0518_));
 sg13g2_a21oi_1 _4788_ (.A1(\main.demo._d___pip_58_1_3___stage___block_3_cx[4] ),
    .A2(net358),
    .Y(_1077_),
    .B1(_1076_));
 sg13g2_nand3_1 _4789_ (.B(net358),
    .C(_1076_),
    .A(\main.demo._d___pip_58_1_3___stage___block_3_cx[4] ),
    .Y(_1078_));
 sg13g2_nand2b_1 _4790_ (.Y(_1079_),
    .B(_1078_),
    .A_N(_1077_));
 sg13g2_nand2_1 _4791_ (.Y(_1080_),
    .A(_0875_),
    .B(_1079_));
 sg13g2_or2_1 _4792_ (.X(_1081_),
    .B(_1079_),
    .A(_0875_));
 sg13g2_nand2_1 _4793_ (.Y(_1082_),
    .A(_1080_),
    .B(_1081_));
 sg13g2_xor2_1 _4794_ (.B(_1082_),
    .A(_0873_),
    .X(_1083_));
 sg13g2_a21oi_1 _4795_ (.A1(_0877_),
    .A2(_0880_),
    .Y(_1084_),
    .B1(_1083_));
 sg13g2_and3_1 _4796_ (.X(_1085_),
    .A(_0877_),
    .B(_0880_),
    .C(_1083_));
 sg13g2_nor2_1 _4797_ (.A(_1084_),
    .B(_1085_),
    .Y(_1086_));
 sg13g2_xnor2_1 _4798_ (.Y(_1087_),
    .A(_1075_),
    .B(_1086_));
 sg13g2_nor2_1 _4799_ (.A(_1074_),
    .B(_1087_),
    .Y(_1088_));
 sg13g2_xor2_1 _4800_ (.B(_1087_),
    .A(_1074_),
    .X(_1089_));
 sg13g2_xor2_1 _4801_ (.B(_1089_),
    .A(_1073_),
    .X(_1090_));
 sg13g2_xor2_1 _4802_ (.B(_1090_),
    .A(_1072_),
    .X(_1091_));
 sg13g2_nor2b_1 _4803_ (.A(_1071_),
    .B_N(_1091_),
    .Y(_1092_));
 sg13g2_xnor2_1 _4804_ (.Y(_1093_),
    .A(_1071_),
    .B(_1091_));
 sg13g2_xnor2_1 _4805_ (.Y(_1094_),
    .A(_0020_),
    .B(_1093_));
 sg13g2_nor2b_1 _4806_ (.A(_1070_),
    .B_N(_1094_),
    .Y(_1095_));
 sg13g2_xnor2_1 _4807_ (.Y(_1096_),
    .A(_1070_),
    .B(_1094_));
 sg13g2_nand3_1 _4808_ (.B(_1068_),
    .C(_1096_),
    .A(net385),
    .Y(_1097_));
 sg13g2_a21o_1 _4809_ (.A2(_1068_),
    .A1(net385),
    .B1(_1096_),
    .X(_1098_));
 sg13g2_nand4_1 _4810_ (.B(net420),
    .C(_0960_),
    .A(net416),
    .Y(_1099_),
    .D(_1096_));
 sg13g2_inv_1 _4811_ (.Y(_1100_),
    .A(_1099_));
 sg13g2_a22oi_1 _4812_ (.Y(_1101_),
    .B1(_1097_),
    .B2(_1098_),
    .A2(_0960_),
    .A1(_0917_));
 sg13g2_nor3_1 _4813_ (.A(_1059_),
    .B(_1100_),
    .C(_1101_),
    .Y(_1102_));
 sg13g2_or3_1 _4814_ (.A(_1059_),
    .B(_1100_),
    .C(_1101_),
    .X(_1103_));
 sg13g2_o21ai_1 _4815_ (.B1(_1059_),
    .Y(_1104_),
    .A1(_1100_),
    .A2(_1101_));
 sg13g2_and3_1 _4816_ (.X(_1105_),
    .A(_1057_),
    .B(_1103_),
    .C(_1104_));
 sg13g2_a21oi_1 _4817_ (.A1(_1103_),
    .A2(_1104_),
    .Y(_1106_),
    .B1(_1057_));
 sg13g2_nor3_1 _4818_ (.A(_1015_),
    .B(_1105_),
    .C(_1106_),
    .Y(_1107_));
 sg13g2_o21ai_1 _4819_ (.B1(_1015_),
    .Y(_1108_),
    .A1(_1105_),
    .A2(_1106_));
 sg13g2_nor2b_1 _4820_ (.A(_1107_),
    .B_N(_1108_),
    .Y(_1109_));
 sg13g2_xnor2_1 _4821_ (.Y(_1110_),
    .A(_1014_),
    .B(_1109_));
 sg13g2_nor2_2 _4822_ (.A(net387),
    .B(_1069_),
    .Y(_1111_));
 sg13g2_xnor2_1 _4823_ (.Y(_1112_),
    .A(_1110_),
    .B(_1111_));
 sg13g2_xnor2_1 _4824_ (.Y(_1113_),
    .A(_1009_),
    .B(_1011_));
 sg13g2_nand2_1 _4825_ (.Y(_1114_),
    .A(net390),
    .B(_0960_));
 sg13g2_xor2_1 _4826_ (.B(_1114_),
    .A(_1113_),
    .X(_1115_));
 sg13g2_nand2_1 _4827_ (.Y(_1116_),
    .A(net390),
    .B(_0915_));
 sg13g2_xnor2_1 _4828_ (.Y(_1117_),
    .A(_0932_),
    .B(_1116_));
 sg13g2_xnor2_1 _4829_ (.Y(_1118_),
    .A(_1006_),
    .B(_1008_));
 sg13g2_nand2_1 _4830_ (.Y(_1119_),
    .A(net390),
    .B(_0943_));
 sg13g2_xnor2_1 _4831_ (.Y(_1120_),
    .A(_1118_),
    .B(_1119_));
 sg13g2_a22oi_1 _4832_ (.Y(_1121_),
    .B1(_1120_),
    .B2(\main.demo._q_th[3] ),
    .A2(_1117_),
    .A1(\main.demo._q_th[2] ));
 sg13g2_nor2_1 _4833_ (.A(\main.demo._q_th[3] ),
    .B(_1120_),
    .Y(_1122_));
 sg13g2_o21ai_1 _4834_ (.B1(_1115_),
    .Y(_1123_),
    .A1(_1121_),
    .A2(_1122_));
 sg13g2_nand2_1 _4835_ (.Y(_1124_),
    .A(net390),
    .B(_0988_));
 sg13g2_xor2_1 _4836_ (.B(_1013_),
    .A(_1012_),
    .X(_1125_));
 sg13g2_xnor2_1 _4837_ (.Y(_1126_),
    .A(_1124_),
    .B(_1125_));
 sg13g2_nand2_1 _4838_ (.Y(_1127_),
    .A(_2611_),
    .B(_1126_));
 sg13g2_nor2_1 _4839_ (.A(_2611_),
    .B(_1126_),
    .Y(_1128_));
 sg13g2_a221oi_1 _4840_ (.B2(_1127_),
    .C1(_1128_),
    .B1(_1123_),
    .A1(_0023_),
    .Y(_1129_),
    .A2(_1112_));
 sg13g2_o21ai_1 _4841_ (.B1(_1129_),
    .Y(_1130_),
    .A1(_0023_),
    .A2(_1112_));
 sg13g2_a22oi_1 _4842_ (.Y(_1131_),
    .B1(_1067_),
    .B2(_1061_),
    .A2(_1066_),
    .A1(_2660_));
 sg13g2_and2_1 _4843_ (.A(\main.demo._q_speed[8] ),
    .B(net388),
    .X(_1132_));
 sg13g2_xor2_1 _4844_ (.B(_1132_),
    .A(\main.demo._d___pip_58_1_3___stage___block_3_a[7] ),
    .X(_1133_));
 sg13g2_nand2b_1 _4845_ (.Y(_1134_),
    .B(_1062_),
    .A_N(_1063_));
 sg13g2_a21oi_1 _4846_ (.A1(_1062_),
    .A2(_1064_),
    .Y(_1135_),
    .B1(_0896_));
 sg13g2_xnor2_1 _4847_ (.Y(_1136_),
    .A(_1133_),
    .B(_1135_));
 sg13g2_o21ai_1 _4848_ (.B1(net389),
    .Y(_1137_),
    .A1(_1131_),
    .A2(_1136_));
 sg13g2_a21o_1 _4849_ (.A2(_1136_),
    .A1(_1131_),
    .B1(_1137_),
    .X(_1138_));
 sg13g2_a21oi_1 _4850_ (.A1(_1014_),
    .A2(_1108_),
    .Y(_1139_),
    .B1(_1107_));
 sg13g2_nor2_1 _4851_ (.A(_1102_),
    .B(_1105_),
    .Y(_1140_));
 sg13g2_nand2_1 _4852_ (.Y(_1141_),
    .A(_0943_),
    .B(_0969_));
 sg13g2_nand2_1 _4853_ (.Y(_1142_),
    .A(_1097_),
    .B(_1099_));
 sg13g2_nand2_1 _4854_ (.Y(_1143_),
    .A(_0982_),
    .B(net342));
 sg13g2_xor2_1 _4855_ (.B(_1143_),
    .A(_0981_),
    .X(_1144_));
 sg13g2_xnor2_1 _4856_ (.Y(_1145_),
    .A(_2657_),
    .B(_1144_));
 sg13g2_nand2_1 _4857_ (.Y(_1146_),
    .A(_0955_),
    .B(net342));
 sg13g2_xor2_1 _4858_ (.B(_1146_),
    .A(_0954_),
    .X(_1147_));
 sg13g2_nor2b_1 _4859_ (.A(_0018_),
    .B_N(_1147_),
    .Y(_1148_));
 sg13g2_nor2b_1 _4860_ (.A(_1147_),
    .B_N(_0018_),
    .Y(_1149_));
 sg13g2_a22oi_1 _4861_ (.Y(_1150_),
    .B1(_1054_),
    .B2(_1051_),
    .A2(_1053_),
    .A1(_2658_));
 sg13g2_a221oi_1 _4862_ (.B2(_1051_),
    .C1(_1148_),
    .B1(_1054_),
    .A1(_2658_),
    .Y(_1151_),
    .A2(_1053_));
 sg13g2_nor3_1 _4863_ (.A(_1145_),
    .B(_1149_),
    .C(_1151_),
    .Y(_1152_));
 sg13g2_a21oi_1 _4864_ (.A1(_2657_),
    .A2(_1144_),
    .Y(_1153_),
    .B1(_1152_));
 sg13g2_nand2_1 _4865_ (.Y(_1154_),
    .A(net342),
    .B(_1063_));
 sg13g2_xor2_1 _4866_ (.B(_1154_),
    .A(_1062_),
    .X(_1155_));
 sg13g2_xor2_1 _4867_ (.B(_1155_),
    .A(\main.demo._d___pip_58_1_3___stage___block_3_a[5] ),
    .X(_1156_));
 sg13g2_inv_1 _4868_ (.Y(_1157_),
    .A(_1156_));
 sg13g2_nand2b_1 _4869_ (.Y(_1158_),
    .B(_1155_),
    .A_N(_0022_));
 sg13g2_o21ai_1 _4870_ (.B1(_1158_),
    .Y(_1159_),
    .A1(_1153_),
    .A2(_1157_));
 sg13g2_nand2_1 _4871_ (.Y(_1160_),
    .A(net342),
    .B(_1134_));
 sg13g2_xnor2_1 _4872_ (.Y(_1161_),
    .A(_1132_),
    .B(_1160_));
 sg13g2_xnor2_1 _4873_ (.Y(_1162_),
    .A(\main.demo._d___pip_58_1_3___stage___block_3_a[6] ),
    .B(_1161_));
 sg13g2_inv_1 _4874_ (.Y(_1163_),
    .A(_1162_));
 sg13g2_a22oi_1 _4875_ (.Y(_1164_),
    .B1(_1163_),
    .B2(_1159_),
    .A2(_1161_),
    .A1(_2660_));
 sg13g2_nand2_1 _4876_ (.Y(_1165_),
    .A(\main.demo._q_speed[9] ),
    .B(net388));
 sg13g2_xnor2_1 _4877_ (.Y(_1166_),
    .A(\main.demo._d___pip_58_1_3___stage___block_3_a[7] ),
    .B(_1165_));
 sg13g2_o21ai_1 _4878_ (.B1(net342),
    .Y(_1167_),
    .A1(_1132_),
    .A2(_1134_));
 sg13g2_xnor2_1 _4879_ (.Y(_1168_),
    .A(_1166_),
    .B(_1167_));
 sg13g2_xnor2_1 _4880_ (.Y(_1169_),
    .A(_1164_),
    .B(_1168_));
 sg13g2_nand2_1 _4881_ (.Y(_1170_),
    .A(net385),
    .B(_1169_));
 sg13g2_nand2_1 _4882_ (.Y(_1171_),
    .A(_0917_),
    .B(_0988_));
 sg13g2_a21oi_1 _4883_ (.A1(_2659_),
    .A2(_1093_),
    .Y(_1172_),
    .B1(_1095_));
 sg13g2_a21oi_1 _4884_ (.A1(_1072_),
    .A2(_1090_),
    .Y(_1173_),
    .B1(_1092_));
 sg13g2_a21oi_1 _4885_ (.A1(_1073_),
    .A2(_1089_),
    .Y(_1174_),
    .B1(_1088_));
 sg13g2_mux2_1 _4886_ (.A0(_1084_),
    .A1(_1085_),
    .S(_1075_),
    .X(_1175_));
 sg13g2_mux2_1 _4887_ (.A0(_1080_),
    .A1(_1081_),
    .S(_0873_),
    .X(_1176_));
 sg13g2_nor3_1 _4888_ (.A(_0009_),
    .B(_0517_),
    .C(_1077_),
    .Y(_1177_));
 sg13g2_a21o_1 _4889_ (.A2(_1077_),
    .A1(_0009_),
    .B1(_1177_),
    .X(_1178_));
 sg13g2_xor2_1 _4890_ (.B(_0531_),
    .A(\main.demo._q_speed[7] ),
    .X(_1179_));
 sg13g2_xnor2_1 _4891_ (.Y(_1180_),
    .A(_1178_),
    .B(_1179_));
 sg13g2_xnor2_1 _4892_ (.Y(_1181_),
    .A(_1176_),
    .B(_1180_));
 sg13g2_xnor2_1 _4893_ (.Y(_1182_),
    .A(_1175_),
    .B(_1181_));
 sg13g2_xnor2_1 _4894_ (.Y(_1183_),
    .A(_1174_),
    .B(_1182_));
 sg13g2_xnor2_1 _4895_ (.Y(_1184_),
    .A(_1173_),
    .B(_1183_));
 sg13g2_xnor2_1 _4896_ (.Y(_1185_),
    .A(_1172_),
    .B(_1184_));
 sg13g2_xnor2_1 _4897_ (.Y(_1186_),
    .A(_1171_),
    .B(_1185_));
 sg13g2_xnor2_1 _4898_ (.Y(_1187_),
    .A(_1170_),
    .B(_1186_));
 sg13g2_xnor2_1 _4899_ (.Y(_1188_),
    .A(_1142_),
    .B(_1187_));
 sg13g2_xnor2_1 _4900_ (.Y(_1189_),
    .A(_1141_),
    .B(_1188_));
 sg13g2_xnor2_1 _4901_ (.Y(_1190_),
    .A(_1140_),
    .B(_1189_));
 sg13g2_xor2_1 _4902_ (.B(_1190_),
    .A(_1139_),
    .X(_1191_));
 sg13g2_xnor2_1 _4903_ (.Y(_1192_),
    .A(_1138_),
    .B(_1191_));
 sg13g2_a22oi_1 _4904_ (.Y(_1193_),
    .B1(_1192_),
    .B2(_2609_),
    .A2(_1112_),
    .A1(_2610_));
 sg13g2_o21ai_1 _4905_ (.B1(net418),
    .Y(_1194_),
    .A1(_2609_),
    .A2(_1191_));
 sg13g2_a21o_2 _4906_ (.A2(_1193_),
    .A1(_1130_),
    .B1(_1194_),
    .X(_1195_));
 sg13g2_xor2_1 _4907_ (.B(_0929_),
    .A(_0927_),
    .X(_1196_));
 sg13g2_o21ai_1 _4908_ (.B1(net390),
    .Y(_1197_),
    .A1(\main.demo._q_speed[1] ),
    .A2(_0909_));
 sg13g2_a21oi_1 _4909_ (.A1(_0900_),
    .A2(_0909_),
    .Y(_1198_),
    .B1(_1197_));
 sg13g2_o21ai_1 _4910_ (.B1(net405),
    .Y(_1199_),
    .A1(_1196_),
    .A2(_1198_));
 sg13g2_a21o_1 _4911_ (.A2(_1198_),
    .A1(_1196_),
    .B1(_1199_),
    .X(_1200_));
 sg13g2_and2_1 _4912_ (.A(_1195_),
    .B(_1200_),
    .X(_1201_));
 sg13g2_nor2_1 _4913_ (.A(net387),
    .B(_1169_),
    .Y(_1202_));
 sg13g2_xor2_1 _4914_ (.B(_1036_),
    .A(_1035_),
    .X(_1203_));
 sg13g2_nor2b_1 _4915_ (.A(_0944_),
    .B_N(_1203_),
    .Y(_1204_));
 sg13g2_nor2_2 _4916_ (.A(_0918_),
    .B(net383),
    .Y(_1205_));
 sg13g2_xnor2_1 _4917_ (.Y(_1206_),
    .A(_0944_),
    .B(_1203_));
 sg13g2_a21o_1 _4918_ (.A2(_1206_),
    .A1(_1205_),
    .B1(_1204_),
    .X(_1207_));
 sg13g2_xnor2_1 _4919_ (.Y(_1208_),
    .A(_0901_),
    .B(_1050_));
 sg13g2_nand2_1 _4920_ (.Y(_1209_),
    .A(_1205_),
    .B(_1208_));
 sg13g2_o21ai_1 _4921_ (.B1(_1145_),
    .Y(_1210_),
    .A1(_1149_),
    .A2(_1151_));
 sg13g2_nor2b_1 _4922_ (.A(_1152_),
    .B_N(_1210_),
    .Y(_1211_));
 sg13g2_nand3b_1 _4923_ (.B(_1210_),
    .C(net386),
    .Y(_1212_),
    .A_N(_1152_));
 sg13g2_xnor2_1 _4924_ (.Y(_1213_),
    .A(_1037_),
    .B(_1038_));
 sg13g2_nor2_1 _4925_ (.A(_1212_),
    .B(_1213_),
    .Y(_1214_));
 sg13g2_xnor2_1 _4926_ (.Y(_1215_),
    .A(_1212_),
    .B(_1213_));
 sg13g2_nor2_1 _4927_ (.A(_1209_),
    .B(_1215_),
    .Y(_1216_));
 sg13g2_xor2_1 _4928_ (.B(_1215_),
    .A(_1209_),
    .X(_1217_));
 sg13g2_nor2_1 _4929_ (.A(net405),
    .B(net381),
    .Y(_1218_));
 sg13g2_nand2_2 _4930_ (.Y(_1219_),
    .A(net418),
    .B(net384));
 sg13g2_xnor2_1 _4931_ (.Y(_1220_),
    .A(_1207_),
    .B(_1217_));
 sg13g2_nor2_2 _4932_ (.A(_1219_),
    .B(_1220_),
    .Y(_1221_));
 sg13g2_a21o_1 _4933_ (.A2(_1217_),
    .A1(_1207_),
    .B1(_1221_),
    .X(_1222_));
 sg13g2_nand2_1 _4934_ (.Y(_1223_),
    .A(_1208_),
    .B(net380));
 sg13g2_or2_1 _4935_ (.X(_1224_),
    .B(_1216_),
    .A(_1214_));
 sg13g2_nand2_1 _4936_ (.Y(_1225_),
    .A(_1055_),
    .B(_1205_));
 sg13g2_inv_1 _4937_ (.Y(_1226_),
    .A(_1225_));
 sg13g2_nand3_1 _4938_ (.B(_0988_),
    .C(net342),
    .A(net385),
    .Y(_1227_));
 sg13g2_a21o_1 _4939_ (.A2(_0988_),
    .A1(net385),
    .B1(net342),
    .X(_1228_));
 sg13g2_nand3_1 _4940_ (.B(_1227_),
    .C(_1228_),
    .A(_1226_),
    .Y(_1229_));
 sg13g2_a21o_1 _4941_ (.A2(_1228_),
    .A1(_1227_),
    .B1(_1226_),
    .X(_1230_));
 sg13g2_and3_1 _4942_ (.X(_1231_),
    .A(_1224_),
    .B(_1229_),
    .C(_1230_));
 sg13g2_a21oi_1 _4943_ (.A1(_1229_),
    .A2(_1230_),
    .Y(_1232_),
    .B1(_1224_));
 sg13g2_or3_1 _4944_ (.A(_1223_),
    .B(_1231_),
    .C(_1232_),
    .X(_1233_));
 sg13g2_o21ai_1 _4945_ (.B1(_1223_),
    .Y(_1234_),
    .A1(_1231_),
    .A2(_1232_));
 sg13g2_nand3_1 _4946_ (.B(_1233_),
    .C(_1234_),
    .A(_1222_),
    .Y(_1235_));
 sg13g2_a21o_1 _4947_ (.A2(_1234_),
    .A1(_1233_),
    .B1(_1222_),
    .X(_1236_));
 sg13g2_nand3_1 _4948_ (.B(_1235_),
    .C(_1236_),
    .A(_0969_),
    .Y(_1237_));
 sg13g2_nand2_1 _4949_ (.Y(_1238_),
    .A(_1235_),
    .B(_1237_));
 sg13g2_nand2b_1 _4950_ (.Y(_1239_),
    .B(_1233_),
    .A_N(_1231_));
 sg13g2_and2_1 _4951_ (.A(_1055_),
    .B(net380),
    .X(_1240_));
 sg13g2_nand2_1 _4952_ (.Y(_1241_),
    .A(_1227_),
    .B(_1229_));
 sg13g2_nor2_1 _4953_ (.A(_1148_),
    .B(_1149_),
    .Y(_1242_));
 sg13g2_xnor2_1 _4954_ (.Y(_1243_),
    .A(_1150_),
    .B(_1242_));
 sg13g2_and2_1 _4955_ (.A(_1205_),
    .B(_1243_),
    .X(_1244_));
 sg13g2_o21ai_1 _4956_ (.B1(_1042_),
    .Y(_1245_),
    .A1(_1039_),
    .A2(_1043_));
 sg13g2_nor2_1 _4957_ (.A(_0891_),
    .B(net382),
    .Y(_1246_));
 sg13g2_a21oi_1 _4958_ (.A1(_0854_),
    .A2(net382),
    .Y(_1247_),
    .B1(_1246_));
 sg13g2_xnor2_1 _4959_ (.Y(_1248_),
    .A(_0020_),
    .B(_1247_));
 sg13g2_nand2b_1 _4960_ (.Y(_1249_),
    .B(_1245_),
    .A_N(_1248_));
 sg13g2_xor2_1 _4961_ (.B(_1248_),
    .A(_1245_),
    .X(_1250_));
 sg13g2_or3_1 _4962_ (.A(_0923_),
    .B(_1069_),
    .C(_1250_),
    .X(_1251_));
 sg13g2_o21ai_1 _4963_ (.B1(_1250_),
    .Y(_1252_),
    .A1(_0923_),
    .A2(_1069_));
 sg13g2_nand3_1 _4964_ (.B(_1251_),
    .C(_1252_),
    .A(_1244_),
    .Y(_1253_));
 sg13g2_a21o_1 _4965_ (.A2(_1252_),
    .A1(_1251_),
    .B1(_1244_),
    .X(_1254_));
 sg13g2_nand3_1 _4966_ (.B(_1253_),
    .C(_1254_),
    .A(_1241_),
    .Y(_1255_));
 sg13g2_a21o_1 _4967_ (.A2(_1254_),
    .A1(_1253_),
    .B1(_1241_),
    .X(_1256_));
 sg13g2_nand3_1 _4968_ (.B(_1255_),
    .C(_1256_),
    .A(_1240_),
    .Y(_1257_));
 sg13g2_a21o_1 _4969_ (.A2(_1256_),
    .A1(_1255_),
    .B1(_1240_),
    .X(_1258_));
 sg13g2_and3_1 _4970_ (.X(_1259_),
    .A(_1239_),
    .B(_1257_),
    .C(_1258_));
 sg13g2_a21oi_1 _4971_ (.A1(_1257_),
    .A2(_1258_),
    .Y(_1260_),
    .B1(_1239_));
 sg13g2_or3_1 _4972_ (.A(_0977_),
    .B(_1259_),
    .C(_1260_),
    .X(_1261_));
 sg13g2_o21ai_1 _4973_ (.B1(_0977_),
    .Y(_1262_),
    .A1(_1259_),
    .A2(_1260_));
 sg13g2_and3_1 _4974_ (.X(_1263_),
    .A(_1238_),
    .B(_1261_),
    .C(_1262_));
 sg13g2_nand3_1 _4975_ (.B(_1261_),
    .C(_1262_),
    .A(_1238_),
    .Y(_1264_));
 sg13g2_xnor2_1 _4976_ (.Y(_1265_),
    .A(_1032_),
    .B(_1034_));
 sg13g2_nand2_1 _4977_ (.Y(_1266_),
    .A(net385),
    .B(_1055_));
 sg13g2_nor2_1 _4978_ (.A(_1265_),
    .B(_1266_),
    .Y(_1267_));
 sg13g2_xnor2_1 _4979_ (.Y(_1268_),
    .A(_1205_),
    .B(_1206_));
 sg13g2_or3_1 _4980_ (.A(_1265_),
    .B(_1266_),
    .C(_1268_),
    .X(_1269_));
 sg13g2_xnor2_1 _4981_ (.Y(_1270_),
    .A(net380),
    .B(_1220_));
 sg13g2_nor2b_1 _4982_ (.A(_1269_),
    .B_N(_1270_),
    .Y(_1271_));
 sg13g2_a21o_1 _4983_ (.A2(_1236_),
    .A1(_1235_),
    .B1(_0969_),
    .X(_1272_));
 sg13g2_and3_1 _4984_ (.X(_1273_),
    .A(_1237_),
    .B(_1271_),
    .C(_1272_));
 sg13g2_xor2_1 _4985_ (.B(_1031_),
    .A(_1030_),
    .X(_1274_));
 sg13g2_and2_1 _4986_ (.A(_0924_),
    .B(_1274_),
    .X(_1275_));
 sg13g2_xor2_1 _4987_ (.B(_1266_),
    .A(_1265_),
    .X(_1276_));
 sg13g2_nand2_1 _4988_ (.Y(_1277_),
    .A(_1275_),
    .B(_1276_));
 sg13g2_xor2_1 _4989_ (.B(_1268_),
    .A(_1267_),
    .X(_1278_));
 sg13g2_nor2_1 _4990_ (.A(_1277_),
    .B(_1278_),
    .Y(_1279_));
 sg13g2_xnor2_1 _4991_ (.Y(_1280_),
    .A(_1269_),
    .B(_1270_));
 sg13g2_and2_1 _4992_ (.A(_1279_),
    .B(_1280_),
    .X(_1281_));
 sg13g2_xnor2_1 _4993_ (.Y(_1282_),
    .A(_0924_),
    .B(_1274_));
 sg13g2_xor2_1 _4994_ (.B(_1029_),
    .A(\main.demo._q_speed[0] ),
    .X(_1283_));
 sg13g2_nand2_1 _4995_ (.Y(_1284_),
    .A(net386),
    .B(_1283_));
 sg13g2_nor2_1 _4996_ (.A(_1282_),
    .B(_1284_),
    .Y(_1285_));
 sg13g2_xor2_1 _4997_ (.B(_1276_),
    .A(_1275_),
    .X(_1286_));
 sg13g2_nand2_2 _4998_ (.Y(_1287_),
    .A(_1285_),
    .B(_1286_));
 sg13g2_xnor2_1 _4999_ (.Y(_1288_),
    .A(_1279_),
    .B(_1280_));
 sg13g2_nor3_2 _5000_ (.A(_1278_),
    .B(_1287_),
    .C(_1288_),
    .Y(_1289_));
 sg13g2_nor2_1 _5001_ (.A(_1281_),
    .B(_1289_),
    .Y(_1290_));
 sg13g2_or2_1 _5002_ (.X(_1291_),
    .B(_1289_),
    .A(_1281_));
 sg13g2_a21oi_1 _5003_ (.A1(_1237_),
    .A2(_1272_),
    .Y(_1292_),
    .B1(_1271_));
 sg13g2_a21o_1 _5004_ (.A2(_1272_),
    .A1(_1237_),
    .B1(_1271_),
    .X(_1293_));
 sg13g2_nor3_1 _5005_ (.A(_1273_),
    .B(_1290_),
    .C(_1292_),
    .Y(_1294_));
 sg13g2_a21oi_2 _5006_ (.B1(_1273_),
    .Y(_1295_),
    .A2(_1293_),
    .A1(_1291_));
 sg13g2_a21oi_1 _5007_ (.A1(_1261_),
    .A2(_1262_),
    .Y(_1296_),
    .B1(_1238_));
 sg13g2_or3_1 _5008_ (.A(_1263_),
    .B(_1295_),
    .C(_1296_),
    .X(_1297_));
 sg13g2_o21ai_1 _5009_ (.B1(_1264_),
    .Y(_1298_),
    .A1(_1295_),
    .A2(_1296_));
 sg13g2_nor2b_1 _5010_ (.A(_1259_),
    .B_N(_1261_),
    .Y(_1299_));
 sg13g2_and2_1 _5011_ (.A(_1255_),
    .B(_1257_),
    .X(_1300_));
 sg13g2_nand2_1 _5012_ (.Y(_1301_),
    .A(net380),
    .B(_1243_));
 sg13g2_and2_1 _5013_ (.A(_1251_),
    .B(_1253_),
    .X(_1302_));
 sg13g2_nand2_1 _5014_ (.Y(_1303_),
    .A(_1205_),
    .B(_1211_));
 sg13g2_o21ai_1 _5015_ (.B1(_1249_),
    .Y(_1304_),
    .A1(_0020_),
    .A2(_1247_));
 sg13g2_nand2_1 _5016_ (.Y(_1305_),
    .A(_0891_),
    .B(net382));
 sg13g2_o21ai_1 _5017_ (.B1(_1305_),
    .Y(_1306_),
    .A1(net382),
    .A2(_1093_));
 sg13g2_xor2_1 _5018_ (.B(_1306_),
    .A(\main.demo._q_speed[7] ),
    .X(_1307_));
 sg13g2_xnor2_1 _5019_ (.Y(_1308_),
    .A(_1304_),
    .B(_1307_));
 sg13g2_xnor2_1 _5020_ (.Y(_1309_),
    .A(_1303_),
    .B(_1308_));
 sg13g2_xnor2_1 _5021_ (.Y(_1310_),
    .A(_1170_),
    .B(_1309_));
 sg13g2_xnor2_1 _5022_ (.Y(_1311_),
    .A(_1302_),
    .B(_1310_));
 sg13g2_xnor2_1 _5023_ (.Y(_1312_),
    .A(_1301_),
    .B(_1311_));
 sg13g2_xnor2_1 _5024_ (.Y(_1313_),
    .A(_1300_),
    .B(_1312_));
 sg13g2_xnor2_1 _5025_ (.Y(_1314_),
    .A(_1057_),
    .B(_1313_));
 sg13g2_xnor2_1 _5026_ (.Y(_1315_),
    .A(_1299_),
    .B(_1314_));
 sg13g2_xnor2_1 _5027_ (.Y(_1316_),
    .A(_1298_),
    .B(_1315_));
 sg13g2_xnor2_1 _5028_ (.Y(_1317_),
    .A(_1202_),
    .B(_1316_));
 sg13g2_o21ai_1 _5029_ (.B1(_1290_),
    .Y(_1318_),
    .A1(_1273_),
    .A2(_1292_));
 sg13g2_nand2b_1 _5030_ (.Y(_1319_),
    .B(_1318_),
    .A_N(_1294_));
 sg13g2_xnor2_1 _5031_ (.Y(_1320_),
    .A(_1153_),
    .B(_1156_));
 sg13g2_nor2_1 _5032_ (.A(net387),
    .B(_1320_),
    .Y(_1321_));
 sg13g2_xnor2_1 _5033_ (.Y(_1322_),
    .A(_1319_),
    .B(_1321_));
 sg13g2_nor2_1 _5034_ (.A(net387),
    .B(_1211_),
    .Y(_1323_));
 sg13g2_o21ai_1 _5035_ (.B1(_1288_),
    .Y(_1324_),
    .A1(_1278_),
    .A2(_1287_));
 sg13g2_nor2b_1 _5036_ (.A(_1289_),
    .B_N(_1324_),
    .Y(_1325_));
 sg13g2_xnor2_1 _5037_ (.Y(_1326_),
    .A(_1323_),
    .B(_1325_));
 sg13g2_xnor2_1 _5038_ (.Y(_1327_),
    .A(_1285_),
    .B(_1286_));
 sg13g2_nor2_1 _5039_ (.A(_0898_),
    .B(_1055_),
    .Y(_1328_));
 sg13g2_xnor2_1 _5040_ (.Y(_1329_),
    .A(_1327_),
    .B(_1328_));
 sg13g2_and2_1 _5041_ (.A(\main.demo._q_th[2] ),
    .B(_1329_),
    .X(_1330_));
 sg13g2_nor2_1 _5042_ (.A(net387),
    .B(_1243_),
    .Y(_1331_));
 sg13g2_nand2_1 _5043_ (.Y(_1332_),
    .A(_1277_),
    .B(_1287_));
 sg13g2_xor2_1 _5044_ (.B(_1332_),
    .A(_1278_),
    .X(_1333_));
 sg13g2_xnor2_1 _5045_ (.Y(_1334_),
    .A(_1331_),
    .B(_1333_));
 sg13g2_a21oi_1 _5046_ (.A1(_1330_),
    .A2(_1334_),
    .Y(_1335_),
    .B1(\main.demo._q_th[3] ));
 sg13g2_nor2_1 _5047_ (.A(_1330_),
    .B(_1334_),
    .Y(_1336_));
 sg13g2_o21ai_1 _5048_ (.B1(_1326_),
    .Y(_1337_),
    .A1(_1335_),
    .A2(_1336_));
 sg13g2_and2_1 _5049_ (.A(\main.demo._q_th[5] ),
    .B(_1337_),
    .X(_1338_));
 sg13g2_nand2b_1 _5050_ (.Y(_1339_),
    .B(_2611_),
    .A_N(_1337_));
 sg13g2_o21ai_1 _5051_ (.B1(_1339_),
    .Y(_1340_),
    .A1(_1322_),
    .A2(_1338_));
 sg13g2_o21ai_1 _5052_ (.B1(_1295_),
    .Y(_1341_),
    .A1(_1263_),
    .A2(_1296_));
 sg13g2_xnor2_1 _5053_ (.Y(_1342_),
    .A(_1159_),
    .B(_1162_));
 sg13g2_nor2_1 _5054_ (.A(net387),
    .B(_1342_),
    .Y(_1343_));
 sg13g2_nand3_1 _5055_ (.B(_1341_),
    .C(_1343_),
    .A(_1297_),
    .Y(_1344_));
 sg13g2_a21o_1 _5056_ (.A2(_1341_),
    .A1(_1297_),
    .B1(_1343_),
    .X(_1345_));
 sg13g2_nand2_1 _5057_ (.Y(_1346_),
    .A(_1344_),
    .B(_1345_));
 sg13g2_nand3_1 _5058_ (.B(_1344_),
    .C(_1345_),
    .A(_2661_),
    .Y(_1347_));
 sg13g2_a21o_1 _5059_ (.A2(_1345_),
    .A1(_1344_),
    .B1(_2661_),
    .X(_1348_));
 sg13g2_nand3_1 _5060_ (.B(_1347_),
    .C(_1348_),
    .A(_1340_),
    .Y(_1349_));
 sg13g2_a22oi_1 _5061_ (.Y(_1350_),
    .B1(_1346_),
    .B2(_2610_),
    .A2(_1317_),
    .A1(_2609_));
 sg13g2_o21ai_1 _5062_ (.B1(net418),
    .Y(_1351_),
    .A1(_2609_),
    .A2(_1317_));
 sg13g2_a21oi_2 _5063_ (.B1(_1351_),
    .Y(_1352_),
    .A2(_1350_),
    .A1(_1349_));
 sg13g2_a21o_2 _5064_ (.A2(_1350_),
    .A1(_1349_),
    .B1(_1351_),
    .X(_1353_));
 sg13g2_nand3_1 _5065_ (.B(net384),
    .C(_1283_),
    .A(net417),
    .Y(_1354_));
 sg13g2_xor2_1 _5066_ (.B(_1284_),
    .A(_1282_),
    .X(_1355_));
 sg13g2_nor2_1 _5067_ (.A(net387),
    .B(_1208_),
    .Y(_1356_));
 sg13g2_xnor2_1 _5068_ (.Y(_1357_),
    .A(_1355_),
    .B(_1356_));
 sg13g2_o21ai_1 _5069_ (.B1(_1354_),
    .Y(_1358_),
    .A1(_1218_),
    .A2(_1357_));
 sg13g2_inv_1 _5070_ (.Y(_1359_),
    .A(_1358_));
 sg13g2_a22oi_1 _5071_ (.Y(_1360_),
    .B1(_1353_),
    .B2(_1359_),
    .A2(_1201_),
    .A1(_0933_));
 sg13g2_and4_1 _5072_ (.A(_0933_),
    .B(_1201_),
    .C(_1353_),
    .D(_1359_),
    .X(_1361_));
 sg13g2_or3_1 _5073_ (.A(net406),
    .B(_1360_),
    .C(_1361_),
    .X(_1362_));
 sg13g2_or2_1 _5074_ (.X(_1363_),
    .B(_1322_),
    .A(_1126_));
 sg13g2_nor2_2 _5075_ (.A(net419),
    .B(_1363_),
    .Y(_1364_));
 sg13g2_nand2_1 _5076_ (.Y(_1365_),
    .A(_1218_),
    .B(_1357_));
 sg13g2_o21ai_1 _5077_ (.B1(_1365_),
    .Y(_1366_),
    .A1(net380),
    .A2(_1329_));
 sg13g2_inv_1 _5078_ (.Y(_1367_),
    .A(_1366_));
 sg13g2_nand2_1 _5079_ (.Y(_1368_),
    .A(_1364_),
    .B(_1366_));
 sg13g2_and2_2 _5080_ (.A(net406),
    .B(_1126_),
    .X(_1369_));
 sg13g2_nand2_1 _5081_ (.Y(_1370_),
    .A(_1201_),
    .B(_1369_));
 sg13g2_nand3_1 _5082_ (.B(_1368_),
    .C(_1370_),
    .A(_1362_),
    .Y(\main.demo._t___block_68_frag[0] ));
 sg13g2_nand2_1 _5083_ (.Y(_1371_),
    .A(net405),
    .B(_1117_));
 sg13g2_nand2_1 _5084_ (.Y(_1372_),
    .A(net418),
    .B(_1118_));
 sg13g2_nand3_1 _5085_ (.B(_1371_),
    .C(_1372_),
    .A(_1195_),
    .Y(_1373_));
 sg13g2_inv_1 _5086_ (.Y(_1374_),
    .A(_1373_));
 sg13g2_nor3_1 _5087_ (.A(_1352_),
    .B(_1367_),
    .C(_1373_),
    .Y(_1375_));
 sg13g2_o21ai_1 _5088_ (.B1(_1373_),
    .Y(_1376_),
    .A1(_1352_),
    .A2(_1367_));
 sg13g2_nand2b_1 _5089_ (.Y(_1377_),
    .B(_1376_),
    .A_N(_1375_));
 sg13g2_xnor2_1 _5090_ (.Y(_1378_),
    .A(_1361_),
    .B(_1377_));
 sg13g2_mux2_1 _5091_ (.A0(_1329_),
    .A1(_1334_),
    .S(_1219_),
    .X(_1379_));
 sg13g2_nor3_1 _5092_ (.A(net419),
    .B(_1334_),
    .C(_1363_),
    .Y(_1380_));
 sg13g2_a221oi_1 _5093_ (.B2(net419),
    .C1(_1380_),
    .B1(_1378_),
    .A1(_1369_),
    .Y(_1381_),
    .A2(_1374_));
 sg13g2_inv_1 _5094_ (.Y(\main.demo._t___block_68_frag[1] ),
    .A(_1381_));
 sg13g2_nand2_1 _5095_ (.Y(_1382_),
    .A(net405),
    .B(_1120_));
 sg13g2_nand2_1 _5096_ (.Y(_1383_),
    .A(net418),
    .B(_1113_));
 sg13g2_nand3_1 _5097_ (.B(_1382_),
    .C(_1383_),
    .A(_1195_),
    .Y(_1384_));
 sg13g2_inv_1 _5098_ (.Y(_1385_),
    .A(_1384_));
 sg13g2_nor3_1 _5099_ (.A(_1352_),
    .B(_1379_),
    .C(_1384_),
    .Y(_1386_));
 sg13g2_o21ai_1 _5100_ (.B1(_1384_),
    .Y(_1387_),
    .A1(_1352_),
    .A2(_1379_));
 sg13g2_nand2b_1 _5101_ (.Y(_1388_),
    .B(_1387_),
    .A_N(_1386_));
 sg13g2_a21oi_1 _5102_ (.A1(_1361_),
    .A2(_1376_),
    .Y(_1389_),
    .B1(_1375_));
 sg13g2_nor2_1 _5103_ (.A(_1388_),
    .B(_1389_),
    .Y(_1390_));
 sg13g2_a21o_1 _5104_ (.A2(_1389_),
    .A1(_1388_),
    .B1(net406),
    .X(_1391_));
 sg13g2_nand2_1 _5105_ (.Y(_1392_),
    .A(_1219_),
    .B(_1326_));
 sg13g2_o21ai_1 _5106_ (.B1(_1392_),
    .Y(_1393_),
    .A1(_1219_),
    .A2(_1334_));
 sg13g2_a22oi_1 _5107_ (.Y(_1394_),
    .B1(_1393_),
    .B2(_1364_),
    .A2(_1385_),
    .A1(_1369_));
 sg13g2_o21ai_1 _5108_ (.B1(_1394_),
    .Y(\main.demo._t___block_68_frag[2] ),
    .A1(_1390_),
    .A2(_1391_));
 sg13g2_mux2_1 _5109_ (.A0(_1115_),
    .A1(_1125_),
    .S(net418),
    .X(_1395_));
 sg13g2_and2_1 _5110_ (.A(_1195_),
    .B(_1395_),
    .X(_1396_));
 sg13g2_a21o_1 _5111_ (.A2(_1393_),
    .A1(_1353_),
    .B1(_1396_),
    .X(_1397_));
 sg13g2_nand3_1 _5112_ (.B(_1393_),
    .C(_1396_),
    .A(_1353_),
    .Y(_1398_));
 sg13g2_nand2_1 _5113_ (.Y(_1399_),
    .A(_1397_),
    .B(_1398_));
 sg13g2_nor2_1 _5114_ (.A(_1386_),
    .B(_1390_),
    .Y(_1400_));
 sg13g2_xnor2_1 _5115_ (.Y(_1401_),
    .A(_1399_),
    .B(_1400_));
 sg13g2_nor2_1 _5116_ (.A(net380),
    .B(_1322_),
    .Y(_1402_));
 sg13g2_o21ai_1 _5117_ (.B1(_1353_),
    .Y(_1403_),
    .A1(_1221_),
    .A2(_1402_));
 sg13g2_nor2_1 _5118_ (.A(_1363_),
    .B(_1403_),
    .Y(_1404_));
 sg13g2_nand2_1 _5119_ (.Y(_1405_),
    .A(_1126_),
    .B(_1396_));
 sg13g2_nor2_1 _5120_ (.A(net418),
    .B(_1404_),
    .Y(_1406_));
 sg13g2_a22oi_1 _5121_ (.Y(\main.demo._t___block_68_frag[3] ),
    .B1(_1405_),
    .B2(_1406_),
    .A2(_1401_),
    .A1(net419));
 sg13g2_nor2b_1 _5122_ (.A(_1386_),
    .B_N(_1398_),
    .Y(_1407_));
 sg13g2_o21ai_1 _5123_ (.B1(_1407_),
    .Y(_1408_),
    .A1(_1388_),
    .A2(_1389_));
 sg13g2_nand2_1 _5124_ (.Y(_1409_),
    .A(_1397_),
    .B(_1408_));
 sg13g2_nor2_1 _5125_ (.A(net405),
    .B(_1110_),
    .Y(_1410_));
 sg13g2_o21ai_1 _5126_ (.B1(_1195_),
    .Y(_1411_),
    .A1(_1369_),
    .A2(_1410_));
 sg13g2_or2_1 _5127_ (.X(_1412_),
    .B(_1411_),
    .A(_1403_));
 sg13g2_xnor2_1 _5128_ (.Y(_1413_),
    .A(_1403_),
    .B(_1411_));
 sg13g2_nand3b_1 _5129_ (.B(_1408_),
    .C(_1397_),
    .Y(_1414_),
    .A_N(_1413_));
 sg13g2_a21oi_1 _5130_ (.A1(_1409_),
    .A2(_1413_),
    .Y(_1415_),
    .B1(net406));
 sg13g2_nor2_1 _5131_ (.A(net380),
    .B(_1346_),
    .Y(_1416_));
 sg13g2_a21oi_2 _5132_ (.B1(_1416_),
    .Y(_1417_),
    .A2(_1322_),
    .A1(net380));
 sg13g2_a221oi_1 _5133_ (.B2(_1364_),
    .C1(_1369_),
    .B1(_1417_),
    .A1(_1414_),
    .Y(_1418_),
    .A2(_1415_));
 sg13g2_inv_1 _5134_ (.Y(\main.demo._t___block_68_frag[4] ),
    .A(_1418_));
 sg13g2_nand2_1 _5135_ (.Y(_1419_),
    .A(_1112_),
    .B(_1369_));
 sg13g2_and2_1 _5136_ (.A(_1412_),
    .B(_1414_),
    .X(_1420_));
 sg13g2_nand2_1 _5137_ (.Y(_1421_),
    .A(_1353_),
    .B(_1417_));
 sg13g2_nand2b_1 _5138_ (.Y(_1422_),
    .B(net419),
    .A_N(_1191_));
 sg13g2_o21ai_1 _5139_ (.B1(_1422_),
    .Y(_1423_),
    .A1(net419),
    .A2(_1112_));
 sg13g2_nand2b_1 _5140_ (.Y(_1424_),
    .B(_1195_),
    .A_N(_1423_));
 sg13g2_xnor2_1 _5141_ (.Y(_1425_),
    .A(_1421_),
    .B(_1424_));
 sg13g2_nor2_1 _5142_ (.A(_1420_),
    .B(_1425_),
    .Y(_1426_));
 sg13g2_a21o_1 _5143_ (.A2(_1425_),
    .A1(_1420_),
    .B1(net406),
    .X(_1427_));
 sg13g2_o21ai_1 _5144_ (.B1(_1419_),
    .Y(\main.demo._t___block_68_frag[5] ),
    .A1(_1426_),
    .A2(_1427_));
 sg13g2_nor3_2 _5145_ (.A(\main.demo.zic._q_squ_env[5] ),
    .B(\main.demo.zic._q_squ_env[4] ),
    .C(\main.demo.zic._q_squ_env[3] ),
    .Y(_1428_));
 sg13g2_nor2_2 _5146_ (.A(\main.demo.zic._q_qpos[12] ),
    .B(_1428_),
    .Y(_1429_));
 sg13g2_or2_2 _5147_ (.X(_1430_),
    .B(_1428_),
    .A(\main.demo.zic._q_qpos[12] ));
 sg13g2_nor2b_2 _5148_ (.A(\main._w_demo_video_vs ),
    .B_N(\main.demo._q_prev_vs ),
    .Y(_1431_));
 sg13g2_nand2b_2 _5149_ (.Y(_1432_),
    .B(\main.demo._q_prev_vs ),
    .A_N(\main._w_demo_video_vs ));
 sg13g2_nand2_1 _5150_ (.Y(_1433_),
    .A(\main.demo._q_frame[1] ),
    .B(\main.demo._q_frame[0] ));
 sg13g2_nand2_1 _5151_ (.Y(_1434_),
    .A(\main.demo._q_frame[0] ),
    .B(_1431_));
 sg13g2_nor3_2 _5152_ (.A(_2634_),
    .B(_1432_),
    .C(_1433_),
    .Y(_1435_));
 sg13g2_and2_1 _5153_ (.A(\main.demo._q_frame[3] ),
    .B(_1435_),
    .X(_1436_));
 sg13g2_and2_1 _5154_ (.A(net435),
    .B(_1436_),
    .X(_1437_));
 sg13g2_and2_1 _5155_ (.A(_2938_),
    .B(_1437_),
    .X(_1438_));
 sg13g2_and2_1 _5156_ (.A(net500),
    .B(_1438_),
    .X(_1439_));
 sg13g2_and2_2 _5157_ (.A(net634),
    .B(_1439_),
    .X(_1440_));
 sg13g2_and2_1 _5158_ (.A(\main.demo._q_frame[9] ),
    .B(_1440_),
    .X(_1441_));
 sg13g2_xor2_1 _5159_ (.B(_1440_),
    .A(net630),
    .X(_1442_));
 sg13g2_nor2_2 _5160_ (.A(net636),
    .B(_1442_),
    .Y(_1443_));
 sg13g2_xnor2_1 _5161_ (.Y(_1444_),
    .A(\main.demo.zic._q_tpos[11] ),
    .B(_1430_));
 sg13g2_nand2_1 _5162_ (.Y(_1445_),
    .A(net530),
    .B(net529));
 sg13g2_xor2_1 _5163_ (.B(\main.demo.zic._q_tpos[10] ),
    .A(\main.demo.zic._q_tpos[11] ),
    .X(_1446_));
 sg13g2_xnor2_1 _5164_ (.Y(_1447_),
    .A(\main.demo.zic._q_tpos[9] ),
    .B(_1446_));
 sg13g2_xnor2_1 _5165_ (.Y(_1448_),
    .A(\main.demo.zic._q_tpos[8] ),
    .B(_1446_));
 sg13g2_xnor2_1 _5166_ (.Y(_1449_),
    .A(\main.demo.zic._q_tpos[7] ),
    .B(_1446_));
 sg13g2_o21ai_1 _5167_ (.B1(\main.demo.zic._q_squ_env[5] ),
    .Y(_1450_),
    .A1(\main.demo.zic._q_squ_env[4] ),
    .A2(\main.demo.zic._q_squ_env[3] ));
 sg13g2_nand2_1 _5168_ (.Y(_1451_),
    .A(_1429_),
    .B(_1450_));
 sg13g2_o21ai_1 _5169_ (.B1(_1451_),
    .Y(_1452_),
    .A1(_2616_),
    .A2(_0025_));
 sg13g2_xnor2_1 _5170_ (.Y(_1453_),
    .A(\main.demo.zic._q_tpos[6] ),
    .B(_1446_));
 sg13g2_inv_1 _5171_ (.Y(_1454_),
    .A(_1453_));
 sg13g2_nand2_1 _5172_ (.Y(_1455_),
    .A(_1452_),
    .B(_1454_));
 sg13g2_xnor2_1 _5173_ (.Y(_1456_),
    .A(_1452_),
    .B(_1453_));
 sg13g2_xnor2_1 _5174_ (.Y(_1457_),
    .A(\main.demo.zic._q_tpos[5] ),
    .B(_1446_));
 sg13g2_xor2_1 _5175_ (.B(\main.demo.zic._q_squ_env[3] ),
    .A(\main.demo.zic._q_squ_env[4] ),
    .X(_1458_));
 sg13g2_nand2_1 _5176_ (.Y(_1459_),
    .A(\main.demo.zic._q_qpos[12] ),
    .B(_0024_));
 sg13g2_o21ai_1 _5177_ (.B1(_1459_),
    .Y(_1460_),
    .A1(\main.demo.zic._q_qpos[12] ),
    .A2(_1458_));
 sg13g2_nor2_1 _5178_ (.A(_1457_),
    .B(_1460_),
    .Y(_1461_));
 sg13g2_xor2_1 _5179_ (.B(_1446_),
    .A(\main.demo.zic._q_tpos[4] ),
    .X(_1462_));
 sg13g2_xor2_1 _5180_ (.B(_1460_),
    .A(_1457_),
    .X(_1463_));
 sg13g2_and3_1 _5181_ (.X(_1464_),
    .A(\main.demo.zic._q_squ_env[3] ),
    .B(_1462_),
    .C(_1463_));
 sg13g2_nor2_1 _5182_ (.A(_1461_),
    .B(_1464_),
    .Y(_1465_));
 sg13g2_nand2b_1 _5183_ (.Y(_1466_),
    .B(_1456_),
    .A_N(_1465_));
 sg13g2_xnor2_1 _5184_ (.Y(_1467_),
    .A(_1430_),
    .B(_1449_));
 sg13g2_a21o_1 _5185_ (.A2(_1466_),
    .A1(_1455_),
    .B1(_1467_),
    .X(_1468_));
 sg13g2_o21ai_1 _5186_ (.B1(_1468_),
    .Y(_1469_),
    .A1(_1430_),
    .A2(_1449_));
 sg13g2_xnor2_1 _5187_ (.Y(_1470_),
    .A(_1430_),
    .B(_1448_));
 sg13g2_nand2b_1 _5188_ (.Y(_1471_),
    .B(_1469_),
    .A_N(_1470_));
 sg13g2_o21ai_1 _5189_ (.B1(_1471_),
    .Y(_1472_),
    .A1(_1430_),
    .A2(_1448_));
 sg13g2_xnor2_1 _5190_ (.Y(_1473_),
    .A(_1430_),
    .B(_1447_));
 sg13g2_nand2b_1 _5191_ (.Y(_1474_),
    .B(_1472_),
    .A_N(_1473_));
 sg13g2_o21ai_1 _5192_ (.B1(_1474_),
    .Y(_1475_),
    .A1(_1430_),
    .A2(_1447_));
 sg13g2_a21oi_1 _5193_ (.A1(_1444_),
    .A2(_1475_),
    .Y(_1476_),
    .B1(_1443_));
 sg13g2_o21ai_1 _5194_ (.B1(_1476_),
    .Y(_1477_),
    .A1(\main.demo.zic._q_tpos[11] ),
    .A2(_1429_));
 sg13g2_nor2_1 _5195_ (.A(_0026_),
    .B(_1477_),
    .Y(_1478_));
 sg13g2_o21ai_1 _5196_ (.B1(_1476_),
    .Y(_1479_),
    .A1(_1444_),
    .A2(_1475_));
 sg13g2_inv_1 _5197_ (.Y(_1480_),
    .A(_1479_));
 sg13g2_xor2_1 _5198_ (.B(_1473_),
    .A(_1472_),
    .X(_1481_));
 sg13g2_or2_1 _5199_ (.X(_1482_),
    .B(_1481_),
    .A(\main.demo.zic._q_clock_count[4] ));
 sg13g2_xor2_1 _5200_ (.B(_1470_),
    .A(_1469_),
    .X(_1483_));
 sg13g2_nor2_1 _5201_ (.A(_2666_),
    .B(_1483_),
    .Y(_1484_));
 sg13g2_a21oi_1 _5202_ (.A1(\main.demo.zic._q_squ_env[3] ),
    .A2(_1462_),
    .Y(_1485_),
    .B1(_1463_));
 sg13g2_nor3_1 _5203_ (.A(\main.demo.zic._q_clock_count[0] ),
    .B(_1464_),
    .C(_1485_),
    .Y(_1486_));
 sg13g2_nand2b_1 _5204_ (.Y(_1487_),
    .B(\main.demo.zic._q_clock_count[1] ),
    .A_N(_1486_));
 sg13g2_nor2b_1 _5205_ (.A(\main.demo.zic._q_clock_count[1] ),
    .B_N(_1486_),
    .Y(_1488_));
 sg13g2_xnor2_1 _5206_ (.Y(_1489_),
    .A(_1456_),
    .B(_1465_));
 sg13g2_o21ai_1 _5207_ (.B1(_1487_),
    .Y(_1490_),
    .A1(_1488_),
    .A2(_1489_));
 sg13g2_nand3_1 _5208_ (.B(_1466_),
    .C(_1467_),
    .A(_1455_),
    .Y(_1491_));
 sg13g2_nand3_1 _5209_ (.B(_1468_),
    .C(_1491_),
    .A(_2638_),
    .Y(_1492_));
 sg13g2_a21oi_1 _5210_ (.A1(_1468_),
    .A2(_1491_),
    .Y(_1493_),
    .B1(_2638_));
 sg13g2_a221oi_1 _5211_ (.B2(_1492_),
    .C1(_1493_),
    .B1(_1490_),
    .A1(_2666_),
    .Y(_1494_),
    .A2(_1483_));
 sg13g2_nand2_1 _5212_ (.Y(_1495_),
    .A(\main.demo.zic._q_clock_count[4] ),
    .B(_1481_));
 sg13g2_o21ai_1 _5213_ (.B1(_1495_),
    .Y(_1496_),
    .A1(_1484_),
    .A2(_1494_));
 sg13g2_a21oi_1 _5214_ (.A1(_1482_),
    .A2(_1496_),
    .Y(_1497_),
    .B1(_1443_));
 sg13g2_o21ai_1 _5215_ (.B1(_1497_),
    .Y(_1498_),
    .A1(net303),
    .A2(_1480_));
 sg13g2_a22oi_1 _5216_ (.Y(_1499_),
    .B1(_1480_),
    .B2(net303),
    .A2(_1477_),
    .A1(_0026_));
 sg13g2_a21oi_1 _5217_ (.A1(_1498_),
    .A2(net304),
    .Y(\main._w_demo_audio1 ),
    .B1(_1478_));
 sg13g2_o21ai_1 _5218_ (.B1(net399),
    .Y(\main.demo._t___pip_58_1_3___block_87_atten_h[2] ),
    .A1(net556),
    .A2(net426));
 sg13g2_a21oi_1 _5219_ (.A1(net551),
    .A2(\main.demo._t___pip_58_1_3___block_87_atten_h[0] ),
    .Y(\main.demo._t___pip_58_1_3___block_87_atten_h[1] ),
    .B1(\main.demo._t___pip_58_1_3___block_87_atten_h[2] ));
 sg13g2_xnor2_1 _5220_ (.Y(_1500_),
    .A(_2676_),
    .B(_2737_));
 sg13g2_nor2_1 _5221_ (.A(_2704_),
    .B(net351),
    .Y(_1501_));
 sg13g2_xnor2_1 _5222_ (.Y(_1502_),
    .A(_2714_),
    .B(_1501_));
 sg13g2_nor2_1 _5223_ (.A(_1500_),
    .B(_1502_),
    .Y(_1503_));
 sg13g2_xor2_1 _5224_ (.B(_1502_),
    .A(_1500_),
    .X(_1504_));
 sg13g2_xnor2_1 _5225_ (.Y(_1505_),
    .A(_2705_),
    .B(_1504_));
 sg13g2_nor3_1 _5226_ (.A(\main.demo._q___pip_58_1_2___stage___block_3_cx[9] ),
    .B(_2761_),
    .C(_2766_),
    .Y(_1506_));
 sg13g2_a21oi_1 _5227_ (.A1(_2761_),
    .A2(_2766_),
    .Y(_1507_),
    .B1(_1506_));
 sg13g2_xnor2_1 _5228_ (.Y(_1508_),
    .A(_0052_),
    .B(_1507_));
 sg13g2_or2_1 _5229_ (.X(_1509_),
    .B(_2778_),
    .A(_2767_));
 sg13g2_o21ai_1 _5230_ (.B1(_1508_),
    .Y(_1510_),
    .A1(net351),
    .A2(_1509_));
 sg13g2_a21oi_1 _5231_ (.A1(_1508_),
    .A2(_1509_),
    .Y(_1511_),
    .B1(net351));
 sg13g2_a21oi_2 _5232_ (.B1(_1511_),
    .Y(_1512_),
    .A2(_1508_),
    .A1(net351));
 sg13g2_inv_1 _5233_ (.Y(_1513_),
    .A(_1512_));
 sg13g2_o21ai_1 _5234_ (.B1(_2797_),
    .Y(_1514_),
    .A1(_0047_),
    .A2(_2784_));
 sg13g2_xnor2_1 _5235_ (.Y(_1515_),
    .A(_2798_),
    .B(_1514_));
 sg13g2_nand2_1 _5236_ (.Y(_1516_),
    .A(_1512_),
    .B(_1515_));
 sg13g2_nor2_1 _5237_ (.A(_1512_),
    .B(_1515_),
    .Y(_1517_));
 sg13g2_xnor2_1 _5238_ (.Y(_1518_),
    .A(_2795_),
    .B(_2796_));
 sg13g2_nor2_1 _5239_ (.A(_1513_),
    .B(_1518_),
    .Y(_1519_));
 sg13g2_xnor2_1 _5240_ (.Y(_1520_),
    .A(_1512_),
    .B(_1518_));
 sg13g2_xnor2_1 _5241_ (.Y(_1521_),
    .A(_2792_),
    .B(_2794_));
 sg13g2_and2_1 _5242_ (.A(_1512_),
    .B(_1521_),
    .X(_1522_));
 sg13g2_xor2_1 _5243_ (.B(_1521_),
    .A(_1512_),
    .X(_1523_));
 sg13g2_o21ai_1 _5244_ (.B1(_1513_),
    .Y(_1524_),
    .A1(_1508_),
    .A2(_1509_));
 sg13g2_xnor2_1 _5245_ (.Y(_1525_),
    .A(_2789_),
    .B(_2791_));
 sg13g2_nand2_1 _5246_ (.Y(_1526_),
    .A(_1524_),
    .B(_1525_));
 sg13g2_a21oi_1 _5247_ (.A1(_2807_),
    .A2(_2830_),
    .Y(_1527_),
    .B1(_2806_));
 sg13g2_xnor2_1 _5248_ (.Y(_1528_),
    .A(_1524_),
    .B(_1525_));
 sg13g2_o21ai_1 _5249_ (.B1(_1526_),
    .Y(_1529_),
    .A1(_1527_),
    .A2(_1528_));
 sg13g2_a21o_1 _5250_ (.A2(_1529_),
    .A1(_1523_),
    .B1(_1522_),
    .X(_1530_));
 sg13g2_a21oi_1 _5251_ (.A1(_1520_),
    .A2(_1530_),
    .Y(_1531_),
    .B1(_1519_));
 sg13g2_a21oi_1 _5252_ (.A1(_1516_),
    .A2(_1531_),
    .Y(_1532_),
    .B1(_1517_));
 sg13g2_xor2_1 _5253_ (.B(_1532_),
    .A(_1510_),
    .X(_1533_));
 sg13g2_nand2_1 _5254_ (.Y(_1534_),
    .A(_2831_),
    .B(_1533_));
 sg13g2_xor2_1 _5255_ (.B(_1528_),
    .A(_1527_),
    .X(_1535_));
 sg13g2_xnor2_1 _5256_ (.Y(_1536_),
    .A(_1534_),
    .B(_1535_));
 sg13g2_inv_1 _5257_ (.Y(_1537_),
    .A(_1536_));
 sg13g2_xor2_1 _5258_ (.B(_1536_),
    .A(_1505_),
    .X(_1538_));
 sg13g2_nor2_1 _5259_ (.A(_2832_),
    .B(_1538_),
    .Y(_1539_));
 sg13g2_xor2_1 _5260_ (.B(_1538_),
    .A(_2832_),
    .X(\main.demo._d___pip_58_1_2___stage___block_3_cx[1] ));
 sg13g2_a21oi_1 _5261_ (.A1(_1505_),
    .A2(_1537_),
    .Y(_1540_),
    .B1(_1539_));
 sg13g2_a21oi_1 _5262_ (.A1(_2706_),
    .A2(_1504_),
    .Y(_1541_),
    .B1(_1503_));
 sg13g2_xor2_1 _5263_ (.B(_2739_),
    .A(_2738_),
    .X(_1542_));
 sg13g2_inv_1 _5264_ (.Y(_1543_),
    .A(_1542_));
 sg13g2_nand2_1 _5265_ (.Y(_1544_),
    .A(_2704_),
    .B(_2714_));
 sg13g2_nand2_1 _5266_ (.Y(_1545_),
    .A(net349),
    .B(_1544_));
 sg13g2_xor2_1 _5267_ (.B(_1545_),
    .A(_1525_),
    .X(_1546_));
 sg13g2_xnor2_1 _5268_ (.Y(_1547_),
    .A(_1542_),
    .B(_1546_));
 sg13g2_nor2b_1 _5269_ (.A(_1541_),
    .B_N(_1547_),
    .Y(_1548_));
 sg13g2_xnor2_1 _5270_ (.Y(_1549_),
    .A(_1541_),
    .B(_1547_));
 sg13g2_nor2_1 _5271_ (.A(_2831_),
    .B(_1535_),
    .Y(_1550_));
 sg13g2_o21ai_1 _5272_ (.B1(_1533_),
    .Y(_1551_),
    .A1(_2831_),
    .A2(_1535_));
 sg13g2_xnor2_1 _5273_ (.Y(_1552_),
    .A(_1523_),
    .B(_1529_));
 sg13g2_xor2_1 _5274_ (.B(_1552_),
    .A(_1551_),
    .X(_1553_));
 sg13g2_inv_1 _5275_ (.Y(_1554_),
    .A(_1553_));
 sg13g2_xor2_1 _5276_ (.B(_1553_),
    .A(_1549_),
    .X(_1555_));
 sg13g2_nor2_1 _5277_ (.A(_1540_),
    .B(_1555_),
    .Y(_1556_));
 sg13g2_xor2_1 _5278_ (.B(_1555_),
    .A(_1540_),
    .X(\main.demo._d___pip_58_1_2___stage___block_3_cx[2] ));
 sg13g2_a21oi_1 _5279_ (.A1(_1549_),
    .A2(_1554_),
    .Y(_1557_),
    .B1(_1556_));
 sg13g2_a21oi_1 _5280_ (.A1(_1543_),
    .A2(_1546_),
    .Y(_1558_),
    .B1(_1548_));
 sg13g2_xor2_1 _5281_ (.B(_2742_),
    .A(_2741_),
    .X(_1559_));
 sg13g2_nor2_1 _5282_ (.A(_1525_),
    .B(_1544_),
    .Y(_1560_));
 sg13g2_nor2_1 _5283_ (.A(net351),
    .B(_1560_),
    .Y(_1561_));
 sg13g2_xnor2_1 _5284_ (.Y(_1562_),
    .A(_1521_),
    .B(_1561_));
 sg13g2_inv_1 _5285_ (.Y(_1563_),
    .A(_1562_));
 sg13g2_xnor2_1 _5286_ (.Y(_1564_),
    .A(_1559_),
    .B(_1562_));
 sg13g2_nand2b_1 _5287_ (.Y(_1565_),
    .B(_1564_),
    .A_N(_1558_));
 sg13g2_xnor2_1 _5288_ (.Y(_1566_),
    .A(_1558_),
    .B(_1564_));
 sg13g2_nand2_1 _5289_ (.Y(_1567_),
    .A(_1550_),
    .B(_1552_));
 sg13g2_nand2_1 _5290_ (.Y(_1568_),
    .A(_1533_),
    .B(_1567_));
 sg13g2_xnor2_1 _5291_ (.Y(_1569_),
    .A(_1520_),
    .B(_1530_));
 sg13g2_xor2_1 _5292_ (.B(_1569_),
    .A(_1568_),
    .X(_1570_));
 sg13g2_inv_1 _5293_ (.Y(_1571_),
    .A(_1570_));
 sg13g2_xor2_1 _5294_ (.B(_1570_),
    .A(_1566_),
    .X(_1572_));
 sg13g2_nor2_1 _5295_ (.A(_1557_),
    .B(_1572_),
    .Y(_1573_));
 sg13g2_xor2_1 _5296_ (.B(_1572_),
    .A(_1557_),
    .X(\main.demo._d___pip_58_1_2___stage___block_3_cx[3] ));
 sg13g2_a21oi_2 _5297_ (.B1(_1573_),
    .Y(_1574_),
    .A2(_1571_),
    .A1(_1566_));
 sg13g2_o21ai_1 _5298_ (.B1(_1565_),
    .Y(_1575_),
    .A1(_1559_),
    .A2(_1563_));
 sg13g2_nand2b_1 _5299_ (.Y(_1576_),
    .B(_1560_),
    .A_N(_1521_));
 sg13g2_nand2_1 _5300_ (.Y(_1577_),
    .A(net349),
    .B(_1576_));
 sg13g2_xor2_1 _5301_ (.B(_1577_),
    .A(_1518_),
    .X(_1578_));
 sg13g2_nor2_1 _5302_ (.A(_2770_),
    .B(_1578_),
    .Y(_1579_));
 sg13g2_xnor2_1 _5303_ (.Y(_1580_),
    .A(_2771_),
    .B(_1578_));
 sg13g2_xnor2_1 _5304_ (.Y(_1581_),
    .A(_1575_),
    .B(_1580_));
 sg13g2_nand2b_1 _5305_ (.Y(_1582_),
    .B(_1569_),
    .A_N(_1567_));
 sg13g2_nand2_1 _5306_ (.Y(_1583_),
    .A(_1533_),
    .B(_1582_));
 sg13g2_xor2_1 _5307_ (.B(_1515_),
    .A(_1512_),
    .X(_1584_));
 sg13g2_xnor2_1 _5308_ (.Y(_1585_),
    .A(_1531_),
    .B(_1584_));
 sg13g2_xnor2_1 _5309_ (.Y(_1586_),
    .A(_1583_),
    .B(_1585_));
 sg13g2_nor2_1 _5310_ (.A(_1581_),
    .B(_1586_),
    .Y(_1587_));
 sg13g2_xor2_1 _5311_ (.B(_1586_),
    .A(_1581_),
    .X(_1588_));
 sg13g2_nor2b_1 _5312_ (.A(_1574_),
    .B_N(_1588_),
    .Y(_1589_));
 sg13g2_xnor2_1 _5313_ (.Y(\main.demo._d___pip_58_1_2___stage___block_3_cx[4] ),
    .A(_1574_),
    .B(_1588_));
 sg13g2_nor2_2 _5314_ (.A(_1587_),
    .B(_1589_),
    .Y(_1590_));
 sg13g2_nor2_1 _5315_ (.A(_1582_),
    .B(_1585_),
    .Y(_1591_));
 sg13g2_nand2_2 _5316_ (.Y(_1592_),
    .A(_1533_),
    .B(_1591_));
 sg13g2_a21oi_2 _5317_ (.B1(_1579_),
    .Y(_1593_),
    .A2(_1580_),
    .A1(_1575_));
 sg13g2_nand2b_1 _5318_ (.Y(_1594_),
    .B(_1518_),
    .A_N(_1576_));
 sg13g2_nand2_1 _5319_ (.Y(_1595_),
    .A(net349),
    .B(_1594_));
 sg13g2_xor2_1 _5320_ (.B(_1595_),
    .A(_1515_),
    .X(_1596_));
 sg13g2_nand2_1 _5321_ (.Y(_1597_),
    .A(_2769_),
    .B(_1596_));
 sg13g2_xnor2_1 _5322_ (.Y(_1598_),
    .A(_2769_),
    .B(_1596_));
 sg13g2_xor2_1 _5323_ (.B(_1598_),
    .A(_1593_),
    .X(_1599_));
 sg13g2_inv_1 _5324_ (.Y(_1600_),
    .A(_1599_));
 sg13g2_xnor2_1 _5325_ (.Y(_1601_),
    .A(net341),
    .B(_1599_));
 sg13g2_xnor2_1 _5326_ (.Y(\main.demo._d___pip_58_1_2___stage___block_3_cx[5] ),
    .A(_1590_),
    .B(_1601_));
 sg13g2_a21oi_1 _5327_ (.A1(net341),
    .A2(_1600_),
    .Y(_1602_),
    .B1(_1590_));
 sg13g2_nor3_2 _5328_ (.A(net351),
    .B(_1515_),
    .C(_1594_),
    .Y(_1603_));
 sg13g2_xnor2_1 _5329_ (.Y(_1604_),
    .A(_2768_),
    .B(_1603_));
 sg13g2_o21ai_1 _5330_ (.B1(_1597_),
    .Y(_1605_),
    .A1(_1593_),
    .A2(_1598_));
 sg13g2_nor2b_1 _5331_ (.A(_1604_),
    .B_N(_1605_),
    .Y(_1606_));
 sg13g2_xor2_1 _5332_ (.B(_1605_),
    .A(_1604_),
    .X(_1607_));
 sg13g2_nor2_1 _5333_ (.A(net341),
    .B(_1607_),
    .Y(_1608_));
 sg13g2_xor2_1 _5334_ (.B(_1607_),
    .A(net341),
    .X(_1609_));
 sg13g2_xor2_1 _5335_ (.B(_1609_),
    .A(_1602_),
    .X(\main.demo._d___pip_58_1_2___stage___block_3_cx[6] ));
 sg13g2_a21oi_1 _5336_ (.A1(_1602_),
    .A2(_1609_),
    .Y(_1610_),
    .B1(_1608_));
 sg13g2_nand2_1 _5337_ (.Y(_1611_),
    .A(_2774_),
    .B(net343));
 sg13g2_xnor2_1 _5338_ (.Y(_1612_),
    .A(_2774_),
    .B(net343));
 sg13g2_a21oi_1 _5339_ (.A1(_2768_),
    .A2(net343),
    .Y(_1613_),
    .B1(_1606_));
 sg13g2_xnor2_1 _5340_ (.Y(_1614_),
    .A(_1612_),
    .B(_1613_));
 sg13g2_nor2_1 _5341_ (.A(net341),
    .B(_1614_),
    .Y(_1615_));
 sg13g2_xor2_1 _5342_ (.B(_1614_),
    .A(_1592_),
    .X(_1616_));
 sg13g2_nor2b_1 _5343_ (.A(_1610_),
    .B_N(_1616_),
    .Y(_1617_));
 sg13g2_xnor2_1 _5344_ (.Y(\main.demo._d___pip_58_1_2___stage___block_3_cx[7] ),
    .A(_1610_),
    .B(_1616_));
 sg13g2_nor2b_1 _5345_ (.A(_2777_),
    .B_N(net343),
    .Y(_1618_));
 sg13g2_xnor2_1 _5346_ (.Y(_1619_),
    .A(_2777_),
    .B(net343));
 sg13g2_o21ai_1 _5347_ (.B1(_1611_),
    .Y(_1620_),
    .A1(_1612_),
    .A2(_1613_));
 sg13g2_xor2_1 _5348_ (.B(_1620_),
    .A(_1619_),
    .X(_1621_));
 sg13g2_inv_1 _5349_ (.Y(_1622_),
    .A(_1621_));
 sg13g2_xnor2_1 _5350_ (.Y(_1623_),
    .A(_1592_),
    .B(_1621_));
 sg13g2_o21ai_1 _5351_ (.B1(_1623_),
    .Y(_1624_),
    .A1(_1615_),
    .A2(_1617_));
 sg13g2_or3_1 _5352_ (.A(_1615_),
    .B(_1617_),
    .C(_1623_),
    .X(_1625_));
 sg13g2_and2_1 _5353_ (.A(_1624_),
    .B(_1625_),
    .X(\main.demo._d___pip_58_1_2___stage___block_3_cx[8] ));
 sg13g2_nor2_1 _5354_ (.A(_2767_),
    .B(net343),
    .Y(_1626_));
 sg13g2_xnor2_1 _5355_ (.Y(_1627_),
    .A(_2767_),
    .B(net343));
 sg13g2_a21oi_1 _5356_ (.A1(_1619_),
    .A2(_1620_),
    .Y(_1628_),
    .B1(_1618_));
 sg13g2_xnor2_1 _5357_ (.Y(_1629_),
    .A(_1627_),
    .B(_1628_));
 sg13g2_xnor2_1 _5358_ (.Y(_1630_),
    .A(net341),
    .B(_1629_));
 sg13g2_o21ai_1 _5359_ (.B1(_1624_),
    .Y(_1631_),
    .A1(net341),
    .A2(_1622_));
 sg13g2_xnor2_1 _5360_ (.Y(\main.demo._d___pip_58_1_2___stage___block_3_cx[9] ),
    .A(_1630_),
    .B(_1631_));
 sg13g2_nand3b_1 _5361_ (.B(_1631_),
    .C(net341),
    .Y(_1632_),
    .A_N(_1629_));
 sg13g2_nor2_1 _5362_ (.A(_1626_),
    .B(_1628_),
    .Y(_1633_));
 sg13g2_xor2_1 _5363_ (.B(net343),
    .A(_1508_),
    .X(_1634_));
 sg13g2_xnor2_1 _5364_ (.Y(_1635_),
    .A(_1633_),
    .B(_1634_));
 sg13g2_xnor2_1 _5365_ (.Y(\main.demo._d___pip_58_1_2___stage___block_3_cx[10] ),
    .A(_1632_),
    .B(_1635_));
 sg13g2_xor2_1 _5366_ (.B(\main.demo._q___pip_58_1_2___stage___block_3_a[1] ),
    .A(net449),
    .X(_1636_));
 sg13g2_nor2b_1 _5367_ (.A(_1533_),
    .B_N(_1636_),
    .Y(_1637_));
 sg13g2_xnor2_1 _5368_ (.Y(\main.demo._d___pip_58_1_2___stage___block_3_a[1] ),
    .A(_1533_),
    .B(_1636_));
 sg13g2_a21oi_2 _5369_ (.B1(\main.demo._q___pip_58_1_2___stage___block_3_a[2] ),
    .Y(_1638_),
    .A2(\main.demo._q___pip_58_1_2___stage___block_3_a[1] ),
    .A1(net449));
 sg13g2_nand3_1 _5370_ (.B(\main.demo._q___pip_58_1_2___stage___block_3_a[1] ),
    .C(\main.demo._q___pip_58_1_2___stage___block_3_a[2] ),
    .A(net449),
    .Y(_1639_));
 sg13g2_nand2b_1 _5371_ (.Y(_1640_),
    .B(_1639_),
    .A_N(_1638_));
 sg13g2_inv_1 _5372_ (.Y(_1641_),
    .A(_1640_));
 sg13g2_xnor2_1 _5373_ (.Y(_1642_),
    .A(net352),
    .B(_1641_));
 sg13g2_xnor2_1 _5374_ (.Y(\main.demo._d___pip_58_1_2___stage___block_3_a[2] ),
    .A(_1637_),
    .B(_1642_));
 sg13g2_nand2b_1 _5375_ (.Y(_1643_),
    .B(_1636_),
    .A_N(_1642_));
 sg13g2_nand2b_1 _5376_ (.Y(_1644_),
    .B(_1533_),
    .A_N(_1643_));
 sg13g2_o21ai_1 _5377_ (.B1(_1643_),
    .Y(_1645_),
    .A1(net352),
    .A2(_1641_));
 sg13g2_nand2_1 _5378_ (.Y(_1646_),
    .A(_2621_),
    .B(\main.demo._q___pip_58_1_2___stage___block_3_a[3] ));
 sg13g2_nor2_1 _5379_ (.A(net404),
    .B(\main.demo._q___pip_58_1_2___stage___block_3_a[3] ),
    .Y(_1647_));
 sg13g2_xnor2_1 _5380_ (.Y(_1648_),
    .A(net450),
    .B(\main.demo._q___pip_58_1_2___stage___block_3_a[3] ));
 sg13g2_xnor2_1 _5381_ (.Y(_1649_),
    .A(_1638_),
    .B(_1648_));
 sg13g2_and2_1 _5382_ (.A(net350),
    .B(_1649_),
    .X(_1650_));
 sg13g2_xnor2_1 _5383_ (.Y(_1651_),
    .A(net352),
    .B(_1649_));
 sg13g2_xor2_1 _5384_ (.B(_1651_),
    .A(_1645_),
    .X(_1652_));
 sg13g2_nand2b_1 _5385_ (.Y(_1653_),
    .B(_1651_),
    .A_N(_1644_));
 sg13g2_xnor2_1 _5386_ (.Y(\main.demo._d___pip_58_1_2___stage___block_3_a[3] ),
    .A(_1644_),
    .B(_1652_));
 sg13g2_xor2_1 _5387_ (.B(\main.demo._q___pip_58_1_2___stage___block_3_a[4] ),
    .A(net449),
    .X(_1654_));
 sg13g2_o21ai_1 _5388_ (.B1(_1646_),
    .Y(_1655_),
    .A1(_1638_),
    .A2(_1647_));
 sg13g2_xnor2_1 _5389_ (.Y(_1656_),
    .A(_1654_),
    .B(_1655_));
 sg13g2_nand2_1 _5390_ (.Y(_1657_),
    .A(net350),
    .B(_1656_));
 sg13g2_nor2_1 _5391_ (.A(net350),
    .B(_1656_),
    .Y(_1658_));
 sg13g2_xnor2_1 _5392_ (.Y(_1659_),
    .A(net352),
    .B(_1656_));
 sg13g2_a21oi_1 _5393_ (.A1(_1645_),
    .A2(_1651_),
    .Y(_1660_),
    .B1(_1650_));
 sg13g2_xnor2_1 _5394_ (.Y(_1661_),
    .A(_1659_),
    .B(_1660_));
 sg13g2_or2_1 _5395_ (.X(_1662_),
    .B(_1661_),
    .A(_1653_));
 sg13g2_xnor2_1 _5396_ (.Y(\main.demo._d___pip_58_1_2___stage___block_3_a[4] ),
    .A(_1653_),
    .B(_1661_));
 sg13g2_o21ai_1 _5397_ (.B1(_1655_),
    .Y(_1663_),
    .A1(net404),
    .A2(\main.demo._q___pip_58_1_2___stage___block_3_a[4] ));
 sg13g2_o21ai_1 _5398_ (.B1(_1663_),
    .Y(_1664_),
    .A1(net449),
    .A2(_2668_));
 sg13g2_a21oi_2 _5399_ (.B1(_1647_),
    .Y(_1665_),
    .A2(_1664_),
    .A1(_1646_));
 sg13g2_nand2_1 _5400_ (.Y(_1666_),
    .A(net350),
    .B(_1665_));
 sg13g2_o21ai_1 _5401_ (.B1(_1657_),
    .Y(_1667_),
    .A1(_1658_),
    .A2(_1660_));
 sg13g2_nand2_1 _5402_ (.Y(_1668_),
    .A(_1666_),
    .B(_1667_));
 sg13g2_o21ai_1 _5403_ (.B1(_1668_),
    .Y(_1669_),
    .A1(net350),
    .A2(_1665_));
 sg13g2_nand2_1 _5404_ (.Y(\main.demo._d___pip_58_1_2___stage___block_3_a[5] ),
    .A(_1662_),
    .B(_1669_));
 sg13g2_xor2_1 _5405_ (.B(\main.demo._q___pip_58_1_2___stage___block_3_a[6] ),
    .A(net449),
    .X(_1670_));
 sg13g2_xnor2_1 _5406_ (.Y(_1671_),
    .A(_1664_),
    .B(_1670_));
 sg13g2_nor2_1 _5407_ (.A(net349),
    .B(_1671_),
    .Y(_1672_));
 sg13g2_xnor2_1 _5408_ (.Y(_1673_),
    .A(net349),
    .B(_1671_));
 sg13g2_xnor2_1 _5409_ (.Y(_1674_),
    .A(_1667_),
    .B(_1673_));
 sg13g2_nor2_1 _5410_ (.A(_1662_),
    .B(_1674_),
    .Y(_1675_));
 sg13g2_xnor2_1 _5411_ (.Y(\main.demo._d___pip_58_1_2___stage___block_3_a[6] ),
    .A(_1662_),
    .B(_1674_));
 sg13g2_o21ai_1 _5412_ (.B1(net349),
    .Y(_1676_),
    .A1(_1665_),
    .A2(_1671_));
 sg13g2_o21ai_1 _5413_ (.B1(_1676_),
    .Y(_1677_),
    .A1(_1668_),
    .A2(_1672_));
 sg13g2_nor3_1 _5414_ (.A(net449),
    .B(\main.demo._q___pip_58_1_2___stage___block_3_a[6] ),
    .C(_1664_),
    .Y(_1678_));
 sg13g2_nand4_1 _5415_ (.B(\main.demo._q___pip_58_1_2___stage___block_3_a[4] ),
    .C(\main.demo._q___pip_58_1_2___stage___block_3_a[6] ),
    .A(net449),
    .Y(_1679_),
    .D(_1655_));
 sg13g2_nor2b_1 _5416_ (.A(_1678_),
    .B_N(_1679_),
    .Y(_1680_));
 sg13g2_xnor2_1 _5417_ (.Y(_1681_),
    .A(\main.demo._q___pip_58_1_2___stage___block_3_a[7] ),
    .B(_1680_));
 sg13g2_xnor2_1 _5418_ (.Y(_1682_),
    .A(net352),
    .B(_1681_));
 sg13g2_xnor2_1 _5419_ (.Y(_1683_),
    .A(_1677_),
    .B(_1682_));
 sg13g2_xnor2_1 _5420_ (.Y(\main.demo._d___pip_58_1_2___stage___block_3_a[7] ),
    .A(_1675_),
    .B(_1683_));
 sg13g2_nor2_1 _5421_ (.A(net433),
    .B(_0068_),
    .Y(_1684_));
 sg13g2_xnor2_1 _5422_ (.Y(\main.demo._d___pip_58_1_1___stage___block_3_a[6] ),
    .A(net433),
    .B(net294));
 sg13g2_xor2_1 _5423_ (.B(_1684_),
    .A(net287),
    .X(\main.demo._d___pip_58_1_1___stage___block_3_a[7] ));
 sg13g2_nor2_1 _5424_ (.A(net347),
    .B(_2905_),
    .Y(_1685_));
 sg13g2_xnor2_1 _5425_ (.Y(_1686_),
    .A(_2923_),
    .B(_1685_));
 sg13g2_xor2_1 _5426_ (.B(_1686_),
    .A(_2909_),
    .X(_1687_));
 sg13g2_nand2_1 _5427_ (.Y(_1688_),
    .A(_2906_),
    .B(_1687_));
 sg13g2_xnor2_1 _5428_ (.Y(_1689_),
    .A(_2906_),
    .B(_1687_));
 sg13g2_nand2_1 _5429_ (.Y(_1690_),
    .A(_2934_),
    .B(_0415_));
 sg13g2_xnor2_1 _5430_ (.Y(_1691_),
    .A(_0398_),
    .B(_0399_));
 sg13g2_xnor2_1 _5431_ (.Y(_1692_),
    .A(_1690_),
    .B(_1691_));
 sg13g2_nor2_1 _5432_ (.A(_1689_),
    .B(_1692_),
    .Y(_1693_));
 sg13g2_xor2_1 _5433_ (.B(_1692_),
    .A(_1689_),
    .X(_1694_));
 sg13g2_xor2_1 _5434_ (.B(_1694_),
    .A(_2935_),
    .X(\main.demo._d___pip_58_1_1___stage___block_3_cx[1] ));
 sg13g2_a21oi_1 _5435_ (.A1(_2935_),
    .A2(_1694_),
    .Y(_1695_),
    .B1(_1693_));
 sg13g2_o21ai_1 _5436_ (.B1(_1688_),
    .Y(_1696_),
    .A1(_2909_),
    .A2(_1686_));
 sg13g2_nand2_1 _5437_ (.Y(_1697_),
    .A(_2905_),
    .B(_2923_));
 sg13g2_nand2_1 _5438_ (.Y(_1698_),
    .A(\main.demo._d___pip_58_1_1___stage___block_3_a[2] ),
    .B(_1697_));
 sg13g2_xor2_1 _5439_ (.B(_1698_),
    .A(_0395_),
    .X(_1699_));
 sg13g2_nor2b_1 _5440_ (.A(_2915_),
    .B_N(_1699_),
    .Y(_1700_));
 sg13g2_xnor2_1 _5441_ (.Y(_1701_),
    .A(_2915_),
    .B(_1699_));
 sg13g2_xnor2_1 _5442_ (.Y(_1702_),
    .A(_1696_),
    .B(_1701_));
 sg13g2_inv_1 _5443_ (.Y(_1703_),
    .A(_1702_));
 sg13g2_nor2_1 _5444_ (.A(_2934_),
    .B(_1691_),
    .Y(_1704_));
 sg13g2_nor2_1 _5445_ (.A(net340),
    .B(_1704_),
    .Y(_1705_));
 sg13g2_xnor2_1 _5446_ (.Y(_1706_),
    .A(_0393_),
    .B(_0401_));
 sg13g2_xor2_1 _5447_ (.B(_1706_),
    .A(_1705_),
    .X(_1707_));
 sg13g2_xnor2_1 _5448_ (.Y(_1708_),
    .A(_1703_),
    .B(_1707_));
 sg13g2_nor2_1 _5449_ (.A(_1695_),
    .B(_1708_),
    .Y(_1709_));
 sg13g2_xor2_1 _5450_ (.B(_1708_),
    .A(_1695_),
    .X(\main.demo._d___pip_58_1_1___stage___block_3_cx[2] ));
 sg13g2_a21oi_1 _5451_ (.A1(_1703_),
    .A2(_1707_),
    .Y(_1710_),
    .B1(_1709_));
 sg13g2_a21o_1 _5452_ (.A2(_1701_),
    .A1(_1696_),
    .B1(_1700_),
    .X(_1711_));
 sg13g2_nor2_1 _5453_ (.A(_0395_),
    .B(_1697_),
    .Y(_1712_));
 sg13g2_nor2_1 _5454_ (.A(net348),
    .B(_1712_),
    .Y(_1713_));
 sg13g2_xnor2_1 _5455_ (.Y(_1714_),
    .A(_0388_),
    .B(_1713_));
 sg13g2_xnor2_1 _5456_ (.Y(_1715_),
    .A(_2929_),
    .B(_1714_));
 sg13g2_nand2_1 _5457_ (.Y(_1716_),
    .A(_1711_),
    .B(_1715_));
 sg13g2_xor2_1 _5458_ (.B(_1715_),
    .A(_1711_),
    .X(_1717_));
 sg13g2_nand2_1 _5459_ (.Y(_1718_),
    .A(_1704_),
    .B(_1706_));
 sg13g2_nand2_1 _5460_ (.Y(_1719_),
    .A(_0415_),
    .B(_1718_));
 sg13g2_xnor2_1 _5461_ (.Y(_1720_),
    .A(_0402_),
    .B(_0403_));
 sg13g2_xnor2_1 _5462_ (.Y(_1721_),
    .A(_1719_),
    .B(_1720_));
 sg13g2_inv_1 _5463_ (.Y(_1722_),
    .A(_1721_));
 sg13g2_xor2_1 _5464_ (.B(_1721_),
    .A(_1717_),
    .X(_1723_));
 sg13g2_nor2_1 _5465_ (.A(_1710_),
    .B(_1723_),
    .Y(_1724_));
 sg13g2_xor2_1 _5466_ (.B(_1723_),
    .A(_1710_),
    .X(\main.demo._d___pip_58_1_1___stage___block_3_cx[3] ));
 sg13g2_a21oi_1 _5467_ (.A1(_1717_),
    .A2(_1722_),
    .Y(_1725_),
    .B1(_1724_));
 sg13g2_o21ai_1 _5468_ (.B1(_1716_),
    .Y(_1726_),
    .A1(_2930_),
    .A2(_1714_));
 sg13g2_nand2_1 _5469_ (.Y(_1727_),
    .A(_0388_),
    .B(_1712_));
 sg13g2_nand2_1 _5470_ (.Y(_1728_),
    .A(net344),
    .B(_1727_));
 sg13g2_xor2_1 _5471_ (.B(_1728_),
    .A(_0384_),
    .X(_1729_));
 sg13g2_nor2b_1 _5472_ (.A(_0331_),
    .B_N(_1729_),
    .Y(_1730_));
 sg13g2_xnor2_1 _5473_ (.Y(_1731_),
    .A(_0331_),
    .B(_1729_));
 sg13g2_xor2_1 _5474_ (.B(_1731_),
    .A(_1726_),
    .X(_1732_));
 sg13g2_nor2_1 _5475_ (.A(_1718_),
    .B(_1720_),
    .Y(_1733_));
 sg13g2_nor2_1 _5476_ (.A(net339),
    .B(_1733_),
    .Y(_1734_));
 sg13g2_xor2_1 _5477_ (.B(_0405_),
    .A(_0381_),
    .X(_1735_));
 sg13g2_xor2_1 _5478_ (.B(_1735_),
    .A(_1734_),
    .X(_1736_));
 sg13g2_xnor2_1 _5479_ (.Y(_1737_),
    .A(_1732_),
    .B(_1736_));
 sg13g2_nor2_1 _5480_ (.A(_1725_),
    .B(_1737_),
    .Y(_1738_));
 sg13g2_xor2_1 _5481_ (.B(_1737_),
    .A(_1725_),
    .X(\main.demo._d___pip_58_1_1___stage___block_3_cx[4] ));
 sg13g2_a21oi_1 _5482_ (.A1(_1732_),
    .A2(_1736_),
    .Y(_1739_),
    .B1(_1738_));
 sg13g2_a21o_1 _5483_ (.A2(_1731_),
    .A1(_1726_),
    .B1(_1730_),
    .X(_1740_));
 sg13g2_nor2_1 _5484_ (.A(_0384_),
    .B(_1727_),
    .Y(_1741_));
 sg13g2_nor2_1 _5485_ (.A(net347),
    .B(_1741_),
    .Y(_1742_));
 sg13g2_xnor2_1 _5486_ (.Y(_1743_),
    .A(_0376_),
    .B(_1742_));
 sg13g2_xnor2_1 _5487_ (.Y(_1744_),
    .A(_0335_),
    .B(_1743_));
 sg13g2_nand2_1 _5488_ (.Y(_1745_),
    .A(_1740_),
    .B(_1744_));
 sg13g2_xor2_1 _5489_ (.B(_1744_),
    .A(_1740_),
    .X(_1746_));
 sg13g2_nand2_1 _5490_ (.Y(_1747_),
    .A(_1733_),
    .B(_1735_));
 sg13g2_nand2_1 _5491_ (.Y(_1748_),
    .A(_0415_),
    .B(_1747_));
 sg13g2_xnor2_1 _5492_ (.Y(_1749_),
    .A(_0406_),
    .B(_0407_));
 sg13g2_xnor2_1 _5493_ (.Y(_1750_),
    .A(_1748_),
    .B(_1749_));
 sg13g2_inv_1 _5494_ (.Y(_1751_),
    .A(_1750_));
 sg13g2_xor2_1 _5495_ (.B(_1750_),
    .A(_1746_),
    .X(_1752_));
 sg13g2_nor2_1 _5496_ (.A(_1739_),
    .B(_1752_),
    .Y(_1753_));
 sg13g2_xor2_1 _5497_ (.B(_1752_),
    .A(_1739_),
    .X(\main.demo._d___pip_58_1_1___stage___block_3_cx[5] ));
 sg13g2_a21oi_1 _5498_ (.A1(_1746_),
    .A2(_1751_),
    .Y(_1754_),
    .B1(_1753_));
 sg13g2_o21ai_1 _5499_ (.B1(_1745_),
    .Y(_1755_),
    .A1(_0336_),
    .A2(_1743_));
 sg13g2_nand2_1 _5500_ (.Y(_1756_),
    .A(_0376_),
    .B(_1741_));
 sg13g2_nand2_1 _5501_ (.Y(_1757_),
    .A(net344),
    .B(_1756_));
 sg13g2_xor2_1 _5502_ (.B(_1757_),
    .A(_0372_),
    .X(_1758_));
 sg13g2_nor2b_1 _5503_ (.A(_0342_),
    .B_N(_1758_),
    .Y(_1759_));
 sg13g2_xnor2_1 _5504_ (.Y(_1760_),
    .A(_0342_),
    .B(_1758_));
 sg13g2_xor2_1 _5505_ (.B(_1760_),
    .A(_1755_),
    .X(_1761_));
 sg13g2_nor2_1 _5506_ (.A(_1747_),
    .B(_1749_),
    .Y(_1762_));
 sg13g2_nor2_1 _5507_ (.A(net339),
    .B(_1762_),
    .Y(_1763_));
 sg13g2_xnor2_1 _5508_ (.Y(_1764_),
    .A(_0409_),
    .B(_0410_));
 sg13g2_xor2_1 _5509_ (.B(_1764_),
    .A(_1763_),
    .X(_1765_));
 sg13g2_xnor2_1 _5510_ (.Y(_1766_),
    .A(_1761_),
    .B(_1765_));
 sg13g2_nor2_1 _5511_ (.A(_1754_),
    .B(_1766_),
    .Y(_1767_));
 sg13g2_xor2_1 _5512_ (.B(_1766_),
    .A(_1754_),
    .X(\main.demo._d___pip_58_1_1___stage___block_3_cx[6] ));
 sg13g2_a21oi_1 _5513_ (.A1(_1761_),
    .A2(_1765_),
    .Y(_1768_),
    .B1(_1767_));
 sg13g2_a21o_1 _5514_ (.A2(_1760_),
    .A1(_1755_),
    .B1(_1759_),
    .X(_1769_));
 sg13g2_nor2_1 _5515_ (.A(_0372_),
    .B(_1756_),
    .Y(_1770_));
 sg13g2_nor2_1 _5516_ (.A(net347),
    .B(_1770_),
    .Y(_1771_));
 sg13g2_xnor2_1 _5517_ (.Y(_1772_),
    .A(_0365_),
    .B(_1771_));
 sg13g2_xor2_1 _5518_ (.B(_1772_),
    .A(_0345_),
    .X(_1773_));
 sg13g2_nand2_1 _5519_ (.Y(_1774_),
    .A(_1769_),
    .B(_1773_));
 sg13g2_xor2_1 _5520_ (.B(_1773_),
    .A(_1769_),
    .X(_1775_));
 sg13g2_nand2_1 _5521_ (.Y(_1776_),
    .A(_1762_),
    .B(_1764_));
 sg13g2_nand2_1 _5522_ (.Y(_1777_),
    .A(_0415_),
    .B(_1776_));
 sg13g2_xnor2_1 _5523_ (.Y(_1778_),
    .A(_0411_),
    .B(_0412_));
 sg13g2_xnor2_1 _5524_ (.Y(_1779_),
    .A(_1777_),
    .B(_1778_));
 sg13g2_inv_1 _5525_ (.Y(_1780_),
    .A(_1779_));
 sg13g2_xor2_1 _5526_ (.B(_1779_),
    .A(_1775_),
    .X(_1781_));
 sg13g2_nor2_1 _5527_ (.A(_1768_),
    .B(_1781_),
    .Y(_1782_));
 sg13g2_xor2_1 _5528_ (.B(_1781_),
    .A(_1768_),
    .X(\main.demo._d___pip_58_1_1___stage___block_3_cx[7] ));
 sg13g2_a21oi_1 _5529_ (.A1(_1775_),
    .A2(_1780_),
    .Y(_1783_),
    .B1(_1782_));
 sg13g2_or3_1 _5530_ (.A(net339),
    .B(_1776_),
    .C(_1778_),
    .X(_1784_));
 sg13g2_o21ai_1 _5531_ (.B1(_1774_),
    .Y(_1785_),
    .A1(_0345_),
    .A2(_1772_));
 sg13g2_a21oi_1 _5532_ (.A1(_0365_),
    .A2(_1770_),
    .Y(_1786_),
    .B1(net347));
 sg13g2_xor2_1 _5533_ (.B(_1786_),
    .A(_0361_),
    .X(_1787_));
 sg13g2_and2_1 _5534_ (.A(_0349_),
    .B(_1787_),
    .X(_1788_));
 sg13g2_xnor2_1 _5535_ (.Y(_1789_),
    .A(_0350_),
    .B(_1787_));
 sg13g2_xor2_1 _5536_ (.B(_1789_),
    .A(_1785_),
    .X(_1790_));
 sg13g2_xnor2_1 _5537_ (.Y(_1791_),
    .A(_1784_),
    .B(_1790_));
 sg13g2_nor2b_1 _5538_ (.A(_1783_),
    .B_N(_1791_),
    .Y(_1792_));
 sg13g2_xnor2_1 _5539_ (.Y(\main.demo._d___pip_58_1_1___stage___block_3_cx[8] ),
    .A(_1783_),
    .B(_1791_));
 sg13g2_nand4_1 _5540_ (.B(_0361_),
    .C(_0365_),
    .A(net344),
    .Y(_1793_),
    .D(_1770_));
 sg13g2_a21oi_1 _5541_ (.A1(_1785_),
    .A2(_1789_),
    .Y(_1794_),
    .B1(_1788_));
 sg13g2_inv_1 _5542_ (.Y(_1795_),
    .A(_1794_));
 sg13g2_xnor2_1 _5543_ (.Y(_1796_),
    .A(_0354_),
    .B(_1794_));
 sg13g2_xnor2_1 _5544_ (.Y(_1797_),
    .A(_1793_),
    .B(_1796_));
 sg13g2_nand3_1 _5545_ (.B(_1792_),
    .C(_1797_),
    .A(_1784_),
    .Y(_1798_));
 sg13g2_a21o_1 _5546_ (.A2(_1792_),
    .A1(_1784_),
    .B1(_1797_),
    .X(_1799_));
 sg13g2_and2_1 _5547_ (.A(_1798_),
    .B(_1799_),
    .X(\main.demo._d___pip_58_1_1___stage___block_3_cx[9] ));
 sg13g2_nand3_1 _5548_ (.B(_1793_),
    .C(_1795_),
    .A(_0354_),
    .Y(_1800_));
 sg13g2_xnor2_1 _5549_ (.Y(_1801_),
    .A(_0357_),
    .B(_1800_));
 sg13g2_xnor2_1 _5550_ (.Y(\main.demo._d___pip_58_1_1___stage___block_3_cx[10] ),
    .A(_1798_),
    .B(_1801_));
 sg13g2_xor2_1 _5551_ (.B(_2909_),
    .A(_2902_),
    .X(_1802_));
 sg13g2_nand2_1 _5552_ (.Y(_1803_),
    .A(_1703_),
    .B(_1802_));
 sg13g2_xnor2_1 _5553_ (.Y(\main.demo._d___pip_58_1_1___stage___block_3_cy[0] ),
    .A(_1702_),
    .B(_1802_));
 sg13g2_xor2_1 _5554_ (.B(_2919_),
    .A(_2918_),
    .X(_1804_));
 sg13g2_nor2_1 _5555_ (.A(net340),
    .B(_1702_),
    .Y(_1805_));
 sg13g2_xor2_1 _5556_ (.B(_1805_),
    .A(_1717_),
    .X(_1806_));
 sg13g2_xor2_1 _5557_ (.B(_1806_),
    .A(_1804_),
    .X(_1807_));
 sg13g2_nor2b_1 _5558_ (.A(_1803_),
    .B_N(_1807_),
    .Y(_1808_));
 sg13g2_xnor2_1 _5559_ (.Y(\main.demo._d___pip_58_1_1___stage___block_3_cy[1] ),
    .A(_1803_),
    .B(_1807_));
 sg13g2_nor2_1 _5560_ (.A(_1703_),
    .B(_1717_),
    .Y(_1809_));
 sg13g2_nor2_1 _5561_ (.A(net340),
    .B(_1809_),
    .Y(_1810_));
 sg13g2_xnor2_1 _5562_ (.Y(_1811_),
    .A(_1732_),
    .B(_1810_));
 sg13g2_nand2b_1 _5563_ (.Y(_1812_),
    .B(_2934_),
    .A_N(_1811_));
 sg13g2_xnor2_1 _5564_ (.Y(_1813_),
    .A(_2934_),
    .B(_1811_));
 sg13g2_inv_1 _5565_ (.Y(_1814_),
    .A(_1813_));
 sg13g2_a21oi_1 _5566_ (.A1(_1804_),
    .A2(_1806_),
    .Y(_1815_),
    .B1(_1808_));
 sg13g2_xnor2_1 _5567_ (.Y(\main.demo._d___pip_58_1_1___stage___block_3_cy[2] ),
    .A(_1813_),
    .B(_1815_));
 sg13g2_o21ai_1 _5568_ (.B1(_1812_),
    .Y(_1816_),
    .A1(_1814_),
    .A2(_1815_));
 sg13g2_nor2b_1 _5569_ (.A(_1732_),
    .B_N(_1809_),
    .Y(_1817_));
 sg13g2_nor2_1 _5570_ (.A(net340),
    .B(_1817_),
    .Y(_1818_));
 sg13g2_xor2_1 _5571_ (.B(_1818_),
    .A(_1746_),
    .X(_1819_));
 sg13g2_xnor2_1 _5572_ (.Y(_1820_),
    .A(_1691_),
    .B(_1819_));
 sg13g2_nor2b_1 _5573_ (.A(_1820_),
    .B_N(_1816_),
    .Y(_1821_));
 sg13g2_xnor2_1 _5574_ (.Y(\main.demo._d___pip_58_1_1___stage___block_3_cy[3] ),
    .A(_1816_),
    .B(_1820_));
 sg13g2_nor2b_1 _5575_ (.A(_1746_),
    .B_N(_1817_),
    .Y(_1822_));
 sg13g2_nor2_1 _5576_ (.A(net339),
    .B(_1822_),
    .Y(_1823_));
 sg13g2_xnor2_1 _5577_ (.Y(_1824_),
    .A(_1761_),
    .B(_1823_));
 sg13g2_nor2_1 _5578_ (.A(_1706_),
    .B(_1824_),
    .Y(_1825_));
 sg13g2_xnor2_1 _5579_ (.Y(_1826_),
    .A(_1706_),
    .B(_1824_));
 sg13g2_inv_1 _5580_ (.Y(_1827_),
    .A(_1826_));
 sg13g2_a21o_1 _5581_ (.A2(_1819_),
    .A1(_1691_),
    .B1(_1821_),
    .X(_1828_));
 sg13g2_xnor2_1 _5582_ (.Y(\main.demo._d___pip_58_1_1___stage___block_3_cy[4] ),
    .A(_1826_),
    .B(_1828_));
 sg13g2_a21oi_1 _5583_ (.A1(_1827_),
    .A2(_1828_),
    .Y(_1829_),
    .B1(_1825_));
 sg13g2_nor2b_1 _5584_ (.A(_1761_),
    .B_N(_1822_),
    .Y(_1830_));
 sg13g2_nor2_1 _5585_ (.A(net339),
    .B(_1830_),
    .Y(_1831_));
 sg13g2_xor2_1 _5586_ (.B(_1831_),
    .A(_1775_),
    .X(_1832_));
 sg13g2_nand2_1 _5587_ (.Y(_1833_),
    .A(_1720_),
    .B(_1832_));
 sg13g2_xnor2_1 _5588_ (.Y(_1834_),
    .A(_1720_),
    .B(_1832_));
 sg13g2_xor2_1 _5589_ (.B(_1834_),
    .A(_1829_),
    .X(\main.demo._d___pip_58_1_1___stage___block_3_cy[5] ));
 sg13g2_nor2b_1 _5590_ (.A(_1775_),
    .B_N(_1830_),
    .Y(_1835_));
 sg13g2_nor2_1 _5591_ (.A(net339),
    .B(_1835_),
    .Y(_1836_));
 sg13g2_xnor2_1 _5592_ (.Y(_1837_),
    .A(_1790_),
    .B(_1836_));
 sg13g2_nor2_1 _5593_ (.A(_1735_),
    .B(_1837_),
    .Y(_1838_));
 sg13g2_nand2_1 _5594_ (.Y(_1839_),
    .A(_1735_),
    .B(_1837_));
 sg13g2_nand2b_1 _5595_ (.Y(_1840_),
    .B(_1839_),
    .A_N(_1838_));
 sg13g2_o21ai_1 _5596_ (.B1(_1833_),
    .Y(_1841_),
    .A1(_1829_),
    .A2(_1834_));
 sg13g2_xnor2_1 _5597_ (.Y(\main.demo._d___pip_58_1_1___stage___block_3_cy[6] ),
    .A(_1840_),
    .B(_1841_));
 sg13g2_a21oi_2 _5598_ (.B1(_1838_),
    .Y(_1842_),
    .A2(_1841_),
    .A1(_1839_));
 sg13g2_nor2b_1 _5599_ (.A(_1790_),
    .B_N(_1835_),
    .Y(_1843_));
 sg13g2_nor2_1 _5600_ (.A(net339),
    .B(_1843_),
    .Y(_1844_));
 sg13g2_xnor2_1 _5601_ (.Y(_1845_),
    .A(_1797_),
    .B(_1844_));
 sg13g2_inv_1 _5602_ (.Y(_1846_),
    .A(_1845_));
 sg13g2_nand2_1 _5603_ (.Y(_1847_),
    .A(_1749_),
    .B(_1846_));
 sg13g2_xor2_1 _5604_ (.B(_1845_),
    .A(_1749_),
    .X(_1848_));
 sg13g2_xor2_1 _5605_ (.B(_1848_),
    .A(_1842_),
    .X(\main.demo._d___pip_58_1_1___stage___block_3_cy[7] ));
 sg13g2_nor2_1 _5606_ (.A(_0415_),
    .B(_1801_),
    .Y(_1849_));
 sg13g2_nor2b_1 _5607_ (.A(_1797_),
    .B_N(_1843_),
    .Y(_1850_));
 sg13g2_o21ai_1 _5608_ (.B1(_0415_),
    .Y(_1851_),
    .A1(_1801_),
    .A2(_1850_));
 sg13g2_nor2b_2 _5609_ (.A(_1849_),
    .B_N(_1851_),
    .Y(_1852_));
 sg13g2_a21oi_1 _5610_ (.A1(_1801_),
    .A2(_1850_),
    .Y(_1853_),
    .B1(_1852_));
 sg13g2_nor2_1 _5611_ (.A(_1764_),
    .B(_1853_),
    .Y(_1854_));
 sg13g2_nand2_1 _5612_ (.Y(_1855_),
    .A(_1764_),
    .B(_1853_));
 sg13g2_nand2b_1 _5613_ (.Y(_1856_),
    .B(_1855_),
    .A_N(_1854_));
 sg13g2_o21ai_1 _5614_ (.B1(_1847_),
    .Y(_1857_),
    .A1(_1842_),
    .A2(_1848_));
 sg13g2_xnor2_1 _5615_ (.Y(\main.demo._d___pip_58_1_1___stage___block_3_cy[8] ),
    .A(_1856_),
    .B(_1857_));
 sg13g2_nand2_1 _5616_ (.Y(_1858_),
    .A(_1778_),
    .B(_1852_));
 sg13g2_nor2_1 _5617_ (.A(_1778_),
    .B(_1852_),
    .Y(_1859_));
 sg13g2_xor2_1 _5618_ (.B(_1852_),
    .A(_1778_),
    .X(_1860_));
 sg13g2_a21oi_1 _5619_ (.A1(_1855_),
    .A2(_1857_),
    .Y(_1861_),
    .B1(_1854_));
 sg13g2_xnor2_1 _5620_ (.Y(\main.demo._d___pip_58_1_1___stage___block_3_cy[9] ),
    .A(_1860_),
    .B(_1861_));
 sg13g2_a21oi_1 _5621_ (.A1(_0415_),
    .A2(_1850_),
    .Y(_1862_),
    .B1(_1801_));
 sg13g2_a21oi_1 _5622_ (.A1(_1858_),
    .A2(_1861_),
    .Y(_1863_),
    .B1(_1859_));
 sg13g2_xor2_1 _5623_ (.B(_1863_),
    .A(_1862_),
    .X(\main.demo._d___pip_58_1_1___stage___block_3_cy[10] ));
 sg13g2_xnor2_1 _5624_ (.Y(_1864_),
    .A(net407),
    .B(\main.demo._t___stage___block_3_x[1] ));
 sg13g2_xnor2_1 _5625_ (.Y(_1865_),
    .A(\main.demo._t___stage___block_3_y[2] ),
    .B(\main.demo._t___stage___block_3_x[2] ));
 sg13g2_nor2b_1 _5626_ (.A(\main.demo._t___stage___block_3_y[2] ),
    .B_N(\main.demo._q_frame[0] ),
    .Y(_1866_));
 sg13g2_o21ai_1 _5627_ (.B1(_1865_),
    .Y(_1867_),
    .A1(\main.demo._q_frame[1] ),
    .A2(_1866_));
 sg13g2_a22oi_1 _5628_ (.Y(_1868_),
    .B1(_1866_),
    .B2(\main.demo._q_frame[1] ),
    .A2(_2641_),
    .A1(\main.demo._q_frame[2] ));
 sg13g2_a22oi_1 _5629_ (.Y(_1869_),
    .B1(_1867_),
    .B2(_1868_),
    .A2(net407),
    .A1(_2634_));
 sg13g2_a21oi_1 _5630_ (.A1(net436),
    .A2(_1864_),
    .Y(_1870_),
    .B1(_1869_));
 sg13g2_nand2b_1 _5631_ (.Y(_1871_),
    .B(\main.demo._t___stage___block_3_y[0] ),
    .A_N(net435));
 sg13g2_o21ai_1 _5632_ (.B1(_1871_),
    .Y(_1872_),
    .A1(net436),
    .A2(_1864_));
 sg13g2_a22oi_1 _5633_ (.Y(_1873_),
    .B1(_1017_),
    .B2(\main.demo._q_frame[5] ),
    .A2(_2640_),
    .A1(net435));
 sg13g2_o21ai_1 _5634_ (.B1(_1873_),
    .Y(_1874_),
    .A1(_1870_),
    .A2(_1872_));
 sg13g2_nand4_1 _5635_ (.B(\main.demo._q_frame[6] ),
    .C(\main.demo._q_go ),
    .A(net500),
    .Y(_1875_),
    .D(net634));
 sg13g2_o21ai_1 _5636_ (.B1(_1874_),
    .Y(_1876_),
    .A1(\main.demo._q_frame[5] ),
    .A2(net381));
 sg13g2_or2_2 _5637_ (.X(_1877_),
    .B(_1876_),
    .A(_1875_));
 sg13g2_nor2b_1 _5638_ (.A(\main.demo._t___stage___block_3_y[2] ),
    .B_N(\main.demo._d___pip_58_1_4___stage___block_3_cx[1] ),
    .Y(_1878_));
 sg13g2_o21ai_1 _5639_ (.B1(_1878_),
    .Y(_1879_),
    .A1(_2644_),
    .A2(\main.demo._d___pip_58_1_4___stage___block_3_cx[2] ));
 sg13g2_a22oi_1 _5640_ (.Y(_1880_),
    .B1(\main.demo._d___pip_58_1_4___stage___block_3_cx[2] ),
    .B2(_1865_),
    .A2(\main.demo._d___pip_58_1_4___stage___block_3_cx[3] ),
    .A1(_2641_));
 sg13g2_a22oi_1 _5641_ (.Y(_1881_),
    .B1(_1879_),
    .B2(_1880_),
    .A2(_2672_),
    .A1(net407));
 sg13g2_o21ai_1 _5642_ (.B1(_1881_),
    .Y(_1882_),
    .A1(\main.demo._d___pip_58_1_4___stage___block_3_cx[4] ),
    .A2(_1864_));
 sg13g2_a22oi_1 _5643_ (.Y(_1883_),
    .B1(\main.demo._d___pip_58_1_4___stage___block_3_cx[4] ),
    .B2(_1864_),
    .A2(\main.demo._d___pip_58_1_4___stage___block_3_cx[5] ),
    .A1(_2640_));
 sg13g2_nand2_1 _5644_ (.Y(_1884_),
    .A(_1882_),
    .B(_1883_));
 sg13g2_a22oi_1 _5645_ (.Y(_1885_),
    .B1(net383),
    .B2(_2670_),
    .A2(_2671_),
    .A1(\main.demo._t___stage___block_3_y[0] ));
 sg13g2_a221oi_1 _5646_ (.B2(_1885_),
    .C1(\main.demo._d___pip_58_1_4___stage___block_3_cx[9] ),
    .B1(_1884_),
    .A1(\main.demo._d___pip_58_1_4___stage___block_3_cx[6] ),
    .Y(_1886_),
    .A2(net381));
 sg13g2_nand2_1 _5647_ (.Y(_1887_),
    .A(\main.demo._d___pip_58_1_4___block_87_atten_l[1] ),
    .B(\main.demo._d___pip_58_1_4___block_68_frag[3] ));
 sg13g2_nand2_1 _5648_ (.Y(_1888_),
    .A(\main.demo._d___pip_58_1_4___block_87_atten_l[0] ),
    .B(\main.demo._d___pip_58_1_4___block_68_frag[4] ));
 sg13g2_nor2_1 _5649_ (.A(_1887_),
    .B(_1888_),
    .Y(_1889_));
 sg13g2_and2_1 _5650_ (.A(\main.demo._d___pip_58_1_4___block_87_atten_l[1] ),
    .B(\main.demo._d___pip_58_1_4___block_68_frag[1] ),
    .X(_1890_));
 sg13g2_nand2_1 _5651_ (.Y(_1891_),
    .A(net423),
    .B(\main.demo._d___pip_58_1_4___block_68_frag[1] ));
 sg13g2_nand2_1 _5652_ (.Y(_1892_),
    .A(net424),
    .B(\main.demo._d___pip_58_1_4___block_68_frag[0] ));
 sg13g2_nor3_1 _5653_ (.A(_2669_),
    .B(_1891_),
    .C(_1892_),
    .Y(_1893_));
 sg13g2_nand2_2 _5654_ (.Y(_1894_),
    .A(net424),
    .B(\main.demo._d___pip_58_1_4___block_68_frag[2] ));
 sg13g2_nor2_1 _5655_ (.A(_1887_),
    .B(_1894_),
    .Y(_1895_));
 sg13g2_nor2_1 _5656_ (.A(_1893_),
    .B(_1895_),
    .Y(_1896_));
 sg13g2_o21ai_1 _5657_ (.B1(_1896_),
    .Y(_1897_),
    .A1(_1891_),
    .A2(_1894_));
 sg13g2_xor2_1 _5658_ (.B(_1888_),
    .A(_1887_),
    .X(_1898_));
 sg13g2_and2_1 _5659_ (.A(_1897_),
    .B(_1898_),
    .X(_1899_));
 sg13g2_nor2_1 _5660_ (.A(_1889_),
    .B(_1899_),
    .Y(_1900_));
 sg13g2_nand2_1 _5661_ (.Y(_1901_),
    .A(net423),
    .B(\main.demo._d___pip_58_1_4___block_68_frag[5] ));
 sg13g2_nor2_1 _5662_ (.A(_1888_),
    .B(_1901_),
    .Y(_1902_));
 sg13g2_a22oi_1 _5663_ (.Y(_1903_),
    .B1(\main.demo._d___pip_58_1_4___block_68_frag[4] ),
    .B2(net423),
    .A2(\main.demo._d___pip_58_1_4___block_68_frag[5] ),
    .A1(net424));
 sg13g2_nor2_1 _5664_ (.A(_1902_),
    .B(_1903_),
    .Y(_1904_));
 sg13g2_xnor2_1 _5665_ (.Y(_1905_),
    .A(_1900_),
    .B(_1904_));
 sg13g2_and2_1 _5666_ (.A(\main.demo._d___pip_58_1_4___block_68_frag[4] ),
    .B(\main.demo._d___pip_58_1_4___block_87_atten_h[0] ),
    .X(_1906_));
 sg13g2_nand2_1 _5667_ (.Y(_1907_),
    .A(\main.demo._d___pip_58_1_4___block_68_frag[2] ),
    .B(\main.demo._d___pip_58_1_4___block_87_atten_h[1] ));
 sg13g2_nand2_1 _5668_ (.Y(_1908_),
    .A(\main.demo._d___pip_58_1_4___block_68_frag[3] ),
    .B(\main.demo._d___pip_58_1_4___block_87_atten_h[2] ));
 sg13g2_or2_1 _5669_ (.X(_1909_),
    .B(_1908_),
    .A(_1907_));
 sg13g2_inv_1 _5670_ (.Y(_1910_),
    .A(_1909_));
 sg13g2_a22oi_1 _5671_ (.Y(_1911_),
    .B1(\main.demo._d___pip_58_1_4___block_87_atten_h[1] ),
    .B2(\main.demo._d___pip_58_1_4___block_68_frag[3] ),
    .A2(\main.demo._d___pip_58_1_4___block_87_atten_h[2] ),
    .A1(\main.demo._d___pip_58_1_4___block_68_frag[2] ));
 sg13g2_nor2_1 _5672_ (.A(_1910_),
    .B(_1911_),
    .Y(_1912_));
 sg13g2_xor2_1 _5673_ (.B(_1912_),
    .A(_1906_),
    .X(_1913_));
 sg13g2_and2_1 _5674_ (.A(\main.demo._d___pip_58_1_4___block_68_frag[1] ),
    .B(\main.demo._d___pip_58_1_4___block_87_atten_h[1] ),
    .X(_1914_));
 sg13g2_nand2_1 _5675_ (.Y(_1915_),
    .A(\main.demo._d___pip_58_1_4___block_68_frag[1] ),
    .B(\main.demo._d___pip_58_1_4___block_87_atten_h[2] ));
 sg13g2_nand2_1 _5676_ (.Y(_1916_),
    .A(\main.demo._d___pip_58_1_4___block_68_frag[3] ),
    .B(\main.demo._d___pip_58_1_4___block_87_atten_h[0] ));
 sg13g2_xor2_1 _5677_ (.B(_1915_),
    .A(_1907_),
    .X(_1917_));
 sg13g2_nand2b_1 _5678_ (.Y(_1918_),
    .B(_1917_),
    .A_N(_1916_));
 sg13g2_o21ai_1 _5679_ (.B1(_1918_),
    .Y(_1919_),
    .A1(_1907_),
    .A2(_1915_));
 sg13g2_nand2_1 _5680_ (.Y(_1920_),
    .A(_1913_),
    .B(_1919_));
 sg13g2_and2_1 _5681_ (.A(\main.demo._d___pip_58_1_4___block_68_frag[0] ),
    .B(_1914_),
    .X(_1921_));
 sg13g2_and2_1 _5682_ (.A(\main.demo._d___pip_58_1_4___block_68_frag[2] ),
    .B(\main.demo._d___pip_58_1_4___block_87_atten_h[0] ),
    .X(_1922_));
 sg13g2_a21oi_1 _5683_ (.A1(\main.demo._d___pip_58_1_4___block_68_frag[0] ),
    .A2(\main.demo._d___pip_58_1_4___block_87_atten_h[2] ),
    .Y(_1923_),
    .B1(_1914_));
 sg13g2_a21oi_1 _5684_ (.A1(\main.demo._d___pip_58_1_4___block_87_atten_h[2] ),
    .A2(_1921_),
    .Y(_1924_),
    .B1(_1923_));
 sg13g2_a22oi_1 _5685_ (.Y(_1925_),
    .B1(_1922_),
    .B2(_1924_),
    .A2(_1921_),
    .A1(\main.demo._d___pip_58_1_4___block_87_atten_h[2] ));
 sg13g2_xnor2_1 _5686_ (.Y(_1926_),
    .A(_1916_),
    .B(_1917_));
 sg13g2_nor2b_1 _5687_ (.A(_1925_),
    .B_N(_1926_),
    .Y(_1927_));
 sg13g2_xor2_1 _5688_ (.B(_1924_),
    .A(_1922_),
    .X(_1928_));
 sg13g2_nand2_1 _5689_ (.Y(_1929_),
    .A(\main.demo._d___pip_58_1_4___block_87_atten_h[0] ),
    .B(_1921_));
 sg13g2_nand3_1 _5690_ (.B(_1921_),
    .C(_1928_),
    .A(\main.demo._d___pip_58_1_4___block_87_atten_h[0] ),
    .Y(_1930_));
 sg13g2_xnor2_1 _5691_ (.Y(_1931_),
    .A(_1925_),
    .B(_1926_));
 sg13g2_nor2b_1 _5692_ (.A(_1930_),
    .B_N(_1931_),
    .Y(_1932_));
 sg13g2_xor2_1 _5693_ (.B(_1919_),
    .A(_1913_),
    .X(_1933_));
 sg13g2_o21ai_1 _5694_ (.B1(_1933_),
    .Y(_1934_),
    .A1(_1927_),
    .A2(_1932_));
 sg13g2_a21oi_1 _5695_ (.A1(_1906_),
    .A2(_1912_),
    .Y(_1935_),
    .B1(_1910_));
 sg13g2_nand2_1 _5696_ (.Y(_1936_),
    .A(\main.demo._d___pip_58_1_4___block_68_frag[5] ),
    .B(\main.demo._d___pip_58_1_4___block_87_atten_h[0] ));
 sg13g2_nand2_1 _5697_ (.Y(_1937_),
    .A(\main.demo._d___pip_58_1_4___block_68_frag[4] ),
    .B(\main.demo._d___pip_58_1_4___block_87_atten_h[2] ));
 sg13g2_nand2_1 _5698_ (.Y(_1938_),
    .A(\main.demo._d___pip_58_1_4___block_68_frag[4] ),
    .B(\main.demo._d___pip_58_1_4___block_87_atten_h[1] ));
 sg13g2_xor2_1 _5699_ (.B(_1938_),
    .A(_1908_),
    .X(_1939_));
 sg13g2_nand2b_1 _5700_ (.Y(_1940_),
    .B(_1939_),
    .A_N(_1936_));
 sg13g2_xnor2_1 _5701_ (.Y(_1941_),
    .A(_1936_),
    .B(_1939_));
 sg13g2_nor2b_1 _5702_ (.A(_1935_),
    .B_N(_1941_),
    .Y(_1942_));
 sg13g2_xor2_1 _5703_ (.B(_1941_),
    .A(_1935_),
    .X(_1943_));
 sg13g2_nand3_1 _5704_ (.B(_1934_),
    .C(_1943_),
    .A(_1920_),
    .Y(_1944_));
 sg13g2_a21oi_1 _5705_ (.A1(_1920_),
    .A2(_1934_),
    .Y(_1945_),
    .B1(_1943_));
 sg13g2_nor2_1 _5706_ (.A(net362),
    .B(_1945_),
    .Y(_1946_));
 sg13g2_a22oi_1 _5707_ (.Y(_1947_),
    .B1(_1944_),
    .B2(_1946_),
    .A2(_1905_),
    .A1(net362));
 sg13g2_and2_1 _5708_ (.A(net384),
    .B(_1947_),
    .X(_1948_));
 sg13g2_nor2_1 _5709_ (.A(net384),
    .B(_1947_),
    .Y(_1949_));
 sg13g2_xor2_1 _5710_ (.B(_1898_),
    .A(_1897_),
    .X(_1950_));
 sg13g2_or3_1 _5711_ (.A(_1927_),
    .B(_1932_),
    .C(_1933_),
    .X(_1951_));
 sg13g2_nor2b_1 _5712_ (.A(net362),
    .B_N(_1934_),
    .Y(_1952_));
 sg13g2_a22oi_1 _5713_ (.Y(_1953_),
    .B1(_1951_),
    .B2(_1952_),
    .A2(_1950_),
    .A1(_1886_));
 sg13g2_a21oi_1 _5714_ (.A1(_1892_),
    .A2(_1894_),
    .Y(_1954_),
    .B1(_1891_));
 sg13g2_a22oi_1 _5715_ (.Y(_1955_),
    .B1(\main.demo._d___pip_58_1_4___block_68_frag[2] ),
    .B2(net423),
    .A2(\main.demo._d___pip_58_1_4___block_68_frag[3] ),
    .A1(net424));
 sg13g2_nor2_1 _5716_ (.A(_1895_),
    .B(_1955_),
    .Y(_1956_));
 sg13g2_xor2_1 _5717_ (.B(_1956_),
    .A(_1954_),
    .X(_1957_));
 sg13g2_nand2_1 _5718_ (.Y(_1958_),
    .A(_1886_),
    .B(_1957_));
 sg13g2_xor2_1 _5719_ (.B(_1931_),
    .A(_1930_),
    .X(_1959_));
 sg13g2_o21ai_1 _5720_ (.B1(_1958_),
    .Y(_1960_),
    .A1(net362),
    .A2(_1959_));
 sg13g2_xnor2_1 _5721_ (.Y(_1961_),
    .A(_0004_),
    .B(_1953_));
 sg13g2_o21ai_1 _5722_ (.B1(_1961_),
    .Y(_1962_),
    .A1(_1864_),
    .A2(_1960_));
 sg13g2_nor3_1 _5723_ (.A(_1948_),
    .B(_1949_),
    .C(_1962_),
    .Y(_1963_));
 sg13g2_nand2_1 _5724_ (.Y(_1964_),
    .A(_1864_),
    .B(_1960_));
 sg13g2_nand3_1 _5725_ (.B(_1892_),
    .C(_1894_),
    .A(_1890_),
    .Y(_1965_));
 sg13g2_a21oi_1 _5726_ (.A1(_1890_),
    .A2(_1892_),
    .Y(_1966_),
    .B1(_1894_));
 sg13g2_nand3b_1 _5727_ (.B(_1886_),
    .C(_1965_),
    .Y(_1967_),
    .A_N(_1966_));
 sg13g2_xnor2_1 _5728_ (.Y(_1968_),
    .A(_1928_),
    .B(_1929_));
 sg13g2_o21ai_1 _5729_ (.B1(_1967_),
    .Y(_1969_),
    .A1(net362),
    .A2(_1968_));
 sg13g2_o21ai_1 _5730_ (.B1(_1964_),
    .Y(_1970_),
    .A1(_2645_),
    .A2(_1969_));
 sg13g2_a21oi_1 _5731_ (.A1(_2645_),
    .A2(_1969_),
    .Y(_1971_),
    .B1(_1970_));
 sg13g2_nand3_1 _5732_ (.B(_1964_),
    .C(_1969_),
    .A(\main.demo._t___stage___block_3_x[1] ),
    .Y(_1972_));
 sg13g2_nand2_1 _5733_ (.Y(_1973_),
    .A(_1963_),
    .B(_1972_));
 sg13g2_nor3_1 _5734_ (.A(\main.demo._t___stage___block_3_x[0] ),
    .B(_1948_),
    .C(_1953_),
    .Y(_1974_));
 sg13g2_nor2_1 _5735_ (.A(_1949_),
    .B(_1974_),
    .Y(_1975_));
 sg13g2_a22oi_1 _5736_ (.Y(_1976_),
    .B1(_1973_),
    .B2(_1975_),
    .A2(_1971_),
    .A1(_1963_));
 sg13g2_nor2b_1 _5737_ (.A(_1903_),
    .B_N(_1899_),
    .Y(_1977_));
 sg13g2_nor3_1 _5738_ (.A(_1889_),
    .B(_1902_),
    .C(_1977_),
    .Y(_1978_));
 sg13g2_o21ai_1 _5739_ (.B1(net362),
    .Y(_1979_),
    .A1(_1901_),
    .A2(_1978_));
 sg13g2_a21oi_1 _5740_ (.A1(_1901_),
    .A2(_1978_),
    .Y(_1980_),
    .B1(_1979_));
 sg13g2_o21ai_1 _5741_ (.B1(_1940_),
    .Y(_1981_),
    .A1(_1908_),
    .A2(_1938_));
 sg13g2_nand2_1 _5742_ (.Y(_1982_),
    .A(\main.demo._d___pip_58_1_4___block_68_frag[5] ),
    .B(\main.demo._d___pip_58_1_4___block_87_atten_h[1] ));
 sg13g2_xor2_1 _5743_ (.B(_1982_),
    .A(_1937_),
    .X(_1983_));
 sg13g2_xor2_1 _5744_ (.B(_1983_),
    .A(_1981_),
    .X(_1984_));
 sg13g2_nor3_1 _5745_ (.A(_1942_),
    .B(_1945_),
    .C(_1984_),
    .Y(_1985_));
 sg13g2_o21ai_1 _5746_ (.B1(_1984_),
    .Y(_1986_),
    .A1(_1942_),
    .A2(_1945_));
 sg13g2_inv_1 _5747_ (.Y(_1987_),
    .A(_1986_));
 sg13g2_nor2_1 _5748_ (.A(net362),
    .B(_1985_),
    .Y(_1988_));
 sg13g2_a21oi_1 _5749_ (.A1(_1986_),
    .A2(_1988_),
    .Y(_1989_),
    .B1(_1980_));
 sg13g2_nor2b_1 _5750_ (.A(_1976_),
    .B_N(_1989_),
    .Y(_1990_));
 sg13g2_nand2b_1 _5751_ (.Y(_1991_),
    .B(_1976_),
    .A_N(_1989_));
 sg13g2_nand3_1 _5752_ (.B(\main.demo._d___pip_58_1_4___block_87_atten_h[2] ),
    .C(_1938_),
    .A(\main.demo._d___pip_58_1_4___block_68_frag[5] ),
    .Y(_1992_));
 sg13g2_a21oi_1 _5753_ (.A1(_1981_),
    .A2(_1983_),
    .Y(_1993_),
    .B1(_1987_));
 sg13g2_xor2_1 _5754_ (.B(_1993_),
    .A(_1992_),
    .X(_1994_));
 sg13g2_o21ai_1 _5755_ (.B1(_1979_),
    .Y(_1995_),
    .A1(net362),
    .A2(_1994_));
 sg13g2_nor2b_1 _5756_ (.A(_1991_),
    .B_N(_1995_),
    .Y(_1996_));
 sg13g2_o21ai_1 _5757_ (.B1(_1877_),
    .Y(\main.demo._d_prev_b[0] ),
    .A1(_1990_),
    .A2(_1996_));
 sg13g2_nor2_1 _5758_ (.A(\main.demo._w_vga_vga_x[5] ),
    .B(\main.demo._w_vga_vga_y[5] ),
    .Y(_1997_));
 sg13g2_nor2_1 _5759_ (.A(_2633_),
    .B(\main.demo._w_vga_vga_y[6] ),
    .Y(_1998_));
 sg13g2_a21oi_1 _5760_ (.A1(\main.demo._w_vga_vga_y[5] ),
    .A2(_1998_),
    .Y(_1999_),
    .B1(_1997_));
 sg13g2_nor2_1 _5761_ (.A(net414),
    .B(_1999_),
    .Y(_2000_));
 sg13g2_nor2_1 _5762_ (.A(net412),
    .B(net413),
    .Y(_2001_));
 sg13g2_a21oi_1 _5763_ (.A1(_2000_),
    .A2(_2001_),
    .Y(_2002_),
    .B1(_2630_));
 sg13g2_and2_1 _5764_ (.A(\main.demo._w_vga_vga_y[6] ),
    .B(\main.demo._w_vga_vga_y[5] ),
    .X(_2003_));
 sg13g2_nand2_1 _5765_ (.Y(_2004_),
    .A(\main.demo._w_vga_vga_y[6] ),
    .B(\main.demo._w_vga_vga_y[5] ));
 sg13g2_nand2_1 _5766_ (.Y(_2005_),
    .A(\main.demo._w_vga_vga_x[5] ),
    .B(_2004_));
 sg13g2_inv_1 _5767_ (.Y(_2006_),
    .A(_2005_));
 sg13g2_nor2_1 _5768_ (.A(\main.demo._w_vga_vga_y[6] ),
    .B(\main.demo._w_vga_vga_y[5] ),
    .Y(_2007_));
 sg13g2_o21ai_1 _5769_ (.B1(\main.demo._w_vga_vga_x[5] ),
    .Y(_2008_),
    .A1(\main.demo._w_vga_vga_y[6] ),
    .A2(\main.demo._w_vga_vga_y[5] ));
 sg13g2_nor2_2 _5770_ (.A(_2003_),
    .B(_2008_),
    .Y(_2009_));
 sg13g2_nand2_1 _5771_ (.Y(_2010_),
    .A(net412),
    .B(net413));
 sg13g2_a22oi_1 _5772_ (.Y(_2011_),
    .B1(_2009_),
    .B2(_2010_),
    .A2(_2006_),
    .A1(\main.demo._w_vga_vga_x[6] ));
 sg13g2_or2_1 _5773_ (.X(_2012_),
    .B(_2011_),
    .A(_2001_));
 sg13g2_nor2_1 _5774_ (.A(_0056_),
    .B(_1998_),
    .Y(_2013_));
 sg13g2_and2_1 _5775_ (.A(_2001_),
    .B(_2004_),
    .X(_2014_));
 sg13g2_a221oi_1 _5776_ (.B2(_2014_),
    .C1(\main.demo._w_vga_vga_x[9] ),
    .B1(_2013_),
    .A1(net412),
    .Y(_2015_),
    .A2(_2000_));
 sg13g2_a21oi_1 _5777_ (.A1(_2012_),
    .A2(_2015_),
    .Y(_2016_),
    .B1(_2002_));
 sg13g2_nand4_1 _5778_ (.B(_0054_),
    .C(_2631_),
    .A(\main.demo._w_vga_vga_x[9] ),
    .Y(_2017_),
    .D(_2632_));
 sg13g2_or2_1 _5779_ (.X(_2018_),
    .B(_1998_),
    .A(_1997_));
 sg13g2_nand2b_1 _5780_ (.Y(_2019_),
    .B(_2018_),
    .A_N(_2017_));
 sg13g2_nand2_1 _5781_ (.Y(_2020_),
    .A(\main.demo._w_vga_vga_x[6] ),
    .B(_2009_));
 sg13g2_a21oi_1 _5782_ (.A1(\main.demo._w_vga_vga_y[6] ),
    .A2(_0063_),
    .Y(_2021_),
    .B1(_1998_));
 sg13g2_o21ai_1 _5783_ (.B1(_2020_),
    .Y(_2022_),
    .A1(net414),
    .A2(_2021_));
 sg13g2_nor2_1 _5784_ (.A(net413),
    .B(_2632_),
    .Y(_2023_));
 sg13g2_nand2_1 _5785_ (.Y(_2024_),
    .A(_2633_),
    .B(_2023_));
 sg13g2_nor3_1 _5786_ (.A(_2003_),
    .B(_2007_),
    .C(_2024_),
    .Y(_2025_));
 sg13g2_a21o_1 _5787_ (.A2(_2022_),
    .A1(net413),
    .B1(_2025_),
    .X(_2026_));
 sg13g2_a21oi_1 _5788_ (.A1(\main.demo._w_vga_vga_x[5] ),
    .A2(\main.demo._w_vga_vga_y[5] ),
    .Y(_2027_),
    .B1(_2018_));
 sg13g2_a21oi_1 _5789_ (.A1(_0057_),
    .A2(_2636_),
    .Y(_2028_),
    .B1(net413));
 sg13g2_a221oi_1 _5790_ (.B2(_2005_),
    .C1(net414),
    .B1(_2028_),
    .A1(net413),
    .Y(_2029_),
    .A2(_2027_));
 sg13g2_nand3b_1 _5791_ (.B(net412),
    .C(_2020_),
    .Y(_2030_),
    .A_N(_2029_));
 sg13g2_o21ai_1 _5792_ (.B1(_2030_),
    .Y(_2031_),
    .A1(net412),
    .A2(_2026_));
 sg13g2_o21ai_1 _5793_ (.B1(_2019_),
    .Y(_2032_),
    .A1(\main.demo._w_vga_vga_x[9] ),
    .A2(_2031_));
 sg13g2_o21ai_1 _5794_ (.B1(_2633_),
    .Y(_2033_),
    .A1(_2003_),
    .A2(_2007_));
 sg13g2_nand3_1 _5795_ (.B(_2005_),
    .C(_2033_),
    .A(net414),
    .Y(_2034_));
 sg13g2_or2_1 _5796_ (.X(_2035_),
    .B(_2008_),
    .A(_2631_));
 sg13g2_mux2_1 _5797_ (.A0(net413),
    .A1(_2035_),
    .S(_2034_),
    .X(_2036_));
 sg13g2_nor2_2 _5798_ (.A(_1997_),
    .B(_2009_),
    .Y(_2037_));
 sg13g2_o21ai_1 _5799_ (.B1(\main.demo._w_vga_vga_x[7] ),
    .Y(_2038_),
    .A1(_2632_),
    .A2(_2008_));
 sg13g2_inv_1 _5800_ (.Y(_2039_),
    .A(_2038_));
 sg13g2_o21ai_1 _5801_ (.B1(_2039_),
    .Y(_2040_),
    .A1(net414),
    .A2(_2037_));
 sg13g2_o21ai_1 _5802_ (.B1(_2008_),
    .Y(_2041_),
    .A1(_2023_),
    .A2(_2028_));
 sg13g2_nand3_1 _5803_ (.B(_2040_),
    .C(_2041_),
    .A(net412),
    .Y(_2042_));
 sg13g2_o21ai_1 _5804_ (.B1(_2042_),
    .Y(_2043_),
    .A1(net412),
    .A2(_2036_));
 sg13g2_nand2_1 _5805_ (.Y(_2044_),
    .A(_2630_),
    .B(_2043_));
 sg13g2_o21ai_1 _5806_ (.B1(_2044_),
    .Y(_2045_),
    .A1(_2017_),
    .A2(_2037_));
 sg13g2_nor2_1 _5807_ (.A(net414),
    .B(\main.demo._w_vga_vga_x[5] ),
    .Y(_2046_));
 sg13g2_a221oi_1 _5808_ (.B2(_2046_),
    .C1(_2000_),
    .B1(\main.demo._w_vga_vga_y[6] ),
    .A1(_2631_),
    .Y(_2047_),
    .A2(_2632_));
 sg13g2_a22oi_1 _5809_ (.Y(_2048_),
    .B1(_2047_),
    .B2(_2020_),
    .A2(_2037_),
    .A1(_2631_));
 sg13g2_nor3_1 _5810_ (.A(net414),
    .B(\main.demo._w_vga_vga_x[5] ),
    .C(_2004_),
    .Y(_2049_));
 sg13g2_nor3_1 _5811_ (.A(_2009_),
    .B(_2038_),
    .C(_2049_),
    .Y(_2050_));
 sg13g2_nor3_1 _5812_ (.A(_0056_),
    .B(\main.demo._w_vga_vga_x[5] ),
    .C(_2007_),
    .Y(_2051_));
 sg13g2_nor2_1 _5813_ (.A(net413),
    .B(_2051_),
    .Y(_2052_));
 sg13g2_nor3_1 _5814_ (.A(\main.demo._w_vga_vga_x[8] ),
    .B(_2050_),
    .C(_2052_),
    .Y(_2053_));
 sg13g2_a21oi_1 _5815_ (.A1(net412),
    .A2(_2048_),
    .Y(_2054_),
    .B1(_2053_));
 sg13g2_a21oi_1 _5816_ (.A1(_2630_),
    .A2(_2054_),
    .Y(_2055_),
    .B1(_2002_));
 sg13g2_nor2_1 _5817_ (.A(_2045_),
    .B(_2055_),
    .Y(_2056_));
 sg13g2_or2_2 _5818_ (.X(_2057_),
    .B(_2045_),
    .A(_2016_));
 sg13g2_xnor2_1 _5819_ (.Y(_2058_),
    .A(\main.demo._w_vga_vga_x[4] ),
    .B(_2057_));
 sg13g2_xnor2_1 _5820_ (.Y(_2059_),
    .A(\main.demo._w_vga_vga_x[3] ),
    .B(_2057_));
 sg13g2_xnor2_1 _5821_ (.Y(_2060_),
    .A(_2644_),
    .B(_2057_));
 sg13g2_xor2_1 _5822_ (.B(_2060_),
    .A(_0003_),
    .X(_2061_));
 sg13g2_xnor2_1 _5823_ (.Y(_2062_),
    .A(\main.demo._t___stage___block_3_x[1] ),
    .B(_2057_));
 sg13g2_nor2_1 _5824_ (.A(net407),
    .B(_2062_),
    .Y(_2063_));
 sg13g2_xnor2_1 _5825_ (.Y(_2064_),
    .A(_0004_),
    .B(_2057_));
 sg13g2_nor3_1 _5826_ (.A(_2640_),
    .B(_2063_),
    .C(_2064_),
    .Y(_2065_));
 sg13g2_a21oi_1 _5827_ (.A1(net407),
    .A2(_2062_),
    .Y(_2066_),
    .B1(_2065_));
 sg13g2_a22oi_1 _5828_ (.Y(_2067_),
    .B1(_2061_),
    .B2(_2066_),
    .A2(_2060_),
    .A1(_2643_));
 sg13g2_a21oi_1 _5829_ (.A1(\main.demo._w_vga_vga_y[3] ),
    .A2(_2059_),
    .Y(_2068_),
    .B1(_2067_));
 sg13g2_nor2_1 _5830_ (.A(\main.demo._w_vga_vga_y[4] ),
    .B(_2058_),
    .Y(_2069_));
 sg13g2_nor2_1 _5831_ (.A(\main.demo._w_vga_vga_y[3] ),
    .B(_2059_),
    .Y(_2070_));
 sg13g2_nor3_1 _5832_ (.A(_2068_),
    .B(_2069_),
    .C(_2070_),
    .Y(_2071_));
 sg13g2_a21oi_1 _5833_ (.A1(\main.demo._w_vga_vga_y[4] ),
    .A2(_2058_),
    .Y(_2072_),
    .B1(_2071_));
 sg13g2_xor2_1 _5834_ (.B(_2072_),
    .A(_2056_),
    .X(_2073_));
 sg13g2_a21oi_1 _5835_ (.A1(_2016_),
    .A2(_2032_),
    .Y(_2074_),
    .B1(_2073_));
 sg13g2_nor3_1 _5836_ (.A(_2032_),
    .B(_2055_),
    .C(_2057_),
    .Y(_2075_));
 sg13g2_nor2b_1 _5837_ (.A(net415),
    .B_N(\main.demo._q_th[1] ),
    .Y(_2076_));
 sg13g2_o21ai_1 _5838_ (.B1(_2076_),
    .Y(_2077_),
    .A1(\main.demo._q_th[2] ),
    .A2(_2642_));
 sg13g2_nor2_1 _5839_ (.A(_2612_),
    .B(\main.demo._w_vga_vga_x[3] ),
    .Y(_2078_));
 sg13g2_a22oi_1 _5840_ (.Y(_2079_),
    .B1(_2644_),
    .B2(\main.demo._q_th[3] ),
    .A2(_2642_),
    .A1(\main.demo._q_th[2] ));
 sg13g2_a22oi_1 _5841_ (.Y(_2080_),
    .B1(_2077_),
    .B2(_2079_),
    .A2(\main.demo._t___stage___block_3_x[2] ),
    .A1(_2613_));
 sg13g2_a22oi_1 _5842_ (.Y(_2081_),
    .B1(\main.demo._w_vga_vga_x[3] ),
    .B2(_2612_),
    .A2(\main.demo._w_vga_vga_x[4] ),
    .A1(_2611_));
 sg13g2_o21ai_1 _5843_ (.B1(_2081_),
    .Y(_2082_),
    .A1(_2078_),
    .A2(_2080_));
 sg13g2_o21ai_1 _5844_ (.B1(_2082_),
    .Y(_2083_),
    .A1(_2611_),
    .A2(\main.demo._w_vga_vga_x[4] ));
 sg13g2_nor4_1 _5845_ (.A(\main.demo._q_th[8] ),
    .B(net312),
    .C(\main.demo._q_th[6] ),
    .D(_2083_),
    .Y(_2084_));
 sg13g2_and2_2 _5846_ (.A(\main.demo._q_go ),
    .B(_0969_),
    .X(_2085_));
 sg13g2_nand2_1 _5847_ (.Y(_2086_),
    .A(\main.demo._q_go ),
    .B(_0969_));
 sg13g2_nor3_1 _5848_ (.A(\main.demo._w_vga_vga_y[10] ),
    .B(\main.demo._w_vga_vga_y[8] ),
    .C(_2086_),
    .Y(_2087_));
 sg13g2_o21ai_1 _5849_ (.B1(_2087_),
    .Y(_2088_),
    .A1(_2635_),
    .A2(\main.demo._w_vga_vga_y[7] ));
 sg13g2_or4_1 _5850_ (.A(_2074_),
    .B(_2075_),
    .C(_2084_),
    .D(_2088_),
    .X(_2089_));
 sg13g2_nand4_1 _5851_ (.B(_1991_),
    .C(_1995_),
    .A(_1877_),
    .Y(\main.demo._d_prev_b[1] ),
    .D(_2089_));
 sg13g2_or2_1 _5852_ (.X(_2090_),
    .B(_0231_),
    .A(net301));
 sg13g2_and2_1 _5853_ (.A(net452),
    .B(net309),
    .X(_2091_));
 sg13g2_nor3_1 _5854_ (.A(net301),
    .B(_3024_),
    .C(_2091_),
    .Y(_0070_));
 sg13g2_and2_1 _5855_ (.A(net316),
    .B(_2091_),
    .X(_2092_));
 sg13g2_nor2_1 _5856_ (.A(net316),
    .B(_2091_),
    .Y(_2093_));
 sg13g2_nor3_1 _5857_ (.A(_2090_),
    .B(_2092_),
    .C(_2093_),
    .Y(_0071_));
 sg13g2_and2_1 _5858_ (.A(net504),
    .B(_2092_),
    .X(_2094_));
 sg13g2_nand2_1 _5859_ (.Y(_2095_),
    .A(\main.demo.vga._q_xcount[3] ),
    .B(_2092_));
 sg13g2_nor2_1 _5860_ (.A(net504),
    .B(_2092_),
    .Y(_2096_));
 sg13g2_nor3_1 _5861_ (.A(_2090_),
    .B(_2094_),
    .C(_2096_),
    .Y(_0072_));
 sg13g2_xnor2_1 _5862_ (.Y(_2097_),
    .A(net456),
    .B(_2094_));
 sg13g2_nor2_1 _5863_ (.A(_2090_),
    .B(_2097_),
    .Y(_0073_));
 sg13g2_and3_1 _5864_ (.X(_2098_),
    .A(net468),
    .B(net488),
    .C(_2094_));
 sg13g2_and3_1 _5865_ (.X(_2099_),
    .A(net482),
    .B(net460),
    .C(_2098_));
 sg13g2_a21oi_1 _5866_ (.A1(net460),
    .A2(_2098_),
    .Y(_2100_),
    .B1(net482));
 sg13g2_nor3_1 _5867_ (.A(_2090_),
    .B(_2099_),
    .C(_2100_),
    .Y(_0074_));
 sg13g2_nand3_1 _5868_ (.B(\main.demo.vga._q_ycount[0] ),
    .C(net374),
    .A(net625),
    .Y(_2101_));
 sg13g2_inv_1 _5869_ (.Y(_2102_),
    .A(_2101_));
 sg13g2_and3_1 _5870_ (.X(_2103_),
    .A(\main.demo.vga._q_ycount[3] ),
    .B(\main.demo.vga._q_ycount[2] ),
    .C(_2102_));
 sg13g2_and3_1 _5871_ (.X(_2104_),
    .A(net319),
    .B(net561),
    .C(_2103_));
 sg13g2_and2_1 _5872_ (.A(net458),
    .B(_2104_),
    .X(_2105_));
 sg13g2_nand2_2 _5873_ (.Y(_2106_),
    .A(net374),
    .B(_0239_));
 sg13g2_nand4_1 _5874_ (.B(\main.demo.vga._q_ycount[7] ),
    .C(\main.demo.vga._q_ycount[6] ),
    .A(net615),
    .Y(_2107_),
    .D(_2104_));
 sg13g2_nand3_1 _5875_ (.B(\main.demo.vga._q_ycount[2] ),
    .C(net465),
    .A(net475),
    .Y(_2108_));
 sg13g2_xor2_1 _5876_ (.B(_2107_),
    .A(net485),
    .X(_2109_));
 sg13g2_a21oi_1 _5877_ (.A1(_2106_),
    .A2(net617),
    .Y(_0075_),
    .B1(net400));
 sg13g2_nor2_1 _5878_ (.A(\main.demo._q_speed[6] ),
    .B(_1432_),
    .Y(_2110_));
 sg13g2_o21ai_1 _5879_ (.B1(_2085_),
    .Y(_2111_),
    .A1(net575),
    .A2(_2110_));
 sg13g2_a21oi_1 _5880_ (.A1(net575),
    .A2(_2110_),
    .Y(_0076_),
    .B1(_2111_));
 sg13g2_nor2_1 _5881_ (.A(_1432_),
    .B(net371),
    .Y(_2112_));
 sg13g2_nand2_2 _5882_ (.Y(_2113_),
    .A(_1431_),
    .B(_2085_));
 sg13g2_nand2_1 _5883_ (.Y(_2114_),
    .A(\main.demo._q_speed[7] ),
    .B(\main.demo._q_speed[1] ));
 sg13g2_xnor2_1 _5884_ (.Y(_2115_),
    .A(\main.demo._q_speed[7] ),
    .B(\main.demo._q_speed[1] ));
 sg13g2_nor2_1 _5885_ (.A(\main.demo._q_speed[0] ),
    .B(\main.demo._q_speed[6] ),
    .Y(_2116_));
 sg13g2_xnor2_1 _5886_ (.Y(_2117_),
    .A(_2115_),
    .B(_2116_));
 sg13g2_nor2_1 _5887_ (.A(_1431_),
    .B(net371),
    .Y(_2118_));
 sg13g2_nor3_1 _5888_ (.A(net623),
    .B(_1431_),
    .C(net373),
    .Y(_2119_));
 sg13g2_xnor2_1 _5889_ (.Y(_2120_),
    .A(net633),
    .B(_1431_));
 sg13g2_a221oi_1 _5890_ (.B2(net373),
    .C1(_2119_),
    .B1(_2120_),
    .A1(net365),
    .Y(_0077_),
    .A2(_2117_));
 sg13g2_nand2_1 _5891_ (.Y(_2121_),
    .A(\main.demo._q_speed[2] ),
    .B(\main.demo._q_speed[8] ));
 sg13g2_xor2_1 _5892_ (.B(\main.demo._q_speed[8] ),
    .A(\main.demo._q_speed[2] ),
    .X(_2122_));
 sg13g2_o21ai_1 _5893_ (.B1(_2114_),
    .Y(_2123_),
    .A1(_2115_),
    .A2(_2116_));
 sg13g2_nand2_1 _5894_ (.Y(_2124_),
    .A(_2122_),
    .B(_2123_));
 sg13g2_or2_1 _5895_ (.X(_2125_),
    .B(_2123_),
    .A(_2122_));
 sg13g2_nand3_1 _5896_ (.B(_2124_),
    .C(_2125_),
    .A(_2085_),
    .Y(_2126_));
 sg13g2_xnor2_1 _5897_ (.Y(_2127_),
    .A(\main.demo._q_frame[1] ),
    .B(_1434_));
 sg13g2_a21oi_1 _5898_ (.A1(net373),
    .A2(_2127_),
    .Y(_2128_),
    .B1(net364));
 sg13g2_a22oi_1 _5899_ (.Y(_0078_),
    .B1(_2126_),
    .B2(_2128_),
    .A2(net364),
    .A1(_2648_));
 sg13g2_nand2_1 _5900_ (.Y(_2129_),
    .A(\main.demo._q_speed[3] ),
    .B(\main.demo._q_speed[9] ));
 sg13g2_xnor2_1 _5901_ (.Y(_2130_),
    .A(\main.demo._q_speed[3] ),
    .B(\main.demo._q_speed[9] ));
 sg13g2_nand3_1 _5902_ (.B(_2124_),
    .C(_2130_),
    .A(_2121_),
    .Y(_2131_));
 sg13g2_a21o_1 _5903_ (.A2(_2124_),
    .A1(_2121_),
    .B1(_2130_),
    .X(_2132_));
 sg13g2_nand3_1 _5904_ (.B(_2131_),
    .C(_2132_),
    .A(_2085_),
    .Y(_2133_));
 sg13g2_o21ai_1 _5905_ (.B1(_2634_),
    .Y(_2134_),
    .A1(_1432_),
    .A2(_1433_));
 sg13g2_nor2b_1 _5906_ (.A(_1435_),
    .B_N(_2134_),
    .Y(_2135_));
 sg13g2_o21ai_1 _5907_ (.B1(_2113_),
    .Y(_2136_),
    .A1(_2085_),
    .A2(_2135_));
 sg13g2_a22oi_1 _5908_ (.Y(_0079_),
    .B1(_2133_),
    .B2(_2136_),
    .A2(net364),
    .A1(_2649_));
 sg13g2_xnor2_1 _5909_ (.Y(_2137_),
    .A(\main.demo._q_speed[10] ),
    .B(net568));
 sg13g2_a21oi_1 _5910_ (.A1(_2129_),
    .A2(_2132_),
    .Y(_2138_),
    .B1(_2137_));
 sg13g2_nand3_1 _5911_ (.B(_2132_),
    .C(_2137_),
    .A(_2129_),
    .Y(_2139_));
 sg13g2_nand2_1 _5912_ (.Y(_2140_),
    .A(net365),
    .B(_2139_));
 sg13g2_xor2_1 _5913_ (.B(_1435_),
    .A(net436),
    .X(_2141_));
 sg13g2_a22oi_1 _5914_ (.Y(_2142_),
    .B1(_2141_),
    .B2(net373),
    .A2(net364),
    .A1(net568));
 sg13g2_o21ai_1 _5915_ (.B1(_2142_),
    .Y(_0080_),
    .A1(_2138_),
    .A2(_2140_));
 sg13g2_a21o_1 _5916_ (.A2(\main.demo._q_speed[4] ),
    .A1(\main.demo._q_speed[10] ),
    .B1(_2138_),
    .X(_2143_));
 sg13g2_xor2_1 _5917_ (.B(\main.demo._q_speed[5] ),
    .A(\main.demo._q_speed[11] ),
    .X(_2144_));
 sg13g2_xnor2_1 _5918_ (.Y(_2145_),
    .A(_2143_),
    .B(_2144_));
 sg13g2_xor2_1 _5919_ (.B(_1436_),
    .A(net602),
    .X(_2146_));
 sg13g2_nand2_1 _5920_ (.Y(_2147_),
    .A(net373),
    .B(_2146_));
 sg13g2_a22oi_1 _5921_ (.Y(_2148_),
    .B1(_2147_),
    .B2(_2113_),
    .A2(_2145_),
    .A1(_2085_));
 sg13g2_a21o_1 _5922_ (.A2(net364),
    .A1(net594),
    .B1(_2148_),
    .X(_0081_));
 sg13g2_nand2_1 _5923_ (.Y(_2149_),
    .A(\main.demo._q_speed[6] ),
    .B(\main.demo._q_speed[12] ));
 sg13g2_xnor2_1 _5924_ (.Y(_2150_),
    .A(\main.demo._q_speed[6] ),
    .B(\main.demo._q_speed[12] ));
 sg13g2_a21o_1 _5925_ (.A2(\main.demo._q_speed[5] ),
    .A1(\main.demo._q_speed[11] ),
    .B1(_2143_),
    .X(_2151_));
 sg13g2_o21ai_1 _5926_ (.B1(_2151_),
    .Y(_2152_),
    .A1(\main.demo._q_speed[11] ),
    .A2(\main.demo._q_speed[5] ));
 sg13g2_xnor2_1 _5927_ (.Y(_2153_),
    .A(_2150_),
    .B(_2152_));
 sg13g2_xor2_1 _5928_ (.B(_1437_),
    .A(net637),
    .X(_2154_));
 sg13g2_a22oi_1 _5929_ (.Y(_2155_),
    .B1(_2154_),
    .B2(net373),
    .A2(net364),
    .A1(net627));
 sg13g2_o21ai_1 _5930_ (.B1(_2155_),
    .Y(_0082_),
    .A1(_2113_),
    .A2(_2153_));
 sg13g2_xor2_1 _5931_ (.B(\main.demo._q_speed[13] ),
    .A(\main.demo._q_speed[7] ),
    .X(_2156_));
 sg13g2_o21ai_1 _5932_ (.B1(_2149_),
    .Y(_2157_),
    .A1(_2150_),
    .A2(_2152_));
 sg13g2_and2_1 _5933_ (.A(_2156_),
    .B(_2157_),
    .X(_2158_));
 sg13g2_o21ai_1 _5934_ (.B1(net365),
    .Y(_2159_),
    .A1(_2156_),
    .A2(_2157_));
 sg13g2_mux2_1 _5935_ (.A0(\main.demo._q_frame[6] ),
    .A1(net392),
    .S(_1437_),
    .X(_2160_));
 sg13g2_a22oi_1 _5936_ (.Y(_2161_),
    .B1(_2160_),
    .B2(net373),
    .A2(net364),
    .A1(net642));
 sg13g2_o21ai_1 _5937_ (.B1(_2161_),
    .Y(_0083_),
    .A1(_2158_),
    .A2(_2159_));
 sg13g2_xnor2_1 _5938_ (.Y(_2162_),
    .A(\main.demo._q_speed[8] ),
    .B(\main.demo._q_speed[14] ));
 sg13g2_a21oi_1 _5939_ (.A1(\main.demo._q_speed[7] ),
    .A2(\main.demo._q_speed[13] ),
    .Y(_2163_),
    .B1(_2158_));
 sg13g2_nor2_1 _5940_ (.A(_2162_),
    .B(_2163_),
    .Y(_2164_));
 sg13g2_a21o_1 _5941_ (.A2(_2163_),
    .A1(_2162_),
    .B1(_2113_),
    .X(_2165_));
 sg13g2_xor2_1 _5942_ (.B(_1438_),
    .A(net434),
    .X(_2166_));
 sg13g2_a22oi_1 _5943_ (.Y(_2167_),
    .B1(_2166_),
    .B2(net371),
    .A2(net363),
    .A1(net622));
 sg13g2_o21ai_1 _5944_ (.B1(_2167_),
    .Y(_0084_),
    .A1(_2164_),
    .A2(_2165_));
 sg13g2_xnor2_1 _5945_ (.Y(_2168_),
    .A(net609),
    .B(_1439_));
 sg13g2_a21oi_1 _5946_ (.A1(\main.demo._q_speed[8] ),
    .A2(\main.demo._q_speed[14] ),
    .Y(_2169_),
    .B1(_2164_));
 sg13g2_nor2_1 _5947_ (.A(\main.demo._q_speed[9] ),
    .B(\main.demo._q_speed[15] ),
    .Y(_2170_));
 sg13g2_or2_1 _5948_ (.X(_2171_),
    .B(\main.demo._q_speed[15] ),
    .A(\main.demo._q_speed[9] ));
 sg13g2_nand2_1 _5949_ (.Y(_2172_),
    .A(\main.demo._q_speed[9] ),
    .B(\main.demo._q_speed[15] ));
 sg13g2_nand3_1 _5950_ (.B(_2171_),
    .C(_2172_),
    .A(_2169_),
    .Y(_2173_));
 sg13g2_a21oi_1 _5951_ (.A1(_2171_),
    .A2(_2172_),
    .Y(_2174_),
    .B1(_2169_));
 sg13g2_nor2_1 _5952_ (.A(net371),
    .B(_2174_),
    .Y(_2175_));
 sg13g2_a221oi_1 _5953_ (.B2(_2175_),
    .C1(net363),
    .B1(_2173_),
    .A1(net371),
    .Y(_2176_),
    .A2(_2168_));
 sg13g2_a21o_1 _5954_ (.A2(net363),
    .A1(net591),
    .B1(_2176_),
    .X(_0085_));
 sg13g2_o21ai_1 _5955_ (.B1(_2172_),
    .Y(_2177_),
    .A1(_2169_),
    .A2(_2170_));
 sg13g2_and2_1 _5956_ (.A(\main.demo._q_speed[10] ),
    .B(_2177_),
    .X(_2178_));
 sg13g2_o21ai_1 _5957_ (.B1(_2112_),
    .Y(_2179_),
    .A1(net583),
    .A2(_2177_));
 sg13g2_a22oi_1 _5958_ (.Y(_2180_),
    .B1(_2118_),
    .B2(net583),
    .A2(net371),
    .A1(_1442_));
 sg13g2_o21ai_1 _5959_ (.B1(_2180_),
    .Y(_0086_),
    .A1(_2178_),
    .A2(_2179_));
 sg13g2_and2_1 _5960_ (.A(\main.demo._q_speed[11] ),
    .B(_2178_),
    .X(_2181_));
 sg13g2_o21ai_1 _5961_ (.B1(net365),
    .Y(_2182_),
    .A1(net597),
    .A2(_2178_));
 sg13g2_xor2_1 _5962_ (.B(_1441_),
    .A(net624),
    .X(_2183_));
 sg13g2_a22oi_1 _5963_ (.Y(_2184_),
    .B1(_2183_),
    .B2(net372),
    .A2(net363),
    .A1(net597));
 sg13g2_o21ai_1 _5964_ (.B1(net598),
    .Y(_0087_),
    .A1(_2181_),
    .A2(_2182_));
 sg13g2_and2_1 _5965_ (.A(net592),
    .B(_2181_),
    .X(_2185_));
 sg13g2_o21ai_1 _5966_ (.B1(net365),
    .Y(_2186_),
    .A1(net592),
    .A2(_2181_));
 sg13g2_a21oi_1 _5967_ (.A1(\main.demo._q_frame[10] ),
    .A2(_1441_),
    .Y(_2187_),
    .B1(net604));
 sg13g2_nand3_1 _5968_ (.B(\main.demo._q_frame[10] ),
    .C(_1441_),
    .A(\main.demo._q_frame[11] ),
    .Y(_2188_));
 sg13g2_nor2b_1 _5969_ (.A(net605),
    .B_N(_2188_),
    .Y(_2189_));
 sg13g2_a22oi_1 _5970_ (.Y(_2190_),
    .B1(_2189_),
    .B2(net372),
    .A2(net363),
    .A1(net592));
 sg13g2_o21ai_1 _5971_ (.B1(net593),
    .Y(_0088_),
    .A1(_2185_),
    .A2(_2186_));
 sg13g2_and2_1 _5972_ (.A(net581),
    .B(_2185_),
    .X(_2191_));
 sg13g2_o21ai_1 _5973_ (.B1(net365),
    .Y(_2192_),
    .A1(net581),
    .A2(_2185_));
 sg13g2_nand4_1 _5974_ (.B(\main.demo._q_frame[10] ),
    .C(\main.demo._q_frame[12] ),
    .A(net604),
    .Y(_2193_),
    .D(_1441_));
 sg13g2_xnor2_1 _5975_ (.Y(_2194_),
    .A(net628),
    .B(_2188_));
 sg13g2_a22oi_1 _5976_ (.Y(_2195_),
    .B1(_2194_),
    .B2(net372),
    .A2(net363),
    .A1(net581));
 sg13g2_o21ai_1 _5977_ (.B1(net582),
    .Y(_0089_),
    .A1(_2191_),
    .A2(_2192_));
 sg13g2_nand2_1 _5978_ (.Y(_2196_),
    .A(\main.demo._q_speed[14] ),
    .B(_2191_));
 sg13g2_nor2_1 _5979_ (.A(net570),
    .B(_2191_),
    .Y(_2197_));
 sg13g2_nand2_1 _5980_ (.Y(_2198_),
    .A(net365),
    .B(_2196_));
 sg13g2_nor2_1 _5981_ (.A(_2647_),
    .B(_2193_),
    .Y(_2199_));
 sg13g2_xnor2_1 _5982_ (.Y(_2200_),
    .A(net613),
    .B(_2193_));
 sg13g2_a22oi_1 _5983_ (.Y(_2201_),
    .B1(_2200_),
    .B2(net371),
    .A2(net363),
    .A1(net570));
 sg13g2_o21ai_1 _5984_ (.B1(net571),
    .Y(_0090_),
    .A1(_2197_),
    .A2(_2198_));
 sg13g2_nand2_1 _5985_ (.Y(_2202_),
    .A(net498),
    .B(net363));
 sg13g2_xor2_1 _5986_ (.B(_2199_),
    .A(net595),
    .X(_2203_));
 sg13g2_a21oi_1 _5987_ (.A1(net371),
    .A2(_2203_),
    .Y(_2204_),
    .B1(net365));
 sg13g2_o21ai_1 _5988_ (.B1(_2085_),
    .Y(_2205_),
    .A1(net498),
    .A2(_2196_));
 sg13g2_a21oi_1 _5989_ (.A1(net498),
    .A2(_2196_),
    .Y(_2206_),
    .B1(_2205_));
 sg13g2_o21ai_1 _5990_ (.B1(_2202_),
    .Y(_0091_),
    .A1(_2204_),
    .A2(_2206_));
 sg13g2_nor2_1 _5991_ (.A(net402),
    .B(_2120_),
    .Y(_0092_));
 sg13g2_and2_1 _5992_ (.A(net443),
    .B(_2127_),
    .X(_0093_));
 sg13g2_and2_1 _5993_ (.A(net442),
    .B(_2135_),
    .X(_0094_));
 sg13g2_and2_1 _5994_ (.A(net442),
    .B(_2141_),
    .X(_0095_));
 sg13g2_and2_1 _5995_ (.A(net442),
    .B(net603),
    .X(_0096_));
 sg13g2_and2_1 _5996_ (.A(net442),
    .B(_2154_),
    .X(_0097_));
 sg13g2_and2_1 _5997_ (.A(net442),
    .B(_2160_),
    .X(_0098_));
 sg13g2_and2_1 _5998_ (.A(net442),
    .B(_2166_),
    .X(_0099_));
 sg13g2_nor2_1 _5999_ (.A(net402),
    .B(_2168_),
    .Y(_0100_));
 sg13g2_and2_1 _6000_ (.A(net443),
    .B(_1442_),
    .X(_0101_));
 sg13g2_and2_1 _6001_ (.A(net443),
    .B(_2183_),
    .X(_0102_));
 sg13g2_and2_1 _6002_ (.A(net443),
    .B(_2189_),
    .X(_0103_));
 sg13g2_and2_1 _6003_ (.A(net443),
    .B(net629),
    .X(_0104_));
 sg13g2_and2_1 _6004_ (.A(net443),
    .B(net614),
    .X(_0105_));
 sg13g2_and2_1 _6005_ (.A(net443),
    .B(net596),
    .X(_0106_));
 sg13g2_nor3_2 _6006_ (.A(\main.demo.zic._q_clock_count[7] ),
    .B(\main.demo.zic._q_clock_count[6] ),
    .C(\main.demo.zic._q_clock_count[8] ),
    .Y(_2207_));
 sg13g2_nor2_1 _6007_ (.A(\main.demo.zic._q_clock_count[1] ),
    .B(net577),
    .Y(_2208_));
 sg13g2_nor4_2 _6008_ (.A(\main.demo.zic._q_clock_count[3] ),
    .B(\main.demo.zic._q_clock_count[2] ),
    .C(\main.demo.zic._q_clock_count[5] ),
    .Y(_2209_),
    .D(\main.demo.zic._q_clock_count[4] ));
 sg13g2_and3_1 _6009_ (.X(_2210_),
    .A(_2207_),
    .B(_2208_),
    .C(_2209_));
 sg13g2_nand3_1 _6010_ (.B(_2208_),
    .C(_2209_),
    .A(_2207_),
    .Y(_2211_));
 sg13g2_nor2b_2 _6011_ (.A(\main.demo.zic._q_idx[5] ),
    .B_N(\main.demo.zic._q_idx[6] ),
    .Y(_2212_));
 sg13g2_and2_1 _6012_ (.A(\main.demo.zic._q_idx[4] ),
    .B(_2212_),
    .X(_2213_));
 sg13g2_nand2_2 _6013_ (.Y(_2214_),
    .A(\main.demo.zic._q_idx[4] ),
    .B(_2212_));
 sg13g2_and2_2 _6014_ (.A(net409),
    .B(net410),
    .X(_2215_));
 sg13g2_nand2_1 _6015_ (.Y(_2216_),
    .A(net408),
    .B(net410));
 sg13g2_nor2_2 _6016_ (.A(\main.demo.zic._q_idx[1] ),
    .B(\main.demo.zic._q_idx[0] ),
    .Y(_2217_));
 sg13g2_nand2_2 _6017_ (.Y(_2218_),
    .A(net410),
    .B(_2217_));
 sg13g2_nand2_2 _6018_ (.Y(_2219_),
    .A(_2215_),
    .B(_2217_));
 sg13g2_nor2b_2 _6019_ (.A(\main.demo.zic._q_idx[1] ),
    .B_N(\main.demo.zic._q_idx[0] ),
    .Y(_2220_));
 sg13g2_nand2_2 _6020_ (.Y(_2221_),
    .A(net411),
    .B(_2220_));
 sg13g2_nor2_1 _6021_ (.A(net408),
    .B(_2221_),
    .Y(_2222_));
 sg13g2_o21ai_1 _6022_ (.B1(_2219_),
    .Y(_2223_),
    .A1(net409),
    .A2(_2221_));
 sg13g2_nand2_1 _6023_ (.Y(_2224_),
    .A(_2213_),
    .B(_2223_));
 sg13g2_nand2_1 _6024_ (.Y(_2225_),
    .A(\main.demo.zic._q_idx[5] ),
    .B(_0035_));
 sg13g2_nand3_1 _6025_ (.B(\main.demo.zic._q_idx[4] ),
    .C(_0035_),
    .A(\main.demo.zic._q_idx[5] ),
    .Y(_2226_));
 sg13g2_o21ai_1 _6026_ (.B1(_2224_),
    .Y(_2227_),
    .A1(_2221_),
    .A2(_2226_));
 sg13g2_nand2_2 _6027_ (.Y(_2228_),
    .A(_2619_),
    .B(_2212_));
 sg13g2_inv_1 _6028_ (.Y(_2229_),
    .A(_2228_));
 sg13g2_nand2b_2 _6029_ (.Y(_2230_),
    .B(\main.demo.zic._q_idx[1] ),
    .A_N(\main.demo.zic._q_idx[0] ));
 sg13g2_nor3_2 _6030_ (.A(net409),
    .B(_2618_),
    .C(_2230_),
    .Y(_2231_));
 sg13g2_nand2_2 _6031_ (.Y(_2232_),
    .A(\main.demo.zic._q_idx[1] ),
    .B(\main.demo.zic._q_idx[0] ));
 sg13g2_nor2_1 _6032_ (.A(net408),
    .B(_2232_),
    .Y(_2233_));
 sg13g2_nor2_2 _6033_ (.A(net408),
    .B(net411),
    .Y(_2234_));
 sg13g2_nor3_2 _6034_ (.A(net408),
    .B(net410),
    .C(_2232_),
    .Y(_2235_));
 sg13g2_nor2_1 _6035_ (.A(_2231_),
    .B(_2235_),
    .Y(_2236_));
 sg13g2_inv_1 _6036_ (.Y(_2237_),
    .A(_2236_));
 sg13g2_nand2_1 _6037_ (.Y(_2238_),
    .A(_2217_),
    .B(_2234_));
 sg13g2_nor2b_2 _6038_ (.A(net410),
    .B_N(net409),
    .Y(_2239_));
 sg13g2_a22oi_1 _6039_ (.Y(_2240_),
    .B1(_2239_),
    .B2(_2220_),
    .A2(_2234_),
    .A1(_2217_));
 sg13g2_a21oi_1 _6040_ (.A1(_2236_),
    .A2(_2240_),
    .Y(_2241_),
    .B1(_2228_));
 sg13g2_nand2b_2 _6041_ (.Y(_2242_),
    .B(_2619_),
    .A_N(_2225_));
 sg13g2_nand2_1 _6042_ (.Y(_2243_),
    .A(_2228_),
    .B(_2242_));
 sg13g2_nand2_1 _6043_ (.Y(_2244_),
    .A(_2222_),
    .B(_2243_));
 sg13g2_o21ai_1 _6044_ (.B1(_2244_),
    .Y(_2245_),
    .A1(_2219_),
    .A2(_2242_));
 sg13g2_nor2b_1 _6045_ (.A(_2232_),
    .B_N(_2239_),
    .Y(_2246_));
 sg13g2_nor2_1 _6046_ (.A(net410),
    .B(_2230_),
    .Y(_2247_));
 sg13g2_nor2b_1 _6047_ (.A(_2230_),
    .B_N(_2234_),
    .Y(_2248_));
 sg13g2_nor2_1 _6048_ (.A(_2246_),
    .B(_2248_),
    .Y(_2249_));
 sg13g2_nand2_1 _6049_ (.Y(_2250_),
    .A(_2217_),
    .B(_2239_));
 sg13g2_nor2b_1 _6050_ (.A(_2231_),
    .B_N(_2250_),
    .Y(_2251_));
 sg13g2_a21oi_1 _6051_ (.A1(_2249_),
    .A2(_2251_),
    .Y(_2252_),
    .B1(_2242_));
 sg13g2_nand2_1 _6052_ (.Y(_2253_),
    .A(_2220_),
    .B(_2234_));
 sg13g2_a21oi_1 _6053_ (.A1(_2214_),
    .A2(_2242_),
    .Y(_2254_),
    .B1(_2253_));
 sg13g2_nor4_2 _6054_ (.A(_2241_),
    .B(_2245_),
    .C(_2252_),
    .Y(_2255_),
    .D(_2254_));
 sg13g2_nand2_1 _6055_ (.Y(_2256_),
    .A(net411),
    .B(_2233_));
 sg13g2_nand2_1 _6056_ (.Y(_2257_),
    .A(_2250_),
    .B(_2256_));
 sg13g2_nor2_1 _6057_ (.A(_2247_),
    .B(_2257_),
    .Y(_2258_));
 sg13g2_a21oi_1 _6058_ (.A1(_2253_),
    .A2(_2258_),
    .Y(_2259_),
    .B1(_2226_));
 sg13g2_or2_1 _6059_ (.X(_2260_),
    .B(_2230_),
    .A(_2216_));
 sg13g2_nor2_1 _6060_ (.A(_2228_),
    .B(_2260_),
    .Y(_2261_));
 sg13g2_nor2_1 _6061_ (.A(_2218_),
    .B(_2226_),
    .Y(_2262_));
 sg13g2_nor3_2 _6062_ (.A(_2259_),
    .B(_2261_),
    .C(_2262_),
    .Y(_2263_));
 sg13g2_nand2_2 _6063_ (.Y(_2264_),
    .A(_2255_),
    .B(_2263_));
 sg13g2_a21oi_1 _6064_ (.A1(\main.demo.zic._q_idx[0] ),
    .A2(_2239_),
    .Y(_2265_),
    .B1(_2237_));
 sg13g2_nand2_1 _6065_ (.Y(_2266_),
    .A(_2214_),
    .B(_2225_));
 sg13g2_o21ai_1 _6066_ (.B1(_2260_),
    .Y(_2267_),
    .A1(_2214_),
    .A2(_2265_));
 sg13g2_nand2_1 _6067_ (.Y(_2268_),
    .A(_2266_),
    .B(_2267_));
 sg13g2_a21oi_1 _6068_ (.A1(_2238_),
    .A2(_2265_),
    .Y(_2269_),
    .B1(_2226_));
 sg13g2_nor2b_1 _6069_ (.A(_2212_),
    .B_N(_2225_),
    .Y(_2270_));
 sg13g2_nor2_2 _6070_ (.A(_2216_),
    .B(_2232_),
    .Y(_2271_));
 sg13g2_or2_1 _6071_ (.X(_2272_),
    .B(_2232_),
    .A(_2216_));
 sg13g2_nor2_1 _6072_ (.A(_2270_),
    .B(_2272_),
    .Y(_2273_));
 sg13g2_nor2_1 _6073_ (.A(_2214_),
    .B(_2258_),
    .Y(_2274_));
 sg13g2_nor3_1 _6074_ (.A(_2269_),
    .B(_2273_),
    .C(_2274_),
    .Y(_2275_));
 sg13g2_and2_1 _6075_ (.A(_2268_),
    .B(_2275_),
    .X(_2276_));
 sg13g2_nand2b_1 _6076_ (.Y(_2277_),
    .B(_2240_),
    .A_N(_2233_));
 sg13g2_o21ai_1 _6077_ (.B1(_2242_),
    .Y(_2278_),
    .A1(_2214_),
    .A2(_2238_));
 sg13g2_nand2_1 _6078_ (.Y(_2279_),
    .A(_2277_),
    .B(_2278_));
 sg13g2_nand3_1 _6079_ (.B(_2249_),
    .C(_2253_),
    .A(_2218_),
    .Y(_2280_));
 sg13g2_o21ai_1 _6080_ (.B1(_2229_),
    .Y(_2281_),
    .A1(_2257_),
    .A2(_2280_));
 sg13g2_inv_1 _6081_ (.Y(_2282_),
    .A(_2281_));
 sg13g2_nor2_1 _6082_ (.A(net408),
    .B(_2218_),
    .Y(_2283_));
 sg13g2_a21oi_1 _6083_ (.A1(_2215_),
    .A2(_2220_),
    .Y(_2284_),
    .B1(_2283_));
 sg13g2_nor2_1 _6084_ (.A(_2214_),
    .B(_2284_),
    .Y(_2285_));
 sg13g2_nor2_1 _6085_ (.A(_2227_),
    .B(_2285_),
    .Y(_2286_));
 sg13g2_or2_1 _6086_ (.X(_2287_),
    .B(\main.demo.zic._q_idx[6] ),
    .A(\main.demo.zic._q_idx[5] ));
 sg13g2_o21ai_1 _6087_ (.B1(_2221_),
    .Y(_2288_),
    .A1(net410),
    .A2(_2230_));
 sg13g2_nand3_1 _6088_ (.B(_2243_),
    .C(_2288_),
    .A(net408),
    .Y(_2289_));
 sg13g2_nand4_1 _6089_ (.B(_2281_),
    .C(_2287_),
    .A(_2279_),
    .Y(_2290_),
    .D(_2289_));
 sg13g2_nor4_1 _6090_ (.A(_2227_),
    .B(_2264_),
    .C(_2285_),
    .D(_2290_),
    .Y(_2291_));
 sg13g2_a21o_1 _6091_ (.A2(_2291_),
    .A1(_2276_),
    .B1(_2227_),
    .X(_2292_));
 sg13g2_nand2_1 _6092_ (.Y(_2293_),
    .A(_2255_),
    .B(_2268_));
 sg13g2_or2_1 _6093_ (.X(_2294_),
    .B(_2293_),
    .A(_2292_));
 sg13g2_a21oi_1 _6094_ (.A1(net376),
    .A2(_2294_),
    .Y(_2295_),
    .B1(net299));
 sg13g2_nand2_1 _6095_ (.Y(_2296_),
    .A(net299),
    .B(_2294_));
 sg13g2_o21ai_1 _6096_ (.B1(net437),
    .Y(_2297_),
    .A1(_2211_),
    .A2(_2296_));
 sg13g2_nor2_1 _6097_ (.A(_2295_),
    .B(_2297_),
    .Y(_0107_));
 sg13g2_nor3_1 _6098_ (.A(_2227_),
    .B(_2245_),
    .C(_2262_),
    .Y(_2298_));
 sg13g2_nand3_1 _6099_ (.B(_2281_),
    .C(_2298_),
    .A(_2276_),
    .Y(_2299_));
 sg13g2_nor2b_1 _6100_ (.A(_0029_),
    .B_N(_2299_),
    .Y(_2300_));
 sg13g2_xor2_1 _6101_ (.B(_2299_),
    .A(_0029_),
    .X(_2301_));
 sg13g2_nor2_1 _6102_ (.A(_2296_),
    .B(_2301_),
    .Y(_2302_));
 sg13g2_xnor2_1 _6103_ (.Y(_2303_),
    .A(_2296_),
    .B(_2301_));
 sg13g2_o21ai_1 _6104_ (.B1(net437),
    .Y(_2304_),
    .A1(net332),
    .A2(net375));
 sg13g2_a21oi_1 _6105_ (.A1(net375),
    .A2(_2303_),
    .Y(_0108_),
    .B1(_2304_));
 sg13g2_or2_1 _6106_ (.X(_2305_),
    .B(_2228_),
    .A(_2218_));
 sg13g2_nand4_1 _6107_ (.B(_2275_),
    .C(_2286_),
    .A(_2263_),
    .Y(_2306_),
    .D(_2305_));
 sg13g2_nand2_1 _6108_ (.Y(_2307_),
    .A(\main.demo.zic._q_qpos[2] ),
    .B(_2306_));
 sg13g2_xor2_1 _6109_ (.B(_2306_),
    .A(\main.demo.zic._q_qpos[2] ),
    .X(_2308_));
 sg13g2_or3_1 _6110_ (.A(_2300_),
    .B(_2302_),
    .C(_2308_),
    .X(_2309_));
 sg13g2_o21ai_1 _6111_ (.B1(_2308_),
    .Y(_2310_),
    .A1(_2300_),
    .A2(_2302_));
 sg13g2_a21oi_1 _6112_ (.A1(_2309_),
    .A2(_2310_),
    .Y(_2311_),
    .B1(_2211_));
 sg13g2_o21ai_1 _6113_ (.B1(net438),
    .Y(_2312_),
    .A1(net546),
    .A2(net375));
 sg13g2_nor2_1 _6114_ (.A(_2311_),
    .B(_2312_),
    .Y(_0109_));
 sg13g2_nand3b_1 _6115_ (.B(_2268_),
    .C(_2263_),
    .Y(_2313_),
    .A_N(_2285_));
 sg13g2_nor2b_1 _6116_ (.A(_0030_),
    .B_N(_2313_),
    .Y(_2314_));
 sg13g2_xor2_1 _6117_ (.B(_2313_),
    .A(_0030_),
    .X(_2315_));
 sg13g2_and3_1 _6118_ (.X(_2316_),
    .A(_2307_),
    .B(_2310_),
    .C(_2315_));
 sg13g2_a21oi_1 _6119_ (.A1(_2307_),
    .A2(_2310_),
    .Y(_2317_),
    .B1(_2315_));
 sg13g2_o21ai_1 _6120_ (.B1(net376),
    .Y(_2318_),
    .A1(_2316_),
    .A2(_2317_));
 sg13g2_o21ai_1 _6121_ (.B1(net438),
    .Y(_2319_),
    .A1(net318),
    .A2(net376));
 sg13g2_nor2b_1 _6122_ (.A(_2319_),
    .B_N(_2318_),
    .Y(_0110_));
 sg13g2_nand2_1 _6123_ (.Y(_2320_),
    .A(_2275_),
    .B(_2279_));
 sg13g2_nor2_1 _6124_ (.A(_2292_),
    .B(_2320_),
    .Y(_2321_));
 sg13g2_o21ai_1 _6125_ (.B1(\main.demo.zic._q_qpos[4] ),
    .Y(_2322_),
    .A1(_2292_),
    .A2(_2320_));
 sg13g2_xnor2_1 _6126_ (.Y(_2323_),
    .A(\main.demo.zic._q_qpos[4] ),
    .B(_2321_));
 sg13g2_or3_1 _6127_ (.A(_2314_),
    .B(_2317_),
    .C(_2323_),
    .X(_2324_));
 sg13g2_o21ai_1 _6128_ (.B1(_2323_),
    .Y(_2325_),
    .A1(_2314_),
    .A2(_2317_));
 sg13g2_a21oi_1 _6129_ (.A1(_2324_),
    .A2(_2325_),
    .Y(_2326_),
    .B1(_2211_));
 sg13g2_o21ai_1 _6130_ (.B1(net437),
    .Y(_2327_),
    .A1(net547),
    .A2(net375));
 sg13g2_nor2_1 _6131_ (.A(_2326_),
    .B(_2327_),
    .Y(_0111_));
 sg13g2_xnor2_1 _6132_ (.Y(_2328_),
    .A(_2667_),
    .B(_2264_));
 sg13g2_and3_1 _6133_ (.X(_2329_),
    .A(_2322_),
    .B(_2325_),
    .C(_2328_));
 sg13g2_a21oi_1 _6134_ (.A1(_2322_),
    .A2(_2325_),
    .Y(_2330_),
    .B1(_2328_));
 sg13g2_o21ai_1 _6135_ (.B1(net379),
    .Y(_2331_),
    .A1(_2329_),
    .A2(_2330_));
 sg13g2_o21ai_1 _6136_ (.B1(net438),
    .Y(_2332_),
    .A1(net317),
    .A2(net379));
 sg13g2_nor2b_1 _6137_ (.A(_2332_),
    .B_N(_2331_),
    .Y(_0112_));
 sg13g2_xor2_1 _6138_ (.B(_2281_),
    .A(\main.demo.zic._q_qpos[6] ),
    .X(_2333_));
 sg13g2_a21oi_1 _6139_ (.A1(_2667_),
    .A2(_2264_),
    .Y(_2334_),
    .B1(_2330_));
 sg13g2_nor2_1 _6140_ (.A(_2333_),
    .B(_2334_),
    .Y(_2335_));
 sg13g2_xnor2_1 _6141_ (.Y(_2336_),
    .A(_2333_),
    .B(_2334_));
 sg13g2_o21ai_1 _6142_ (.B1(net438),
    .Y(_2337_),
    .A1(net564),
    .A2(net376));
 sg13g2_a21oi_1 _6143_ (.A1(net376),
    .A2(_2336_),
    .Y(_0113_),
    .B1(_2337_));
 sg13g2_a21oi_2 _6144_ (.B1(_2335_),
    .Y(_2338_),
    .A2(_2282_),
    .A1(\main.demo.zic._q_qpos[6] ));
 sg13g2_nor3_2 _6145_ (.A(_0032_),
    .B(_2211_),
    .C(_2338_),
    .Y(_2339_));
 sg13g2_and3_1 _6146_ (.X(_2340_),
    .A(_0032_),
    .B(net378),
    .C(_2338_));
 sg13g2_o21ai_1 _6147_ (.B1(net439),
    .Y(_2341_),
    .A1(net329),
    .A2(net377));
 sg13g2_nor3_1 _6148_ (.A(_2339_),
    .B(_2340_),
    .C(net330),
    .Y(_0114_));
 sg13g2_and2_1 _6149_ (.A(net462),
    .B(_2339_),
    .X(_2342_));
 sg13g2_o21ai_1 _6150_ (.B1(net439),
    .Y(_2343_),
    .A1(net462),
    .A2(_2339_));
 sg13g2_nor2_1 _6151_ (.A(_2342_),
    .B(net463),
    .Y(_0115_));
 sg13g2_nand2_1 _6152_ (.Y(_2344_),
    .A(net545),
    .B(_2342_));
 sg13g2_o21ai_1 _6153_ (.B1(net441),
    .Y(_2345_),
    .A1(net545),
    .A2(_2342_));
 sg13g2_nor2b_1 _6154_ (.A(_2345_),
    .B_N(_2344_),
    .Y(_0116_));
 sg13g2_nand3_1 _6155_ (.B(net545),
    .C(_2342_),
    .A(net310),
    .Y(_2346_));
 sg13g2_nand2_1 _6156_ (.Y(_2347_),
    .A(net441),
    .B(_2346_));
 sg13g2_a21oi_1 _6157_ (.A1(_2617_),
    .A2(_2344_),
    .Y(_0117_),
    .B1(_2347_));
 sg13g2_nand2b_1 _6158_ (.Y(_2348_),
    .B(_2346_),
    .A_N(net479));
 sg13g2_nand4_1 _6159_ (.B(net310),
    .C(\main.demo.zic._q_qpos[9] ),
    .A(net479),
    .Y(_2349_),
    .D(_2342_));
 sg13g2_and3_1 _6160_ (.X(_0118_),
    .A(net441),
    .B(_2348_),
    .C(net480));
 sg13g2_o21ai_1 _6161_ (.B1(net441),
    .Y(_2350_),
    .A1(_2616_),
    .A2(net480));
 sg13g2_a21oi_1 _6162_ (.A1(_2616_),
    .A2(net480),
    .Y(_0119_),
    .B1(_2350_));
 sg13g2_a21oi_1 _6163_ (.A1(_0917_),
    .A2(_1440_),
    .Y(_2351_),
    .B1(_2194_));
 sg13g2_o21ai_1 _6164_ (.B1(net444),
    .Y(_2352_),
    .A1(net296),
    .A2(_2351_));
 sg13g2_a21oi_1 _6165_ (.A1(_2615_),
    .A2(_2351_),
    .Y(_0120_),
    .B1(net297));
 sg13g2_mux2_1 _6166_ (.A0(net421),
    .A1(net541),
    .S(_1440_),
    .X(_2353_));
 sg13g2_and3_1 _6167_ (.X(_0121_),
    .A(net442),
    .B(\main.demo._q_go ),
    .C(_2353_));
 sg13g2_nand3_1 _6168_ (.B(net636),
    .C(_0970_),
    .A(net442),
    .Y(_2354_));
 sg13g2_a21oi_1 _6169_ (.A1(net386),
    .A2(_1440_),
    .Y(_2355_),
    .B1(_2354_));
 sg13g2_o21ai_1 _6170_ (.B1(_2355_),
    .Y(_0122_),
    .A1(net405),
    .A2(_1440_));
 sg13g2_nand4_1 _6171_ (.B(net435),
    .C(net436),
    .A(net434),
    .Y(_2356_),
    .D(_2938_));
 sg13g2_nand4_1 _6172_ (.B(\main.demo._q_frame[1] ),
    .C(\main.demo._q_frame[0] ),
    .A(\main.demo._q_frame[2] ),
    .Y(_2357_),
    .D(\main.demo._q_frame[8] ));
 sg13g2_o21ai_1 _6173_ (.B1(\main.demo._q_go ),
    .Y(_2358_),
    .A1(_2356_),
    .A2(_2357_));
 sg13g2_nand2_1 _6174_ (.Y(_2359_),
    .A(\main.demo._q_th[0] ),
    .B(_1432_));
 sg13g2_nand2_1 _6175_ (.Y(_2360_),
    .A(net289),
    .B(_1431_));
 sg13g2_a21oi_1 _6176_ (.A1(_2359_),
    .A2(net290),
    .Y(_0123_),
    .B1(net370));
 sg13g2_and3_1 _6177_ (.X(_2361_),
    .A(net306),
    .B(\main.demo._q_th[0] ),
    .C(_1431_));
 sg13g2_a21oi_1 _6178_ (.A1(\main.demo._q_th[0] ),
    .A2(_1431_),
    .Y(_2362_),
    .B1(net306));
 sg13g2_nor3_1 _6179_ (.A(net370),
    .B(_2361_),
    .C(net307),
    .Y(_0124_));
 sg13g2_and2_1 _6180_ (.A(net573),
    .B(_2361_),
    .X(_2363_));
 sg13g2_nor2_1 _6181_ (.A(net573),
    .B(_2361_),
    .Y(_2364_));
 sg13g2_nor3_1 _6182_ (.A(net370),
    .B(_2363_),
    .C(net574),
    .Y(_0125_));
 sg13g2_nor2_1 _6183_ (.A(net608),
    .B(_2363_),
    .Y(_2365_));
 sg13g2_and2_1 _6184_ (.A(net608),
    .B(_2363_),
    .X(_2366_));
 sg13g2_nor3_1 _6185_ (.A(net370),
    .B(_2365_),
    .C(_2366_),
    .Y(_0126_));
 sg13g2_nor2_1 _6186_ (.A(net523),
    .B(_2366_),
    .Y(_2367_));
 sg13g2_and2_1 _6187_ (.A(net523),
    .B(_2366_),
    .X(_2368_));
 sg13g2_nor3_1 _6188_ (.A(net370),
    .B(_2367_),
    .C(_2368_),
    .Y(_0127_));
 sg13g2_nor2_1 _6189_ (.A(net539),
    .B(_2368_),
    .Y(_2369_));
 sg13g2_and2_1 _6190_ (.A(net539),
    .B(_2368_),
    .X(_2370_));
 sg13g2_nor3_1 _6191_ (.A(net370),
    .B(_2369_),
    .C(_2370_),
    .Y(_0128_));
 sg13g2_xnor2_1 _6192_ (.Y(_2371_),
    .A(net527),
    .B(_2370_));
 sg13g2_nor2_1 _6193_ (.A(net370),
    .B(net528),
    .Y(_0129_));
 sg13g2_and2_1 _6194_ (.A(_2661_),
    .B(_2370_),
    .X(_2372_));
 sg13g2_xnor2_1 _6195_ (.Y(_2373_),
    .A(net312),
    .B(_2372_));
 sg13g2_nor2_1 _6196_ (.A(net370),
    .B(_2373_),
    .Y(_0130_));
 sg13g2_nand3_1 _6197_ (.B(\main.demo._q_th[6] ),
    .C(_2370_),
    .A(net312),
    .Y(_2374_));
 sg13g2_xor2_1 _6198_ (.B(net313),
    .A(\main.demo._q_th[8] ),
    .X(_2375_));
 sg13g2_nor2_1 _6199_ (.A(_2358_),
    .B(net314),
    .Y(_0131_));
 sg13g2_mux4_1 _6200_ (.S0(net424),
    .A0(net467),
    .A1(net283),
    .A2(net281),
    .A3(\main.demo._d_prev_b[3] ),
    .S1(net423),
    .X(_2376_));
 sg13g2_and2_1 _6201_ (.A(net457),
    .B(_2376_),
    .X(_0132_));
 sg13g2_and2_1 _6202_ (.A(net457),
    .B(\main.demo._d_prev_b[1] ),
    .X(_0133_));
 sg13g2_mux4_1 _6203_ (.S0(net424),
    .A0(net285),
    .A1(net281),
    .A2(net283),
    .A3(net467),
    .S1(net423),
    .X(_2377_));
 sg13g2_and2_1 _6204_ (.A(net457),
    .B(_2377_),
    .X(_0134_));
 sg13g2_mux4_1 _6205_ (.S0(net424),
    .A0(net497),
    .A1(net280),
    .A2(net279),
    .A3(net282),
    .S1(net423),
    .X(_2378_));
 sg13g2_and2_1 _6206_ (.A(net457),
    .B(_2378_),
    .X(_0135_));
 sg13g2_and2_1 _6207_ (.A(net457),
    .B(\main.demo._d_prev_b[0] ),
    .X(_0136_));
 sg13g2_mux4_1 _6208_ (.S0(net424),
    .A0(net282),
    .A1(net279),
    .A2(net280),
    .A3(net497),
    .S1(net423),
    .X(_2379_));
 sg13g2_and2_1 _6209_ (.A(net457),
    .B(_2379_),
    .X(_0137_));
 sg13g2_nand2b_1 _6210_ (.Y(_2380_),
    .B(\main.demo.zic._q_rythm_count[12] ),
    .A_N(\main.demo.zic._q_rythm_count[11] ));
 sg13g2_nor4_2 _6211_ (.A(_2607_),
    .B(\main.demo.zic._q_rythm_count[9] ),
    .C(\main.demo.zic._q_rythm_count[8] ),
    .Y(_2381_),
    .D(_2380_));
 sg13g2_or4_2 _6212_ (.A(_2607_),
    .B(\main.demo.zic._q_rythm_count[9] ),
    .C(\main.demo.zic._q_rythm_count[8] ),
    .D(_2380_),
    .X(_2382_));
 sg13g2_nor4_1 _6213_ (.A(\main.demo.zic._q_rythm_count[7] ),
    .B(\main.demo.zic._q_rythm_count[6] ),
    .C(\main.demo.zic._q_rythm_count[5] ),
    .D(\main.demo.zic._q_rythm_count[4] ),
    .Y(_2383_));
 sg13g2_nor4_1 _6214_ (.A(\main.demo.zic._q_rythm_count[3] ),
    .B(\main.demo.zic._q_rythm_count[2] ),
    .C(\main.demo.zic._q_rythm_count[1] ),
    .D(\main.demo.zic._q_rythm_count[0] ),
    .Y(_2384_));
 sg13g2_and2_2 _6215_ (.A(_2383_),
    .B(_2384_),
    .X(_2385_));
 sg13g2_a21oi_2 _6216_ (.B1(_2381_),
    .Y(_2386_),
    .A2(_2385_),
    .A1(net379));
 sg13g2_a21oi_2 _6217_ (.B1(_2382_),
    .Y(_2387_),
    .A2(_2271_),
    .A1(_2213_));
 sg13g2_nand3_1 _6218_ (.B(\main.demo.zic._q_idx[4] ),
    .C(_2271_),
    .A(\main.demo.zic._q_idx[5] ),
    .Y(_2388_));
 sg13g2_xor2_1 _6219_ (.B(_2388_),
    .A(_0035_),
    .X(_2389_));
 sg13g2_a22oi_1 _6220_ (.Y(_2390_),
    .B1(_2387_),
    .B2(_2389_),
    .A2(_2382_),
    .A1(net589));
 sg13g2_inv_1 _6221_ (.Y(_2391_),
    .A(_2390_));
 sg13g2_nor2_1 _6222_ (.A(_0034_),
    .B(_2272_),
    .Y(_2392_));
 sg13g2_xnor2_1 _6223_ (.Y(_2393_),
    .A(\main.demo.zic._q_idx[5] ),
    .B(_2392_));
 sg13g2_a22oi_1 _6224_ (.Y(_2394_),
    .B1(_2387_),
    .B2(_2393_),
    .A2(_2382_),
    .A1(net619));
 sg13g2_nand2_1 _6225_ (.Y(_2395_),
    .A(_2390_),
    .B(_2394_));
 sg13g2_nor2_2 _6226_ (.A(_2232_),
    .B(_2382_),
    .Y(_2396_));
 sg13g2_nor2_1 _6227_ (.A(net411),
    .B(_2396_),
    .Y(_2397_));
 sg13g2_nand2_2 _6228_ (.Y(_2398_),
    .A(net411),
    .B(_2396_));
 sg13g2_nor2b_1 _6229_ (.A(_2397_),
    .B_N(_2398_),
    .Y(_2399_));
 sg13g2_nand2b_2 _6230_ (.Y(_2400_),
    .B(_2398_),
    .A_N(_2397_));
 sg13g2_and2_1 _6231_ (.A(net409),
    .B(_2399_),
    .X(_2401_));
 sg13g2_xnor2_1 _6232_ (.Y(_2402_),
    .A(\main.demo.zic._q_idx[0] ),
    .B(_2382_));
 sg13g2_nand2_1 _6233_ (.Y(_2403_),
    .A(\main.demo.zic._q_idx[1] ),
    .B(_2402_));
 sg13g2_nand2_1 _6234_ (.Y(_2404_),
    .A(_0034_),
    .B(_2272_));
 sg13g2_nand3b_1 _6235_ (.B(_2404_),
    .C(_2387_),
    .Y(_2405_),
    .A_N(_2392_));
 sg13g2_o21ai_1 _6236_ (.B1(_2405_),
    .Y(_2406_),
    .A1(_2619_),
    .A2(_2381_));
 sg13g2_nor2_1 _6237_ (.A(_2403_),
    .B(_2406_),
    .Y(_2407_));
 sg13g2_or2_1 _6238_ (.X(_2408_),
    .B(_2407_),
    .A(_2220_));
 sg13g2_xnor2_1 _6239_ (.Y(_2409_),
    .A(net409),
    .B(_2398_));
 sg13g2_nor2_1 _6240_ (.A(net409),
    .B(_2400_),
    .Y(_2410_));
 sg13g2_a21oi_1 _6241_ (.A1(\main.demo.zic._q_idx[0] ),
    .A2(_2381_),
    .Y(_2411_),
    .B1(net640));
 sg13g2_or2_2 _6242_ (.X(_2412_),
    .B(_2411_),
    .A(_2396_));
 sg13g2_nor2_1 _6243_ (.A(_2402_),
    .B(_2412_),
    .Y(_2413_));
 sg13g2_nand2_1 _6244_ (.Y(_2414_),
    .A(_2239_),
    .B(_2413_));
 sg13g2_o21ai_1 _6245_ (.B1(_2413_),
    .Y(_2415_),
    .A1(_2239_),
    .A2(_2410_));
 sg13g2_nand3b_1 _6246_ (.B(_2413_),
    .C(_2400_),
    .Y(_2416_),
    .A_N(_2409_));
 sg13g2_nand3_1 _6247_ (.B(_2415_),
    .C(_2416_),
    .A(_2403_),
    .Y(_2417_));
 sg13g2_a22oi_1 _6248_ (.Y(_2418_),
    .B1(_2417_),
    .B2(_2406_),
    .A2(_2408_),
    .A1(_2401_));
 sg13g2_or2_1 _6249_ (.X(_2419_),
    .B(_2418_),
    .A(_2395_));
 sg13g2_or3_1 _6250_ (.A(_2390_),
    .B(_2394_),
    .C(_2412_),
    .X(_2420_));
 sg13g2_nor2_1 _6251_ (.A(_2391_),
    .B(_2394_),
    .Y(_2421_));
 sg13g2_nand3_1 _6252_ (.B(_2403_),
    .C(_2409_),
    .A(_2400_),
    .Y(_2422_));
 sg13g2_o21ai_1 _6253_ (.B1(_2412_),
    .Y(_2423_),
    .A1(_2399_),
    .A2(_2409_));
 sg13g2_nand2b_1 _6254_ (.Y(_2424_),
    .B(_2422_),
    .A_N(_2423_));
 sg13g2_nor3_1 _6255_ (.A(_2215_),
    .B(_2395_),
    .C(_2412_),
    .Y(_2425_));
 sg13g2_a21oi_1 _6256_ (.A1(_2410_),
    .A2(_2421_),
    .Y(_2426_),
    .B1(_2425_));
 sg13g2_o21ai_1 _6257_ (.B1(_2381_),
    .Y(_2427_),
    .A1(_2406_),
    .A2(_2426_));
 sg13g2_a21oi_1 _6258_ (.A1(_2421_),
    .A2(_2424_),
    .Y(_2428_),
    .B1(_2427_));
 sg13g2_nand3_1 _6259_ (.B(_2420_),
    .C(_2428_),
    .A(_2419_),
    .Y(_2429_));
 sg13g2_nor3_1 _6260_ (.A(\main.demo.zic._q_drum_inc[0] ),
    .B(\main.demo.zic._q_drum_inc[1] ),
    .C(\main.demo.zic._q_drum_inc[2] ),
    .Y(_2430_));
 sg13g2_a21oi_1 _6261_ (.A1(_2664_),
    .A2(_2430_),
    .Y(_2431_),
    .B1(_2381_));
 sg13g2_a21oi_1 _6262_ (.A1(_2662_),
    .A2(_2431_),
    .Y(_2432_),
    .B1(net369));
 sg13g2_a22oi_1 _6263_ (.Y(_0138_),
    .B1(_2429_),
    .B2(_2432_),
    .A2(net369),
    .A1(_2662_));
 sg13g2_xnor2_1 _6264_ (.Y(_2433_),
    .A(\main.demo.zic._q_drum_inc[0] ),
    .B(net607));
 sg13g2_a21oi_1 _6265_ (.A1(_2431_),
    .A2(_2433_),
    .Y(_2434_),
    .B1(net369));
 sg13g2_a22oi_1 _6266_ (.Y(_0139_),
    .B1(_2429_),
    .B2(_2434_),
    .A2(net369),
    .A1(_2663_));
 sg13g2_o21ai_1 _6267_ (.B1(\main.demo.zic._q_drum_inc[2] ),
    .Y(_2435_),
    .A1(\main.demo.zic._q_drum_inc[0] ),
    .A2(net644));
 sg13g2_nand2b_1 _6268_ (.Y(_2436_),
    .B(_2435_),
    .A_N(_2430_));
 sg13g2_a21oi_1 _6269_ (.A1(_2431_),
    .A2(_2436_),
    .Y(_2437_),
    .B1(net369));
 sg13g2_a22oi_1 _6270_ (.Y(_0140_),
    .B1(_2429_),
    .B2(_2437_),
    .A2(net369),
    .A1(_2665_));
 sg13g2_nor3_1 _6271_ (.A(_2664_),
    .B(_2381_),
    .C(_2430_),
    .Y(_2438_));
 sg13g2_nor2_1 _6272_ (.A(net369),
    .B(_2438_),
    .Y(_2439_));
 sg13g2_a22oi_1 _6273_ (.Y(_0141_),
    .B1(_2429_),
    .B2(_2439_),
    .A2(net369),
    .A1(_2664_));
 sg13g2_and2_1 _6274_ (.A(net309),
    .B(net366),
    .X(_0142_));
 sg13g2_and2_1 _6275_ (.A(net452),
    .B(net367),
    .X(_0143_));
 sg13g2_and2_1 _6276_ (.A(net316),
    .B(net367),
    .X(_0144_));
 sg13g2_and2_1 _6277_ (.A(net504),
    .B(net367),
    .X(_0145_));
 sg13g2_and2_1 _6278_ (.A(net456),
    .B(net367),
    .X(_0146_));
 sg13g2_and2_1 _6279_ (.A(net468),
    .B(net366),
    .X(_0147_));
 sg13g2_and2_1 _6280_ (.A(net460),
    .B(net366),
    .X(_0148_));
 sg13g2_and2_1 _6281_ (.A(net482),
    .B(net366),
    .X(_0149_));
 sg13g2_and2_1 _6282_ (.A(net489),
    .B(net366),
    .X(_0150_));
 sg13g2_and2_1 _6283_ (.A(net540),
    .B(net366),
    .X(_0151_));
 sg13g2_and2_1 _6284_ (.A(net516),
    .B(net366),
    .X(_0152_));
 sg13g2_nor2_1 _6285_ (.A(net401),
    .B(_0243_),
    .Y(_0153_));
 sg13g2_nand4_1 _6286_ (.B(\main.demo.vga._q_ycount[6] ),
    .C(_2608_),
    .A(\main.demo.vga._q_ycount[7] ),
    .Y(_2440_),
    .D(\main.demo.vga._q_ycount[4] ));
 sg13g2_nand2_1 _6287_ (.Y(_2441_),
    .A(net469),
    .B(net531));
 sg13g2_nor4_1 _6288_ (.A(net521),
    .B(_2108_),
    .C(_2440_),
    .D(_2441_),
    .Y(_2442_));
 sg13g2_nor2_1 _6289_ (.A(net286),
    .B(net532),
    .Y(_2443_));
 sg13g2_nand3_1 _6290_ (.B(\main.demo.vga._q_ycount[2] ),
    .C(\main.demo.vga._q_ycount[0] ),
    .A(net475),
    .Y(_2444_));
 sg13g2_nor4_1 _6291_ (.A(net465),
    .B(_2440_),
    .C(_2441_),
    .D(_2444_),
    .Y(_2445_));
 sg13g2_nor3_1 _6292_ (.A(net301),
    .B(_2443_),
    .C(_2445_),
    .Y(_0154_));
 sg13g2_nand4_1 _6293_ (.B(\main.demo.vga._q_xcount[9] ),
    .C(\main.demo.vga._q_xcount[8] ),
    .A(\main.demo.vga._q_xcount[6] ),
    .Y(_2446_),
    .D(\main.demo.vga._q_xcount[10] ));
 sg13g2_nor2_1 _6294_ (.A(_2095_),
    .B(_2446_),
    .Y(_2447_));
 sg13g2_a21oi_1 _6295_ (.A1(_3027_),
    .A2(_2447_),
    .Y(_2448_),
    .B1(net278));
 sg13g2_nand3_1 _6296_ (.B(\main.demo.vga._q_xcount[4] ),
    .C(_3025_),
    .A(\main.demo.vga._q_xcount[5] ),
    .Y(_2449_));
 sg13g2_nor3_1 _6297_ (.A(\main.demo.vga._q_xcount[7] ),
    .B(_2446_),
    .C(_2449_),
    .Y(_2450_));
 sg13g2_nor3_1 _6298_ (.A(net301),
    .B(_2448_),
    .C(_2450_),
    .Y(_0155_));
 sg13g2_nor2_1 _6299_ (.A(net400),
    .B(_0235_),
    .Y(_0156_));
 sg13g2_nor2_1 _6300_ (.A(net402),
    .B(net309),
    .Y(_0157_));
 sg13g2_a21oi_1 _6301_ (.A1(net456),
    .A2(_2094_),
    .Y(_2451_),
    .B1(net468));
 sg13g2_nor2_1 _6302_ (.A(_2098_),
    .B(_2451_),
    .Y(_2452_));
 sg13g2_o21ai_1 _6303_ (.B1(net441),
    .Y(_2453_),
    .A1(net374),
    .A2(_2452_));
 sg13g2_inv_1 _6304_ (.Y(_0158_),
    .A(_2453_));
 sg13g2_xor2_1 _6305_ (.B(_2098_),
    .A(net460),
    .X(_2454_));
 sg13g2_o21ai_1 _6306_ (.B1(net440),
    .Y(_2455_),
    .A1(net374),
    .A2(_2454_));
 sg13g2_inv_1 _6307_ (.Y(_0159_),
    .A(_2455_));
 sg13g2_and2_1 _6308_ (.A(net489),
    .B(_2099_),
    .X(_2456_));
 sg13g2_xor2_1 _6309_ (.B(_2099_),
    .A(net489),
    .X(_2457_));
 sg13g2_o21ai_1 _6310_ (.B1(net440),
    .Y(_2458_),
    .A1(net374),
    .A2(_2457_));
 sg13g2_inv_1 _6311_ (.Y(_0160_),
    .A(_2458_));
 sg13g2_nand2_1 _6312_ (.Y(_2459_),
    .A(net540),
    .B(_2456_));
 sg13g2_o21ai_1 _6313_ (.B1(net440),
    .Y(_2460_),
    .A1(net540),
    .A2(_2456_));
 sg13g2_nor2b_1 _6314_ (.A(_2460_),
    .B_N(_2459_),
    .Y(_0161_));
 sg13g2_or2_1 _6315_ (.X(_2461_),
    .B(_2459_),
    .A(net516));
 sg13g2_a21oi_1 _6316_ (.A1(net516),
    .A2(_2459_),
    .Y(_2462_),
    .B1(net374));
 sg13g2_a21oi_1 _6317_ (.A1(_2461_),
    .A2(_2462_),
    .Y(_0162_),
    .B1(net400));
 sg13g2_nand2_1 _6318_ (.Y(_2463_),
    .A(net440),
    .B(_2106_));
 sg13g2_xnor2_1 _6319_ (.Y(_2464_),
    .A(net521),
    .B(net374));
 sg13g2_nor2_1 _6320_ (.A(_2463_),
    .B(_2464_),
    .Y(_0163_));
 sg13g2_a21oi_1 _6321_ (.A1(net521),
    .A2(net374),
    .Y(_2465_),
    .B1(net465));
 sg13g2_nor3_1 _6322_ (.A(net400),
    .B(_2102_),
    .C(_2465_),
    .Y(_0164_));
 sg13g2_xor2_1 _6323_ (.B(net626),
    .A(net513),
    .X(_2466_));
 sg13g2_a21oi_1 _6324_ (.A1(_2106_),
    .A2(_2466_),
    .Y(_0165_),
    .B1(net401));
 sg13g2_a21oi_1 _6325_ (.A1(net513),
    .A2(_2102_),
    .Y(_2467_),
    .B1(net475));
 sg13g2_nor3_1 _6326_ (.A(net400),
    .B(_2103_),
    .C(net514),
    .Y(_0166_));
 sg13g2_xnor2_1 _6327_ (.Y(_2468_),
    .A(net501),
    .B(_2103_));
 sg13g2_a21oi_1 _6328_ (.A1(_2106_),
    .A2(_2468_),
    .Y(_0167_),
    .B1(net400));
 sg13g2_a21oi_1 _6329_ (.A1(\main.demo.vga._q_ycount[4] ),
    .A2(_2103_),
    .Y(_2469_),
    .B1(net319));
 sg13g2_nor3_1 _6330_ (.A(_2104_),
    .B(_2463_),
    .C(net320),
    .Y(_0168_));
 sg13g2_o21ai_1 _6331_ (.B1(net440),
    .Y(_2470_),
    .A1(net458),
    .A2(_2104_));
 sg13g2_nor2_1 _6332_ (.A(_2105_),
    .B(_2470_),
    .Y(_0169_));
 sg13g2_o21ai_1 _6333_ (.B1(net441),
    .Y(_2471_),
    .A1(net548),
    .A2(_2105_));
 sg13g2_a21oi_1 _6334_ (.A1(net548),
    .A2(_2105_),
    .Y(_0170_),
    .B1(_2471_));
 sg13g2_a21o_1 _6335_ (.A2(_2105_),
    .A1(net548),
    .B1(net469),
    .X(_2472_));
 sg13g2_and3_1 _6336_ (.X(_0171_),
    .A(net441),
    .B(net616),
    .C(_2472_));
 sg13g2_nor2_1 _6337_ (.A(net402),
    .B(_1443_),
    .Y(_0172_));
 sg13g2_or2_2 _6338_ (.X(_2473_),
    .B(_1443_),
    .A(net505));
 sg13g2_nand2b_1 _6339_ (.Y(_2474_),
    .B(_2382_),
    .A_N(_2473_));
 sg13g2_nand2_1 _6340_ (.Y(_2475_),
    .A(\main.demo.zic._q_rythm_count[0] ),
    .B(_2211_));
 sg13g2_nand2_1 _6341_ (.Y(_2476_),
    .A(net292),
    .B(net375));
 sg13g2_a21oi_1 _6342_ (.A1(_2475_),
    .A2(_2476_),
    .Y(_0173_),
    .B1(net360));
 sg13g2_a21oi_1 _6343_ (.A1(\main.demo.zic._q_rythm_count[0] ),
    .A2(net375),
    .Y(_2477_),
    .B1(net326));
 sg13g2_and3_1 _6344_ (.X(_2478_),
    .A(net326),
    .B(\main.demo.zic._q_rythm_count[0] ),
    .C(net375));
 sg13g2_nor3_1 _6345_ (.A(net359),
    .B(net327),
    .C(_2478_),
    .Y(_0174_));
 sg13g2_and4_1 _6346_ (.A(\main.demo.zic._q_rythm_count[2] ),
    .B(net326),
    .C(\main.demo.zic._q_rythm_count[0] ),
    .D(net375),
    .X(_2479_));
 sg13g2_nor2_1 _6347_ (.A(net492),
    .B(_2478_),
    .Y(_2480_));
 sg13g2_and2_1 _6348_ (.A(net492),
    .B(_2478_),
    .X(_2481_));
 sg13g2_nor3_1 _6349_ (.A(net360),
    .B(net493),
    .C(_2481_),
    .Y(_0175_));
 sg13g2_nor2_1 _6350_ (.A(net483),
    .B(_2479_),
    .Y(_2482_));
 sg13g2_and2_1 _6351_ (.A(net483),
    .B(_2481_),
    .X(_2483_));
 sg13g2_nor3_1 _6352_ (.A(net360),
    .B(net484),
    .C(_2483_),
    .Y(_0176_));
 sg13g2_and3_1 _6353_ (.X(_2484_),
    .A(net487),
    .B(net483),
    .C(_2479_));
 sg13g2_nor2_1 _6354_ (.A(net487),
    .B(_2483_),
    .Y(_2485_));
 sg13g2_nor3_1 _6355_ (.A(net360),
    .B(_2484_),
    .C(_2485_),
    .Y(_0177_));
 sg13g2_nor2_1 _6356_ (.A(net490),
    .B(_2484_),
    .Y(_2486_));
 sg13g2_and3_1 _6357_ (.X(_2487_),
    .A(net490),
    .B(net487),
    .C(_2483_));
 sg13g2_nor3_1 _6358_ (.A(net360),
    .B(_2486_),
    .C(_2487_),
    .Y(_0178_));
 sg13g2_nor2_1 _6359_ (.A(net323),
    .B(_2487_),
    .Y(_2488_));
 sg13g2_and3_1 _6360_ (.X(_2489_),
    .A(net323),
    .B(\main.demo.zic._q_rythm_count[5] ),
    .C(_2484_));
 sg13g2_nor3_1 _6361_ (.A(net359),
    .B(net324),
    .C(_2489_),
    .Y(_0179_));
 sg13g2_and2_1 _6362_ (.A(net338),
    .B(_2489_),
    .X(_2490_));
 sg13g2_nor2_1 _6363_ (.A(net338),
    .B(_2489_),
    .Y(_2491_));
 sg13g2_nor3_1 _6364_ (.A(net359),
    .B(_2490_),
    .C(net451),
    .Y(_0180_));
 sg13g2_and2_1 _6365_ (.A(net491),
    .B(_2490_),
    .X(_2492_));
 sg13g2_nor2_1 _6366_ (.A(net491),
    .B(_2490_),
    .Y(_2493_));
 sg13g2_nor3_1 _6367_ (.A(net359),
    .B(_2492_),
    .C(_2493_),
    .Y(_0181_));
 sg13g2_nor2_1 _6368_ (.A(net495),
    .B(_2492_),
    .Y(_2494_));
 sg13g2_and2_1 _6369_ (.A(net495),
    .B(_2492_),
    .X(_2495_));
 sg13g2_nor3_1 _6370_ (.A(net359),
    .B(_2494_),
    .C(_2495_),
    .Y(_0182_));
 sg13g2_nor2_1 _6371_ (.A(net334),
    .B(_2495_),
    .Y(_2496_));
 sg13g2_and2_1 _6372_ (.A(net334),
    .B(_2495_),
    .X(_2497_));
 sg13g2_nor3_1 _6373_ (.A(net359),
    .B(net335),
    .C(_2497_),
    .Y(_0183_));
 sg13g2_nor2_1 _6374_ (.A(net461),
    .B(_2497_),
    .Y(_2498_));
 sg13g2_and2_1 _6375_ (.A(net461),
    .B(_2497_),
    .X(_2499_));
 sg13g2_nor3_1 _6376_ (.A(net359),
    .B(_2498_),
    .C(_2499_),
    .Y(_0184_));
 sg13g2_a21oi_1 _6377_ (.A1(net506),
    .A2(_2499_),
    .Y(_2500_),
    .B1(net359));
 sg13g2_o21ai_1 _6378_ (.B1(_2500_),
    .Y(_2501_),
    .A1(net506),
    .A2(_2499_));
 sg13g2_inv_1 _6379_ (.Y(_0185_),
    .A(_2501_));
 sg13g2_and2_1 _6380_ (.A(net437),
    .B(_2402_),
    .X(_0186_));
 sg13g2_nor2_1 _6381_ (.A(net403),
    .B(_2412_),
    .Y(_0187_));
 sg13g2_nor2_1 _6382_ (.A(net403),
    .B(_2400_),
    .Y(_0188_));
 sg13g2_and2_1 _6383_ (.A(net437),
    .B(_2409_),
    .X(_0189_));
 sg13g2_and2_1 _6384_ (.A(net437),
    .B(_2406_),
    .X(_0190_));
 sg13g2_and2_1 _6385_ (.A(net437),
    .B(_2394_),
    .X(_0191_));
 sg13g2_nor2_1 _6386_ (.A(net403),
    .B(net590),
    .Y(_0192_));
 sg13g2_nor2b_1 _6387_ (.A(_0243_),
    .B_N(net521),
    .Y(_0193_));
 sg13g2_nor2b_1 _6388_ (.A(_0243_),
    .B_N(net465),
    .Y(_0194_));
 sg13g2_nor2b_1 _6389_ (.A(_0243_),
    .B_N(net513),
    .Y(_0195_));
 sg13g2_nor2b_1 _6390_ (.A(_0243_),
    .B_N(net475),
    .Y(_0196_));
 sg13g2_and2_1 _6391_ (.A(net501),
    .B(_0240_),
    .X(_0197_));
 sg13g2_nor2_1 _6392_ (.A(_2608_),
    .B(_0243_),
    .Y(_0198_));
 sg13g2_and2_1 _6393_ (.A(net458),
    .B(_0240_),
    .X(_0199_));
 sg13g2_and2_1 _6394_ (.A(net548),
    .B(_0240_),
    .X(_0200_));
 sg13g2_nor2b_1 _6395_ (.A(_0243_),
    .B_N(net469),
    .Y(_0201_));
 sg13g2_and2_1 _6396_ (.A(net485),
    .B(_0240_),
    .X(_0202_));
 sg13g2_nand3b_1 _6397_ (.B(_2401_),
    .C(_2402_),
    .Y(_2502_),
    .A_N(\main.demo.zic._q_idx[1] ));
 sg13g2_a221oi_1 _6398_ (.B2(_2502_),
    .C1(_2406_),
    .B1(_2414_),
    .A1(_2391_),
    .Y(_2503_),
    .A2(_2394_));
 sg13g2_or3_2 _6399_ (.A(_2382_),
    .B(_2421_),
    .C(_2503_),
    .X(_2504_));
 sg13g2_nor3_2 _6400_ (.A(\main.demo.zic._q_squ_env[2] ),
    .B(\main.demo.zic._q_squ_env[1] ),
    .C(\main.demo.zic._q_squ_env[0] ),
    .Y(_2505_));
 sg13g2_nor2b_1 _6401_ (.A(\main.demo.zic._q_squ_env[3] ),
    .B_N(_2505_),
    .Y(_2506_));
 sg13g2_nor2b_1 _6402_ (.A(\main.demo.zic._q_squ_env[4] ),
    .B_N(_2506_),
    .Y(_2507_));
 sg13g2_a21oi_1 _6403_ (.A1(_1428_),
    .A2(_2505_),
    .Y(_2508_),
    .B1(_2381_));
 sg13g2_a21oi_1 _6404_ (.A1(_2606_),
    .A2(_2508_),
    .Y(_2509_),
    .B1(net368));
 sg13g2_a221oi_1 _6405_ (.B2(_2509_),
    .C1(net403),
    .B1(_2504_),
    .A1(_2606_),
    .Y(_0203_),
    .A2(_2386_));
 sg13g2_xnor2_1 _6406_ (.Y(_2510_),
    .A(\main.demo.zic._q_squ_env[1] ),
    .B(\main.demo.zic._q_squ_env[0] ));
 sg13g2_a21oi_1 _6407_ (.A1(_2508_),
    .A2(_2510_),
    .Y(_2511_),
    .B1(net368));
 sg13g2_a221oi_1 _6408_ (.B2(_2511_),
    .C1(net403),
    .B1(_2504_),
    .A1(_2605_),
    .Y(_0204_),
    .A2(net368));
 sg13g2_o21ai_1 _6409_ (.B1(net557),
    .Y(_2512_),
    .A1(\main.demo.zic._q_squ_env[1] ),
    .A2(\main.demo.zic._q_squ_env[0] ));
 sg13g2_nand2b_1 _6410_ (.Y(_2513_),
    .B(_2512_),
    .A_N(_2505_));
 sg13g2_nor2b_2 _6411_ (.A(net368),
    .B_N(_2508_),
    .Y(_2514_));
 sg13g2_a22oi_1 _6412_ (.Y(_2515_),
    .B1(_2513_),
    .B2(_2514_),
    .A2(net368),
    .A1(net557));
 sg13g2_a21oi_1 _6413_ (.A1(_2504_),
    .A2(_2515_),
    .Y(_0205_),
    .B1(net403));
 sg13g2_xor2_1 _6414_ (.B(_2505_),
    .A(\main.demo.zic._q_squ_env[3] ),
    .X(_2516_));
 sg13g2_a22oi_1 _6415_ (.Y(_2517_),
    .B1(_2514_),
    .B2(_2516_),
    .A2(net368),
    .A1(net635));
 sg13g2_a21oi_1 _6416_ (.A1(_2504_),
    .A2(_2517_),
    .Y(_0206_),
    .B1(net401));
 sg13g2_xnor2_1 _6417_ (.Y(_2518_),
    .A(net585),
    .B(_2506_));
 sg13g2_a22oi_1 _6418_ (.Y(_2519_),
    .B1(_2514_),
    .B2(_2518_),
    .A2(net368),
    .A1(\main.demo.zic._q_squ_env[4] ));
 sg13g2_a21oi_1 _6419_ (.A1(_2504_),
    .A2(net586),
    .Y(_0207_),
    .B1(net401));
 sg13g2_xnor2_1 _6420_ (.Y(_2520_),
    .A(_0025_),
    .B(_2507_));
 sg13g2_a22oi_1 _6421_ (.Y(_2521_),
    .B1(_2514_),
    .B2(_2520_),
    .A2(net368),
    .A1(net554));
 sg13g2_a21oi_1 _6422_ (.A1(_2504_),
    .A2(net555),
    .Y(_0208_),
    .B1(net401));
 sg13g2_nor2_1 _6423_ (.A(_2673_),
    .B(net361),
    .Y(_0209_));
 sg13g2_and2_1 _6424_ (.A(\main.demo.zic._q_clock_count[1] ),
    .B(net577),
    .X(_2522_));
 sg13g2_nor3_1 _6425_ (.A(net578),
    .B(_2473_),
    .C(_2522_),
    .Y(_0210_));
 sg13g2_and2_1 _6426_ (.A(net477),
    .B(_2522_),
    .X(_2523_));
 sg13g2_nor2_1 _6427_ (.A(net477),
    .B(_2522_),
    .Y(_2524_));
 sg13g2_nor3_1 _6428_ (.A(net361),
    .B(_2523_),
    .C(net478),
    .Y(_0211_));
 sg13g2_and2_1 _6429_ (.A(net453),
    .B(_2523_),
    .X(_2525_));
 sg13g2_nor2_1 _6430_ (.A(net453),
    .B(_2523_),
    .Y(_2526_));
 sg13g2_nor3_1 _6431_ (.A(net361),
    .B(_2525_),
    .C(net454),
    .Y(_0212_));
 sg13g2_and2_1 _6432_ (.A(net503),
    .B(_2525_),
    .X(_2527_));
 sg13g2_nor2_1 _6433_ (.A(net503),
    .B(_2525_),
    .Y(_2528_));
 sg13g2_nor3_1 _6434_ (.A(net361),
    .B(_2527_),
    .C(_2528_),
    .Y(_0213_));
 sg13g2_and2_1 _6435_ (.A(net471),
    .B(_2527_),
    .X(_2529_));
 sg13g2_nor2_1 _6436_ (.A(net471),
    .B(_2527_),
    .Y(_2530_));
 sg13g2_nor3_1 _6437_ (.A(net361),
    .B(_2529_),
    .C(net472),
    .Y(_0214_));
 sg13g2_xnor2_1 _6438_ (.Y(_2531_),
    .A(net496),
    .B(_2529_));
 sg13g2_nor2_1 _6439_ (.A(net361),
    .B(_2531_),
    .Y(_0215_));
 sg13g2_nor2b_1 _6440_ (.A(net524),
    .B_N(_2529_),
    .Y(_2532_));
 sg13g2_xnor2_1 _6441_ (.Y(_2533_),
    .A(\main.demo.zic._q_clock_count[7] ),
    .B(_2532_));
 sg13g2_nor2_1 _6442_ (.A(net361),
    .B(net525),
    .Y(_0216_));
 sg13g2_nand3_1 _6443_ (.B(net496),
    .C(_2529_),
    .A(\main.demo.zic._q_clock_count[7] ),
    .Y(_2534_));
 sg13g2_xor2_1 _6444_ (.B(_2534_),
    .A(net507),
    .X(_2535_));
 sg13g2_nor2_1 _6445_ (.A(net361),
    .B(net508),
    .Y(_0217_));
 sg13g2_nand2_1 _6446_ (.Y(_2536_),
    .A(_0034_),
    .B(\main.demo.zic._q_idx[4] ));
 sg13g2_nand2_1 _6447_ (.Y(_2537_),
    .A(_2240_),
    .B(_2260_));
 sg13g2_nor2_1 _6448_ (.A(_0034_),
    .B(\main.demo.zic._q_idx[4] ),
    .Y(_2538_));
 sg13g2_nor3_1 _6449_ (.A(\main.demo.zic._q_idx[3] ),
    .B(_2221_),
    .C(_2538_),
    .Y(_2539_));
 sg13g2_a21oi_1 _6450_ (.A1(_2536_),
    .A2(_2537_),
    .Y(_2540_),
    .B1(_2539_));
 sg13g2_inv_1 _6451_ (.Y(_2541_),
    .A(_2540_));
 sg13g2_nor3_1 _6452_ (.A(net408),
    .B(_2218_),
    .C(_2538_),
    .Y(_2542_));
 sg13g2_a21oi_1 _6453_ (.A1(_2215_),
    .A2(_2220_),
    .Y(_2543_),
    .B1(_2246_));
 sg13g2_a22oi_1 _6454_ (.Y(_2544_),
    .B1(_2256_),
    .B2(_2543_),
    .A2(\main.demo.zic._q_idx[4] ),
    .A1(_0034_));
 sg13g2_nor4_2 _6455_ (.A(_2248_),
    .B(_2541_),
    .C(_2542_),
    .Y(_2545_),
    .D(_2544_));
 sg13g2_nand2_1 _6456_ (.Y(_2546_),
    .A(\main.demo.zic._q_tpos[0] ),
    .B(_2545_));
 sg13g2_xor2_1 _6457_ (.B(_2545_),
    .A(net536),
    .X(_2547_));
 sg13g2_nand2_1 _6458_ (.Y(_2548_),
    .A(\main.demo.zic._q_drum_inc[0] ),
    .B(_2547_));
 sg13g2_xnor2_1 _6459_ (.Y(_2549_),
    .A(\main.demo.zic._q_drum_inc[0] ),
    .B(_2547_));
 sg13g2_o21ai_1 _6460_ (.B1(net439),
    .Y(_2550_),
    .A1(net536),
    .A2(net376));
 sg13g2_a21oi_1 _6461_ (.A1(net376),
    .A2(_2549_),
    .Y(_0218_),
    .B1(net537));
 sg13g2_o21ai_1 _6462_ (.B1(_2536_),
    .Y(_2551_),
    .A1(_2231_),
    .A2(_2271_));
 sg13g2_and2_2 _6463_ (.A(_2540_),
    .B(_2551_),
    .X(_2552_));
 sg13g2_inv_1 _6464_ (.Y(_2553_),
    .A(_2552_));
 sg13g2_nor2b_1 _6465_ (.A(_2219_),
    .B_N(_2536_),
    .Y(_2554_));
 sg13g2_nor2_1 _6466_ (.A(_2250_),
    .B(_2538_),
    .Y(_2555_));
 sg13g2_nor4_2 _6467_ (.A(_2235_),
    .B(_2553_),
    .C(_2554_),
    .Y(_2556_),
    .D(_2555_));
 sg13g2_xnor2_1 _6468_ (.Y(_2557_),
    .A(\main.demo.zic._q_tpos[1] ),
    .B(_2556_));
 sg13g2_nor2_1 _6469_ (.A(_2663_),
    .B(_2557_),
    .Y(_2558_));
 sg13g2_xnor2_1 _6470_ (.Y(_2559_),
    .A(_2663_),
    .B(_2557_));
 sg13g2_nand2_1 _6471_ (.Y(_2560_),
    .A(_2546_),
    .B(_2548_));
 sg13g2_nor2b_1 _6472_ (.A(_2559_),
    .B_N(_2560_),
    .Y(_2561_));
 sg13g2_xor2_1 _6473_ (.B(_2560_),
    .A(_2559_),
    .X(_2562_));
 sg13g2_o21ai_1 _6474_ (.B1(net439),
    .Y(_2563_),
    .A1(net518),
    .A2(net377));
 sg13g2_a21oi_1 _6475_ (.A1(net377),
    .A2(_2562_),
    .Y(_0219_),
    .B1(net519));
 sg13g2_a21oi_1 _6476_ (.A1(\main.demo.zic._q_tpos[1] ),
    .A2(_2556_),
    .Y(_2564_),
    .B1(_2558_));
 sg13g2_and2_1 _6477_ (.A(\main.demo.zic._q_tpos[2] ),
    .B(_2552_),
    .X(_2565_));
 sg13g2_xor2_1 _6478_ (.B(_2552_),
    .A(\main.demo.zic._q_tpos[2] ),
    .X(_2566_));
 sg13g2_xnor2_1 _6479_ (.Y(_2567_),
    .A(\main.demo.zic._q_drum_inc[2] ),
    .B(_2566_));
 sg13g2_xor2_1 _6480_ (.B(_2567_),
    .A(_2564_),
    .X(_2568_));
 sg13g2_nand2_1 _6481_ (.Y(_2569_),
    .A(_2561_),
    .B(_2568_));
 sg13g2_xnor2_1 _6482_ (.Y(_2570_),
    .A(_2561_),
    .B(_2568_));
 sg13g2_o21ai_1 _6483_ (.B1(net439),
    .Y(_2571_),
    .A1(net509),
    .A2(net377));
 sg13g2_a21oi_1 _6484_ (.A1(net377),
    .A2(_2570_),
    .Y(_0220_),
    .B1(net510));
 sg13g2_o21ai_1 _6485_ (.B1(_2569_),
    .Y(_2572_),
    .A1(_2564_),
    .A2(_2567_));
 sg13g2_a21oi_1 _6486_ (.A1(\main.demo.zic._q_drum_inc[2] ),
    .A2(_2566_),
    .Y(_2573_),
    .B1(_2565_));
 sg13g2_nor2b_1 _6487_ (.A(_2552_),
    .B_N(\main.demo.zic._q_tpos[3] ),
    .Y(_2574_));
 sg13g2_xnor2_1 _6488_ (.Y(_2575_),
    .A(\main.demo.zic._q_tpos[3] ),
    .B(_2552_));
 sg13g2_xnor2_1 _6489_ (.Y(_2576_),
    .A(\main.demo.zic._q_drum_inc[3] ),
    .B(_2575_));
 sg13g2_nor2_1 _6490_ (.A(_2573_),
    .B(_2576_),
    .Y(_2577_));
 sg13g2_xnor2_1 _6491_ (.Y(_2578_),
    .A(_2573_),
    .B(_2576_));
 sg13g2_nor2b_1 _6492_ (.A(_2578_),
    .B_N(_2572_),
    .Y(_2579_));
 sg13g2_xor2_1 _6493_ (.B(_2578_),
    .A(_2572_),
    .X(_2580_));
 sg13g2_o21ai_1 _6494_ (.B1(net439),
    .Y(_2581_),
    .A1(net534),
    .A2(net377));
 sg13g2_a21oi_1 _6495_ (.A1(net377),
    .A2(_2580_),
    .Y(_0221_),
    .B1(net535));
 sg13g2_a21oi_1 _6496_ (.A1(\main.demo.zic._q_drum_inc[3] ),
    .A2(_2575_),
    .Y(_2582_),
    .B1(_2574_));
 sg13g2_nor2b_1 _6497_ (.A(_2582_),
    .B_N(\main.demo.zic._q_tpos[4] ),
    .Y(_2583_));
 sg13g2_xnor2_1 _6498_ (.Y(_2584_),
    .A(\main.demo.zic._q_tpos[4] ),
    .B(_2582_));
 sg13g2_or3_1 _6499_ (.A(_2577_),
    .B(_2579_),
    .C(_2584_),
    .X(_2585_));
 sg13g2_o21ai_1 _6500_ (.B1(_2584_),
    .Y(_2586_),
    .A1(_2577_),
    .A2(_2579_));
 sg13g2_a21oi_1 _6501_ (.A1(_2585_),
    .A2(_2586_),
    .Y(_2587_),
    .B1(_2211_));
 sg13g2_o21ai_1 _6502_ (.B1(net439),
    .Y(_2588_),
    .A1(net606),
    .A2(net377));
 sg13g2_nor2_1 _6503_ (.A(_2587_),
    .B(_2588_),
    .Y(_0222_));
 sg13g2_nor2b_1 _6504_ (.A(_2583_),
    .B_N(_2586_),
    .Y(_2589_));
 sg13g2_nor3_2 _6505_ (.A(net511),
    .B(_2211_),
    .C(_2589_),
    .Y(_2590_));
 sg13g2_nand3_1 _6506_ (.B(net378),
    .C(_2589_),
    .A(net511),
    .Y(_2591_));
 sg13g2_o21ai_1 _6507_ (.B1(_2591_),
    .Y(_2592_),
    .A1(\main.demo.zic._q_tpos[5] ),
    .A2(net378));
 sg13g2_nor3_1 _6508_ (.A(net401),
    .B(_2590_),
    .C(net512),
    .Y(_0223_));
 sg13g2_o21ai_1 _6509_ (.B1(net440),
    .Y(_2593_),
    .A1(net558),
    .A2(_2590_));
 sg13g2_and2_1 _6510_ (.A(net558),
    .B(_2590_),
    .X(_2594_));
 sg13g2_nor2_1 _6511_ (.A(_2593_),
    .B(_2594_),
    .Y(_0224_));
 sg13g2_nor2_1 _6512_ (.A(net473),
    .B(_2594_),
    .Y(_2595_));
 sg13g2_and2_2 _6513_ (.A(net473),
    .B(_2594_),
    .X(_2596_));
 sg13g2_nor3_1 _6514_ (.A(net400),
    .B(net474),
    .C(_2596_),
    .Y(_0225_));
 sg13g2_o21ai_1 _6515_ (.B1(net441),
    .Y(_2597_),
    .A1(net336),
    .A2(_2596_));
 sg13g2_a21oi_1 _6516_ (.A1(net336),
    .A2(_2596_),
    .Y(_0226_),
    .B1(_2597_));
 sg13g2_a21oi_1 _6517_ (.A1(\main.demo.zic._q_tpos[8] ),
    .A2(_2596_),
    .Y(_2598_),
    .B1(net321));
 sg13g2_nand3_1 _6518_ (.B(net336),
    .C(_2596_),
    .A(net321),
    .Y(_2599_));
 sg13g2_inv_1 _6519_ (.Y(_2600_),
    .A(_2599_));
 sg13g2_nor3_1 _6520_ (.A(net400),
    .B(net322),
    .C(_2600_),
    .Y(_0227_));
 sg13g2_o21ai_1 _6521_ (.B1(net440),
    .Y(_2601_),
    .A1(_2604_),
    .A2(_2599_));
 sg13g2_a21oi_1 _6522_ (.A1(_2604_),
    .A2(_2599_),
    .Y(_0228_),
    .B1(_2601_));
 sg13g2_a21oi_1 _6523_ (.A1(net529),
    .A2(_2600_),
    .Y(_2602_),
    .B1(net530));
 sg13g2_o21ai_1 _6524_ (.B1(net440),
    .Y(_2603_),
    .A1(_1445_),
    .A2(_2599_));
 sg13g2_nor2_1 _6525_ (.A(_2602_),
    .B(_2603_),
    .Y(_0229_));
 sg13g2_xor2_1 _6526_ (.B(_0414_),
    .A(_0358_),
    .X(\main.demo._d___pip_58_1_1___stage___block_3_a[4] ));
 sg13g2_dfrbp_1 _6527_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net18),
    .D(\main.demo._d___pip_58_1_1___stage___block_3_cy[2] ),
    .Q_N(_3150_),
    .Q(\main.demo._q___pip_58_1_2___stage___block_3_cy[2] ));
 sg13g2_dfrbp_1 _6528_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net19),
    .D(\main.demo._d___pip_58_1_1___stage___block_3_cy[3] ),
    .Q_N(_0039_),
    .Q(\main.demo._q___pip_58_1_2___stage___block_3_cy[3] ));
 sg13g2_dfrbp_1 _6529_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net20),
    .D(\main.demo._d___pip_58_1_1___stage___block_3_cy[4] ),
    .Q_N(_0051_),
    .Q(\main.demo._q___pip_58_1_2___stage___block_3_cy[4] ));
 sg13g2_dfrbp_1 _6530_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net21),
    .D(\main.demo._d___pip_58_1_1___stage___block_3_cy[5] ),
    .Q_N(_0050_),
    .Q(\main.demo._q___pip_58_1_2___stage___block_3_cy[5] ));
 sg13g2_dfrbp_1 _6531_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net22),
    .D(\main.demo._d___pip_58_1_1___stage___block_3_cy[6] ),
    .Q_N(_0049_),
    .Q(\main.demo._q___pip_58_1_2___stage___block_3_cy[6] ));
 sg13g2_dfrbp_1 _6532_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net23),
    .D(\main.demo._d___pip_58_1_1___stage___block_3_cy[7] ),
    .Q_N(_0048_),
    .Q(\main.demo._q___pip_58_1_2___stage___block_3_cy[7] ));
 sg13g2_dfrbp_1 _6533_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net24),
    .D(\main.demo._d___pip_58_1_1___stage___block_3_cy[8] ),
    .Q_N(_0047_),
    .Q(\main.demo._q___pip_58_1_2___stage___block_3_cy[8] ));
 sg13g2_dfrbp_1 _6534_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net25),
    .D(\main.demo._d___pip_58_1_1___stage___block_3_cy[9] ),
    .Q_N(_0046_),
    .Q(\main.demo._q___pip_58_1_2___stage___block_3_cy[9] ));
 sg13g2_dfrbp_1 _6535_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net26),
    .D(\main.demo._d___pip_58_1_1___stage___block_3_cy[10] ),
    .Q_N(_0044_),
    .Q(\main.demo._q___pip_58_1_2___stage___block_3_cy[10] ));
 sg13g2_dfrbp_1 _6536_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net27),
    .D(net1),
    .Q_N(_0002_),
    .Q(rst_n_q));
 sg13g2_dfrbp_1 _6537_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net34),
    .D(net356),
    .Q_N(_3151_),
    .Q(_0068_));
 sg13g2_dfrbp_1 _6538_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net17),
    .D(\main.demo._t___pip_58_1_0___stage___block_3_a[7] ),
    .Q_N(_3149_),
    .Q(_0069_));
 sg13g2_dfrbp_1 _6539_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net225),
    .D(_0070_),
    .Q_N(_3148_),
    .Q(\main.demo.vga._q_xcount[1] ));
 sg13g2_dfrbp_1 _6540_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net224),
    .D(_0071_),
    .Q_N(_3147_),
    .Q(\main.demo.vga._q_xcount[2] ));
 sg13g2_dfrbp_1 _6541_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net223),
    .D(_0072_),
    .Q_N(_3146_),
    .Q(\main.demo.vga._q_xcount[3] ));
 sg13g2_dfrbp_1 _6542_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net222),
    .D(_0073_),
    .Q_N(_3145_),
    .Q(\main.demo.vga._q_xcount[4] ));
 sg13g2_dfrbp_1 _6543_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net221),
    .D(_0074_),
    .Q_N(_3144_),
    .Q(\main.demo.vga._q_xcount[7] ));
 sg13g2_dfrbp_1 _6544_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net66),
    .D(net618),
    .Q_N(_3152_),
    .Q(\main.demo.vga._d_vblank ));
 sg13g2_dfrbp_1 _6545_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net220),
    .D(net305),
    .Q_N(_3143_),
    .Q(uio_out[7]));
 sg13g2_dfrbp_1 _6546_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net218),
    .D(net576),
    .Q_N(_3142_),
    .Q(\main.demo._q_speed[0] ));
 sg13g2_dfrbp_1 _6547_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net216),
    .D(_0077_),
    .Q_N(_0016_),
    .Q(\main.demo._q_speed[1] ));
 sg13g2_dfrbp_1 _6548_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net215),
    .D(_0078_),
    .Q_N(_0015_),
    .Q(\main.demo._q_speed[2] ));
 sg13g2_dfrbp_1 _6549_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net214),
    .D(_0079_),
    .Q_N(_0014_),
    .Q(\main.demo._q_speed[3] ));
 sg13g2_dfrbp_1 _6550_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net213),
    .D(net569),
    .Q_N(_0013_),
    .Q(\main.demo._q_speed[4] ));
 sg13g2_dfrbp_1 _6551_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net212),
    .D(_0081_),
    .Q_N(_0007_),
    .Q(\main.demo._q_speed[5] ));
 sg13g2_dfrbp_1 _6552_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net211),
    .D(_0082_),
    .Q_N(_0020_),
    .Q(\main.demo._q_speed[6] ));
 sg13g2_dfrbp_1 _6553_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net210),
    .D(_0083_),
    .Q_N(_3141_),
    .Q(\main.demo._q_speed[7] ));
 sg13g2_dfrbp_1 _6554_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net209),
    .D(_0084_),
    .Q_N(_3140_),
    .Q(\main.demo._q_speed[8] ));
 sg13g2_dfrbp_1 _6555_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net208),
    .D(_0085_),
    .Q_N(_3139_),
    .Q(\main.demo._q_speed[9] ));
 sg13g2_dfrbp_1 _6556_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net207),
    .D(net584),
    .Q_N(_3138_),
    .Q(\main.demo._q_speed[10] ));
 sg13g2_dfrbp_1 _6557_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net206),
    .D(net599),
    .Q_N(_3137_),
    .Q(\main.demo._q_speed[11] ));
 sg13g2_dfrbp_1 _6558_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net205),
    .D(_0088_),
    .Q_N(_3136_),
    .Q(\main.demo._q_speed[12] ));
 sg13g2_dfrbp_1 _6559_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net204),
    .D(_0089_),
    .Q_N(_3135_),
    .Q(\main.demo._q_speed[13] ));
 sg13g2_dfrbp_1 _6560_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net203),
    .D(net572),
    .Q_N(_3134_),
    .Q(\main.demo._q_speed[14] ));
 sg13g2_dfrbp_1 _6561_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net202),
    .D(net499),
    .Q_N(_3133_),
    .Q(\main.demo._q_speed[15] ));
 sg13g2_dfrbp_1 _6562_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net201),
    .D(_0092_),
    .Q_N(_3132_),
    .Q(\main.demo._q_frame[0] ));
 sg13g2_dfrbp_1 _6563_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net200),
    .D(_0093_),
    .Q_N(_3131_),
    .Q(\main.demo._q_frame[1] ));
 sg13g2_dfrbp_1 _6564_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net199),
    .D(_0094_),
    .Q_N(_3130_),
    .Q(\main.demo._q_frame[2] ));
 sg13g2_dfrbp_1 _6565_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net197),
    .D(_0095_),
    .Q_N(_3129_),
    .Q(\main.demo._q_frame[3] ));
 sg13g2_dfrbp_1 _6566_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net196),
    .D(_0096_),
    .Q_N(_3128_),
    .Q(\main.demo._q_frame[4] ));
 sg13g2_dfrbp_1 _6567_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net195),
    .D(_0097_),
    .Q_N(_3127_),
    .Q(\main.demo._q_frame[5] ));
 sg13g2_dfrbp_1 _6568_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net194),
    .D(_0098_),
    .Q_N(_3126_),
    .Q(\main.demo._q_frame[6] ));
 sg13g2_dfrbp_1 _6569_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net193),
    .D(_0099_),
    .Q_N(_3125_),
    .Q(\main.demo._q_frame[7] ));
 sg13g2_dfrbp_1 _6570_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net192),
    .D(_0100_),
    .Q_N(_3124_),
    .Q(\main.demo._q_frame[8] ));
 sg13g2_dfrbp_1 _6571_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net191),
    .D(_0101_),
    .Q_N(_3123_),
    .Q(\main.demo._q_frame[9] ));
 sg13g2_dfrbp_1 _6572_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net190),
    .D(_0102_),
    .Q_N(_3122_),
    .Q(\main.demo._q_frame[10] ));
 sg13g2_dfrbp_1 _6573_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net189),
    .D(_0103_),
    .Q_N(_3121_),
    .Q(\main.demo._q_frame[11] ));
 sg13g2_dfrbp_1 _6574_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net188),
    .D(_0104_),
    .Q_N(_3120_),
    .Q(\main.demo._q_frame[12] ));
 sg13g2_dfrbp_1 _6575_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net187),
    .D(_0105_),
    .Q_N(_3119_),
    .Q(\main.demo._q_frame[13] ));
 sg13g2_dfrbp_1 _6576_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net67),
    .D(_0106_),
    .Q_N(_3153_),
    .Q(\main.demo._q_frame[14] ));
 sg13g2_dfrbp_1 _6577_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net68),
    .D(\main.demo._t___pip_58_1_0___stage___block_3_cy[0] ),
    .Q_N(_3154_),
    .Q(\main.demo._q___pip_58_1_1___stage___block_3_cy[0] ));
 sg13g2_dfrbp_1 _6578_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net69),
    .D(\main.demo._t___pip_58_1_0___stage___block_3_cy[1] ),
    .Q_N(_3155_),
    .Q(\main.demo._q___pip_58_1_1___stage___block_3_cy[1] ));
 sg13g2_dfrbp_1 _6579_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net70),
    .D(\main.demo._t___pip_58_1_0___stage___block_3_cy[2] ),
    .Q_N(_3156_),
    .Q(\main.demo._q___pip_58_1_1___stage___block_3_cy[2] ));
 sg13g2_dfrbp_1 _6580_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net71),
    .D(\main.demo._t___pip_58_1_0___stage___block_3_cy[3] ),
    .Q_N(_3157_),
    .Q(\main.demo._q___pip_58_1_1___stage___block_3_cy[3] ));
 sg13g2_dfrbp_1 _6581_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net72),
    .D(\main.demo._t___pip_58_1_0___stage___block_3_cy[4] ),
    .Q_N(_3158_),
    .Q(\main.demo._q___pip_58_1_1___stage___block_3_cy[4] ));
 sg13g2_dfrbp_1 _6582_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net73),
    .D(\main.demo._t___pip_58_1_0___stage___block_3_cy[5] ),
    .Q_N(_3159_),
    .Q(\main.demo._q___pip_58_1_1___stage___block_3_cy[5] ));
 sg13g2_dfrbp_1 _6583_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net74),
    .D(\main.demo._t___pip_58_1_0___stage___block_3_cy[6] ),
    .Q_N(_3160_),
    .Q(\main.demo._q___pip_58_1_1___stage___block_3_cy[6] ));
 sg13g2_dfrbp_1 _6584_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net75),
    .D(\main.demo._t___pip_58_1_0___stage___block_3_cy[7] ),
    .Q_N(_3161_),
    .Q(\main.demo._q___pip_58_1_1___stage___block_3_cy[7] ));
 sg13g2_dfrbp_1 _6585_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net76),
    .D(\main.demo._t___pip_58_1_0___stage___block_3_cy[8] ),
    .Q_N(_3162_),
    .Q(\main.demo._q___pip_58_1_1___stage___block_3_cy[8] ));
 sg13g2_dfrbp_1 _6586_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net90),
    .D(\main.demo._t___pip_58_1_0___stage___block_3_cy[9] ),
    .Q_N(_3163_),
    .Q(\main.demo._q___pip_58_1_1___stage___block_3_cy[9] ));
 sg13g2_dfrbp_1 _6587_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net186),
    .D(\main.demo._t___pip_58_1_0___stage___block_3_cy[10] ),
    .Q_N(_3118_),
    .Q(\main.demo._q___pip_58_1_1___stage___block_3_cy[10] ));
 sg13g2_dfrbp_1 _6588_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net185),
    .D(_0107_),
    .Q_N(_3117_),
    .Q(\main.demo.zic._q_qpos[0] ));
 sg13g2_dfrbp_1 _6589_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net183),
    .D(net333),
    .Q_N(_0029_),
    .Q(\main.demo.zic._q_qpos[1] ));
 sg13g2_dfrbp_1 _6590_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net175),
    .D(_0109_),
    .Q_N(_3116_),
    .Q(\main.demo.zic._q_qpos[2] ));
 sg13g2_dfrbp_1 _6591_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net173),
    .D(_0110_),
    .Q_N(_0030_),
    .Q(\main.demo.zic._q_qpos[3] ));
 sg13g2_dfrbp_1 _6592_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net171),
    .D(_0111_),
    .Q_N(_3115_),
    .Q(\main.demo.zic._q_qpos[4] ));
 sg13g2_dfrbp_1 _6593_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net159),
    .D(_0112_),
    .Q_N(_0031_),
    .Q(\main.demo.zic._q_qpos[5] ));
 sg13g2_dfrbp_1 _6594_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net157),
    .D(net565),
    .Q_N(_3114_),
    .Q(\main.demo.zic._q_qpos[6] ));
 sg13g2_dfrbp_1 _6595_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net155),
    .D(net331),
    .Q_N(_0032_),
    .Q(\main.demo.zic._q_qpos[7] ));
 sg13g2_dfrbp_1 _6596_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net153),
    .D(net464),
    .Q_N(_3113_),
    .Q(\main.demo.zic._q_qpos[8] ));
 sg13g2_dfrbp_1 _6597_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net151),
    .D(_0116_),
    .Q_N(_3112_),
    .Q(\main.demo.zic._q_qpos[9] ));
 sg13g2_dfrbp_1 _6598_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net149),
    .D(net311),
    .Q_N(_3111_),
    .Q(\main.demo.zic._q_qpos[10] ));
 sg13g2_dfrbp_1 _6599_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net89),
    .D(_0118_),
    .Q_N(_3110_),
    .Q(\main.demo.zic._q_qpos[11] ));
 sg13g2_dfrbp_1 _6600_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net91),
    .D(net481),
    .Q_N(_3164_),
    .Q(\main.demo.zic._q_qpos[12] ));
 sg13g2_dfrbp_1 _6601_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net92),
    .D(net428),
    .Q_N(_3165_),
    .Q(\main.demo._d___pip_58_1_4___stage___block_3_cx[1] ));
 sg13g2_dfrbp_1 _6602_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net93),
    .D(net526),
    .Q_N(_3166_),
    .Q(\main.demo._d___pip_58_1_4___stage___block_3_cx[2] ));
 sg13g2_dfrbp_1 _6603_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net94),
    .D(net562),
    .Q_N(_3167_),
    .Q(\main.demo._d___pip_58_1_4___stage___block_3_cx[3] ));
 sg13g2_dfrbp_1 _6604_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net95),
    .D(net455),
    .Q_N(_3168_),
    .Q(\main.demo._d___pip_58_1_4___stage___block_3_cx[4] ));
 sg13g2_dfrbp_1 _6605_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net96),
    .D(net427),
    .Q_N(_3169_),
    .Q(\main.demo._d___pip_58_1_4___stage___block_3_cx[5] ));
 sg13g2_dfrbp_1 _6606_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net97),
    .D(net300),
    .Q_N(_3170_),
    .Q(\main.demo._d___pip_58_1_4___stage___block_3_cx[6] ));
 sg13g2_dfrbp_1 _6607_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net98),
    .D(net425),
    .Q_N(_3171_),
    .Q(\main.demo._d___pip_58_1_4___stage___block_3_cx[9] ));
 sg13g2_dfrbp_1 _6608_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net99),
    .D(\main.demo._d___pip_58_1_2___stage___block_3_cx[0] ),
    .Q_N(_0012_),
    .Q(\main.demo._d___pip_58_1_3___stage___block_3_cx[0] ));
 sg13g2_dfrbp_1 _6609_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net100),
    .D(\main.demo._d___pip_58_1_2___stage___block_3_cx[1] ),
    .Q_N(_0010_),
    .Q(\main.demo._d___pip_58_1_3___stage___block_3_cx[1] ));
 sg13g2_dfrbp_1 _6610_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net101),
    .D(\main.demo._d___pip_58_1_2___stage___block_3_cx[2] ),
    .Q_N(_0011_),
    .Q(\main.demo._d___pip_58_1_3___stage___block_3_cx[2] ));
 sg13g2_dfrbp_1 _6611_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net102),
    .D(\main.demo._d___pip_58_1_2___stage___block_3_cx[3] ),
    .Q_N(_0008_),
    .Q(\main.demo._d___pip_58_1_3___stage___block_3_cx[3] ));
 sg13g2_dfrbp_1 _6612_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net103),
    .D(\main.demo._d___pip_58_1_2___stage___block_3_cx[4] ),
    .Q_N(_0009_),
    .Q(\main.demo._d___pip_58_1_3___stage___block_3_cx[4] ));
 sg13g2_dfrbp_1 _6613_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net104),
    .D(\main.demo._d___pip_58_1_2___stage___block_3_cx[5] ),
    .Q_N(_3172_),
    .Q(\main.demo._d___pip_58_1_3___stage___block_3_cx[5] ));
 sg13g2_dfrbp_1 _6614_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net105),
    .D(\main.demo._d___pip_58_1_2___stage___block_3_cx[6] ),
    .Q_N(_3173_),
    .Q(\main.demo._d___pip_58_1_3___stage___block_3_cx[6] ));
 sg13g2_dfrbp_1 _6615_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net106),
    .D(\main.demo._d___pip_58_1_2___stage___block_3_cx[7] ),
    .Q_N(_0037_),
    .Q(\main.demo._d___pip_58_1_3___stage___block_3_cx[7] ));
 sg13g2_dfrbp_1 _6616_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net107),
    .D(\main.demo._d___pip_58_1_2___stage___block_3_cx[8] ),
    .Q_N(_0006_),
    .Q(\main.demo._d___pip_58_1_3___stage___block_3_cx[8] ));
 sg13g2_dfrbp_1 _6617_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net108),
    .D(\main.demo._d___pip_58_1_2___stage___block_3_cx[9] ),
    .Q_N(_3174_),
    .Q(\main.demo._d___pip_58_1_3___stage___block_3_cx[9] ));
 sg13g2_dfrbp_1 _6618_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net109),
    .D(\main.demo._d___pip_58_1_2___stage___block_3_cx[10] ),
    .Q_N(_3175_),
    .Q(\main.demo._d___pip_58_1_3___stage___block_3_cx[10] ));
 sg13g2_dfrbp_1 _6619_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net110),
    .D(\main.demo._d___pip_58_1_1___stage___block_3_cx[0] ),
    .Q_N(_3176_),
    .Q(\main.demo._q___pip_58_1_2___stage___block_3_cx[0] ));
 sg13g2_dfrbp_1 _6620_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net111),
    .D(\main.demo._d___pip_58_1_1___stage___block_3_cx[1] ),
    .Q_N(_3177_),
    .Q(\main.demo._q___pip_58_1_2___stage___block_3_cx[1] ));
 sg13g2_dfrbp_1 _6621_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net112),
    .D(\main.demo._d___pip_58_1_1___stage___block_3_cx[2] ),
    .Q_N(_3178_),
    .Q(\main.demo._q___pip_58_1_2___stage___block_3_cx[2] ));
 sg13g2_dfrbp_1 _6622_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net113),
    .D(\main.demo._d___pip_58_1_1___stage___block_3_cx[3] ),
    .Q_N(_3179_),
    .Q(\main.demo._q___pip_58_1_2___stage___block_3_cx[3] ));
 sg13g2_dfrbp_1 _6623_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net114),
    .D(\main.demo._d___pip_58_1_1___stage___block_3_cx[4] ),
    .Q_N(_0042_),
    .Q(\main.demo._q___pip_58_1_2___stage___block_3_cx[4] ));
 sg13g2_dfrbp_1 _6624_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net115),
    .D(\main.demo._d___pip_58_1_1___stage___block_3_cx[5] ),
    .Q_N(_0041_),
    .Q(\main.demo._q___pip_58_1_2___stage___block_3_cx[5] ));
 sg13g2_dfrbp_1 _6625_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net116),
    .D(\main.demo._d___pip_58_1_1___stage___block_3_cx[6] ),
    .Q_N(_0040_),
    .Q(\main.demo._q___pip_58_1_2___stage___block_3_cx[6] ));
 sg13g2_dfrbp_1 _6626_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net117),
    .D(\main.demo._d___pip_58_1_1___stage___block_3_cx[7] ),
    .Q_N(_0038_),
    .Q(\main.demo._q___pip_58_1_2___stage___block_3_cx[7] ));
 sg13g2_dfrbp_1 _6627_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net118),
    .D(\main.demo._d___pip_58_1_1___stage___block_3_cx[8] ),
    .Q_N(_0045_),
    .Q(\main.demo._q___pip_58_1_2___stage___block_3_cx[8] ));
 sg13g2_dfrbp_1 _6628_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net119),
    .D(\main.demo._d___pip_58_1_1___stage___block_3_cx[9] ),
    .Q_N(_0043_),
    .Q(\main.demo._q___pip_58_1_2___stage___block_3_cx[9] ));
 sg13g2_dfrbp_1 _6629_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net120),
    .D(\main.demo._d___pip_58_1_1___stage___block_3_cx[10] ),
    .Q_N(_0052_),
    .Q(\main.demo._q___pip_58_1_2___stage___block_3_cx[10] ));
 sg13g2_dfrbp_1 _6630_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net121),
    .D(net601),
    .Q_N(_3180_),
    .Q(\main.demo._q___pip_58_1_1___stage___block_3_cx[0] ));
 sg13g2_dfrbp_1 _6631_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net122),
    .D(\main.demo._t___pip_58_1_0___stage___block_3_cx[1] ),
    .Q_N(_3181_),
    .Q(\main.demo._q___pip_58_1_1___stage___block_3_cx[1] ));
 sg13g2_dfrbp_1 _6632_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net123),
    .D(net588),
    .Q_N(_3182_),
    .Q(\main.demo._q___pip_58_1_1___stage___block_3_cx[2] ));
 sg13g2_dfrbp_1 _6633_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net124),
    .D(\main.demo._t___pip_58_1_0___stage___block_3_cx[3] ),
    .Q_N(_3183_),
    .Q(\main.demo._q___pip_58_1_1___stage___block_3_cx[3] ));
 sg13g2_dfrbp_1 _6634_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net125),
    .D(\main.demo._t___pip_58_1_0___stage___block_3_cx[4] ),
    .Q_N(_3184_),
    .Q(\main.demo._q___pip_58_1_1___stage___block_3_cx[4] ));
 sg13g2_dfrbp_1 _6635_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net126),
    .D(\main.demo._t___pip_58_1_0___stage___block_3_cx[5] ),
    .Q_N(_3185_),
    .Q(\main.demo._q___pip_58_1_1___stage___block_3_cx[5] ));
 sg13g2_dfrbp_1 _6636_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net127),
    .D(\main.demo._t___pip_58_1_0___stage___block_3_cx[6] ),
    .Q_N(_3186_),
    .Q(\main.demo._q___pip_58_1_1___stage___block_3_cx[6] ));
 sg13g2_dfrbp_1 _6637_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net128),
    .D(\main.demo._t___pip_58_1_0___stage___block_3_cx[7] ),
    .Q_N(_3187_),
    .Q(\main.demo._q___pip_58_1_1___stage___block_3_cx[7] ));
 sg13g2_dfrbp_1 _6638_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net129),
    .D(\main.demo._t___pip_58_1_0___stage___block_3_cx[8] ),
    .Q_N(_3188_),
    .Q(\main.demo._q___pip_58_1_1___stage___block_3_cx[8] ));
 sg13g2_dfrbp_1 _6639_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net130),
    .D(\main.demo._t___pip_58_1_0___stage___block_3_cx[9] ),
    .Q_N(_3189_),
    .Q(\main.demo._q___pip_58_1_1___stage___block_3_cx[9] ));
 sg13g2_dfrbp_1 _6640_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net131),
    .D(\main.demo._t___pip_58_1_0___stage___block_3_cx[10] ),
    .Q_N(_3190_),
    .Q(\main.demo._q___pip_58_1_1___stage___block_3_cx[10] ));
 sg13g2_dfrbp_1 _6641_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net132),
    .D(\main.demo._d___pip_58_1_2___stage___block_3_a[1] ),
    .Q_N(_3191_),
    .Q(\main.demo._d___pip_58_1_3___stage___block_3_a[1] ));
 sg13g2_dfrbp_1 _6642_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net133),
    .D(\main.demo._d___pip_58_1_2___stage___block_3_a[2] ),
    .Q_N(_0019_),
    .Q(\main.demo._d___pip_58_1_3___stage___block_3_a[2] ));
 sg13g2_dfrbp_1 _6643_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net134),
    .D(\main.demo._d___pip_58_1_2___stage___block_3_a[3] ),
    .Q_N(_0018_),
    .Q(\main.demo._d___pip_58_1_3___stage___block_3_a[3] ));
 sg13g2_dfrbp_1 _6644_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net135),
    .D(\main.demo._d___pip_58_1_2___stage___block_3_a[4] ),
    .Q_N(_0017_),
    .Q(\main.demo._d___pip_58_1_3___stage___block_3_a[4] ));
 sg13g2_dfrbp_1 _6645_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net136),
    .D(\main.demo._d___pip_58_1_2___stage___block_3_a[5] ),
    .Q_N(_0022_),
    .Q(\main.demo._d___pip_58_1_3___stage___block_3_a[5] ));
 sg13g2_dfrbp_1 _6646_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net137),
    .D(\main.demo._d___pip_58_1_2___stage___block_3_a[6] ),
    .Q_N(_0021_),
    .Q(\main.demo._d___pip_58_1_3___stage___block_3_a[6] ));
 sg13g2_dfrbp_1 _6647_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net138),
    .D(\main.demo._d___pip_58_1_2___stage___block_3_a[7] ),
    .Q_N(_3192_),
    .Q(\main.demo._d___pip_58_1_3___stage___block_3_a[7] ));
 sg13g2_dfrbp_1 _6648_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net139),
    .D(\main.demo._t___pip_58_1_3___block_87_atten_l[0] ),
    .Q_N(_3193_),
    .Q(\main.demo._d___pip_58_1_4___block_87_atten_l[0] ));
 sg13g2_dfrbp_1 _6649_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net140),
    .D(\main.demo._t___pip_58_1_3___block_87_atten_l[1] ),
    .Q_N(_3194_),
    .Q(\main.demo._d___pip_58_1_4___block_87_atten_l[1] ));
 sg13g2_dfrbp_1 _6650_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net141),
    .D(\main.demo._t___pip_58_1_3___block_87_atten_h[0] ),
    .Q_N(_3195_),
    .Q(\main.demo._d___pip_58_1_4___block_87_atten_h[0] ));
 sg13g2_dfrbp_1 _6651_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net142),
    .D(net552),
    .Q_N(_3196_),
    .Q(\main.demo._d___pip_58_1_4___block_87_atten_h[1] ));
 sg13g2_dfrbp_1 _6652_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net143),
    .D(\main.demo._t___pip_58_1_3___block_87_atten_h[2] ),
    .Q_N(_3197_),
    .Q(\main.demo._d___pip_58_1_4___block_87_atten_h[2] ));
 sg13g2_dfrbp_1 _6653_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net144),
    .D(\main.demo._t___block_68_frag[0] ),
    .Q_N(_3198_),
    .Q(\main.demo._d___pip_58_1_4___block_68_frag[0] ));
 sg13g2_dfrbp_1 _6654_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net145),
    .D(\main.demo._t___block_68_frag[1] ),
    .Q_N(_3199_),
    .Q(\main.demo._d___pip_58_1_4___block_68_frag[1] ));
 sg13g2_dfrbp_1 _6655_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net146),
    .D(\main.demo._t___block_68_frag[2] ),
    .Q_N(_3200_),
    .Q(\main.demo._d___pip_58_1_4___block_68_frag[2] ));
 sg13g2_dfrbp_1 _6656_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net147),
    .D(\main.demo._t___block_68_frag[3] ),
    .Q_N(_3201_),
    .Q(\main.demo._d___pip_58_1_4___block_68_frag[3] ));
 sg13g2_dfrbp_1 _6657_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net160),
    .D(\main.demo._t___block_68_frag[4] ),
    .Q_N(_3202_),
    .Q(\main.demo._d___pip_58_1_4___block_68_frag[4] ));
 sg13g2_dfrbp_1 _6658_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net87),
    .D(\main.demo._t___block_68_frag[5] ),
    .Q_N(_3109_),
    .Q(\main.demo._d___pip_58_1_4___block_68_frag[5] ));
 sg13g2_dfrbp_1 _6659_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net85),
    .D(net298),
    .Q_N(_0000_),
    .Q(\main.demo._q_rot_en ));
 sg13g2_dfrbp_1 _6660_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net83),
    .D(net542),
    .Q_N(_0067_),
    .Q(\main.demo._q_effect[0] ));
 sg13g2_dfrbp_1 _6661_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net81),
    .D(_0122_),
    .Q_N(_3108_),
    .Q(\main.demo._q_effect[1] ));
 sg13g2_dfrbp_1 _6662_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net79),
    .D(net291),
    .Q_N(_0066_),
    .Q(\main.demo._q_th[0] ));
 sg13g2_dfrbp_1 _6663_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net77),
    .D(net308),
    .Q_N(_3107_),
    .Q(\main.demo._q_th[1] ));
 sg13g2_dfrbp_1 _6664_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net64),
    .D(_0125_),
    .Q_N(_3106_),
    .Q(\main.demo._q_th[2] ));
 sg13g2_dfrbp_1 _6665_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net62),
    .D(_0126_),
    .Q_N(_3105_),
    .Q(\main.demo._q_th[3] ));
 sg13g2_dfrbp_1 _6666_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net60),
    .D(_0127_),
    .Q_N(_3104_),
    .Q(\main.demo._q_th[4] ));
 sg13g2_dfrbp_1 _6667_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net58),
    .D(_0128_),
    .Q_N(_3103_),
    .Q(\main.demo._q_th[5] ));
 sg13g2_dfrbp_1 _6668_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net56),
    .D(_0129_),
    .Q_N(_0023_),
    .Q(\main.demo._q_th[6] ));
 sg13g2_dfrbp_1 _6669_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net54),
    .D(_0130_),
    .Q_N(_3102_),
    .Q(\main.demo._q_th[7] ));
 sg13g2_dfrbp_1 _6670_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net161),
    .D(net315),
    .Q_N(_3203_),
    .Q(\main.demo._q_th[8] ));
 sg13g2_dfrbp_1 _6671_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net162),
    .D(\main.demo._d_prev_b[0] ),
    .Q_N(_3204_),
    .Q(\main.demo._d_prev_b[2] ));
 sg13g2_dfrbp_1 _6672_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net163),
    .D(\main.demo._d_prev_b[1] ),
    .Q_N(_3205_),
    .Q(\main.demo._d_prev_b[3] ));
 sg13g2_dfrbp_1 _6673_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net164),
    .D(net282),
    .Q_N(_3206_),
    .Q(\main.demo._d_prev_b[4] ));
 sg13g2_dfrbp_1 _6674_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net165),
    .D(net285),
    .Q_N(_3207_),
    .Q(\main.demo._d_prev_b[5] ));
 sg13g2_dfrbp_1 _6675_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net166),
    .D(net279),
    .Q_N(_3208_),
    .Q(\main.demo._d_prev_b[6] ));
 sg13g2_dfrbp_1 _6676_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net167),
    .D(net281),
    .Q_N(_3209_),
    .Q(\main.demo._d_prev_b[7] ));
 sg13g2_dfrbp_1 _6677_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net168),
    .D(net280),
    .Q_N(_3210_),
    .Q(\main.demo._q_prev_b[6] ));
 sg13g2_dfrbp_1 _6678_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net169),
    .D(net283),
    .Q_N(_3211_),
    .Q(\main.demo._q_prev_b[7] ));
 sg13g2_dfrbp_1 _6679_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net176),
    .D(net286),
    .Q_N(_3212_),
    .Q(\main.demo._q_prev_vs ));
 sg13g2_dfrbp_1 _6680_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net52),
    .D(net278),
    .Q_N(_3101_),
    .Q(uo_out[7]));
 sg13g2_dfrbp_1 _6681_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net50),
    .D(_0132_),
    .Q_N(_3100_),
    .Q(uo_out[0]));
 sg13g2_dfrbp_1 _6682_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net49),
    .D(_0133_),
    .Q_N(_3099_),
    .Q(uo_out[1]));
 sg13g2_dfrbp_1 _6683_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net48),
    .D(_0134_),
    .Q_N(_3098_),
    .Q(uo_out[2]));
 sg13g2_dfrbp_1 _6684_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net47),
    .D(_0135_),
    .Q_N(_3097_),
    .Q(uo_out[4]));
 sg13g2_dfrbp_1 _6685_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net46),
    .D(_0136_),
    .Q_N(_3096_),
    .Q(uo_out[5]));
 sg13g2_dfrbp_1 _6686_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net177),
    .D(_0137_),
    .Q_N(_3213_),
    .Q(uo_out[6]));
 sg13g2_dfrbp_1 _6687_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net178),
    .D(net340),
    .Q_N(_3214_),
    .Q(\main.demo._q___pip_58_1_2___stage___block_3_a[1] ));
 sg13g2_dfrbp_1 _6688_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net179),
    .D(net344),
    .Q_N(_3215_),
    .Q(\main.demo._q___pip_58_1_2___stage___block_3_a[2] ));
 sg13g2_dfrbp_1 _6689_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net180),
    .D(net348),
    .Q_N(_3216_),
    .Q(\main.demo._q___pip_58_1_2___stage___block_3_a[3] ));
 sg13g2_dfrbp_1 _6690_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net181),
    .D(\main.demo._d___pip_58_1_1___stage___block_3_a[4] ),
    .Q_N(_3217_),
    .Q(\main.demo._q___pip_58_1_2___stage___block_3_a[4] ));
 sg13g2_dfrbp_1 _6691_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net198),
    .D(net295),
    .Q_N(_3218_),
    .Q(\main.demo._q___pip_58_1_2___stage___block_3_a[6] ));
 sg13g2_dfrbp_1 _6692_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net45),
    .D(net288),
    .Q_N(_3095_),
    .Q(\main.demo._q___pip_58_1_2___stage___block_3_a[7] ));
 sg13g2_dfrbp_1 _6693_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net44),
    .D(_0138_),
    .Q_N(_3094_),
    .Q(\main.demo.zic._q_drum_inc[0] ));
 sg13g2_dfrbp_1 _6694_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net43),
    .D(_0139_),
    .Q_N(_3093_),
    .Q(\main.demo.zic._q_drum_inc[1] ));
 sg13g2_dfrbp_1 _6695_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net42),
    .D(_0140_),
    .Q_N(_3092_),
    .Q(\main.demo.zic._q_drum_inc[2] ));
 sg13g2_dfrbp_1 _6696_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net41),
    .D(_0141_),
    .Q_N(_3091_),
    .Q(\main.demo.zic._q_drum_inc[3] ));
 sg13g2_dfrbp_1 _6697_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net40),
    .D(_0142_),
    .Q_N(_0004_),
    .Q(\main.demo._t___stage___block_3_x[0] ));
 sg13g2_dfrbp_1 _6698_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net39),
    .D(_0143_),
    .Q_N(_0005_),
    .Q(\main.demo._t___stage___block_3_x[1] ));
 sg13g2_dfrbp_1 _6699_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net38),
    .D(_0144_),
    .Q_N(_3090_),
    .Q(\main.demo._t___stage___block_3_x[2] ));
 sg13g2_dfrbp_1 _6700_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net37),
    .D(_0145_),
    .Q_N(_0059_),
    .Q(\main.demo._w_vga_vga_x[3] ));
 sg13g2_dfrbp_1 _6701_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net36),
    .D(_0146_),
    .Q_N(_0058_),
    .Q(\main.demo._w_vga_vga_x[4] ));
 sg13g2_dfrbp_1 _6702_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net35),
    .D(_0147_),
    .Q_N(_0057_),
    .Q(\main.demo._w_vga_vga_x[5] ));
 sg13g2_dfrbp_1 _6703_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net33),
    .D(_0148_),
    .Q_N(_0056_),
    .Q(\main.demo._w_vga_vga_x[6] ));
 sg13g2_dfrbp_1 _6704_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net32),
    .D(_0149_),
    .Q_N(_0055_),
    .Q(\main.demo._w_vga_vga_x[7] ));
 sg13g2_dfrbp_1 _6705_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net31),
    .D(_0150_),
    .Q_N(_0054_),
    .Q(\main.demo._w_vga_vga_x[8] ));
 sg13g2_dfrbp_1 _6706_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net30),
    .D(_0151_),
    .Q_N(_0053_),
    .Q(\main.demo._w_vga_vga_x[9] ));
 sg13g2_dfrbp_1 _6707_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net29),
    .D(_0152_),
    .Q_N(_3089_),
    .Q(\main.demo._w_vga_vga_x[10] ));
 sg13g2_dfrbp_1 _6708_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net275),
    .D(_0153_),
    .Q_N(_3219_),
    .Q(\main.demo.vga._q_active_v ));
 sg13g2_dfrbp_1 _6709_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net28),
    .D(\main.demo.vga._d_active ),
    .Q_N(_3088_),
    .Q(\main.demo._w_vga_active ));
 sg13g2_dfrbp_1 _6710_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net16),
    .D(net533),
    .Q_N(_3087_),
    .Q(\main._w_demo_video_vs ));
 sg13g2_dfrbp_1 _6711_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net273),
    .D(net302),
    .Q_N(_3086_),
    .Q(\main._w_demo_video_hs ));
 sg13g2_dfrbp_1 _6712_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net271),
    .D(_0156_),
    .Q_N(_3085_),
    .Q(\main.demo.vga._q_active_h ));
 sg13g2_dfrbp_1 _6713_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net270),
    .D(_0157_),
    .Q_N(_3084_),
    .Q(\main.demo.vga._q_xcount[0] ));
 sg13g2_dfrbp_1 _6714_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net269),
    .D(_0158_),
    .Q_N(_3083_),
    .Q(\main.demo.vga._q_xcount[5] ));
 sg13g2_dfrbp_1 _6715_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net268),
    .D(_0159_),
    .Q_N(_3082_),
    .Q(\main.demo.vga._q_xcount[6] ));
 sg13g2_dfrbp_1 _6716_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net267),
    .D(_0160_),
    .Q_N(_3081_),
    .Q(\main.demo.vga._q_xcount[8] ));
 sg13g2_dfrbp_1 _6717_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net266),
    .D(_0161_),
    .Q_N(_3080_),
    .Q(\main.demo.vga._q_xcount[9] ));
 sg13g2_dfrbp_1 _6718_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net265),
    .D(_0162_),
    .Q_N(_3079_),
    .Q(\main.demo.vga._q_xcount[10] ));
 sg13g2_dfrbp_1 _6719_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net264),
    .D(_0163_),
    .Q_N(_3078_),
    .Q(\main.demo.vga._q_ycount[0] ));
 sg13g2_dfrbp_1 _6720_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net262),
    .D(net522),
    .Q_N(_3077_),
    .Q(\main.demo.vga._q_ycount[1] ));
 sg13g2_dfrbp_1 _6721_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net260),
    .D(_0165_),
    .Q_N(_3076_),
    .Q(\main.demo.vga._q_ycount[2] ));
 sg13g2_dfrbp_1 _6722_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net258),
    .D(net515),
    .Q_N(_3075_),
    .Q(\main.demo.vga._q_ycount[3] ));
 sg13g2_dfrbp_1 _6723_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net256),
    .D(_0167_),
    .Q_N(_3074_),
    .Q(\main.demo.vga._q_ycount[4] ));
 sg13g2_dfrbp_1 _6724_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net254),
    .D(_0168_),
    .Q_N(_3073_),
    .Q(\main.demo.vga._q_ycount[5] ));
 sg13g2_dfrbp_1 _6725_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net252),
    .D(_0169_),
    .Q_N(_3072_),
    .Q(\main.demo.vga._q_ycount[6] ));
 sg13g2_dfrbp_1 _6726_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net250),
    .D(_0170_),
    .Q_N(_3071_),
    .Q(\main.demo.vga._q_ycount[7] ));
 sg13g2_dfrbp_1 _6727_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net248),
    .D(_0171_),
    .Q_N(_3070_),
    .Q(\main.demo.vga._q_ycount[8] ));
 sg13g2_dfrbp_1 _6728_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net246),
    .D(_0172_),
    .Q_N(_3069_),
    .Q(\main.demo._q_go ));
 sg13g2_dfrbp_1 _6729_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net245),
    .D(net293),
    .Q_N(_0065_),
    .Q(\main.demo.zic._q_rythm_count[0] ));
 sg13g2_dfrbp_1 _6730_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net243),
    .D(net328),
    .Q_N(_3068_),
    .Q(\main.demo.zic._q_rythm_count[1] ));
 sg13g2_dfrbp_1 _6731_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net241),
    .D(_0175_),
    .Q_N(_3067_),
    .Q(\main.demo.zic._q_rythm_count[2] ));
 sg13g2_dfrbp_1 _6732_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net239),
    .D(_0176_),
    .Q_N(_3066_),
    .Q(\main.demo.zic._q_rythm_count[3] ));
 sg13g2_dfrbp_1 _6733_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net237),
    .D(_0177_),
    .Q_N(_3065_),
    .Q(\main.demo.zic._q_rythm_count[4] ));
 sg13g2_dfrbp_1 _6734_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net235),
    .D(_0178_),
    .Q_N(_3064_),
    .Q(\main.demo.zic._q_rythm_count[5] ));
 sg13g2_dfrbp_1 _6735_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net233),
    .D(net325),
    .Q_N(_3063_),
    .Q(\main.demo.zic._q_rythm_count[6] ));
 sg13g2_dfrbp_1 _6736_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net231),
    .D(_0180_),
    .Q_N(_3062_),
    .Q(\main.demo.zic._q_rythm_count[7] ));
 sg13g2_dfrbp_1 _6737_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net229),
    .D(_0181_),
    .Q_N(_3061_),
    .Q(\main.demo.zic._q_rythm_count[8] ));
 sg13g2_dfrbp_1 _6738_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net227),
    .D(_0182_),
    .Q_N(_3060_),
    .Q(\main.demo.zic._q_rythm_count[9] ));
 sg13g2_dfrbp_1 _6739_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net219),
    .D(_0183_),
    .Q_N(_3059_),
    .Q(\main.demo.zic._q_rythm_count[10] ));
 sg13g2_dfrbp_1 _6740_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net184),
    .D(_0184_),
    .Q_N(_3058_),
    .Q(\main.demo.zic._q_rythm_count[11] ));
 sg13g2_dfrbp_1 _6741_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net174),
    .D(_0185_),
    .Q_N(_3057_),
    .Q(\main.demo.zic._q_rythm_count[12] ));
 sg13g2_dfrbp_1 _6742_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net170),
    .D(_0186_),
    .Q_N(_3056_),
    .Q(\main.demo.zic._q_idx[0] ));
 sg13g2_dfrbp_1 _6743_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net158),
    .D(_0187_),
    .Q_N(_3055_),
    .Q(\main.demo.zic._q_idx[1] ));
 sg13g2_dfrbp_1 _6744_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net156),
    .D(_0188_),
    .Q_N(_3054_),
    .Q(\main.demo.zic._q_idx[2] ));
 sg13g2_dfrbp_1 _6745_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net154),
    .D(_0189_),
    .Q_N(_3053_),
    .Q(\main.demo.zic._q_idx[3] ));
 sg13g2_dfrbp_1 _6746_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net152),
    .D(_0190_),
    .Q_N(_0034_),
    .Q(\main.demo.zic._q_idx[4] ));
 sg13g2_dfrbp_1 _6747_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net150),
    .D(_0191_),
    .Q_N(_0036_),
    .Q(\main.demo.zic._q_idx[5] ));
 sg13g2_dfrbp_1 _6748_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net148),
    .D(_0192_),
    .Q_N(_0035_),
    .Q(\main.demo.zic._q_idx[6] ));
 sg13g2_dfrbp_1 _6749_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net88),
    .D(_0193_),
    .Q_N(_3052_),
    .Q(\main.demo._t___stage___block_3_y[0] ));
 sg13g2_dfrbp_1 _6750_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net86),
    .D(net466),
    .Q_N(_3051_),
    .Q(\main.demo._t___stage___block_3_y[1] ));
 sg13g2_dfrbp_1 _6751_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net84),
    .D(_0195_),
    .Q_N(_0003_),
    .Q(\main.demo._t___stage___block_3_y[2] ));
 sg13g2_dfrbp_1 _6752_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net82),
    .D(net476),
    .Q_N(_0001_),
    .Q(\main.demo._w_vga_vga_y[3] ));
 sg13g2_dfrbp_1 _6753_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net80),
    .D(net502),
    .Q_N(_3050_),
    .Q(\main.demo._w_vga_vga_y[4] ));
 sg13g2_dfrbp_1 _6754_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net78),
    .D(_0198_),
    .Q_N(_0063_),
    .Q(\main.demo._w_vga_vga_y[5] ));
 sg13g2_dfrbp_1 _6755_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net65),
    .D(net459),
    .Q_N(_0062_),
    .Q(\main.demo._w_vga_vga_y[6] ));
 sg13g2_dfrbp_1 _6756_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net63),
    .D(net549),
    .Q_N(_0061_),
    .Q(\main.demo._w_vga_vga_y[7] ));
 sg13g2_dfrbp_1 _6757_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net61),
    .D(net470),
    .Q_N(_3049_),
    .Q(\main.demo._w_vga_vga_y[8] ));
 sg13g2_dfrbp_1 _6758_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net59),
    .D(net486),
    .Q_N(_0060_),
    .Q(\main.demo._w_vga_vga_y[10] ));
 sg13g2_dfrbp_1 _6759_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net57),
    .D(_0203_),
    .Q_N(_3048_),
    .Q(\main.demo.zic._q_squ_env[0] ));
 sg13g2_dfrbp_1 _6760_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net53),
    .D(net544),
    .Q_N(_3047_),
    .Q(\main.demo.zic._q_squ_env[1] ));
 sg13g2_dfrbp_1 _6761_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net274),
    .D(_0205_),
    .Q_N(_3046_),
    .Q(\main.demo.zic._q_squ_env[2] ));
 sg13g2_dfrbp_1 _6762_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net263),
    .D(_0206_),
    .Q_N(_3045_),
    .Q(\main.demo.zic._q_squ_env[3] ));
 sg13g2_dfrbp_1 _6763_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net259),
    .D(_0207_),
    .Q_N(_0024_),
    .Q(\main.demo.zic._q_squ_env[4] ));
 sg13g2_dfrbp_1 _6764_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net255),
    .D(_0208_),
    .Q_N(_0025_),
    .Q(\main.demo.zic._q_squ_env[5] ));
 sg13g2_dfrbp_1 _6765_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net251),
    .D(_0209_),
    .Q_N(_0064_),
    .Q(\main.demo.zic._q_clock_count[0] ));
 sg13g2_dfrbp_1 _6766_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net249),
    .D(net579),
    .Q_N(_3044_),
    .Q(\main.demo.zic._q_clock_count[1] ));
 sg13g2_dfrbp_1 _6767_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net247),
    .D(_0211_),
    .Q_N(_3043_),
    .Q(\main.demo.zic._q_clock_count[2] ));
 sg13g2_dfrbp_1 _6768_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net244),
    .D(_0212_),
    .Q_N(_0028_),
    .Q(\main.demo.zic._q_clock_count[3] ));
 sg13g2_dfrbp_1 _6769_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net242),
    .D(_0213_),
    .Q_N(_3042_),
    .Q(\main.demo.zic._q_clock_count[4] ));
 sg13g2_dfrbp_1 _6770_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net240),
    .D(_0214_),
    .Q_N(_0027_),
    .Q(\main.demo.zic._q_clock_count[5] ));
 sg13g2_dfrbp_1 _6771_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net238),
    .D(_0215_),
    .Q_N(_0026_),
    .Q(\main.demo.zic._q_clock_count[6] ));
 sg13g2_dfrbp_1 _6772_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net236),
    .D(_0216_),
    .Q_N(_3041_),
    .Q(\main.demo.zic._q_clock_count[7] ));
 sg13g2_dfrbp_1 _6773_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net234),
    .D(_0217_),
    .Q_N(_3040_),
    .Q(\main.demo.zic._q_clock_count[8] ));
 sg13g2_dfrbp_1 _6774_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net232),
    .D(net538),
    .Q_N(_3039_),
    .Q(\main.demo.zic._q_tpos[0] ));
 sg13g2_dfrbp_1 _6775_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net228),
    .D(net520),
    .Q_N(_3038_),
    .Q(\main.demo.zic._q_tpos[1] ));
 sg13g2_dfrbp_1 _6776_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net217),
    .D(_0220_),
    .Q_N(_3037_),
    .Q(\main.demo.zic._q_tpos[2] ));
 sg13g2_dfrbp_1 _6777_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net172),
    .D(_0221_),
    .Q_N(_3036_),
    .Q(\main.demo.zic._q_tpos[3] ));
 sg13g2_dfrbp_1 _6778_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net51),
    .D(_0222_),
    .Q_N(_3035_),
    .Q(\main.demo.zic._q_tpos[4] ));
 sg13g2_dfrbp_1 _6779_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net261),
    .D(_0223_),
    .Q_N(_0033_),
    .Q(\main.demo.zic._q_tpos[5] ));
 sg13g2_dfrbp_1 _6780_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net253),
    .D(_0224_),
    .Q_N(_3034_),
    .Q(\main.demo.zic._q_tpos[6] ));
 sg13g2_dfrbp_1 _6781_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net226),
    .D(_0225_),
    .Q_N(_3033_),
    .Q(\main.demo.zic._q_tpos[7] ));
 sg13g2_dfrbp_1 _6782_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net55),
    .D(net337),
    .Q_N(_3032_),
    .Q(\main.demo.zic._q_tpos[8] ));
 sg13g2_dfrbp_1 _6783_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net257),
    .D(_0227_),
    .Q_N(_3031_),
    .Q(\main.demo.zic._q_tpos[9] ));
 sg13g2_dfrbp_1 _6784_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net182),
    .D(_0228_),
    .Q_N(_3030_),
    .Q(\main.demo.zic._q_tpos[10] ));
 sg13g2_dfrbp_1 _6785_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net276),
    .D(_0229_),
    .Q_N(_3220_),
    .Q(\main.demo.zic._q_tpos[11] ));
 sg13g2_dfrbp_1 _6786_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net272),
    .D(\main.demo._d___pip_58_1_1___stage___block_3_cy[0] ),
    .Q_N(_3221_),
    .Q(\main.demo._q___pip_58_1_2___stage___block_3_cy[0] ));
 sg13g2_dfrbp_1 _6787_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net230),
    .D(\main.demo._d___pip_58_1_1___stage___block_3_cy[1] ),
    .Q_N(_3029_),
    .Q(\main.demo._q___pip_58_1_2___stage___block_3_cy[1] ));
 sg13g2_tiehi _6538__17 (.L_HI(net17));
 sg13g2_tiehi _6527__18 (.L_HI(net18));
 sg13g2_tiehi _6528__19 (.L_HI(net19));
 sg13g2_tiehi _6529__20 (.L_HI(net20));
 sg13g2_tiehi _6530__21 (.L_HI(net21));
 sg13g2_tiehi _6531__22 (.L_HI(net22));
 sg13g2_tiehi _6532__23 (.L_HI(net23));
 sg13g2_tiehi _6533__24 (.L_HI(net24));
 sg13g2_tiehi _6534__25 (.L_HI(net25));
 sg13g2_tiehi _6535__26 (.L_HI(net26));
 sg13g2_tiehi _6536__27 (.L_HI(net27));
 sg13g2_tiehi _6709__28 (.L_HI(net28));
 sg13g2_tiehi _6707__29 (.L_HI(net29));
 sg13g2_tiehi _6706__30 (.L_HI(net30));
 sg13g2_tiehi _6705__31 (.L_HI(net31));
 sg13g2_tiehi _6704__32 (.L_HI(net32));
 sg13g2_tiehi _6703__33 (.L_HI(net33));
 sg13g2_tiehi _6537__34 (.L_HI(net34));
 sg13g2_tiehi _6702__35 (.L_HI(net35));
 sg13g2_tiehi _6701__36 (.L_HI(net36));
 sg13g2_tiehi _6700__37 (.L_HI(net37));
 sg13g2_tiehi _6699__38 (.L_HI(net38));
 sg13g2_tiehi _6698__39 (.L_HI(net39));
 sg13g2_tiehi _6697__40 (.L_HI(net40));
 sg13g2_tiehi _6696__41 (.L_HI(net41));
 sg13g2_tiehi _6695__42 (.L_HI(net42));
 sg13g2_tiehi _6694__43 (.L_HI(net43));
 sg13g2_tiehi _6693__44 (.L_HI(net44));
 sg13g2_tiehi _6692__45 (.L_HI(net45));
 sg13g2_tiehi _6685__46 (.L_HI(net46));
 sg13g2_tiehi _6684__47 (.L_HI(net47));
 sg13g2_tiehi _6683__48 (.L_HI(net48));
 sg13g2_tiehi _6682__49 (.L_HI(net49));
 sg13g2_tiehi _6681__50 (.L_HI(net50));
 sg13g2_tiehi _6778__51 (.L_HI(net51));
 sg13g2_tiehi _6680__52 (.L_HI(net52));
 sg13g2_tiehi _6760__53 (.L_HI(net53));
 sg13g2_tiehi _6669__54 (.L_HI(net54));
 sg13g2_tiehi _6782__55 (.L_HI(net55));
 sg13g2_tiehi _6668__56 (.L_HI(net56));
 sg13g2_tiehi _6759__57 (.L_HI(net57));
 sg13g2_tiehi _6667__58 (.L_HI(net58));
 sg13g2_tiehi _6758__59 (.L_HI(net59));
 sg13g2_tiehi _6666__60 (.L_HI(net60));
 sg13g2_tiehi _6757__61 (.L_HI(net61));
 sg13g2_tiehi _6665__62 (.L_HI(net62));
 sg13g2_tiehi _6756__63 (.L_HI(net63));
 sg13g2_tiehi _6664__64 (.L_HI(net64));
 sg13g2_tiehi _6755__65 (.L_HI(net65));
 sg13g2_tiehi _6544__66 (.L_HI(net66));
 sg13g2_tiehi _6576__67 (.L_HI(net67));
 sg13g2_tiehi _6577__68 (.L_HI(net68));
 sg13g2_tiehi _6578__69 (.L_HI(net69));
 sg13g2_tiehi _6579__70 (.L_HI(net70));
 sg13g2_tiehi _6580__71 (.L_HI(net71));
 sg13g2_tiehi _6581__72 (.L_HI(net72));
 sg13g2_tiehi _6582__73 (.L_HI(net73));
 sg13g2_tiehi _6583__74 (.L_HI(net74));
 sg13g2_tiehi _6584__75 (.L_HI(net75));
 sg13g2_tiehi _6585__76 (.L_HI(net76));
 sg13g2_tiehi _6663__77 (.L_HI(net77));
 sg13g2_tiehi _6754__78 (.L_HI(net78));
 sg13g2_tiehi _6662__79 (.L_HI(net79));
 sg13g2_tiehi _6753__80 (.L_HI(net80));
 sg13g2_tiehi _6661__81 (.L_HI(net81));
 sg13g2_tiehi _6752__82 (.L_HI(net82));
 sg13g2_tiehi _6660__83 (.L_HI(net83));
 sg13g2_tiehi _6751__84 (.L_HI(net84));
 sg13g2_tiehi _6659__85 (.L_HI(net85));
 sg13g2_tiehi _6750__86 (.L_HI(net86));
 sg13g2_tiehi _6658__87 (.L_HI(net87));
 sg13g2_tiehi _6749__88 (.L_HI(net88));
 sg13g2_tiehi _6599__89 (.L_HI(net89));
 sg13g2_tiehi _6586__90 (.L_HI(net90));
 sg13g2_tiehi _6600__91 (.L_HI(net91));
 sg13g2_tiehi _6601__92 (.L_HI(net92));
 sg13g2_tiehi _6602__93 (.L_HI(net93));
 sg13g2_tiehi _6603__94 (.L_HI(net94));
 sg13g2_tiehi _6604__95 (.L_HI(net95));
 sg13g2_tiehi _6605__96 (.L_HI(net96));
 sg13g2_tiehi _6606__97 (.L_HI(net97));
 sg13g2_tiehi _6607__98 (.L_HI(net98));
 sg13g2_tiehi _6608__99 (.L_HI(net99));
 sg13g2_tiehi _6609__100 (.L_HI(net100));
 sg13g2_tiehi _6610__101 (.L_HI(net101));
 sg13g2_tiehi _6611__102 (.L_HI(net102));
 sg13g2_tiehi _6612__103 (.L_HI(net103));
 sg13g2_tiehi _6613__104 (.L_HI(net104));
 sg13g2_tiehi _6614__105 (.L_HI(net105));
 sg13g2_tiehi _6615__106 (.L_HI(net106));
 sg13g2_tiehi _6616__107 (.L_HI(net107));
 sg13g2_tiehi _6617__108 (.L_HI(net108));
 sg13g2_tiehi _6618__109 (.L_HI(net109));
 sg13g2_tiehi _6619__110 (.L_HI(net110));
 sg13g2_tiehi _6620__111 (.L_HI(net111));
 sg13g2_tiehi _6621__112 (.L_HI(net112));
 sg13g2_tiehi _6622__113 (.L_HI(net113));
 sg13g2_tiehi _6623__114 (.L_HI(net114));
 sg13g2_tiehi _6624__115 (.L_HI(net115));
 sg13g2_tiehi _6625__116 (.L_HI(net116));
 sg13g2_tiehi _6626__117 (.L_HI(net117));
 sg13g2_tiehi _6627__118 (.L_HI(net118));
 sg13g2_tiehi _6628__119 (.L_HI(net119));
 sg13g2_tiehi _6629__120 (.L_HI(net120));
 sg13g2_tiehi _6630__121 (.L_HI(net121));
 sg13g2_tiehi _6631__122 (.L_HI(net122));
 sg13g2_tiehi _6632__123 (.L_HI(net123));
 sg13g2_tiehi _6633__124 (.L_HI(net124));
 sg13g2_tiehi _6634__125 (.L_HI(net125));
 sg13g2_tiehi _6635__126 (.L_HI(net126));
 sg13g2_tiehi _6636__127 (.L_HI(net127));
 sg13g2_tiehi _6637__128 (.L_HI(net128));
 sg13g2_tiehi _6638__129 (.L_HI(net129));
 sg13g2_tiehi _6639__130 (.L_HI(net130));
 sg13g2_tiehi _6640__131 (.L_HI(net131));
 sg13g2_tiehi _6641__132 (.L_HI(net132));
 sg13g2_tiehi _6642__133 (.L_HI(net133));
 sg13g2_tiehi _6643__134 (.L_HI(net134));
 sg13g2_tiehi _6644__135 (.L_HI(net135));
 sg13g2_tiehi _6645__136 (.L_HI(net136));
 sg13g2_tiehi _6646__137 (.L_HI(net137));
 sg13g2_tiehi _6647__138 (.L_HI(net138));
 sg13g2_tiehi _6648__139 (.L_HI(net139));
 sg13g2_tiehi _6649__140 (.L_HI(net140));
 sg13g2_tiehi _6650__141 (.L_HI(net141));
 sg13g2_tiehi _6651__142 (.L_HI(net142));
 sg13g2_tiehi _6652__143 (.L_HI(net143));
 sg13g2_tiehi _6653__144 (.L_HI(net144));
 sg13g2_tiehi _6654__145 (.L_HI(net145));
 sg13g2_tiehi _6655__146 (.L_HI(net146));
 sg13g2_tiehi _6656__147 (.L_HI(net147));
 sg13g2_tiehi _6748__148 (.L_HI(net148));
 sg13g2_tiehi _6598__149 (.L_HI(net149));
 sg13g2_tiehi _6747__150 (.L_HI(net150));
 sg13g2_tiehi _6597__151 (.L_HI(net151));
 sg13g2_tiehi _6746__152 (.L_HI(net152));
 sg13g2_tiehi _6596__153 (.L_HI(net153));
 sg13g2_tiehi _6745__154 (.L_HI(net154));
 sg13g2_tiehi _6595__155 (.L_HI(net155));
 sg13g2_tiehi _6744__156 (.L_HI(net156));
 sg13g2_tiehi _6594__157 (.L_HI(net157));
 sg13g2_tiehi _6743__158 (.L_HI(net158));
 sg13g2_tiehi _6593__159 (.L_HI(net159));
 sg13g2_tiehi _6657__160 (.L_HI(net160));
 sg13g2_tiehi _6670__161 (.L_HI(net161));
 sg13g2_tiehi _6671__162 (.L_HI(net162));
 sg13g2_tiehi _6672__163 (.L_HI(net163));
 sg13g2_tiehi _6673__164 (.L_HI(net164));
 sg13g2_tiehi _6674__165 (.L_HI(net165));
 sg13g2_tiehi _6675__166 (.L_HI(net166));
 sg13g2_tiehi _6676__167 (.L_HI(net167));
 sg13g2_tiehi _6677__168 (.L_HI(net168));
 sg13g2_tiehi _6678__169 (.L_HI(net169));
 sg13g2_tiehi _6742__170 (.L_HI(net170));
 sg13g2_tiehi _6592__171 (.L_HI(net171));
 sg13g2_tiehi _6777__172 (.L_HI(net172));
 sg13g2_tiehi _6591__173 (.L_HI(net173));
 sg13g2_tiehi _6741__174 (.L_HI(net174));
 sg13g2_tiehi _6590__175 (.L_HI(net175));
 sg13g2_tiehi _6679__176 (.L_HI(net176));
 sg13g2_tiehi _6686__177 (.L_HI(net177));
 sg13g2_tiehi _6687__178 (.L_HI(net178));
 sg13g2_tiehi _6688__179 (.L_HI(net179));
 sg13g2_tiehi _6689__180 (.L_HI(net180));
 sg13g2_tiehi _6690__181 (.L_HI(net181));
 sg13g2_tiehi _6784__182 (.L_HI(net182));
 sg13g2_tiehi _6589__183 (.L_HI(net183));
 sg13g2_tiehi _6740__184 (.L_HI(net184));
 sg13g2_tiehi _6588__185 (.L_HI(net185));
 sg13g2_tiehi _6587__186 (.L_HI(net186));
 sg13g2_tiehi _6575__187 (.L_HI(net187));
 sg13g2_tiehi _6574__188 (.L_HI(net188));
 sg13g2_tiehi _6573__189 (.L_HI(net189));
 sg13g2_tiehi _6572__190 (.L_HI(net190));
 sg13g2_tiehi _6571__191 (.L_HI(net191));
 sg13g2_tiehi _6570__192 (.L_HI(net192));
 sg13g2_tiehi _6569__193 (.L_HI(net193));
 sg13g2_tiehi _6568__194 (.L_HI(net194));
 sg13g2_tiehi _6567__195 (.L_HI(net195));
 sg13g2_tiehi _6566__196 (.L_HI(net196));
 sg13g2_tiehi _6565__197 (.L_HI(net197));
 sg13g2_tiehi _6691__198 (.L_HI(net198));
 sg13g2_tiehi _6564__199 (.L_HI(net199));
 sg13g2_tiehi _6563__200 (.L_HI(net200));
 sg13g2_tiehi _6562__201 (.L_HI(net201));
 sg13g2_tiehi _6561__202 (.L_HI(net202));
 sg13g2_tiehi _6560__203 (.L_HI(net203));
 sg13g2_tiehi _6559__204 (.L_HI(net204));
 sg13g2_tiehi _6558__205 (.L_HI(net205));
 sg13g2_tiehi _6557__206 (.L_HI(net206));
 sg13g2_tiehi _6556__207 (.L_HI(net207));
 sg13g2_tiehi _6555__208 (.L_HI(net208));
 sg13g2_tiehi _6554__209 (.L_HI(net209));
 sg13g2_tiehi _6553__210 (.L_HI(net210));
 sg13g2_tiehi _6552__211 (.L_HI(net211));
 sg13g2_tiehi _6551__212 (.L_HI(net212));
 sg13g2_tiehi _6550__213 (.L_HI(net213));
 sg13g2_tiehi _6549__214 (.L_HI(net214));
 sg13g2_tiehi _6548__215 (.L_HI(net215));
 sg13g2_tiehi _6547__216 (.L_HI(net216));
 sg13g2_tiehi _6776__217 (.L_HI(net217));
 sg13g2_tiehi _6546__218 (.L_HI(net218));
 sg13g2_tiehi _6739__219 (.L_HI(net219));
 sg13g2_tiehi _6545__220 (.L_HI(net220));
 sg13g2_tiehi _6543__221 (.L_HI(net221));
 sg13g2_tiehi _6542__222 (.L_HI(net222));
 sg13g2_tiehi _6541__223 (.L_HI(net223));
 sg13g2_tiehi _6540__224 (.L_HI(net224));
 sg13g2_tiehi _6539__225 (.L_HI(net225));
 sg13g2_tiehi _6781__226 (.L_HI(net226));
 sg13g2_tiehi _6738__227 (.L_HI(net227));
 sg13g2_tiehi _6775__228 (.L_HI(net228));
 sg13g2_tiehi _6737__229 (.L_HI(net229));
 sg13g2_tiehi _6787__230 (.L_HI(net230));
 sg13g2_tiehi _6736__231 (.L_HI(net231));
 sg13g2_tiehi _6774__232 (.L_HI(net232));
 sg13g2_tiehi _6735__233 (.L_HI(net233));
 sg13g2_tiehi _6773__234 (.L_HI(net234));
 sg13g2_tiehi _6734__235 (.L_HI(net235));
 sg13g2_tiehi _6772__236 (.L_HI(net236));
 sg13g2_tiehi _6733__237 (.L_HI(net237));
 sg13g2_tiehi _6771__238 (.L_HI(net238));
 sg13g2_tiehi _6732__239 (.L_HI(net239));
 sg13g2_tiehi _6770__240 (.L_HI(net240));
 sg13g2_tiehi _6731__241 (.L_HI(net241));
 sg13g2_tiehi _6769__242 (.L_HI(net242));
 sg13g2_tiehi _6730__243 (.L_HI(net243));
 sg13g2_tiehi _6768__244 (.L_HI(net244));
 sg13g2_tiehi _6729__245 (.L_HI(net245));
 sg13g2_tiehi _6728__246 (.L_HI(net246));
 sg13g2_tiehi _6767__247 (.L_HI(net247));
 sg13g2_tiehi _6727__248 (.L_HI(net248));
 sg13g2_tiehi _6766__249 (.L_HI(net249));
 sg13g2_tiehi _6726__250 (.L_HI(net250));
 sg13g2_tiehi _6765__251 (.L_HI(net251));
 sg13g2_tiehi _6725__252 (.L_HI(net252));
 sg13g2_tiehi _6780__253 (.L_HI(net253));
 sg13g2_tiehi _6724__254 (.L_HI(net254));
 sg13g2_tiehi _6764__255 (.L_HI(net255));
 sg13g2_tiehi _6723__256 (.L_HI(net256));
 sg13g2_tiehi _6783__257 (.L_HI(net257));
 sg13g2_tiehi _6722__258 (.L_HI(net258));
 sg13g2_tiehi _6763__259 (.L_HI(net259));
 sg13g2_tiehi _6721__260 (.L_HI(net260));
 sg13g2_tiehi _6779__261 (.L_HI(net261));
 sg13g2_tiehi _6720__262 (.L_HI(net262));
 sg13g2_tiehi _6762__263 (.L_HI(net263));
 sg13g2_tiehi _6719__264 (.L_HI(net264));
 sg13g2_tiehi _6718__265 (.L_HI(net265));
 sg13g2_tiehi _6717__266 (.L_HI(net266));
 sg13g2_tiehi _6716__267 (.L_HI(net267));
 sg13g2_tiehi _6715__268 (.L_HI(net268));
 sg13g2_tiehi _6714__269 (.L_HI(net269));
 sg13g2_tiehi _6713__270 (.L_HI(net270));
 sg13g2_tiehi _6712__271 (.L_HI(net271));
 sg13g2_tiehi _6786__272 (.L_HI(net272));
 sg13g2_tiehi _6711__273 (.L_HI(net273));
 sg13g2_tiehi _6761__274 (.L_HI(net274));
 sg13g2_tiehi _6708__275 (.L_HI(net275));
 sg13g2_tiehi _6785__276 (.L_HI(net276));
 sg13g2_tiehi tt_um_warp_277 (.L_HI(net277));
 sg13g2_buf_2 clkbuf_leaf_0_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_tielo tt_um_warp_3 (.L_LO(net3));
 sg13g2_tielo tt_um_warp_4 (.L_LO(net4));
 sg13g2_tielo tt_um_warp_5 (.L_LO(net5));
 sg13g2_tielo tt_um_warp_6 (.L_LO(net6));
 sg13g2_tielo tt_um_warp_7 (.L_LO(net7));
 sg13g2_tielo tt_um_warp_8 (.L_LO(net8));
 sg13g2_tielo tt_um_warp_9 (.L_LO(net9));
 sg13g2_tielo tt_um_warp_10 (.L_LO(net10));
 sg13g2_tielo tt_um_warp_11 (.L_LO(net11));
 sg13g2_tielo tt_um_warp_12 (.L_LO(net12));
 sg13g2_tielo tt_um_warp_13 (.L_LO(net13));
 sg13g2_tielo tt_um_warp_14 (.L_LO(net14));
 sg13g2_tielo tt_um_warp_15 (.L_LO(net15));
 sg13g2_tiehi _6710__16 (.L_HI(net16));
 sg13g2_buf_1 _7064_ (.A(\main.demo._q_prev_vs ),
    .X(uo_out[3]));
 sg13g2_buf_2 fanout339 (.A(\main.demo._d___pip_58_1_1___stage___block_3_a[1] ),
    .X(net339));
 sg13g2_buf_1 fanout340 (.A(\main.demo._d___pip_58_1_1___stage___block_3_a[1] ),
    .X(net340));
 sg13g2_buf_2 fanout341 (.A(_1592_),
    .X(net341));
 sg13g2_buf_2 fanout342 (.A(_1044_),
    .X(net342));
 sg13g2_buf_2 fanout343 (.A(_1603_),
    .X(net343));
 sg13g2_buf_4 fanout344 (.X(net344),
    .A(\main.demo._d___pip_58_1_1___stage___block_3_a[2] ));
 sg13g2_buf_2 fanout345 (.A(_0277_),
    .X(net345));
 sg13g2_buf_2 fanout346 (.A(_3023_),
    .X(net346));
 sg13g2_buf_2 fanout347 (.A(\main.demo._d___pip_58_1_1___stage___block_3_a[3] ),
    .X(net347));
 sg13g2_buf_1 fanout348 (.A(\main.demo._d___pip_58_1_1___stage___block_3_a[3] ),
    .X(net348));
 sg13g2_buf_4 fanout349 (.X(net349),
    .A(_2803_));
 sg13g2_buf_2 fanout350 (.A(_2803_),
    .X(net350));
 sg13g2_buf_2 fanout351 (.A(net352),
    .X(net351));
 sg13g2_buf_4 fanout352 (.X(net352),
    .A(_2802_));
 sg13g2_buf_2 fanout353 (.A(net357),
    .X(net353));
 sg13g2_buf_2 fanout354 (.A(net357),
    .X(net354));
 sg13g2_buf_2 fanout355 (.A(net356),
    .X(net355));
 sg13g2_buf_2 fanout356 (.A(net357),
    .X(net356));
 sg13g2_buf_1 fanout357 (.A(\main.demo._t___pip_58_1_0___stage___block_3_a[6] ),
    .X(net357));
 sg13g2_buf_2 fanout358 (.A(_0704_),
    .X(net358));
 sg13g2_buf_2 fanout359 (.A(_2474_),
    .X(net359));
 sg13g2_buf_1 fanout360 (.A(_2474_),
    .X(net360));
 sg13g2_buf_2 fanout361 (.A(_2473_),
    .X(net361));
 sg13g2_buf_2 fanout362 (.A(_1886_),
    .X(net362));
 sg13g2_buf_2 fanout363 (.A(net364),
    .X(net363));
 sg13g2_buf_2 fanout364 (.A(_2118_),
    .X(net364));
 sg13g2_buf_2 fanout365 (.A(_2112_),
    .X(net365));
 sg13g2_buf_2 fanout366 (.A(_0234_),
    .X(net366));
 sg13g2_buf_1 fanout367 (.A(_0234_),
    .X(net367));
 sg13g2_buf_2 fanout368 (.A(_2386_),
    .X(net368));
 sg13g2_buf_2 fanout369 (.A(_2386_),
    .X(net369));
 sg13g2_buf_2 fanout370 (.A(_2358_),
    .X(net370));
 sg13g2_buf_2 fanout371 (.A(net372),
    .X(net371));
 sg13g2_buf_1 fanout372 (.A(net373),
    .X(net372));
 sg13g2_buf_2 fanout373 (.A(_2086_),
    .X(net373));
 sg13g2_buf_2 fanout374 (.A(_0231_),
    .X(net374));
 sg13g2_buf_2 fanout375 (.A(net376),
    .X(net375));
 sg13g2_buf_4 fanout376 (.X(net376),
    .A(net379));
 sg13g2_buf_2 fanout377 (.A(net378),
    .X(net377));
 sg13g2_buf_2 fanout378 (.A(net379),
    .X(net378));
 sg13g2_buf_4 fanout379 (.X(net379),
    .A(_2210_));
 sg13g2_buf_4 fanout380 (.X(net380),
    .A(_1218_));
 sg13g2_buf_4 fanout381 (.X(net381),
    .A(_1017_));
 sg13g2_buf_2 fanout382 (.A(net383),
    .X(net382));
 sg13g2_buf_4 fanout383 (.X(net383),
    .A(net384));
 sg13g2_buf_4 fanout384 (.X(net384),
    .A(_1016_));
 sg13g2_buf_2 fanout385 (.A(net386),
    .X(net385));
 sg13g2_buf_2 fanout386 (.A(_0922_),
    .X(net386));
 sg13g2_buf_2 fanout387 (.A(_0898_),
    .X(net387));
 sg13g2_buf_4 fanout388 (.X(net388),
    .A(net389));
 sg13g2_buf_2 fanout389 (.A(net390),
    .X(net389));
 sg13g2_buf_2 fanout390 (.A(_0897_),
    .X(net390));
 sg13g2_buf_2 fanout391 (.A(net392),
    .X(net391));
 sg13g2_buf_1 fanout392 (.A(_2939_),
    .X(net392));
 sg13g2_buf_4 fanout393 (.X(net393),
    .A(_2675_));
 sg13g2_buf_2 fanout394 (.A(_2675_),
    .X(net394));
 sg13g2_buf_2 fanout395 (.A(net397),
    .X(net395));
 sg13g2_buf_2 fanout396 (.A(net397),
    .X(net396));
 sg13g2_buf_1 fanout397 (.A(net398),
    .X(net397));
 sg13g2_buf_4 fanout398 (.X(net398),
    .A(net399));
 sg13g2_buf_1 fanout399 (.A(_2674_),
    .X(net399));
 sg13g2_buf_2 fanout400 (.A(net401),
    .X(net400));
 sg13g2_buf_2 fanout401 (.A(net402),
    .X(net401));
 sg13g2_buf_4 fanout402 (.X(net402),
    .A(net403));
 sg13g2_buf_4 fanout403 (.X(net403),
    .A(_2637_));
 sg13g2_buf_4 fanout404 (.X(net404),
    .A(_2621_));
 sg13g2_buf_4 fanout405 (.X(net405),
    .A(_2614_));
 sg13g2_buf_1 fanout406 (.A(_2614_),
    .X(net406));
 sg13g2_buf_2 fanout407 (.A(\main.demo._t___stage___block_3_y[1] ),
    .X(net407));
 sg13g2_buf_2 fanout408 (.A(net409),
    .X(net408));
 sg13g2_buf_2 fanout409 (.A(\main.demo.zic._q_idx[3] ),
    .X(net409));
 sg13g2_buf_2 fanout410 (.A(net411),
    .X(net410));
 sg13g2_buf_2 fanout411 (.A(net638),
    .X(net411));
 sg13g2_buf_2 fanout412 (.A(\main.demo._w_vga_vga_x[8] ),
    .X(net412));
 sg13g2_buf_2 fanout413 (.A(\main.demo._w_vga_vga_x[7] ),
    .X(net413));
 sg13g2_buf_2 fanout414 (.A(\main.demo._w_vga_vga_x[6] ),
    .X(net414));
 sg13g2_buf_4 fanout415 (.X(net415),
    .A(net611));
 sg13g2_buf_2 fanout416 (.A(net417),
    .X(net416));
 sg13g2_buf_1 fanout417 (.A(\main.demo._q_effect[1] ),
    .X(net417));
 sg13g2_buf_2 fanout418 (.A(\main.demo._q_effect[1] ),
    .X(net418));
 sg13g2_buf_2 fanout419 (.A(net639),
    .X(net419));
 sg13g2_buf_2 fanout420 (.A(net421),
    .X(net420));
 sg13g2_buf_1 fanout421 (.A(\main.demo._q_effect[0] ),
    .X(net421));
 sg13g2_buf_4 fanout422 (.X(net422),
    .A(\main.demo._q_rot_en ));
 sg13g2_buf_4 fanout423 (.X(net423),
    .A(\main.demo._d___pip_58_1_4___block_87_atten_l[1] ));
 sg13g2_buf_4 fanout424 (.X(net424),
    .A(\main.demo._d___pip_58_1_4___block_87_atten_l[0] ));
 sg13g2_buf_4 fanout425 (.X(net425),
    .A(net494));
 sg13g2_buf_4 fanout426 (.X(net426),
    .A(_0006_));
 sg13g2_buf_2 fanout427 (.A(net563),
    .X(net427));
 sg13g2_buf_4 fanout428 (.X(net428),
    .A(net580));
 sg13g2_buf_2 fanout429 (.A(net430),
    .X(net429));
 sg13g2_buf_1 fanout430 (.A(net431),
    .X(net430));
 sg13g2_buf_2 fanout431 (.A(\main.demo._q___pip_58_1_1___stage___block_3_cy[10] ),
    .X(net431));
 sg13g2_buf_2 fanout432 (.A(\main.demo._q___pip_58_1_1___stage___block_3_cy[10] ),
    .X(net432));
 sg13g2_buf_2 fanout433 (.A(\main.demo._q___pip_58_1_1___stage___block_3_cy[10] ),
    .X(net433));
 sg13g2_buf_4 fanout434 (.X(net434),
    .A(\main.demo._q_frame[7] ));
 sg13g2_buf_2 fanout435 (.A(\main.demo._q_frame[4] ),
    .X(net435));
 sg13g2_buf_2 fanout436 (.A(\main.demo._q_frame[3] ),
    .X(net436));
 sg13g2_buf_2 fanout437 (.A(net438),
    .X(net437));
 sg13g2_buf_2 fanout438 (.A(net439),
    .X(net438));
 sg13g2_buf_2 fanout439 (.A(net559),
    .X(net439));
 sg13g2_buf_4 fanout440 (.X(net440),
    .A(net560));
 sg13g2_buf_4 fanout441 (.X(net441),
    .A(net560));
 sg13g2_buf_2 fanout442 (.A(net443),
    .X(net442));
 sg13g2_buf_2 fanout443 (.A(net444),
    .X(net443));
 sg13g2_buf_2 fanout444 (.A(rst_n_q),
    .X(net444));
 sg13g2_buf_2 fanout445 (.A(net446),
    .X(net445));
 sg13g2_buf_1 fanout446 (.A(net447),
    .X(net446));
 sg13g2_buf_2 fanout447 (.A(net448),
    .X(net447));
 sg13g2_buf_2 fanout448 (.A(net450),
    .X(net448));
 sg13g2_buf_2 fanout449 (.A(net450),
    .X(net449));
 sg13g2_buf_2 fanout450 (.A(\main.demo._q___pip_58_1_2___stage___block_3_cy[10] ),
    .X(net450));
 sg13g2_buf_2 input1 (.A(rst_n),
    .X(net1));
 sg13g2_tielo tt_um_warp_2 (.L_LO(net2));
 sg13g2_buf_2 clkbuf_leaf_1_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_2 clkbuf_leaf_2_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_2 clkbuf_leaf_3_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_2 clkbuf_leaf_4_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_2 clkbuf_leaf_5_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_2 clkbuf_leaf_6_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_2 clkbuf_leaf_7_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_2 clkbuf_leaf_8_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_2 clkbuf_leaf_9_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_2 clkbuf_leaf_10_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_2 clkbuf_leaf_11_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_2 clkbuf_leaf_12_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_2 clkbuf_leaf_13_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_2 clkbuf_leaf_14_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_2 clkbuf_leaf_15_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_2 clkbuf_leaf_16_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_2 clkbuf_leaf_17_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_2 clkbuf_leaf_18_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_2 clkbuf_leaf_19_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_2 clkbuf_leaf_20_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_2 clkbuf_leaf_21_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_2 clkbuf_leaf_22_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_2 clkbuf_leaf_23_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_2 clkbuf_leaf_24_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_2 clkbuf_leaf_26_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_2 clkbuf_leaf_27_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_2 clkbuf_leaf_28_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_2 clkbuf_leaf_29_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_2 clkbuf_leaf_30_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_2 clkbuf_leaf_31_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_31_clk));
 sg13g2_buf_2 clkbuf_leaf_32_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_32_clk));
 sg13g2_buf_2 clkbuf_leaf_33_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_33_clk));
 sg13g2_buf_2 clkbuf_leaf_34_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_34_clk));
 sg13g2_buf_2 clkbuf_leaf_36_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_36_clk));
 sg13g2_buf_2 clkbuf_leaf_37_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_37_clk));
 sg13g2_buf_2 clkbuf_leaf_38_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_38_clk));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_2 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sg13g2_buf_2 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sg13g2_buf_2 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sg13g2_buf_2 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sg13g2_buf_2 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sg13g2_buf_2 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sg13g2_buf_2 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sg13g2_buf_2 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sg13g2_buf_1 clkload0 (.A(clknet_3_0__leaf_clk));
 sg13g2_buf_1 clkload1 (.A(clknet_3_1__leaf_clk));
 sg13g2_buf_1 clkload2 (.A(clknet_3_3__leaf_clk));
 sg13g2_buf_1 clkload3 (.A(clknet_3_4__leaf_clk));
 sg13g2_buf_1 clkload4 (.A(clknet_3_5__leaf_clk));
 sg13g2_buf_1 clkload5 (.A(clknet_3_6__leaf_clk));
 sg13g2_buf_2 clkload6 (.A(clknet_3_7__leaf_clk));
 sg13g2_inv_8 clkload7 (.A(clknet_leaf_1_clk));
 sg13g2_inv_1 clkload8 (.A(clknet_leaf_38_clk));
 sg13g2_inv_4 clkload9 (.A(clknet_leaf_2_clk));
 sg13g2_inv_4 clkload10 (.A(clknet_leaf_3_clk));
 sg13g2_inv_8 clkload11 (.A(clknet_leaf_4_clk));
 sg13g2_inv_1 clkload12 (.A(clknet_leaf_31_clk));
 sg13g2_inv_4 clkload13 (.A(clknet_leaf_6_clk));
 sg13g2_inv_2 clkload14 (.A(clknet_leaf_30_clk));
 sg13g2_inv_1 clkload15 (.A(clknet_leaf_11_clk));
 sg13g2_inv_1 clkload16 (.A(clknet_leaf_16_clk));
 sg13g2_inv_1 clkload17 (.A(clknet_leaf_17_clk));
 sg13g2_inv_4 clkload18 (.A(clknet_leaf_20_clk));
 sg13g2_inv_2 clkload19 (.A(clknet_leaf_27_clk));
 sg13g2_inv_2 clkload20 (.A(clknet_leaf_26_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\main._w_demo_video_hs ),
    .X(net278));
 sg13g2_dlygate4sd3_1 hold2 (.A(\main.demo._d_prev_b[4] ),
    .X(net279));
 sg13g2_dlygate4sd3_1 hold3 (.A(\main.demo._d_prev_b[6] ),
    .X(net280));
 sg13g2_dlygate4sd3_1 hold4 (.A(\main.demo._d_prev_b[5] ),
    .X(net281));
 sg13g2_dlygate4sd3_1 hold5 (.A(\main.demo._d_prev_b[2] ),
    .X(net282));
 sg13g2_dlygate4sd3_1 hold6 (.A(\main.demo._d_prev_b[7] ),
    .X(net283));
 sg13g2_dlygate4sd3_1 hold7 (.A(_0064_),
    .X(net284));
 sg13g2_dlygate4sd3_1 hold8 (.A(\main.demo._d_prev_b[3] ),
    .X(net285));
 sg13g2_dlygate4sd3_1 hold9 (.A(\main._w_demo_video_vs ),
    .X(net286));
 sg13g2_dlygate4sd3_1 hold10 (.A(_0069_),
    .X(net287));
 sg13g2_dlygate4sd3_1 hold11 (.A(\main.demo._d___pip_58_1_1___stage___block_3_a[7] ),
    .X(net288));
 sg13g2_dlygate4sd3_1 hold12 (.A(_0066_),
    .X(net289));
 sg13g2_dlygate4sd3_1 hold13 (.A(_2360_),
    .X(net290));
 sg13g2_dlygate4sd3_1 hold14 (.A(_0123_),
    .X(net291));
 sg13g2_dlygate4sd3_1 hold15 (.A(_0065_),
    .X(net292));
 sg13g2_dlygate4sd3_1 hold16 (.A(_0173_),
    .X(net293));
 sg13g2_dlygate4sd3_1 hold17 (.A(_0068_),
    .X(net294));
 sg13g2_dlygate4sd3_1 hold18 (.A(\main.demo._d___pip_58_1_1___stage___block_3_a[6] ),
    .X(net295));
 sg13g2_dlygate4sd3_1 hold19 (.A(_0000_),
    .X(net296));
 sg13g2_dlygate4sd3_1 hold20 (.A(_2352_),
    .X(net297));
 sg13g2_dlygate4sd3_1 hold21 (.A(_0120_),
    .X(net298));
 sg13g2_dlygate4sd3_1 hold22 (.A(\main.demo.zic._q_qpos[0] ),
    .X(net299));
 sg13g2_dlygate4sd3_1 hold23 (.A(\main.demo._d___pip_58_1_3___stage___block_3_cx[6] ),
    .X(net300));
 sg13g2_dlygate4sd3_1 hold24 (.A(_0002_),
    .X(net301));
 sg13g2_dlygate4sd3_1 hold25 (.A(_0155_),
    .X(net302));
 sg13g2_dlygate4sd3_1 hold26 (.A(_0027_),
    .X(net303));
 sg13g2_dlygate4sd3_1 hold27 (.A(_1499_),
    .X(net304));
 sg13g2_dlygate4sd3_1 hold28 (.A(\main._w_demo_audio1 ),
    .X(net305));
 sg13g2_dlygate4sd3_1 hold29 (.A(\main.demo._q_th[1] ),
    .X(net306));
 sg13g2_dlygate4sd3_1 hold30 (.A(_2362_),
    .X(net307));
 sg13g2_dlygate4sd3_1 hold31 (.A(_0124_),
    .X(net308));
 sg13g2_dlygate4sd3_1 hold32 (.A(\main.demo.vga._q_xcount[0] ),
    .X(net309));
 sg13g2_dlygate4sd3_1 hold33 (.A(\main.demo.zic._q_qpos[10] ),
    .X(net310));
 sg13g2_dlygate4sd3_1 hold34 (.A(_0117_),
    .X(net311));
 sg13g2_dlygate4sd3_1 hold35 (.A(\main.demo._q_th[7] ),
    .X(net312));
 sg13g2_dlygate4sd3_1 hold36 (.A(_2374_),
    .X(net313));
 sg13g2_dlygate4sd3_1 hold37 (.A(_2375_),
    .X(net314));
 sg13g2_dlygate4sd3_1 hold38 (.A(_0131_),
    .X(net315));
 sg13g2_dlygate4sd3_1 hold39 (.A(\main.demo.vga._q_xcount[2] ),
    .X(net316));
 sg13g2_dlygate4sd3_1 hold40 (.A(\main.demo.zic._q_qpos[5] ),
    .X(net317));
 sg13g2_dlygate4sd3_1 hold41 (.A(\main.demo.zic._q_qpos[3] ),
    .X(net318));
 sg13g2_dlygate4sd3_1 hold42 (.A(\main.demo.vga._q_ycount[5] ),
    .X(net319));
 sg13g2_dlygate4sd3_1 hold43 (.A(_2469_),
    .X(net320));
 sg13g2_dlygate4sd3_1 hold44 (.A(\main.demo.zic._q_tpos[9] ),
    .X(net321));
 sg13g2_dlygate4sd3_1 hold45 (.A(_2598_),
    .X(net322));
 sg13g2_dlygate4sd3_1 hold46 (.A(\main.demo.zic._q_rythm_count[6] ),
    .X(net323));
 sg13g2_dlygate4sd3_1 hold47 (.A(_2488_),
    .X(net324));
 sg13g2_dlygate4sd3_1 hold48 (.A(_0179_),
    .X(net325));
 sg13g2_dlygate4sd3_1 hold49 (.A(\main.demo.zic._q_rythm_count[1] ),
    .X(net326));
 sg13g2_dlygate4sd3_1 hold50 (.A(_2477_),
    .X(net327));
 sg13g2_dlygate4sd3_1 hold51 (.A(_0174_),
    .X(net328));
 sg13g2_dlygate4sd3_1 hold52 (.A(\main.demo.zic._q_qpos[7] ),
    .X(net329));
 sg13g2_dlygate4sd3_1 hold53 (.A(_2341_),
    .X(net330));
 sg13g2_dlygate4sd3_1 hold54 (.A(_0114_),
    .X(net331));
 sg13g2_dlygate4sd3_1 hold55 (.A(\main.demo.zic._q_qpos[1] ),
    .X(net332));
 sg13g2_dlygate4sd3_1 hold56 (.A(_0108_),
    .X(net333));
 sg13g2_dlygate4sd3_1 hold57 (.A(\main.demo.zic._q_rythm_count[10] ),
    .X(net334));
 sg13g2_dlygate4sd3_1 hold58 (.A(_2496_),
    .X(net335));
 sg13g2_dlygate4sd3_1 hold59 (.A(\main.demo.zic._q_tpos[8] ),
    .X(net336));
 sg13g2_dlygate4sd3_1 hold60 (.A(_0226_),
    .X(net337));
 sg13g2_dlygate4sd3_1 hold61 (.A(\main.demo.zic._q_rythm_count[7] ),
    .X(net338));
 sg13g2_dlygate4sd3_1 hold62 (.A(_2491_),
    .X(net451));
 sg13g2_dlygate4sd3_1 hold63 (.A(\main.demo.vga._q_xcount[1] ),
    .X(net452));
 sg13g2_dlygate4sd3_1 hold64 (.A(\main.demo.zic._q_clock_count[3] ),
    .X(net453));
 sg13g2_dlygate4sd3_1 hold65 (.A(_2526_),
    .X(net454));
 sg13g2_dlygate4sd3_1 hold66 (.A(\main.demo._d___pip_58_1_3___stage___block_3_cx[4] ),
    .X(net455));
 sg13g2_dlygate4sd3_1 hold67 (.A(\main.demo.vga._q_xcount[4] ),
    .X(net456));
 sg13g2_dlygate4sd3_1 hold68 (.A(\main.demo._w_vga_active ),
    .X(net457));
 sg13g2_dlygate4sd3_1 hold69 (.A(\main.demo.vga._q_ycount[6] ),
    .X(net458));
 sg13g2_dlygate4sd3_1 hold70 (.A(_0199_),
    .X(net459));
 sg13g2_dlygate4sd3_1 hold71 (.A(\main.demo.vga._q_xcount[6] ),
    .X(net460));
 sg13g2_dlygate4sd3_1 hold72 (.A(\main.demo.zic._q_rythm_count[11] ),
    .X(net461));
 sg13g2_dlygate4sd3_1 hold73 (.A(\main.demo.zic._q_qpos[8] ),
    .X(net462));
 sg13g2_dlygate4sd3_1 hold74 (.A(_2343_),
    .X(net463));
 sg13g2_dlygate4sd3_1 hold75 (.A(_0115_),
    .X(net464));
 sg13g2_dlygate4sd3_1 hold76 (.A(\main.demo.vga._q_ycount[1] ),
    .X(net465));
 sg13g2_dlygate4sd3_1 hold77 (.A(_0194_),
    .X(net466));
 sg13g2_dlygate4sd3_1 hold78 (.A(\main.demo._q_prev_b[7] ),
    .X(net467));
 sg13g2_dlygate4sd3_1 hold79 (.A(\main.demo.vga._q_xcount[5] ),
    .X(net468));
 sg13g2_dlygate4sd3_1 hold80 (.A(\main.demo.vga._q_ycount[8] ),
    .X(net469));
 sg13g2_dlygate4sd3_1 hold81 (.A(_0201_),
    .X(net470));
 sg13g2_dlygate4sd3_1 hold82 (.A(\main.demo.zic._q_clock_count[5] ),
    .X(net471));
 sg13g2_dlygate4sd3_1 hold83 (.A(_2530_),
    .X(net472));
 sg13g2_dlygate4sd3_1 hold84 (.A(\main.demo.zic._q_tpos[7] ),
    .X(net473));
 sg13g2_dlygate4sd3_1 hold85 (.A(_2595_),
    .X(net474));
 sg13g2_dlygate4sd3_1 hold86 (.A(\main.demo.vga._q_ycount[3] ),
    .X(net475));
 sg13g2_dlygate4sd3_1 hold87 (.A(_0196_),
    .X(net476));
 sg13g2_dlygate4sd3_1 hold88 (.A(\main.demo.zic._q_clock_count[2] ),
    .X(net477));
 sg13g2_dlygate4sd3_1 hold89 (.A(_2524_),
    .X(net478));
 sg13g2_dlygate4sd3_1 hold90 (.A(\main.demo.zic._q_qpos[11] ),
    .X(net479));
 sg13g2_dlygate4sd3_1 hold91 (.A(_2349_),
    .X(net480));
 sg13g2_dlygate4sd3_1 hold92 (.A(_0119_),
    .X(net481));
 sg13g2_dlygate4sd3_1 hold93 (.A(\main.demo.vga._q_xcount[7] ),
    .X(net482));
 sg13g2_dlygate4sd3_1 hold94 (.A(\main.demo.zic._q_rythm_count[3] ),
    .X(net483));
 sg13g2_dlygate4sd3_1 hold95 (.A(_2482_),
    .X(net484));
 sg13g2_dlygate4sd3_1 hold96 (.A(\main.demo.vga._d_vblank ),
    .X(net485));
 sg13g2_dlygate4sd3_1 hold97 (.A(_0202_),
    .X(net486));
 sg13g2_dlygate4sd3_1 hold98 (.A(\main.demo.zic._q_rythm_count[4] ),
    .X(net487));
 sg13g2_dlygate4sd3_1 hold99 (.A(\main.demo.vga._q_xcount[4] ),
    .X(net488));
 sg13g2_dlygate4sd3_1 hold100 (.A(\main.demo.vga._q_xcount[8] ),
    .X(net489));
 sg13g2_dlygate4sd3_1 hold101 (.A(\main.demo.zic._q_rythm_count[5] ),
    .X(net490));
 sg13g2_dlygate4sd3_1 hold102 (.A(\main.demo.zic._q_rythm_count[8] ),
    .X(net491));
 sg13g2_dlygate4sd3_1 hold103 (.A(\main.demo.zic._q_rythm_count[2] ),
    .X(net492));
 sg13g2_dlygate4sd3_1 hold104 (.A(_2480_),
    .X(net493));
 sg13g2_dlygate4sd3_1 hold105 (.A(\main.demo._d___pip_58_1_3___stage___block_3_cx[9] ),
    .X(net494));
 sg13g2_dlygate4sd3_1 hold106 (.A(\main.demo.zic._q_rythm_count[9] ),
    .X(net495));
 sg13g2_dlygate4sd3_1 hold107 (.A(\main.demo.zic._q_clock_count[6] ),
    .X(net496));
 sg13g2_dlygate4sd3_1 hold108 (.A(\main.demo._q_prev_b[6] ),
    .X(net497));
 sg13g2_dlygate4sd3_1 hold109 (.A(\main.demo._q_speed[15] ),
    .X(net498));
 sg13g2_dlygate4sd3_1 hold110 (.A(_0091_),
    .X(net499));
 sg13g2_dlygate4sd3_1 hold111 (.A(\main.demo._q_frame[7] ),
    .X(net500));
 sg13g2_dlygate4sd3_1 hold112 (.A(\main.demo.vga._q_ycount[4] ),
    .X(net501));
 sg13g2_dlygate4sd3_1 hold113 (.A(_0197_),
    .X(net502));
 sg13g2_dlygate4sd3_1 hold114 (.A(\main.demo.zic._q_clock_count[4] ),
    .X(net503));
 sg13g2_dlygate4sd3_1 hold115 (.A(\main.demo.vga._q_xcount[3] ),
    .X(net504));
 sg13g2_dlygate4sd3_1 hold116 (.A(_0002_),
    .X(net505));
 sg13g2_dlygate4sd3_1 hold117 (.A(\main.demo.zic._q_rythm_count[12] ),
    .X(net506));
 sg13g2_dlygate4sd3_1 hold118 (.A(\main.demo.zic._q_clock_count[8] ),
    .X(net507));
 sg13g2_dlygate4sd3_1 hold119 (.A(_2535_),
    .X(net508));
 sg13g2_dlygate4sd3_1 hold120 (.A(\main.demo.zic._q_tpos[2] ),
    .X(net509));
 sg13g2_dlygate4sd3_1 hold121 (.A(_2571_),
    .X(net510));
 sg13g2_dlygate4sd3_1 hold122 (.A(_0033_),
    .X(net511));
 sg13g2_dlygate4sd3_1 hold123 (.A(_2592_),
    .X(net512));
 sg13g2_dlygate4sd3_1 hold124 (.A(\main.demo.vga._q_ycount[2] ),
    .X(net513));
 sg13g2_dlygate4sd3_1 hold125 (.A(_2467_),
    .X(net514));
 sg13g2_dlygate4sd3_1 hold126 (.A(_0166_),
    .X(net515));
 sg13g2_dlygate4sd3_1 hold127 (.A(\main.demo.vga._q_xcount[10] ),
    .X(net516));
 sg13g2_dlygate4sd3_1 hold128 (.A(_0005_),
    .X(net517));
 sg13g2_dlygate4sd3_1 hold129 (.A(\main.demo.zic._q_tpos[1] ),
    .X(net518));
 sg13g2_dlygate4sd3_1 hold130 (.A(_2563_),
    .X(net519));
 sg13g2_dlygate4sd3_1 hold131 (.A(_0219_),
    .X(net520));
 sg13g2_dlygate4sd3_1 hold132 (.A(\main.demo.vga._q_ycount[0] ),
    .X(net521));
 sg13g2_dlygate4sd3_1 hold133 (.A(_0164_),
    .X(net522));
 sg13g2_dlygate4sd3_1 hold134 (.A(\main.demo._q_th[4] ),
    .X(net523));
 sg13g2_dlygate4sd3_1 hold135 (.A(_0026_),
    .X(net524));
 sg13g2_dlygate4sd3_1 hold136 (.A(_2533_),
    .X(net525));
 sg13g2_dlygate4sd3_1 hold137 (.A(\main.demo._d___pip_58_1_3___stage___block_3_cx[2] ),
    .X(net526));
 sg13g2_dlygate4sd3_1 hold138 (.A(\main.demo._q_th[6] ),
    .X(net527));
 sg13g2_dlygate4sd3_1 hold139 (.A(_2371_),
    .X(net528));
 sg13g2_dlygate4sd3_1 hold140 (.A(\main.demo.zic._q_tpos[10] ),
    .X(net529));
 sg13g2_dlygate4sd3_1 hold141 (.A(\main.demo.zic._q_tpos[11] ),
    .X(net530));
 sg13g2_dlygate4sd3_1 hold142 (.A(\main.demo.vga._d_vblank ),
    .X(net531));
 sg13g2_dlygate4sd3_1 hold143 (.A(_2442_),
    .X(net532));
 sg13g2_dlygate4sd3_1 hold144 (.A(_0154_),
    .X(net533));
 sg13g2_dlygate4sd3_1 hold145 (.A(\main.demo.zic._q_tpos[3] ),
    .X(net534));
 sg13g2_dlygate4sd3_1 hold146 (.A(_2581_),
    .X(net535));
 sg13g2_dlygate4sd3_1 hold147 (.A(\main.demo.zic._q_tpos[0] ),
    .X(net536));
 sg13g2_dlygate4sd3_1 hold148 (.A(_2550_),
    .X(net537));
 sg13g2_dlygate4sd3_1 hold149 (.A(_0218_),
    .X(net538));
 sg13g2_dlygate4sd3_1 hold150 (.A(\main.demo._q_th[5] ),
    .X(net539));
 sg13g2_dlygate4sd3_1 hold151 (.A(\main.demo.vga._q_xcount[9] ),
    .X(net540));
 sg13g2_dlygate4sd3_1 hold152 (.A(_0067_),
    .X(net541));
 sg13g2_dlygate4sd3_1 hold153 (.A(_0121_),
    .X(net542));
 sg13g2_dlygate4sd3_1 hold154 (.A(\main.demo.zic._q_squ_env[1] ),
    .X(net543));
 sg13g2_dlygate4sd3_1 hold155 (.A(_0204_),
    .X(net544));
 sg13g2_dlygate4sd3_1 hold156 (.A(\main.demo.zic._q_qpos[9] ),
    .X(net545));
 sg13g2_dlygate4sd3_1 hold157 (.A(\main.demo.zic._q_qpos[2] ),
    .X(net546));
 sg13g2_dlygate4sd3_1 hold158 (.A(\main.demo.zic._q_qpos[4] ),
    .X(net547));
 sg13g2_dlygate4sd3_1 hold159 (.A(\main.demo.vga._q_ycount[7] ),
    .X(net548));
 sg13g2_dlygate4sd3_1 hold160 (.A(_0200_),
    .X(net549));
 sg13g2_dlygate4sd3_1 hold161 (.A(\main.demo.zic._q_drum_inc[2] ),
    .X(net550));
 sg13g2_dlygate4sd3_1 hold162 (.A(_0006_),
    .X(net551));
 sg13g2_dlygate4sd3_1 hold163 (.A(\main.demo._t___pip_58_1_3___block_87_atten_h[1] ),
    .X(net552));
 sg13g2_dlygate4sd3_1 hold164 (.A(\main.demo.vga._q_active_v ),
    .X(net553));
 sg13g2_dlygate4sd3_1 hold165 (.A(\main.demo.zic._q_squ_env[5] ),
    .X(net554));
 sg13g2_dlygate4sd3_1 hold166 (.A(_2521_),
    .X(net555));
 sg13g2_dlygate4sd3_1 hold167 (.A(_0037_),
    .X(net556));
 sg13g2_dlygate4sd3_1 hold168 (.A(\main.demo.zic._q_squ_env[2] ),
    .X(net557));
 sg13g2_dlygate4sd3_1 hold169 (.A(\main.demo.zic._q_tpos[6] ),
    .X(net558));
 sg13g2_dlygate4sd3_1 hold170 (.A(rst_n_q),
    .X(net559));
 sg13g2_dlygate4sd3_1 hold171 (.A(net444),
    .X(net560));
 sg13g2_dlygate4sd3_1 hold172 (.A(\main.demo.vga._q_ycount[4] ),
    .X(net561));
 sg13g2_dlygate4sd3_1 hold173 (.A(\main.demo._d___pip_58_1_3___stage___block_3_cx[3] ),
    .X(net562));
 sg13g2_dlygate4sd3_1 hold174 (.A(\main.demo._d___pip_58_1_3___stage___block_3_cx[5] ),
    .X(net563));
 sg13g2_dlygate4sd3_1 hold175 (.A(\main.demo.zic._q_qpos[6] ),
    .X(net564));
 sg13g2_dlygate4sd3_1 hold176 (.A(_0113_),
    .X(net565));
 sg13g2_dlygate4sd3_1 hold177 (.A(\main.demo.zic._q_squ_env[0] ),
    .X(net566));
 sg13g2_dlygate4sd3_1 hold178 (.A(\main.demo.zic._q_drum_inc[3] ),
    .X(net567));
 sg13g2_dlygate4sd3_1 hold179 (.A(\main.demo._q_speed[4] ),
    .X(net568));
 sg13g2_dlygate4sd3_1 hold180 (.A(_0080_),
    .X(net569));
 sg13g2_dlygate4sd3_1 hold181 (.A(\main.demo._q_speed[14] ),
    .X(net570));
 sg13g2_dlygate4sd3_1 hold182 (.A(_2201_),
    .X(net571));
 sg13g2_dlygate4sd3_1 hold183 (.A(_0090_),
    .X(net572));
 sg13g2_dlygate4sd3_1 hold184 (.A(\main.demo._q_th[2] ),
    .X(net573));
 sg13g2_dlygate4sd3_1 hold185 (.A(_2364_),
    .X(net574));
 sg13g2_dlygate4sd3_1 hold186 (.A(\main.demo._q_speed[0] ),
    .X(net575));
 sg13g2_dlygate4sd3_1 hold187 (.A(_0076_),
    .X(net576));
 sg13g2_dlygate4sd3_1 hold188 (.A(\main.demo.zic._q_clock_count[0] ),
    .X(net577));
 sg13g2_dlygate4sd3_1 hold189 (.A(_2208_),
    .X(net578));
 sg13g2_dlygate4sd3_1 hold190 (.A(_0210_),
    .X(net579));
 sg13g2_dlygate4sd3_1 hold191 (.A(\main.demo._d___pip_58_1_3___stage___block_3_cx[1] ),
    .X(net580));
 sg13g2_dlygate4sd3_1 hold192 (.A(\main.demo._q_speed[13] ),
    .X(net581));
 sg13g2_dlygate4sd3_1 hold193 (.A(_2195_),
    .X(net582));
 sg13g2_dlygate4sd3_1 hold194 (.A(\main.demo._q_speed[10] ),
    .X(net583));
 sg13g2_dlygate4sd3_1 hold195 (.A(_0086_),
    .X(net584));
 sg13g2_dlygate4sd3_1 hold196 (.A(_0024_),
    .X(net585));
 sg13g2_dlygate4sd3_1 hold197 (.A(_2519_),
    .X(net586));
 sg13g2_dlygate4sd3_1 hold198 (.A(\main.demo._t___stage___block_3_y[2] ),
    .X(net587));
 sg13g2_dlygate4sd3_1 hold199 (.A(\main.demo._t___pip_58_1_0___stage___block_3_cx[2] ),
    .X(net588));
 sg13g2_dlygate4sd3_1 hold200 (.A(\main.demo.zic._q_idx[6] ),
    .X(net589));
 sg13g2_dlygate4sd3_1 hold201 (.A(_2390_),
    .X(net590));
 sg13g2_dlygate4sd3_1 hold202 (.A(\main.demo._q_speed[9] ),
    .X(net591));
 sg13g2_dlygate4sd3_1 hold203 (.A(\main.demo._q_speed[12] ),
    .X(net592));
 sg13g2_dlygate4sd3_1 hold204 (.A(_2190_),
    .X(net593));
 sg13g2_dlygate4sd3_1 hold205 (.A(\main.demo._q_speed[5] ),
    .X(net594));
 sg13g2_dlygate4sd3_1 hold206 (.A(\main.demo._q_frame[14] ),
    .X(net595));
 sg13g2_dlygate4sd3_1 hold207 (.A(_2203_),
    .X(net596));
 sg13g2_dlygate4sd3_1 hold208 (.A(\main.demo._q_speed[11] ),
    .X(net597));
 sg13g2_dlygate4sd3_1 hold209 (.A(_2184_),
    .X(net598));
 sg13g2_dlygate4sd3_1 hold210 (.A(_0087_),
    .X(net599));
 sg13g2_dlygate4sd3_1 hold211 (.A(_0004_),
    .X(net600));
 sg13g2_dlygate4sd3_1 hold212 (.A(\main.demo._t___pip_58_1_0___stage___block_3_cx[0] ),
    .X(net601));
 sg13g2_dlygate4sd3_1 hold213 (.A(\main.demo._q_frame[4] ),
    .X(net602));
 sg13g2_dlygate4sd3_1 hold214 (.A(_2146_),
    .X(net603));
 sg13g2_dlygate4sd3_1 hold215 (.A(\main.demo._q_frame[11] ),
    .X(net604));
 sg13g2_dlygate4sd3_1 hold216 (.A(_2187_),
    .X(net605));
 sg13g2_dlygate4sd3_1 hold217 (.A(\main.demo.zic._q_tpos[4] ),
    .X(net606));
 sg13g2_dlygate4sd3_1 hold218 (.A(\main.demo.zic._q_drum_inc[1] ),
    .X(net607));
 sg13g2_dlygate4sd3_1 hold219 (.A(\main.demo._q_th[3] ),
    .X(net608));
 sg13g2_dlygate4sd3_1 hold220 (.A(\main.demo._q_frame[8] ),
    .X(net609));
 sg13g2_dlygate4sd3_1 hold221 (.A(\main.demo._q_speed[3] ),
    .X(net610));
 sg13g2_dlygate4sd3_1 hold222 (.A(\main.demo._t___stage___block_3_x[0] ),
    .X(net611));
 sg13g2_dlygate4sd3_1 hold223 (.A(\main.demo.zic._q_drum_inc[0] ),
    .X(net612));
 sg13g2_dlygate4sd3_1 hold224 (.A(\main.demo._q_frame[13] ),
    .X(net613));
 sg13g2_dlygate4sd3_1 hold225 (.A(_2200_),
    .X(net614));
 sg13g2_dlygate4sd3_1 hold226 (.A(\main.demo.vga._q_ycount[8] ),
    .X(net615));
 sg13g2_dlygate4sd3_1 hold227 (.A(_2107_),
    .X(net616));
 sg13g2_dlygate4sd3_1 hold228 (.A(_2109_),
    .X(net617));
 sg13g2_dlygate4sd3_1 hold229 (.A(_0075_),
    .X(net618));
 sg13g2_dlygate4sd3_1 hold230 (.A(_0036_),
    .X(net619));
 sg13g2_dlygate4sd3_1 hold231 (.A(\main.demo.vga._q_ycount[7] ),
    .X(net620));
 sg13g2_dlygate4sd3_1 hold232 (.A(_0236_),
    .X(net621));
 sg13g2_dlygate4sd3_1 hold233 (.A(\main.demo._q_speed[8] ),
    .X(net622));
 sg13g2_dlygate4sd3_1 hold234 (.A(\main.demo._q_speed[1] ),
    .X(net623));
 sg13g2_dlygate4sd3_1 hold235 (.A(\main.demo._q_frame[10] ),
    .X(net624));
 sg13g2_dlygate4sd3_1 hold236 (.A(\main.demo.vga._q_ycount[1] ),
    .X(net625));
 sg13g2_dlygate4sd3_1 hold237 (.A(_2101_),
    .X(net626));
 sg13g2_dlygate4sd3_1 hold238 (.A(\main.demo._q_speed[6] ),
    .X(net627));
 sg13g2_dlygate4sd3_1 hold239 (.A(\main.demo._q_frame[12] ),
    .X(net628));
 sg13g2_dlygate4sd3_1 hold240 (.A(_2194_),
    .X(net629));
 sg13g2_dlygate4sd3_1 hold241 (.A(\main.demo._q_frame[9] ),
    .X(net630));
 sg13g2_dlygate4sd3_1 hold242 (.A(\main.demo._q___pip_58_1_1___stage___block_3_cx[10] ),
    .X(net631));
 sg13g2_dlygate4sd3_1 hold243 (.A(_0003_),
    .X(net632));
 sg13g2_dlygate4sd3_1 hold244 (.A(\main.demo._q_frame[0] ),
    .X(net633));
 sg13g2_dlygate4sd3_1 hold245 (.A(\main.demo._q_frame[8] ),
    .X(net634));
 sg13g2_dlygate4sd3_1 hold246 (.A(\main.demo.zic._q_squ_env[3] ),
    .X(net635));
 sg13g2_dlygate4sd3_1 hold247 (.A(\main.demo._q_go ),
    .X(net636));
 sg13g2_dlygate4sd3_1 hold248 (.A(\main.demo._q_frame[5] ),
    .X(net637));
 sg13g2_dlygate4sd3_1 hold249 (.A(\main.demo.zic._q_idx[2] ),
    .X(net638));
 sg13g2_dlygate4sd3_1 hold250 (.A(\main.demo._q_effect[1] ),
    .X(net639));
 sg13g2_dlygate4sd3_1 hold251 (.A(\main.demo.zic._q_idx[1] ),
    .X(net640));
 sg13g2_dlygate4sd3_1 hold252 (.A(\main.demo._q_speed[2] ),
    .X(net641));
 sg13g2_dlygate4sd3_1 hold253 (.A(\main.demo._q_speed[7] ),
    .X(net642));
 sg13g2_dlygate4sd3_1 hold254 (.A(_0001_),
    .X(net643));
 sg13g2_dlygate4sd3_1 hold255 (.A(\main.demo.zic._q_drum_inc[1] ),
    .X(net644));
 sg13g2_dlygate4sd3_1 hold256 (.A(\main.demo.vga._q_ycount[1] ),
    .X(net645));
 sg13g2_antennanp ANTENNA_1 (.A(clk));
 sg13g2_antennanp ANTENNA_2 (.A(clk));
 sg13g2_fill_2 FILLER_0_40 ();
 sg13g2_fill_1 FILLER_0_42 ();
 sg13g2_fill_2 FILLER_0_58 ();
 sg13g2_fill_1 FILLER_0_69 ();
 sg13g2_decap_8 FILLER_0_86 ();
 sg13g2_decap_8 FILLER_0_93 ();
 sg13g2_decap_8 FILLER_0_100 ();
 sg13g2_decap_8 FILLER_0_107 ();
 sg13g2_decap_8 FILLER_0_114 ();
 sg13g2_decap_8 FILLER_0_121 ();
 sg13g2_decap_8 FILLER_0_128 ();
 sg13g2_decap_8 FILLER_0_135 ();
 sg13g2_decap_8 FILLER_0_142 ();
 sg13g2_decap_4 FILLER_0_149 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_187 ();
 sg13g2_decap_4 FILLER_0_194 ();
 sg13g2_fill_2 FILLER_0_198 ();
 sg13g2_decap_8 FILLER_0_205 ();
 sg13g2_decap_8 FILLER_0_212 ();
 sg13g2_decap_8 FILLER_0_219 ();
 sg13g2_fill_1 FILLER_0_226 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_4 FILLER_0_238 ();
 sg13g2_fill_1 FILLER_0_242 ();
 sg13g2_fill_2 FILLER_0_247 ();
 sg13g2_fill_1 FILLER_0_249 ();
 sg13g2_decap_8 FILLER_0_255 ();
 sg13g2_decap_8 FILLER_0_262 ();
 sg13g2_decap_8 FILLER_0_269 ();
 sg13g2_decap_8 FILLER_0_276 ();
 sg13g2_decap_8 FILLER_0_283 ();
 sg13g2_decap_8 FILLER_0_290 ();
 sg13g2_decap_8 FILLER_0_297 ();
 sg13g2_fill_2 FILLER_0_304 ();
 sg13g2_decap_8 FILLER_0_310 ();
 sg13g2_decap_4 FILLER_0_317 ();
 sg13g2_fill_2 FILLER_0_321 ();
 sg13g2_decap_8 FILLER_0_327 ();
 sg13g2_decap_8 FILLER_0_334 ();
 sg13g2_fill_2 FILLER_0_341 ();
 sg13g2_fill_1 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_351 ();
 sg13g2_decap_4 FILLER_0_358 ();
 sg13g2_fill_2 FILLER_0_362 ();
 sg13g2_decap_8 FILLER_0_376 ();
 sg13g2_decap_8 FILLER_0_383 ();
 sg13g2_decap_8 FILLER_0_390 ();
 sg13g2_decap_8 FILLER_0_397 ();
 sg13g2_decap_4 FILLER_0_404 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_fill_2 FILLER_1_74 ();
 sg13g2_fill_2 FILLER_1_80 ();
 sg13g2_fill_1 FILLER_1_82 ();
 sg13g2_fill_1 FILLER_1_87 ();
 sg13g2_fill_2 FILLER_1_96 ();
 sg13g2_fill_1 FILLER_1_98 ();
 sg13g2_decap_4 FILLER_1_109 ();
 sg13g2_fill_2 FILLER_1_199 ();
 sg13g2_fill_1 FILLER_1_206 ();
 sg13g2_fill_1 FILLER_1_215 ();
 sg13g2_fill_2 FILLER_1_237 ();
 sg13g2_fill_1 FILLER_1_253 ();
 sg13g2_fill_1 FILLER_1_270 ();
 sg13g2_fill_1 FILLER_1_372 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_fill_1 FILLER_2_0 ();
 sg13g2_fill_2 FILLER_2_215 ();
 sg13g2_fill_1 FILLER_2_217 ();
 sg13g2_fill_1 FILLER_2_226 ();
 sg13g2_fill_1 FILLER_2_337 ();
 sg13g2_fill_2 FILLER_2_343 ();
 sg13g2_fill_2 FILLER_2_376 ();
 sg13g2_decap_8 FILLER_2_400 ();
 sg13g2_fill_2 FILLER_2_407 ();
 sg13g2_fill_1 FILLER_3_0 ();
 sg13g2_fill_1 FILLER_3_70 ();
 sg13g2_fill_2 FILLER_3_93 ();
 sg13g2_fill_2 FILLER_3_147 ();
 sg13g2_fill_1 FILLER_3_149 ();
 sg13g2_fill_1 FILLER_3_199 ();
 sg13g2_fill_1 FILLER_3_216 ();
 sg13g2_fill_1 FILLER_3_242 ();
 sg13g2_fill_1 FILLER_3_335 ();
 sg13g2_fill_1 FILLER_3_349 ();
 sg13g2_fill_2 FILLER_3_363 ();
 sg13g2_fill_1 FILLER_3_365 ();
 sg13g2_decap_4 FILLER_3_404 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_fill_2 FILLER_4_0 ();
 sg13g2_fill_1 FILLER_4_53 ();
 sg13g2_decap_4 FILLER_4_121 ();
 sg13g2_fill_1 FILLER_4_134 ();
 sg13g2_decap_8 FILLER_4_143 ();
 sg13g2_fill_2 FILLER_4_150 ();
 sg13g2_fill_1 FILLER_4_152 ();
 sg13g2_fill_1 FILLER_4_170 ();
 sg13g2_fill_2 FILLER_4_195 ();
 sg13g2_decap_8 FILLER_4_202 ();
 sg13g2_decap_8 FILLER_4_209 ();
 sg13g2_decap_4 FILLER_4_228 ();
 sg13g2_fill_1 FILLER_4_232 ();
 sg13g2_fill_2 FILLER_4_238 ();
 sg13g2_fill_1 FILLER_4_240 ();
 sg13g2_fill_1 FILLER_4_251 ();
 sg13g2_fill_2 FILLER_4_259 ();
 sg13g2_fill_1 FILLER_4_318 ();
 sg13g2_decap_8 FILLER_4_400 ();
 sg13g2_fill_2 FILLER_4_407 ();
 sg13g2_fill_1 FILLER_5_0 ();
 sg13g2_fill_1 FILLER_5_55 ();
 sg13g2_fill_2 FILLER_5_95 ();
 sg13g2_fill_1 FILLER_5_107 ();
 sg13g2_decap_4 FILLER_5_112 ();
 sg13g2_fill_2 FILLER_5_116 ();
 sg13g2_decap_8 FILLER_5_144 ();
 sg13g2_fill_2 FILLER_5_151 ();
 sg13g2_fill_2 FILLER_5_166 ();
 sg13g2_decap_4 FILLER_5_187 ();
 sg13g2_fill_1 FILLER_5_191 ();
 sg13g2_decap_8 FILLER_5_201 ();
 sg13g2_decap_8 FILLER_5_208 ();
 sg13g2_fill_2 FILLER_5_215 ();
 sg13g2_fill_1 FILLER_5_217 ();
 sg13g2_fill_1 FILLER_5_225 ();
 sg13g2_decap_4 FILLER_5_236 ();
 sg13g2_fill_1 FILLER_5_240 ();
 sg13g2_fill_2 FILLER_5_258 ();
 sg13g2_fill_1 FILLER_5_260 ();
 sg13g2_decap_8 FILLER_5_304 ();
 sg13g2_decap_8 FILLER_5_311 ();
 sg13g2_decap_4 FILLER_5_318 ();
 sg13g2_fill_1 FILLER_5_322 ();
 sg13g2_fill_2 FILLER_5_326 ();
 sg13g2_fill_2 FILLER_5_348 ();
 sg13g2_fill_1 FILLER_5_380 ();
 sg13g2_fill_2 FILLER_5_386 ();
 sg13g2_fill_1 FILLER_5_388 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_fill_2 FILLER_6_100 ();
 sg13g2_decap_8 FILLER_6_111 ();
 sg13g2_fill_2 FILLER_6_118 ();
 sg13g2_fill_2 FILLER_6_178 ();
 sg13g2_fill_1 FILLER_6_180 ();
 sg13g2_fill_1 FILLER_6_186 ();
 sg13g2_fill_2 FILLER_6_195 ();
 sg13g2_decap_4 FILLER_6_210 ();
 sg13g2_fill_1 FILLER_6_214 ();
 sg13g2_fill_2 FILLER_6_251 ();
 sg13g2_fill_2 FILLER_6_261 ();
 sg13g2_fill_1 FILLER_6_263 ();
 sg13g2_decap_8 FILLER_6_272 ();
 sg13g2_decap_8 FILLER_6_279 ();
 sg13g2_fill_2 FILLER_6_286 ();
 sg13g2_fill_1 FILLER_6_288 ();
 sg13g2_fill_2 FILLER_6_307 ();
 sg13g2_fill_1 FILLER_6_309 ();
 sg13g2_fill_1 FILLER_6_317 ();
 sg13g2_decap_4 FILLER_6_346 ();
 sg13g2_fill_2 FILLER_6_354 ();
 sg13g2_decap_8 FILLER_6_360 ();
 sg13g2_fill_2 FILLER_6_367 ();
 sg13g2_decap_4 FILLER_6_377 ();
 sg13g2_fill_2 FILLER_6_381 ();
 sg13g2_fill_1 FILLER_7_50 ();
 sg13g2_fill_2 FILLER_7_89 ();
 sg13g2_fill_1 FILLER_7_91 ();
 sg13g2_fill_1 FILLER_7_125 ();
 sg13g2_fill_2 FILLER_7_165 ();
 sg13g2_fill_1 FILLER_7_172 ();
 sg13g2_decap_4 FILLER_7_215 ();
 sg13g2_fill_2 FILLER_7_219 ();
 sg13g2_decap_4 FILLER_7_239 ();
 sg13g2_decap_8 FILLER_7_251 ();
 sg13g2_decap_4 FILLER_7_258 ();
 sg13g2_decap_4 FILLER_7_282 ();
 sg13g2_fill_2 FILLER_7_286 ();
 sg13g2_decap_8 FILLER_7_291 ();
 sg13g2_fill_2 FILLER_7_298 ();
 sg13g2_fill_1 FILLER_7_300 ();
 sg13g2_fill_2 FILLER_7_309 ();
 sg13g2_decap_8 FILLER_7_337 ();
 sg13g2_decap_4 FILLER_7_344 ();
 sg13g2_decap_8 FILLER_7_353 ();
 sg13g2_fill_1 FILLER_7_360 ();
 sg13g2_fill_2 FILLER_7_378 ();
 sg13g2_fill_1 FILLER_7_380 ();
 sg13g2_fill_1 FILLER_7_394 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_fill_2 FILLER_8_26 ();
 sg13g2_fill_2 FILLER_8_66 ();
 sg13g2_fill_1 FILLER_8_114 ();
 sg13g2_fill_2 FILLER_8_128 ();
 sg13g2_fill_1 FILLER_8_130 ();
 sg13g2_fill_1 FILLER_8_139 ();
 sg13g2_fill_1 FILLER_8_149 ();
 sg13g2_decap_8 FILLER_8_173 ();
 sg13g2_fill_1 FILLER_8_180 ();
 sg13g2_fill_2 FILLER_8_224 ();
 sg13g2_fill_1 FILLER_8_226 ();
 sg13g2_fill_2 FILLER_8_230 ();
 sg13g2_fill_1 FILLER_8_232 ();
 sg13g2_fill_1 FILLER_8_238 ();
 sg13g2_fill_2 FILLER_8_262 ();
 sg13g2_fill_2 FILLER_8_303 ();
 sg13g2_fill_2 FILLER_8_313 ();
 sg13g2_fill_2 FILLER_8_331 ();
 sg13g2_fill_2 FILLER_8_344 ();
 sg13g2_decap_4 FILLER_8_359 ();
 sg13g2_fill_2 FILLER_8_363 ();
 sg13g2_decap_8 FILLER_8_382 ();
 sg13g2_decap_4 FILLER_8_389 ();
 sg13g2_decap_4 FILLER_8_405 ();
 sg13g2_fill_2 FILLER_9_0 ();
 sg13g2_fill_1 FILLER_9_2 ();
 sg13g2_fill_1 FILLER_9_72 ();
 sg13g2_fill_2 FILLER_9_87 ();
 sg13g2_fill_1 FILLER_9_89 ();
 sg13g2_fill_2 FILLER_9_122 ();
 sg13g2_fill_1 FILLER_9_124 ();
 sg13g2_decap_8 FILLER_9_151 ();
 sg13g2_decap_8 FILLER_9_158 ();
 sg13g2_fill_2 FILLER_9_177 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_fill_2 FILLER_9_224 ();
 sg13g2_fill_2 FILLER_9_250 ();
 sg13g2_decap_4 FILLER_9_314 ();
 sg13g2_fill_1 FILLER_9_326 ();
 sg13g2_fill_1 FILLER_9_335 ();
 sg13g2_decap_4 FILLER_9_383 ();
 sg13g2_decap_8 FILLER_9_400 ();
 sg13g2_fill_2 FILLER_9_407 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_fill_2 FILLER_10_14 ();
 sg13g2_fill_2 FILLER_10_43 ();
 sg13g2_fill_2 FILLER_10_59 ();
 sg13g2_fill_1 FILLER_10_61 ();
 sg13g2_fill_2 FILLER_10_87 ();
 sg13g2_fill_1 FILLER_10_108 ();
 sg13g2_decap_4 FILLER_10_118 ();
 sg13g2_fill_1 FILLER_10_122 ();
 sg13g2_decap_8 FILLER_10_128 ();
 sg13g2_fill_2 FILLER_10_135 ();
 sg13g2_fill_2 FILLER_10_181 ();
 sg13g2_fill_1 FILLER_10_188 ();
 sg13g2_decap_8 FILLER_10_197 ();
 sg13g2_fill_2 FILLER_10_204 ();
 sg13g2_fill_1 FILLER_10_227 ();
 sg13g2_fill_2 FILLER_10_244 ();
 sg13g2_fill_1 FILLER_10_258 ();
 sg13g2_fill_2 FILLER_10_277 ();
 sg13g2_fill_1 FILLER_10_279 ();
 sg13g2_fill_2 FILLER_10_318 ();
 sg13g2_fill_1 FILLER_10_320 ();
 sg13g2_fill_1 FILLER_10_341 ();
 sg13g2_fill_1 FILLER_10_351 ();
 sg13g2_fill_2 FILLER_10_357 ();
 sg13g2_fill_2 FILLER_10_368 ();
 sg13g2_decap_4 FILLER_10_375 ();
 sg13g2_decap_4 FILLER_11_26 ();
 sg13g2_fill_2 FILLER_11_30 ();
 sg13g2_fill_1 FILLER_11_36 ();
 sg13g2_fill_2 FILLER_11_133 ();
 sg13g2_fill_1 FILLER_11_135 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_fill_1 FILLER_11_147 ();
 sg13g2_fill_2 FILLER_11_152 ();
 sg13g2_fill_1 FILLER_11_154 ();
 sg13g2_decap_4 FILLER_11_159 ();
 sg13g2_fill_1 FILLER_11_163 ();
 sg13g2_fill_2 FILLER_11_168 ();
 sg13g2_fill_1 FILLER_11_170 ();
 sg13g2_fill_2 FILLER_11_176 ();
 sg13g2_fill_1 FILLER_11_178 ();
 sg13g2_decap_8 FILLER_11_236 ();
 sg13g2_fill_1 FILLER_11_243 ();
 sg13g2_decap_8 FILLER_11_251 ();
 sg13g2_decap_8 FILLER_11_258 ();
 sg13g2_decap_4 FILLER_11_265 ();
 sg13g2_decap_8 FILLER_11_278 ();
 sg13g2_fill_1 FILLER_11_285 ();
 sg13g2_fill_2 FILLER_11_295 ();
 sg13g2_fill_1 FILLER_11_297 ();
 sg13g2_fill_1 FILLER_11_328 ();
 sg13g2_decap_4 FILLER_11_355 ();
 sg13g2_fill_2 FILLER_11_359 ();
 sg13g2_fill_1 FILLER_11_374 ();
 sg13g2_decap_4 FILLER_12_38 ();
 sg13g2_fill_2 FILLER_12_42 ();
 sg13g2_fill_1 FILLER_12_108 ();
 sg13g2_decap_4 FILLER_12_125 ();
 sg13g2_decap_8 FILLER_12_134 ();
 sg13g2_fill_2 FILLER_12_141 ();
 sg13g2_fill_1 FILLER_12_143 ();
 sg13g2_fill_1 FILLER_12_188 ();
 sg13g2_fill_2 FILLER_12_197 ();
 sg13g2_fill_1 FILLER_12_199 ();
 sg13g2_decap_4 FILLER_12_212 ();
 sg13g2_decap_8 FILLER_12_219 ();
 sg13g2_decap_4 FILLER_12_230 ();
 sg13g2_fill_2 FILLER_12_234 ();
 sg13g2_decap_8 FILLER_12_263 ();
 sg13g2_fill_2 FILLER_12_270 ();
 sg13g2_decap_4 FILLER_12_302 ();
 sg13g2_decap_8 FILLER_12_310 ();
 sg13g2_decap_8 FILLER_12_321 ();
 sg13g2_decap_8 FILLER_12_328 ();
 sg13g2_decap_4 FILLER_12_335 ();
 sg13g2_fill_1 FILLER_12_339 ();
 sg13g2_decap_8 FILLER_12_344 ();
 sg13g2_fill_1 FILLER_12_358 ();
 sg13g2_fill_1 FILLER_12_369 ();
 sg13g2_fill_2 FILLER_12_386 ();
 sg13g2_fill_1 FILLER_12_388 ();
 sg13g2_fill_2 FILLER_13_0 ();
 sg13g2_fill_2 FILLER_13_20 ();
 sg13g2_fill_1 FILLER_13_53 ();
 sg13g2_fill_2 FILLER_13_58 ();
 sg13g2_fill_2 FILLER_13_77 ();
 sg13g2_fill_1 FILLER_13_79 ();
 sg13g2_fill_2 FILLER_13_99 ();
 sg13g2_fill_1 FILLER_13_101 ();
 sg13g2_fill_2 FILLER_13_110 ();
 sg13g2_fill_2 FILLER_13_117 ();
 sg13g2_fill_1 FILLER_13_161 ();
 sg13g2_fill_1 FILLER_13_182 ();
 sg13g2_fill_2 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_4 FILLER_13_210 ();
 sg13g2_fill_1 FILLER_13_214 ();
 sg13g2_fill_2 FILLER_13_235 ();
 sg13g2_decap_4 FILLER_13_269 ();
 sg13g2_fill_2 FILLER_13_273 ();
 sg13g2_fill_1 FILLER_13_292 ();
 sg13g2_decap_8 FILLER_13_330 ();
 sg13g2_fill_2 FILLER_13_337 ();
 sg13g2_fill_1 FILLER_13_372 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_fill_1 FILLER_14_0 ();
 sg13g2_fill_2 FILLER_14_10 ();
 sg13g2_fill_1 FILLER_14_103 ();
 sg13g2_decap_8 FILLER_14_135 ();
 sg13g2_decap_4 FILLER_14_142 ();
 sg13g2_fill_2 FILLER_14_150 ();
 sg13g2_fill_2 FILLER_14_178 ();
 sg13g2_fill_1 FILLER_14_185 ();
 sg13g2_decap_8 FILLER_14_194 ();
 sg13g2_fill_2 FILLER_14_209 ();
 sg13g2_decap_4 FILLER_14_234 ();
 sg13g2_fill_2 FILLER_14_243 ();
 sg13g2_decap_4 FILLER_14_261 ();
 sg13g2_fill_1 FILLER_14_320 ();
 sg13g2_fill_2 FILLER_14_332 ();
 sg13g2_fill_2 FILLER_14_345 ();
 sg13g2_fill_1 FILLER_14_347 ();
 sg13g2_decap_8 FILLER_14_353 ();
 sg13g2_decap_4 FILLER_14_360 ();
 sg13g2_fill_1 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_370 ();
 sg13g2_fill_2 FILLER_14_377 ();
 sg13g2_fill_1 FILLER_14_379 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_4 FILLER_14_392 ();
 sg13g2_fill_1 FILLER_14_396 ();
 sg13g2_fill_2 FILLER_14_406 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_fill_1 FILLER_15_0 ();
 sg13g2_fill_2 FILLER_15_27 ();
 sg13g2_fill_1 FILLER_15_67 ();
 sg13g2_fill_1 FILLER_15_73 ();
 sg13g2_fill_2 FILLER_15_101 ();
 sg13g2_decap_8 FILLER_15_124 ();
 sg13g2_decap_4 FILLER_15_131 ();
 sg13g2_fill_2 FILLER_15_135 ();
 sg13g2_decap_8 FILLER_15_149 ();
 sg13g2_decap_8 FILLER_15_156 ();
 sg13g2_decap_8 FILLER_15_167 ();
 sg13g2_decap_8 FILLER_15_174 ();
 sg13g2_fill_2 FILLER_15_181 ();
 sg13g2_decap_4 FILLER_15_197 ();
 sg13g2_fill_2 FILLER_15_209 ();
 sg13g2_fill_1 FILLER_15_211 ();
 sg13g2_fill_1 FILLER_15_242 ();
 sg13g2_decap_4 FILLER_15_248 ();
 sg13g2_fill_1 FILLER_15_252 ();
 sg13g2_fill_1 FILLER_15_275 ();
 sg13g2_decap_4 FILLER_15_280 ();
 sg13g2_fill_2 FILLER_15_284 ();
 sg13g2_fill_2 FILLER_15_301 ();
 sg13g2_fill_1 FILLER_15_303 ();
 sg13g2_fill_1 FILLER_15_327 ();
 sg13g2_fill_2 FILLER_15_338 ();
 sg13g2_fill_1 FILLER_15_340 ();
 sg13g2_fill_2 FILLER_15_351 ();
 sg13g2_fill_2 FILLER_15_378 ();
 sg13g2_fill_1 FILLER_15_380 ();
 sg13g2_fill_2 FILLER_15_386 ();
 sg13g2_fill_1 FILLER_15_388 ();
 sg13g2_fill_2 FILLER_16_44 ();
 sg13g2_fill_2 FILLER_16_56 ();
 sg13g2_fill_1 FILLER_16_58 ();
 sg13g2_fill_2 FILLER_16_109 ();
 sg13g2_fill_1 FILLER_16_111 ();
 sg13g2_fill_2 FILLER_16_116 ();
 sg13g2_fill_2 FILLER_16_130 ();
 sg13g2_fill_1 FILLER_16_132 ();
 sg13g2_fill_2 FILLER_16_228 ();
 sg13g2_fill_2 FILLER_16_253 ();
 sg13g2_decap_8 FILLER_16_276 ();
 sg13g2_decap_4 FILLER_16_283 ();
 sg13g2_fill_2 FILLER_16_287 ();
 sg13g2_fill_2 FILLER_16_294 ();
 sg13g2_fill_2 FILLER_16_314 ();
 sg13g2_fill_1 FILLER_16_316 ();
 sg13g2_fill_1 FILLER_16_323 ();
 sg13g2_fill_2 FILLER_16_347 ();
 sg13g2_fill_1 FILLER_16_349 ();
 sg13g2_decap_4 FILLER_16_383 ();
 sg13g2_fill_2 FILLER_17_15 ();
 sg13g2_fill_2 FILLER_17_40 ();
 sg13g2_fill_2 FILLER_17_62 ();
 sg13g2_fill_1 FILLER_17_64 ();
 sg13g2_fill_2 FILLER_17_83 ();
 sg13g2_fill_1 FILLER_17_85 ();
 sg13g2_decap_8 FILLER_17_90 ();
 sg13g2_decap_8 FILLER_17_97 ();
 sg13g2_fill_1 FILLER_17_128 ();
 sg13g2_decap_8 FILLER_17_145 ();
 sg13g2_fill_1 FILLER_17_152 ();
 sg13g2_fill_1 FILLER_17_210 ();
 sg13g2_fill_2 FILLER_17_222 ();
 sg13g2_fill_1 FILLER_17_224 ();
 sg13g2_decap_8 FILLER_17_274 ();
 sg13g2_fill_2 FILLER_17_281 ();
 sg13g2_fill_1 FILLER_17_305 ();
 sg13g2_fill_1 FILLER_17_374 ();
 sg13g2_fill_2 FILLER_17_386 ();
 sg13g2_fill_2 FILLER_18_45 ();
 sg13g2_decap_8 FILLER_18_51 ();
 sg13g2_fill_1 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_79 ();
 sg13g2_decap_8 FILLER_18_86 ();
 sg13g2_fill_2 FILLER_18_101 ();
 sg13g2_fill_1 FILLER_18_103 ();
 sg13g2_fill_2 FILLER_18_114 ();
 sg13g2_fill_2 FILLER_18_124 ();
 sg13g2_decap_8 FILLER_18_147 ();
 sg13g2_fill_2 FILLER_18_154 ();
 sg13g2_fill_1 FILLER_18_156 ();
 sg13g2_fill_2 FILLER_18_166 ();
 sg13g2_fill_1 FILLER_18_176 ();
 sg13g2_fill_1 FILLER_18_205 ();
 sg13g2_fill_2 FILLER_18_214 ();
 sg13g2_fill_2 FILLER_18_224 ();
 sg13g2_fill_2 FILLER_18_234 ();
 sg13g2_fill_1 FILLER_18_236 ();
 sg13g2_fill_2 FILLER_18_250 ();
 sg13g2_fill_1 FILLER_18_257 ();
 sg13g2_fill_2 FILLER_18_275 ();
 sg13g2_fill_2 FILLER_18_303 ();
 sg13g2_fill_1 FILLER_18_319 ();
 sg13g2_fill_1 FILLER_18_385 ();
 sg13g2_fill_1 FILLER_18_393 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_fill_2 FILLER_19_14 ();
 sg13g2_fill_1 FILLER_19_16 ();
 sg13g2_decap_4 FILLER_19_32 ();
 sg13g2_fill_1 FILLER_19_50 ();
 sg13g2_fill_1 FILLER_19_66 ();
 sg13g2_decap_8 FILLER_19_82 ();
 sg13g2_fill_1 FILLER_19_89 ();
 sg13g2_fill_2 FILLER_19_98 ();
 sg13g2_fill_1 FILLER_19_100 ();
 sg13g2_fill_2 FILLER_19_117 ();
 sg13g2_fill_1 FILLER_19_119 ();
 sg13g2_fill_2 FILLER_19_133 ();
 sg13g2_fill_1 FILLER_19_135 ();
 sg13g2_decap_8 FILLER_19_179 ();
 sg13g2_decap_8 FILLER_19_186 ();
 sg13g2_decap_8 FILLER_19_193 ();
 sg13g2_decap_4 FILLER_19_200 ();
 sg13g2_fill_1 FILLER_19_204 ();
 sg13g2_decap_4 FILLER_19_237 ();
 sg13g2_decap_4 FILLER_19_265 ();
 sg13g2_fill_1 FILLER_19_269 ();
 sg13g2_fill_2 FILLER_19_330 ();
 sg13g2_fill_1 FILLER_19_368 ();
 sg13g2_fill_1 FILLER_19_395 ();
 sg13g2_decap_4 FILLER_20_0 ();
 sg13g2_fill_1 FILLER_20_25 ();
 sg13g2_fill_1 FILLER_20_44 ();
 sg13g2_fill_1 FILLER_20_50 ();
 sg13g2_fill_2 FILLER_20_56 ();
 sg13g2_fill_1 FILLER_20_98 ();
 sg13g2_fill_1 FILLER_20_111 ();
 sg13g2_fill_1 FILLER_20_117 ();
 sg13g2_fill_1 FILLER_20_122 ();
 sg13g2_decap_8 FILLER_20_155 ();
 sg13g2_decap_4 FILLER_20_162 ();
 sg13g2_fill_1 FILLER_20_166 ();
 sg13g2_decap_8 FILLER_20_193 ();
 sg13g2_decap_8 FILLER_20_200 ();
 sg13g2_decap_4 FILLER_20_207 ();
 sg13g2_decap_8 FILLER_20_228 ();
 sg13g2_decap_8 FILLER_20_235 ();
 sg13g2_decap_8 FILLER_20_242 ();
 sg13g2_decap_4 FILLER_20_253 ();
 sg13g2_fill_2 FILLER_20_257 ();
 sg13g2_fill_2 FILLER_20_263 ();
 sg13g2_fill_2 FILLER_20_293 ();
 sg13g2_fill_1 FILLER_20_318 ();
 sg13g2_fill_2 FILLER_20_330 ();
 sg13g2_fill_1 FILLER_20_332 ();
 sg13g2_fill_2 FILLER_20_345 ();
 sg13g2_fill_1 FILLER_20_347 ();
 sg13g2_fill_2 FILLER_20_370 ();
 sg13g2_fill_1 FILLER_20_372 ();
 sg13g2_fill_1 FILLER_20_378 ();
 sg13g2_decap_4 FILLER_20_388 ();
 sg13g2_fill_2 FILLER_20_392 ();
 sg13g2_decap_4 FILLER_20_403 ();
 sg13g2_fill_2 FILLER_20_407 ();
 sg13g2_fill_1 FILLER_21_0 ();
 sg13g2_fill_1 FILLER_21_28 ();
 sg13g2_fill_2 FILLER_21_42 ();
 sg13g2_fill_1 FILLER_21_44 ();
 sg13g2_fill_2 FILLER_21_55 ();
 sg13g2_fill_2 FILLER_21_101 ();
 sg13g2_fill_1 FILLER_21_111 ();
 sg13g2_fill_2 FILLER_21_125 ();
 sg13g2_fill_1 FILLER_21_127 ();
 sg13g2_fill_1 FILLER_21_144 ();
 sg13g2_fill_2 FILLER_21_162 ();
 sg13g2_fill_1 FILLER_21_181 ();
 sg13g2_decap_8 FILLER_21_208 ();
 sg13g2_decap_8 FILLER_21_215 ();
 sg13g2_decap_4 FILLER_21_222 ();
 sg13g2_fill_2 FILLER_21_226 ();
 sg13g2_decap_8 FILLER_21_233 ();
 sg13g2_decap_8 FILLER_21_240 ();
 sg13g2_fill_1 FILLER_21_247 ();
 sg13g2_decap_4 FILLER_21_274 ();
 sg13g2_fill_1 FILLER_21_278 ();
 sg13g2_fill_1 FILLER_21_294 ();
 sg13g2_fill_2 FILLER_21_304 ();
 sg13g2_fill_2 FILLER_21_318 ();
 sg13g2_fill_1 FILLER_21_320 ();
 sg13g2_decap_4 FILLER_21_366 ();
 sg13g2_fill_2 FILLER_21_370 ();
 sg13g2_fill_2 FILLER_21_380 ();
 sg13g2_fill_1 FILLER_21_382 ();
 sg13g2_decap_4 FILLER_21_405 ();
 sg13g2_fill_2 FILLER_22_37 ();
 sg13g2_fill_1 FILLER_22_39 ();
 sg13g2_fill_2 FILLER_22_54 ();
 sg13g2_fill_1 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_81 ();
 sg13g2_decap_8 FILLER_22_96 ();
 sg13g2_fill_1 FILLER_22_103 ();
 sg13g2_fill_1 FILLER_22_112 ();
 sg13g2_decap_4 FILLER_22_121 ();
 sg13g2_fill_2 FILLER_22_125 ();
 sg13g2_decap_8 FILLER_22_248 ();
 sg13g2_decap_8 FILLER_22_255 ();
 sg13g2_decap_8 FILLER_22_262 ();
 sg13g2_decap_4 FILLER_22_269 ();
 sg13g2_fill_1 FILLER_22_273 ();
 sg13g2_fill_2 FILLER_22_298 ();
 sg13g2_fill_1 FILLER_22_313 ();
 sg13g2_fill_2 FILLER_22_328 ();
 sg13g2_fill_2 FILLER_22_345 ();
 sg13g2_fill_1 FILLER_22_347 ();
 sg13g2_fill_1 FILLER_22_365 ();
 sg13g2_fill_2 FILLER_22_384 ();
 sg13g2_fill_2 FILLER_22_407 ();
 sg13g2_fill_1 FILLER_23_0 ();
 sg13g2_fill_1 FILLER_23_19 ();
 sg13g2_fill_2 FILLER_23_50 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_4 FILLER_23_77 ();
 sg13g2_fill_2 FILLER_23_81 ();
 sg13g2_fill_2 FILLER_23_103 ();
 sg13g2_decap_8 FILLER_23_110 ();
 sg13g2_decap_4 FILLER_23_117 ();
 sg13g2_decap_8 FILLER_23_129 ();
 sg13g2_fill_2 FILLER_23_136 ();
 sg13g2_fill_1 FILLER_23_138 ();
 sg13g2_fill_1 FILLER_23_147 ();
 sg13g2_fill_2 FILLER_23_165 ();
 sg13g2_decap_4 FILLER_23_265 ();
 sg13g2_fill_2 FILLER_23_269 ();
 sg13g2_fill_1 FILLER_23_298 ();
 sg13g2_fill_2 FILLER_23_314 ();
 sg13g2_fill_1 FILLER_23_339 ();
 sg13g2_fill_2 FILLER_23_353 ();
 sg13g2_fill_1 FILLER_23_386 ();
 sg13g2_fill_2 FILLER_23_407 ();
 sg13g2_decap_4 FILLER_24_0 ();
 sg13g2_fill_1 FILLER_24_4 ();
 sg13g2_decap_4 FILLER_24_28 ();
 sg13g2_fill_2 FILLER_24_56 ();
 sg13g2_decap_4 FILLER_24_70 ();
 sg13g2_fill_2 FILLER_24_74 ();
 sg13g2_fill_2 FILLER_24_140 ();
 sg13g2_fill_1 FILLER_24_142 ();
 sg13g2_decap_8 FILLER_24_151 ();
 sg13g2_decap_8 FILLER_24_158 ();
 sg13g2_fill_2 FILLER_24_165 ();
 sg13g2_fill_1 FILLER_24_167 ();
 sg13g2_fill_1 FILLER_24_176 ();
 sg13g2_decap_8 FILLER_24_181 ();
 sg13g2_decap_8 FILLER_24_188 ();
 sg13g2_fill_1 FILLER_24_195 ();
 sg13g2_decap_4 FILLER_24_200 ();
 sg13g2_fill_2 FILLER_24_230 ();
 sg13g2_fill_1 FILLER_24_232 ();
 sg13g2_decap_4 FILLER_24_237 ();
 sg13g2_fill_2 FILLER_24_241 ();
 sg13g2_fill_2 FILLER_24_296 ();
 sg13g2_fill_1 FILLER_24_298 ();
 sg13g2_fill_2 FILLER_24_308 ();
 sg13g2_fill_2 FILLER_24_338 ();
 sg13g2_fill_2 FILLER_24_349 ();
 sg13g2_fill_1 FILLER_24_351 ();
 sg13g2_fill_2 FILLER_24_392 ();
 sg13g2_fill_1 FILLER_24_394 ();
 sg13g2_fill_2 FILLER_24_407 ();
 sg13g2_decap_4 FILLER_25_0 ();
 sg13g2_fill_1 FILLER_25_4 ();
 sg13g2_fill_2 FILLER_25_21 ();
 sg13g2_fill_2 FILLER_25_46 ();
 sg13g2_decap_8 FILLER_25_66 ();
 sg13g2_decap_4 FILLER_25_78 ();
 sg13g2_decap_8 FILLER_25_107 ();
 sg13g2_fill_1 FILLER_25_129 ();
 sg13g2_decap_8 FILLER_25_151 ();
 sg13g2_decap_4 FILLER_25_158 ();
 sg13g2_fill_2 FILLER_25_162 ();
 sg13g2_decap_4 FILLER_25_210 ();
 sg13g2_fill_1 FILLER_25_214 ();
 sg13g2_decap_8 FILLER_25_219 ();
 sg13g2_fill_2 FILLER_25_226 ();
 sg13g2_decap_4 FILLER_25_246 ();
 sg13g2_fill_2 FILLER_25_284 ();
 sg13g2_fill_1 FILLER_25_286 ();
 sg13g2_fill_2 FILLER_25_325 ();
 sg13g2_fill_1 FILLER_25_339 ();
 sg13g2_decap_4 FILLER_25_381 ();
 sg13g2_fill_1 FILLER_25_394 ();
 sg13g2_fill_2 FILLER_26_0 ();
 sg13g2_fill_1 FILLER_26_89 ();
 sg13g2_fill_2 FILLER_26_101 ();
 sg13g2_decap_8 FILLER_26_107 ();
 sg13g2_decap_8 FILLER_26_114 ();
 sg13g2_decap_8 FILLER_26_121 ();
 sg13g2_fill_2 FILLER_26_140 ();
 sg13g2_fill_1 FILLER_26_186 ();
 sg13g2_decap_4 FILLER_26_213 ();
 sg13g2_fill_1 FILLER_26_217 ();
 sg13g2_decap_4 FILLER_26_223 ();
 sg13g2_fill_1 FILLER_26_227 ();
 sg13g2_fill_1 FILLER_26_241 ();
 sg13g2_fill_1 FILLER_26_267 ();
 sg13g2_fill_2 FILLER_26_291 ();
 sg13g2_fill_2 FILLER_26_311 ();
 sg13g2_fill_1 FILLER_26_319 ();
 sg13g2_decap_8 FILLER_26_356 ();
 sg13g2_fill_2 FILLER_26_363 ();
 sg13g2_decap_8 FILLER_26_370 ();
 sg13g2_decap_8 FILLER_26_377 ();
 sg13g2_decap_4 FILLER_26_384 ();
 sg13g2_fill_2 FILLER_26_388 ();
 sg13g2_fill_1 FILLER_26_408 ();
 sg13g2_fill_2 FILLER_27_0 ();
 sg13g2_fill_1 FILLER_27_2 ();
 sg13g2_fill_1 FILLER_27_88 ();
 sg13g2_fill_2 FILLER_27_108 ();
 sg13g2_fill_2 FILLER_27_136 ();
 sg13g2_fill_1 FILLER_27_138 ();
 sg13g2_fill_1 FILLER_27_147 ();
 sg13g2_fill_1 FILLER_27_161 ();
 sg13g2_decap_8 FILLER_27_191 ();
 sg13g2_decap_4 FILLER_27_206 ();
 sg13g2_fill_2 FILLER_27_210 ();
 sg13g2_fill_1 FILLER_27_271 ();
 sg13g2_decap_4 FILLER_27_289 ();
 sg13g2_fill_1 FILLER_27_334 ();
 sg13g2_decap_4 FILLER_27_348 ();
 sg13g2_decap_8 FILLER_27_356 ();
 sg13g2_fill_2 FILLER_27_367 ();
 sg13g2_fill_1 FILLER_27_376 ();
 sg13g2_fill_2 FILLER_27_381 ();
 sg13g2_fill_2 FILLER_28_40 ();
 sg13g2_fill_1 FILLER_28_42 ();
 sg13g2_fill_2 FILLER_28_54 ();
 sg13g2_fill_1 FILLER_28_56 ();
 sg13g2_fill_2 FILLER_28_92 ();
 sg13g2_fill_1 FILLER_28_94 ();
 sg13g2_fill_1 FILLER_28_131 ();
 sg13g2_fill_2 FILLER_28_147 ();
 sg13g2_fill_1 FILLER_28_149 ();
 sg13g2_fill_1 FILLER_28_163 ();
 sg13g2_decap_8 FILLER_28_177 ();
 sg13g2_decap_4 FILLER_28_184 ();
 sg13g2_decap_4 FILLER_28_214 ();
 sg13g2_fill_1 FILLER_28_222 ();
 sg13g2_decap_4 FILLER_28_232 ();
 sg13g2_fill_2 FILLER_28_236 ();
 sg13g2_decap_4 FILLER_28_248 ();
 sg13g2_fill_2 FILLER_28_265 ();
 sg13g2_fill_1 FILLER_28_267 ();
 sg13g2_fill_1 FILLER_28_281 ();
 sg13g2_decap_4 FILLER_28_337 ();
 sg13g2_fill_1 FILLER_28_341 ();
 sg13g2_fill_2 FILLER_28_347 ();
 sg13g2_fill_1 FILLER_28_349 ();
 sg13g2_fill_2 FILLER_28_358 ();
 sg13g2_fill_1 FILLER_28_360 ();
 sg13g2_decap_8 FILLER_28_385 ();
 sg13g2_fill_2 FILLER_28_392 ();
 sg13g2_fill_2 FILLER_28_407 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_fill_2 FILLER_29_33 ();
 sg13g2_fill_2 FILLER_29_65 ();
 sg13g2_fill_1 FILLER_29_67 ();
 sg13g2_decap_8 FILLER_29_76 ();
 sg13g2_fill_1 FILLER_29_83 ();
 sg13g2_fill_1 FILLER_29_105 ();
 sg13g2_fill_2 FILLER_29_135 ();
 sg13g2_decap_8 FILLER_29_141 ();
 sg13g2_fill_1 FILLER_29_152 ();
 sg13g2_fill_2 FILLER_29_160 ();
 sg13g2_decap_4 FILLER_29_170 ();
 sg13g2_decap_8 FILLER_29_178 ();
 sg13g2_decap_4 FILLER_29_185 ();
 sg13g2_decap_4 FILLER_29_215 ();
 sg13g2_fill_1 FILLER_29_219 ();
 sg13g2_decap_4 FILLER_29_233 ();
 sg13g2_fill_1 FILLER_29_237 ();
 sg13g2_fill_1 FILLER_29_256 ();
 sg13g2_decap_8 FILLER_29_291 ();
 sg13g2_decap_8 FILLER_29_298 ();
 sg13g2_fill_2 FILLER_29_305 ();
 sg13g2_fill_1 FILLER_29_307 ();
 sg13g2_decap_8 FILLER_29_324 ();
 sg13g2_decap_8 FILLER_29_331 ();
 sg13g2_fill_2 FILLER_29_351 ();
 sg13g2_fill_2 FILLER_29_361 ();
 sg13g2_fill_1 FILLER_29_363 ();
 sg13g2_decap_8 FILLER_29_398 ();
 sg13g2_decap_4 FILLER_29_405 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_4 FILLER_30_7 ();
 sg13g2_fill_2 FILLER_30_15 ();
 sg13g2_fill_1 FILLER_30_17 ();
 sg13g2_fill_2 FILLER_30_33 ();
 sg13g2_fill_1 FILLER_30_35 ();
 sg13g2_fill_2 FILLER_30_52 ();
 sg13g2_decap_8 FILLER_30_80 ();
 sg13g2_fill_1 FILLER_30_92 ();
 sg13g2_fill_2 FILLER_30_126 ();
 sg13g2_fill_2 FILLER_30_140 ();
 sg13g2_fill_2 FILLER_30_163 ();
 sg13g2_decap_8 FILLER_30_186 ();
 sg13g2_decap_4 FILLER_30_193 ();
 sg13g2_fill_2 FILLER_30_202 ();
 sg13g2_fill_2 FILLER_30_212 ();
 sg13g2_fill_2 FILLER_30_235 ();
 sg13g2_fill_1 FILLER_30_237 ();
 sg13g2_decap_8 FILLER_30_252 ();
 sg13g2_decap_8 FILLER_30_259 ();
 sg13g2_fill_2 FILLER_30_266 ();
 sg13g2_decap_4 FILLER_30_272 ();
 sg13g2_decap_8 FILLER_30_293 ();
 sg13g2_decap_8 FILLER_30_300 ();
 sg13g2_decap_8 FILLER_30_307 ();
 sg13g2_decap_8 FILLER_30_322 ();
 sg13g2_fill_2 FILLER_30_342 ();
 sg13g2_fill_2 FILLER_30_367 ();
 sg13g2_fill_1 FILLER_30_369 ();
 sg13g2_fill_2 FILLER_30_375 ();
 sg13g2_fill_1 FILLER_30_408 ();
 sg13g2_fill_2 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_15 ();
 sg13g2_decap_8 FILLER_31_22 ();
 sg13g2_decap_4 FILLER_31_98 ();
 sg13g2_fill_2 FILLER_31_102 ();
 sg13g2_fill_1 FILLER_31_169 ();
 sg13g2_fill_1 FILLER_31_183 ();
 sg13g2_decap_4 FILLER_31_192 ();
 sg13g2_fill_2 FILLER_31_196 ();
 sg13g2_decap_8 FILLER_31_202 ();
 sg13g2_fill_2 FILLER_31_209 ();
 sg13g2_fill_2 FILLER_31_214 ();
 sg13g2_fill_1 FILLER_31_216 ();
 sg13g2_fill_2 FILLER_31_265 ();
 sg13g2_fill_1 FILLER_31_267 ();
 sg13g2_decap_4 FILLER_31_351 ();
 sg13g2_fill_2 FILLER_31_355 ();
 sg13g2_fill_2 FILLER_31_362 ();
 sg13g2_decap_8 FILLER_31_372 ();
 sg13g2_decap_4 FILLER_31_379 ();
 sg13g2_fill_2 FILLER_31_383 ();
 sg13g2_fill_2 FILLER_31_406 ();
 sg13g2_fill_1 FILLER_31_408 ();
 sg13g2_decap_4 FILLER_32_83 ();
 sg13g2_decap_8 FILLER_32_103 ();
 sg13g2_decap_8 FILLER_32_110 ();
 sg13g2_decap_8 FILLER_32_117 ();
 sg13g2_fill_2 FILLER_32_124 ();
 sg13g2_fill_1 FILLER_32_126 ();
 sg13g2_fill_2 FILLER_32_177 ();
 sg13g2_fill_1 FILLER_32_226 ();
 sg13g2_fill_1 FILLER_32_237 ();
 sg13g2_decap_8 FILLER_32_322 ();
 sg13g2_decap_8 FILLER_32_329 ();
 sg13g2_decap_8 FILLER_32_336 ();
 sg13g2_fill_2 FILLER_32_343 ();
 sg13g2_fill_2 FILLER_32_349 ();
 sg13g2_fill_1 FILLER_32_351 ();
 sg13g2_fill_1 FILLER_32_362 ();
 sg13g2_decap_8 FILLER_32_381 ();
 sg13g2_decap_4 FILLER_32_388 ();
 sg13g2_fill_2 FILLER_32_392 ();
 sg13g2_fill_2 FILLER_33_0 ();
 sg13g2_fill_2 FILLER_33_42 ();
 sg13g2_fill_2 FILLER_33_70 ();
 sg13g2_fill_1 FILLER_33_72 ();
 sg13g2_decap_4 FILLER_33_107 ();
 sg13g2_fill_2 FILLER_33_111 ();
 sg13g2_fill_1 FILLER_33_117 ();
 sg13g2_decap_8 FILLER_33_123 ();
 sg13g2_decap_8 FILLER_33_130 ();
 sg13g2_decap_8 FILLER_33_137 ();
 sg13g2_decap_8 FILLER_33_144 ();
 sg13g2_decap_8 FILLER_33_151 ();
 sg13g2_decap_4 FILLER_33_158 ();
 sg13g2_decap_4 FILLER_33_167 ();
 sg13g2_fill_2 FILLER_33_171 ();
 sg13g2_fill_2 FILLER_33_194 ();
 sg13g2_fill_2 FILLER_33_271 ();
 sg13g2_decap_8 FILLER_33_277 ();
 sg13g2_fill_2 FILLER_33_297 ();
 sg13g2_decap_8 FILLER_33_325 ();
 sg13g2_fill_2 FILLER_33_360 ();
 sg13g2_fill_1 FILLER_33_362 ();
 sg13g2_fill_1 FILLER_33_388 ();
 sg13g2_decap_4 FILLER_33_403 ();
 sg13g2_fill_2 FILLER_33_407 ();
 sg13g2_fill_2 FILLER_34_26 ();
 sg13g2_fill_1 FILLER_34_41 ();
 sg13g2_fill_1 FILLER_34_106 ();
 sg13g2_decap_4 FILLER_34_132 ();
 sg13g2_fill_1 FILLER_34_136 ();
 sg13g2_decap_4 FILLER_34_146 ();
 sg13g2_decap_8 FILLER_34_155 ();
 sg13g2_fill_2 FILLER_34_162 ();
 sg13g2_fill_1 FILLER_34_172 ();
 sg13g2_fill_2 FILLER_34_185 ();
 sg13g2_decap_4 FILLER_34_217 ();
 sg13g2_fill_2 FILLER_34_229 ();
 sg13g2_decap_8 FILLER_34_247 ();
 sg13g2_fill_1 FILLER_34_254 ();
 sg13g2_decap_4 FILLER_34_285 ();
 sg13g2_fill_1 FILLER_34_289 ();
 sg13g2_decap_8 FILLER_34_316 ();
 sg13g2_fill_1 FILLER_34_323 ();
 sg13g2_fill_1 FILLER_34_408 ();
 sg13g2_fill_2 FILLER_35_23 ();
 sg13g2_fill_2 FILLER_35_34 ();
 sg13g2_fill_2 FILLER_35_44 ();
 sg13g2_fill_1 FILLER_35_99 ();
 sg13g2_fill_1 FILLER_35_132 ();
 sg13g2_fill_2 FILLER_35_138 ();
 sg13g2_fill_1 FILLER_35_140 ();
 sg13g2_decap_8 FILLER_35_239 ();
 sg13g2_decap_8 FILLER_35_246 ();
 sg13g2_decap_8 FILLER_35_253 ();
 sg13g2_decap_8 FILLER_35_260 ();
 sg13g2_fill_2 FILLER_35_267 ();
 sg13g2_fill_1 FILLER_35_269 ();
 sg13g2_decap_8 FILLER_35_274 ();
 sg13g2_decap_8 FILLER_35_281 ();
 sg13g2_decap_8 FILLER_35_288 ();
 sg13g2_decap_4 FILLER_35_295 ();
 sg13g2_fill_2 FILLER_35_299 ();
 sg13g2_decap_4 FILLER_35_305 ();
 sg13g2_fill_1 FILLER_35_309 ();
 sg13g2_decap_8 FILLER_35_314 ();
 sg13g2_fill_2 FILLER_35_346 ();
 sg13g2_fill_2 FILLER_35_353 ();
 sg13g2_fill_2 FILLER_35_373 ();
 sg13g2_fill_2 FILLER_35_383 ();
 sg13g2_fill_1 FILLER_35_385 ();
 sg13g2_fill_2 FILLER_35_394 ();
 sg13g2_fill_2 FILLER_36_14 ();
 sg13g2_fill_1 FILLER_36_26 ();
 sg13g2_fill_1 FILLER_36_42 ();
 sg13g2_fill_2 FILLER_36_51 ();
 sg13g2_fill_1 FILLER_36_121 ();
 sg13g2_fill_2 FILLER_36_144 ();
 sg13g2_fill_1 FILLER_36_162 ();
 sg13g2_fill_2 FILLER_36_168 ();
 sg13g2_fill_2 FILLER_36_227 ();
 sg13g2_fill_2 FILLER_36_285 ();
 sg13g2_fill_1 FILLER_36_287 ();
 sg13g2_decap_4 FILLER_36_293 ();
 sg13g2_decap_8 FILLER_36_301 ();
 sg13g2_decap_8 FILLER_36_321 ();
 sg13g2_decap_4 FILLER_36_328 ();
 sg13g2_fill_1 FILLER_36_332 ();
 sg13g2_decap_8 FILLER_36_341 ();
 sg13g2_decap_8 FILLER_36_348 ();
 sg13g2_decap_8 FILLER_36_355 ();
 sg13g2_decap_4 FILLER_36_362 ();
 sg13g2_decap_4 FILLER_36_370 ();
 sg13g2_fill_1 FILLER_36_374 ();
 sg13g2_fill_2 FILLER_36_382 ();
 sg13g2_fill_2 FILLER_36_406 ();
 sg13g2_fill_1 FILLER_36_408 ();
 sg13g2_fill_1 FILLER_37_0 ();
 sg13g2_fill_2 FILLER_37_49 ();
 sg13g2_decap_4 FILLER_37_86 ();
 sg13g2_fill_2 FILLER_37_102 ();
 sg13g2_fill_1 FILLER_37_104 ();
 sg13g2_decap_4 FILLER_37_110 ();
 sg13g2_fill_1 FILLER_37_122 ();
 sg13g2_fill_1 FILLER_37_135 ();
 sg13g2_fill_2 FILLER_37_174 ();
 sg13g2_fill_1 FILLER_37_200 ();
 sg13g2_fill_2 FILLER_37_244 ();
 sg13g2_fill_1 FILLER_37_251 ();
 sg13g2_fill_1 FILLER_37_256 ();
 sg13g2_fill_1 FILLER_37_297 ();
 sg13g2_decap_4 FILLER_37_324 ();
 sg13g2_fill_1 FILLER_37_328 ();
 sg13g2_fill_1 FILLER_37_342 ();
 sg13g2_fill_2 FILLER_37_372 ();
 sg13g2_decap_8 FILLER_37_401 ();
 sg13g2_fill_1 FILLER_37_408 ();
 sg13g2_fill_1 FILLER_38_42 ();
 sg13g2_fill_1 FILLER_38_49 ();
 sg13g2_fill_1 FILLER_38_76 ();
 sg13g2_fill_2 FILLER_38_106 ();
 sg13g2_fill_2 FILLER_38_139 ();
 sg13g2_decap_4 FILLER_38_156 ();
 sg13g2_fill_2 FILLER_38_218 ();
 sg13g2_fill_1 FILLER_38_224 ();
 sg13g2_fill_1 FILLER_38_257 ();
 sg13g2_fill_1 FILLER_38_265 ();
 sg13g2_decap_8 FILLER_38_338 ();
 sg13g2_fill_2 FILLER_38_345 ();
 sg13g2_fill_1 FILLER_38_347 ();
 sg13g2_fill_2 FILLER_38_356 ();
 sg13g2_fill_2 FILLER_38_395 ();
 sg13g2_fill_1 FILLER_38_397 ();
 sg13g2_fill_2 FILLER_38_406 ();
 sg13g2_fill_1 FILLER_38_408 ();
 sg13g2_fill_1 FILLER_39_30 ();
 sg13g2_fill_2 FILLER_39_51 ();
 sg13g2_fill_1 FILLER_39_53 ();
 sg13g2_fill_2 FILLER_39_64 ();
 sg13g2_fill_1 FILLER_39_66 ();
 sg13g2_fill_2 FILLER_39_95 ();
 sg13g2_fill_1 FILLER_39_97 ();
 sg13g2_fill_1 FILLER_39_120 ();
 sg13g2_fill_1 FILLER_39_146 ();
 sg13g2_decap_8 FILLER_39_165 ();
 sg13g2_decap_8 FILLER_39_172 ();
 sg13g2_decap_8 FILLER_39_179 ();
 sg13g2_fill_2 FILLER_39_186 ();
 sg13g2_decap_8 FILLER_39_192 ();
 sg13g2_decap_4 FILLER_39_199 ();
 sg13g2_fill_2 FILLER_39_206 ();
 sg13g2_fill_1 FILLER_39_208 ();
 sg13g2_fill_2 FILLER_39_244 ();
 sg13g2_fill_1 FILLER_39_246 ();
 sg13g2_fill_1 FILLER_39_270 ();
 sg13g2_fill_1 FILLER_39_327 ();
 sg13g2_fill_1 FILLER_39_333 ();
 sg13g2_decap_8 FILLER_39_342 ();
 sg13g2_fill_2 FILLER_39_349 ();
 sg13g2_decap_4 FILLER_39_356 ();
 sg13g2_fill_2 FILLER_39_375 ();
 sg13g2_fill_1 FILLER_39_377 ();
 sg13g2_fill_2 FILLER_39_385 ();
 sg13g2_fill_2 FILLER_39_407 ();
 sg13g2_decap_4 FILLER_40_0 ();
 sg13g2_fill_2 FILLER_40_4 ();
 sg13g2_fill_2 FILLER_40_46 ();
 sg13g2_fill_1 FILLER_40_48 ();
 sg13g2_fill_2 FILLER_40_67 ();
 sg13g2_fill_2 FILLER_40_78 ();
 sg13g2_fill_1 FILLER_40_80 ();
 sg13g2_fill_2 FILLER_40_96 ();
 sg13g2_fill_2 FILLER_40_113 ();
 sg13g2_decap_8 FILLER_40_136 ();
 sg13g2_decap_8 FILLER_40_143 ();
 sg13g2_decap_8 FILLER_40_150 ();
 sg13g2_decap_8 FILLER_40_157 ();
 sg13g2_decap_8 FILLER_40_164 ();
 sg13g2_fill_2 FILLER_40_171 ();
 sg13g2_fill_1 FILLER_40_173 ();
 sg13g2_decap_8 FILLER_40_212 ();
 sg13g2_decap_8 FILLER_40_219 ();
 sg13g2_fill_2 FILLER_40_226 ();
 sg13g2_fill_1 FILLER_40_228 ();
 sg13g2_decap_8 FILLER_40_233 ();
 sg13g2_fill_1 FILLER_40_240 ();
 sg13g2_fill_2 FILLER_40_317 ();
 sg13g2_fill_1 FILLER_40_334 ();
 sg13g2_decap_8 FILLER_40_363 ();
 sg13g2_fill_2 FILLER_40_370 ();
 sg13g2_fill_1 FILLER_40_372 ();
 sg13g2_fill_2 FILLER_40_382 ();
 sg13g2_decap_4 FILLER_41_0 ();
 sg13g2_fill_1 FILLER_41_23 ();
 sg13g2_decap_8 FILLER_41_89 ();
 sg13g2_decap_8 FILLER_41_96 ();
 sg13g2_decap_8 FILLER_41_103 ();
 sg13g2_decap_8 FILLER_41_110 ();
 sg13g2_fill_2 FILLER_41_117 ();
 sg13g2_decap_8 FILLER_41_145 ();
 sg13g2_decap_8 FILLER_41_152 ();
 sg13g2_decap_4 FILLER_41_159 ();
 sg13g2_fill_1 FILLER_41_163 ();
 sg13g2_fill_2 FILLER_41_190 ();
 sg13g2_fill_1 FILLER_41_218 ();
 sg13g2_decap_8 FILLER_41_231 ();
 sg13g2_decap_8 FILLER_41_238 ();
 sg13g2_decap_8 FILLER_41_245 ();
 sg13g2_fill_2 FILLER_41_252 ();
 sg13g2_fill_1 FILLER_41_254 ();
 sg13g2_fill_2 FILLER_41_264 ();
 sg13g2_fill_2 FILLER_41_274 ();
 sg13g2_fill_1 FILLER_41_311 ();
 sg13g2_fill_1 FILLER_41_323 ();
 sg13g2_fill_1 FILLER_41_348 ();
 sg13g2_fill_2 FILLER_41_406 ();
 sg13g2_fill_1 FILLER_41_408 ();
 sg13g2_decap_4 FILLER_42_64 ();
 sg13g2_decap_8 FILLER_42_94 ();
 sg13g2_decap_4 FILLER_42_101 ();
 sg13g2_decap_8 FILLER_42_109 ();
 sg13g2_decap_4 FILLER_42_116 ();
 sg13g2_fill_1 FILLER_42_120 ();
 sg13g2_fill_2 FILLER_42_147 ();
 sg13g2_decap_8 FILLER_42_188 ();
 sg13g2_decap_4 FILLER_42_195 ();
 sg13g2_fill_2 FILLER_42_307 ();
 sg13g2_fill_1 FILLER_42_323 ();
 sg13g2_fill_1 FILLER_42_345 ();
 sg13g2_fill_2 FILLER_42_357 ();
 sg13g2_fill_2 FILLER_42_373 ();
 sg13g2_fill_1 FILLER_42_375 ();
 sg13g2_fill_2 FILLER_42_389 ();
 sg13g2_fill_2 FILLER_42_395 ();
 sg13g2_fill_1 FILLER_42_397 ();
 sg13g2_fill_1 FILLER_42_408 ();
 sg13g2_fill_1 FILLER_43_26 ();
 sg13g2_fill_2 FILLER_43_51 ();
 sg13g2_fill_2 FILLER_43_64 ();
 sg13g2_fill_1 FILLER_43_66 ();
 sg13g2_fill_1 FILLER_43_179 ();
 sg13g2_decap_4 FILLER_43_206 ();
 sg13g2_fill_2 FILLER_43_210 ();
 sg13g2_fill_2 FILLER_43_289 ();
 sg13g2_fill_2 FILLER_43_313 ();
 sg13g2_fill_1 FILLER_43_342 ();
 sg13g2_fill_1 FILLER_43_351 ();
 sg13g2_decap_8 FILLER_43_369 ();
 sg13g2_decap_8 FILLER_43_376 ();
 sg13g2_decap_8 FILLER_43_383 ();
 sg13g2_fill_1 FILLER_43_390 ();
 sg13g2_fill_2 FILLER_43_406 ();
 sg13g2_fill_1 FILLER_43_408 ();
 sg13g2_decap_4 FILLER_44_0 ();
 sg13g2_fill_2 FILLER_44_24 ();
 sg13g2_fill_2 FILLER_44_43 ();
 sg13g2_fill_2 FILLER_44_94 ();
 sg13g2_fill_1 FILLER_44_96 ();
 sg13g2_fill_2 FILLER_44_123 ();
 sg13g2_fill_2 FILLER_44_140 ();
 sg13g2_fill_1 FILLER_44_142 ();
 sg13g2_decap_8 FILLER_44_204 ();
 sg13g2_decap_8 FILLER_44_211 ();
 sg13g2_fill_2 FILLER_44_218 ();
 sg13g2_fill_2 FILLER_44_280 ();
 sg13g2_fill_1 FILLER_44_282 ();
 sg13g2_fill_2 FILLER_44_315 ();
 sg13g2_fill_2 FILLER_44_329 ();
 sg13g2_fill_2 FILLER_44_348 ();
 sg13g2_fill_2 FILLER_44_361 ();
 sg13g2_fill_1 FILLER_44_363 ();
 sg13g2_fill_2 FILLER_44_372 ();
 sg13g2_fill_1 FILLER_44_374 ();
 sg13g2_fill_2 FILLER_44_387 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_fill_2 FILLER_45_71 ();
 sg13g2_decap_8 FILLER_45_112 ();
 sg13g2_decap_8 FILLER_45_119 ();
 sg13g2_fill_2 FILLER_45_126 ();
 sg13g2_decap_4 FILLER_45_132 ();
 sg13g2_decap_8 FILLER_45_144 ();
 sg13g2_decap_8 FILLER_45_155 ();
 sg13g2_decap_4 FILLER_45_162 ();
 sg13g2_fill_1 FILLER_45_166 ();
 sg13g2_fill_1 FILLER_45_171 ();
 sg13g2_fill_2 FILLER_45_185 ();
 sg13g2_fill_1 FILLER_45_187 ();
 sg13g2_fill_2 FILLER_45_214 ();
 sg13g2_fill_1 FILLER_45_216 ();
 sg13g2_decap_4 FILLER_45_222 ();
 sg13g2_decap_8 FILLER_45_239 ();
 sg13g2_fill_2 FILLER_45_246 ();
 sg13g2_fill_1 FILLER_45_248 ();
 sg13g2_fill_1 FILLER_45_262 ();
 sg13g2_fill_1 FILLER_45_286 ();
 sg13g2_fill_1 FILLER_45_296 ();
 sg13g2_fill_2 FILLER_45_303 ();
 sg13g2_fill_2 FILLER_45_320 ();
 sg13g2_fill_1 FILLER_45_322 ();
 sg13g2_fill_2 FILLER_45_358 ();
 sg13g2_fill_2 FILLER_45_370 ();
 sg13g2_fill_1 FILLER_45_372 ();
 sg13g2_fill_2 FILLER_45_386 ();
 sg13g2_fill_1 FILLER_45_388 ();
 sg13g2_fill_2 FILLER_45_406 ();
 sg13g2_fill_1 FILLER_45_408 ();
 sg13g2_fill_2 FILLER_46_0 ();
 sg13g2_fill_1 FILLER_46_2 ();
 sg13g2_fill_1 FILLER_46_53 ();
 sg13g2_decap_4 FILLER_46_97 ();
 sg13g2_fill_1 FILLER_46_113 ();
 sg13g2_fill_1 FILLER_46_124 ();
 sg13g2_fill_1 FILLER_46_135 ();
 sg13g2_fill_2 FILLER_46_146 ();
 sg13g2_fill_1 FILLER_46_158 ();
 sg13g2_fill_2 FILLER_46_164 ();
 sg13g2_fill_1 FILLER_46_166 ();
 sg13g2_fill_2 FILLER_46_184 ();
 sg13g2_fill_1 FILLER_46_186 ();
 sg13g2_fill_2 FILLER_46_204 ();
 sg13g2_decap_8 FILLER_46_246 ();
 sg13g2_decap_4 FILLER_46_253 ();
 sg13g2_fill_2 FILLER_46_261 ();
 sg13g2_fill_1 FILLER_46_303 ();
 sg13g2_fill_2 FILLER_46_317 ();
 sg13g2_fill_1 FILLER_46_319 ();
 sg13g2_fill_2 FILLER_46_328 ();
 sg13g2_fill_1 FILLER_46_330 ();
 sg13g2_decap_4 FILLER_46_347 ();
 sg13g2_fill_1 FILLER_46_375 ();
 sg13g2_fill_1 FILLER_46_408 ();
 sg13g2_fill_1 FILLER_47_34 ();
 sg13g2_fill_2 FILLER_47_98 ();
 sg13g2_fill_1 FILLER_47_100 ();
 sg13g2_fill_1 FILLER_47_127 ();
 sg13g2_fill_1 FILLER_47_164 ();
 sg13g2_fill_1 FILLER_47_176 ();
 sg13g2_fill_1 FILLER_47_206 ();
 sg13g2_fill_1 FILLER_47_273 ();
 sg13g2_fill_2 FILLER_47_286 ();
 sg13g2_fill_1 FILLER_47_302 ();
 sg13g2_fill_1 FILLER_47_307 ();
 sg13g2_fill_2 FILLER_47_363 ();
 sg13g2_fill_2 FILLER_48_0 ();
 sg13g2_fill_1 FILLER_48_38 ();
 sg13g2_fill_1 FILLER_48_127 ();
 sg13g2_fill_2 FILLER_48_136 ();
 sg13g2_fill_1 FILLER_48_138 ();
 sg13g2_fill_1 FILLER_48_147 ();
 sg13g2_fill_2 FILLER_48_156 ();
 sg13g2_fill_1 FILLER_48_158 ();
 sg13g2_fill_2 FILLER_48_167 ();
 sg13g2_fill_1 FILLER_48_200 ();
 sg13g2_fill_1 FILLER_48_251 ();
 sg13g2_fill_1 FILLER_48_267 ();
 sg13g2_decap_8 FILLER_48_289 ();
 sg13g2_fill_2 FILLER_48_296 ();
 sg13g2_fill_2 FILLER_48_307 ();
 sg13g2_fill_2 FILLER_48_314 ();
 sg13g2_fill_2 FILLER_48_328 ();
 sg13g2_fill_1 FILLER_48_330 ();
 sg13g2_decap_8 FILLER_48_336 ();
 sg13g2_decap_4 FILLER_48_343 ();
 sg13g2_fill_2 FILLER_48_347 ();
 sg13g2_decap_8 FILLER_48_353 ();
 sg13g2_fill_2 FILLER_48_360 ();
 sg13g2_fill_2 FILLER_48_365 ();
 sg13g2_fill_2 FILLER_48_371 ();
 sg13g2_fill_2 FILLER_48_380 ();
 sg13g2_fill_1 FILLER_48_382 ();
 sg13g2_fill_2 FILLER_48_406 ();
 sg13g2_fill_1 FILLER_48_408 ();
 sg13g2_fill_1 FILLER_49_99 ();
 sg13g2_fill_1 FILLER_49_131 ();
 sg13g2_fill_2 FILLER_49_153 ();
 sg13g2_fill_1 FILLER_49_155 ();
 sg13g2_fill_1 FILLER_49_178 ();
 sg13g2_decap_4 FILLER_49_204 ();
 sg13g2_fill_1 FILLER_49_222 ();
 sg13g2_fill_2 FILLER_49_228 ();
 sg13g2_fill_2 FILLER_49_243 ();
 sg13g2_fill_1 FILLER_49_280 ();
 sg13g2_fill_2 FILLER_49_305 ();
 sg13g2_decap_8 FILLER_49_334 ();
 sg13g2_decap_8 FILLER_49_341 ();
 sg13g2_decap_8 FILLER_49_348 ();
 sg13g2_fill_2 FILLER_49_360 ();
 sg13g2_fill_1 FILLER_49_367 ();
 sg13g2_fill_2 FILLER_49_373 ();
 sg13g2_fill_1 FILLER_49_375 ();
 sg13g2_fill_2 FILLER_49_385 ();
 sg13g2_decap_4 FILLER_49_392 ();
 sg13g2_fill_1 FILLER_49_396 ();
 sg13g2_fill_2 FILLER_49_406 ();
 sg13g2_fill_1 FILLER_49_408 ();
 sg13g2_fill_2 FILLER_50_0 ();
 sg13g2_fill_2 FILLER_50_67 ();
 sg13g2_fill_1 FILLER_50_69 ();
 sg13g2_fill_2 FILLER_50_88 ();
 sg13g2_fill_1 FILLER_50_98 ();
 sg13g2_fill_2 FILLER_50_121 ();
 sg13g2_fill_2 FILLER_50_143 ();
 sg13g2_fill_1 FILLER_50_145 ();
 sg13g2_fill_2 FILLER_50_163 ();
 sg13g2_fill_1 FILLER_50_165 ();
 sg13g2_fill_2 FILLER_50_170 ();
 sg13g2_decap_4 FILLER_50_197 ();
 sg13g2_decap_8 FILLER_50_205 ();
 sg13g2_decap_4 FILLER_50_212 ();
 sg13g2_fill_2 FILLER_50_216 ();
 sg13g2_fill_1 FILLER_50_226 ();
 sg13g2_decap_8 FILLER_50_239 ();
 sg13g2_fill_2 FILLER_50_246 ();
 sg13g2_fill_2 FILLER_50_305 ();
 sg13g2_fill_2 FILLER_50_315 ();
 sg13g2_decap_4 FILLER_50_343 ();
 sg13g2_fill_1 FILLER_50_347 ();
 sg13g2_fill_1 FILLER_50_359 ();
 sg13g2_fill_2 FILLER_50_406 ();
 sg13g2_fill_1 FILLER_50_408 ();
 sg13g2_fill_2 FILLER_51_0 ();
 sg13g2_fill_1 FILLER_51_2 ();
 sg13g2_fill_2 FILLER_51_40 ();
 sg13g2_fill_1 FILLER_51_42 ();
 sg13g2_fill_2 FILLER_51_78 ();
 sg13g2_fill_1 FILLER_51_110 ();
 sg13g2_fill_1 FILLER_51_132 ();
 sg13g2_decap_8 FILLER_51_162 ();
 sg13g2_decap_4 FILLER_51_169 ();
 sg13g2_fill_1 FILLER_51_173 ();
 sg13g2_fill_1 FILLER_51_195 ();
 sg13g2_fill_1 FILLER_51_206 ();
 sg13g2_fill_1 FILLER_51_220 ();
 sg13g2_fill_2 FILLER_51_224 ();
 sg13g2_fill_1 FILLER_51_226 ();
 sg13g2_decap_8 FILLER_51_232 ();
 sg13g2_decap_4 FILLER_51_239 ();
 sg13g2_fill_2 FILLER_51_243 ();
 sg13g2_fill_1 FILLER_51_265 ();
 sg13g2_fill_1 FILLER_51_280 ();
 sg13g2_fill_1 FILLER_51_327 ();
 sg13g2_fill_1 FILLER_51_344 ();
 sg13g2_fill_2 FILLER_51_349 ();
 sg13g2_fill_1 FILLER_51_351 ();
 sg13g2_fill_1 FILLER_51_377 ();
 sg13g2_fill_2 FILLER_51_388 ();
 sg13g2_fill_2 FILLER_51_406 ();
 sg13g2_fill_1 FILLER_51_408 ();
 sg13g2_fill_2 FILLER_52_71 ();
 sg13g2_fill_1 FILLER_52_73 ();
 sg13g2_fill_2 FILLER_52_109 ();
 sg13g2_fill_1 FILLER_52_111 ();
 sg13g2_fill_2 FILLER_52_128 ();
 sg13g2_fill_1 FILLER_52_130 ();
 sg13g2_decap_8 FILLER_52_135 ();
 sg13g2_fill_1 FILLER_52_142 ();
 sg13g2_decap_8 FILLER_52_160 ();
 sg13g2_fill_2 FILLER_52_182 ();
 sg13g2_fill_1 FILLER_52_199 ();
 sg13g2_fill_2 FILLER_52_248 ();
 sg13g2_fill_1 FILLER_52_250 ();
 sg13g2_fill_2 FILLER_52_290 ();
 sg13g2_fill_1 FILLER_52_323 ();
 sg13g2_fill_1 FILLER_52_408 ();
 sg13g2_fill_1 FILLER_53_100 ();
 sg13g2_decap_8 FILLER_53_135 ();
 sg13g2_decap_8 FILLER_53_142 ();
 sg13g2_fill_2 FILLER_53_183 ();
 sg13g2_fill_2 FILLER_53_193 ();
 sg13g2_fill_1 FILLER_53_215 ();
 sg13g2_decap_4 FILLER_53_237 ();
 sg13g2_fill_1 FILLER_53_262 ();
 sg13g2_fill_1 FILLER_53_289 ();
 sg13g2_fill_2 FILLER_53_304 ();
 sg13g2_fill_1 FILLER_53_306 ();
 sg13g2_decap_4 FILLER_53_327 ();
 sg13g2_decap_8 FILLER_53_347 ();
 sg13g2_fill_2 FILLER_53_354 ();
 sg13g2_fill_1 FILLER_53_356 ();
 sg13g2_fill_2 FILLER_53_406 ();
 sg13g2_fill_1 FILLER_53_408 ();
 sg13g2_fill_2 FILLER_54_40 ();
 sg13g2_fill_2 FILLER_54_68 ();
 sg13g2_fill_2 FILLER_54_91 ();
 sg13g2_fill_2 FILLER_54_164 ();
 sg13g2_fill_1 FILLER_54_166 ();
 sg13g2_fill_2 FILLER_54_173 ();
 sg13g2_fill_1 FILLER_54_175 ();
 sg13g2_decap_4 FILLER_54_191 ();
 sg13g2_decap_8 FILLER_54_208 ();
 sg13g2_decap_4 FILLER_54_215 ();
 sg13g2_fill_2 FILLER_54_235 ();
 sg13g2_fill_1 FILLER_54_237 ();
 sg13g2_fill_2 FILLER_54_345 ();
 sg13g2_fill_2 FILLER_54_353 ();
 sg13g2_fill_1 FILLER_54_355 ();
 sg13g2_fill_2 FILLER_54_359 ();
 sg13g2_fill_1 FILLER_54_361 ();
 sg13g2_fill_1 FILLER_54_373 ();
 sg13g2_decap_4 FILLER_54_404 ();
 sg13g2_fill_1 FILLER_54_408 ();
 sg13g2_fill_2 FILLER_55_38 ();
 sg13g2_fill_1 FILLER_55_50 ();
 sg13g2_fill_1 FILLER_55_61 ();
 sg13g2_fill_2 FILLER_55_93 ();
 sg13g2_fill_1 FILLER_55_95 ();
 sg13g2_fill_1 FILLER_55_114 ();
 sg13g2_fill_2 FILLER_55_148 ();
 sg13g2_fill_1 FILLER_55_155 ();
 sg13g2_fill_2 FILLER_55_168 ();
 sg13g2_fill_1 FILLER_55_170 ();
 sg13g2_decap_8 FILLER_55_179 ();
 sg13g2_fill_2 FILLER_55_186 ();
 sg13g2_fill_2 FILLER_55_193 ();
 sg13g2_fill_2 FILLER_55_199 ();
 sg13g2_fill_1 FILLER_55_201 ();
 sg13g2_fill_1 FILLER_55_221 ();
 sg13g2_fill_1 FILLER_55_243 ();
 sg13g2_fill_1 FILLER_55_313 ();
 sg13g2_fill_1 FILLER_55_322 ();
 sg13g2_decap_4 FILLER_55_342 ();
 sg13g2_fill_1 FILLER_55_346 ();
 sg13g2_fill_2 FILLER_55_358 ();
 sg13g2_decap_8 FILLER_55_370 ();
 sg13g2_decap_4 FILLER_55_377 ();
 sg13g2_fill_1 FILLER_55_381 ();
 sg13g2_decap_4 FILLER_55_387 ();
 sg13g2_decap_4 FILLER_55_405 ();
 sg13g2_fill_1 FILLER_56_0 ();
 sg13g2_fill_2 FILLER_56_45 ();
 sg13g2_fill_2 FILLER_56_51 ();
 sg13g2_fill_1 FILLER_56_122 ();
 sg13g2_fill_2 FILLER_56_161 ();
 sg13g2_decap_4 FILLER_56_168 ();
 sg13g2_fill_1 FILLER_56_172 ();
 sg13g2_fill_2 FILLER_56_188 ();
 sg13g2_fill_1 FILLER_56_190 ();
 sg13g2_fill_1 FILLER_56_262 ();
 sg13g2_fill_2 FILLER_56_272 ();
 sg13g2_fill_1 FILLER_56_274 ();
 sg13g2_fill_2 FILLER_56_284 ();
 sg13g2_fill_1 FILLER_56_286 ();
 sg13g2_decap_4 FILLER_56_332 ();
 sg13g2_fill_2 FILLER_56_336 ();
 sg13g2_decap_8 FILLER_56_365 ();
 sg13g2_fill_2 FILLER_56_393 ();
 sg13g2_fill_1 FILLER_56_395 ();
 sg13g2_fill_2 FILLER_57_26 ();
 sg13g2_fill_1 FILLER_57_57 ();
 sg13g2_fill_1 FILLER_57_62 ();
 sg13g2_fill_2 FILLER_57_88 ();
 sg13g2_fill_1 FILLER_57_137 ();
 sg13g2_decap_8 FILLER_57_156 ();
 sg13g2_fill_1 FILLER_57_163 ();
 sg13g2_fill_2 FILLER_57_168 ();
 sg13g2_fill_1 FILLER_57_170 ();
 sg13g2_fill_2 FILLER_57_181 ();
 sg13g2_fill_2 FILLER_57_188 ();
 sg13g2_fill_2 FILLER_57_195 ();
 sg13g2_fill_1 FILLER_57_197 ();
 sg13g2_fill_1 FILLER_57_217 ();
 sg13g2_fill_2 FILLER_57_256 ();
 sg13g2_fill_1 FILLER_57_267 ();
 sg13g2_fill_1 FILLER_57_274 ();
 sg13g2_fill_1 FILLER_57_343 ();
 sg13g2_fill_2 FILLER_57_360 ();
 sg13g2_fill_1 FILLER_57_367 ();
 sg13g2_fill_1 FILLER_57_408 ();
 sg13g2_fill_2 FILLER_58_0 ();
 sg13g2_fill_1 FILLER_58_34 ();
 sg13g2_fill_1 FILLER_58_66 ();
 sg13g2_fill_2 FILLER_58_92 ();
 sg13g2_fill_1 FILLER_58_155 ();
 sg13g2_fill_2 FILLER_58_169 ();
 sg13g2_fill_2 FILLER_58_189 ();
 sg13g2_fill_2 FILLER_58_201 ();
 sg13g2_fill_2 FILLER_58_239 ();
 sg13g2_fill_1 FILLER_58_241 ();
 sg13g2_fill_2 FILLER_58_260 ();
 sg13g2_fill_1 FILLER_58_277 ();
 sg13g2_fill_1 FILLER_58_304 ();
 sg13g2_fill_2 FILLER_58_315 ();
 sg13g2_fill_1 FILLER_58_317 ();
 sg13g2_fill_1 FILLER_58_324 ();
 sg13g2_fill_1 FILLER_58_336 ();
 sg13g2_fill_1 FILLER_58_342 ();
 sg13g2_fill_1 FILLER_58_408 ();
 sg13g2_fill_2 FILLER_59_85 ();
 sg13g2_fill_1 FILLER_59_144 ();
 sg13g2_fill_1 FILLER_59_171 ();
 sg13g2_fill_2 FILLER_59_180 ();
 sg13g2_fill_1 FILLER_59_182 ();
 sg13g2_fill_2 FILLER_59_197 ();
 sg13g2_fill_2 FILLER_59_248 ();
 sg13g2_fill_2 FILLER_59_261 ();
 sg13g2_fill_1 FILLER_59_263 ();
 sg13g2_fill_2 FILLER_59_368 ();
 sg13g2_fill_1 FILLER_59_387 ();
 sg13g2_fill_1 FILLER_60_43 ();
 sg13g2_fill_2 FILLER_60_49 ();
 sg13g2_fill_2 FILLER_60_74 ();
 sg13g2_fill_2 FILLER_60_113 ();
 sg13g2_fill_2 FILLER_60_165 ();
 sg13g2_fill_1 FILLER_60_167 ();
 sg13g2_fill_2 FILLER_60_223 ();
 sg13g2_fill_1 FILLER_60_250 ();
 sg13g2_fill_2 FILLER_60_261 ();
 sg13g2_fill_1 FILLER_60_283 ();
 sg13g2_fill_2 FILLER_60_293 ();
 sg13g2_fill_1 FILLER_60_295 ();
 sg13g2_fill_2 FILLER_60_325 ();
 sg13g2_fill_2 FILLER_60_342 ();
 sg13g2_fill_2 FILLER_60_357 ();
 sg13g2_fill_1 FILLER_60_391 ();
 sg13g2_decap_8 FILLER_60_400 ();
 sg13g2_fill_2 FILLER_60_407 ();
 sg13g2_fill_1 FILLER_61_44 ();
 sg13g2_fill_2 FILLER_61_221 ();
 sg13g2_fill_2 FILLER_61_249 ();
 sg13g2_fill_2 FILLER_61_307 ();
 sg13g2_fill_2 FILLER_61_318 ();
 sg13g2_fill_1 FILLER_61_320 ();
 sg13g2_fill_2 FILLER_61_327 ();
 sg13g2_fill_1 FILLER_61_341 ();
 sg13g2_fill_2 FILLER_61_357 ();
 sg13g2_fill_1 FILLER_61_359 ();
 sg13g2_fill_2 FILLER_61_387 ();
 sg13g2_decap_4 FILLER_61_393 ();
 sg13g2_fill_1 FILLER_61_397 ();
 sg13g2_decap_8 FILLER_61_402 ();
 sg13g2_fill_1 FILLER_62_32 ();
 sg13g2_fill_2 FILLER_62_62 ();
 sg13g2_fill_1 FILLER_62_86 ();
 sg13g2_fill_2 FILLER_62_145 ();
 sg13g2_decap_4 FILLER_62_182 ();
 sg13g2_fill_2 FILLER_62_212 ();
 sg13g2_fill_1 FILLER_62_214 ();
 sg13g2_fill_1 FILLER_62_233 ();
 sg13g2_fill_2 FILLER_62_260 ();
 sg13g2_fill_2 FILLER_62_335 ();
 sg13g2_fill_1 FILLER_62_337 ();
 sg13g2_fill_2 FILLER_62_350 ();
 sg13g2_decap_8 FILLER_62_371 ();
 sg13g2_decap_4 FILLER_62_378 ();
 sg13g2_fill_1 FILLER_62_382 ();
 sg13g2_fill_1 FILLER_62_408 ();
 sg13g2_fill_1 FILLER_63_107 ();
 sg13g2_fill_1 FILLER_63_138 ();
 sg13g2_fill_2 FILLER_63_152 ();
 sg13g2_fill_2 FILLER_63_193 ();
 sg13g2_fill_2 FILLER_63_203 ();
 sg13g2_fill_1 FILLER_63_205 ();
 sg13g2_decap_8 FILLER_63_210 ();
 sg13g2_decap_4 FILLER_63_217 ();
 sg13g2_fill_2 FILLER_63_221 ();
 sg13g2_fill_1 FILLER_63_258 ();
 sg13g2_fill_2 FILLER_63_290 ();
 sg13g2_fill_2 FILLER_63_322 ();
 sg13g2_fill_1 FILLER_63_324 ();
 sg13g2_fill_1 FILLER_63_341 ();
 sg13g2_fill_1 FILLER_63_355 ();
 sg13g2_decap_4 FILLER_63_368 ();
 sg13g2_fill_1 FILLER_63_372 ();
 sg13g2_fill_1 FILLER_64_0 ();
 sg13g2_fill_2 FILLER_64_25 ();
 sg13g2_fill_1 FILLER_64_32 ();
 sg13g2_fill_1 FILLER_64_175 ();
 sg13g2_fill_1 FILLER_64_193 ();
 sg13g2_fill_2 FILLER_64_263 ();
 sg13g2_decap_8 FILLER_64_363 ();
 sg13g2_fill_2 FILLER_64_370 ();
 sg13g2_fill_1 FILLER_64_372 ();
 sg13g2_fill_2 FILLER_64_383 ();
 sg13g2_fill_2 FILLER_64_406 ();
 sg13g2_fill_1 FILLER_64_408 ();
 sg13g2_fill_1 FILLER_65_54 ();
 sg13g2_fill_2 FILLER_65_138 ();
 sg13g2_fill_1 FILLER_65_140 ();
 sg13g2_fill_1 FILLER_65_188 ();
 sg13g2_fill_2 FILLER_65_197 ();
 sg13g2_fill_2 FILLER_65_280 ();
 sg13g2_fill_1 FILLER_65_305 ();
 sg13g2_decap_4 FILLER_65_352 ();
 sg13g2_fill_1 FILLER_65_380 ();
 sg13g2_decap_8 FILLER_65_401 ();
 sg13g2_fill_1 FILLER_65_408 ();
 sg13g2_fill_1 FILLER_66_46 ();
 sg13g2_fill_2 FILLER_66_56 ();
 sg13g2_fill_1 FILLER_66_84 ();
 sg13g2_fill_2 FILLER_66_139 ();
 sg13g2_fill_1 FILLER_66_161 ();
 sg13g2_fill_1 FILLER_66_186 ();
 sg13g2_fill_1 FILLER_66_208 ();
 sg13g2_fill_2 FILLER_66_213 ();
 sg13g2_fill_1 FILLER_66_215 ();
 sg13g2_fill_1 FILLER_66_223 ();
 sg13g2_fill_1 FILLER_66_249 ();
 sg13g2_fill_1 FILLER_66_278 ();
 sg13g2_fill_2 FILLER_66_335 ();
 sg13g2_fill_1 FILLER_66_337 ();
 sg13g2_decap_4 FILLER_66_353 ();
 sg13g2_fill_2 FILLER_66_377 ();
 sg13g2_fill_2 FILLER_66_388 ();
 sg13g2_fill_2 FILLER_66_406 ();
 sg13g2_fill_1 FILLER_66_408 ();
 sg13g2_fill_2 FILLER_67_0 ();
 sg13g2_fill_1 FILLER_67_2 ();
 sg13g2_fill_2 FILLER_67_57 ();
 sg13g2_fill_1 FILLER_67_142 ();
 sg13g2_decap_8 FILLER_67_178 ();
 sg13g2_decap_4 FILLER_67_185 ();
 sg13g2_fill_2 FILLER_67_189 ();
 sg13g2_fill_1 FILLER_67_250 ();
 sg13g2_fill_1 FILLER_67_260 ();
 sg13g2_fill_1 FILLER_67_300 ();
 sg13g2_fill_2 FILLER_67_379 ();
 sg13g2_fill_2 FILLER_67_386 ();
 sg13g2_fill_2 FILLER_68_58 ();
 sg13g2_fill_1 FILLER_68_60 ();
 sg13g2_fill_2 FILLER_68_160 ();
 sg13g2_fill_1 FILLER_68_162 ();
 sg13g2_decap_4 FILLER_68_168 ();
 sg13g2_fill_1 FILLER_68_172 ();
 sg13g2_decap_4 FILLER_68_176 ();
 sg13g2_fill_1 FILLER_68_180 ();
 sg13g2_fill_2 FILLER_68_202 ();
 sg13g2_fill_1 FILLER_68_204 ();
 sg13g2_fill_2 FILLER_68_238 ();
 sg13g2_fill_1 FILLER_68_254 ();
 sg13g2_fill_1 FILLER_68_330 ();
 sg13g2_fill_1 FILLER_68_338 ();
 sg13g2_fill_1 FILLER_68_342 ();
 sg13g2_fill_2 FILLER_68_364 ();
 sg13g2_fill_1 FILLER_68_366 ();
 sg13g2_fill_1 FILLER_69_0 ();
 sg13g2_fill_2 FILLER_69_107 ();
 sg13g2_fill_1 FILLER_69_128 ();
 sg13g2_fill_2 FILLER_69_134 ();
 sg13g2_decap_8 FILLER_69_156 ();
 sg13g2_fill_2 FILLER_69_163 ();
 sg13g2_fill_1 FILLER_69_165 ();
 sg13g2_fill_2 FILLER_69_180 ();
 sg13g2_fill_2 FILLER_69_187 ();
 sg13g2_fill_1 FILLER_69_225 ();
 sg13g2_fill_1 FILLER_69_235 ();
 sg13g2_decap_8 FILLER_69_329 ();
 sg13g2_decap_8 FILLER_69_336 ();
 sg13g2_decap_4 FILLER_69_343 ();
 sg13g2_fill_1 FILLER_69_347 ();
 sg13g2_fill_1 FILLER_69_353 ();
 sg13g2_fill_2 FILLER_69_368 ();
 sg13g2_fill_1 FILLER_69_370 ();
 sg13g2_fill_1 FILLER_69_388 ();
 sg13g2_fill_2 FILLER_70_0 ();
 sg13g2_fill_2 FILLER_70_28 ();
 sg13g2_fill_2 FILLER_70_56 ();
 sg13g2_fill_2 FILLER_70_84 ();
 sg13g2_fill_1 FILLER_70_96 ();
 sg13g2_fill_1 FILLER_70_158 ();
 sg13g2_fill_2 FILLER_70_209 ();
 sg13g2_fill_1 FILLER_70_211 ();
 sg13g2_fill_1 FILLER_70_249 ();
 sg13g2_fill_1 FILLER_70_268 ();
 sg13g2_decap_8 FILLER_70_340 ();
 sg13g2_decap_4 FILLER_70_347 ();
 sg13g2_fill_1 FILLER_70_351 ();
 sg13g2_fill_1 FILLER_70_365 ();
 sg13g2_fill_2 FILLER_70_388 ();
 sg13g2_fill_1 FILLER_70_395 ();
 sg13g2_fill_2 FILLER_71_0 ();
 sg13g2_fill_1 FILLER_71_2 ();
 sg13g2_fill_2 FILLER_71_187 ();
 sg13g2_fill_2 FILLER_71_223 ();
 sg13g2_fill_2 FILLER_71_264 ();
 sg13g2_fill_1 FILLER_71_275 ();
 sg13g2_decap_4 FILLER_71_349 ();
 sg13g2_fill_1 FILLER_71_353 ();
 sg13g2_fill_2 FILLER_71_385 ();
 sg13g2_fill_1 FILLER_72_0 ();
 sg13g2_fill_2 FILLER_72_13 ();
 sg13g2_fill_1 FILLER_72_34 ();
 sg13g2_fill_2 FILLER_72_56 ();
 sg13g2_fill_1 FILLER_72_159 ();
 sg13g2_fill_2 FILLER_72_189 ();
 sg13g2_fill_1 FILLER_72_191 ();
 sg13g2_fill_1 FILLER_72_218 ();
 sg13g2_fill_2 FILLER_72_275 ();
 sg13g2_fill_1 FILLER_72_318 ();
 sg13g2_decap_4 FILLER_72_358 ();
 sg13g2_fill_2 FILLER_72_362 ();
 sg13g2_fill_1 FILLER_72_376 ();
 sg13g2_fill_1 FILLER_72_408 ();
 sg13g2_fill_2 FILLER_73_66 ();
 sg13g2_fill_1 FILLER_73_68 ();
 sg13g2_fill_1 FILLER_73_83 ();
 sg13g2_fill_1 FILLER_73_93 ();
 sg13g2_fill_2 FILLER_73_141 ();
 sg13g2_fill_1 FILLER_73_143 ();
 sg13g2_fill_2 FILLER_73_152 ();
 sg13g2_fill_1 FILLER_73_154 ();
 sg13g2_fill_2 FILLER_73_173 ();
 sg13g2_fill_1 FILLER_73_181 ();
 sg13g2_decap_4 FILLER_73_197 ();
 sg13g2_fill_1 FILLER_73_201 ();
 sg13g2_fill_1 FILLER_73_229 ();
 sg13g2_fill_1 FILLER_73_240 ();
 sg13g2_fill_1 FILLER_73_305 ();
 sg13g2_fill_2 FILLER_73_337 ();
 sg13g2_fill_1 FILLER_73_339 ();
 sg13g2_fill_1 FILLER_73_365 ();
 sg13g2_fill_1 FILLER_73_384 ();
 sg13g2_fill_1 FILLER_73_392 ();
 sg13g2_fill_1 FILLER_73_408 ();
 sg13g2_fill_1 FILLER_74_0 ();
 sg13g2_fill_1 FILLER_74_70 ();
 sg13g2_fill_2 FILLER_74_88 ();
 sg13g2_fill_2 FILLER_74_110 ();
 sg13g2_fill_1 FILLER_74_112 ();
 sg13g2_fill_1 FILLER_74_136 ();
 sg13g2_fill_1 FILLER_74_167 ();
 sg13g2_decap_4 FILLER_74_205 ();
 sg13g2_fill_1 FILLER_74_209 ();
 sg13g2_fill_2 FILLER_74_261 ();
 sg13g2_fill_1 FILLER_74_301 ();
 sg13g2_fill_1 FILLER_74_317 ();
 sg13g2_decap_8 FILLER_74_323 ();
 sg13g2_fill_2 FILLER_74_330 ();
 sg13g2_fill_1 FILLER_74_332 ();
 sg13g2_fill_2 FILLER_74_338 ();
 sg13g2_fill_1 FILLER_74_340 ();
 sg13g2_decap_8 FILLER_74_363 ();
 sg13g2_decap_8 FILLER_74_379 ();
 sg13g2_fill_1 FILLER_74_386 ();
 sg13g2_decap_4 FILLER_74_404 ();
 sg13g2_fill_1 FILLER_74_408 ();
 sg13g2_fill_1 FILLER_75_48 ();
 sg13g2_fill_1 FILLER_75_92 ();
 sg13g2_fill_2 FILLER_75_116 ();
 sg13g2_fill_2 FILLER_75_178 ();
 sg13g2_fill_2 FILLER_75_194 ();
 sg13g2_fill_2 FILLER_75_248 ();
 sg13g2_fill_2 FILLER_75_297 ();
 sg13g2_fill_1 FILLER_75_307 ();
 sg13g2_decap_8 FILLER_75_326 ();
 sg13g2_decap_4 FILLER_75_333 ();
 sg13g2_fill_1 FILLER_75_346 ();
 sg13g2_decap_8 FILLER_75_360 ();
 sg13g2_decap_8 FILLER_75_367 ();
 sg13g2_decap_8 FILLER_75_374 ();
 sg13g2_fill_2 FILLER_75_381 ();
 sg13g2_fill_2 FILLER_76_0 ();
 sg13g2_fill_1 FILLER_76_2 ();
 sg13g2_fill_1 FILLER_76_7 ();
 sg13g2_fill_1 FILLER_76_29 ();
 sg13g2_fill_1 FILLER_76_112 ();
 sg13g2_fill_1 FILLER_76_118 ();
 sg13g2_fill_1 FILLER_76_131 ();
 sg13g2_fill_2 FILLER_76_204 ();
 sg13g2_fill_1 FILLER_76_221 ();
 sg13g2_fill_1 FILLER_76_236 ();
 sg13g2_fill_1 FILLER_76_254 ();
 sg13g2_fill_2 FILLER_76_290 ();
 sg13g2_fill_1 FILLER_76_326 ();
 sg13g2_fill_1 FILLER_76_333 ();
 sg13g2_fill_2 FILLER_76_360 ();
 sg13g2_decap_4 FILLER_76_388 ();
 sg13g2_fill_2 FILLER_76_392 ();
 sg13g2_decap_8 FILLER_76_398 ();
 sg13g2_decap_4 FILLER_76_405 ();
 sg13g2_fill_2 FILLER_77_70 ();
 sg13g2_fill_1 FILLER_77_91 ();
 sg13g2_fill_2 FILLER_77_143 ();
 sg13g2_fill_1 FILLER_77_169 ();
 sg13g2_fill_2 FILLER_77_226 ();
 sg13g2_fill_1 FILLER_77_228 ();
 sg13g2_decap_8 FILLER_77_281 ();
 sg13g2_fill_1 FILLER_77_288 ();
 sg13g2_decap_8 FILLER_77_293 ();
 sg13g2_fill_1 FILLER_77_300 ();
 sg13g2_fill_1 FILLER_77_338 ();
 sg13g2_decap_4 FILLER_77_403 ();
 sg13g2_fill_2 FILLER_77_407 ();
 sg13g2_fill_2 FILLER_78_119 ();
 sg13g2_fill_1 FILLER_78_174 ();
 sg13g2_fill_2 FILLER_78_189 ();
 sg13g2_fill_1 FILLER_78_191 ();
 sg13g2_fill_1 FILLER_78_270 ();
 sg13g2_fill_2 FILLER_78_276 ();
 sg13g2_fill_2 FILLER_78_320 ();
 sg13g2_fill_1 FILLER_78_322 ();
 sg13g2_fill_2 FILLER_78_381 ();
 sg13g2_fill_2 FILLER_79_0 ();
 sg13g2_fill_2 FILLER_79_28 ();
 sg13g2_fill_1 FILLER_79_34 ();
 sg13g2_fill_1 FILLER_79_44 ();
 sg13g2_fill_2 FILLER_79_136 ();
 sg13g2_fill_1 FILLER_79_138 ();
 sg13g2_fill_1 FILLER_79_182 ();
 sg13g2_fill_2 FILLER_79_209 ();
 sg13g2_fill_1 FILLER_79_211 ();
 sg13g2_fill_2 FILLER_79_242 ();
 sg13g2_fill_1 FILLER_79_244 ();
 sg13g2_fill_2 FILLER_79_271 ();
 sg13g2_fill_2 FILLER_79_307 ();
 sg13g2_fill_2 FILLER_79_317 ();
 sg13g2_fill_1 FILLER_79_339 ();
 sg13g2_fill_1 FILLER_79_363 ();
 sg13g2_fill_2 FILLER_79_406 ();
 sg13g2_fill_1 FILLER_79_408 ();
 sg13g2_fill_1 FILLER_80_0 ();
 sg13g2_fill_1 FILLER_80_79 ();
 sg13g2_fill_2 FILLER_80_94 ();
 sg13g2_fill_1 FILLER_80_106 ();
 sg13g2_fill_1 FILLER_80_115 ();
 sg13g2_fill_2 FILLER_80_121 ();
 sg13g2_fill_1 FILLER_80_123 ();
 sg13g2_fill_2 FILLER_80_157 ();
 sg13g2_fill_1 FILLER_80_159 ();
 sg13g2_fill_2 FILLER_80_192 ();
 sg13g2_fill_1 FILLER_80_206 ();
 sg13g2_fill_2 FILLER_80_220 ();
 sg13g2_decap_8 FILLER_80_226 ();
 sg13g2_fill_2 FILLER_80_233 ();
 sg13g2_fill_1 FILLER_80_235 ();
 sg13g2_fill_2 FILLER_80_244 ();
 sg13g2_decap_8 FILLER_80_303 ();
 sg13g2_decap_8 FILLER_80_310 ();
 sg13g2_decap_4 FILLER_80_317 ();
 sg13g2_fill_2 FILLER_80_321 ();
 sg13g2_decap_8 FILLER_80_335 ();
 sg13g2_decap_8 FILLER_80_342 ();
 sg13g2_decap_8 FILLER_80_358 ();
 sg13g2_decap_8 FILLER_80_365 ();
 sg13g2_fill_1 FILLER_80_372 ();
 sg13g2_fill_2 FILLER_80_381 ();
 assign uio_oe[0] = net2;
 assign uio_oe[1] = net3;
 assign uio_oe[2] = net4;
 assign uio_oe[3] = net5;
 assign uio_oe[4] = net6;
 assign uio_oe[5] = net7;
 assign uio_oe[6] = net8;
 assign uio_oe[7] = net277;
 assign uio_out[0] = net9;
 assign uio_out[1] = net10;
 assign uio_out[2] = net11;
 assign uio_out[3] = net12;
 assign uio_out[4] = net13;
 assign uio_out[5] = net14;
 assign uio_out[6] = net15;
endmodule

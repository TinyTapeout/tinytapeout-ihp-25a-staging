module tt_um_patater_demokit (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire net29;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire clknet_0_clk;
 wire \frame[0] ;
 wire \frame[1] ;
 wire \frame[2] ;
 wire \frame[3] ;
 wire \frame[4] ;
 wire \frame[5] ;
 wire \frame[6] ;
 wire \hpos[0] ;
 wire \hpos[1] ;
 wire \hpos[2] ;
 wire \hpos[3] ;
 wire \hpos[4] ;
 wire \hpos[5] ;
 wire \hpos[6] ;
 wire \hpos[7] ;
 wire \hpos[8] ;
 wire \hpos[9] ;
 wire hsync;
 wire \hvsync_gen.vpos[0] ;
 wire \hvsync_gen.vpos[1] ;
 wire \hvsync_gen.vpos[2] ;
 wire \hvsync_gen.vpos[3] ;
 wire \hvsync_gen.vpos[4] ;
 wire \hvsync_gen.vpos[5] ;
 wire \hvsync_gen.vpos[6] ;
 wire \hvsync_gen.vpos[7] ;
 wire \hvsync_gen.vpos[8] ;
 wire \hvsync_gen.vpos[9] ;
 wire \hvsync_gen.vsync ;
 wire \palette_inst.palette[0] ;
 wire \palette_inst.palette[1] ;
 wire \palette_inst.palette[2] ;
 wire \palette_inst.palette[3] ;
 wire \palette_inst.palette[4] ;
 wire \palette_inst.palette[5] ;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire \waggle_demo.p0[1] ;
 wire \waggle_demo.p0[2] ;
 wire \waggle_demo.p0[3] ;
 wire \waggle_demo.p0[4] ;
 wire \waggle_demo.p0[5] ;
 wire \waggle_demo.p0[6] ;
 wire \waggle_demo.p0[7] ;
 wire \waggle_demo.p0[8] ;
 wire \waggle_demo.p0[9] ;
 wire \waggle_demo.p1[0] ;
 wire \waggle_demo.p1[1] ;
 wire \waggle_demo.p1[2] ;
 wire \waggle_demo.p1[3] ;
 wire \waggle_demo.p1[4] ;
 wire \waggle_demo.p1[5] ;
 wire \waggle_demo.p1[6] ;
 wire \waggle_demo.p1[7] ;
 wire \waggle_demo.p1[8] ;
 wire \waggle_demo.p1[9] ;
 wire \waggle_demo.xpos[0] ;
 wire \waggle_demo.xpos[1] ;
 wire \waggle_demo.xpos[2] ;
 wire \waggle_demo.xpos[3] ;
 wire \waggle_demo.xpos[4] ;
 wire \waggle_demo.xpos[5] ;
 wire \waggle_demo.xpos[6] ;
 wire \waggle_demo.xpos[7] ;
 wire \waggle_demo.ypos[1] ;
 wire \waggle_demo.ypos[2] ;
 wire \waggle_demo.ypos[3] ;
 wire \waggle_demo.ypos[4] ;
 wire \waggle_demo.ypos[5] ;
 wire \waggle_demo.ypos[6] ;
 wire \waggle_demo.ypos[7] ;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;

 sg13g2_a221oi_1 _1142_ (.B2(_0387_),
    .C1(net302),
    .B1(_0380_),
    .A1(_0337_),
    .Y(_0510_),
    .A2(_0338_));
 sg13g2_o21ai_1 _1143_ (.B1(_0341_),
    .Y(_0511_),
    .A1(net281),
    .A2(net280));
 sg13g2_nand2b_1 _1144_ (.Y(_0512_),
    .B(_0510_),
    .A_N(_0479_));
 sg13g2_o21ai_1 _1145_ (.B1(net296),
    .Y(_0513_),
    .A1(net290),
    .A2(_0355_));
 sg13g2_a21oi_1 _1146_ (.A1(net304),
    .A2(_0450_),
    .Y(_0514_),
    .B1(_0339_));
 sg13g2_nor3_1 _1147_ (.A(_0329_),
    .B(_0411_),
    .C(_0514_),
    .Y(_0515_));
 sg13g2_a221oi_1 _1148_ (.B2(_0515_),
    .C1(_0326_),
    .B1(_0512_),
    .A1(_0507_),
    .Y(_0516_),
    .A2(_0509_));
 sg13g2_nor2_1 _1149_ (.A(_0501_),
    .B(_0516_),
    .Y(_0517_));
 sg13g2_o21ai_1 _1150_ (.B1(_0366_),
    .Y(_0518_),
    .A1(_0501_),
    .A2(_0516_));
 sg13g2_nor2b_1 _1151_ (.A(_0486_),
    .B_N(_0518_),
    .Y(_0519_));
 sg13g2_o21ai_1 _1152_ (.B1(net293),
    .Y(_0520_),
    .A1(net287),
    .A2(net281));
 sg13g2_nand3_1 _1153_ (.B(_0435_),
    .C(_0520_),
    .A(net298),
    .Y(_0521_));
 sg13g2_a221oi_1 _1154_ (.B2(_0387_),
    .C1(net301),
    .B1(_0385_),
    .A1(net293),
    .Y(_0522_),
    .A2(_0381_));
 sg13g2_o21ai_1 _1155_ (.B1(_0521_),
    .Y(_0523_),
    .A1(_0341_),
    .A2(_0522_));
 sg13g2_nor2_1 _1156_ (.A(net304),
    .B(_0395_),
    .Y(_0524_));
 sg13g2_a221oi_1 _1157_ (.B2(_0524_),
    .C1(net306),
    .B1(_0478_),
    .A1(net296),
    .Y(_0525_),
    .A2(_0411_));
 sg13g2_o21ai_1 _1158_ (.B1(_0404_),
    .Y(_0526_),
    .A1(net281),
    .A2(net280));
 sg13g2_a221oi_1 _1159_ (.B2(_0341_),
    .C1(_0329_),
    .B1(_0526_),
    .A1(net280),
    .Y(_0527_),
    .A2(_0402_));
 sg13g2_a21o_1 _1160_ (.A2(_0525_),
    .A1(_0523_),
    .B1(_0527_),
    .X(_0528_));
 sg13g2_o21ai_1 _1161_ (.B1(_0510_),
    .Y(_0529_),
    .A1(net290),
    .A2(net287));
 sg13g2_o21ai_1 _1162_ (.B1(_0392_),
    .Y(_0530_),
    .A1(_0357_),
    .A2(_0382_));
 sg13g2_a22oi_1 _1163_ (.Y(_0531_),
    .B1(_0434_),
    .B2(_0391_),
    .A2(_0395_),
    .A1(_0381_));
 sg13g2_nand2b_1 _1164_ (.Y(_0532_),
    .B(_0402_),
    .A_N(_0531_));
 sg13g2_nor2_1 _1165_ (.A(net304),
    .B(net297),
    .Y(_0533_));
 sg13g2_nand2_1 _1166_ (.Y(_0534_),
    .A(net301),
    .B(net298));
 sg13g2_mux2_1 _1167_ (.A0(_0367_),
    .A1(_0534_),
    .S(_0530_),
    .X(_0535_));
 sg13g2_nand4_1 _1168_ (.B(_0529_),
    .C(_0532_),
    .A(net306),
    .Y(_0536_),
    .D(_0535_));
 sg13g2_xnor2_1 _1169_ (.Y(_0537_),
    .A(_0355_),
    .B(net282));
 sg13g2_o21ai_1 _1170_ (.B1(_0477_),
    .Y(_0538_),
    .A1(net292),
    .A2(_0537_));
 sg13g2_a221oi_1 _1171_ (.B2(_0416_),
    .C1(net304),
    .B1(_0475_),
    .A1(net291),
    .Y(_0539_),
    .A2(_0426_));
 sg13g2_o21ai_1 _1172_ (.B1(_0538_),
    .Y(_0540_),
    .A1(_0533_),
    .A2(_0539_));
 sg13g2_a221oi_1 _1173_ (.B2(_0357_),
    .C1(_0537_),
    .B1(net300),
    .A1(_0332_),
    .Y(_0541_),
    .A2(_0333_));
 sg13g2_nor2_1 _1174_ (.A(net307),
    .B(_0541_),
    .Y(_0542_));
 sg13g2_a21oi_1 _1175_ (.A1(_0540_),
    .A2(_0542_),
    .Y(_0543_),
    .B1(_0325_));
 sg13g2_a22oi_1 _1176_ (.Y(_0544_),
    .B1(_0536_),
    .B2(_0543_),
    .A2(_0528_),
    .A1(net308));
 sg13g2_or2_1 _1177_ (.X(_0545_),
    .B(_0544_),
    .A(_0365_));
 sg13g2_nand3b_1 _1178_ (.B(_0518_),
    .C(_0545_),
    .Y(_0546_),
    .A_N(_0486_));
 sg13g2_a21oi_1 _1179_ (.A1(net295),
    .A2(_0409_),
    .Y(_0547_),
    .B1(_0415_));
 sg13g2_nor2_1 _1180_ (.A(_0454_),
    .B(_0547_),
    .Y(_0548_));
 sg13g2_nand3_1 _1181_ (.B(net298),
    .C(_0435_),
    .A(net308),
    .Y(_0549_));
 sg13g2_a221oi_1 _1182_ (.B2(_0349_),
    .C1(_0548_),
    .B1(_0549_),
    .A1(net307),
    .Y(_0550_),
    .A2(_0511_));
 sg13g2_nor2_1 _1183_ (.A(_0387_),
    .B(_0420_),
    .Y(_0551_));
 sg13g2_a22oi_1 _1184_ (.Y(_0552_),
    .B1(_0551_),
    .B2(_0404_),
    .A2(_0435_),
    .A1(_0400_));
 sg13g2_nand2b_1 _1185_ (.Y(_0553_),
    .B(net296),
    .A_N(_0404_));
 sg13g2_nor2_1 _1186_ (.A(net301),
    .B(_0382_),
    .Y(_0554_));
 sg13g2_a21oi_1 _1187_ (.A1(_0553_),
    .A2(_0554_),
    .Y(_0555_),
    .B1(net306));
 sg13g2_o21ai_1 _1188_ (.B1(_0555_),
    .Y(_0556_),
    .A1(net303),
    .A2(_0552_));
 sg13g2_nand2b_1 _1189_ (.Y(_0557_),
    .B(_0392_),
    .A_N(_0513_));
 sg13g2_nand4_1 _1190_ (.B(net295),
    .C(_0392_),
    .A(net303),
    .Y(_0558_),
    .D(_0396_));
 sg13g2_nand2_1 _1191_ (.Y(_0559_),
    .A(net306),
    .B(_0558_));
 sg13g2_a221oi_1 _1192_ (.B2(_0384_),
    .C1(_0559_),
    .B1(_0557_),
    .A1(_0358_),
    .Y(_0560_),
    .A2(_0510_));
 sg13g2_nor2_1 _1193_ (.A(net308),
    .B(_0560_),
    .Y(_0561_));
 sg13g2_a21oi_1 _1194_ (.A1(_0556_),
    .A2(_0561_),
    .Y(_0562_),
    .B1(_0550_));
 sg13g2_and2_1 _1195_ (.A(_0366_),
    .B(_0562_),
    .X(_0563_));
 sg13g2_nor3_1 _1196_ (.A(_0414_),
    .B(_0546_),
    .C(_0563_),
    .Y(_0564_));
 sg13g2_o21ai_1 _1197_ (.B1(net306),
    .Y(_0565_),
    .A1(_0359_),
    .A2(_0384_));
 sg13g2_nor2_1 _1198_ (.A(_0399_),
    .B(_0454_),
    .Y(_0566_));
 sg13g2_nor2_1 _1199_ (.A(net308),
    .B(_0566_),
    .Y(_0567_));
 sg13g2_a22oi_1 _1200_ (.Y(_0568_),
    .B1(_0565_),
    .B2(_0567_),
    .A2(_0348_),
    .A1(net308));
 sg13g2_nor2_1 _1201_ (.A(_0365_),
    .B(_0564_),
    .Y(_0569_));
 sg13g2_a21o_2 _1202_ (.A2(_0568_),
    .A1(_0366_),
    .B1(_0569_),
    .X(_0570_));
 sg13g2_xnor2_1 _1203_ (.Y(_0571_),
    .A(_0361_),
    .B(_0570_));
 sg13g2_a21o_1 _1204_ (.A2(_0571_),
    .A1(_0272_),
    .B1(_0271_),
    .X(_0572_));
 sg13g2_nor2b_1 _1205_ (.A(\waggle_demo.ypos[6] ),
    .B_N(net346),
    .Y(_0573_));
 sg13g2_nand2b_1 _1206_ (.Y(_0574_),
    .B(\waggle_demo.ypos[6] ),
    .A_N(net346));
 sg13g2_nand2b_1 _1207_ (.Y(_0575_),
    .B(_0574_),
    .A_N(_0573_));
 sg13g2_nand2_1 _1208_ (.Y(_0576_),
    .A(_0349_),
    .B(_0570_));
 sg13g2_o21ai_1 _1209_ (.B1(_0576_),
    .Y(_0577_),
    .A1(_0349_),
    .A2(_0366_));
 sg13g2_xnor2_1 _1210_ (.Y(_0578_),
    .A(_0575_),
    .B(_0577_));
 sg13g2_and2_1 _1211_ (.A(_0572_),
    .B(_0578_),
    .X(_0579_));
 sg13g2_xor2_1 _1212_ (.B(_0578_),
    .A(_0572_),
    .X(_0580_));
 sg13g2_nand2_1 _1213_ (.Y(_0581_),
    .A(net349),
    .B(_0259_));
 sg13g2_xor2_1 _1214_ (.B(\waggle_demo.ypos[4] ),
    .A(net349),
    .X(_0582_));
 sg13g2_xnor2_1 _1215_ (.Y(_0583_),
    .A(_0568_),
    .B(_0569_));
 sg13g2_o21ai_1 _1216_ (.B1(_0581_),
    .Y(_0584_),
    .A1(_0582_),
    .A2(_0583_));
 sg13g2_xnor2_1 _1217_ (.Y(_0585_),
    .A(_0273_),
    .B(_0571_));
 sg13g2_nand2_1 _1218_ (.Y(_0586_),
    .A(_0584_),
    .B(_0585_));
 sg13g2_nand2b_1 _1219_ (.Y(_0587_),
    .B(net351),
    .A_N(\waggle_demo.ypos[3] ));
 sg13g2_xor2_1 _1220_ (.B(\waggle_demo.ypos[3] ),
    .A(net351),
    .X(_0588_));
 sg13g2_o21ai_1 _1221_ (.B1(_0414_),
    .Y(_0589_),
    .A1(_0546_),
    .A2(_0563_));
 sg13g2_nand2b_1 _1222_ (.Y(_0590_),
    .B(_0589_),
    .A_N(_0564_));
 sg13g2_o21ai_1 _1223_ (.B1(_0587_),
    .Y(_0591_),
    .A1(_0588_),
    .A2(_0590_));
 sg13g2_xor2_1 _1224_ (.B(_0583_),
    .A(_0582_),
    .X(_0592_));
 sg13g2_and2_1 _1225_ (.A(_0591_),
    .B(_0592_),
    .X(_0593_));
 sg13g2_nor2b_1 _1226_ (.A(\waggle_demo.ypos[2] ),
    .B_N(net352),
    .Y(_0594_));
 sg13g2_xnor2_1 _1227_ (.Y(_0595_),
    .A(net352),
    .B(\waggle_demo.ypos[2] ));
 sg13g2_xor2_1 _1228_ (.B(_0562_),
    .A(_0546_),
    .X(_0596_));
 sg13g2_a21oi_1 _1229_ (.A1(_0595_),
    .A2(_0596_),
    .Y(_0597_),
    .B1(_0594_));
 sg13g2_xnor2_1 _1230_ (.Y(_0598_),
    .A(_0588_),
    .B(_0590_));
 sg13g2_or2_1 _1231_ (.X(_0599_),
    .B(_0598_),
    .A(_0597_));
 sg13g2_nand2b_1 _1232_ (.Y(_0600_),
    .B(net353),
    .A_N(\waggle_demo.ypos[1] ));
 sg13g2_xor2_1 _1233_ (.B(\waggle_demo.ypos[1] ),
    .A(net353),
    .X(_0601_));
 sg13g2_xnor2_1 _1234_ (.Y(_0602_),
    .A(_0519_),
    .B(_0544_));
 sg13g2_o21ai_1 _1235_ (.B1(_0600_),
    .Y(_0603_),
    .A1(_0601_),
    .A2(_0602_));
 sg13g2_xor2_1 _1236_ (.B(_0596_),
    .A(_0595_),
    .X(_0604_));
 sg13g2_and2_1 _1237_ (.A(_0603_),
    .B(_0604_),
    .X(_0605_));
 sg13g2_xnor2_1 _1238_ (.Y(_0606_),
    .A(_0486_),
    .B(_0517_));
 sg13g2_nand2_1 _1239_ (.Y(_0607_),
    .A(net355),
    .B(_0606_));
 sg13g2_xnor2_1 _1240_ (.Y(_0608_),
    .A(_0601_),
    .B(_0602_));
 sg13g2_nand2_1 _1241_ (.Y(_0609_),
    .A(_0607_),
    .B(_0608_));
 sg13g2_xor2_1 _1242_ (.B(_0604_),
    .A(_0603_),
    .X(_0610_));
 sg13g2_a21oi_1 _1243_ (.A1(_0609_),
    .A2(_0610_),
    .Y(_0611_),
    .B1(_0605_));
 sg13g2_xnor2_1 _1244_ (.Y(_0612_),
    .A(_0597_),
    .B(_0598_));
 sg13g2_o21ai_1 _1245_ (.B1(_0599_),
    .Y(_0613_),
    .A1(_0611_),
    .A2(_0612_));
 sg13g2_xor2_1 _1246_ (.B(_0592_),
    .A(_0591_),
    .X(_0614_));
 sg13g2_a21oi_1 _1247_ (.A1(_0613_),
    .A2(_0614_),
    .Y(_0615_),
    .B1(_0593_));
 sg13g2_nor2_1 _1248_ (.A(_0584_),
    .B(_0585_),
    .Y(_0616_));
 sg13g2_a21oi_1 _1249_ (.A1(_0586_),
    .A2(_0615_),
    .Y(_0617_),
    .B1(_0616_));
 sg13g2_xnor2_1 _1250_ (.Y(_0618_),
    .A(_0580_),
    .B(_0617_));
 sg13g2_nor2b_1 _1251_ (.A(\waggle_demo.xpos[5] ),
    .B_N(net338),
    .Y(_0619_));
 sg13g2_nand2b_1 _1252_ (.Y(_0620_),
    .B(\waggle_demo.xpos[5] ),
    .A_N(net338));
 sg13g2_nand2b_1 _1253_ (.Y(_0621_),
    .B(_0620_),
    .A_N(_0619_));
 sg13g2_and2_1 _1254_ (.A(net354),
    .B(net1),
    .X(_0622_));
 sg13g2_nand2_2 _1255_ (.Y(_0623_),
    .A(net354),
    .B(net1));
 sg13g2_xnor2_1 _1256_ (.Y(_0624_),
    .A(\hvsync_gen.vpos[4] ),
    .B(\waggle_demo.p0[4] ));
 sg13g2_nor2_2 _1257_ (.A(net351),
    .B(\waggle_demo.p0[3] ),
    .Y(_0625_));
 sg13g2_and2_1 _1258_ (.A(net352),
    .B(\waggle_demo.p0[2] ),
    .X(_0626_));
 sg13g2_and2_1 _1259_ (.A(\hvsync_gen.vpos[1] ),
    .B(\waggle_demo.p0[1] ),
    .X(_0627_));
 sg13g2_xor2_1 _1260_ (.B(\waggle_demo.p0[2] ),
    .A(net352),
    .X(_0628_));
 sg13g2_a21oi_1 _1261_ (.A1(_0627_),
    .A2(_0628_),
    .Y(_0629_),
    .B1(_0626_));
 sg13g2_a221oi_1 _1262_ (.B2(_0628_),
    .C1(_0626_),
    .B1(_0627_),
    .A1(net350),
    .Y(_0630_),
    .A2(\waggle_demo.p0[3] ));
 sg13g2_nor3_1 _1263_ (.A(_0624_),
    .B(_0625_),
    .C(_0630_),
    .Y(_0631_));
 sg13g2_nor2_1 _1264_ (.A(net347),
    .B(\waggle_demo.p0[5] ),
    .Y(_0632_));
 sg13g2_xor2_1 _1265_ (.B(\waggle_demo.p0[5] ),
    .A(net347),
    .X(_0633_));
 sg13g2_and2_1 _1266_ (.A(\hvsync_gen.vpos[6] ),
    .B(\waggle_demo.p0[6] ),
    .X(_0634_));
 sg13g2_xor2_1 _1267_ (.B(\waggle_demo.p0[6] ),
    .A(net346),
    .X(_0635_));
 sg13g2_or2_1 _1268_ (.X(_0636_),
    .B(\waggle_demo.p0[7] ),
    .A(net345));
 sg13g2_and2_1 _1269_ (.A(net345),
    .B(\waggle_demo.p0[7] ),
    .X(_0637_));
 sg13g2_xor2_1 _1270_ (.B(\waggle_demo.p0[7] ),
    .A(net345),
    .X(_0638_));
 sg13g2_and2_1 _1271_ (.A(_0635_),
    .B(_0638_),
    .X(_0639_));
 sg13g2_nand3_1 _1272_ (.B(_0635_),
    .C(_0638_),
    .A(_0633_),
    .Y(_0640_));
 sg13g2_nor4_2 _1273_ (.A(_0624_),
    .B(_0625_),
    .C(_0630_),
    .Y(_0641_),
    .D(_0640_));
 sg13g2_or4_1 _1274_ (.A(_0624_),
    .B(_0625_),
    .C(_0630_),
    .D(_0640_),
    .X(_0642_));
 sg13g2_a21o_1 _1275_ (.A2(_0636_),
    .A1(_0634_),
    .B1(_0637_),
    .X(_0643_));
 sg13g2_a22oi_1 _1276_ (.Y(_0644_),
    .B1(\waggle_demo.p0[4] ),
    .B2(net349),
    .A2(\waggle_demo.p0[5] ),
    .A1(net347));
 sg13g2_nor2_1 _1277_ (.A(_0632_),
    .B(_0644_),
    .Y(_0645_));
 sg13g2_a221oi_1 _1278_ (.B2(_0645_),
    .C1(_0637_),
    .B1(_0639_),
    .A1(_0634_),
    .Y(_0646_),
    .A2(_0636_));
 sg13g2_a21o_1 _1279_ (.A2(_0645_),
    .A1(_0639_),
    .B1(_0643_),
    .X(_0647_));
 sg13g2_xor2_1 _1280_ (.B(\waggle_demo.p0[8] ),
    .A(\hvsync_gen.vpos[8] ),
    .X(_0648_));
 sg13g2_xnor2_1 _1281_ (.Y(_0649_),
    .A(\hvsync_gen.vpos[8] ),
    .B(\waggle_demo.p0[8] ));
 sg13g2_a21oi_1 _1282_ (.A1(_0642_),
    .A2(_0646_),
    .Y(_0650_),
    .B1(_0649_));
 sg13g2_o21ai_1 _1283_ (.B1(_0648_),
    .Y(_0651_),
    .A1(_0641_),
    .A2(_0647_));
 sg13g2_nor3_2 _1284_ (.A(_0641_),
    .B(_0647_),
    .C(_0648_),
    .Y(_0652_));
 sg13g2_nand3_1 _1285_ (.B(_0646_),
    .C(_0649_),
    .A(_0642_),
    .Y(_0653_));
 sg13g2_nand2_2 _1286_ (.Y(_0654_),
    .A(net336),
    .B(net335));
 sg13g2_a21oi_1 _1287_ (.A1(net349),
    .A2(\waggle_demo.p0[4] ),
    .Y(_0655_),
    .B1(_0631_));
 sg13g2_xor2_1 _1288_ (.B(_0655_),
    .A(_0633_),
    .X(_0656_));
 sg13g2_xor2_1 _1289_ (.B(_0656_),
    .A(_0654_),
    .X(_0657_));
 sg13g2_xnor2_1 _1290_ (.Y(_0658_),
    .A(_0654_),
    .B(_0656_));
 sg13g2_o21ai_1 _1291_ (.B1(_0624_),
    .Y(_0659_),
    .A1(_0625_),
    .A2(_0630_));
 sg13g2_nand2b_1 _1292_ (.Y(_0660_),
    .B(_0659_),
    .A_N(_0631_));
 sg13g2_o21ai_1 _1293_ (.B1(_0660_),
    .Y(_0661_),
    .A1(net337),
    .A2(_0652_));
 sg13g2_nand3b_1 _1294_ (.B(net335),
    .C(net336),
    .Y(_0662_),
    .A_N(_0660_));
 sg13g2_and2_1 _1295_ (.A(_0661_),
    .B(_0662_),
    .X(_0663_));
 sg13g2_nand2_1 _1296_ (.Y(_0664_),
    .A(_0661_),
    .B(_0662_));
 sg13g2_xor2_1 _1297_ (.B(\waggle_demo.p0[3] ),
    .A(net350),
    .X(_0665_));
 sg13g2_xnor2_1 _1298_ (.Y(_0666_),
    .A(_0629_),
    .B(_0665_));
 sg13g2_o21ai_1 _1299_ (.B1(_0666_),
    .Y(_0667_),
    .A1(net337),
    .A2(_0652_));
 sg13g2_or3_1 _1300_ (.A(net337),
    .B(_0652_),
    .C(_0666_),
    .X(_0668_));
 sg13g2_nand2_1 _1301_ (.Y(_0669_),
    .A(_0667_),
    .B(_0668_));
 sg13g2_and2_1 _1302_ (.A(_0667_),
    .B(_0668_),
    .X(_0670_));
 sg13g2_xor2_1 _1303_ (.B(\waggle_demo.p0[1] ),
    .A(\hvsync_gen.vpos[1] ),
    .X(_0671_));
 sg13g2_xnor2_1 _1304_ (.Y(_0672_),
    .A(\hvsync_gen.vpos[1] ),
    .B(\waggle_demo.p0[1] ));
 sg13g2_o21ai_1 _1305_ (.B1(_0672_),
    .Y(_0673_),
    .A1(net337),
    .A2(_0652_));
 sg13g2_nand3_1 _1306_ (.B(net335),
    .C(_0671_),
    .A(net336),
    .Y(_0674_));
 sg13g2_nand3_1 _1307_ (.B(net335),
    .C(_0672_),
    .A(net336),
    .Y(_0675_));
 sg13g2_o21ai_1 _1308_ (.B1(_0671_),
    .Y(_0676_),
    .A1(net337),
    .A2(_0652_));
 sg13g2_nand2_2 _1309_ (.Y(_0677_),
    .A(_0675_),
    .B(_0676_));
 sg13g2_nand2_2 _1310_ (.Y(_0678_),
    .A(_0673_),
    .B(_0674_));
 sg13g2_xor2_1 _1311_ (.B(_0628_),
    .A(_0627_),
    .X(_0679_));
 sg13g2_xnor2_1 _1312_ (.Y(_0680_),
    .A(_0627_),
    .B(_0628_));
 sg13g2_nand3_1 _1313_ (.B(net335),
    .C(_0679_),
    .A(net336),
    .Y(_0681_));
 sg13g2_o21ai_1 _1314_ (.B1(_0680_),
    .Y(_0682_),
    .A1(net337),
    .A2(_0652_));
 sg13g2_o21ai_1 _1315_ (.B1(_0679_),
    .Y(_0683_),
    .A1(net337),
    .A2(_0652_));
 sg13g2_nand3_1 _1316_ (.B(net335),
    .C(_0680_),
    .A(net336),
    .Y(_0684_));
 sg13g2_nand2_2 _1317_ (.Y(_0685_),
    .A(_0683_),
    .B(_0684_));
 sg13g2_nand2_2 _1318_ (.Y(_0686_),
    .A(_0681_),
    .B(_0682_));
 sg13g2_o21ai_1 _1319_ (.B1(net355),
    .Y(_0687_),
    .A1(net337),
    .A2(_0652_));
 sg13g2_nand3b_1 _1320_ (.B(_0651_),
    .C(_0653_),
    .Y(_0688_),
    .A_N(net355));
 sg13g2_a21o_1 _1321_ (.A2(net335),
    .A1(net336),
    .B1(net354),
    .X(_0689_));
 sg13g2_nand3_1 _1322_ (.B(net336),
    .C(net335),
    .A(net354),
    .Y(_0690_));
 sg13g2_nand2_1 _1323_ (.Y(_0691_),
    .A(_0689_),
    .B(_0690_));
 sg13g2_nand2_2 _1324_ (.Y(_0692_),
    .A(_0687_),
    .B(_0688_));
 sg13g2_nand4_1 _1325_ (.B(_0684_),
    .C(_0687_),
    .A(_0683_),
    .Y(_0693_),
    .D(_0688_));
 sg13g2_a22oi_1 _1326_ (.Y(_0694_),
    .B1(_0681_),
    .B2(_0682_),
    .A2(_0674_),
    .A1(_0673_));
 sg13g2_nand4_1 _1327_ (.B(_0676_),
    .C(_0683_),
    .A(_0675_),
    .Y(_0695_),
    .D(_0684_));
 sg13g2_nor2_2 _1328_ (.A(_0692_),
    .B(_0695_),
    .Y(_0696_));
 sg13g2_nand2_1 _1329_ (.Y(_0697_),
    .A(net314),
    .B(_0694_));
 sg13g2_a21oi_2 _1330_ (.B1(net316),
    .Y(_0698_),
    .A2(_0694_),
    .A1(net314));
 sg13g2_o21ai_1 _1331_ (.B1(net332),
    .Y(_0699_),
    .A1(net329),
    .A2(_0698_));
 sg13g2_a22oi_1 _1332_ (.Y(_0700_),
    .B1(_0687_),
    .B2(_0688_),
    .A2(_0676_),
    .A1(_0675_));
 sg13g2_nand4_1 _1333_ (.B(_0674_),
    .C(_0689_),
    .A(_0673_),
    .Y(_0701_),
    .D(_0690_));
 sg13g2_nand2_1 _1334_ (.Y(_0702_),
    .A(net320),
    .B(net315));
 sg13g2_nand3_1 _1335_ (.B(net315),
    .C(_0700_),
    .A(net320),
    .Y(_0703_));
 sg13g2_nor2_1 _1336_ (.A(net323),
    .B(_0703_),
    .Y(_0704_));
 sg13g2_nor2b_1 _1337_ (.A(_0631_),
    .B_N(_0644_),
    .Y(_0705_));
 sg13g2_nor2_1 _1338_ (.A(_0632_),
    .B(_0705_),
    .Y(_0706_));
 sg13g2_xnor2_1 _1339_ (.Y(_0707_),
    .A(_0635_),
    .B(_0706_));
 sg13g2_xor2_1 _1340_ (.B(_0707_),
    .A(_0654_),
    .X(_0708_));
 sg13g2_xnor2_1 _1341_ (.Y(_0709_),
    .A(_0654_),
    .B(_0707_));
 sg13g2_nor2_2 _1342_ (.A(net320),
    .B(net315),
    .Y(_0710_));
 sg13g2_a21oi_1 _1343_ (.A1(net323),
    .A2(_0710_),
    .Y(_0711_),
    .B1(net332));
 sg13g2_a22oi_1 _1344_ (.Y(_0712_),
    .B1(_0683_),
    .B2(_0684_),
    .A2(_0676_),
    .A1(_0675_));
 sg13g2_or2_1 _1345_ (.X(_0713_),
    .B(_0712_),
    .A(net320));
 sg13g2_inv_1 _1346_ (.Y(_0714_),
    .A(_0713_));
 sg13g2_nand2_1 _1347_ (.Y(_0715_),
    .A(net329),
    .B(_0713_));
 sg13g2_a21oi_1 _1348_ (.A1(_0711_),
    .A2(_0715_),
    .Y(_0716_),
    .B1(net312));
 sg13g2_o21ai_1 _1349_ (.B1(_0716_),
    .Y(_0717_),
    .A1(_0699_),
    .A2(_0704_));
 sg13g2_nand2_2 _1350_ (.Y(_0718_),
    .A(net332),
    .B(net312));
 sg13g2_nor2_1 _1351_ (.A(net320),
    .B(_0697_),
    .Y(_0719_));
 sg13g2_nand2_1 _1352_ (.Y(_0720_),
    .A(net316),
    .B(_0696_));
 sg13g2_nand2_2 _1353_ (.Y(_0721_),
    .A(net323),
    .B(net316));
 sg13g2_nor2_1 _1354_ (.A(_0697_),
    .B(_0721_),
    .Y(_0722_));
 sg13g2_or2_1 _1355_ (.X(_0723_),
    .B(_0721_),
    .A(_0697_));
 sg13g2_a21oi_1 _1356_ (.A1(net316),
    .A2(_0694_),
    .Y(_0724_),
    .B1(net323));
 sg13g2_nor2_1 _1357_ (.A(_0722_),
    .B(_0724_),
    .Y(_0725_));
 sg13g2_nor2_1 _1358_ (.A(_0718_),
    .B(_0725_),
    .Y(_0726_));
 sg13g2_a21oi_1 _1359_ (.A1(_0635_),
    .A2(_0706_),
    .Y(_0727_),
    .B1(_0634_));
 sg13g2_xnor2_1 _1360_ (.Y(_0728_),
    .A(_0638_),
    .B(_0654_));
 sg13g2_xnor2_1 _1361_ (.Y(_0729_),
    .A(_0727_),
    .B(_0728_));
 sg13g2_inv_2 _1362_ (.Y(_0730_),
    .A(net311));
 sg13g2_nor2_2 _1363_ (.A(net333),
    .B(net325),
    .Y(_0731_));
 sg13g2_nand2_1 _1364_ (.Y(_0732_),
    .A(net312),
    .B(_0731_));
 sg13g2_o21ai_1 _1365_ (.B1(_0730_),
    .Y(_0733_),
    .A1(_0719_),
    .A2(_0732_));
 sg13g2_nor2_1 _1366_ (.A(_0726_),
    .B(_0733_),
    .Y(_0734_));
 sg13g2_nand4_1 _1367_ (.B(_0682_),
    .C(_0689_),
    .A(_0681_),
    .Y(_0735_),
    .D(_0690_));
 sg13g2_nor2_2 _1368_ (.A(_0686_),
    .B(_0701_),
    .Y(_0736_));
 sg13g2_nand2_1 _1369_ (.Y(_0737_),
    .A(net315),
    .B(_0700_));
 sg13g2_a21oi_2 _1370_ (.B1(net320),
    .Y(_0738_),
    .A2(_0700_),
    .A1(net315));
 sg13g2_nor2_1 _1371_ (.A(net330),
    .B(_0738_),
    .Y(_0739_));
 sg13g2_nand2_1 _1372_ (.Y(_0740_),
    .A(net312),
    .B(_0729_));
 sg13g2_o21ai_1 _1373_ (.B1(net330),
    .Y(_0741_),
    .A1(net324),
    .A2(net316));
 sg13g2_a21oi_1 _1374_ (.A1(net329),
    .A2(_0739_),
    .Y(_0742_),
    .B1(_0740_));
 sg13g2_a22oi_1 _1375_ (.Y(_0743_),
    .B1(_0741_),
    .B2(_0742_),
    .A2(_0734_),
    .A1(_0717_));
 sg13g2_a21oi_1 _1376_ (.A1(\hvsync_gen.vpos[8] ),
    .A2(\waggle_demo.p0[8] ),
    .Y(_0744_),
    .B1(_0650_));
 sg13g2_xnor2_1 _1377_ (.Y(_0745_),
    .A(\hvsync_gen.vpos[9] ),
    .B(\waggle_demo.p0[9] ));
 sg13g2_xnor2_1 _1378_ (.Y(_0746_),
    .A(_0744_),
    .B(_0745_));
 sg13g2_inv_1 _1379_ (.Y(_0747_),
    .A(_0746_));
 sg13g2_a21oi_1 _1380_ (.A1(net326),
    .A2(net316),
    .Y(_0748_),
    .B1(_0677_));
 sg13g2_xor2_1 _1381_ (.B(_0654_),
    .A(_0064_),
    .X(_0749_));
 sg13g2_nor3_1 _1382_ (.A(net328),
    .B(_0678_),
    .C(_0749_),
    .Y(_0750_));
 sg13g2_nor4_1 _1383_ (.A(net328),
    .B(net322),
    .C(_0678_),
    .D(_0749_),
    .Y(_0751_));
 sg13g2_o21ai_1 _1384_ (.B1(_0686_),
    .Y(_0752_),
    .A1(_0748_),
    .A2(_0751_));
 sg13g2_and2_1 _1385_ (.A(net320),
    .B(_0712_),
    .X(_0753_));
 sg13g2_nand4_1 _1386_ (.B(_0662_),
    .C(_0667_),
    .A(_0661_),
    .Y(_0754_),
    .D(_0668_));
 sg13g2_nand4_1 _1387_ (.B(_0676_),
    .C(_0681_),
    .A(_0675_),
    .Y(_0755_),
    .D(_0682_));
 sg13g2_nand2_1 _1388_ (.Y(_0756_),
    .A(net326),
    .B(_0692_));
 sg13g2_a21oi_1 _1389_ (.A1(net329),
    .A2(_0753_),
    .Y(_0757_),
    .B1(net314));
 sg13g2_nand2b_1 _1390_ (.Y(_0758_),
    .B(_0754_),
    .A_N(_0755_));
 sg13g2_a21oi_1 _1391_ (.A1(net322),
    .A2(_0677_),
    .Y(_0759_),
    .B1(net328));
 sg13g2_o21ai_1 _1392_ (.B1(net317),
    .Y(_0760_),
    .A1(_0692_),
    .A2(_0755_));
 sg13g2_a22oi_1 _1393_ (.Y(_0761_),
    .B1(_0681_),
    .B2(_0682_),
    .A2(_0668_),
    .A1(_0667_));
 sg13g2_nor2_1 _1394_ (.A(net318),
    .B(_0693_),
    .Y(_0762_));
 sg13g2_nor2b_1 _1395_ (.A(_0712_),
    .B_N(_0735_),
    .Y(_0763_));
 sg13g2_nand2b_1 _1396_ (.Y(_0764_),
    .B(_0735_),
    .A_N(_0712_));
 sg13g2_xnor2_1 _1397_ (.Y(_0765_),
    .A(net354),
    .B(_0671_));
 sg13g2_inv_1 _1398_ (.Y(_0766_),
    .A(_0765_));
 sg13g2_nand3_1 _1399_ (.B(_0682_),
    .C(_0766_),
    .A(_0681_),
    .Y(_0767_));
 sg13g2_nor2_1 _1400_ (.A(net315),
    .B(_0766_),
    .Y(_0768_));
 sg13g2_nand3_1 _1401_ (.B(_0684_),
    .C(_0765_),
    .A(_0683_),
    .Y(_0769_));
 sg13g2_nand4_1 _1402_ (.B(_0674_),
    .C(_0683_),
    .A(_0673_),
    .Y(_0770_),
    .D(_0684_));
 sg13g2_a22oi_1 _1403_ (.Y(_0771_),
    .B1(_0758_),
    .B2(net314),
    .A2(_0757_),
    .A1(_0752_));
 sg13g2_xnor2_1 _1404_ (.Y(_0772_),
    .A(_0666_),
    .B(_0679_));
 sg13g2_a21oi_1 _1405_ (.A1(net326),
    .A2(_0695_),
    .Y(_0773_),
    .B1(net314));
 sg13g2_nand2_1 _1406_ (.Y(_0774_),
    .A(_0663_),
    .B(_0677_));
 sg13g2_a221oi_1 _1407_ (.B2(_0762_),
    .C1(net333),
    .B1(_0774_),
    .A1(_0772_),
    .Y(_0775_),
    .A2(_0773_));
 sg13g2_nor2_1 _1408_ (.A(net312),
    .B(_0775_),
    .Y(_0776_));
 sg13g2_o21ai_1 _1409_ (.B1(_0776_),
    .Y(_0777_),
    .A1(net330),
    .A2(_0771_));
 sg13g2_nand4_1 _1410_ (.B(_0684_),
    .C(_0689_),
    .A(_0683_),
    .Y(_0778_),
    .D(_0690_));
 sg13g2_nand3_1 _1411_ (.B(_0767_),
    .C(_0778_),
    .A(net317),
    .Y(_0779_));
 sg13g2_a21oi_1 _1412_ (.A1(net322),
    .A2(_0749_),
    .Y(_0780_),
    .B1(_0663_));
 sg13g2_nor3_1 _1413_ (.A(net324),
    .B(net319),
    .C(net314),
    .Y(_0781_));
 sg13g2_nand2b_1 _1414_ (.Y(_0782_),
    .B(_0692_),
    .A_N(_0755_));
 sg13g2_a21oi_1 _1415_ (.A1(_0686_),
    .A2(_0749_),
    .Y(_0783_),
    .B1(_0754_));
 sg13g2_a221oi_1 _1416_ (.B2(_0783_),
    .C1(_0781_),
    .B1(_0782_),
    .A1(_0779_),
    .Y(_0784_),
    .A2(_0780_));
 sg13g2_o21ai_1 _1417_ (.B1(net324),
    .Y(_0785_),
    .A1(net320),
    .A2(_0712_));
 sg13g2_a221oi_1 _1418_ (.B2(_0678_),
    .C1(net318),
    .B1(net314),
    .A1(_0683_),
    .Y(_0786_),
    .A2(_0684_));
 sg13g2_o21ai_1 _1419_ (.B1(_0785_),
    .Y(_0787_),
    .A1(_0738_),
    .A2(_0786_));
 sg13g2_o21ai_1 _1420_ (.B1(net333),
    .Y(_0788_),
    .A1(_0784_),
    .A2(_0787_));
 sg13g2_nor2_1 _1421_ (.A(net332),
    .B(_0781_),
    .Y(_0789_));
 sg13g2_a21oi_1 _1422_ (.A1(_0723_),
    .A2(_0789_),
    .Y(_0790_),
    .B1(_0708_));
 sg13g2_a21oi_1 _1423_ (.A1(_0788_),
    .A2(_0790_),
    .Y(_0791_),
    .B1(net311));
 sg13g2_nand3_1 _1424_ (.B(_0735_),
    .C(_0770_),
    .A(_0693_),
    .Y(_0792_));
 sg13g2_nand3_1 _1425_ (.B(_0695_),
    .C(_0767_),
    .A(net328),
    .Y(_0793_));
 sg13g2_xnor2_1 _1426_ (.Y(_0794_),
    .A(net321),
    .B(_0792_));
 sg13g2_nor2_1 _1427_ (.A(net331),
    .B(_0750_),
    .Y(_0795_));
 sg13g2_o21ai_1 _1428_ (.B1(_0795_),
    .Y(_0796_),
    .A1(_0793_),
    .A2(_0794_));
 sg13g2_a21oi_1 _1429_ (.A1(net315),
    .A2(_0749_),
    .Y(_0797_),
    .B1(_0754_));
 sg13g2_nand3_1 _1430_ (.B(_0677_),
    .C(net314),
    .A(net328),
    .Y(_0798_));
 sg13g2_nand2_1 _1431_ (.Y(_0799_),
    .A(net318),
    .B(_0677_));
 sg13g2_nor2_2 _1432_ (.A(net332),
    .B(net329),
    .Y(_0800_));
 sg13g2_nand2_1 _1433_ (.Y(_0801_),
    .A(net331),
    .B(net325));
 sg13g2_nand4_1 _1434_ (.B(_0756_),
    .C(_0798_),
    .A(_0693_),
    .Y(_0802_),
    .D(_0799_));
 sg13g2_o21ai_1 _1435_ (.B1(net313),
    .Y(_0803_),
    .A1(_0677_),
    .A2(_0797_));
 sg13g2_o21ai_1 _1436_ (.B1(_0718_),
    .Y(_0804_),
    .A1(_0802_),
    .A2(_0803_));
 sg13g2_a21oi_1 _1437_ (.A1(_0691_),
    .A2(_0694_),
    .Y(_0805_),
    .B1(net321));
 sg13g2_nand2_1 _1438_ (.Y(_0806_),
    .A(_0697_),
    .B(_0738_));
 sg13g2_and2_1 _1439_ (.A(_0702_),
    .B(_0759_),
    .X(_0807_));
 sg13g2_a21o_1 _1440_ (.A2(_0807_),
    .A1(_0806_),
    .B1(net330),
    .X(_0808_));
 sg13g2_nand4_1 _1441_ (.B(_0693_),
    .C(_0767_),
    .A(net317),
    .Y(_0809_),
    .D(_0770_));
 sg13g2_nand4_1 _1442_ (.B(_0678_),
    .C(_0685_),
    .A(net321),
    .Y(_0810_),
    .D(_0692_));
 sg13g2_nand3_1 _1443_ (.B(_0809_),
    .C(_0810_),
    .A(_0800_),
    .Y(_0811_));
 sg13g2_nand3_1 _1444_ (.B(_0770_),
    .C(_0778_),
    .A(net317),
    .Y(_0812_));
 sg13g2_nand4_1 _1445_ (.B(_0701_),
    .C(_0770_),
    .A(net318),
    .Y(_0813_),
    .D(_0778_));
 sg13g2_nand2b_1 _1446_ (.Y(_0814_),
    .B(net326),
    .A_N(_0813_));
 sg13g2_a21oi_1 _1447_ (.A1(_0731_),
    .A2(_0755_),
    .Y(_0815_),
    .B1(net313));
 sg13g2_and3_1 _1448_ (.X(_0816_),
    .A(_0811_),
    .B(_0814_),
    .C(_0815_));
 sg13g2_a221oi_1 _1449_ (.B2(_0816_),
    .C1(_0730_),
    .B1(_0808_),
    .A1(_0796_),
    .Y(_0817_),
    .A2(_0804_));
 sg13g2_a21oi_1 _1450_ (.A1(_0777_),
    .A2(_0791_),
    .Y(_0818_),
    .B1(_0817_));
 sg13g2_a21o_1 _1451_ (.A2(_0791_),
    .A1(_0777_),
    .B1(_0817_),
    .X(_0819_));
 sg13g2_o21ai_1 _1452_ (.B1(net321),
    .Y(_0820_),
    .A1(_0685_),
    .A2(_0700_));
 sg13g2_or2_1 _1453_ (.X(_0821_),
    .B(_0820_),
    .A(_0736_));
 sg13g2_o21ai_1 _1454_ (.B1(_0812_),
    .Y(_0822_),
    .A1(_0736_),
    .A2(_0820_));
 sg13g2_or2_1 _1455_ (.X(_0823_),
    .B(_0820_),
    .A(_0712_));
 sg13g2_nand2b_1 _1456_ (.Y(_0824_),
    .B(_0770_),
    .A_N(_0760_));
 sg13g2_nand3_1 _1457_ (.B(_0823_),
    .C(_0824_),
    .A(_0800_),
    .Y(_0825_));
 sg13g2_a21o_1 _1458_ (.A2(_0737_),
    .A1(_0695_),
    .B1(_0754_),
    .X(_0826_));
 sg13g2_and3_1 _1459_ (.X(_0827_),
    .A(net325),
    .B(_0755_),
    .C(_0770_));
 sg13g2_nand3_1 _1460_ (.B(_0755_),
    .C(_0770_),
    .A(net325),
    .Y(_0828_));
 sg13g2_nor3_1 _1461_ (.A(net325),
    .B(net317),
    .C(_0685_),
    .Y(_0829_));
 sg13g2_nor3_1 _1462_ (.A(net330),
    .B(_0827_),
    .C(_0829_),
    .Y(_0830_));
 sg13g2_a221oi_1 _1463_ (.B2(_0830_),
    .C1(_0708_),
    .B1(_0826_),
    .A1(_0731_),
    .Y(_0831_),
    .A2(_0822_));
 sg13g2_nand2b_2 _1464_ (.Y(_0832_),
    .B(_0800_),
    .A_N(_0786_));
 sg13g2_nand2b_1 _1465_ (.Y(_0833_),
    .B(_0806_),
    .A_N(_0832_));
 sg13g2_a21oi_1 _1466_ (.A1(net330),
    .A2(_0772_),
    .Y(_0834_),
    .B1(net324));
 sg13g2_nor3_1 _1467_ (.A(net313),
    .B(_0739_),
    .C(_0834_),
    .Y(_0835_));
 sg13g2_nand3_1 _1468_ (.B(_0695_),
    .C(_0765_),
    .A(net321),
    .Y(_0836_));
 sg13g2_nand3_1 _1469_ (.B(_0755_),
    .C(_0769_),
    .A(net317),
    .Y(_0837_));
 sg13g2_a21oi_1 _1470_ (.A1(net325),
    .A2(_0770_),
    .Y(_0838_),
    .B1(net333));
 sg13g2_nand3_1 _1471_ (.B(_0837_),
    .C(_0838_),
    .A(_0836_),
    .Y(_0839_));
 sg13g2_a21oi_1 _1472_ (.A1(net321),
    .A2(_0700_),
    .Y(_0840_),
    .B1(net331));
 sg13g2_o21ai_1 _1473_ (.B1(_0761_),
    .Y(_0841_),
    .A1(_0677_),
    .A2(_0692_));
 sg13g2_nand3_1 _1474_ (.B(net317),
    .C(_0694_),
    .A(net325),
    .Y(_0842_));
 sg13g2_nand4_1 _1475_ (.B(_0840_),
    .C(_0841_),
    .A(_0813_),
    .Y(_0843_),
    .D(_0842_));
 sg13g2_a21o_1 _1476_ (.A2(_0837_),
    .A1(_0836_),
    .B1(_0801_),
    .X(_0844_));
 sg13g2_nand3_1 _1477_ (.B(_0843_),
    .C(_0844_),
    .A(_0839_),
    .Y(_0845_));
 sg13g2_o21ai_1 _1478_ (.B1(_0759_),
    .Y(_0846_),
    .A1(_0760_),
    .A2(_0768_));
 sg13g2_a21oi_1 _1479_ (.A1(net321),
    .A2(_0765_),
    .Y(_0847_),
    .B1(net326));
 sg13g2_a21oi_1 _1480_ (.A1(_0799_),
    .A2(_0847_),
    .Y(_0848_),
    .B1(net331));
 sg13g2_nand3_1 _1481_ (.B(_0765_),
    .C(_0842_),
    .A(net313),
    .Y(_0849_));
 sg13g2_a22oi_1 _1482_ (.Y(_0850_),
    .B1(_0849_),
    .B2(_0718_),
    .A2(_0848_),
    .A1(_0846_));
 sg13g2_a221oi_1 _1483_ (.B2(_0835_),
    .C1(_0730_),
    .B1(_0833_),
    .A1(_0825_),
    .Y(_0851_),
    .A2(_0831_));
 sg13g2_a21o_1 _1484_ (.A2(_0845_),
    .A1(_0708_),
    .B1(_0850_),
    .X(_0852_));
 sg13g2_a21oi_2 _1485_ (.B1(_0851_),
    .Y(_0853_),
    .A2(_0852_),
    .A1(_0730_));
 sg13g2_a21oi_1 _1486_ (.A1(_0818_),
    .A2(_0853_),
    .Y(_0854_),
    .B1(_0746_));
 sg13g2_nand2_1 _1487_ (.Y(_0855_),
    .A(net317),
    .B(_0763_));
 sg13g2_a22oi_1 _1488_ (.Y(_0856_),
    .B1(_0828_),
    .B2(_0721_),
    .A2(_0805_),
    .A1(_0763_));
 sg13g2_nor3_1 _1489_ (.A(net321),
    .B(_0678_),
    .C(_0686_),
    .Y(_0857_));
 sg13g2_or4_1 _1490_ (.A(_0694_),
    .B(_0736_),
    .C(_0762_),
    .D(_0857_),
    .X(_0858_));
 sg13g2_a21oi_1 _1491_ (.A1(net328),
    .A2(_0858_),
    .Y(_0859_),
    .B1(_0856_));
 sg13g2_o21ai_1 _1492_ (.B1(_0711_),
    .Y(_0860_),
    .A1(_0696_),
    .A2(_0764_));
 sg13g2_nand2_1 _1493_ (.Y(_0861_),
    .A(net329),
    .B(_0738_));
 sg13g2_o21ai_1 _1494_ (.B1(net323),
    .Y(_0862_),
    .A1(_0714_),
    .A2(_0753_));
 sg13g2_nand3_1 _1495_ (.B(_0861_),
    .C(_0862_),
    .A(net332),
    .Y(_0863_));
 sg13g2_nand3_1 _1496_ (.B(_0820_),
    .C(_0855_),
    .A(net325),
    .Y(_0864_));
 sg13g2_o21ai_1 _1497_ (.B1(net328),
    .Y(_0865_),
    .A1(_0736_),
    .A2(_0805_));
 sg13g2_nand3_1 _1498_ (.B(_0864_),
    .C(_0865_),
    .A(net331),
    .Y(_0866_));
 sg13g2_nand3_1 _1499_ (.B(_0863_),
    .C(_0866_),
    .A(net311),
    .Y(_0867_));
 sg13g2_o21ai_1 _1500_ (.B1(_0860_),
    .Y(_0868_),
    .A1(net330),
    .A2(_0859_));
 sg13g2_a21oi_1 _1501_ (.A1(_0730_),
    .A2(_0868_),
    .Y(_0869_),
    .B1(_0708_));
 sg13g2_o21ai_1 _1502_ (.B1(_0737_),
    .Y(_0870_),
    .A1(_0698_),
    .A2(_0710_));
 sg13g2_xnor2_1 _1503_ (.Y(_0871_),
    .A(net323),
    .B(_0870_));
 sg13g2_a21oi_1 _1504_ (.A1(net316),
    .A2(net315),
    .Y(_0872_),
    .B1(_0832_));
 sg13g2_o21ai_1 _1505_ (.B1(_0821_),
    .Y(_0873_),
    .A1(_0696_),
    .A2(_0713_));
 sg13g2_a221oi_1 _1506_ (.B2(_0731_),
    .C1(_0872_),
    .B1(_0873_),
    .A1(net332),
    .Y(_0874_),
    .A2(_0871_));
 sg13g2_or2_1 _1507_ (.X(_0875_),
    .B(_0874_),
    .A(net311));
 sg13g2_or2_1 _1508_ (.X(_0876_),
    .B(_0786_),
    .A(_0719_));
 sg13g2_a221oi_1 _1509_ (.B2(_0876_),
    .C1(_0730_),
    .B1(_0800_),
    .A1(_0702_),
    .Y(_0877_),
    .A2(_0731_));
 sg13g2_nor2_1 _1510_ (.A(net312),
    .B(_0877_),
    .Y(_0878_));
 sg13g2_a22oi_1 _1511_ (.Y(_0879_),
    .B1(_0875_),
    .B2(_0878_),
    .A2(_0869_),
    .A1(_0867_));
 sg13g2_a21oi_1 _1512_ (.A1(_0747_),
    .A2(_0879_),
    .Y(_0880_),
    .B1(_0854_));
 sg13g2_nand3_1 _1513_ (.B(net316),
    .C(_0686_),
    .A(net328),
    .Y(_0881_));
 sg13g2_o21ai_1 _1514_ (.B1(_0698_),
    .Y(_0882_),
    .A1(net323),
    .A2(_0736_));
 sg13g2_a21oi_1 _1515_ (.A1(_0881_),
    .A2(_0882_),
    .Y(_0883_),
    .B1(net330));
 sg13g2_and3_1 _1516_ (.X(_0884_),
    .A(_0703_),
    .B(_0713_),
    .C(_0731_));
 sg13g2_o21ai_1 _1517_ (.B1(_0708_),
    .Y(_0885_),
    .A1(_0710_),
    .A2(_0832_));
 sg13g2_nor3_1 _1518_ (.A(_0883_),
    .B(_0884_),
    .C(_0885_),
    .Y(_0886_));
 sg13g2_a221oi_1 _1519_ (.B2(_0724_),
    .C1(_0718_),
    .B1(_0820_),
    .A1(_0720_),
    .Y(_0887_),
    .A2(_0807_));
 sg13g2_a21oi_1 _1520_ (.A1(net329),
    .A2(_0719_),
    .Y(_0888_),
    .B1(_0698_));
 sg13g2_nor3_1 _1521_ (.A(net332),
    .B(_0708_),
    .C(_0888_),
    .Y(_0889_));
 sg13g2_nor4_1 _1522_ (.A(net311),
    .B(_0886_),
    .C(_0887_),
    .D(_0889_),
    .Y(_0890_));
 sg13g2_o21ai_1 _1523_ (.B1(net311),
    .Y(_0891_),
    .A1(_0708_),
    .A2(_0741_));
 sg13g2_nand3_1 _1524_ (.B(net311),
    .C(_0820_),
    .A(net323),
    .Y(_0892_));
 sg13g2_a21oi_1 _1525_ (.A1(_0785_),
    .A2(_0861_),
    .Y(_0893_),
    .B1(_0718_));
 sg13g2_a221oi_1 _1526_ (.B2(_0892_),
    .C1(_0893_),
    .B1(_0891_),
    .A1(_0708_),
    .Y(_0894_),
    .A2(_0832_));
 sg13g2_or2_1 _1527_ (.X(_0895_),
    .B(_0894_),
    .A(_0890_));
 sg13g2_o21ai_1 _1528_ (.B1(_0880_),
    .Y(_0896_),
    .A1(_0746_),
    .A2(_0895_));
 sg13g2_xor2_1 _1529_ (.B(_0896_),
    .A(_0743_),
    .X(_0897_));
 sg13g2_a21o_1 _1530_ (.A2(_0819_),
    .A1(_0747_),
    .B1(_0853_),
    .X(_0898_));
 sg13g2_nand3_1 _1531_ (.B(_0819_),
    .C(_0853_),
    .A(_0747_),
    .Y(_0899_));
 sg13g2_and2_1 _1532_ (.A(_0898_),
    .B(_0899_),
    .X(_0900_));
 sg13g2_a21oi_1 _1533_ (.A1(_0898_),
    .A2(_0899_),
    .Y(_0901_),
    .B1(_0623_));
 sg13g2_xnor2_1 _1534_ (.Y(_0902_),
    .A(_0854_),
    .B(_0879_));
 sg13g2_a21oi_1 _1535_ (.A1(_0900_),
    .A2(_0902_),
    .Y(_0903_),
    .B1(_0623_));
 sg13g2_xnor2_1 _1536_ (.Y(_0904_),
    .A(_0880_),
    .B(_0895_));
 sg13g2_nor2b_1 _1537_ (.A(_0903_),
    .B_N(_0904_),
    .Y(_0905_));
 sg13g2_nor2_1 _1538_ (.A(_0623_),
    .B(_0905_),
    .Y(_0906_));
 sg13g2_a21oi_1 _1539_ (.A1(_0622_),
    .A2(_0897_),
    .Y(_0907_),
    .B1(_0906_));
 sg13g2_nand2_1 _1540_ (.Y(_0908_),
    .A(_0710_),
    .B(_0800_));
 sg13g2_a21oi_1 _1541_ (.A1(_0699_),
    .A2(_0908_),
    .Y(_0909_),
    .B1(net312));
 sg13g2_o21ai_1 _1542_ (.B1(_0730_),
    .Y(_0910_),
    .A1(_0718_),
    .A2(_0722_));
 sg13g2_o21ai_1 _1543_ (.B1(_0891_),
    .Y(_0911_),
    .A1(_0909_),
    .A2(_0910_));
 sg13g2_o21ai_1 _1544_ (.B1(_0747_),
    .Y(_0912_),
    .A1(_0743_),
    .A2(_0896_));
 sg13g2_xnor2_1 _1545_ (.Y(_0913_),
    .A(_0911_),
    .B(_0912_));
 sg13g2_o21ai_1 _1546_ (.B1(_0907_),
    .Y(_0914_),
    .A1(_0623_),
    .A2(_0913_));
 sg13g2_a21oi_1 _1547_ (.A1(_0710_),
    .A2(_0800_),
    .Y(_0915_),
    .B1(net312));
 sg13g2_o21ai_1 _1548_ (.B1(_0891_),
    .Y(_0916_),
    .A1(net311),
    .A2(_0915_));
 sg13g2_or2_1 _1549_ (.X(_0917_),
    .B(_0911_),
    .A(_0746_));
 sg13g2_and2_1 _1550_ (.A(_0912_),
    .B(_0917_),
    .X(_0918_));
 sg13g2_xor2_1 _1551_ (.B(_0918_),
    .A(_0916_),
    .X(_0919_));
 sg13g2_nor2_1 _1552_ (.A(_0914_),
    .B(_0919_),
    .Y(_0920_));
 sg13g2_xor2_1 _1553_ (.B(_0919_),
    .A(_0914_),
    .X(_0921_));
 sg13g2_a21oi_1 _1554_ (.A1(_0620_),
    .A2(_0921_),
    .Y(_0922_),
    .B1(_0619_));
 sg13g2_xnor2_1 _1555_ (.Y(_0923_),
    .A(\hpos[6] ),
    .B(\waggle_demo.xpos[6] ));
 sg13g2_nor2_1 _1556_ (.A(_0623_),
    .B(_0920_),
    .Y(_0924_));
 sg13g2_nor2_1 _1557_ (.A(_0891_),
    .B(_0912_),
    .Y(_0925_));
 sg13g2_a21oi_1 _1558_ (.A1(_0891_),
    .A2(_0918_),
    .Y(_0926_),
    .B1(_0925_));
 sg13g2_xnor2_1 _1559_ (.Y(_0927_),
    .A(_0924_),
    .B(_0926_));
 sg13g2_nor2b_1 _1560_ (.A(_0927_),
    .B_N(_0923_),
    .Y(_0928_));
 sg13g2_xor2_1 _1561_ (.B(_0927_),
    .A(_0923_),
    .X(_0929_));
 sg13g2_nor2_1 _1562_ (.A(_0922_),
    .B(_0929_),
    .Y(_0930_));
 sg13g2_xor2_1 _1563_ (.B(_0929_),
    .A(_0922_),
    .X(_0931_));
 sg13g2_nor2b_1 _1564_ (.A(\waggle_demo.xpos[4] ),
    .B_N(\hpos[4] ),
    .Y(_0932_));
 sg13g2_xor2_1 _1565_ (.B(\waggle_demo.xpos[4] ),
    .A(\hpos[4] ),
    .X(_0933_));
 sg13g2_xnor2_1 _1566_ (.Y(_0934_),
    .A(_0907_),
    .B(_0913_));
 sg13g2_nor2_1 _1567_ (.A(_0933_),
    .B(_0934_),
    .Y(_0935_));
 sg13g2_xnor2_1 _1568_ (.Y(_0936_),
    .A(_0621_),
    .B(_0921_));
 sg13g2_nor3_1 _1569_ (.A(_0932_),
    .B(_0935_),
    .C(_0936_),
    .Y(_0937_));
 sg13g2_o21ai_1 _1570_ (.B1(_0936_),
    .Y(_0938_),
    .A1(_0932_),
    .A2(_0935_));
 sg13g2_xor2_1 _1571_ (.B(\waggle_demo.xpos[3] ),
    .A(\hpos[3] ),
    .X(_0939_));
 sg13g2_xnor2_1 _1572_ (.Y(_0940_),
    .A(_0897_),
    .B(_0906_));
 sg13g2_nor2_1 _1573_ (.A(_0939_),
    .B(_0940_),
    .Y(_0941_));
 sg13g2_a21oi_1 _1574_ (.A1(\hpos[3] ),
    .A2(_0254_),
    .Y(_0942_),
    .B1(_0941_));
 sg13g2_xor2_1 _1575_ (.B(_0934_),
    .A(_0933_),
    .X(_0943_));
 sg13g2_nand2b_1 _1576_ (.Y(_0944_),
    .B(_0943_),
    .A_N(_0942_));
 sg13g2_xor2_1 _1577_ (.B(\waggle_demo.xpos[2] ),
    .A(\hpos[2] ),
    .X(_0945_));
 sg13g2_xor2_1 _1578_ (.B(_0904_),
    .A(_0903_),
    .X(_0946_));
 sg13g2_nor2_1 _1579_ (.A(_0945_),
    .B(_0946_),
    .Y(_0947_));
 sg13g2_a21oi_2 _1580_ (.B1(_0947_),
    .Y(_0948_),
    .A2(_0255_),
    .A1(\hpos[2] ));
 sg13g2_xnor2_1 _1581_ (.Y(_0949_),
    .A(_0939_),
    .B(_0940_));
 sg13g2_nor2_1 _1582_ (.A(_0948_),
    .B(_0949_),
    .Y(_0950_));
 sg13g2_nor2b_1 _1583_ (.A(\waggle_demo.xpos[1] ),
    .B_N(\hpos[1] ),
    .Y(_0951_));
 sg13g2_xnor2_1 _1584_ (.Y(_0952_),
    .A(\hpos[1] ),
    .B(\waggle_demo.xpos[1] ));
 sg13g2_xnor2_1 _1585_ (.Y(_0953_),
    .A(_0901_),
    .B(_0902_));
 sg13g2_a21o_1 _1586_ (.A2(_0953_),
    .A1(_0952_),
    .B1(_0951_),
    .X(_0954_));
 sg13g2_xor2_1 _1587_ (.B(_0946_),
    .A(_0945_),
    .X(_0955_));
 sg13g2_nand2_1 _1588_ (.Y(_0956_),
    .A(\waggle_demo.xpos[0] ),
    .B(_0900_));
 sg13g2_xnor2_1 _1589_ (.Y(_0957_),
    .A(_0952_),
    .B(_0953_));
 sg13g2_nand2b_1 _1590_ (.Y(_0958_),
    .B(_0956_),
    .A_N(_0957_));
 sg13g2_xor2_1 _1591_ (.B(_0900_),
    .A(_0066_),
    .X(_0959_));
 sg13g2_nand2_1 _1592_ (.Y(_0960_),
    .A(\hpos[0] ),
    .B(_0959_));
 sg13g2_xnor2_1 _1593_ (.Y(_0961_),
    .A(_0956_),
    .B(_0957_));
 sg13g2_nand2b_1 _1594_ (.Y(_0962_),
    .B(_0961_),
    .A_N(_0960_));
 sg13g2_xnor2_1 _1595_ (.Y(_0963_),
    .A(_0954_),
    .B(_0955_));
 sg13g2_a21oi_1 _1596_ (.A1(_0958_),
    .A2(_0962_),
    .Y(_0964_),
    .B1(_0963_));
 sg13g2_a21o_1 _1597_ (.A2(_0955_),
    .A1(_0954_),
    .B1(_0964_),
    .X(_0965_));
 sg13g2_xor2_1 _1598_ (.B(_0949_),
    .A(_0948_),
    .X(_0966_));
 sg13g2_a21oi_1 _1599_ (.A1(_0965_),
    .A2(_0966_),
    .Y(_0967_),
    .B1(_0950_));
 sg13g2_xor2_1 _1600_ (.B(_0943_),
    .A(_0942_),
    .X(_0968_));
 sg13g2_o21ai_1 _1601_ (.B1(_0944_),
    .Y(_0969_),
    .A1(_0967_),
    .A2(_0968_));
 sg13g2_nor2b_1 _1602_ (.A(_0969_),
    .B_N(_0938_),
    .Y(_0970_));
 sg13g2_nor2_1 _1603_ (.A(_0937_),
    .B(_0970_),
    .Y(_0971_));
 sg13g2_xnor2_1 _1604_ (.Y(_0972_),
    .A(_0931_),
    .B(_0971_));
 sg13g2_xnor2_1 _1605_ (.Y(_0973_),
    .A(_0618_),
    .B(_0972_));
 sg13g2_xnor2_1 _1606_ (.Y(_0974_),
    .A(_0613_),
    .B(_0614_));
 sg13g2_xnor2_1 _1607_ (.Y(_0975_),
    .A(_0967_),
    .B(_0968_));
 sg13g2_xor2_1 _1608_ (.B(_0975_),
    .A(_0974_),
    .X(_0976_));
 sg13g2_nor2b_1 _1609_ (.A(_0009_),
    .B_N(_0976_),
    .Y(_0977_));
 sg13g2_xnor2_1 _1610_ (.Y(_0978_),
    .A(_0611_),
    .B(_0612_));
 sg13g2_xnor2_1 _1611_ (.Y(_0979_),
    .A(_0965_),
    .B(_0966_));
 sg13g2_xnor2_1 _1612_ (.Y(_0980_),
    .A(_0978_),
    .B(_0979_));
 sg13g2_or2_1 _1613_ (.X(_0981_),
    .B(_0980_),
    .A(_0016_));
 sg13g2_xnor2_1 _1614_ (.Y(_0982_),
    .A(_0609_),
    .B(_0610_));
 sg13g2_nand3_1 _1615_ (.B(_0962_),
    .C(_0963_),
    .A(_0958_),
    .Y(_0983_));
 sg13g2_nor2b_1 _1616_ (.A(_0964_),
    .B_N(_0983_),
    .Y(_0984_));
 sg13g2_xnor2_1 _1617_ (.Y(_0985_),
    .A(_0982_),
    .B(_0984_));
 sg13g2_nor2b_1 _1618_ (.A(_0024_),
    .B_N(_0985_),
    .Y(_0986_));
 sg13g2_xnor2_1 _1619_ (.Y(_0987_),
    .A(_0960_),
    .B(_0961_));
 sg13g2_xor2_1 _1620_ (.B(_0608_),
    .A(_0607_),
    .X(_0988_));
 sg13g2_xnor2_1 _1621_ (.Y(_0989_),
    .A(_0987_),
    .B(_0988_));
 sg13g2_nor2b_1 _1622_ (.A(_0065_),
    .B_N(_0989_),
    .Y(_0990_));
 sg13g2_xnor2_1 _1623_ (.Y(_0991_),
    .A(_0024_),
    .B(_0985_));
 sg13g2_a21oi_1 _1624_ (.A1(_0990_),
    .A2(_0991_),
    .Y(_0992_),
    .B1(_0986_));
 sg13g2_and2_1 _1625_ (.A(_0016_),
    .B(_0980_),
    .X(_0993_));
 sg13g2_xor2_1 _1626_ (.B(_0980_),
    .A(_0016_),
    .X(_0994_));
 sg13g2_o21ai_1 _1627_ (.B1(_0981_),
    .Y(_0995_),
    .A1(_0992_),
    .A2(_0993_));
 sg13g2_xnor2_1 _1628_ (.Y(_0996_),
    .A(_0009_),
    .B(_0976_));
 sg13g2_a21oi_2 _1629_ (.B1(_0977_),
    .Y(_0997_),
    .A2(_0996_),
    .A1(_0995_));
 sg13g2_nand2b_1 _1630_ (.Y(_0998_),
    .B(_0938_),
    .A_N(_0937_));
 sg13g2_xnor2_1 _1631_ (.Y(_0999_),
    .A(_0615_),
    .B(_0998_));
 sg13g2_xnor2_1 _1632_ (.Y(_1000_),
    .A(_0584_),
    .B(_0585_));
 sg13g2_xnor2_1 _1633_ (.Y(_1001_),
    .A(_0969_),
    .B(_1000_));
 sg13g2_xnor2_1 _1634_ (.Y(_1002_),
    .A(_0999_),
    .B(_1001_));
 sg13g2_xnor2_1 _1635_ (.Y(_1003_),
    .A(\frame[4] ),
    .B(_1002_));
 sg13g2_nor2_1 _1636_ (.A(_0997_),
    .B(_1003_),
    .Y(_1004_));
 sg13g2_xnor2_1 _1637_ (.Y(_1005_),
    .A(\frame[5] ),
    .B(_0973_));
 sg13g2_nand2_1 _1638_ (.Y(_1006_),
    .A(_0010_),
    .B(_0973_));
 sg13g2_nand2b_1 _1639_ (.Y(_1007_),
    .B(_1002_),
    .A_N(_0011_));
 sg13g2_o21ai_1 _1640_ (.B1(_1007_),
    .Y(_1008_),
    .A1(_0010_),
    .A2(_0973_));
 sg13g2_a22oi_1 _1641_ (.Y(_1009_),
    .B1(_1006_),
    .B2(_1008_),
    .A2(_1005_),
    .A1(_1004_));
 sg13g2_a21oi_1 _1642_ (.A1(_0580_),
    .A2(_0617_),
    .Y(_1010_),
    .B1(_0579_));
 sg13g2_xor2_1 _1643_ (.B(_1010_),
    .A(\frame[6] ),
    .X(_1011_));
 sg13g2_a21oi_1 _1644_ (.A1(_0931_),
    .A2(_0971_),
    .Y(_1012_),
    .B1(_0930_));
 sg13g2_a21oi_1 _1645_ (.A1(\hpos[6] ),
    .A2(_0260_),
    .Y(_1013_),
    .B1(_0928_));
 sg13g2_a21oi_1 _1646_ (.A1(_0622_),
    .A2(_0926_),
    .Y(_1014_),
    .B1(_0924_));
 sg13g2_xor2_1 _1647_ (.B(\waggle_demo.ypos[7] ),
    .A(net345),
    .X(_1015_));
 sg13g2_xnor2_1 _1648_ (.Y(_1016_),
    .A(\hpos[7] ),
    .B(\waggle_demo.xpos[7] ));
 sg13g2_xnor2_1 _1649_ (.Y(_1017_),
    .A(_1015_),
    .B(_1016_));
 sg13g2_xnor2_1 _1650_ (.Y(_1018_),
    .A(_0918_),
    .B(_1017_));
 sg13g2_xnor2_1 _1651_ (.Y(_1019_),
    .A(_0570_),
    .B(_1018_));
 sg13g2_xnor2_1 _1652_ (.Y(_1020_),
    .A(_1014_),
    .B(_1019_));
 sg13g2_a21oi_1 _1653_ (.A1(_0574_),
    .A2(_0577_),
    .Y(_1021_),
    .B1(_0573_));
 sg13g2_xnor2_1 _1654_ (.Y(_1022_),
    .A(_1020_),
    .B(_1021_));
 sg13g2_xnor2_1 _1655_ (.Y(_1023_),
    .A(_1013_),
    .B(_1022_));
 sg13g2_xnor2_1 _1656_ (.Y(_1024_),
    .A(_1012_),
    .B(_1023_));
 sg13g2_xor2_1 _1657_ (.B(_1024_),
    .A(_1011_),
    .X(_1025_));
 sg13g2_xnor2_1 _1658_ (.Y(_1026_),
    .A(_1009_),
    .B(_1025_));
 sg13g2_xor2_1 _1659_ (.B(_1025_),
    .A(_1009_),
    .X(_1027_));
 sg13g2_xor2_1 _1660_ (.B(_1003_),
    .A(_0997_),
    .X(_1028_));
 sg13g2_xnor2_1 _1661_ (.Y(_1029_),
    .A(_0997_),
    .B(_1003_));
 sg13g2_xnor2_1 _1662_ (.Y(_1030_),
    .A(_0995_),
    .B(_0996_));
 sg13g2_inv_1 _1663_ (.Y(_1031_),
    .A(_1030_));
 sg13g2_xnor2_1 _1664_ (.Y(_1032_),
    .A(_0992_),
    .B(_0994_));
 sg13g2_xor2_1 _1665_ (.B(_0991_),
    .A(_0990_),
    .X(_1033_));
 sg13g2_xnor2_1 _1666_ (.Y(_1034_),
    .A(\frame[0] ),
    .B(_0989_));
 sg13g2_inv_1 _1667_ (.Y(_1035_),
    .A(_1034_));
 sg13g2_xor2_1 _1668_ (.B(_0959_),
    .A(\hpos[0] ),
    .X(_1036_));
 sg13g2_xor2_1 _1669_ (.B(_0606_),
    .A(net355),
    .X(_1037_));
 sg13g2_xnor2_1 _1670_ (.Y(_1038_),
    .A(_1036_),
    .B(_1037_));
 sg13g2_nand2_1 _1671_ (.Y(_1039_),
    .A(_1034_),
    .B(_1038_));
 sg13g2_a21o_1 _1672_ (.A2(_1039_),
    .A1(_1033_),
    .B1(_1032_),
    .X(_1040_));
 sg13g2_a21oi_1 _1673_ (.A1(_1031_),
    .A2(_1040_),
    .Y(_1041_),
    .B1(_1028_));
 sg13g2_xor2_1 _1674_ (.B(_0973_),
    .A(_0010_),
    .X(_1042_));
 sg13g2_o21ai_1 _1675_ (.B1(_1007_),
    .Y(_1043_),
    .A1(_0997_),
    .A2(_1003_));
 sg13g2_xor2_1 _1676_ (.B(_1043_),
    .A(_1042_),
    .X(_1044_));
 sg13g2_xnor2_1 _1677_ (.Y(_1045_),
    .A(_1042_),
    .B(_1043_));
 sg13g2_nor2_1 _1678_ (.A(_1034_),
    .B(_1038_),
    .Y(_1046_));
 sg13g2_a21oi_1 _1679_ (.A1(_1033_),
    .A2(_1046_),
    .Y(_1047_),
    .B1(_1032_));
 sg13g2_nand3_1 _1680_ (.B(_1030_),
    .C(_1047_),
    .A(_1029_),
    .Y(_1048_));
 sg13g2_nand2_1 _1681_ (.Y(_1049_),
    .A(_1044_),
    .B(_1048_));
 sg13g2_nand3_1 _1682_ (.B(_1044_),
    .C(_1048_),
    .A(_1041_),
    .Y(_1050_));
 sg13g2_or2_1 _1683_ (.X(_1051_),
    .B(_1033_),
    .A(_1032_));
 sg13g2_or2_1 _1684_ (.X(_1052_),
    .B(_1051_),
    .A(_1035_));
 sg13g2_nand3_1 _1685_ (.B(_1031_),
    .C(_1052_),
    .A(_1028_),
    .Y(_1053_));
 sg13g2_nor2_1 _1686_ (.A(_1045_),
    .B(_1053_),
    .Y(_1054_));
 sg13g2_nor2b_1 _1687_ (.A(_1051_),
    .B_N(_1030_),
    .Y(_1055_));
 sg13g2_nor2_1 _1688_ (.A(_1029_),
    .B(_1055_),
    .Y(_1056_));
 sg13g2_or3_1 _1689_ (.A(_1041_),
    .B(_1045_),
    .C(_1056_),
    .X(_1057_));
 sg13g2_nand2b_1 _1690_ (.Y(_1058_),
    .B(_1057_),
    .A_N(_1054_));
 sg13g2_nand2_1 _1691_ (.Y(_1059_),
    .A(net279),
    .B(_1054_));
 sg13g2_a21o_1 _1692_ (.A2(_1057_),
    .A1(_1050_),
    .B1(_1026_),
    .X(_1060_));
 sg13g2_and3_1 _1693_ (.X(_1061_),
    .A(_1044_),
    .B(_1053_),
    .C(_1056_));
 sg13g2_nand2_1 _1694_ (.Y(_1062_),
    .A(_1026_),
    .B(_1061_));
 sg13g2_nand2_1 _1695_ (.Y(_1063_),
    .A(_1027_),
    .B(_1049_));
 sg13g2_and4_1 _1696_ (.A(_1059_),
    .B(_1060_),
    .C(_1062_),
    .D(_1063_),
    .X(_0002_));
 sg13g2_and2_1 _1697_ (.A(_1032_),
    .B(_1033_),
    .X(_1064_));
 sg13g2_a21oi_2 _1698_ (.B1(_1028_),
    .Y(_1065_),
    .A2(_1064_),
    .A1(_1031_));
 sg13g2_o21ai_1 _1699_ (.B1(_1032_),
    .Y(_1066_),
    .A1(_1033_),
    .A2(_1046_));
 sg13g2_a21oi_2 _1700_ (.B1(_1029_),
    .Y(_1067_),
    .A2(_1066_),
    .A1(_1030_));
 sg13g2_nor3_1 _1701_ (.A(_1044_),
    .B(_1065_),
    .C(_1067_),
    .Y(_1068_));
 sg13g2_or2_1 _1702_ (.X(_1069_),
    .B(_1039_),
    .A(_1033_));
 sg13g2_nand4_1 _1703_ (.B(_1031_),
    .C(_1032_),
    .A(_1028_),
    .Y(_1070_),
    .D(_1069_));
 sg13g2_and3_1 _1704_ (.X(_0087_),
    .A(_1045_),
    .B(_1067_),
    .C(_1070_));
 sg13g2_nand3_1 _1705_ (.B(_1067_),
    .C(_1070_),
    .A(_1045_),
    .Y(_0088_));
 sg13g2_nand2_1 _1706_ (.Y(_0089_),
    .A(_1050_),
    .B(_0088_));
 sg13g2_o21ai_1 _1707_ (.B1(_1026_),
    .Y(_0090_),
    .A1(_1068_),
    .A2(_0089_));
 sg13g2_nand3_1 _1708_ (.B(_1045_),
    .C(_1065_),
    .A(_1026_),
    .Y(_0091_));
 sg13g2_and3_1 _1709_ (.X(_0092_),
    .A(_1059_),
    .B(_1062_),
    .C(_0091_));
 sg13g2_mux2_1 _1710_ (.A0(_1048_),
    .A1(_1070_),
    .S(_1045_),
    .X(_0093_));
 sg13g2_a21o_1 _1711_ (.A2(_0093_),
    .A1(_1057_),
    .B1(net279),
    .X(_0094_));
 sg13g2_nand3_1 _1712_ (.B(_0092_),
    .C(_0094_),
    .A(_0090_),
    .Y(_0003_));
 sg13g2_nand2_1 _1713_ (.Y(_0095_),
    .A(net279),
    .B(_1061_));
 sg13g2_o21ai_1 _1714_ (.B1(net279),
    .Y(_0096_),
    .A1(_1061_),
    .A2(_0087_));
 sg13g2_nand2b_1 _1715_ (.Y(_0097_),
    .B(net279),
    .A_N(_0093_));
 sg13g2_and4_1 _1716_ (.A(_1059_),
    .B(_1060_),
    .C(_0096_),
    .D(_0097_),
    .X(_0098_));
 sg13g2_nand3_1 _1717_ (.B(_1033_),
    .C(_1035_),
    .A(_1032_),
    .Y(_0099_));
 sg13g2_nand3_1 _1718_ (.B(_1030_),
    .C(_0099_),
    .A(_1029_),
    .Y(_0100_));
 sg13g2_nand4_1 _1719_ (.B(_1045_),
    .C(_1065_),
    .A(net279),
    .Y(_0101_),
    .D(_0100_));
 sg13g2_o21ai_1 _1720_ (.B1(_0100_),
    .Y(_0102_),
    .A1(_1065_),
    .A2(_1067_));
 sg13g2_nand3_1 _1721_ (.B(_1045_),
    .C(_0102_),
    .A(_1026_),
    .Y(_0103_));
 sg13g2_nand3_1 _1722_ (.B(_0101_),
    .C(_0103_),
    .A(_0098_),
    .Y(_0004_));
 sg13g2_nand2_1 _1723_ (.Y(_0104_),
    .A(net279),
    .B(_1068_));
 sg13g2_nand3_1 _1724_ (.B(_0098_),
    .C(_0104_),
    .A(_0091_),
    .Y(_0005_));
 sg13g2_and2_1 _1725_ (.A(_0091_),
    .B(_0095_),
    .X(_0105_));
 sg13g2_nand2_1 _1726_ (.Y(_0106_),
    .A(_1027_),
    .B(_1058_));
 sg13g2_and4_1 _1727_ (.A(_0090_),
    .B(_0097_),
    .C(_0105_),
    .D(_0106_),
    .X(_0006_));
 sg13g2_xnor2_1 _1728_ (.Y(_0007_),
    .A(net279),
    .B(_1049_));
 sg13g2_nor2_1 _1729_ (.A(net3),
    .B(net2),
    .Y(_0107_));
 sg13g2_nor3_2 _1730_ (.A(net359),
    .B(net3),
    .C(net2),
    .Y(_0108_));
 sg13g2_nand2_1 _1731_ (.Y(_0109_),
    .A(\waggle_demo.p0[1] ),
    .B(_0108_));
 sg13g2_nor2b_1 _1732_ (.A(net3),
    .B_N(net2),
    .Y(_0110_));
 sg13g2_nor2b_1 _1733_ (.A(net359),
    .B_N(_0110_),
    .Y(_0111_));
 sg13g2_nand2_1 _1734_ (.Y(_0112_),
    .A(\waggle_demo.p0[2] ),
    .B(_0111_));
 sg13g2_xnor2_1 _1735_ (.Y(_0113_),
    .A(\waggle_demo.p0[2] ),
    .B(_0111_));
 sg13g2_xor2_1 _1736_ (.B(_0113_),
    .A(_0109_),
    .X(_0032_));
 sg13g2_o21ai_1 _1737_ (.B1(_0112_),
    .Y(_0114_),
    .A1(_0109_),
    .A2(_0113_));
 sg13g2_nor2b_1 _1738_ (.A(net2),
    .B_N(net3),
    .Y(_0115_));
 sg13g2_nand2b_1 _1739_ (.Y(_0116_),
    .B(net3),
    .A_N(net2));
 sg13g2_nor3_1 _1740_ (.A(net359),
    .B(_0012_),
    .C(_0116_),
    .Y(_0117_));
 sg13g2_o21ai_1 _1741_ (.B1(_0012_),
    .Y(_0118_),
    .A1(net359),
    .A2(_0116_));
 sg13g2_nor2b_1 _1742_ (.A(_0117_),
    .B_N(_0118_),
    .Y(_0119_));
 sg13g2_xor2_1 _1743_ (.B(_0119_),
    .A(_0114_),
    .X(_0033_));
 sg13g2_a21oi_1 _1744_ (.A1(_0114_),
    .A2(_0119_),
    .Y(_0120_),
    .B1(_0117_));
 sg13g2_nand2_1 _1745_ (.Y(_0121_),
    .A(net3),
    .B(net2));
 sg13g2_nor2_1 _1746_ (.A(net358),
    .B(_0121_),
    .Y(_0122_));
 sg13g2_xor2_1 _1747_ (.B(_0122_),
    .A(\waggle_demo.p0[4] ),
    .X(_0123_));
 sg13g2_nor2b_1 _1748_ (.A(_0120_),
    .B_N(_0123_),
    .Y(_0124_));
 sg13g2_xnor2_1 _1749_ (.Y(_0034_),
    .A(_0120_),
    .B(_0123_));
 sg13g2_a21o_1 _1750_ (.A2(_0122_),
    .A1(\waggle_demo.p0[4] ),
    .B1(_0124_),
    .X(_0125_));
 sg13g2_nand2_1 _1751_ (.Y(_0126_),
    .A(net358),
    .B(_0107_));
 sg13g2_nor2_1 _1752_ (.A(_0013_),
    .B(_0126_),
    .Y(_0127_));
 sg13g2_xor2_1 _1753_ (.B(_0126_),
    .A(_0013_),
    .X(_0128_));
 sg13g2_xor2_1 _1754_ (.B(_0128_),
    .A(_0125_),
    .X(_0035_));
 sg13g2_a21oi_1 _1755_ (.A1(_0125_),
    .A2(_0128_),
    .Y(_0129_),
    .B1(_0127_));
 sg13g2_nand3_1 _1756_ (.B(net358),
    .C(_0110_),
    .A(\waggle_demo.p0[6] ),
    .Y(_0130_));
 sg13g2_a21o_1 _1757_ (.A2(_0110_),
    .A1(net358),
    .B1(\waggle_demo.p0[6] ),
    .X(_0131_));
 sg13g2_and2_1 _1758_ (.A(_0130_),
    .B(_0131_),
    .X(_0132_));
 sg13g2_nand2b_1 _1759_ (.Y(_0133_),
    .B(_0132_),
    .A_N(_0129_));
 sg13g2_xnor2_1 _1760_ (.Y(_0036_),
    .A(_0129_),
    .B(_0132_));
 sg13g2_and2_1 _1761_ (.A(_0130_),
    .B(_0133_),
    .X(_0134_));
 sg13g2_nand3_1 _1762_ (.B(net358),
    .C(_0115_),
    .A(\waggle_demo.p0[7] ),
    .Y(_0135_));
 sg13g2_a21o_1 _1763_ (.A2(_0115_),
    .A1(net358),
    .B1(\waggle_demo.p0[7] ),
    .X(_0136_));
 sg13g2_and2_1 _1764_ (.A(_0135_),
    .B(_0136_),
    .X(_0137_));
 sg13g2_nand2b_1 _1765_ (.Y(_0138_),
    .B(_0137_),
    .A_N(_0134_));
 sg13g2_xnor2_1 _1766_ (.Y(_0037_),
    .A(_0134_),
    .B(_0137_));
 sg13g2_and2_1 _1767_ (.A(_0135_),
    .B(_0138_),
    .X(_0139_));
 sg13g2_nand3_1 _1768_ (.B(net3),
    .C(net2),
    .A(net358),
    .Y(_0140_));
 sg13g2_nand4_1 _1769_ (.B(net358),
    .C(net3),
    .A(\waggle_demo.p0[8] ),
    .Y(_0141_),
    .D(net2));
 sg13g2_xor2_1 _1770_ (.B(_0140_),
    .A(\waggle_demo.p0[8] ),
    .X(_0142_));
 sg13g2_xor2_1 _1771_ (.B(_0142_),
    .A(_0139_),
    .X(_0038_));
 sg13g2_o21ai_1 _1772_ (.B1(_0141_),
    .Y(_0143_),
    .A1(_0139_),
    .A2(_0142_));
 sg13g2_xor2_1 _1773_ (.B(_0143_),
    .A(\waggle_demo.p0[9] ),
    .X(_0039_));
 sg13g2_xor2_1 _1774_ (.B(_0108_),
    .A(\waggle_demo.p0[1] ),
    .X(_0031_));
 sg13g2_nand2_1 _1775_ (.Y(_0144_),
    .A(\frame[1] ),
    .B(\frame[0] ));
 sg13g2_xor2_1 _1776_ (.B(\frame[0] ),
    .A(\frame[1] ),
    .X(_0025_));
 sg13g2_xnor2_1 _1777_ (.Y(_0026_),
    .A(\frame[2] ),
    .B(_0144_));
 sg13g2_nor2_1 _1778_ (.A(_0016_),
    .B(_0144_),
    .Y(_0145_));
 sg13g2_xor2_1 _1779_ (.B(_0145_),
    .A(\frame[3] ),
    .X(_0027_));
 sg13g2_nand4_1 _1780_ (.B(\frame[1] ),
    .C(\frame[0] ),
    .A(\frame[2] ),
    .Y(_0146_),
    .D(\frame[3] ));
 sg13g2_inv_1 _1781_ (.Y(_0147_),
    .A(_0146_));
 sg13g2_xnor2_1 _1782_ (.Y(_0028_),
    .A(\frame[4] ),
    .B(_0146_));
 sg13g2_nor2_1 _1783_ (.A(_0011_),
    .B(_0146_),
    .Y(_0148_));
 sg13g2_xor2_1 _1784_ (.B(_0148_),
    .A(\frame[5] ),
    .X(_0029_));
 sg13g2_nand3_1 _1785_ (.B(\frame[5] ),
    .C(_0147_),
    .A(\frame[4] ),
    .Y(_0149_));
 sg13g2_xnor2_1 _1786_ (.Y(_0030_),
    .A(\frame[6] ),
    .B(_0149_));
 sg13g2_xor2_1 _1787_ (.B(\waggle_demo.ypos[1] ),
    .A(\waggle_demo.ypos[2] ),
    .X(_0057_));
 sg13g2_nand3_1 _1788_ (.B(\waggle_demo.ypos[2] ),
    .C(\waggle_demo.ypos[1] ),
    .A(\waggle_demo.ypos[3] ),
    .Y(_0150_));
 sg13g2_a21o_1 _1789_ (.A2(\waggle_demo.ypos[1] ),
    .A1(\waggle_demo.ypos[2] ),
    .B1(\waggle_demo.ypos[3] ),
    .X(_0151_));
 sg13g2_and2_1 _1790_ (.A(_0150_),
    .B(_0151_),
    .X(_0058_));
 sg13g2_nor2_2 _1791_ (.A(_0259_),
    .B(_0150_),
    .Y(_0152_));
 sg13g2_xnor2_1 _1792_ (.Y(_0059_),
    .A(\waggle_demo.ypos[4] ),
    .B(_0150_));
 sg13g2_xor2_1 _1793_ (.B(_0152_),
    .A(\waggle_demo.ypos[5] ),
    .X(_0060_));
 sg13g2_nand3_1 _1794_ (.B(\waggle_demo.ypos[6] ),
    .C(_0152_),
    .A(\waggle_demo.ypos[5] ),
    .Y(_0153_));
 sg13g2_a21o_1 _1795_ (.A2(_0152_),
    .A1(\waggle_demo.ypos[5] ),
    .B1(\waggle_demo.ypos[6] ),
    .X(_0154_));
 sg13g2_and2_1 _1796_ (.A(_0153_),
    .B(_0154_),
    .X(_0061_));
 sg13g2_xnor2_1 _1797_ (.Y(_0062_),
    .A(\waggle_demo.ypos[7] ),
    .B(_0153_));
 sg13g2_xor2_1 _1798_ (.B(\waggle_demo.xpos[0] ),
    .A(\waggle_demo.xpos[1] ),
    .X(_0050_));
 sg13g2_nand3_1 _1799_ (.B(\waggle_demo.xpos[1] ),
    .C(\waggle_demo.xpos[0] ),
    .A(\waggle_demo.xpos[2] ),
    .Y(_0155_));
 sg13g2_a21o_1 _1800_ (.A2(\waggle_demo.xpos[0] ),
    .A1(\waggle_demo.xpos[1] ),
    .B1(\waggle_demo.xpos[2] ),
    .X(_0156_));
 sg13g2_and2_1 _1801_ (.A(_0155_),
    .B(_0156_),
    .X(_0051_));
 sg13g2_nor2_2 _1802_ (.A(_0254_),
    .B(_0155_),
    .Y(_0157_));
 sg13g2_xnor2_1 _1803_ (.Y(_0052_),
    .A(\waggle_demo.xpos[3] ),
    .B(_0155_));
 sg13g2_xor2_1 _1804_ (.B(_0157_),
    .A(\waggle_demo.xpos[4] ),
    .X(_0053_));
 sg13g2_nand3_1 _1805_ (.B(\waggle_demo.xpos[4] ),
    .C(_0157_),
    .A(\waggle_demo.xpos[5] ),
    .Y(_0158_));
 sg13g2_a21o_1 _1806_ (.A2(_0157_),
    .A1(\waggle_demo.xpos[4] ),
    .B1(\waggle_demo.xpos[5] ),
    .X(_0159_));
 sg13g2_and2_1 _1807_ (.A(_0158_),
    .B(_0159_),
    .X(_0054_));
 sg13g2_nand4_1 _1808_ (.B(\waggle_demo.xpos[4] ),
    .C(\waggle_demo.xpos[6] ),
    .A(\waggle_demo.xpos[5] ),
    .Y(_0160_),
    .D(_0157_));
 sg13g2_xnor2_1 _1809_ (.Y(_0055_),
    .A(\waggle_demo.xpos[6] ),
    .B(_0158_));
 sg13g2_xnor2_1 _1810_ (.Y(_0056_),
    .A(\waggle_demo.xpos[7] ),
    .B(_0160_));
 sg13g2_nor2_1 _1811_ (.A(net356),
    .B(net357),
    .Y(_0161_));
 sg13g2_nor3_2 _1812_ (.A(net356),
    .B(net4),
    .C(net357),
    .Y(_0162_));
 sg13g2_xor2_1 _1813_ (.B(_0162_),
    .A(\waggle_demo.p1[0] ),
    .X(_0040_));
 sg13g2_nor2b_1 _1814_ (.A(_0023_),
    .B_N(_0162_),
    .Y(_0163_));
 sg13g2_nor2b_1 _1815_ (.A(_0163_),
    .B_N(_0161_),
    .Y(_0164_));
 sg13g2_xnor2_1 _1816_ (.Y(_0041_),
    .A(_0257_),
    .B(_0164_));
 sg13g2_a22oi_1 _1817_ (.Y(_0165_),
    .B1(_0163_),
    .B2(_0257_),
    .A2(_0161_),
    .A1(_0258_));
 sg13g2_and2_1 _1818_ (.A(net4),
    .B(net357),
    .X(_0166_));
 sg13g2_nor2_1 _1819_ (.A(net356),
    .B(_0166_),
    .Y(_0167_));
 sg13g2_o21ai_1 _1820_ (.B1(_0167_),
    .Y(_0168_),
    .A1(net4),
    .A2(net357));
 sg13g2_xor2_1 _1821_ (.B(_0168_),
    .A(_0020_),
    .X(_0169_));
 sg13g2_nand2b_1 _1822_ (.Y(_0170_),
    .B(_0169_),
    .A_N(_0165_));
 sg13g2_xnor2_1 _1823_ (.Y(_0042_),
    .A(_0165_),
    .B(_0169_));
 sg13g2_o21ai_1 _1824_ (.B1(_0170_),
    .Y(_0171_),
    .A1(_0256_),
    .A2(_0168_));
 sg13g2_nor2b_1 _1825_ (.A(net356),
    .B_N(net357),
    .Y(_0172_));
 sg13g2_nor2b_1 _1826_ (.A(_0014_),
    .B_N(_0172_),
    .Y(_0173_));
 sg13g2_xnor2_1 _1827_ (.Y(_0174_),
    .A(_0014_),
    .B(_0172_));
 sg13g2_and2_1 _1828_ (.A(_0171_),
    .B(_0174_),
    .X(_0175_));
 sg13g2_xor2_1 _1829_ (.B(_0174_),
    .A(_0171_),
    .X(_0043_));
 sg13g2_o21ai_1 _1830_ (.B1(net356),
    .Y(_0176_),
    .A1(net4),
    .A2(net357));
 sg13g2_o21ai_1 _1831_ (.B1(_0176_),
    .Y(_0177_),
    .A1(net356),
    .A2(_0166_));
 sg13g2_xnor2_1 _1832_ (.Y(_0178_),
    .A(\waggle_demo.p1[4] ),
    .B(_0177_));
 sg13g2_o21ai_1 _1833_ (.B1(_0178_),
    .Y(_0179_),
    .A1(_0173_),
    .A2(_0175_));
 sg13g2_or3_1 _1834_ (.A(_0173_),
    .B(_0175_),
    .C(_0178_),
    .X(_0180_));
 sg13g2_and2_1 _1835_ (.A(_0179_),
    .B(_0180_),
    .X(_0044_));
 sg13g2_o21ai_1 _1836_ (.B1(_0179_),
    .Y(_0181_),
    .A1(_0018_),
    .A2(_0177_));
 sg13g2_nor2b_1 _1837_ (.A(net357),
    .B_N(net356),
    .Y(_0182_));
 sg13g2_nor2b_1 _1838_ (.A(_0015_),
    .B_N(_0182_),
    .Y(_0183_));
 sg13g2_xnor2_1 _1839_ (.Y(_0184_),
    .A(_0015_),
    .B(_0182_));
 sg13g2_and2_1 _1840_ (.A(_0181_),
    .B(_0184_),
    .X(_0185_));
 sg13g2_xor2_1 _1841_ (.B(_0184_),
    .A(_0181_),
    .X(_0045_));
 sg13g2_nor2_1 _1842_ (.A(_0166_),
    .B(_0176_),
    .Y(_0186_));
 sg13g2_xnor2_1 _1843_ (.Y(_0187_),
    .A(_0017_),
    .B(_0186_));
 sg13g2_o21ai_1 _1844_ (.B1(_0187_),
    .Y(_0188_),
    .A1(_0183_),
    .A2(_0185_));
 sg13g2_or3_1 _1845_ (.A(_0183_),
    .B(_0185_),
    .C(_0187_),
    .X(_0189_));
 sg13g2_and2_1 _1846_ (.A(_0188_),
    .B(_0189_),
    .X(_0046_));
 sg13g2_nand2_1 _1847_ (.Y(_0190_),
    .A(\waggle_demo.p1[6] ),
    .B(_0186_));
 sg13g2_nand2_1 _1848_ (.Y(_0191_),
    .A(_0188_),
    .B(_0190_));
 sg13g2_inv_1 _1849_ (.Y(_0192_),
    .A(_0191_));
 sg13g2_nand3_1 _1850_ (.B(net6),
    .C(net5),
    .A(\waggle_demo.p1[7] ),
    .Y(_0193_));
 sg13g2_a21o_1 _1851_ (.A2(net357),
    .A1(net6),
    .B1(\waggle_demo.p1[7] ),
    .X(_0194_));
 sg13g2_nand2_1 _1852_ (.Y(_0195_),
    .A(_0193_),
    .B(_0194_));
 sg13g2_xnor2_1 _1853_ (.Y(_0047_),
    .A(_0191_),
    .B(_0195_));
 sg13g2_o21ai_1 _1854_ (.B1(_0193_),
    .Y(_0196_),
    .A1(_0192_),
    .A2(_0195_));
 sg13g2_and2_1 _1855_ (.A(net356),
    .B(_0166_),
    .X(_0197_));
 sg13g2_xnor2_1 _1856_ (.Y(_0198_),
    .A(_0022_),
    .B(_0197_));
 sg13g2_xor2_1 _1857_ (.B(_0198_),
    .A(_0196_),
    .X(_0048_));
 sg13g2_a22oi_1 _1858_ (.Y(_0199_),
    .B1(_0198_),
    .B2(_0196_),
    .A2(_0197_),
    .A1(\waggle_demo.p1[8] ));
 sg13g2_xor2_1 _1859_ (.B(_0199_),
    .A(_0021_),
    .X(_0049_));
 sg13g2_nor3_1 _1860_ (.A(net347),
    .B(net349),
    .C(\hvsync_gen.vpos[8] ),
    .Y(_0200_));
 sg13g2_nand2_1 _1861_ (.Y(_0201_),
    .A(\hvsync_gen.vpos[9] ),
    .B(_0200_));
 sg13g2_nor4_1 _1862_ (.A(net353),
    .B(net354),
    .C(net345),
    .D(net346),
    .Y(_0202_));
 sg13g2_nand3_1 _1863_ (.B(net352),
    .C(_0202_),
    .A(net350),
    .Y(_0203_));
 sg13g2_o21ai_1 _1864_ (.B1(net368),
    .Y(_0204_),
    .A1(_0201_),
    .A2(_0203_));
 sg13g2_and3_1 _1865_ (.X(_0205_),
    .A(net85),
    .B(\hpos[0] ),
    .C(net67));
 sg13g2_and2_1 _1866_ (.A(net79),
    .B(_0205_),
    .X(_0206_));
 sg13g2_and2_1 _1867_ (.A(\hpos[4] ),
    .B(_0206_),
    .X(_0207_));
 sg13g2_nor3_1 _1868_ (.A(\hpos[7] ),
    .B(\hpos[6] ),
    .C(\hpos[5] ),
    .Y(_0208_));
 sg13g2_and4_2 _1869_ (.A(\hpos[9] ),
    .B(net61),
    .C(_0207_),
    .D(_0208_),
    .X(_0209_));
 sg13g2_nor2b_2 _1870_ (.A(_0204_),
    .B_N(_0209_),
    .Y(_0210_));
 sg13g2_nor2_2 _1871_ (.A(_0253_),
    .B(_0209_),
    .Y(_0211_));
 sg13g2_nand2b_1 _1872_ (.Y(_0212_),
    .B(net368),
    .A_N(_0209_));
 sg13g2_a22oi_1 _1873_ (.Y(_0213_),
    .B1(_0211_),
    .B2(net354),
    .A2(_0210_),
    .A1(net58));
 sg13g2_inv_1 _1874_ (.Y(_0067_),
    .A(net59));
 sg13g2_and3_1 _1875_ (.X(_0214_),
    .A(net353),
    .B(net355),
    .C(net334));
 sg13g2_a21oi_1 _1876_ (.A1(net355),
    .A2(_0209_),
    .Y(_0215_),
    .B1(net353));
 sg13g2_nor3_1 _1877_ (.A(_0253_),
    .B(_0214_),
    .C(net81),
    .Y(_0068_));
 sg13g2_and3_1 _1878_ (.X(_0216_),
    .A(net353),
    .B(net354),
    .C(net352));
 sg13g2_o21ai_1 _1879_ (.B1(_0212_),
    .Y(_0217_),
    .A1(_0204_),
    .A2(_0216_));
 sg13g2_o21ai_1 _1880_ (.B1(_0217_),
    .Y(_0218_),
    .A1(net63),
    .A2(_0214_));
 sg13g2_inv_1 _1881_ (.Y(_0069_),
    .A(_0218_));
 sg13g2_nand2_1 _1882_ (.Y(_0219_),
    .A(net350),
    .B(_0217_));
 sg13g2_nand2_1 _1883_ (.Y(_0220_),
    .A(_0210_),
    .B(_0216_));
 sg13g2_o21ai_1 _1884_ (.B1(_0219_),
    .Y(_0070_),
    .A1(net350),
    .A2(_0220_));
 sg13g2_and3_1 _1885_ (.X(_0221_),
    .A(net350),
    .B(net349),
    .C(_0216_));
 sg13g2_nor2_1 _1886_ (.A(_0204_),
    .B(_0221_),
    .Y(_0222_));
 sg13g2_nor2_1 _1887_ (.A(_0211_),
    .B(_0222_),
    .Y(_0223_));
 sg13g2_nand3_1 _1888_ (.B(net334),
    .C(_0216_),
    .A(net350),
    .Y(_0224_));
 sg13g2_a21oi_1 _1889_ (.A1(_0251_),
    .A2(_0224_),
    .Y(_0071_),
    .B1(_0223_));
 sg13g2_nand2_1 _1890_ (.Y(_0225_),
    .A(_0210_),
    .B(_0221_));
 sg13g2_o21ai_1 _1891_ (.B1(net347),
    .Y(_0226_),
    .A1(_0211_),
    .A2(_0222_));
 sg13g2_o21ai_1 _1892_ (.B1(_0226_),
    .Y(_0072_),
    .A1(net348),
    .A2(_0225_));
 sg13g2_nand3_1 _1893_ (.B(net347),
    .C(_0221_),
    .A(net346),
    .Y(_0227_));
 sg13g2_inv_1 _1894_ (.Y(_0228_),
    .A(_0227_));
 sg13g2_o21ai_1 _1895_ (.B1(net334),
    .Y(_0229_),
    .A1(_0204_),
    .A2(_0228_));
 sg13g2_and3_1 _1896_ (.X(_0230_),
    .A(net347),
    .B(net334),
    .C(_0221_));
 sg13g2_o21ai_1 _1897_ (.B1(_0229_),
    .Y(_0231_),
    .A1(net64),
    .A2(_0230_));
 sg13g2_inv_1 _1898_ (.Y(_0073_),
    .A(_0231_));
 sg13g2_nor2_1 _1899_ (.A(net60),
    .B(_0227_),
    .Y(_0232_));
 sg13g2_a22oi_1 _1900_ (.Y(_0233_),
    .B1(_0232_),
    .B2(_0210_),
    .A2(_0229_),
    .A1(net60));
 sg13g2_inv_1 _1901_ (.Y(_0074_),
    .A(_0233_));
 sg13g2_nand2b_1 _1902_ (.Y(_0234_),
    .B(_0267_),
    .A_N(_0204_));
 sg13g2_nand2_1 _1903_ (.Y(_0235_),
    .A(_0223_),
    .B(_0234_));
 sg13g2_nand3_1 _1904_ (.B(net346),
    .C(_0230_),
    .A(net345),
    .Y(_0236_));
 sg13g2_a22oi_1 _1905_ (.Y(_0075_),
    .B1(_0236_),
    .B2(_0252_),
    .A2(_0234_),
    .A1(_0223_));
 sg13g2_nand2_1 _1906_ (.Y(_0237_),
    .A(net69),
    .B(_0235_));
 sg13g2_or2_1 _1907_ (.X(_0238_),
    .B(_0236_),
    .A(_0204_));
 sg13g2_o21ai_1 _1908_ (.B1(_0237_),
    .Y(_0076_),
    .A1(_0262_),
    .A2(_0238_));
 sg13g2_and2_1 _1909_ (.A(net57),
    .B(_0211_),
    .X(_0077_));
 sg13g2_o21ai_1 _1910_ (.B1(_0211_),
    .Y(_0239_),
    .A1(net75),
    .A2(\hpos[0] ));
 sg13g2_a21oi_1 _1911_ (.A1(net75),
    .A2(\hpos[0] ),
    .Y(_0078_),
    .B1(_0239_));
 sg13g2_a21oi_1 _1912_ (.A1(\hpos[1] ),
    .A2(\hpos[0] ),
    .Y(_0240_),
    .B1(net67));
 sg13g2_nor3_1 _1913_ (.A(_0253_),
    .B(_0205_),
    .C(net68),
    .Y(_0079_));
 sg13g2_o21ai_1 _1914_ (.B1(net364),
    .Y(_0241_),
    .A1(net79),
    .A2(_0205_));
 sg13g2_nor2_1 _1915_ (.A(_0206_),
    .B(_0241_),
    .Y(_0080_));
 sg13g2_o21ai_1 _1916_ (.B1(net364),
    .Y(_0242_),
    .A1(net84),
    .A2(_0206_));
 sg13g2_nor2_1 _1917_ (.A(_0207_),
    .B(_0242_),
    .Y(_0081_));
 sg13g2_o21ai_1 _1918_ (.B1(_0211_),
    .Y(_0243_),
    .A1(net338),
    .A2(_0207_));
 sg13g2_a21oi_1 _1919_ (.A1(net338),
    .A2(_0207_),
    .Y(_0082_),
    .B1(_0243_));
 sg13g2_a21oi_1 _1920_ (.A1(net338),
    .A2(_0207_),
    .Y(_0244_),
    .B1(net71));
 sg13g2_and2_1 _1921_ (.A(_0264_),
    .B(_0206_),
    .X(_0245_));
 sg13g2_nor3_1 _1922_ (.A(net334),
    .B(net72),
    .C(_0245_),
    .Y(_0083_));
 sg13g2_xnor2_1 _1923_ (.Y(_0246_),
    .A(net65),
    .B(_0245_));
 sg13g2_nor2_1 _1924_ (.A(net334),
    .B(_0246_),
    .Y(_0084_));
 sg13g2_a21oi_1 _1925_ (.A1(net65),
    .A2(_0245_),
    .Y(_0247_),
    .B1(net61));
 sg13g2_and3_1 _1926_ (.X(_0248_),
    .A(net61),
    .B(\hpos[7] ),
    .C(_0245_));
 sg13g2_nor3_1 _1927_ (.A(net334),
    .B(_0247_),
    .C(_0248_),
    .Y(_0085_));
 sg13g2_a21oi_1 _1928_ (.A1(net77),
    .A2(_0248_),
    .Y(_0249_),
    .B1(net334));
 sg13g2_o21ai_1 _1929_ (.B1(_0249_),
    .Y(_0250_),
    .A1(net77),
    .A2(_0248_));
 sg13g2_inv_1 _1930_ (.Y(_0086_),
    .A(_0250_));
 sg13g2_inv_1 _1931_ (.Y(_0251_),
    .A(net349));
 sg13g2_inv_1 _1932_ (.Y(_0252_),
    .A(net73));
 sg13g2_inv_1 _1933_ (.Y(_0253_),
    .A(net368));
 sg13g2_inv_1 _1934_ (.Y(_0254_),
    .A(\waggle_demo.xpos[3] ));
 sg13g2_inv_1 _1935_ (.Y(_0255_),
    .A(\waggle_demo.xpos[2] ));
 sg13g2_inv_1 _1936_ (.Y(_0256_),
    .A(\waggle_demo.p1[2] ));
 sg13g2_inv_1 _1937_ (.Y(_0257_),
    .A(\waggle_demo.p1[1] ));
 sg13g2_inv_1 _1938_ (.Y(_0258_),
    .A(_0019_));
 sg13g2_inv_1 _1939_ (.Y(_0259_),
    .A(\waggle_demo.ypos[4] ));
 sg13g2_inv_1 _1940_ (.Y(_0260_),
    .A(\waggle_demo.xpos[6] ));
 sg13g2_nand3_1 _1941_ (.B(net346),
    .C(net347),
    .A(net345),
    .Y(_0261_));
 sg13g2_nand2b_1 _1942_ (.Y(_0262_),
    .B(net73),
    .A_N(net69));
 sg13g2_nand3b_1 _1943_ (.B(net350),
    .C(net353),
    .Y(_0263_),
    .A_N(net352));
 sg13g2_nor4_1 _1944_ (.A(net349),
    .B(_0261_),
    .C(_0262_),
    .D(_0263_),
    .Y(_0001_));
 sg13g2_and3_1 _1945_ (.X(_0264_),
    .A(\hpos[6] ),
    .B(net338),
    .C(\hpos[4] ));
 sg13g2_nand2_1 _1946_ (.Y(_0265_),
    .A(\hpos[9] ),
    .B(\hpos[7] ));
 sg13g2_nor3_1 _1947_ (.A(\hpos[6] ),
    .B(net338),
    .C(\hpos[4] ),
    .Y(_0266_));
 sg13g2_nor4_1 _1948_ (.A(net61),
    .B(_0264_),
    .C(_0265_),
    .D(_0266_),
    .Y(_0000_));
 sg13g2_or2_1 _1949_ (.X(_0267_),
    .B(_0261_),
    .A(_0252_));
 sg13g2_o21ai_1 _1950_ (.B1(\hpos[9] ),
    .Y(_0268_),
    .A1(\hpos[8] ),
    .A2(\hpos[7] ));
 sg13g2_nand2_1 _1951_ (.Y(_0269_),
    .A(_0267_),
    .B(_0268_));
 sg13g2_nor2_2 _1952_ (.A(\hvsync_gen.vpos[9] ),
    .B(_0269_),
    .Y(_0270_));
 sg13g2_and2_1 _1953_ (.A(\palette_inst.palette[4] ),
    .B(_0270_),
    .X(uo_out[4]));
 sg13g2_and2_1 _1954_ (.A(\palette_inst.palette[5] ),
    .B(_0270_),
    .X(uo_out[0]));
 sg13g2_and2_1 _1955_ (.A(\palette_inst.palette[2] ),
    .B(_0270_),
    .X(uo_out[5]));
 sg13g2_and2_1 _1956_ (.A(\palette_inst.palette[3] ),
    .B(_0270_),
    .X(uo_out[1]));
 sg13g2_and2_1 _1957_ (.A(\palette_inst.palette[0] ),
    .B(_0270_),
    .X(uo_out[6]));
 sg13g2_and2_1 _1958_ (.A(\palette_inst.palette[1] ),
    .B(_0270_),
    .X(uo_out[2]));
 sg13g2_nor2b_1 _1959_ (.A(\waggle_demo.ypos[5] ),
    .B_N(net348),
    .Y(_0271_));
 sg13g2_nand2b_1 _1960_ (.Y(_0272_),
    .B(\waggle_demo.ypos[5] ),
    .A_N(net348));
 sg13g2_nand2b_1 _1961_ (.Y(_0273_),
    .B(_0272_),
    .A_N(_0271_));
 sg13g2_mux2_1 _1962_ (.A0(net351),
    .A1(\hpos[3] ),
    .S(net360),
    .X(_0274_));
 sg13g2_nand2_1 _1963_ (.Y(_0275_),
    .A(\waggle_demo.p1[3] ),
    .B(_0274_));
 sg13g2_mux2_1 _1964_ (.A0(net352),
    .A1(\hpos[2] ),
    .S(net360),
    .X(_0276_));
 sg13g2_mux2_1 _1965_ (.A0(net353),
    .A1(\hpos[1] ),
    .S(net360),
    .X(_0277_));
 sg13g2_nand2_1 _1966_ (.Y(_0278_),
    .A(_0258_),
    .B(_0277_));
 sg13g2_mux2_1 _1967_ (.A0(net355),
    .A1(\hpos[0] ),
    .S(net360),
    .X(_0279_));
 sg13g2_nand2_1 _1968_ (.Y(_0280_),
    .A(\waggle_demo.p1[0] ),
    .B(_0279_));
 sg13g2_xnor2_1 _1969_ (.Y(_0281_),
    .A(\waggle_demo.p1[1] ),
    .B(_0277_));
 sg13g2_o21ai_1 _1970_ (.B1(_0278_),
    .Y(_0282_),
    .A1(_0280_),
    .A2(_0281_));
 sg13g2_xnor2_1 _1971_ (.Y(_0283_),
    .A(_0020_),
    .B(_0276_));
 sg13g2_a22oi_1 _1972_ (.Y(_0284_),
    .B1(_0282_),
    .B2(_0283_),
    .A2(_0276_),
    .A1(\waggle_demo.p1[2] ));
 sg13g2_xnor2_1 _1973_ (.Y(_0285_),
    .A(\waggle_demo.p1[3] ),
    .B(_0274_));
 sg13g2_o21ai_1 _1974_ (.B1(_0275_),
    .Y(_0286_),
    .A1(_0284_),
    .A2(_0285_));
 sg13g2_mux2_2 _1975_ (.A0(net348),
    .A1(net338),
    .S(net360),
    .X(_0287_));
 sg13g2_nor2_1 _1976_ (.A(\waggle_demo.p1[5] ),
    .B(_0287_),
    .Y(_0288_));
 sg13g2_xnor2_1 _1977_ (.Y(_0289_),
    .A(\waggle_demo.p1[5] ),
    .B(_0287_));
 sg13g2_nand2_1 _1978_ (.Y(_0290_),
    .A(\hpos[4] ),
    .B(net361));
 sg13g2_o21ai_1 _1979_ (.B1(_0290_),
    .Y(_0291_),
    .A1(_0251_),
    .A2(net360));
 sg13g2_xnor2_1 _1980_ (.Y(_0292_),
    .A(_0018_),
    .B(_0291_));
 sg13g2_nor2b_1 _1981_ (.A(_0289_),
    .B_N(_0292_),
    .Y(_0293_));
 sg13g2_mux2_1 _1982_ (.A0(net345),
    .A1(\hpos[7] ),
    .S(net361),
    .X(_0294_));
 sg13g2_nand2_1 _1983_ (.Y(_0295_),
    .A(\waggle_demo.p1[7] ),
    .B(_0294_));
 sg13g2_or2_1 _1984_ (.X(_0296_),
    .B(_0294_),
    .A(\waggle_demo.p1[7] ));
 sg13g2_mux2_1 _1985_ (.A0(net346),
    .A1(\hpos[6] ),
    .S(net361),
    .X(_0297_));
 sg13g2_nand2_1 _1986_ (.Y(_0298_),
    .A(\waggle_demo.p1[6] ),
    .B(_0297_));
 sg13g2_nand2_1 _1987_ (.Y(_0299_),
    .A(_0295_),
    .B(_0298_));
 sg13g2_nand2_1 _1988_ (.Y(_0300_),
    .A(_0296_),
    .B(_0299_));
 sg13g2_a22oi_1 _1989_ (.Y(_0301_),
    .B1(_0291_),
    .B2(\waggle_demo.p1[4] ),
    .A2(_0287_),
    .A1(\waggle_demo.p1[5] ));
 sg13g2_nor2_1 _1990_ (.A(_0288_),
    .B(_0301_),
    .Y(_0302_));
 sg13g2_nand2b_1 _1991_ (.Y(_0303_),
    .B(_0300_),
    .A_N(_0302_));
 sg13g2_a21oi_1 _1992_ (.A1(_0286_),
    .A2(_0293_),
    .Y(_0304_),
    .B1(_0303_));
 sg13g2_a21o_1 _1993_ (.A2(_0293_),
    .A1(_0286_),
    .B1(_0303_),
    .X(_0305_));
 sg13g2_xnor2_1 _1994_ (.Y(_0306_),
    .A(_0017_),
    .B(_0297_));
 sg13g2_inv_1 _1995_ (.Y(_0307_),
    .A(_0306_));
 sg13g2_nand2_1 _1996_ (.Y(_0308_),
    .A(_0296_),
    .B(_0306_));
 sg13g2_o21ai_1 _1997_ (.B1(_0296_),
    .Y(_0309_),
    .A1(_0299_),
    .A2(_0306_));
 sg13g2_nand2_1 _1998_ (.Y(_0310_),
    .A(_0300_),
    .B(_0308_));
 sg13g2_nand2_1 _1999_ (.Y(_0311_),
    .A(\hpos[8] ),
    .B(net361));
 sg13g2_o21ai_1 _2000_ (.B1(_0311_),
    .Y(_0312_),
    .A1(_0252_),
    .A2(net360));
 sg13g2_inv_1 _2001_ (.Y(_0313_),
    .A(_0312_));
 sg13g2_xnor2_1 _2002_ (.Y(_0314_),
    .A(\waggle_demo.p1[8] ),
    .B(_0312_));
 sg13g2_xor2_1 _2003_ (.B(_0312_),
    .A(\waggle_demo.p1[8] ),
    .X(_0315_));
 sg13g2_nor3_2 _2004_ (.A(_0304_),
    .B(_0309_),
    .C(_0314_),
    .Y(_0316_));
 sg13g2_nand3_1 _2005_ (.B(_0310_),
    .C(_0315_),
    .A(_0305_),
    .Y(_0317_));
 sg13g2_a21oi_2 _2006_ (.B1(_0315_),
    .Y(_0318_),
    .A2(_0310_),
    .A1(_0305_));
 sg13g2_o21ai_1 _2007_ (.B1(_0314_),
    .Y(_0319_),
    .A1(_0304_),
    .A2(_0309_));
 sg13g2_nand2_2 _2008_ (.Y(_0320_),
    .A(_0317_),
    .B(_0319_));
 sg13g2_nand2_1 _2009_ (.Y(_0321_),
    .A(_0295_),
    .B(_0296_));
 sg13g2_a21oi_1 _2010_ (.A1(_0286_),
    .A2(_0293_),
    .Y(_0322_),
    .B1(_0302_));
 sg13g2_o21ai_1 _2011_ (.B1(_0298_),
    .Y(_0323_),
    .A1(_0307_),
    .A2(_0322_));
 sg13g2_xor2_1 _2012_ (.B(_0323_),
    .A(_0321_),
    .X(_0324_));
 sg13g2_xor2_1 _2013_ (.B(_0324_),
    .A(_0320_),
    .X(_0325_));
 sg13g2_xnor2_1 _2014_ (.Y(_0326_),
    .A(_0320_),
    .B(_0324_));
 sg13g2_xnor2_1 _2015_ (.Y(_0327_),
    .A(_0306_),
    .B(_0322_));
 sg13g2_xnor2_1 _2016_ (.Y(_0328_),
    .A(_0320_),
    .B(_0327_));
 sg13g2_xor2_1 _2017_ (.B(_0327_),
    .A(_0320_),
    .X(_0329_));
 sg13g2_a22oi_1 _2018_ (.Y(_0330_),
    .B1(_0292_),
    .B2(_0286_),
    .A2(_0291_),
    .A1(\waggle_demo.p1[4] ));
 sg13g2_xnor2_1 _2019_ (.Y(_0331_),
    .A(_0289_),
    .B(_0330_));
 sg13g2_o21ai_1 _2020_ (.B1(_0331_),
    .Y(_0332_),
    .A1(_0316_),
    .A2(_0318_));
 sg13g2_nand3b_1 _2021_ (.B(net309),
    .C(_0317_),
    .Y(_0333_),
    .A_N(_0331_));
 sg13g2_nand2_1 _2022_ (.Y(_0334_),
    .A(_0332_),
    .B(_0333_));
 sg13g2_and2_1 _2023_ (.A(_0332_),
    .B(_0333_),
    .X(_0335_));
 sg13g2_xor2_1 _2024_ (.B(_0292_),
    .A(_0286_),
    .X(_0336_));
 sg13g2_nand3_1 _2025_ (.B(net309),
    .C(_0336_),
    .A(net310),
    .Y(_0337_));
 sg13g2_a21o_1 _2026_ (.A2(net309),
    .A1(net310),
    .B1(_0336_),
    .X(_0338_));
 sg13g2_nand2_1 _2027_ (.Y(_0339_),
    .A(_0337_),
    .B(_0338_));
 sg13g2_and2_1 _2028_ (.A(_0337_),
    .B(_0338_),
    .X(_0340_));
 sg13g2_nor2_2 _2029_ (.A(net302),
    .B(net296),
    .Y(_0341_));
 sg13g2_xor2_1 _2030_ (.B(_0285_),
    .A(_0284_),
    .X(_0342_));
 sg13g2_nand3_1 _2031_ (.B(net309),
    .C(_0342_),
    .A(net310),
    .Y(_0343_));
 sg13g2_a21o_1 _2032_ (.A2(net309),
    .A1(net310),
    .B1(_0342_),
    .X(_0344_));
 sg13g2_nand2_1 _2033_ (.Y(_0345_),
    .A(_0343_),
    .B(_0344_));
 sg13g2_and2_1 _2034_ (.A(_0343_),
    .B(_0344_),
    .X(_0346_));
 sg13g2_a21oi_2 _2035_ (.B1(_0335_),
    .Y(_0347_),
    .A2(net291),
    .A1(net297));
 sg13g2_nand2_1 _2036_ (.Y(_0348_),
    .A(net305),
    .B(_0347_));
 sg13g2_nand2_2 _2037_ (.Y(_0349_),
    .A(net308),
    .B(_0348_));
 sg13g2_xor2_1 _2038_ (.B(_0283_),
    .A(_0282_),
    .X(_0350_));
 sg13g2_xnor2_1 _2039_ (.Y(_0351_),
    .A(_0282_),
    .B(_0283_));
 sg13g2_nand3_1 _2040_ (.B(net309),
    .C(_0350_),
    .A(net310),
    .Y(_0352_));
 sg13g2_o21ai_1 _2041_ (.B1(_0351_),
    .Y(_0353_),
    .A1(_0316_),
    .A2(_0318_));
 sg13g2_nand2_2 _2042_ (.Y(_0354_),
    .A(_0352_),
    .B(_0353_));
 sg13g2_and2_2 _2043_ (.A(_0352_),
    .B(_0353_),
    .X(_0355_));
 sg13g2_nand2_1 _2044_ (.Y(_0356_),
    .A(net298),
    .B(net288));
 sg13g2_nor2_2 _2045_ (.A(net290),
    .B(_0355_),
    .Y(_0357_));
 sg13g2_inv_1 _2046_ (.Y(_0358_),
    .A(_0357_));
 sg13g2_and2_1 _2047_ (.A(_0341_),
    .B(_0357_),
    .X(_0359_));
 sg13g2_nor2_1 _2048_ (.A(net305),
    .B(_0359_),
    .Y(_0360_));
 sg13g2_o21ai_1 _2049_ (.B1(_0349_),
    .Y(_0361_),
    .A1(net308),
    .A2(_0360_));
 sg13g2_o21ai_1 _2050_ (.B1(net310),
    .Y(_0362_),
    .A1(_0022_),
    .A2(_0313_));
 sg13g2_mux2_2 _2051_ (.A0(\hvsync_gen.vpos[9] ),
    .A1(\hpos[9] ),
    .S(net360),
    .X(_0363_));
 sg13g2_xnor2_1 _2052_ (.Y(_0364_),
    .A(_0021_),
    .B(_0363_));
 sg13g2_xnor2_1 _2053_ (.Y(_0365_),
    .A(_0362_),
    .B(_0364_));
 sg13g2_xor2_1 _2054_ (.B(_0364_),
    .A(_0362_),
    .X(_0366_));
 sg13g2_nand2_1 _2055_ (.Y(_0367_),
    .A(net301),
    .B(net295));
 sg13g2_xor2_1 _2056_ (.B(_0279_),
    .A(_0023_),
    .X(_0368_));
 sg13g2_o21ai_1 _2057_ (.B1(_0368_),
    .Y(_0369_),
    .A1(_0316_),
    .A2(_0318_));
 sg13g2_or3_2 _2058_ (.A(_0316_),
    .B(_0318_),
    .C(_0368_),
    .X(_0370_));
 sg13g2_nand2_1 _2059_ (.Y(_0371_),
    .A(_0369_),
    .B(_0370_));
 sg13g2_and2_1 _2060_ (.A(_0369_),
    .B(_0370_),
    .X(_0372_));
 sg13g2_xor2_1 _2061_ (.B(_0281_),
    .A(_0280_),
    .X(_0373_));
 sg13g2_nand3_1 _2062_ (.B(net309),
    .C(_0373_),
    .A(net310),
    .Y(_0374_));
 sg13g2_a21o_2 _2063_ (.A2(net309),
    .A1(net310),
    .B1(_0373_),
    .X(_0375_));
 sg13g2_nand2_2 _2064_ (.Y(_0376_),
    .A(_0374_),
    .B(_0375_));
 sg13g2_and2_2 _2065_ (.A(_0374_),
    .B(_0375_),
    .X(_0377_));
 sg13g2_nand2_1 _2066_ (.Y(_0378_),
    .A(_0354_),
    .B(net283));
 sg13g2_a22oi_1 _2067_ (.Y(_0379_),
    .B1(_0374_),
    .B2(_0375_),
    .A2(_0370_),
    .A1(_0369_));
 sg13g2_nand2_1 _2068_ (.Y(_0380_),
    .A(net286),
    .B(_0376_));
 sg13g2_nand2_1 _2069_ (.Y(_0381_),
    .A(net287),
    .B(net281));
 sg13g2_a21oi_1 _2070_ (.A1(net287),
    .A2(net281),
    .Y(_0382_),
    .B1(net293));
 sg13g2_nor2_1 _2071_ (.A(net296),
    .B(_0382_),
    .Y(_0383_));
 sg13g2_nor2_1 _2072_ (.A(net303),
    .B(_0383_),
    .Y(_0384_));
 sg13g2_and4_2 _2073_ (.A(_0369_),
    .B(_0370_),
    .C(_0374_),
    .D(_0375_),
    .X(_0385_));
 sg13g2_nand4_1 _2074_ (.B(_0370_),
    .C(_0374_),
    .A(_0369_),
    .Y(_0386_),
    .D(_0375_));
 sg13g2_nor2_1 _2075_ (.A(net293),
    .B(net288),
    .Y(_0387_));
 sg13g2_nand4_1 _2076_ (.B(_0344_),
    .C(_0352_),
    .A(_0343_),
    .Y(_0388_),
    .D(_0353_));
 sg13g2_and4_2 _2077_ (.A(_0352_),
    .B(_0353_),
    .C(_0374_),
    .D(_0375_),
    .X(_0389_));
 sg13g2_nand4_1 _2078_ (.B(_0353_),
    .C(_0374_),
    .A(_0352_),
    .Y(_0390_),
    .D(_0375_));
 sg13g2_nand2_1 _2079_ (.Y(_0391_),
    .A(net284),
    .B(_0389_));
 sg13g2_or2_1 _2080_ (.X(_0392_),
    .B(net280),
    .A(_0386_));
 sg13g2_o21ai_1 _2081_ (.B1(_0384_),
    .Y(_0393_),
    .A1(net299),
    .A2(_0392_));
 sg13g2_a21oi_1 _2082_ (.A1(net299),
    .A2(_0357_),
    .Y(_0394_),
    .B1(net301));
 sg13g2_nor2_2 _2083_ (.A(net289),
    .B(_0389_),
    .Y(_0395_));
 sg13g2_nand2_1 _2084_ (.Y(_0396_),
    .A(net293),
    .B(_0390_));
 sg13g2_o21ai_1 _2085_ (.B1(_0394_),
    .Y(_0397_),
    .A1(net299),
    .A2(_0395_));
 sg13g2_nand3_1 _2086_ (.B(_0357_),
    .C(_0376_),
    .A(_0339_),
    .Y(_0398_));
 sg13g2_nor2_1 _2087_ (.A(net284),
    .B(_0398_),
    .Y(_0399_));
 sg13g2_a21oi_1 _2088_ (.A1(_0357_),
    .A2(net283),
    .Y(_0400_),
    .B1(net299));
 sg13g2_o21ai_1 _2089_ (.B1(net301),
    .Y(_0401_),
    .A1(_0399_),
    .A2(_0400_));
 sg13g2_nor2_2 _2090_ (.A(net301),
    .B(net298),
    .Y(_0402_));
 sg13g2_nand2_1 _2091_ (.Y(_0403_),
    .A(net303),
    .B(net295));
 sg13g2_nand3_1 _2092_ (.B(net287),
    .C(net281),
    .A(net293),
    .Y(_0404_));
 sg13g2_nand2_1 _2093_ (.Y(_0405_),
    .A(_0402_),
    .B(_0404_));
 sg13g2_nand3_1 _2094_ (.B(_0393_),
    .C(_0397_),
    .A(net306),
    .Y(_0406_));
 sg13g2_a21oi_1 _2095_ (.A1(_0401_),
    .A2(_0405_),
    .Y(_0407_),
    .B1(net307));
 sg13g2_nor2_1 _2096_ (.A(net308),
    .B(_0407_),
    .Y(_0408_));
 sg13g2_a21oi_2 _2097_ (.B1(net289),
    .Y(_0409_),
    .A2(_0389_),
    .A1(net284));
 sg13g2_o21ai_1 _2098_ (.B1(net293),
    .Y(_0410_),
    .A1(net286),
    .A2(_0390_));
 sg13g2_nor2_1 _2099_ (.A(net303),
    .B(_0409_),
    .Y(_0411_));
 sg13g2_a21oi_1 _2100_ (.A1(net295),
    .A2(_0411_),
    .Y(_0412_),
    .B1(net306));
 sg13g2_nor2_1 _2101_ (.A(_0326_),
    .B(_0347_),
    .Y(_0413_));
 sg13g2_a22oi_1 _2102_ (.Y(_0414_),
    .B1(_0412_),
    .B2(_0413_),
    .A2(_0408_),
    .A1(_0406_));
 sg13g2_nor2_1 _2103_ (.A(net295),
    .B(_0395_),
    .Y(_0415_));
 sg13g2_nand2_1 _2104_ (.Y(_0416_),
    .A(net291),
    .B(_0371_));
 sg13g2_a21o_1 _2105_ (.A2(net281),
    .A1(net289),
    .B1(net306),
    .X(_0417_));
 sg13g2_a221oi_1 _2106_ (.B2(net280),
    .C1(_0417_),
    .B1(_0410_),
    .A1(net298),
    .Y(_0418_),
    .A2(_0396_));
 sg13g2_nand2_1 _2107_ (.Y(_0419_),
    .A(net291),
    .B(_0377_));
 sg13g2_o21ai_1 _2108_ (.B1(net298),
    .Y(_0420_),
    .A1(net294),
    .A2(net283));
 sg13g2_inv_1 _2109_ (.Y(_0421_),
    .A(_0420_));
 sg13g2_nor2_1 _2110_ (.A(net288),
    .B(net282),
    .Y(_0422_));
 sg13g2_nor2_1 _2111_ (.A(_0355_),
    .B(_0385_),
    .Y(_0423_));
 sg13g2_o21ai_1 _2112_ (.B1(net294),
    .Y(_0424_),
    .A1(_0422_),
    .A2(_0423_));
 sg13g2_xnor2_1 _2113_ (.Y(_0425_),
    .A(_0368_),
    .B(_0373_));
 sg13g2_nor2_1 _2114_ (.A(net288),
    .B(net285),
    .Y(_0426_));
 sg13g2_a21oi_2 _2115_ (.B1(net289),
    .Y(_0427_),
    .A2(net286),
    .A1(_0355_));
 sg13g2_nand3_1 _2116_ (.B(_0390_),
    .C(_0425_),
    .A(net294),
    .Y(_0428_));
 sg13g2_o21ai_1 _2117_ (.B1(net289),
    .Y(_0429_),
    .A1(_0355_),
    .A2(net283));
 sg13g2_nor2_1 _2118_ (.A(net284),
    .B(_0390_),
    .Y(_0430_));
 sg13g2_o21ai_1 _2119_ (.B1(_0428_),
    .Y(_0431_),
    .A1(_0429_),
    .A2(_0430_));
 sg13g2_a221oi_1 _2120_ (.B2(net297),
    .C1(_0418_),
    .B1(_0431_),
    .A1(_0421_),
    .Y(_0432_),
    .A2(_0424_));
 sg13g2_nor2_1 _2121_ (.A(_0354_),
    .B(_0425_),
    .Y(_0433_));
 sg13g2_a21oi_1 _2122_ (.A1(net287),
    .A2(_0386_),
    .Y(_0434_),
    .B1(net293));
 sg13g2_o21ai_1 _2123_ (.B1(net290),
    .Y(_0435_),
    .A1(_0355_),
    .A2(_0385_));
 sg13g2_nor2_1 _2124_ (.A(net298),
    .B(net289),
    .Y(_0436_));
 sg13g2_nand3_1 _2125_ (.B(net284),
    .C(net283),
    .A(net287),
    .Y(_0437_));
 sg13g2_a221oi_1 _2126_ (.B2(_0437_),
    .C1(_0434_),
    .B1(_0436_),
    .A1(net289),
    .Y(_0438_),
    .A2(net281));
 sg13g2_xnor2_1 _2127_ (.Y(_0439_),
    .A(_0350_),
    .B(_0368_));
 sg13g2_nand4_1 _2128_ (.B(net294),
    .C(_0380_),
    .A(net300),
    .Y(_0440_),
    .D(_0439_));
 sg13g2_o21ai_1 _2129_ (.B1(_0440_),
    .Y(_0441_),
    .A1(_0433_),
    .A2(_0438_));
 sg13g2_a21o_1 _2130_ (.A2(_0441_),
    .A1(net307),
    .B1(_0432_),
    .X(_0442_));
 sg13g2_a21oi_1 _2131_ (.A1(net286),
    .A2(_0398_),
    .Y(_0443_),
    .B1(net307));
 sg13g2_o21ai_1 _2132_ (.B1(_0347_),
    .Y(_0444_),
    .A1(net285),
    .A2(_0398_));
 sg13g2_o21ai_1 _2133_ (.B1(_0444_),
    .Y(_0445_),
    .A1(net302),
    .A2(_0443_));
 sg13g2_nand2_1 _2134_ (.Y(_0446_),
    .A(net291),
    .B(_0439_));
 sg13g2_a21oi_1 _2135_ (.A1(_0427_),
    .A2(_0437_),
    .Y(_0447_),
    .B1(_0356_));
 sg13g2_nand2_1 _2136_ (.Y(_0448_),
    .A(_0446_),
    .B(_0447_));
 sg13g2_nand2_1 _2137_ (.Y(_0449_),
    .A(net291),
    .B(_0354_));
 sg13g2_nand2b_1 _2138_ (.Y(_0450_),
    .B(net280),
    .A_N(_0357_));
 sg13g2_a21oi_1 _2139_ (.A1(net286),
    .A2(_0449_),
    .Y(_0451_),
    .B1(net300));
 sg13g2_o21ai_1 _2140_ (.B1(_0451_),
    .Y(_0452_),
    .A1(net282),
    .A2(_0450_));
 sg13g2_a21o_1 _2141_ (.A2(_0452_),
    .A1(_0448_),
    .B1(net305),
    .X(_0453_));
 sg13g2_nand2_1 _2142_ (.Y(_0454_),
    .A(net305),
    .B(net301));
 sg13g2_nand3_1 _2143_ (.B(net285),
    .C(_0390_),
    .A(_0345_),
    .Y(_0455_));
 sg13g2_a21oi_1 _2144_ (.A1(net286),
    .A2(_0389_),
    .Y(_0456_),
    .B1(net297));
 sg13g2_nand3_1 _2145_ (.B(_0455_),
    .C(_0456_),
    .A(_0416_),
    .Y(_0457_));
 sg13g2_a21o_1 _2146_ (.A2(_0455_),
    .A1(_0416_),
    .B1(net300),
    .X(_0458_));
 sg13g2_and3_1 _2147_ (.X(_0459_),
    .A(_0418_),
    .B(_0457_),
    .C(_0458_));
 sg13g2_o21ai_1 _2148_ (.B1(_0326_),
    .Y(_0460_),
    .A1(_0454_),
    .A2(_0459_));
 sg13g2_a221oi_1 _2149_ (.B2(_0453_),
    .C1(_0460_),
    .B1(_0445_),
    .A1(net302),
    .Y(_0461_),
    .A2(_0442_));
 sg13g2_a21oi_1 _2150_ (.A1(net303),
    .A2(net280),
    .Y(_0462_),
    .B1(net284));
 sg13g2_a22oi_1 _2151_ (.Y(_0463_),
    .B1(_0462_),
    .B2(_0367_),
    .A2(_0427_),
    .A1(net295));
 sg13g2_nor3_1 _2152_ (.A(net284),
    .B(_0377_),
    .C(_0388_),
    .Y(_0464_));
 sg13g2_o21ai_1 _2153_ (.B1(net295),
    .Y(_0465_),
    .A1(net303),
    .A2(_0464_));
 sg13g2_o21ai_1 _2154_ (.B1(_0465_),
    .Y(_0466_),
    .A1(net283),
    .A2(_0463_));
 sg13g2_xnor2_1 _2155_ (.Y(_0467_),
    .A(_0425_),
    .B(_0427_));
 sg13g2_a22oi_1 _2156_ (.Y(_0468_),
    .B1(_0427_),
    .B2(_0437_),
    .A2(net286),
    .A1(net290));
 sg13g2_a21o_1 _2157_ (.A2(_0468_),
    .A1(_0467_),
    .B1(_0403_),
    .X(_0469_));
 sg13g2_nand3_1 _2158_ (.B(_0466_),
    .C(_0469_),
    .A(net305),
    .Y(_0470_));
 sg13g2_o21ai_1 _2159_ (.B1(net288),
    .Y(_0471_),
    .A1(net284),
    .A2(_0377_));
 sg13g2_nand2_1 _2160_ (.Y(_0472_),
    .A(_0355_),
    .B(net283));
 sg13g2_and2_1 _2161_ (.A(_0386_),
    .B(_0471_),
    .X(_0473_));
 sg13g2_a21o_1 _2162_ (.A2(_0471_),
    .A1(_0386_),
    .B1(net289),
    .X(_0474_));
 sg13g2_xnor2_1 _2163_ (.Y(_0475_),
    .A(_0351_),
    .B(_0373_));
 sg13g2_xnor2_1 _2164_ (.Y(_0476_),
    .A(_0350_),
    .B(_0373_));
 sg13g2_a21oi_1 _2165_ (.A1(net291),
    .A2(_0476_),
    .Y(_0477_),
    .B1(net297));
 sg13g2_nand2_1 _2166_ (.Y(_0478_),
    .A(_0356_),
    .B(_0420_));
 sg13g2_and2_1 _2167_ (.A(_0381_),
    .B(_0409_),
    .X(_0479_));
 sg13g2_a221oi_1 _2168_ (.B2(_0477_),
    .C1(_0479_),
    .B1(_0474_),
    .A1(_0356_),
    .Y(_0480_),
    .A2(_0420_));
 sg13g2_nand2_1 _2169_ (.Y(_0481_),
    .A(net294),
    .B(_0475_));
 sg13g2_nand4_1 _2170_ (.B(_0419_),
    .C(_0449_),
    .A(net285),
    .Y(_0482_),
    .D(_0481_));
 sg13g2_a221oi_1 _2171_ (.B2(_0341_),
    .C1(net305),
    .B1(_0482_),
    .A1(_0402_),
    .Y(_0483_),
    .A2(_0472_));
 sg13g2_o21ai_1 _2172_ (.B1(_0483_),
    .Y(_0484_),
    .A1(net303),
    .A2(_0480_));
 sg13g2_a21oi_1 _2173_ (.A1(_0470_),
    .A2(_0484_),
    .Y(_0485_),
    .B1(_0326_));
 sg13g2_nor3_2 _2174_ (.A(_0365_),
    .B(_0461_),
    .C(_0485_),
    .Y(_0486_));
 sg13g2_a221oi_1 _2175_ (.B2(_0385_),
    .C1(net282),
    .B1(net288),
    .A1(_0343_),
    .Y(_0487_),
    .A2(_0344_));
 sg13g2_a21o_1 _2176_ (.A2(_0377_),
    .A1(net291),
    .B1(_0487_),
    .X(_0488_));
 sg13g2_a21oi_1 _2177_ (.A1(_0458_),
    .A2(_0488_),
    .Y(_0489_),
    .B1(net304));
 sg13g2_o21ai_1 _2178_ (.B1(_0489_),
    .Y(_0490_),
    .A1(_0458_),
    .A2(_0488_));
 sg13g2_nor2_1 _2179_ (.A(net302),
    .B(_0425_),
    .Y(_0491_));
 sg13g2_a21oi_1 _2180_ (.A1(_0398_),
    .A2(_0491_),
    .Y(_0492_),
    .B1(net307));
 sg13g2_nor2_1 _2181_ (.A(_0345_),
    .B(_0425_),
    .Y(_0493_));
 sg13g2_a22oi_1 _2182_ (.Y(_0494_),
    .B1(_0493_),
    .B2(_0378_),
    .A2(_0487_),
    .A1(_0472_));
 sg13g2_a21oi_1 _2183_ (.A1(net288),
    .A2(_0377_),
    .Y(_0495_),
    .B1(net297));
 sg13g2_o21ai_1 _2184_ (.B1(net304),
    .Y(_0496_),
    .A1(net300),
    .A2(_0494_));
 sg13g2_a21o_1 _2185_ (.A2(_0495_),
    .A1(_0494_),
    .B1(_0496_),
    .X(_0497_));
 sg13g2_xnor2_1 _2186_ (.Y(_0498_),
    .A(net292),
    .B(_0473_));
 sg13g2_and2_1 _2187_ (.A(net302),
    .B(_0398_),
    .X(_0499_));
 sg13g2_a21oi_1 _2188_ (.A1(_0498_),
    .A2(_0499_),
    .Y(_0500_),
    .B1(net305));
 sg13g2_a221oi_1 _2189_ (.B2(_0500_),
    .C1(_0325_),
    .B1(_0497_),
    .A1(_0490_),
    .Y(_0501_),
    .A2(_0492_));
 sg13g2_a22oi_1 _2190_ (.Y(_0502_),
    .B1(_0471_),
    .B2(net294),
    .A2(_0434_),
    .A1(_0391_));
 sg13g2_o21ai_1 _2191_ (.B1(_0446_),
    .Y(_0503_),
    .A1(net286),
    .A2(_0377_));
 sg13g2_a221oi_1 _2192_ (.B2(_0410_),
    .C1(_0367_),
    .B1(net280),
    .A1(net287),
    .Y(_0504_),
    .A2(net283));
 sg13g2_a21oi_1 _2193_ (.A1(net304),
    .A2(_0503_),
    .Y(_0505_),
    .B1(_0476_));
 sg13g2_nor3_1 _2194_ (.A(net302),
    .B(net294),
    .C(_0475_),
    .Y(_0506_));
 sg13g2_o21ai_1 _2195_ (.B1(net300),
    .Y(_0507_),
    .A1(_0505_),
    .A2(_0506_));
 sg13g2_o21ai_1 _2196_ (.B1(net305),
    .Y(_0508_),
    .A1(_0403_),
    .A2(_0502_));
 sg13g2_nor2_1 _2197_ (.A(_0504_),
    .B(_0508_),
    .Y(_0509_));
 sg13g2_dfrbp_1 _2198_ (.CLK(net339),
    .RESET_B(net362),
    .D(_1071_),
    .Q_N(_1071_),
    .Q(\waggle_demo.ypos[1] ));
 sg13g2_dfrbp_1 _2199_ (.CLK(net339),
    .RESET_B(net362),
    .D(_0057_),
    .Q_N(_1090_),
    .Q(\waggle_demo.ypos[2] ));
 sg13g2_dfrbp_1 _2200_ (.CLK(net339),
    .RESET_B(net362),
    .D(_0058_),
    .Q_N(_1091_),
    .Q(\waggle_demo.ypos[3] ));
 sg13g2_dfrbp_1 _2201_ (.CLK(net340),
    .RESET_B(net363),
    .D(_0059_),
    .Q_N(_1092_),
    .Q(\waggle_demo.ypos[4] ));
 sg13g2_dfrbp_1 _2202_ (.CLK(net340),
    .RESET_B(net363),
    .D(_0060_),
    .Q_N(_1093_),
    .Q(\waggle_demo.ypos[5] ));
 sg13g2_dfrbp_1 _2203_ (.CLK(net341),
    .RESET_B(net364),
    .D(_0061_),
    .Q_N(_1094_),
    .Q(\waggle_demo.ypos[6] ));
 sg13g2_dfrbp_1 _2204_ (.CLK(net341),
    .RESET_B(net364),
    .D(_0062_),
    .Q_N(_1095_),
    .Q(\waggle_demo.ypos[7] ));
 sg13g2_dfrbp_1 _2205_ (.CLK(net340),
    .RESET_B(net363),
    .D(_0065_),
    .Q_N(_0065_),
    .Q(\frame[0] ));
 sg13g2_dfrbp_1 _2206_ (.CLK(net340),
    .RESET_B(net363),
    .D(_0025_),
    .Q_N(_0024_),
    .Q(\frame[1] ));
 sg13g2_dfrbp_1 _2207_ (.CLK(net340),
    .RESET_B(net363),
    .D(_0026_),
    .Q_N(_0016_),
    .Q(\frame[2] ));
 sg13g2_dfrbp_1 _2208_ (.CLK(net340),
    .RESET_B(net365),
    .D(_0027_),
    .Q_N(_0009_),
    .Q(\frame[3] ));
 sg13g2_dfrbp_1 _2209_ (.CLK(net341),
    .RESET_B(net363),
    .D(_0028_),
    .Q_N(_0011_),
    .Q(\frame[4] ));
 sg13g2_dfrbp_1 _2210_ (.CLK(net340),
    .RESET_B(net363),
    .D(_0029_),
    .Q_N(_0010_),
    .Q(\frame[5] ));
 sg13g2_dfrbp_1 _2211_ (.CLK(net340),
    .RESET_B(net363),
    .D(_0030_),
    .Q_N(_1096_),
    .Q(\frame[6] ));
 sg13g2_dfrbp_1 _2212_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net29),
    .D(net62),
    .Q_N(_1089_),
    .Q(hsync));
 sg13g2_dfrbp_1 _2213_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net53),
    .D(_0067_),
    .Q_N(_0064_),
    .Q(\hvsync_gen.vpos[0] ));
 sg13g2_dfrbp_1 _2214_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net51),
    .D(_0068_),
    .Q_N(_1088_),
    .Q(\hvsync_gen.vpos[1] ));
 sg13g2_dfrbp_1 _2215_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net49),
    .D(_0069_),
    .Q_N(_1087_),
    .Q(\hvsync_gen.vpos[2] ));
 sg13g2_dfrbp_1 _2216_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net47),
    .D(_0070_),
    .Q_N(_1086_),
    .Q(\hvsync_gen.vpos[3] ));
 sg13g2_dfrbp_1 _2217_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net45),
    .D(_0071_),
    .Q_N(_1085_),
    .Q(\hvsync_gen.vpos[4] ));
 sg13g2_dfrbp_1 _2218_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net37),
    .D(_0072_),
    .Q_N(_1084_),
    .Q(\hvsync_gen.vpos[5] ));
 sg13g2_dfrbp_1 _2219_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net35),
    .D(_0073_),
    .Q_N(_1083_),
    .Q(\hvsync_gen.vpos[6] ));
 sg13g2_dfrbp_1 _2220_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net33),
    .D(_0074_),
    .Q_N(_1082_),
    .Q(\hvsync_gen.vpos[7] ));
 sg13g2_dfrbp_1 _2221_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net31),
    .D(_0075_),
    .Q_N(_1081_),
    .Q(\hvsync_gen.vpos[8] ));
 sg13g2_dfrbp_1 _2222_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net55),
    .D(net70),
    .Q_N(_1097_),
    .Q(\hvsync_gen.vpos[9] ));
 sg13g2_dfrbp_1 _2223_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net30),
    .D(net74),
    .Q_N(_1080_),
    .Q(\hvsync_gen.vsync ));
 sg13g2_dllrq_1 _2224_ (.D(_0002_),
    .GATE_N(net23),
    .RESET_B(net39),
    .Q(\palette_inst.palette[0] ));
 sg13g2_dllrq_1 _2225_ (.D(_0003_),
    .GATE_N(net24),
    .RESET_B(net40),
    .Q(\palette_inst.palette[1] ));
 sg13g2_dllrq_1 _2226_ (.D(_0004_),
    .GATE_N(net25),
    .RESET_B(net41),
    .Q(\palette_inst.palette[2] ));
 sg13g2_dllrq_1 _2227_ (.D(_0005_),
    .GATE_N(net26),
    .RESET_B(net42),
    .Q(\palette_inst.palette[3] ));
 sg13g2_dllrq_1 _2228_ (.D(_0006_),
    .GATE_N(net27),
    .RESET_B(net43),
    .Q(\palette_inst.palette[4] ));
 sg13g2_dllrq_1 _2229_ (.D(_0007_),
    .GATE_N(net28),
    .RESET_B(net44),
    .Q(\palette_inst.palette[5] ));
 sg13g2_dfrbp_1 _2230_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net54),
    .D(_0077_),
    .Q_N(_0063_),
    .Q(\hpos[0] ));
 sg13g2_dfrbp_1 _2231_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net52),
    .D(net76),
    .Q_N(_1079_),
    .Q(\hpos[1] ));
 sg13g2_dfrbp_1 _2232_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net50),
    .D(_0079_),
    .Q_N(_1078_),
    .Q(\hpos[2] ));
 sg13g2_dfrbp_1 _2233_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net48),
    .D(_0080_),
    .Q_N(_1077_),
    .Q(\hpos[3] ));
 sg13g2_dfrbp_1 _2234_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net46),
    .D(_0081_),
    .Q_N(_1076_),
    .Q(\hpos[4] ));
 sg13g2_dfrbp_1 _2235_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net38),
    .D(_0082_),
    .Q_N(_1075_),
    .Q(\hpos[5] ));
 sg13g2_dfrbp_1 _2236_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net36),
    .D(_0083_),
    .Q_N(_1074_),
    .Q(\hpos[6] ));
 sg13g2_dfrbp_1 _2237_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net34),
    .D(_0084_),
    .Q_N(_1073_),
    .Q(\hpos[7] ));
 sg13g2_dfrbp_1 _2238_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net32),
    .D(net66),
    .Q_N(_1072_),
    .Q(\hpos[8] ));
 sg13g2_dfrbp_1 _2239_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net56),
    .D(_0086_),
    .Q_N(_1098_),
    .Q(\hpos[9] ));
 sg13g2_dfrbp_1 _2240_ (.CLK(net342),
    .RESET_B(net366),
    .D(_0066_),
    .Q_N(_0066_),
    .Q(\waggle_demo.xpos[0] ));
 sg13g2_dfrbp_1 _2241_ (.CLK(net339),
    .RESET_B(net362),
    .D(_0050_),
    .Q_N(_1099_),
    .Q(\waggle_demo.xpos[1] ));
 sg13g2_dfrbp_1 _2242_ (.CLK(net339),
    .RESET_B(net362),
    .D(_0051_),
    .Q_N(_1100_),
    .Q(\waggle_demo.xpos[2] ));
 sg13g2_dfrbp_1 _2243_ (.CLK(net342),
    .RESET_B(net364),
    .D(_0052_),
    .Q_N(_1101_),
    .Q(\waggle_demo.xpos[3] ));
 sg13g2_dfrbp_1 _2244_ (.CLK(net341),
    .RESET_B(net365),
    .D(_0053_),
    .Q_N(_1102_),
    .Q(\waggle_demo.xpos[4] ));
 sg13g2_dfrbp_1 _2245_ (.CLK(net341),
    .RESET_B(net364),
    .D(_0054_),
    .Q_N(_1103_),
    .Q(\waggle_demo.xpos[5] ));
 sg13g2_dfrbp_1 _2246_ (.CLK(net341),
    .RESET_B(net364),
    .D(_0055_),
    .Q_N(_1104_),
    .Q(\waggle_demo.xpos[6] ));
 sg13g2_dfrbp_1 _2247_ (.CLK(net341),
    .RESET_B(net364),
    .D(_0056_),
    .Q_N(_1105_),
    .Q(\waggle_demo.xpos[7] ));
 sg13g2_dfrbp_1 _2248_ (.CLK(net343),
    .RESET_B(net368),
    .D(_0031_),
    .Q_N(_1106_),
    .Q(\waggle_demo.p0[1] ));
 sg13g2_dfrbp_1 _2249_ (.CLK(net344),
    .RESET_B(net367),
    .D(_0032_),
    .Q_N(_1107_),
    .Q(\waggle_demo.p0[2] ));
 sg13g2_dfrbp_1 _2250_ (.CLK(net343),
    .RESET_B(net367),
    .D(_0033_),
    .Q_N(_0012_),
    .Q(\waggle_demo.p0[3] ));
 sg13g2_dfrbp_1 _2251_ (.CLK(net343),
    .RESET_B(net367),
    .D(_0034_),
    .Q_N(_1108_),
    .Q(\waggle_demo.p0[4] ));
 sg13g2_dfrbp_1 _2252_ (.CLK(net343),
    .RESET_B(net367),
    .D(_0035_),
    .Q_N(_0013_),
    .Q(\waggle_demo.p0[5] ));
 sg13g2_dfrbp_1 _2253_ (.CLK(net343),
    .RESET_B(net367),
    .D(_0036_),
    .Q_N(_1109_),
    .Q(\waggle_demo.p0[6] ));
 sg13g2_dfrbp_1 _2254_ (.CLK(net343),
    .RESET_B(net367),
    .D(_0037_),
    .Q_N(_1110_),
    .Q(\waggle_demo.p0[7] ));
 sg13g2_dfrbp_1 _2255_ (.CLK(net343),
    .RESET_B(net367),
    .D(_0038_),
    .Q_N(_1111_),
    .Q(\waggle_demo.p0[8] ));
 sg13g2_dfrbp_1 _2256_ (.CLK(net343),
    .RESET_B(net367),
    .D(_0039_),
    .Q_N(_1112_),
    .Q(\waggle_demo.p0[9] ));
 sg13g2_dfrbp_1 _2257_ (.CLK(net339),
    .RESET_B(net362),
    .D(_0040_),
    .Q_N(_0023_),
    .Q(\waggle_demo.p1[0] ));
 sg13g2_dfrbp_1 _2258_ (.CLK(net344),
    .RESET_B(net369),
    .D(_0041_),
    .Q_N(_0019_),
    .Q(\waggle_demo.p1[1] ));
 sg13g2_dfrbp_1 _2259_ (.CLK(net339),
    .RESET_B(net362),
    .D(_0042_),
    .Q_N(_0020_),
    .Q(\waggle_demo.p1[2] ));
 sg13g2_dfrbp_1 _2260_ (.CLK(net344),
    .RESET_B(net369),
    .D(_0043_),
    .Q_N(_0014_),
    .Q(\waggle_demo.p1[3] ));
 sg13g2_dfrbp_1 _2261_ (.CLK(net344),
    .RESET_B(net369),
    .D(_0044_),
    .Q_N(_0018_),
    .Q(\waggle_demo.p1[4] ));
 sg13g2_dfrbp_1 _2262_ (.CLK(net344),
    .RESET_B(net369),
    .D(_0045_),
    .Q_N(_0015_),
    .Q(\waggle_demo.p1[5] ));
 sg13g2_dfrbp_1 _2263_ (.CLK(net344),
    .RESET_B(net369),
    .D(_0046_),
    .Q_N(_0017_),
    .Q(\waggle_demo.p1[6] ));
 sg13g2_dfrbp_1 _2264_ (.CLK(net344),
    .RESET_B(net369),
    .D(_0047_),
    .Q_N(_1113_),
    .Q(\waggle_demo.p1[7] ));
 sg13g2_dfrbp_1 _2265_ (.CLK(net342),
    .RESET_B(net366),
    .D(_0048_),
    .Q_N(_0022_),
    .Q(\waggle_demo.p1[8] ));
 sg13g2_dfrbp_1 _2266_ (.CLK(net339),
    .RESET_B(net362),
    .D(_0049_),
    .Q_N(_0021_),
    .Q(\waggle_demo.p1[9] ));
 sg13g2_tiehi _2223__30 (.L_HI(net30));
 sg13g2_tiehi _2221__31 (.L_HI(net31));
 sg13g2_tiehi _2238__32 (.L_HI(net32));
 sg13g2_tiehi _2220__33 (.L_HI(net33));
 sg13g2_tiehi _2237__34 (.L_HI(net34));
 sg13g2_tiehi _2219__35 (.L_HI(net35));
 sg13g2_tiehi _2236__36 (.L_HI(net36));
 sg13g2_tiehi _2218__37 (.L_HI(net37));
 sg13g2_tiehi _2235__38 (.L_HI(net38));
 sg13g2_tiehi _2224__39 (.L_HI(net39));
 sg13g2_tiehi _2225__40 (.L_HI(net40));
 sg13g2_tiehi _2226__41 (.L_HI(net41));
 sg13g2_tiehi _2227__42 (.L_HI(net42));
 sg13g2_tiehi _2228__43 (.L_HI(net43));
 sg13g2_tiehi _2229__44 (.L_HI(net44));
 sg13g2_tiehi _2217__45 (.L_HI(net45));
 sg13g2_tiehi _2234__46 (.L_HI(net46));
 sg13g2_tiehi _2216__47 (.L_HI(net47));
 sg13g2_tiehi _2233__48 (.L_HI(net48));
 sg13g2_tiehi _2215__49 (.L_HI(net49));
 sg13g2_tiehi _2232__50 (.L_HI(net50));
 sg13g2_tiehi _2214__51 (.L_HI(net51));
 sg13g2_tiehi _2231__52 (.L_HI(net52));
 sg13g2_tiehi _2213__53 (.L_HI(net53));
 sg13g2_tiehi _2230__54 (.L_HI(net54));
 sg13g2_tiehi _2222__55 (.L_HI(net55));
 sg13g2_tiehi _2239__56 (.L_HI(net56));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_patater_demokit_8 (.L_LO(net8));
 sg13g2_tielo tt_um_patater_demokit_9 (.L_LO(net9));
 sg13g2_tielo tt_um_patater_demokit_10 (.L_LO(net10));
 sg13g2_tielo tt_um_patater_demokit_11 (.L_LO(net11));
 sg13g2_tielo tt_um_patater_demokit_12 (.L_LO(net12));
 sg13g2_tielo tt_um_patater_demokit_13 (.L_LO(net13));
 sg13g2_tielo tt_um_patater_demokit_14 (.L_LO(net14));
 sg13g2_tielo tt_um_patater_demokit_15 (.L_LO(net15));
 sg13g2_tielo tt_um_patater_demokit_16 (.L_LO(net16));
 sg13g2_tielo tt_um_patater_demokit_17 (.L_LO(net17));
 sg13g2_tielo tt_um_patater_demokit_18 (.L_LO(net18));
 sg13g2_tielo tt_um_patater_demokit_19 (.L_LO(net19));
 sg13g2_tielo tt_um_patater_demokit_20 (.L_LO(net20));
 sg13g2_tielo tt_um_patater_demokit_21 (.L_LO(net21));
 sg13g2_tielo tt_um_patater_demokit_22 (.L_LO(net22));
 sg13g2_tielo _2224__23 (.L_LO(net23));
 sg13g2_tiehi _2212__29 (.L_HI(net29));
 sg13g2_buf_1 _2312_ (.A(\hvsync_gen.vsync ),
    .X(uo_out[3]));
 sg13g2_buf_1 _2313_ (.A(hsync),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout279 (.A(_1027_),
    .X(net279));
 sg13g2_buf_2 fanout280 (.A(_0388_),
    .X(net280));
 sg13g2_buf_2 fanout281 (.A(_0379_),
    .X(net281));
 sg13g2_buf_2 fanout282 (.A(_0379_),
    .X(net282));
 sg13g2_buf_4 fanout283 (.X(net283),
    .A(_0376_));
 sg13g2_buf_2 fanout284 (.A(_0372_),
    .X(net284));
 sg13g2_buf_1 fanout285 (.A(_0372_),
    .X(net285));
 sg13g2_buf_2 fanout286 (.A(_0371_),
    .X(net286));
 sg13g2_buf_2 fanout287 (.A(net288),
    .X(net287));
 sg13g2_buf_2 fanout288 (.A(_0354_),
    .X(net288));
 sg13g2_buf_2 fanout289 (.A(net290),
    .X(net289));
 sg13g2_buf_2 fanout290 (.A(net292),
    .X(net290));
 sg13g2_buf_2 fanout291 (.A(net292),
    .X(net291));
 sg13g2_buf_1 fanout292 (.A(_0346_),
    .X(net292));
 sg13g2_buf_2 fanout293 (.A(net294),
    .X(net293));
 sg13g2_buf_2 fanout294 (.A(_0345_),
    .X(net294));
 sg13g2_buf_2 fanout295 (.A(net297),
    .X(net295));
 sg13g2_buf_2 fanout296 (.A(net297),
    .X(net296));
 sg13g2_buf_2 fanout297 (.A(_0340_),
    .X(net297));
 sg13g2_buf_2 fanout298 (.A(net300),
    .X(net298));
 sg13g2_buf_1 fanout299 (.A(net300),
    .X(net299));
 sg13g2_buf_2 fanout300 (.A(_0339_),
    .X(net300));
 sg13g2_buf_2 fanout301 (.A(net302),
    .X(net301));
 sg13g2_buf_2 fanout302 (.A(_0335_),
    .X(net302));
 sg13g2_buf_2 fanout303 (.A(net304),
    .X(net303));
 sg13g2_buf_2 fanout304 (.A(_0334_),
    .X(net304));
 sg13g2_buf_2 fanout305 (.A(_0329_),
    .X(net305));
 sg13g2_buf_2 fanout306 (.A(net307),
    .X(net306));
 sg13g2_buf_2 fanout307 (.A(_0328_),
    .X(net307));
 sg13g2_buf_2 fanout308 (.A(_0325_),
    .X(net308));
 sg13g2_buf_2 fanout309 (.A(_0319_),
    .X(net309));
 sg13g2_buf_2 fanout310 (.A(_0317_),
    .X(net310));
 sg13g2_buf_2 fanout311 (.A(_0729_),
    .X(net311));
 sg13g2_buf_2 fanout312 (.A(net313),
    .X(net312));
 sg13g2_buf_2 fanout313 (.A(_0709_),
    .X(net313));
 sg13g2_buf_2 fanout314 (.A(_0691_),
    .X(net314));
 sg13g2_buf_2 fanout315 (.A(_0685_),
    .X(net315));
 sg13g2_buf_2 fanout316 (.A(net319),
    .X(net316));
 sg13g2_buf_2 fanout317 (.A(net319),
    .X(net317));
 sg13g2_buf_1 fanout318 (.A(net319),
    .X(net318));
 sg13g2_buf_1 fanout319 (.A(_0670_),
    .X(net319));
 sg13g2_buf_2 fanout320 (.A(net322),
    .X(net320));
 sg13g2_buf_2 fanout321 (.A(net322),
    .X(net321));
 sg13g2_buf_1 fanout322 (.A(_0669_),
    .X(net322));
 sg13g2_buf_2 fanout323 (.A(net327),
    .X(net323));
 sg13g2_buf_1 fanout324 (.A(net327),
    .X(net324));
 sg13g2_buf_2 fanout325 (.A(net327),
    .X(net325));
 sg13g2_buf_1 fanout326 (.A(net327),
    .X(net326));
 sg13g2_buf_1 fanout327 (.A(_0664_),
    .X(net327));
 sg13g2_buf_2 fanout328 (.A(net329),
    .X(net328));
 sg13g2_buf_4 fanout329 (.X(net329),
    .A(_0663_));
 sg13g2_buf_2 fanout330 (.A(_0658_),
    .X(net330));
 sg13g2_buf_2 fanout331 (.A(_0658_),
    .X(net331));
 sg13g2_buf_2 fanout332 (.A(net333),
    .X(net332));
 sg13g2_buf_2 fanout333 (.A(_0657_),
    .X(net333));
 sg13g2_buf_2 fanout334 (.A(_0212_),
    .X(net334));
 sg13g2_buf_2 fanout335 (.A(_0653_),
    .X(net335));
 sg13g2_buf_2 fanout336 (.A(_0651_),
    .X(net336));
 sg13g2_buf_2 fanout337 (.A(_0650_),
    .X(net337));
 sg13g2_buf_2 fanout338 (.A(net82),
    .X(net338));
 sg13g2_buf_4 fanout339 (.X(net339),
    .A(net342));
 sg13g2_buf_2 fanout340 (.A(net341),
    .X(net340));
 sg13g2_buf_2 fanout341 (.A(net342),
    .X(net341));
 sg13g2_buf_2 fanout342 (.A(\hvsync_gen.vsync ),
    .X(net342));
 sg13g2_buf_2 fanout343 (.A(net344),
    .X(net343));
 sg13g2_buf_4 fanout344 (.X(net344),
    .A(\hvsync_gen.vsync ));
 sg13g2_buf_2 fanout345 (.A(net60),
    .X(net345));
 sg13g2_buf_4 fanout346 (.X(net346),
    .A(net64));
 sg13g2_buf_2 fanout347 (.A(net348),
    .X(net347));
 sg13g2_buf_2 fanout348 (.A(net78),
    .X(net348));
 sg13g2_buf_4 fanout349 (.X(net349),
    .A(net83));
 sg13g2_buf_2 fanout350 (.A(net351),
    .X(net350));
 sg13g2_buf_4 fanout351 (.X(net351),
    .A(\hvsync_gen.vpos[3] ));
 sg13g2_buf_4 fanout352 (.X(net352),
    .A(net63));
 sg13g2_buf_4 fanout353 (.X(net353),
    .A(\hvsync_gen.vpos[1] ));
 sg13g2_buf_4 fanout354 (.X(net354),
    .A(net355));
 sg13g2_buf_4 fanout355 (.X(net355),
    .A(net80));
 sg13g2_buf_2 fanout356 (.A(net6),
    .X(net356));
 sg13g2_buf_2 fanout357 (.A(net5),
    .X(net357));
 sg13g2_buf_2 fanout358 (.A(ui_in[4]),
    .X(net358));
 sg13g2_buf_1 fanout359 (.A(ui_in[4]),
    .X(net359));
 sg13g2_buf_4 fanout360 (.X(net360),
    .A(ui_in[1]));
 sg13g2_buf_2 fanout361 (.A(ui_in[1]),
    .X(net361));
 sg13g2_buf_4 fanout362 (.X(net362),
    .A(net366));
 sg13g2_buf_4 fanout363 (.X(net363),
    .A(net365));
 sg13g2_buf_4 fanout364 (.X(net364),
    .A(net365));
 sg13g2_buf_2 fanout365 (.A(net366),
    .X(net365));
 sg13g2_buf_2 fanout366 (.A(rst_n),
    .X(net366));
 sg13g2_buf_4 fanout367 (.X(net367),
    .A(net368));
 sg13g2_buf_2 fanout368 (.A(net369),
    .X(net368));
 sg13g2_buf_4 fanout369 (.X(net369),
    .A(rst_n));
 sg13g2_buf_2 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_2 input2 (.A(ui_in[2]),
    .X(net2));
 sg13g2_buf_2 input3 (.A(ui_in[3]),
    .X(net3));
 sg13g2_buf_2 input4 (.A(ui_in[5]),
    .X(net4));
 sg13g2_buf_2 input5 (.A(ui_in[6]),
    .X(net5));
 sg13g2_buf_2 input6 (.A(ui_in[7]),
    .X(net6));
 sg13g2_tielo tt_um_patater_demokit_7 (.L_LO(net7));
 sg13g2_tielo _2225__24 (.L_LO(net24));
 sg13g2_tielo _2226__25 (.L_LO(net25));
 sg13g2_tielo _2227__26 (.L_LO(net26));
 sg13g2_tielo _2228__27 (.L_LO(net27));
 sg13g2_tielo _2229__28 (.L_LO(net28));
 sg13g2_buf_2 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .X(clknet_2_0__leaf_clk));
 sg13g2_buf_2 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .X(clknet_2_1__leaf_clk));
 sg13g2_buf_2 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .X(clknet_2_2__leaf_clk));
 sg13g2_buf_2 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .X(clknet_2_3__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_2_1__leaf_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_2_3__leaf_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(_0063_),
    .X(net57));
 sg13g2_dlygate4sd3_1 hold2 (.A(_0064_),
    .X(net58));
 sg13g2_dlygate4sd3_1 hold3 (.A(_0213_),
    .X(net59));
 sg13g2_dlygate4sd3_1 hold4 (.A(\hvsync_gen.vpos[7] ),
    .X(net60));
 sg13g2_dlygate4sd3_1 hold5 (.A(\hpos[8] ),
    .X(net61));
 sg13g2_dlygate4sd3_1 hold6 (.A(_0000_),
    .X(net62));
 sg13g2_dlygate4sd3_1 hold7 (.A(\hvsync_gen.vpos[2] ),
    .X(net63));
 sg13g2_dlygate4sd3_1 hold8 (.A(\hvsync_gen.vpos[6] ),
    .X(net64));
 sg13g2_dlygate4sd3_1 hold9 (.A(\hpos[7] ),
    .X(net65));
 sg13g2_dlygate4sd3_1 hold10 (.A(_0085_),
    .X(net66));
 sg13g2_dlygate4sd3_1 hold11 (.A(\hpos[2] ),
    .X(net67));
 sg13g2_dlygate4sd3_1 hold12 (.A(_0240_),
    .X(net68));
 sg13g2_dlygate4sd3_1 hold13 (.A(\hvsync_gen.vpos[9] ),
    .X(net69));
 sg13g2_dlygate4sd3_1 hold14 (.A(_0076_),
    .X(net70));
 sg13g2_dlygate4sd3_1 hold15 (.A(\hpos[6] ),
    .X(net71));
 sg13g2_dlygate4sd3_1 hold16 (.A(_0244_),
    .X(net72));
 sg13g2_dlygate4sd3_1 hold17 (.A(\hvsync_gen.vpos[8] ),
    .X(net73));
 sg13g2_dlygate4sd3_1 hold18 (.A(_0001_),
    .X(net74));
 sg13g2_dlygate4sd3_1 hold19 (.A(\hpos[1] ),
    .X(net75));
 sg13g2_dlygate4sd3_1 hold20 (.A(_0078_),
    .X(net76));
 sg13g2_dlygate4sd3_1 hold21 (.A(\hpos[9] ),
    .X(net77));
 sg13g2_dlygate4sd3_1 hold22 (.A(\hvsync_gen.vpos[5] ),
    .X(net78));
 sg13g2_dlygate4sd3_1 hold23 (.A(\hpos[3] ),
    .X(net79));
 sg13g2_dlygate4sd3_1 hold24 (.A(\hvsync_gen.vpos[0] ),
    .X(net80));
 sg13g2_dlygate4sd3_1 hold25 (.A(_0215_),
    .X(net81));
 sg13g2_dlygate4sd3_1 hold26 (.A(\hpos[5] ),
    .X(net82));
 sg13g2_dlygate4sd3_1 hold27 (.A(\hvsync_gen.vpos[4] ),
    .X(net83));
 sg13g2_dlygate4sd3_1 hold28 (.A(\hpos[4] ),
    .X(net84));
 sg13g2_dlygate4sd3_1 hold29 (.A(\hpos[1] ),
    .X(net85));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_fill_1 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_48 ();
 sg13g2_decap_8 FILLER_3_55 ();
 sg13g2_decap_8 FILLER_3_62 ();
 sg13g2_decap_8 FILLER_3_69 ();
 sg13g2_decap_4 FILLER_3_76 ();
 sg13g2_fill_2 FILLER_3_80 ();
 sg13g2_fill_2 FILLER_3_87 ();
 sg13g2_decap_8 FILLER_3_94 ();
 sg13g2_fill_1 FILLER_3_101 ();
 sg13g2_fill_2 FILLER_3_106 ();
 sg13g2_fill_1 FILLER_3_108 ();
 sg13g2_decap_8 FILLER_3_114 ();
 sg13g2_decap_4 FILLER_3_121 ();
 sg13g2_decap_4 FILLER_3_136 ();
 sg13g2_fill_2 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_146 ();
 sg13g2_fill_2 FILLER_3_153 ();
 sg13g2_fill_1 FILLER_3_155 ();
 sg13g2_decap_8 FILLER_3_162 ();
 sg13g2_decap_8 FILLER_3_169 ();
 sg13g2_decap_8 FILLER_3_176 ();
 sg13g2_decap_8 FILLER_3_183 ();
 sg13g2_decap_8 FILLER_3_190 ();
 sg13g2_decap_8 FILLER_3_197 ();
 sg13g2_decap_8 FILLER_3_204 ();
 sg13g2_decap_8 FILLER_3_211 ();
 sg13g2_decap_8 FILLER_3_218 ();
 sg13g2_decap_8 FILLER_3_225 ();
 sg13g2_decap_8 FILLER_3_232 ();
 sg13g2_decap_8 FILLER_3_239 ();
 sg13g2_decap_8 FILLER_3_246 ();
 sg13g2_decap_8 FILLER_3_253 ();
 sg13g2_decap_8 FILLER_3_260 ();
 sg13g2_decap_8 FILLER_3_267 ();
 sg13g2_decap_8 FILLER_3_274 ();
 sg13g2_decap_8 FILLER_3_281 ();
 sg13g2_decap_8 FILLER_3_288 ();
 sg13g2_decap_8 FILLER_3_295 ();
 sg13g2_decap_8 FILLER_3_302 ();
 sg13g2_decap_8 FILLER_3_309 ();
 sg13g2_decap_8 FILLER_3_316 ();
 sg13g2_decap_8 FILLER_3_323 ();
 sg13g2_decap_8 FILLER_3_330 ();
 sg13g2_decap_8 FILLER_3_337 ();
 sg13g2_decap_8 FILLER_3_344 ();
 sg13g2_decap_8 FILLER_3_351 ();
 sg13g2_decap_8 FILLER_3_358 ();
 sg13g2_decap_8 FILLER_3_365 ();
 sg13g2_decap_8 FILLER_3_372 ();
 sg13g2_decap_8 FILLER_3_379 ();
 sg13g2_decap_8 FILLER_3_386 ();
 sg13g2_decap_8 FILLER_3_393 ();
 sg13g2_decap_8 FILLER_3_400 ();
 sg13g2_fill_2 FILLER_3_407 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_fill_2 FILLER_4_21 ();
 sg13g2_fill_2 FILLER_4_28 ();
 sg13g2_fill_1 FILLER_4_30 ();
 sg13g2_fill_1 FILLER_4_39 ();
 sg13g2_fill_1 FILLER_4_55 ();
 sg13g2_fill_2 FILLER_4_62 ();
 sg13g2_fill_1 FILLER_4_64 ();
 sg13g2_fill_1 FILLER_4_87 ();
 sg13g2_decap_4 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_177 ();
 sg13g2_decap_8 FILLER_4_184 ();
 sg13g2_decap_8 FILLER_4_191 ();
 sg13g2_decap_8 FILLER_4_198 ();
 sg13g2_decap_8 FILLER_4_205 ();
 sg13g2_decap_8 FILLER_4_212 ();
 sg13g2_decap_8 FILLER_4_219 ();
 sg13g2_decap_8 FILLER_4_226 ();
 sg13g2_decap_8 FILLER_4_233 ();
 sg13g2_decap_8 FILLER_4_240 ();
 sg13g2_decap_8 FILLER_4_247 ();
 sg13g2_decap_8 FILLER_4_254 ();
 sg13g2_decap_8 FILLER_4_261 ();
 sg13g2_decap_8 FILLER_4_268 ();
 sg13g2_decap_8 FILLER_4_275 ();
 sg13g2_decap_8 FILLER_4_282 ();
 sg13g2_decap_8 FILLER_4_289 ();
 sg13g2_decap_8 FILLER_4_296 ();
 sg13g2_decap_8 FILLER_4_303 ();
 sg13g2_decap_8 FILLER_4_310 ();
 sg13g2_decap_8 FILLER_4_317 ();
 sg13g2_decap_8 FILLER_4_324 ();
 sg13g2_decap_8 FILLER_4_331 ();
 sg13g2_decap_8 FILLER_4_338 ();
 sg13g2_decap_8 FILLER_4_345 ();
 sg13g2_decap_8 FILLER_4_352 ();
 sg13g2_decap_8 FILLER_4_359 ();
 sg13g2_decap_8 FILLER_4_366 ();
 sg13g2_decap_8 FILLER_4_373 ();
 sg13g2_decap_8 FILLER_4_380 ();
 sg13g2_decap_8 FILLER_4_387 ();
 sg13g2_decap_8 FILLER_4_394 ();
 sg13g2_decap_8 FILLER_4_401 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_4 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_31 ();
 sg13g2_fill_1 FILLER_5_38 ();
 sg13g2_fill_2 FILLER_5_48 ();
 sg13g2_fill_1 FILLER_5_60 ();
 sg13g2_fill_1 FILLER_5_65 ();
 sg13g2_fill_1 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_78 ();
 sg13g2_fill_2 FILLER_5_85 ();
 sg13g2_fill_1 FILLER_5_87 ();
 sg13g2_decap_8 FILLER_5_92 ();
 sg13g2_decap_8 FILLER_5_109 ();
 sg13g2_decap_8 FILLER_5_116 ();
 sg13g2_decap_4 FILLER_5_123 ();
 sg13g2_decap_4 FILLER_5_138 ();
 sg13g2_fill_1 FILLER_5_142 ();
 sg13g2_decap_4 FILLER_5_148 ();
 sg13g2_fill_1 FILLER_5_152 ();
 sg13g2_decap_4 FILLER_5_159 ();
 sg13g2_fill_1 FILLER_5_163 ();
 sg13g2_decap_8 FILLER_5_190 ();
 sg13g2_decap_8 FILLER_5_197 ();
 sg13g2_decap_8 FILLER_5_204 ();
 sg13g2_decap_8 FILLER_5_211 ();
 sg13g2_decap_8 FILLER_5_218 ();
 sg13g2_decap_8 FILLER_5_225 ();
 sg13g2_decap_8 FILLER_5_232 ();
 sg13g2_decap_8 FILLER_5_239 ();
 sg13g2_decap_8 FILLER_5_246 ();
 sg13g2_decap_8 FILLER_5_253 ();
 sg13g2_decap_8 FILLER_5_260 ();
 sg13g2_decap_8 FILLER_5_267 ();
 sg13g2_decap_8 FILLER_5_274 ();
 sg13g2_decap_8 FILLER_5_281 ();
 sg13g2_decap_8 FILLER_5_288 ();
 sg13g2_decap_8 FILLER_5_295 ();
 sg13g2_decap_8 FILLER_5_302 ();
 sg13g2_decap_8 FILLER_5_309 ();
 sg13g2_decap_8 FILLER_5_316 ();
 sg13g2_decap_8 FILLER_5_323 ();
 sg13g2_decap_8 FILLER_5_330 ();
 sg13g2_decap_8 FILLER_5_337 ();
 sg13g2_decap_8 FILLER_5_344 ();
 sg13g2_decap_8 FILLER_5_351 ();
 sg13g2_decap_8 FILLER_5_358 ();
 sg13g2_decap_8 FILLER_5_365 ();
 sg13g2_decap_8 FILLER_5_372 ();
 sg13g2_decap_8 FILLER_5_379 ();
 sg13g2_decap_8 FILLER_5_386 ();
 sg13g2_decap_8 FILLER_5_393 ();
 sg13g2_decap_8 FILLER_5_400 ();
 sg13g2_fill_2 FILLER_5_407 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_4 FILLER_6_7 ();
 sg13g2_fill_1 FILLER_6_26 ();
 sg13g2_fill_1 FILLER_6_60 ();
 sg13g2_fill_2 FILLER_6_66 ();
 sg13g2_decap_4 FILLER_6_85 ();
 sg13g2_decap_4 FILLER_6_110 ();
 sg13g2_fill_1 FILLER_6_114 ();
 sg13g2_fill_2 FILLER_6_134 ();
 sg13g2_fill_1 FILLER_6_146 ();
 sg13g2_fill_2 FILLER_6_155 ();
 sg13g2_fill_2 FILLER_6_167 ();
 sg13g2_decap_8 FILLER_6_179 ();
 sg13g2_decap_8 FILLER_6_186 ();
 sg13g2_decap_8 FILLER_6_193 ();
 sg13g2_decap_8 FILLER_6_200 ();
 sg13g2_decap_8 FILLER_6_207 ();
 sg13g2_decap_8 FILLER_6_214 ();
 sg13g2_decap_8 FILLER_6_221 ();
 sg13g2_decap_8 FILLER_6_228 ();
 sg13g2_decap_8 FILLER_6_235 ();
 sg13g2_decap_8 FILLER_6_242 ();
 sg13g2_decap_8 FILLER_6_249 ();
 sg13g2_decap_8 FILLER_6_256 ();
 sg13g2_decap_8 FILLER_6_263 ();
 sg13g2_decap_8 FILLER_6_270 ();
 sg13g2_decap_8 FILLER_6_277 ();
 sg13g2_decap_8 FILLER_6_284 ();
 sg13g2_decap_8 FILLER_6_291 ();
 sg13g2_decap_8 FILLER_6_298 ();
 sg13g2_decap_8 FILLER_6_305 ();
 sg13g2_decap_8 FILLER_6_312 ();
 sg13g2_decap_8 FILLER_6_319 ();
 sg13g2_decap_8 FILLER_6_326 ();
 sg13g2_decap_8 FILLER_6_333 ();
 sg13g2_decap_8 FILLER_6_340 ();
 sg13g2_decap_8 FILLER_6_347 ();
 sg13g2_decap_8 FILLER_6_354 ();
 sg13g2_decap_8 FILLER_6_361 ();
 sg13g2_decap_8 FILLER_6_368 ();
 sg13g2_decap_8 FILLER_6_375 ();
 sg13g2_decap_8 FILLER_6_382 ();
 sg13g2_decap_8 FILLER_6_389 ();
 sg13g2_decap_8 FILLER_6_396 ();
 sg13g2_decap_4 FILLER_6_403 ();
 sg13g2_fill_2 FILLER_6_407 ();
 sg13g2_decap_4 FILLER_7_0 ();
 sg13g2_fill_2 FILLER_7_4 ();
 sg13g2_fill_2 FILLER_7_19 ();
 sg13g2_decap_8 FILLER_7_30 ();
 sg13g2_decap_4 FILLER_7_37 ();
 sg13g2_fill_1 FILLER_7_54 ();
 sg13g2_decap_8 FILLER_7_60 ();
 sg13g2_decap_4 FILLER_7_67 ();
 sg13g2_fill_1 FILLER_7_71 ();
 sg13g2_fill_1 FILLER_7_77 ();
 sg13g2_fill_2 FILLER_7_88 ();
 sg13g2_fill_1 FILLER_7_90 ();
 sg13g2_decap_4 FILLER_7_102 ();
 sg13g2_decap_4 FILLER_7_149 ();
 sg13g2_fill_1 FILLER_7_153 ();
 sg13g2_decap_8 FILLER_7_179 ();
 sg13g2_decap_8 FILLER_7_186 ();
 sg13g2_decap_8 FILLER_7_193 ();
 sg13g2_decap_4 FILLER_7_200 ();
 sg13g2_fill_2 FILLER_7_204 ();
 sg13g2_decap_8 FILLER_7_218 ();
 sg13g2_decap_8 FILLER_7_225 ();
 sg13g2_decap_8 FILLER_7_232 ();
 sg13g2_decap_8 FILLER_7_239 ();
 sg13g2_decap_8 FILLER_7_246 ();
 sg13g2_decap_8 FILLER_7_253 ();
 sg13g2_decap_8 FILLER_7_260 ();
 sg13g2_decap_8 FILLER_7_267 ();
 sg13g2_decap_8 FILLER_7_274 ();
 sg13g2_decap_8 FILLER_7_281 ();
 sg13g2_decap_8 FILLER_7_288 ();
 sg13g2_decap_8 FILLER_7_295 ();
 sg13g2_decap_8 FILLER_7_302 ();
 sg13g2_decap_8 FILLER_7_309 ();
 sg13g2_decap_8 FILLER_7_316 ();
 sg13g2_decap_8 FILLER_7_323 ();
 sg13g2_decap_8 FILLER_7_330 ();
 sg13g2_decap_8 FILLER_7_337 ();
 sg13g2_decap_8 FILLER_7_344 ();
 sg13g2_decap_8 FILLER_7_351 ();
 sg13g2_decap_8 FILLER_7_358 ();
 sg13g2_decap_8 FILLER_7_365 ();
 sg13g2_decap_8 FILLER_7_372 ();
 sg13g2_decap_8 FILLER_7_379 ();
 sg13g2_decap_8 FILLER_7_386 ();
 sg13g2_decap_8 FILLER_7_393 ();
 sg13g2_decap_8 FILLER_7_400 ();
 sg13g2_fill_2 FILLER_7_407 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_fill_2 FILLER_8_56 ();
 sg13g2_fill_1 FILLER_8_58 ();
 sg13g2_fill_2 FILLER_8_73 ();
 sg13g2_fill_1 FILLER_8_75 ();
 sg13g2_decap_4 FILLER_8_89 ();
 sg13g2_fill_2 FILLER_8_114 ();
 sg13g2_fill_1 FILLER_8_121 ();
 sg13g2_fill_2 FILLER_8_133 ();
 sg13g2_fill_1 FILLER_8_145 ();
 sg13g2_fill_2 FILLER_8_158 ();
 sg13g2_decap_4 FILLER_8_180 ();
 sg13g2_fill_2 FILLER_8_184 ();
 sg13g2_fill_2 FILLER_8_220 ();
 sg13g2_fill_1 FILLER_8_222 ();
 sg13g2_fill_1 FILLER_8_228 ();
 sg13g2_decap_8 FILLER_8_240 ();
 sg13g2_decap_8 FILLER_8_247 ();
 sg13g2_fill_1 FILLER_8_254 ();
 sg13g2_decap_8 FILLER_8_258 ();
 sg13g2_decap_8 FILLER_8_265 ();
 sg13g2_decap_8 FILLER_8_272 ();
 sg13g2_decap_8 FILLER_8_279 ();
 sg13g2_decap_8 FILLER_8_286 ();
 sg13g2_decap_8 FILLER_8_293 ();
 sg13g2_decap_8 FILLER_8_300 ();
 sg13g2_decap_8 FILLER_8_307 ();
 sg13g2_decap_8 FILLER_8_314 ();
 sg13g2_decap_8 FILLER_8_321 ();
 sg13g2_decap_8 FILLER_8_328 ();
 sg13g2_decap_8 FILLER_8_335 ();
 sg13g2_decap_8 FILLER_8_342 ();
 sg13g2_decap_8 FILLER_8_349 ();
 sg13g2_decap_8 FILLER_8_356 ();
 sg13g2_decap_8 FILLER_8_363 ();
 sg13g2_decap_8 FILLER_8_370 ();
 sg13g2_decap_8 FILLER_8_377 ();
 sg13g2_decap_8 FILLER_8_384 ();
 sg13g2_decap_8 FILLER_8_391 ();
 sg13g2_decap_8 FILLER_8_398 ();
 sg13g2_decap_4 FILLER_8_405 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_fill_2 FILLER_9_7 ();
 sg13g2_fill_1 FILLER_9_9 ();
 sg13g2_fill_2 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_fill_2 FILLER_9_42 ();
 sg13g2_fill_2 FILLER_9_73 ();
 sg13g2_fill_1 FILLER_9_75 ();
 sg13g2_decap_8 FILLER_9_94 ();
 sg13g2_decap_8 FILLER_9_106 ();
 sg13g2_fill_2 FILLER_9_118 ();
 sg13g2_fill_1 FILLER_9_120 ();
 sg13g2_fill_2 FILLER_9_153 ();
 sg13g2_fill_1 FILLER_9_155 ();
 sg13g2_decap_8 FILLER_9_165 ();
 sg13g2_decap_8 FILLER_9_172 ();
 sg13g2_decap_4 FILLER_9_195 ();
 sg13g2_fill_2 FILLER_9_207 ();
 sg13g2_fill_1 FILLER_9_209 ();
 sg13g2_fill_1 FILLER_9_215 ();
 sg13g2_decap_8 FILLER_9_265 ();
 sg13g2_decap_8 FILLER_9_272 ();
 sg13g2_decap_8 FILLER_9_279 ();
 sg13g2_decap_8 FILLER_9_286 ();
 sg13g2_decap_8 FILLER_9_293 ();
 sg13g2_decap_8 FILLER_9_300 ();
 sg13g2_decap_8 FILLER_9_307 ();
 sg13g2_decap_8 FILLER_9_314 ();
 sg13g2_decap_8 FILLER_9_321 ();
 sg13g2_decap_8 FILLER_9_328 ();
 sg13g2_decap_8 FILLER_9_335 ();
 sg13g2_decap_8 FILLER_9_342 ();
 sg13g2_decap_8 FILLER_9_349 ();
 sg13g2_decap_8 FILLER_9_356 ();
 sg13g2_decap_8 FILLER_9_363 ();
 sg13g2_decap_8 FILLER_9_370 ();
 sg13g2_decap_8 FILLER_9_377 ();
 sg13g2_decap_8 FILLER_9_384 ();
 sg13g2_decap_8 FILLER_9_391 ();
 sg13g2_decap_8 FILLER_9_398 ();
 sg13g2_decap_4 FILLER_9_405 ();
 sg13g2_decap_4 FILLER_10_0 ();
 sg13g2_fill_2 FILLER_10_4 ();
 sg13g2_fill_2 FILLER_10_37 ();
 sg13g2_fill_2 FILLER_10_51 ();
 sg13g2_fill_1 FILLER_10_53 ();
 sg13g2_fill_1 FILLER_10_74 ();
 sg13g2_fill_2 FILLER_10_86 ();
 sg13g2_fill_2 FILLER_10_118 ();
 sg13g2_decap_8 FILLER_10_132 ();
 sg13g2_decap_8 FILLER_10_139 ();
 sg13g2_fill_2 FILLER_10_146 ();
 sg13g2_fill_2 FILLER_10_158 ();
 sg13g2_decap_8 FILLER_10_165 ();
 sg13g2_decap_8 FILLER_10_172 ();
 sg13g2_fill_1 FILLER_10_221 ();
 sg13g2_decap_4 FILLER_10_238 ();
 sg13g2_fill_2 FILLER_10_242 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_fill_2 FILLER_11_14 ();
 sg13g2_decap_4 FILLER_11_27 ();
 sg13g2_fill_1 FILLER_11_36 ();
 sg13g2_fill_2 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_53 ();
 sg13g2_fill_2 FILLER_11_60 ();
 sg13g2_fill_1 FILLER_11_62 ();
 sg13g2_decap_4 FILLER_11_77 ();
 sg13g2_fill_2 FILLER_11_81 ();
 sg13g2_fill_2 FILLER_11_88 ();
 sg13g2_fill_1 FILLER_11_95 ();
 sg13g2_decap_8 FILLER_11_103 ();
 sg13g2_decap_8 FILLER_11_110 ();
 sg13g2_fill_1 FILLER_11_117 ();
 sg13g2_fill_1 FILLER_11_132 ();
 sg13g2_fill_1 FILLER_11_149 ();
 sg13g2_fill_2 FILLER_11_155 ();
 sg13g2_fill_1 FILLER_11_157 ();
 sg13g2_fill_2 FILLER_11_163 ();
 sg13g2_decap_8 FILLER_11_177 ();
 sg13g2_fill_2 FILLER_11_201 ();
 sg13g2_fill_1 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_fill_2 FILLER_11_217 ();
 sg13g2_fill_2 FILLER_11_236 ();
 sg13g2_decap_8 FILLER_11_277 ();
 sg13g2_decap_8 FILLER_11_284 ();
 sg13g2_decap_8 FILLER_11_291 ();
 sg13g2_decap_8 FILLER_11_298 ();
 sg13g2_decap_8 FILLER_11_305 ();
 sg13g2_decap_8 FILLER_11_312 ();
 sg13g2_decap_8 FILLER_11_319 ();
 sg13g2_decap_8 FILLER_11_326 ();
 sg13g2_decap_8 FILLER_11_333 ();
 sg13g2_decap_8 FILLER_11_340 ();
 sg13g2_decap_8 FILLER_11_347 ();
 sg13g2_decap_8 FILLER_11_354 ();
 sg13g2_decap_8 FILLER_11_361 ();
 sg13g2_decap_8 FILLER_11_368 ();
 sg13g2_decap_8 FILLER_11_375 ();
 sg13g2_decap_8 FILLER_11_382 ();
 sg13g2_decap_8 FILLER_11_389 ();
 sg13g2_decap_8 FILLER_11_396 ();
 sg13g2_decap_4 FILLER_11_403 ();
 sg13g2_fill_2 FILLER_11_407 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_4 FILLER_12_34 ();
 sg13g2_fill_2 FILLER_12_53 ();
 sg13g2_fill_2 FILLER_12_64 ();
 sg13g2_fill_1 FILLER_12_66 ();
 sg13g2_decap_4 FILLER_12_71 ();
 sg13g2_fill_2 FILLER_12_84 ();
 sg13g2_fill_1 FILLER_12_92 ();
 sg13g2_fill_2 FILLER_12_101 ();
 sg13g2_fill_1 FILLER_12_103 ();
 sg13g2_fill_1 FILLER_12_108 ();
 sg13g2_fill_1 FILLER_12_114 ();
 sg13g2_fill_2 FILLER_12_130 ();
 sg13g2_fill_1 FILLER_12_137 ();
 sg13g2_fill_2 FILLER_12_143 ();
 sg13g2_decap_8 FILLER_12_181 ();
 sg13g2_fill_2 FILLER_12_188 ();
 sg13g2_fill_2 FILLER_12_198 ();
 sg13g2_decap_8 FILLER_12_208 ();
 sg13g2_decap_8 FILLER_12_215 ();
 sg13g2_fill_1 FILLER_12_222 ();
 sg13g2_fill_2 FILLER_12_242 ();
 sg13g2_fill_1 FILLER_12_244 ();
 sg13g2_decap_8 FILLER_12_267 ();
 sg13g2_decap_8 FILLER_12_274 ();
 sg13g2_decap_8 FILLER_12_281 ();
 sg13g2_decap_8 FILLER_12_288 ();
 sg13g2_decap_8 FILLER_12_295 ();
 sg13g2_decap_8 FILLER_12_302 ();
 sg13g2_decap_8 FILLER_12_309 ();
 sg13g2_decap_8 FILLER_12_316 ();
 sg13g2_decap_8 FILLER_12_323 ();
 sg13g2_decap_8 FILLER_12_330 ();
 sg13g2_decap_8 FILLER_12_337 ();
 sg13g2_decap_8 FILLER_12_344 ();
 sg13g2_decap_8 FILLER_12_351 ();
 sg13g2_decap_8 FILLER_12_358 ();
 sg13g2_decap_8 FILLER_12_365 ();
 sg13g2_decap_8 FILLER_12_372 ();
 sg13g2_decap_8 FILLER_12_379 ();
 sg13g2_decap_8 FILLER_12_386 ();
 sg13g2_decap_8 FILLER_12_393 ();
 sg13g2_decap_8 FILLER_12_400 ();
 sg13g2_fill_2 FILLER_12_407 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_4 FILLER_13_28 ();
 sg13g2_fill_2 FILLER_13_32 ();
 sg13g2_fill_1 FILLER_13_52 ();
 sg13g2_decap_4 FILLER_13_78 ();
 sg13g2_fill_2 FILLER_13_82 ();
 sg13g2_decap_8 FILLER_13_92 ();
 sg13g2_fill_1 FILLER_13_99 ();
 sg13g2_fill_1 FILLER_13_110 ();
 sg13g2_decap_4 FILLER_13_128 ();
 sg13g2_fill_1 FILLER_13_132 ();
 sg13g2_decap_8 FILLER_13_145 ();
 sg13g2_decap_4 FILLER_13_152 ();
 sg13g2_fill_1 FILLER_13_156 ();
 sg13g2_decap_4 FILLER_13_180 ();
 sg13g2_fill_1 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_216 ();
 sg13g2_fill_2 FILLER_13_242 ();
 sg13g2_fill_1 FILLER_13_244 ();
 sg13g2_fill_2 FILLER_13_258 ();
 sg13g2_decap_8 FILLER_13_286 ();
 sg13g2_decap_8 FILLER_13_293 ();
 sg13g2_decap_8 FILLER_13_300 ();
 sg13g2_decap_8 FILLER_13_307 ();
 sg13g2_decap_8 FILLER_13_314 ();
 sg13g2_decap_8 FILLER_13_321 ();
 sg13g2_decap_8 FILLER_13_328 ();
 sg13g2_decap_8 FILLER_13_335 ();
 sg13g2_decap_8 FILLER_13_342 ();
 sg13g2_decap_8 FILLER_13_349 ();
 sg13g2_decap_8 FILLER_13_356 ();
 sg13g2_decap_8 FILLER_13_363 ();
 sg13g2_decap_8 FILLER_13_370 ();
 sg13g2_decap_8 FILLER_13_377 ();
 sg13g2_decap_8 FILLER_13_384 ();
 sg13g2_decap_8 FILLER_13_391 ();
 sg13g2_decap_8 FILLER_13_398 ();
 sg13g2_decap_4 FILLER_13_405 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_4 FILLER_14_35 ();
 sg13g2_fill_1 FILLER_14_39 ();
 sg13g2_fill_2 FILLER_14_44 ();
 sg13g2_decap_8 FILLER_14_50 ();
 sg13g2_fill_2 FILLER_14_57 ();
 sg13g2_fill_1 FILLER_14_64 ();
 sg13g2_decap_8 FILLER_14_74 ();
 sg13g2_fill_1 FILLER_14_81 ();
 sg13g2_fill_1 FILLER_14_88 ();
 sg13g2_fill_2 FILLER_14_98 ();
 sg13g2_fill_2 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_fill_1 FILLER_14_126 ();
 sg13g2_decap_4 FILLER_14_151 ();
 sg13g2_fill_2 FILLER_14_155 ();
 sg13g2_decap_8 FILLER_14_170 ();
 sg13g2_fill_2 FILLER_14_177 ();
 sg13g2_fill_1 FILLER_14_179 ();
 sg13g2_fill_1 FILLER_14_188 ();
 sg13g2_fill_1 FILLER_14_199 ();
 sg13g2_decap_8 FILLER_14_218 ();
 sg13g2_fill_2 FILLER_14_230 ();
 sg13g2_fill_1 FILLER_14_232 ();
 sg13g2_decap_8 FILLER_14_242 ();
 sg13g2_fill_1 FILLER_14_249 ();
 sg13g2_fill_2 FILLER_14_258 ();
 sg13g2_fill_1 FILLER_14_260 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_fill_2 FILLER_14_406 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_4 FILLER_15_49 ();
 sg13g2_fill_1 FILLER_15_53 ();
 sg13g2_fill_2 FILLER_15_97 ();
 sg13g2_fill_1 FILLER_15_99 ();
 sg13g2_decap_4 FILLER_15_124 ();
 sg13g2_fill_1 FILLER_15_128 ();
 sg13g2_decap_8 FILLER_15_142 ();
 sg13g2_fill_2 FILLER_15_149 ();
 sg13g2_decap_4 FILLER_15_175 ();
 sg13g2_decap_4 FILLER_15_201 ();
 sg13g2_fill_1 FILLER_15_205 ();
 sg13g2_decap_4 FILLER_15_210 ();
 sg13g2_fill_1 FILLER_15_214 ();
 sg13g2_fill_2 FILLER_15_237 ();
 sg13g2_fill_1 FILLER_15_239 ();
 sg13g2_decap_8 FILLER_15_267 ();
 sg13g2_decap_8 FILLER_15_274 ();
 sg13g2_decap_8 FILLER_15_281 ();
 sg13g2_decap_8 FILLER_15_288 ();
 sg13g2_fill_1 FILLER_15_295 ();
 sg13g2_decap_8 FILLER_15_301 ();
 sg13g2_decap_8 FILLER_15_308 ();
 sg13g2_decap_8 FILLER_15_315 ();
 sg13g2_decap_8 FILLER_15_322 ();
 sg13g2_decap_8 FILLER_15_329 ();
 sg13g2_decap_8 FILLER_15_336 ();
 sg13g2_decap_8 FILLER_15_343 ();
 sg13g2_decap_8 FILLER_15_350 ();
 sg13g2_decap_8 FILLER_15_357 ();
 sg13g2_decap_8 FILLER_15_364 ();
 sg13g2_decap_8 FILLER_15_371 ();
 sg13g2_decap_8 FILLER_15_378 ();
 sg13g2_decap_8 FILLER_15_385 ();
 sg13g2_decap_8 FILLER_15_392 ();
 sg13g2_decap_8 FILLER_15_399 ();
 sg13g2_fill_2 FILLER_15_406 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_fill_1 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_55 ();
 sg13g2_fill_2 FILLER_16_62 ();
 sg13g2_fill_1 FILLER_16_64 ();
 sg13g2_fill_1 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_79 ();
 sg13g2_fill_1 FILLER_16_86 ();
 sg13g2_fill_1 FILLER_16_108 ();
 sg13g2_fill_2 FILLER_16_135 ();
 sg13g2_fill_2 FILLER_16_177 ();
 sg13g2_fill_2 FILLER_16_191 ();
 sg13g2_fill_1 FILLER_16_202 ();
 sg13g2_fill_1 FILLER_16_215 ();
 sg13g2_decap_8 FILLER_16_228 ();
 sg13g2_fill_2 FILLER_16_247 ();
 sg13g2_decap_8 FILLER_16_261 ();
 sg13g2_fill_1 FILLER_16_287 ();
 sg13g2_fill_1 FILLER_16_317 ();
 sg13g2_decap_8 FILLER_16_328 ();
 sg13g2_fill_2 FILLER_16_335 ();
 sg13g2_fill_1 FILLER_16_337 ();
 sg13g2_decap_8 FILLER_16_363 ();
 sg13g2_decap_4 FILLER_16_370 ();
 sg13g2_fill_1 FILLER_16_374 ();
 sg13g2_fill_2 FILLER_16_384 ();
 sg13g2_decap_8 FILLER_16_391 ();
 sg13g2_decap_8 FILLER_16_398 ();
 sg13g2_decap_4 FILLER_16_405 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_50 ();
 sg13g2_fill_2 FILLER_17_57 ();
 sg13g2_fill_1 FILLER_17_59 ();
 sg13g2_decap_4 FILLER_17_68 ();
 sg13g2_decap_8 FILLER_17_85 ();
 sg13g2_fill_1 FILLER_17_92 ();
 sg13g2_decap_8 FILLER_17_106 ();
 sg13g2_decap_8 FILLER_17_113 ();
 sg13g2_decap_4 FILLER_17_120 ();
 sg13g2_fill_1 FILLER_17_124 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_4 FILLER_17_154 ();
 sg13g2_fill_2 FILLER_17_158 ();
 sg13g2_decap_8 FILLER_17_193 ();
 sg13g2_fill_2 FILLER_17_200 ();
 sg13g2_decap_4 FILLER_17_207 ();
 sg13g2_fill_2 FILLER_17_211 ();
 sg13g2_decap_8 FILLER_17_221 ();
 sg13g2_fill_2 FILLER_17_228 ();
 sg13g2_decap_8 FILLER_17_256 ();
 sg13g2_fill_1 FILLER_17_289 ();
 sg13g2_decap_4 FILLER_17_306 ();
 sg13g2_fill_1 FILLER_17_310 ();
 sg13g2_decap_4 FILLER_17_364 ();
 sg13g2_fill_2 FILLER_17_378 ();
 sg13g2_fill_1 FILLER_17_380 ();
 sg13g2_decap_8 FILLER_17_402 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_4 FILLER_18_35 ();
 sg13g2_fill_2 FILLER_18_46 ();
 sg13g2_fill_1 FILLER_18_48 ();
 sg13g2_decap_4 FILLER_18_75 ();
 sg13g2_fill_1 FILLER_18_87 ();
 sg13g2_fill_1 FILLER_18_109 ();
 sg13g2_fill_1 FILLER_18_169 ();
 sg13g2_fill_2 FILLER_18_204 ();
 sg13g2_fill_1 FILLER_18_214 ();
 sg13g2_fill_2 FILLER_18_241 ();
 sg13g2_decap_8 FILLER_18_248 ();
 sg13g2_decap_4 FILLER_18_255 ();
 sg13g2_fill_1 FILLER_18_259 ();
 sg13g2_decap_8 FILLER_18_279 ();
 sg13g2_fill_2 FILLER_18_286 ();
 sg13g2_decap_8 FILLER_18_308 ();
 sg13g2_fill_2 FILLER_18_315 ();
 sg13g2_decap_8 FILLER_18_330 ();
 sg13g2_decap_4 FILLER_18_337 ();
 sg13g2_decap_4 FILLER_18_356 ();
 sg13g2_fill_2 FILLER_18_360 ();
 sg13g2_decap_4 FILLER_18_382 ();
 sg13g2_decap_4 FILLER_18_405 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_4 FILLER_19_21 ();
 sg13g2_fill_1 FILLER_19_25 ();
 sg13g2_fill_2 FILLER_19_57 ();
 sg13g2_fill_1 FILLER_19_59 ();
 sg13g2_decap_8 FILLER_19_65 ();
 sg13g2_fill_1 FILLER_19_72 ();
 sg13g2_fill_1 FILLER_19_78 ();
 sg13g2_fill_2 FILLER_19_89 ();
 sg13g2_fill_1 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_122 ();
 sg13g2_fill_1 FILLER_19_137 ();
 sg13g2_decap_4 FILLER_19_143 ();
 sg13g2_fill_2 FILLER_19_147 ();
 sg13g2_decap_8 FILLER_19_168 ();
 sg13g2_fill_1 FILLER_19_175 ();
 sg13g2_decap_8 FILLER_19_184 ();
 sg13g2_fill_1 FILLER_19_191 ();
 sg13g2_fill_2 FILLER_19_222 ();
 sg13g2_decap_8 FILLER_19_229 ();
 sg13g2_fill_2 FILLER_19_236 ();
 sg13g2_decap_8 FILLER_19_248 ();
 sg13g2_decap_4 FILLER_19_255 ();
 sg13g2_fill_2 FILLER_19_259 ();
 sg13g2_fill_1 FILLER_19_266 ();
 sg13g2_decap_4 FILLER_19_288 ();
 sg13g2_fill_1 FILLER_19_306 ();
 sg13g2_fill_2 FILLER_19_317 ();
 sg13g2_fill_1 FILLER_19_319 ();
 sg13g2_fill_1 FILLER_19_342 ();
 sg13g2_decap_4 FILLER_19_354 ();
 sg13g2_decap_4 FILLER_19_374 ();
 sg13g2_decap_8 FILLER_19_402 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_fill_1 FILLER_20_47 ();
 sg13g2_decap_4 FILLER_20_69 ();
 sg13g2_fill_1 FILLER_20_81 ();
 sg13g2_fill_2 FILLER_20_90 ();
 sg13g2_fill_1 FILLER_20_92 ();
 sg13g2_fill_1 FILLER_20_101 ();
 sg13g2_fill_2 FILLER_20_118 ();
 sg13g2_fill_1 FILLER_20_120 ();
 sg13g2_decap_4 FILLER_20_154 ();
 sg13g2_decap_8 FILLER_20_166 ();
 sg13g2_fill_2 FILLER_20_173 ();
 sg13g2_decap_8 FILLER_20_198 ();
 sg13g2_decap_8 FILLER_20_205 ();
 sg13g2_fill_1 FILLER_20_212 ();
 sg13g2_decap_4 FILLER_20_226 ();
 sg13g2_fill_2 FILLER_20_258 ();
 sg13g2_fill_1 FILLER_20_260 ();
 sg13g2_decap_4 FILLER_20_274 ();
 sg13g2_fill_2 FILLER_20_278 ();
 sg13g2_fill_2 FILLER_20_284 ();
 sg13g2_fill_1 FILLER_20_286 ();
 sg13g2_fill_1 FILLER_20_321 ();
 sg13g2_decap_8 FILLER_20_330 ();
 sg13g2_fill_2 FILLER_20_344 ();
 sg13g2_fill_2 FILLER_20_351 ();
 sg13g2_fill_1 FILLER_20_353 ();
 sg13g2_decap_4 FILLER_20_364 ();
 sg13g2_fill_1 FILLER_20_379 ();
 sg13g2_fill_1 FILLER_20_392 ();
 sg13g2_decap_4 FILLER_20_404 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_4 FILLER_21_42 ();
 sg13g2_fill_1 FILLER_21_46 ();
 sg13g2_fill_2 FILLER_21_51 ();
 sg13g2_fill_1 FILLER_21_69 ();
 sg13g2_fill_2 FILLER_21_83 ();
 sg13g2_fill_1 FILLER_21_85 ();
 sg13g2_fill_2 FILLER_21_94 ();
 sg13g2_decap_8 FILLER_21_108 ();
 sg13g2_fill_1 FILLER_21_115 ();
 sg13g2_decap_8 FILLER_21_121 ();
 sg13g2_fill_1 FILLER_21_128 ();
 sg13g2_decap_8 FILLER_21_137 ();
 sg13g2_decap_4 FILLER_21_144 ();
 sg13g2_fill_1 FILLER_21_148 ();
 sg13g2_decap_8 FILLER_21_161 ();
 sg13g2_decap_8 FILLER_21_168 ();
 sg13g2_fill_2 FILLER_21_175 ();
 sg13g2_fill_1 FILLER_21_177 ();
 sg13g2_decap_8 FILLER_21_206 ();
 sg13g2_decap_8 FILLER_21_231 ();
 sg13g2_fill_2 FILLER_21_238 ();
 sg13g2_fill_1 FILLER_21_240 ();
 sg13g2_decap_8 FILLER_21_249 ();
 sg13g2_fill_2 FILLER_21_256 ();
 sg13g2_fill_1 FILLER_21_258 ();
 sg13g2_decap_8 FILLER_21_264 ();
 sg13g2_fill_1 FILLER_21_271 ();
 sg13g2_fill_2 FILLER_21_290 ();
 sg13g2_fill_2 FILLER_21_305 ();
 sg13g2_fill_1 FILLER_21_307 ();
 sg13g2_decap_4 FILLER_21_319 ();
 sg13g2_fill_1 FILLER_21_323 ();
 sg13g2_decap_8 FILLER_21_332 ();
 sg13g2_decap_4 FILLER_21_354 ();
 sg13g2_fill_2 FILLER_21_358 ();
 sg13g2_decap_8 FILLER_21_376 ();
 sg13g2_fill_1 FILLER_21_383 ();
 sg13g2_decap_4 FILLER_21_404 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_fill_2 FILLER_22_28 ();
 sg13g2_fill_1 FILLER_22_30 ();
 sg13g2_decap_4 FILLER_22_39 ();
 sg13g2_fill_2 FILLER_22_51 ();
 sg13g2_decap_4 FILLER_22_58 ();
 sg13g2_fill_1 FILLER_22_62 ();
 sg13g2_decap_8 FILLER_22_68 ();
 sg13g2_decap_8 FILLER_22_75 ();
 sg13g2_fill_1 FILLER_22_82 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_fill_2 FILLER_22_126 ();
 sg13g2_decap_4 FILLER_22_145 ();
 sg13g2_fill_1 FILLER_22_149 ();
 sg13g2_fill_2 FILLER_22_156 ();
 sg13g2_fill_2 FILLER_22_163 ();
 sg13g2_fill_1 FILLER_22_185 ();
 sg13g2_decap_8 FILLER_22_196 ();
 sg13g2_decap_8 FILLER_22_203 ();
 sg13g2_fill_2 FILLER_22_210 ();
 sg13g2_decap_8 FILLER_22_229 ();
 sg13g2_decap_4 FILLER_22_252 ();
 sg13g2_fill_2 FILLER_22_268 ();
 sg13g2_fill_2 FILLER_22_280 ();
 sg13g2_fill_1 FILLER_22_282 ();
 sg13g2_decap_4 FILLER_22_292 ();
 sg13g2_fill_2 FILLER_22_301 ();
 sg13g2_decap_4 FILLER_22_311 ();
 sg13g2_fill_1 FILLER_22_315 ();
 sg13g2_decap_4 FILLER_22_325 ();
 sg13g2_fill_2 FILLER_22_329 ();
 sg13g2_fill_2 FILLER_22_356 ();
 sg13g2_fill_1 FILLER_22_363 ();
 sg13g2_fill_1 FILLER_22_380 ();
 sg13g2_fill_2 FILLER_22_386 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_fill_1 FILLER_23_14 ();
 sg13g2_fill_2 FILLER_23_50 ();
 sg13g2_fill_1 FILLER_23_52 ();
 sg13g2_fill_2 FILLER_23_101 ();
 sg13g2_fill_1 FILLER_23_103 ();
 sg13g2_decap_8 FILLER_23_112 ();
 sg13g2_fill_2 FILLER_23_119 ();
 sg13g2_fill_2 FILLER_23_126 ();
 sg13g2_fill_1 FILLER_23_128 ();
 sg13g2_fill_1 FILLER_23_141 ();
 sg13g2_decap_8 FILLER_23_176 ();
 sg13g2_decap_4 FILLER_23_207 ();
 sg13g2_fill_2 FILLER_23_224 ();
 sg13g2_fill_1 FILLER_23_226 ();
 sg13g2_fill_2 FILLER_23_233 ();
 sg13g2_fill_1 FILLER_23_259 ();
 sg13g2_decap_4 FILLER_23_265 ();
 sg13g2_decap_4 FILLER_23_290 ();
 sg13g2_fill_1 FILLER_23_294 ();
 sg13g2_fill_2 FILLER_23_314 ();
 sg13g2_fill_1 FILLER_23_316 ();
 sg13g2_decap_8 FILLER_23_326 ();
 sg13g2_fill_2 FILLER_23_333 ();
 sg13g2_fill_1 FILLER_23_335 ();
 sg13g2_decap_4 FILLER_23_356 ();
 sg13g2_fill_2 FILLER_23_360 ();
 sg13g2_decap_8 FILLER_23_372 ();
 sg13g2_fill_1 FILLER_23_379 ();
 sg13g2_fill_2 FILLER_23_389 ();
 sg13g2_fill_1 FILLER_23_391 ();
 sg13g2_decap_4 FILLER_23_404 ();
 sg13g2_fill_1 FILLER_23_408 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_fill_2 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_45 ();
 sg13g2_fill_2 FILLER_24_52 ();
 sg13g2_decap_8 FILLER_24_81 ();
 sg13g2_decap_4 FILLER_24_88 ();
 sg13g2_fill_2 FILLER_24_92 ();
 sg13g2_fill_1 FILLER_24_102 ();
 sg13g2_decap_4 FILLER_24_113 ();
 sg13g2_fill_1 FILLER_24_117 ();
 sg13g2_fill_2 FILLER_24_133 ();
 sg13g2_fill_2 FILLER_24_151 ();
 sg13g2_fill_1 FILLER_24_153 ();
 sg13g2_decap_8 FILLER_24_157 ();
 sg13g2_fill_1 FILLER_24_169 ();
 sg13g2_fill_2 FILLER_24_175 ();
 sg13g2_fill_2 FILLER_24_186 ();
 sg13g2_decap_4 FILLER_24_195 ();
 sg13g2_fill_2 FILLER_24_210 ();
 sg13g2_fill_1 FILLER_24_212 ();
 sg13g2_decap_8 FILLER_24_238 ();
 sg13g2_decap_8 FILLER_24_257 ();
 sg13g2_decap_8 FILLER_24_264 ();
 sg13g2_decap_8 FILLER_24_271 ();
 sg13g2_fill_1 FILLER_24_306 ();
 sg13g2_fill_1 FILLER_24_317 ();
 sg13g2_fill_2 FILLER_24_347 ();
 sg13g2_fill_1 FILLER_24_349 ();
 sg13g2_decap_8 FILLER_24_381 ();
 sg13g2_fill_2 FILLER_24_388 ();
 sg13g2_fill_1 FILLER_24_390 ();
 sg13g2_decap_4 FILLER_24_403 ();
 sg13g2_fill_2 FILLER_24_407 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_40 ();
 sg13g2_decap_4 FILLER_25_47 ();
 sg13g2_fill_2 FILLER_25_77 ();
 sg13g2_fill_1 FILLER_25_79 ();
 sg13g2_decap_8 FILLER_25_97 ();
 sg13g2_decap_8 FILLER_25_114 ();
 sg13g2_fill_2 FILLER_25_121 ();
 sg13g2_decap_4 FILLER_25_131 ();
 sg13g2_fill_2 FILLER_25_135 ();
 sg13g2_decap_4 FILLER_25_152 ();
 sg13g2_fill_1 FILLER_25_156 ();
 sg13g2_fill_1 FILLER_25_222 ();
 sg13g2_decap_8 FILLER_25_232 ();
 sg13g2_fill_2 FILLER_25_268 ();
 sg13g2_decap_8 FILLER_25_278 ();
 sg13g2_decap_8 FILLER_25_285 ();
 sg13g2_fill_2 FILLER_25_292 ();
 sg13g2_fill_1 FILLER_25_294 ();
 sg13g2_fill_1 FILLER_25_300 ();
 sg13g2_decap_4 FILLER_25_310 ();
 sg13g2_fill_2 FILLER_25_314 ();
 sg13g2_decap_8 FILLER_25_326 ();
 sg13g2_decap_4 FILLER_25_355 ();
 sg13g2_fill_1 FILLER_25_363 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_4 FILLER_26_7 ();
 sg13g2_fill_1 FILLER_26_37 ();
 sg13g2_fill_2 FILLER_26_43 ();
 sg13g2_decap_8 FILLER_26_53 ();
 sg13g2_fill_2 FILLER_26_60 ();
 sg13g2_fill_1 FILLER_26_62 ();
 sg13g2_decap_8 FILLER_26_71 ();
 sg13g2_fill_2 FILLER_26_86 ();
 sg13g2_fill_2 FILLER_26_114 ();
 sg13g2_fill_1 FILLER_26_116 ();
 sg13g2_decap_4 FILLER_26_138 ();
 sg13g2_fill_2 FILLER_26_147 ();
 sg13g2_fill_1 FILLER_26_149 ();
 sg13g2_decap_4 FILLER_26_158 ();
 sg13g2_fill_2 FILLER_26_162 ();
 sg13g2_fill_2 FILLER_26_182 ();
 sg13g2_fill_1 FILLER_26_184 ();
 sg13g2_decap_4 FILLER_26_221 ();
 sg13g2_fill_1 FILLER_26_225 ();
 sg13g2_decap_8 FILLER_26_232 ();
 sg13g2_fill_1 FILLER_26_239 ();
 sg13g2_fill_2 FILLER_26_336 ();
 sg13g2_fill_2 FILLER_26_353 ();
 sg13g2_fill_1 FILLER_26_355 ();
 sg13g2_fill_2 FILLER_26_361 ();
 sg13g2_decap_8 FILLER_26_369 ();
 sg13g2_decap_8 FILLER_26_376 ();
 sg13g2_decap_8 FILLER_26_383 ();
 sg13g2_decap_4 FILLER_26_405 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_fill_2 FILLER_27_36 ();
 sg13g2_fill_1 FILLER_27_38 ();
 sg13g2_fill_2 FILLER_27_65 ();
 sg13g2_fill_1 FILLER_27_67 ();
 sg13g2_fill_2 FILLER_27_141 ();
 sg13g2_fill_1 FILLER_27_143 ();
 sg13g2_fill_2 FILLER_27_189 ();
 sg13g2_fill_1 FILLER_27_222 ();
 sg13g2_fill_1 FILLER_27_275 ();
 sg13g2_decap_8 FILLER_27_289 ();
 sg13g2_decap_4 FILLER_27_296 ();
 sg13g2_fill_2 FILLER_27_300 ();
 sg13g2_fill_2 FILLER_27_310 ();
 sg13g2_fill_1 FILLER_27_312 ();
 sg13g2_decap_8 FILLER_27_321 ();
 sg13g2_fill_2 FILLER_27_328 ();
 sg13g2_fill_2 FILLER_27_346 ();
 sg13g2_fill_1 FILLER_27_348 ();
 sg13g2_decap_8 FILLER_27_364 ();
 sg13g2_fill_1 FILLER_27_408 ();
 sg13g2_decap_4 FILLER_28_0 ();
 sg13g2_fill_1 FILLER_28_4 ();
 sg13g2_fill_2 FILLER_28_53 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_fill_2 FILLER_28_75 ();
 sg13g2_fill_2 FILLER_28_92 ();
 sg13g2_decap_8 FILLER_28_102 ();
 sg13g2_decap_8 FILLER_28_109 ();
 sg13g2_decap_8 FILLER_28_116 ();
 sg13g2_fill_2 FILLER_28_123 ();
 sg13g2_fill_1 FILLER_28_138 ();
 sg13g2_decap_8 FILLER_28_144 ();
 sg13g2_decap_8 FILLER_28_161 ();
 sg13g2_decap_4 FILLER_28_168 ();
 sg13g2_fill_2 FILLER_28_172 ();
 sg13g2_fill_2 FILLER_28_238 ();
 sg13g2_fill_1 FILLER_28_247 ();
 sg13g2_fill_1 FILLER_28_301 ();
 sg13g2_fill_1 FILLER_28_310 ();
 sg13g2_decap_8 FILLER_28_319 ();
 sg13g2_decap_4 FILLER_28_326 ();
 sg13g2_fill_1 FILLER_28_336 ();
 sg13g2_decap_4 FILLER_28_373 ();
 sg13g2_fill_2 FILLER_28_377 ();
 sg13g2_fill_1 FILLER_28_384 ();
 sg13g2_decap_4 FILLER_28_405 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_4 FILLER_29_28 ();
 sg13g2_fill_1 FILLER_29_32 ();
 sg13g2_fill_2 FILLER_29_67 ();
 sg13g2_fill_1 FILLER_29_69 ();
 sg13g2_fill_2 FILLER_29_78 ();
 sg13g2_decap_8 FILLER_29_96 ();
 sg13g2_decap_4 FILLER_29_129 ();
 sg13g2_fill_2 FILLER_29_133 ();
 sg13g2_decap_4 FILLER_29_190 ();
 sg13g2_fill_2 FILLER_29_231 ();
 sg13g2_fill_1 FILLER_29_233 ();
 sg13g2_fill_2 FILLER_29_252 ();
 sg13g2_fill_1 FILLER_29_254 ();
 sg13g2_decap_8 FILLER_29_284 ();
 sg13g2_decap_8 FILLER_29_291 ();
 sg13g2_decap_4 FILLER_29_319 ();
 sg13g2_fill_1 FILLER_29_328 ();
 sg13g2_decap_8 FILLER_29_344 ();
 sg13g2_decap_4 FILLER_29_351 ();
 sg13g2_fill_1 FILLER_29_355 ();
 sg13g2_decap_8 FILLER_29_364 ();
 sg13g2_decap_4 FILLER_29_371 ();
 sg13g2_fill_1 FILLER_29_375 ();
 sg13g2_fill_1 FILLER_29_408 ();
 sg13g2_decap_4 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_4 FILLER_30_63 ();
 sg13g2_fill_2 FILLER_30_67 ();
 sg13g2_fill_2 FILLER_30_90 ();
 sg13g2_fill_1 FILLER_30_92 ();
 sg13g2_fill_2 FILLER_30_116 ();
 sg13g2_fill_1 FILLER_30_118 ();
 sg13g2_decap_4 FILLER_30_127 ();
 sg13g2_fill_1 FILLER_30_131 ();
 sg13g2_decap_4 FILLER_30_137 ();
 sg13g2_fill_1 FILLER_30_175 ();
 sg13g2_decap_8 FILLER_30_181 ();
 sg13g2_decap_4 FILLER_30_192 ();
 sg13g2_fill_2 FILLER_30_213 ();
 sg13g2_fill_1 FILLER_30_218 ();
 sg13g2_decap_8 FILLER_30_223 ();
 sg13g2_decap_8 FILLER_30_230 ();
 sg13g2_fill_1 FILLER_30_237 ();
 sg13g2_decap_8 FILLER_30_243 ();
 sg13g2_fill_2 FILLER_30_250 ();
 sg13g2_fill_1 FILLER_30_252 ();
 sg13g2_fill_2 FILLER_30_265 ();
 sg13g2_fill_1 FILLER_30_267 ();
 sg13g2_fill_1 FILLER_30_308 ();
 sg13g2_decap_4 FILLER_30_350 ();
 sg13g2_decap_4 FILLER_30_375 ();
 sg13g2_decap_4 FILLER_30_384 ();
 sg13g2_fill_2 FILLER_30_388 ();
 sg13g2_decap_8 FILLER_30_395 ();
 sg13g2_decap_8 FILLER_30_402 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_4 FILLER_31_14 ();
 sg13g2_fill_1 FILLER_31_18 ();
 sg13g2_decap_8 FILLER_31_74 ();
 sg13g2_decap_8 FILLER_31_81 ();
 sg13g2_fill_1 FILLER_31_93 ();
 sg13g2_decap_8 FILLER_31_117 ();
 sg13g2_decap_4 FILLER_31_150 ();
 sg13g2_decap_8 FILLER_31_159 ();
 sg13g2_fill_2 FILLER_31_166 ();
 sg13g2_fill_1 FILLER_31_168 ();
 sg13g2_fill_2 FILLER_31_205 ();
 sg13g2_fill_1 FILLER_31_207 ();
 sg13g2_fill_1 FILLER_31_239 ();
 sg13g2_fill_2 FILLER_31_245 ();
 sg13g2_fill_1 FILLER_31_247 ();
 sg13g2_fill_2 FILLER_31_262 ();
 sg13g2_fill_1 FILLER_31_264 ();
 sg13g2_decap_4 FILLER_31_283 ();
 sg13g2_fill_1 FILLER_31_287 ();
 sg13g2_fill_2 FILLER_31_301 ();
 sg13g2_fill_1 FILLER_31_303 ();
 sg13g2_fill_2 FILLER_31_330 ();
 sg13g2_fill_1 FILLER_31_332 ();
 sg13g2_decap_4 FILLER_31_345 ();
 sg13g2_fill_1 FILLER_31_349 ();
 sg13g2_fill_2 FILLER_31_368 ();
 sg13g2_fill_1 FILLER_31_408 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_fill_1 FILLER_32_21 ();
 sg13g2_fill_2 FILLER_32_56 ();
 sg13g2_fill_1 FILLER_32_58 ();
 sg13g2_fill_2 FILLER_32_88 ();
 sg13g2_decap_4 FILLER_32_106 ();
 sg13g2_decap_8 FILLER_32_134 ();
 sg13g2_decap_4 FILLER_32_141 ();
 sg13g2_fill_1 FILLER_32_184 ();
 sg13g2_decap_4 FILLER_32_248 ();
 sg13g2_fill_1 FILLER_32_252 ();
 sg13g2_fill_2 FILLER_32_264 ();
 sg13g2_fill_1 FILLER_32_266 ();
 sg13g2_fill_2 FILLER_32_293 ();
 sg13g2_fill_1 FILLER_32_295 ();
 sg13g2_fill_2 FILLER_32_305 ();
 sg13g2_decap_4 FILLER_32_323 ();
 sg13g2_decap_4 FILLER_32_351 ();
 sg13g2_fill_1 FILLER_32_355 ();
 sg13g2_fill_1 FILLER_32_364 ();
 sg13g2_fill_2 FILLER_32_407 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_4 FILLER_33_49 ();
 sg13g2_fill_1 FILLER_33_53 ();
 sg13g2_decap_8 FILLER_33_73 ();
 sg13g2_fill_1 FILLER_33_80 ();
 sg13g2_fill_2 FILLER_33_113 ();
 sg13g2_fill_1 FILLER_33_115 ();
 sg13g2_fill_1 FILLER_33_121 ();
 sg13g2_decap_8 FILLER_33_127 ();
 sg13g2_decap_8 FILLER_33_134 ();
 sg13g2_fill_2 FILLER_33_141 ();
 sg13g2_fill_1 FILLER_33_143 ();
 sg13g2_decap_8 FILLER_33_148 ();
 sg13g2_fill_2 FILLER_33_164 ();
 sg13g2_fill_2 FILLER_33_205 ();
 sg13g2_fill_1 FILLER_33_212 ();
 sg13g2_decap_4 FILLER_33_218 ();
 sg13g2_fill_2 FILLER_33_222 ();
 sg13g2_fill_2 FILLER_33_229 ();
 sg13g2_fill_1 FILLER_33_231 ();
 sg13g2_decap_4 FILLER_33_256 ();
 sg13g2_fill_1 FILLER_33_260 ();
 sg13g2_decap_8 FILLER_33_291 ();
 sg13g2_fill_2 FILLER_33_345 ();
 sg13g2_fill_1 FILLER_33_347 ();
 sg13g2_decap_8 FILLER_33_353 ();
 sg13g2_fill_2 FILLER_33_360 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_4 FILLER_34_56 ();
 sg13g2_fill_1 FILLER_34_60 ();
 sg13g2_fill_2 FILLER_34_69 ();
 sg13g2_fill_1 FILLER_34_71 ();
 sg13g2_decap_4 FILLER_34_88 ();
 sg13g2_fill_2 FILLER_34_101 ();
 sg13g2_fill_1 FILLER_34_103 ();
 sg13g2_fill_2 FILLER_34_114 ();
 sg13g2_fill_1 FILLER_34_132 ();
 sg13g2_fill_2 FILLER_34_138 ();
 sg13g2_fill_1 FILLER_34_140 ();
 sg13g2_decap_4 FILLER_34_166 ();
 sg13g2_fill_2 FILLER_34_170 ();
 sg13g2_decap_4 FILLER_34_233 ();
 sg13g2_fill_2 FILLER_34_262 ();
 sg13g2_fill_1 FILLER_34_264 ();
 sg13g2_fill_2 FILLER_34_283 ();
 sg13g2_decap_4 FILLER_34_293 ();
 sg13g2_fill_2 FILLER_34_305 ();
 sg13g2_decap_8 FILLER_34_319 ();
 sg13g2_decap_8 FILLER_34_326 ();
 sg13g2_decap_8 FILLER_34_333 ();
 sg13g2_fill_1 FILLER_34_340 ();
 sg13g2_fill_2 FILLER_34_349 ();
 sg13g2_fill_1 FILLER_34_359 ();
 sg13g2_decap_8 FILLER_34_389 ();
 sg13g2_decap_8 FILLER_34_396 ();
 sg13g2_decap_4 FILLER_34_403 ();
 sg13g2_fill_2 FILLER_34_407 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_4 FILLER_35_77 ();
 sg13g2_fill_1 FILLER_35_112 ();
 sg13g2_fill_2 FILLER_35_126 ();
 sg13g2_fill_1 FILLER_35_182 ();
 sg13g2_fill_1 FILLER_35_191 ();
 sg13g2_fill_2 FILLER_35_197 ();
 sg13g2_fill_1 FILLER_35_239 ();
 sg13g2_fill_1 FILLER_35_299 ();
 sg13g2_fill_2 FILLER_35_326 ();
 sg13g2_fill_2 FILLER_35_336 ();
 sg13g2_decap_4 FILLER_35_353 ();
 sg13g2_fill_2 FILLER_35_357 ();
 sg13g2_fill_1 FILLER_35_364 ();
 sg13g2_fill_1 FILLER_35_370 ();
 sg13g2_fill_2 FILLER_35_381 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_fill_2 FILLER_36_98 ();
 sg13g2_fill_1 FILLER_36_124 ();
 sg13g2_decap_8 FILLER_36_140 ();
 sg13g2_fill_1 FILLER_36_147 ();
 sg13g2_fill_2 FILLER_36_152 ();
 sg13g2_fill_1 FILLER_36_154 ();
 sg13g2_decap_4 FILLER_36_176 ();
 sg13g2_fill_2 FILLER_36_237 ();
 sg13g2_decap_8 FILLER_36_355 ();
 sg13g2_fill_1 FILLER_36_382 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_fill_1 FILLER_37_98 ();
 sg13g2_fill_2 FILLER_37_116 ();
 sg13g2_fill_1 FILLER_37_118 ();
 sg13g2_fill_2 FILLER_37_140 ();
 sg13g2_decap_8 FILLER_37_187 ();
 sg13g2_fill_1 FILLER_37_194 ();
 sg13g2_fill_1 FILLER_37_199 ();
 sg13g2_fill_1 FILLER_37_235 ();
 sg13g2_decap_8 FILLER_37_240 ();
 sg13g2_fill_2 FILLER_37_247 ();
 sg13g2_decap_4 FILLER_37_264 ();
 sg13g2_decap_4 FILLER_37_323 ();
 sg13g2_fill_2 FILLER_37_355 ();
 sg13g2_decap_8 FILLER_37_394 ();
 sg13g2_decap_8 FILLER_37_401 ();
 sg13g2_fill_1 FILLER_37_408 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_4 FILLER_38_60 ();
 sg13g2_decap_4 FILLER_38_68 ();
 sg13g2_decap_4 FILLER_38_76 ();
 sg13g2_decap_4 FILLER_38_84 ();
 sg13g2_fill_1 FILLER_38_108 ();
 sg13g2_fill_2 FILLER_38_130 ();
 sg13g2_fill_2 FILLER_38_161 ();
 sg13g2_fill_1 FILLER_38_163 ();
 sg13g2_decap_4 FILLER_38_193 ();
 sg13g2_fill_1 FILLER_38_197 ();
 sg13g2_fill_1 FILLER_38_224 ();
 sg13g2_fill_2 FILLER_38_260 ();
 sg13g2_decap_8 FILLER_38_292 ();
 sg13g2_decap_8 FILLER_38_299 ();
 sg13g2_decap_4 FILLER_38_306 ();
 sg13g2_fill_2 FILLER_38_310 ();
 sg13g2_fill_2 FILLER_38_317 ();
 sg13g2_fill_1 FILLER_38_319 ();
 sg13g2_fill_2 FILLER_38_325 ();
 sg13g2_fill_1 FILLER_38_327 ();
 sg13g2_fill_2 FILLER_38_333 ();
 sg13g2_fill_1 FILLER_38_343 ();
 sg13g2_fill_2 FILLER_38_349 ();
 sg13g2_fill_1 FILLER_38_351 ();
 sg13g2_fill_1 FILLER_38_357 ();
 sg13g2_fill_1 FILLER_38_373 ();
 sg13g2_fill_1 FILLER_38_382 ();
 assign uio_oe[0] = net7;
 assign uio_oe[1] = net8;
 assign uio_oe[2] = net9;
 assign uio_oe[3] = net10;
 assign uio_oe[4] = net11;
 assign uio_oe[5] = net12;
 assign uio_oe[6] = net13;
 assign uio_oe[7] = net14;
 assign uio_out[0] = net15;
 assign uio_out[1] = net16;
 assign uio_out[2] = net17;
 assign uio_out[3] = net18;
 assign uio_out[4] = net19;
 assign uio_out[5] = net20;
 assign uio_out[6] = net21;
 assign uio_out[7] = net22;
endmodule

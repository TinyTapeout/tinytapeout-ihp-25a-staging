module tt_um_purdue_socet_uart (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire \uart_proj.bg.rate[0] ;
 wire \uart_proj.bg.rate[10] ;
 wire \uart_proj.bg.rate[11] ;
 wire \uart_proj.bg.rate[1] ;
 wire \uart_proj.bg.rate[2] ;
 wire \uart_proj.bg.rate[5] ;
 wire \uart_proj.bg.rate[7] ;
 wire \uart_proj.bg.rate[8] ;
 wire \uart_proj.bg.rxCount[0] ;
 wire \uart_proj.bg.rxCount[10] ;
 wire \uart_proj.bg.rxCount[11] ;
 wire \uart_proj.bg.rxCount[12] ;
 wire \uart_proj.bg.rxCount[13] ;
 wire \uart_proj.bg.rxCount[14] ;
 wire \uart_proj.bg.rxCount[15] ;
 wire \uart_proj.bg.rxCount[1] ;
 wire \uart_proj.bg.rxCount[2] ;
 wire \uart_proj.bg.rxCount[3] ;
 wire \uart_proj.bg.rxCount[4] ;
 wire \uart_proj.bg.rxCount[5] ;
 wire \uart_proj.bg.rxCount[6] ;
 wire \uart_proj.bg.rxCount[7] ;
 wire \uart_proj.bg.rxCount[8] ;
 wire \uart_proj.bg.rxCount[9] ;
 wire \uart_proj.bg.txCount[0] ;
 wire \uart_proj.bg.txCount[10] ;
 wire \uart_proj.bg.txCount[11] ;
 wire \uart_proj.bg.txCount[12] ;
 wire \uart_proj.bg.txCount[13] ;
 wire \uart_proj.bg.txCount[14] ;
 wire \uart_proj.bg.txCount[15] ;
 wire \uart_proj.bg.txCount[16] ;
 wire \uart_proj.bg.txCount[17] ;
 wire \uart_proj.bg.txCount[18] ;
 wire \uart_proj.bg.txCount[19] ;
 wire \uart_proj.bg.txCount[1] ;
 wire \uart_proj.bg.txCount[2] ;
 wire \uart_proj.bg.txCount[3] ;
 wire \uart_proj.bg.txCount[4] ;
 wire \uart_proj.bg.txCount[5] ;
 wire \uart_proj.bg.txCount[6] ;
 wire \uart_proj.bg.txCount[7] ;
 wire \uart_proj.bg.txCount[8] ;
 wire \uart_proj.bg.txCount[9] ;
 wire \uart_proj.err ;
 wire \uart_proj.fifoRx.WEN ;
 wire \uart_proj.fifoRx.count[0] ;
 wire \uart_proj.fifoRx.count[1] ;
 wire \uart_proj.fifoRx.count[2] ;
 wire \uart_proj.fifoRx.count[3] ;
 wire \uart_proj.fifoRx.count_next[0] ;
 wire \uart_proj.fifoRx.count_next[1] ;
 wire \uart_proj.fifoRx.count_next[2] ;
 wire \uart_proj.fifoRx.count_next[3] ;
 wire \uart_proj.fifoRx.empty ;
 wire \uart_proj.fifoRx.fifo[0] ;
 wire \uart_proj.fifoRx.fifo[10] ;
 wire \uart_proj.fifoRx.fifo[11] ;
 wire \uart_proj.fifoRx.fifo[12] ;
 wire \uart_proj.fifoRx.fifo[13] ;
 wire \uart_proj.fifoRx.fifo[14] ;
 wire \uart_proj.fifoRx.fifo[15] ;
 wire \uart_proj.fifoRx.fifo[16] ;
 wire \uart_proj.fifoRx.fifo[17] ;
 wire \uart_proj.fifoRx.fifo[18] ;
 wire \uart_proj.fifoRx.fifo[19] ;
 wire \uart_proj.fifoRx.fifo[1] ;
 wire \uart_proj.fifoRx.fifo[20] ;
 wire \uart_proj.fifoRx.fifo[21] ;
 wire \uart_proj.fifoRx.fifo[22] ;
 wire \uart_proj.fifoRx.fifo[23] ;
 wire \uart_proj.fifoRx.fifo[24] ;
 wire \uart_proj.fifoRx.fifo[25] ;
 wire \uart_proj.fifoRx.fifo[26] ;
 wire \uart_proj.fifoRx.fifo[27] ;
 wire \uart_proj.fifoRx.fifo[28] ;
 wire \uart_proj.fifoRx.fifo[29] ;
 wire \uart_proj.fifoRx.fifo[2] ;
 wire \uart_proj.fifoRx.fifo[30] ;
 wire \uart_proj.fifoRx.fifo[31] ;
 wire \uart_proj.fifoRx.fifo[32] ;
 wire \uart_proj.fifoRx.fifo[33] ;
 wire \uart_proj.fifoRx.fifo[34] ;
 wire \uart_proj.fifoRx.fifo[35] ;
 wire \uart_proj.fifoRx.fifo[36] ;
 wire \uart_proj.fifoRx.fifo[37] ;
 wire \uart_proj.fifoRx.fifo[38] ;
 wire \uart_proj.fifoRx.fifo[39] ;
 wire \uart_proj.fifoRx.fifo[3] ;
 wire \uart_proj.fifoRx.fifo[40] ;
 wire \uart_proj.fifoRx.fifo[41] ;
 wire \uart_proj.fifoRx.fifo[42] ;
 wire \uart_proj.fifoRx.fifo[43] ;
 wire \uart_proj.fifoRx.fifo[44] ;
 wire \uart_proj.fifoRx.fifo[45] ;
 wire \uart_proj.fifoRx.fifo[46] ;
 wire \uart_proj.fifoRx.fifo[47] ;
 wire \uart_proj.fifoRx.fifo[48] ;
 wire \uart_proj.fifoRx.fifo[49] ;
 wire \uart_proj.fifoRx.fifo[4] ;
 wire \uart_proj.fifoRx.fifo[50] ;
 wire \uart_proj.fifoRx.fifo[51] ;
 wire \uart_proj.fifoRx.fifo[52] ;
 wire \uart_proj.fifoRx.fifo[53] ;
 wire \uart_proj.fifoRx.fifo[54] ;
 wire \uart_proj.fifoRx.fifo[55] ;
 wire \uart_proj.fifoRx.fifo[56] ;
 wire \uart_proj.fifoRx.fifo[57] ;
 wire \uart_proj.fifoRx.fifo[58] ;
 wire \uart_proj.fifoRx.fifo[59] ;
 wire \uart_proj.fifoRx.fifo[5] ;
 wire \uart_proj.fifoRx.fifo[60] ;
 wire \uart_proj.fifoRx.fifo[61] ;
 wire \uart_proj.fifoRx.fifo[62] ;
 wire \uart_proj.fifoRx.fifo[63] ;
 wire \uart_proj.fifoRx.fifo[6] ;
 wire \uart_proj.fifoRx.fifo[7] ;
 wire \uart_proj.fifoRx.fifo[8] ;
 wire \uart_proj.fifoRx.fifo[9] ;
 wire \uart_proj.fifoRx.full ;
 wire \uart_proj.fifoRx.overrun ;
 wire \uart_proj.fifoRx.read_ptr[0] ;
 wire \uart_proj.fifoRx.read_ptr[1] ;
 wire \uart_proj.fifoRx.read_ptr[2] ;
 wire \uart_proj.fifoRx.wdata[0] ;
 wire \uart_proj.fifoRx.wdata[1] ;
 wire \uart_proj.fifoRx.wdata[2] ;
 wire \uart_proj.fifoRx.wdata[3] ;
 wire \uart_proj.fifoRx.wdata[4] ;
 wire \uart_proj.fifoRx.wdata[5] ;
 wire \uart_proj.fifoRx.wdata[6] ;
 wire \uart_proj.fifoRx.wdata[7] ;
 wire \uart_proj.fifoRx.write_ptr[0] ;
 wire \uart_proj.fifoRx.write_ptr[1] ;
 wire \uart_proj.fifoRx.write_ptr[2] ;
 wire \uart_proj.fifoTx.REN ;
 wire \uart_proj.fifoTx.count[0] ;
 wire \uart_proj.fifoTx.count[1] ;
 wire \uart_proj.fifoTx.count[2] ;
 wire \uart_proj.fifoTx.count[3] ;
 wire \uart_proj.fifoTx.count_next[0] ;
 wire \uart_proj.fifoTx.count_next[1] ;
 wire \uart_proj.fifoTx.count_next[2] ;
 wire \uart_proj.fifoTx.count_next[3] ;
 wire \uart_proj.fifoTx.fifo[0] ;
 wire \uart_proj.fifoTx.fifo[10] ;
 wire \uart_proj.fifoTx.fifo[11] ;
 wire \uart_proj.fifoTx.fifo[12] ;
 wire \uart_proj.fifoTx.fifo[13] ;
 wire \uart_proj.fifoTx.fifo[14] ;
 wire \uart_proj.fifoTx.fifo[15] ;
 wire \uart_proj.fifoTx.fifo[16] ;
 wire \uart_proj.fifoTx.fifo[17] ;
 wire \uart_proj.fifoTx.fifo[18] ;
 wire \uart_proj.fifoTx.fifo[19] ;
 wire \uart_proj.fifoTx.fifo[1] ;
 wire \uart_proj.fifoTx.fifo[20] ;
 wire \uart_proj.fifoTx.fifo[21] ;
 wire \uart_proj.fifoTx.fifo[22] ;
 wire \uart_proj.fifoTx.fifo[23] ;
 wire \uart_proj.fifoTx.fifo[24] ;
 wire \uart_proj.fifoTx.fifo[25] ;
 wire \uart_proj.fifoTx.fifo[26] ;
 wire \uart_proj.fifoTx.fifo[27] ;
 wire \uart_proj.fifoTx.fifo[28] ;
 wire \uart_proj.fifoTx.fifo[29] ;
 wire \uart_proj.fifoTx.fifo[2] ;
 wire \uart_proj.fifoTx.fifo[30] ;
 wire \uart_proj.fifoTx.fifo[31] ;
 wire \uart_proj.fifoTx.fifo[32] ;
 wire \uart_proj.fifoTx.fifo[33] ;
 wire \uart_proj.fifoTx.fifo[34] ;
 wire \uart_proj.fifoTx.fifo[35] ;
 wire \uart_proj.fifoTx.fifo[36] ;
 wire \uart_proj.fifoTx.fifo[37] ;
 wire \uart_proj.fifoTx.fifo[38] ;
 wire \uart_proj.fifoTx.fifo[39] ;
 wire \uart_proj.fifoTx.fifo[3] ;
 wire \uart_proj.fifoTx.fifo[40] ;
 wire \uart_proj.fifoTx.fifo[41] ;
 wire \uart_proj.fifoTx.fifo[42] ;
 wire \uart_proj.fifoTx.fifo[43] ;
 wire \uart_proj.fifoTx.fifo[44] ;
 wire \uart_proj.fifoTx.fifo[45] ;
 wire \uart_proj.fifoTx.fifo[46] ;
 wire \uart_proj.fifoTx.fifo[47] ;
 wire \uart_proj.fifoTx.fifo[48] ;
 wire \uart_proj.fifoTx.fifo[49] ;
 wire \uart_proj.fifoTx.fifo[4] ;
 wire \uart_proj.fifoTx.fifo[50] ;
 wire \uart_proj.fifoTx.fifo[51] ;
 wire \uart_proj.fifoTx.fifo[52] ;
 wire \uart_proj.fifoTx.fifo[53] ;
 wire \uart_proj.fifoTx.fifo[54] ;
 wire \uart_proj.fifoTx.fifo[55] ;
 wire \uart_proj.fifoTx.fifo[56] ;
 wire \uart_proj.fifoTx.fifo[57] ;
 wire \uart_proj.fifoTx.fifo[58] ;
 wire \uart_proj.fifoTx.fifo[59] ;
 wire \uart_proj.fifoTx.fifo[5] ;
 wire \uart_proj.fifoTx.fifo[60] ;
 wire \uart_proj.fifoTx.fifo[61] ;
 wire \uart_proj.fifoTx.fifo[62] ;
 wire \uart_proj.fifoTx.fifo[63] ;
 wire \uart_proj.fifoTx.fifo[6] ;
 wire \uart_proj.fifoTx.fifo[7] ;
 wire \uart_proj.fifoTx.fifo[8] ;
 wire \uart_proj.fifoTx.fifo[9] ;
 wire \uart_proj.fifoTx.full ;
 wire \uart_proj.fifoTx.read_ptr[0] ;
 wire \uart_proj.fifoTx.read_ptr[1] ;
 wire \uart_proj.fifoTx.read_ptr[2] ;
 wire \uart_proj.fifoTx.write_ptr[0] ;
 wire \uart_proj.fifoTx.write_ptr[1] ;
 wire \uart_proj.fifoTx.write_ptr[2] ;
 wire \uart_proj.new_rate[11] ;
 wire \uart_proj.new_rate[5] ;
 wire \uart_proj.new_rate[7] ;
 wire \uart_proj.new_rate[8] ;
 wire \uart_proj.prev_ren_wen[0] ;
 wire \uart_proj.prev_ren_wen[1] ;
 wire \uart_proj.ren_wen_nidle[0] ;
 wire \uart_proj.ren_wen_nidle[1] ;
 wire \uart_proj.rxData[0] ;
 wire \uart_proj.rxData[1] ;
 wire \uart_proj.rxData[2] ;
 wire \uart_proj.rxData[3] ;
 wire \uart_proj.rxData[4] ;
 wire \uart_proj.rxData[5] ;
 wire \uart_proj.rxData[6] ;
 wire \uart_proj.rxData[7] ;
 wire \uart_proj.tx ;
 wire \uart_proj.txData[0] ;
 wire \uart_proj.txData[1] ;
 wire \uart_proj.txData[2] ;
 wire \uart_proj.txData[3] ;
 wire \uart_proj.txData[4] ;
 wire \uart_proj.txData[5] ;
 wire \uart_proj.txData[6] ;
 wire \uart_proj.txData[7] ;
 wire \uart_proj.uartRx.cmp ;
 wire \uart_proj.uartRx.curState[0] ;
 wire \uart_proj.uartRx.curState[1] ;
 wire \uart_proj.uartRx.curState[2] ;
 wire \uart_proj.uartRx.edgeCmp ;
 wire \uart_proj.uartRx.readBuf[0] ;
 wire \uart_proj.uartRx.readBuf[1] ;
 wire \uart_proj.uartRx.readBuf[2] ;
 wire \uart_proj.uartRx.readBuf[3] ;
 wire \uart_proj.uartRx.readBuf[4] ;
 wire \uart_proj.uartRx.readBuf[5] ;
 wire \uart_proj.uartRx.readBuf[6] ;
 wire \uart_proj.uartRx.readBuf[7] ;
 wire \uart_proj.uartRx.readCount[0] ;
 wire \uart_proj.uartRx.readCount[1] ;
 wire \uart_proj.uartRx.readCount[2] ;
 wire \uart_proj.uartRx.readCount[3] ;
 wire \uart_proj.uartRx.sampleCount[0] ;
 wire \uart_proj.uartRx.sampleCount[1] ;
 wire \uart_proj.uartRx.sampleCount[2] ;
 wire \uart_proj.uartRx.sampleCount[3] ;
 wire \uart_proj.uartTx.curState[0] ;
 wire \uart_proj.uartTx.curState[1] ;
 wire \uart_proj.uartTx.curState[2] ;
 wire \uart_proj.uartTx.curState[3] ;
 wire \uart_proj.uartTx.enterStart ;
 wire \uart_proj.uartTx.hasData ;
 wire \uart_proj.uartTx.writeBuf[0] ;
 wire \uart_proj.uartTx.writeBuf[1] ;
 wire \uart_proj.uartTx.writeBuf[2] ;
 wire \uart_proj.uartTx.writeBuf[3] ;
 wire \uart_proj.uartTx.writeBuf[4] ;
 wire \uart_proj.uartTx.writeBuf[5] ;
 wire \uart_proj.uartTx.writeBuf[6] ;
 wire \uart_proj.uartTx.writeBuf[7] ;
 wire \uart_proj.uartTx.writeCount[0] ;
 wire \uart_proj.uartTx.writeCount[1] ;
 wire \uart_proj.uartTx.writeCount[2] ;
 wire \uart_proj.uartTx.writeCount[3] ;
 wire net16;
 wire net17;
 wire clknet_leaf_0_clk;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_34_clk;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;

 sg13g2_inv_1 _1373_ (.Y(_0900_),
    .A(net1));
 sg13g2_inv_2 _1374_ (.Y(_0901_),
    .A(net478));
 sg13g2_inv_2 _1375_ (.Y(_0902_),
    .A(\uart_proj.bg.rate[10] ));
 sg13g2_inv_2 _1376_ (.Y(_0903_),
    .A(net475));
 sg13g2_inv_1 _1377_ (.Y(_0904_),
    .A(net480));
 sg13g2_inv_1 _1378_ (.Y(_0905_),
    .A(\uart_proj.bg.txCount[15] ));
 sg13g2_inv_1 _1379_ (.Y(_0906_),
    .A(\uart_proj.bg.txCount[12] ));
 sg13g2_inv_1 _1380_ (.Y(_0907_),
    .A(_0112_));
 sg13g2_inv_1 _1381_ (.Y(_0908_),
    .A(\uart_proj.bg.txCount[7] ));
 sg13g2_inv_1 _1382_ (.Y(_0909_),
    .A(net546));
 sg13g2_inv_1 _1383_ (.Y(_0910_),
    .A(\uart_proj.bg.txCount[3] ));
 sg13g2_inv_1 _1384_ (.Y(_0911_),
    .A(\uart_proj.bg.txCount[1] ));
 sg13g2_inv_1 _1385_ (.Y(_0912_),
    .A(net535));
 sg13g2_inv_1 _1386_ (.Y(_0913_),
    .A(_0124_));
 sg13g2_inv_1 _1387_ (.Y(_0914_),
    .A(net215));
 sg13g2_inv_1 _1388_ (.Y(_0915_),
    .A(net349));
 sg13g2_inv_1 _1389_ (.Y(_0916_),
    .A(_0026_));
 sg13g2_inv_1 _1390_ (.Y(_0917_),
    .A(_0031_));
 sg13g2_inv_1 _1391_ (.Y(_0918_),
    .A(net236));
 sg13g2_inv_1 _1392_ (.Y(_0919_),
    .A(\uart_proj.fifoRx.count[2] ));
 sg13g2_inv_1 _1393_ (.Y(_0920_),
    .A(net536));
 sg13g2_inv_1 _1394_ (.Y(_0921_),
    .A(net20));
 sg13g2_inv_2 _1395_ (.Y(_0922_),
    .A(\uart_proj.fifoTx.read_ptr[2] ));
 sg13g2_inv_1 _1396_ (.Y(_0923_),
    .A(net473));
 sg13g2_inv_1 _1397_ (.Y(_0924_),
    .A(net545));
 sg13g2_inv_1 _1398_ (.Y(_0925_),
    .A(net2));
 sg13g2_inv_1 _1399_ (.Y(_0926_),
    .A(_0082_));
 sg13g2_or2_1 _1400_ (.X(_0161_),
    .B(net3),
    .A(net4));
 sg13g2_nor2b_1 _1401_ (.A(net4),
    .B_N(net3),
    .Y(_0160_));
 sg13g2_and2_1 _1402_ (.A(net4),
    .B(net3),
    .X(_0159_));
 sg13g2_nor2_1 _1403_ (.A(\uart_proj.bg.txCount[17] ),
    .B(\uart_proj.bg.txCount[16] ),
    .Y(_0927_));
 sg13g2_nor2_1 _1404_ (.A(\uart_proj.bg.txCount[19] ),
    .B(\uart_proj.bg.txCount[18] ),
    .Y(_0928_));
 sg13g2_or2_1 _1405_ (.X(_0929_),
    .B(\uart_proj.bg.txCount[18] ),
    .A(\uart_proj.bg.txCount[19] ));
 sg13g2_or2_1 _1406_ (.X(_0930_),
    .B(\uart_proj.bg.txCount[14] ),
    .A(\uart_proj.bg.txCount[15] ));
 sg13g2_nor3_1 _1407_ (.A(\uart_proj.bg.txCount[11] ),
    .B(\uart_proj.bg.txCount[10] ),
    .C(_0930_),
    .Y(_0931_));
 sg13g2_nand3_1 _1408_ (.B(_0928_),
    .C(_0931_),
    .A(_0927_),
    .Y(_0932_));
 sg13g2_nor4_1 _1409_ (.A(\uart_proj.bg.txCount[3] ),
    .B(\uart_proj.bg.txCount[2] ),
    .C(\uart_proj.bg.txCount[1] ),
    .D(\uart_proj.bg.txCount[0] ),
    .Y(_0933_));
 sg13g2_nor4_1 _1410_ (.A(\uart_proj.bg.txCount[7] ),
    .B(\uart_proj.bg.txCount[6] ),
    .C(\uart_proj.bg.txCount[5] ),
    .D(\uart_proj.bg.txCount[4] ),
    .Y(_0934_));
 sg13g2_nor4_2 _1411_ (.A(\uart_proj.bg.txCount[13] ),
    .B(\uart_proj.bg.txCount[12] ),
    .C(\uart_proj.bg.txCount[9] ),
    .Y(_0935_),
    .D(\uart_proj.bg.txCount[8] ));
 sg13g2_nand3_1 _1412_ (.B(_0934_),
    .C(_0935_),
    .A(_0933_),
    .Y(_0936_));
 sg13g2_nor2_1 _1413_ (.A(_0932_),
    .B(_0936_),
    .Y(_0937_));
 sg13g2_xor2_1 _1414_ (.B(\uart_proj.bg.rate[2] ),
    .A(net480),
    .X(_0938_));
 sg13g2_nor2_1 _1415_ (.A(net476),
    .B(_0904_),
    .Y(_0939_));
 sg13g2_nand2b_1 _1416_ (.Y(_0940_),
    .B(net481),
    .A_N(net476));
 sg13g2_nor3_1 _1417_ (.A(net475),
    .B(\uart_proj.bg.rate[8] ),
    .C(\uart_proj.bg.rate[7] ),
    .Y(_0941_));
 sg13g2_nor3_1 _1418_ (.A(\uart_proj.bg.rate[0] ),
    .B(\uart_proj.bg.rate[10] ),
    .C(net479),
    .Y(_0942_));
 sg13g2_nand2_2 _1419_ (.Y(_0943_),
    .A(_0941_),
    .B(_0942_));
 sg13g2_nor3_1 _1420_ (.A(_0938_),
    .B(_0939_),
    .C(_0943_),
    .Y(_0944_));
 sg13g2_nor3_2 _1421_ (.A(_0932_),
    .B(_0936_),
    .C(_0944_),
    .Y(_0945_));
 sg13g2_nand2b_2 _1422_ (.Y(_0946_),
    .B(net428),
    .A_N(_0944_));
 sg13g2_nor2_1 _1423_ (.A(\uart_proj.uartTx.curState[3] ),
    .B(net18),
    .Y(_0947_));
 sg13g2_and2_1 _1424_ (.A(net329),
    .B(_0945_),
    .X(_0948_));
 sg13g2_nor2_1 _1425_ (.A(_0947_),
    .B(_0948_),
    .Y(_0949_));
 sg13g2_o21ai_1 _1426_ (.B1(_0949_),
    .Y(_0158_),
    .A1(net18),
    .A2(_0945_));
 sg13g2_nand2_1 _1427_ (.Y(_0950_),
    .A(_0901_),
    .B(net428));
 sg13g2_o21ai_1 _1428_ (.B1(_0950_),
    .Y(_0126_),
    .A1(_0912_),
    .A2(net428));
 sg13g2_and2_1 _1429_ (.A(net351),
    .B(_0946_),
    .X(_0951_));
 sg13g2_nor3_2 _1430_ (.A(\uart_proj.uartTx.writeCount[0] ),
    .B(net280),
    .C(net282),
    .Y(_0952_));
 sg13g2_nand2b_2 _1431_ (.Y(_0953_),
    .B(_0952_),
    .A_N(\uart_proj.uartTx.writeCount[3] ));
 sg13g2_nor2_1 _1432_ (.A(_0946_),
    .B(_0953_),
    .Y(_0954_));
 sg13g2_a21o_1 _1433_ (.A2(_0954_),
    .A1(net335),
    .B1(_0951_),
    .X(_0002_));
 sg13g2_nand2b_1 _1434_ (.Y(_0955_),
    .B(_0948_),
    .A_N(_0947_));
 sg13g2_o21ai_1 _1435_ (.B1(_0955_),
    .Y(_0001_),
    .A1(net41),
    .A2(_0945_));
 sg13g2_a21oi_1 _1436_ (.A1(\uart_proj.uartTx.curState[2] ),
    .A2(_0945_),
    .Y(_0956_),
    .B1(net335));
 sg13g2_nor3_1 _1437_ (.A(\uart_proj.uartTx.curState[2] ),
    .B(_0946_),
    .C(_0953_),
    .Y(_0957_));
 sg13g2_nor2_1 _1438_ (.A(net336),
    .B(_0957_),
    .Y(_0000_));
 sg13g2_a21oi_1 _1439_ (.A1(net347),
    .A2(_0946_),
    .Y(_0958_),
    .B1(_0002_));
 sg13g2_nand2_1 _1440_ (.Y(_0024_),
    .A(_0955_),
    .B(_0958_));
 sg13g2_nand2b_1 _1441_ (.Y(_0025_),
    .B(net336),
    .A_N(_0951_));
 sg13g2_nor3_1 _1442_ (.A(\uart_proj.fifoTx.count[1] ),
    .B(\uart_proj.fifoTx.count[0] ),
    .C(\uart_proj.fifoTx.count[2] ),
    .Y(_0959_));
 sg13g2_or3_1 _1443_ (.A(\uart_proj.fifoTx.count[1] ),
    .B(\uart_proj.fifoTx.count[0] ),
    .C(\uart_proj.fifoTx.count[2] ),
    .X(_0960_));
 sg13g2_nand2_2 _1444_ (.Y(_0961_),
    .A(\uart_proj.fifoTx.count[3] ),
    .B(_0959_));
 sg13g2_inv_1 _1445_ (.Y(\uart_proj.fifoTx.full ),
    .A(_0961_));
 sg13g2_nor3_2 _1446_ (.A(\uart_proj.fifoRx.count[1] ),
    .B(\uart_proj.fifoRx.count[0] ),
    .C(\uart_proj.fifoRx.count[2] ),
    .Y(_0962_));
 sg13g2_nand2_2 _1447_ (.Y(_0963_),
    .A(net398),
    .B(_0962_));
 sg13g2_inv_1 _1448_ (.Y(\uart_proj.fifoRx.full ),
    .A(_0963_));
 sg13g2_nor2b_1 _1449_ (.A(\uart_proj.fifoRx.count[3] ),
    .B_N(_0962_),
    .Y(\uart_proj.fifoRx.empty ));
 sg13g2_nor2b_2 _1450_ (.A(net5),
    .B_N(net6),
    .Y(uio_oe[7]));
 sg13g2_nand3_1 _1451_ (.B(net480),
    .C(\uart_proj.bg.rate[2] ),
    .A(net476),
    .Y(_0964_));
 sg13g2_nand2_1 _1452_ (.Y(_0965_),
    .A(net475),
    .B(_0964_));
 sg13g2_xor2_1 _1453_ (.B(_0965_),
    .A(_0121_),
    .X(_0966_));
 sg13g2_and2_1 _1454_ (.A(_0910_),
    .B(_0966_),
    .X(_0967_));
 sg13g2_xnor2_1 _1455_ (.Y(_0968_),
    .A(net478),
    .B(_0117_));
 sg13g2_nor2_1 _1456_ (.A(_0116_),
    .B(\uart_proj.bg.txCount[7] ),
    .Y(_0969_));
 sg13g2_and2_1 _1457_ (.A(_0116_),
    .B(\uart_proj.bg.txCount[7] ),
    .X(_0970_));
 sg13g2_nor3_1 _1458_ (.A(_0968_),
    .B(_0969_),
    .C(_0970_),
    .Y(_0971_));
 sg13g2_xnor2_1 _1459_ (.Y(_0972_),
    .A(_0118_),
    .B(_0119_));
 sg13g2_nor2_1 _1460_ (.A(net480),
    .B(_0120_),
    .Y(_0973_));
 sg13g2_xor2_1 _1461_ (.B(_0120_),
    .A(net480),
    .X(_0974_));
 sg13g2_nand3_1 _1462_ (.B(_0972_),
    .C(_0974_),
    .A(_0971_),
    .Y(_0975_));
 sg13g2_mux2_2 _1463_ (.A0(\uart_proj.bg.rate[2] ),
    .A1(_0938_),
    .S(_0940_),
    .X(_0976_));
 sg13g2_xnor2_1 _1464_ (.Y(_0977_),
    .A(_0903_),
    .B(_0964_));
 sg13g2_xor2_1 _1465_ (.B(_0977_),
    .A(_0122_),
    .X(_0978_));
 sg13g2_a21oi_1 _1466_ (.A1(_0911_),
    .A2(_0976_),
    .Y(_0979_),
    .B1(_0978_));
 sg13g2_nand2b_1 _1467_ (.Y(_0980_),
    .B(\uart_proj.bg.txCount[1] ),
    .A_N(_0976_));
 sg13g2_xnor2_1 _1468_ (.Y(_0981_),
    .A(net476),
    .B(net481));
 sg13g2_nand3b_1 _1469_ (.B(_0123_),
    .C(_0980_),
    .Y(_0982_),
    .A_N(_0981_));
 sg13g2_nor2_1 _1470_ (.A(_0910_),
    .B(_0966_),
    .Y(_0983_));
 sg13g2_a221oi_1 _1471_ (.B2(_0982_),
    .C1(_0983_),
    .B1(_0979_),
    .A1(\uart_proj.bg.txCount[2] ),
    .Y(_0984_),
    .A2(_0977_));
 sg13g2_nor3_1 _1472_ (.A(_0967_),
    .B(_0975_),
    .C(_0984_),
    .Y(_0985_));
 sg13g2_a21oi_1 _1473_ (.A1(_0901_),
    .A2(\uart_proj.bg.txCount[6] ),
    .Y(_0986_),
    .B1(_0970_));
 sg13g2_a22oi_1 _1474_ (.Y(_0987_),
    .B1(_0972_),
    .B2(_0973_),
    .A2(\uart_proj.bg.txCount[5] ),
    .A1(_0118_));
 sg13g2_inv_1 _1475_ (.Y(_0988_),
    .A(_0987_));
 sg13g2_a21oi_1 _1476_ (.A1(_0971_),
    .A2(_0988_),
    .Y(_0989_),
    .B1(_0985_));
 sg13g2_o21ai_1 _1477_ (.B1(_0989_),
    .Y(_0990_),
    .A1(_0969_),
    .A2(_0986_));
 sg13g2_xor2_1 _1478_ (.B(_0114_),
    .A(_0115_),
    .X(_0991_));
 sg13g2_nor2_1 _1479_ (.A(\uart_proj.bg.txCount[14] ),
    .B(\uart_proj.bg.txCount[13] ),
    .Y(_0992_));
 sg13g2_nor2_1 _1480_ (.A(net478),
    .B(_0906_),
    .Y(_0993_));
 sg13g2_a22oi_1 _1481_ (.Y(_0994_),
    .B1(_0111_),
    .B2(net474),
    .A2(_0906_),
    .A1(net478));
 sg13g2_nor2_1 _1482_ (.A(net474),
    .B(_0111_),
    .Y(_0995_));
 sg13g2_xnor2_1 _1483_ (.Y(_0996_),
    .A(\uart_proj.bg.rate[10] ),
    .B(\uart_proj.bg.txCount[10] ));
 sg13g2_nand3b_1 _1484_ (.B(_0927_),
    .C(_0105_),
    .Y(_0997_),
    .A_N(\uart_proj.bg.txCount[18] ));
 sg13g2_xnor2_1 _1485_ (.Y(_0998_),
    .A(net474),
    .B(\uart_proj.bg.txCount[9] ));
 sg13g2_nand2_1 _1486_ (.Y(_0999_),
    .A(_0105_),
    .B(_0106_));
 sg13g2_nand2b_1 _1487_ (.Y(_1000_),
    .B(\uart_proj.bg.txCount[16] ),
    .A_N(\uart_proj.bg.txCount[17] ));
 sg13g2_a21oi_1 _1488_ (.A1(_0107_),
    .A2(_1000_),
    .Y(_1001_),
    .B1(\uart_proj.bg.txCount[18] ));
 sg13g2_nand3b_1 _1489_ (.B(_0998_),
    .C(_0115_),
    .Y(_1002_),
    .A_N(_0114_));
 sg13g2_o21ai_1 _1490_ (.B1(_1002_),
    .Y(_1003_),
    .A1(net474),
    .A2(_0113_));
 sg13g2_a221oi_1 _1491_ (.B2(_1003_),
    .C1(_0995_),
    .B1(_0996_),
    .A1(_0902_),
    .Y(_1004_),
    .A2(_0907_));
 sg13g2_nor2b_1 _1492_ (.A(_1004_),
    .B_N(_0994_),
    .Y(_1005_));
 sg13g2_o21ai_1 _1493_ (.B1(_0992_),
    .Y(_1006_),
    .A1(_0993_),
    .A2(_1005_));
 sg13g2_or2_1 _1494_ (.X(_1007_),
    .B(_0110_),
    .A(\uart_proj.bg.txCount[14] ));
 sg13g2_nand4_1 _1495_ (.B(_0109_),
    .C(_1006_),
    .A(_0108_),
    .Y(_1008_),
    .D(_1007_));
 sg13g2_nand3_1 _1496_ (.B(_0992_),
    .C(_0998_),
    .A(_0108_),
    .Y(_1009_));
 sg13g2_nor4_1 _1497_ (.A(_0991_),
    .B(_0993_),
    .C(_0995_),
    .D(_1009_),
    .Y(_1010_));
 sg13g2_and3_1 _1498_ (.X(_1011_),
    .A(_0994_),
    .B(_0996_),
    .C(_1010_));
 sg13g2_a21oi_1 _1499_ (.A1(_0990_),
    .A2(_1011_),
    .Y(_1012_),
    .B1(_1008_));
 sg13g2_nor2_1 _1500_ (.A(_0997_),
    .B(_1012_),
    .Y(_1013_));
 sg13g2_nor3_1 _1501_ (.A(_0999_),
    .B(_1001_),
    .C(_1013_),
    .Y(_1014_));
 sg13g2_xnor2_1 _1502_ (.Y(_1015_),
    .A(\uart_proj.bg.txCount[0] ),
    .B(_0981_));
 sg13g2_nor3_1 _1503_ (.A(_0975_),
    .B(_0997_),
    .C(_1015_),
    .Y(_1016_));
 sg13g2_nand3_1 _1504_ (.B(_1011_),
    .C(_1016_),
    .A(_0980_),
    .Y(_1017_));
 sg13g2_nor3_1 _1505_ (.A(_0967_),
    .B(_0983_),
    .C(_1017_),
    .Y(_1018_));
 sg13g2_a21oi_2 _1506_ (.B1(_1014_),
    .Y(_1019_),
    .A2(_1018_),
    .A1(_0979_));
 sg13g2_inv_1 _1507_ (.Y(_1020_),
    .A(_1019_));
 sg13g2_nor3_1 _1508_ (.A(net477),
    .B(net479),
    .C(net481),
    .Y(_1021_));
 sg13g2_nor2b_1 _1509_ (.A(\uart_proj.bg.rate[7] ),
    .B_N(_1021_),
    .Y(_1022_));
 sg13g2_nand2b_2 _1510_ (.Y(_1023_),
    .B(_1022_),
    .A_N(\uart_proj.bg.rate[8] ));
 sg13g2_xnor2_1 _1511_ (.Y(_1024_),
    .A(_0903_),
    .B(_1023_));
 sg13g2_xnor2_1 _1512_ (.Y(_1025_),
    .A(\uart_proj.bg.rate[8] ),
    .B(_1022_));
 sg13g2_mux2_1 _1513_ (.A0(_0121_),
    .A1(_1025_),
    .S(_0965_),
    .X(_1026_));
 sg13g2_inv_1 _1514_ (.Y(_1027_),
    .A(_1026_));
 sg13g2_nand2_1 _1515_ (.Y(_1028_),
    .A(_1024_),
    .B(_1027_));
 sg13g2_xnor2_1 _1516_ (.Y(_1029_),
    .A(\uart_proj.bg.rate[7] ),
    .B(_1021_));
 sg13g2_nor2b_1 _1517_ (.A(_1029_),
    .B_N(_0977_),
    .Y(_1030_));
 sg13g2_xnor2_1 _1518_ (.Y(_1031_),
    .A(_0977_),
    .B(_1029_));
 sg13g2_a21oi_1 _1519_ (.A1(\uart_proj.bg.rate[2] ),
    .A2(_1031_),
    .Y(_1032_),
    .B1(_1030_));
 sg13g2_nor2b_1 _1520_ (.A(net475),
    .B_N(_0121_),
    .Y(_1033_));
 sg13g2_a21oi_1 _1521_ (.A1(net475),
    .A2(_0966_),
    .Y(_1034_),
    .B1(_1033_));
 sg13g2_xnor2_1 _1522_ (.Y(_1035_),
    .A(_1025_),
    .B(_1034_));
 sg13g2_nor2_1 _1523_ (.A(_1032_),
    .B(_1035_),
    .Y(_1036_));
 sg13g2_nand2b_1 _1524_ (.Y(_1037_),
    .B(net479),
    .A_N(net476));
 sg13g2_o21ai_1 _1525_ (.B1(_1037_),
    .Y(_1038_),
    .A1(net479),
    .A2(_0981_));
 sg13g2_nor2_1 _1526_ (.A(_0976_),
    .B(_1038_),
    .Y(_1039_));
 sg13g2_xor2_1 _1527_ (.B(_1038_),
    .A(_0976_),
    .X(_1040_));
 sg13g2_a21o_1 _1528_ (.A2(_1040_),
    .A1(net477),
    .B1(_1039_),
    .X(_1041_));
 sg13g2_xnor2_1 _1529_ (.Y(_1042_),
    .A(\uart_proj.bg.rate[2] ),
    .B(_1031_));
 sg13g2_nand2b_1 _1530_ (.Y(_1043_),
    .B(_1041_),
    .A_N(_1042_));
 sg13g2_or2_1 _1531_ (.X(_1044_),
    .B(_1040_),
    .A(net476));
 sg13g2_nand3_1 _1532_ (.B(net479),
    .C(_0904_),
    .A(net476),
    .Y(_1045_));
 sg13g2_o21ai_1 _1533_ (.B1(_1045_),
    .Y(_1046_),
    .A1(net479),
    .A2(_0940_));
 sg13g2_a21oi_1 _1534_ (.A1(net476),
    .A2(_1040_),
    .Y(_1047_),
    .B1(_1046_));
 sg13g2_and2_1 _1535_ (.A(_1044_),
    .B(_1047_),
    .X(_1048_));
 sg13g2_a21oi_1 _1536_ (.A1(\uart_proj.bg.rate[2] ),
    .A2(_1046_),
    .Y(_1049_),
    .B1(_1048_));
 sg13g2_a221oi_1 _1537_ (.B2(_1044_),
    .C1(_0904_),
    .B1(_1047_),
    .A1(\uart_proj.bg.rate[2] ),
    .Y(_1050_),
    .A2(_1046_));
 sg13g2_xnor2_1 _1538_ (.Y(_1051_),
    .A(_1041_),
    .B(_1042_));
 sg13g2_o21ai_1 _1539_ (.B1(_1051_),
    .Y(_1052_),
    .A1(_1048_),
    .A2(_1050_));
 sg13g2_xnor2_1 _1540_ (.Y(_1053_),
    .A(_1032_),
    .B(_1035_));
 sg13g2_a21oi_1 _1541_ (.A1(_1043_),
    .A2(_1052_),
    .Y(_1054_),
    .B1(_1053_));
 sg13g2_nor2_1 _1542_ (.A(_1036_),
    .B(_1054_),
    .Y(_1055_));
 sg13g2_xor2_1 _1543_ (.B(_1026_),
    .A(_1024_),
    .X(_1056_));
 sg13g2_inv_1 _1544_ (.Y(_1057_),
    .A(_1056_));
 sg13g2_o21ai_1 _1545_ (.B1(_1057_),
    .Y(_1058_),
    .A1(_1036_),
    .A2(_1054_));
 sg13g2_nand2_1 _1546_ (.Y(_1059_),
    .A(_1028_),
    .B(_1058_));
 sg13g2_nand2_1 _1547_ (.Y(_1060_),
    .A(_0902_),
    .B(net474));
 sg13g2_nor2_1 _1548_ (.A(\uart_proj.bg.rate[10] ),
    .B(_1023_),
    .Y(_1061_));
 sg13g2_nor2_2 _1549_ (.A(net475),
    .B(_1061_),
    .Y(_1062_));
 sg13g2_nand2_1 _1550_ (.Y(_1063_),
    .A(\uart_proj.bg.rate[10] ),
    .B(_1023_));
 sg13g2_a22oi_1 _1551_ (.Y(_1064_),
    .B1(_1062_),
    .B2(_1063_),
    .A2(net474),
    .A1(_0902_));
 sg13g2_xnor2_1 _1552_ (.Y(_1065_),
    .A(\uart_proj.bg.rate[5] ),
    .B(_0118_));
 sg13g2_xnor2_1 _1553_ (.Y(_1066_),
    .A(_1064_),
    .B(_1065_));
 sg13g2_nand2b_1 _1554_ (.Y(_1067_),
    .B(_1066_),
    .A_N(_1024_));
 sg13g2_nand2b_1 _1555_ (.Y(_1068_),
    .B(_1024_),
    .A_N(_1066_));
 sg13g2_nand2_1 _1556_ (.Y(_1069_),
    .A(_1067_),
    .B(_1068_));
 sg13g2_xor2_1 _1557_ (.B(_1069_),
    .A(_1059_),
    .X(_1070_));
 sg13g2_nand2_1 _1558_ (.Y(_1071_),
    .A(\uart_proj.bg.txCount[5] ),
    .B(_1070_));
 sg13g2_xnor2_1 _1559_ (.Y(_1072_),
    .A(_1055_),
    .B(_1057_));
 sg13g2_nand2_1 _1560_ (.Y(_1073_),
    .A(_0120_),
    .B(_1072_));
 sg13g2_nand3_1 _1561_ (.B(_1052_),
    .C(_1053_),
    .A(_1043_),
    .Y(_1074_));
 sg13g2_nand2b_1 _1562_ (.Y(_1075_),
    .B(_1074_),
    .A_N(_1054_));
 sg13g2_nor2_1 _1563_ (.A(\uart_proj.bg.txCount[3] ),
    .B(_1075_),
    .Y(_1076_));
 sg13g2_or3_1 _1564_ (.A(_1048_),
    .B(_1050_),
    .C(_1051_),
    .X(_1077_));
 sg13g2_nand2_1 _1565_ (.Y(_1078_),
    .A(_1052_),
    .B(_1077_));
 sg13g2_xnor2_1 _1566_ (.Y(_1079_),
    .A(net477),
    .B(net479));
 sg13g2_nand3_1 _1567_ (.B(_0123_),
    .C(_1079_),
    .A(_0911_),
    .Y(_1080_));
 sg13g2_a21oi_1 _1568_ (.A1(_0123_),
    .A2(_1079_),
    .Y(_1081_),
    .B1(_0911_));
 sg13g2_xnor2_1 _1569_ (.Y(_1082_),
    .A(net480),
    .B(_1049_));
 sg13g2_a21o_1 _1570_ (.A2(_1082_),
    .A1(_1080_),
    .B1(_1081_),
    .X(_1083_));
 sg13g2_xnor2_1 _1571_ (.Y(_1084_),
    .A(_0122_),
    .B(_1078_));
 sg13g2_a22oi_1 _1572_ (.Y(_1085_),
    .B1(_1083_),
    .B2(_1084_),
    .A2(_1078_),
    .A1(\uart_proj.bg.txCount[2] ));
 sg13g2_nor2_1 _1573_ (.A(_0120_),
    .B(_1072_),
    .Y(_1086_));
 sg13g2_nand2_1 _1574_ (.Y(_1087_),
    .A(\uart_proj.bg.txCount[3] ),
    .B(_1075_));
 sg13g2_o21ai_1 _1575_ (.B1(_1087_),
    .Y(_1088_),
    .A1(_1076_),
    .A2(_1085_));
 sg13g2_a21oi_1 _1576_ (.A1(_1073_),
    .A2(_1088_),
    .Y(_1089_),
    .B1(_1086_));
 sg13g2_xor2_1 _1577_ (.B(_1070_),
    .A(_0119_),
    .X(_1090_));
 sg13g2_o21ai_1 _1578_ (.B1(_1071_),
    .Y(_1091_),
    .A1(_1089_),
    .A2(_1090_));
 sg13g2_nand3_1 _1579_ (.B(_0903_),
    .C(_1023_),
    .A(\uart_proj.bg.rate[10] ),
    .Y(_1092_));
 sg13g2_nand2_1 _1580_ (.Y(_1093_),
    .A(_1060_),
    .B(_1092_));
 sg13g2_nand3_1 _1581_ (.B(_1058_),
    .C(_1067_),
    .A(_1028_),
    .Y(_1094_));
 sg13g2_nand2_1 _1582_ (.Y(_1095_),
    .A(_1068_),
    .B(_1094_));
 sg13g2_nand4_1 _1583_ (.B(_1068_),
    .C(_1092_),
    .A(_1060_),
    .Y(_1096_),
    .D(_1094_));
 sg13g2_xor2_1 _1584_ (.B(_1095_),
    .A(_1093_),
    .X(_1097_));
 sg13g2_xnor2_1 _1585_ (.Y(_1098_),
    .A(_0909_),
    .B(_1097_));
 sg13g2_nor2_2 _1586_ (.A(net481),
    .B(_0943_),
    .Y(_1099_));
 sg13g2_nor2_1 _1587_ (.A(net478),
    .B(_1099_),
    .Y(_1100_));
 sg13g2_xnor2_1 _1588_ (.Y(_1101_),
    .A(\uart_proj.bg.rate[7] ),
    .B(_0116_));
 sg13g2_xnor2_1 _1589_ (.Y(_1102_),
    .A(_1100_),
    .B(_1101_));
 sg13g2_xnor2_1 _1590_ (.Y(_1103_),
    .A(_1062_),
    .B(_1102_));
 sg13g2_xor2_1 _1591_ (.B(_1102_),
    .A(_1062_),
    .X(_1104_));
 sg13g2_a21oi_1 _1592_ (.A1(_1092_),
    .A2(_1096_),
    .Y(_1105_),
    .B1(_1104_));
 sg13g2_and3_1 _1593_ (.X(_1106_),
    .A(_1092_),
    .B(_1096_),
    .C(_1104_));
 sg13g2_nor2_1 _1594_ (.A(_1105_),
    .B(_1106_),
    .Y(_1107_));
 sg13g2_nor2b_1 _1595_ (.A(_1097_),
    .B_N(\uart_proj.bg.txCount[6] ),
    .Y(_1108_));
 sg13g2_a221oi_1 _1596_ (.B2(\uart_proj.bg.txCount[7] ),
    .C1(_1108_),
    .B1(_1107_),
    .A1(_1091_),
    .Y(_1109_),
    .A2(_1098_));
 sg13g2_a21o_1 _1597_ (.A2(_1063_),
    .A1(_1062_),
    .B1(_1102_),
    .X(_1110_));
 sg13g2_o21ai_1 _1598_ (.B1(_1110_),
    .Y(_1111_),
    .A1(_1096_),
    .A2(_1103_));
 sg13g2_xnor2_1 _1599_ (.Y(_1112_),
    .A(\uart_proj.bg.rate[8] ),
    .B(_0115_));
 sg13g2_xnor2_1 _1600_ (.Y(_1113_),
    .A(net478),
    .B(_1112_));
 sg13g2_xnor2_1 _1601_ (.Y(_1114_),
    .A(_1111_),
    .B(_1113_));
 sg13g2_o21ai_1 _1602_ (.B1(_0908_),
    .Y(_1115_),
    .A1(_1105_),
    .A2(_1106_));
 sg13g2_o21ai_1 _1603_ (.B1(_1115_),
    .Y(_1116_),
    .A1(\uart_proj.bg.txCount[8] ),
    .A2(_1114_));
 sg13g2_nand2_1 _1604_ (.Y(_1117_),
    .A(\uart_proj.bg.txCount[8] ),
    .B(_1114_));
 sg13g2_o21ai_1 _1605_ (.B1(_1117_),
    .Y(_1118_),
    .A1(_1109_),
    .A2(_1116_));
 sg13g2_nand2_1 _1606_ (.Y(_1119_),
    .A(_1099_),
    .B(_1112_));
 sg13g2_o21ai_1 _1607_ (.B1(_1119_),
    .Y(_1120_),
    .A1(_0901_),
    .A2(_1112_));
 sg13g2_a21oi_2 _1608_ (.B1(_1120_),
    .Y(_1121_),
    .A2(_1113_),
    .A1(_1111_));
 sg13g2_nor2_1 _1609_ (.A(_0113_),
    .B(_1121_),
    .Y(_1122_));
 sg13g2_nor2_1 _1610_ (.A(\uart_proj.bg.txCount[11] ),
    .B(_0907_),
    .Y(_1123_));
 sg13g2_nand2b_1 _1611_ (.Y(_1124_),
    .B(_1123_),
    .A_N(_1121_));
 sg13g2_nand3b_1 _1612_ (.B(\uart_proj.bg.txCount[11] ),
    .C(_0907_),
    .Y(_1125_),
    .A_N(_0113_));
 sg13g2_a21oi_1 _1613_ (.A1(_1124_),
    .A2(_1125_),
    .Y(_1126_),
    .B1(_1122_));
 sg13g2_nand3b_1 _1614_ (.B(_1123_),
    .C(\uart_proj.bg.txCount[9] ),
    .Y(_1127_),
    .A_N(_1121_));
 sg13g2_a21oi_1 _1615_ (.A1(_0109_),
    .A2(\uart_proj.bg.txCount[13] ),
    .Y(_1128_),
    .B1(_0930_));
 sg13g2_nand2_1 _1616_ (.Y(_1129_),
    .A(_0109_),
    .B(_0110_));
 sg13g2_o21ai_1 _1617_ (.B1(_1128_),
    .Y(_1130_),
    .A1(_0125_),
    .A2(_1129_));
 sg13g2_nor3_1 _1618_ (.A(\uart_proj.bg.txCount[11] ),
    .B(\uart_proj.bg.txCount[10] ),
    .C(_1130_),
    .Y(_1131_));
 sg13g2_a21oi_1 _1619_ (.A1(_1127_),
    .A2(_1131_),
    .Y(_1132_),
    .B1(_1121_));
 sg13g2_a21o_1 _1620_ (.A2(_1126_),
    .A1(_1118_),
    .B1(_1132_),
    .X(_1133_));
 sg13g2_a221oi_1 _1621_ (.B2(_1113_),
    .C1(_1120_),
    .B1(_1111_),
    .A1(_0903_),
    .Y(_1134_),
    .A2(_1061_));
 sg13g2_xnor2_1 _1622_ (.Y(_1135_),
    .A(_0107_),
    .B(_1134_));
 sg13g2_nor4_1 _1623_ (.A(_0905_),
    .B(_0109_),
    .C(_0110_),
    .D(_0125_),
    .Y(_1136_));
 sg13g2_a21oi_1 _1624_ (.A1(_1128_),
    .A2(_1129_),
    .Y(_1137_),
    .B1(_1121_));
 sg13g2_a21oi_1 _1625_ (.A1(_1121_),
    .A2(_1136_),
    .Y(_1138_),
    .B1(_1137_));
 sg13g2_xnor2_1 _1626_ (.Y(_1139_),
    .A(_1099_),
    .B(_1121_));
 sg13g2_and2_1 _1627_ (.A(_0913_),
    .B(_1139_),
    .X(_1140_));
 sg13g2_nor2b_1 _1628_ (.A(_0106_),
    .B_N(\uart_proj.bg.txCount[19] ),
    .Y(_1141_));
 sg13g2_nor2b_1 _1629_ (.A(\uart_proj.bg.txCount[19] ),
    .B_N(_0106_),
    .Y(_1142_));
 sg13g2_mux2_1 _1630_ (.A0(_1142_),
    .A1(_1141_),
    .S(_1134_),
    .X(_1143_));
 sg13g2_o21ai_1 _1631_ (.B1(_1143_),
    .Y(_1144_),
    .A1(_0913_),
    .A2(_1139_));
 sg13g2_nor4_2 _1632_ (.A(_1135_),
    .B(_1138_),
    .C(_1140_),
    .Y(_1145_),
    .D(_1144_));
 sg13g2_a21oi_1 _1633_ (.A1(\uart_proj.bg.txCount[17] ),
    .A2(_1143_),
    .Y(_1146_),
    .B1(_0929_));
 sg13g2_nand4_1 _1634_ (.B(_0913_),
    .C(_1139_),
    .A(_0107_),
    .Y(_1147_),
    .D(_1143_));
 sg13g2_o21ai_1 _1635_ (.B1(_1147_),
    .Y(_1148_),
    .A1(_1134_),
    .A2(_1146_));
 sg13g2_a21oi_2 _1636_ (.B1(_1148_),
    .Y(_1149_),
    .A2(_1145_),
    .A1(_1133_));
 sg13g2_a21o_1 _1637_ (.A2(_1145_),
    .A1(_1133_),
    .B1(_1148_),
    .X(_1150_));
 sg13g2_nor4_1 _1638_ (.A(\uart_proj.bg.rxCount[3] ),
    .B(\uart_proj.bg.rxCount[2] ),
    .C(\uart_proj.bg.rxCount[5] ),
    .D(\uart_proj.bg.rxCount[4] ),
    .Y(_1151_));
 sg13g2_nor4_1 _1639_ (.A(\uart_proj.bg.rxCount[13] ),
    .B(\uart_proj.bg.rxCount[12] ),
    .C(\uart_proj.bg.rxCount[15] ),
    .D(\uart_proj.bg.rxCount[14] ),
    .Y(_1152_));
 sg13g2_nor4_1 _1640_ (.A(\uart_proj.bg.rxCount[7] ),
    .B(\uart_proj.bg.rxCount[6] ),
    .C(\uart_proj.bg.rxCount[11] ),
    .D(\uart_proj.bg.rxCount[10] ),
    .Y(_1153_));
 sg13g2_nor4_1 _1641_ (.A(\uart_proj.bg.rxCount[1] ),
    .B(\uart_proj.bg.rxCount[0] ),
    .C(\uart_proj.bg.rxCount[9] ),
    .D(\uart_proj.bg.rxCount[8] ),
    .Y(_1154_));
 sg13g2_and4_1 _1642_ (.A(_1151_),
    .B(_1152_),
    .C(_1153_),
    .D(_1154_),
    .X(_1155_));
 sg13g2_and2_1 _1643_ (.A(_0943_),
    .B(net432),
    .X(_1156_));
 sg13g2_nand2_1 _1644_ (.Y(_1157_),
    .A(_0943_),
    .B(net431));
 sg13g2_nor3_2 _1645_ (.A(_1019_),
    .B(_1149_),
    .C(_1157_),
    .Y(_1158_));
 sg13g2_inv_2 _1646_ (.Y(_1159_),
    .A(_1158_));
 sg13g2_nor2b_1 _1647_ (.A(net1),
    .B_N(\uart_proj.uartRx.cmp ),
    .Y(_1160_));
 sg13g2_xnor2_1 _1648_ (.Y(_1161_),
    .A(net1),
    .B(\uart_proj.uartRx.cmp ));
 sg13g2_nor4_2 _1649_ (.A(_1019_),
    .B(_1149_),
    .C(_1157_),
    .Y(_1162_),
    .D(_1161_));
 sg13g2_nand2b_1 _1650_ (.Y(_1163_),
    .B(net406),
    .A_N(_1161_));
 sg13g2_and2_1 _1651_ (.A(\uart_proj.uartRx.sampleCount[3] ),
    .B(\uart_proj.uartRx.edgeCmp ),
    .X(_1164_));
 sg13g2_nor2_1 _1652_ (.A(\uart_proj.uartRx.sampleCount[0] ),
    .B(\uart_proj.uartRx.sampleCount[1] ),
    .Y(_1165_));
 sg13g2_nor3_2 _1653_ (.A(\uart_proj.uartRx.sampleCount[0] ),
    .B(\uart_proj.uartRx.sampleCount[1] ),
    .C(\uart_proj.uartRx.sampleCount[2] ),
    .Y(_1166_));
 sg13g2_nand2b_2 _1654_ (.Y(_1167_),
    .B(_1165_),
    .A_N(\uart_proj.uartRx.sampleCount[2] ));
 sg13g2_a21oi_2 _1655_ (.B1(\uart_proj.uartRx.sampleCount[3] ),
    .Y(_1168_),
    .A2(_1167_),
    .A1(_1161_));
 sg13g2_nand4_1 _1656_ (.B(_1150_),
    .C(_1156_),
    .A(_1020_),
    .Y(_1169_),
    .D(_1168_));
 sg13g2_a22oi_1 _1657_ (.Y(_1170_),
    .B1(_1169_),
    .B2(\uart_proj.uartRx.curState[0] ),
    .A2(_1164_),
    .A1(_1162_));
 sg13g2_nor2_1 _1658_ (.A(\uart_proj.uartRx.curState[1] ),
    .B(\uart_proj.uartRx.curState[0] ),
    .Y(_1171_));
 sg13g2_o21ai_1 _1659_ (.B1(_0029_),
    .Y(_1172_),
    .A1(\uart_proj.uartRx.curState[1] ),
    .A2(\uart_proj.uartRx.curState[0] ));
 sg13g2_nand2_1 _1660_ (.Y(_1173_),
    .A(\uart_proj.uartRx.curState[2] ),
    .B(_1171_));
 sg13g2_a21oi_1 _1661_ (.A1(_1172_),
    .A2(_1173_),
    .Y(_1174_),
    .B1(_1170_));
 sg13g2_nand2_1 _1662_ (.Y(_1175_),
    .A(\uart_proj.uartRx.sampleCount[3] ),
    .B(_1166_));
 sg13g2_nand3_1 _1663_ (.B(net406),
    .C(_1166_),
    .A(\uart_proj.uartRx.sampleCount[3] ),
    .Y(_1176_));
 sg13g2_nand4_1 _1664_ (.B(\uart_proj.uartRx.sampleCount[3] ),
    .C(net406),
    .A(_0900_),
    .Y(_1177_),
    .D(_1166_));
 sg13g2_nand3b_1 _1665_ (.B(net406),
    .C(_1160_),
    .Y(_1178_),
    .A_N(\uart_proj.uartRx.sampleCount[3] ));
 sg13g2_a21oi_1 _1666_ (.A1(_1177_),
    .A2(_1178_),
    .Y(_1179_),
    .B1(_1173_));
 sg13g2_nor3_2 _1667_ (.A(net241),
    .B(\uart_proj.uartRx.readCount[1] ),
    .C(net21),
    .Y(_1180_));
 sg13g2_nor2b_2 _1668_ (.A(\uart_proj.uartRx.readCount[3] ),
    .B_N(_1180_),
    .Y(_1181_));
 sg13g2_and2_1 _1669_ (.A(\uart_proj.uartRx.curState[1] ),
    .B(_0029_),
    .X(_1182_));
 sg13g2_nand2_1 _1670_ (.Y(_1183_),
    .A(\uart_proj.uartRx.curState[1] ),
    .B(_0029_));
 sg13g2_nor4_1 _1671_ (.A(\uart_proj.uartRx.curState[0] ),
    .B(_1169_),
    .C(_1181_),
    .D(_1183_),
    .Y(_1184_));
 sg13g2_nand2_1 _1672_ (.Y(_1185_),
    .A(_0029_),
    .B(_1171_));
 sg13g2_and3_1 _1673_ (.X(_1186_),
    .A(_0029_),
    .B(_1160_),
    .C(_1171_));
 sg13g2_nor4_2 _1674_ (.A(_1174_),
    .B(_1179_),
    .C(_1184_),
    .Y(_1187_),
    .D(_1186_));
 sg13g2_nand3b_1 _1675_ (.B(\uart_proj.uartRx.curState[0] ),
    .C(_0029_),
    .Y(_1188_),
    .A_N(\uart_proj.uartRx.curState[1] ));
 sg13g2_and2_1 _1676_ (.A(net406),
    .B(_1181_),
    .X(_1189_));
 sg13g2_nand2_1 _1677_ (.Y(_1190_),
    .A(_1168_),
    .B(net403));
 sg13g2_nand4_1 _1678_ (.B(_1168_),
    .C(_1181_),
    .A(net407),
    .Y(_1191_),
    .D(_1188_));
 sg13g2_a221oi_1 _1679_ (.B2(net331),
    .C1(_1172_),
    .B1(_1169_),
    .A1(_1162_),
    .Y(_1192_),
    .A2(_1164_));
 sg13g2_nor3_1 _1680_ (.A(net331),
    .B(_1160_),
    .C(_1185_),
    .Y(_1193_));
 sg13g2_a21oi_2 _1681_ (.B1(net332),
    .Y(_1194_),
    .A2(_1192_),
    .A1(_1191_));
 sg13g2_a22oi_1 _1682_ (.Y(_1195_),
    .B1(_1169_),
    .B2(\uart_proj.uartRx.curState[2] ),
    .A2(_1164_),
    .A1(_1162_));
 sg13g2_nand4_1 _1683_ (.B(_1168_),
    .C(_1181_),
    .A(net406),
    .Y(_1196_),
    .D(_1182_));
 sg13g2_o21ai_1 _1684_ (.B1(_1196_),
    .Y(_1197_),
    .A1(_1172_),
    .A2(_1195_));
 sg13g2_a21oi_2 _1685_ (.B1(_1173_),
    .Y(_1198_),
    .A2(_1195_),
    .A1(_1177_));
 sg13g2_or2_1 _1686_ (.X(_1199_),
    .B(_1198_),
    .A(_1197_));
 sg13g2_nand3b_1 _1687_ (.B(_1194_),
    .C(_1199_),
    .Y(_1200_),
    .A_N(_1187_));
 sg13g2_nand2b_1 _1688_ (.Y(_0003_),
    .B(_1200_),
    .A_N(net88));
 sg13g2_and2_2 _1689_ (.A(net445),
    .B(net444),
    .X(_1201_));
 sg13g2_nand2_1 _1690_ (.Y(_1202_),
    .A(net445),
    .B(net444));
 sg13g2_nor2b_1 _1691_ (.A(\uart_proj.ren_wen_nidle[1] ),
    .B_N(\uart_proj.ren_wen_nidle[0] ),
    .Y(_1203_));
 sg13g2_nand2b_2 _1692_ (.Y(_1204_),
    .B(net445),
    .A_N(net444));
 sg13g2_xnor2_1 _1693_ (.Y(_1205_),
    .A(_0033_),
    .B(net441));
 sg13g2_nor2_2 _1694_ (.A(\uart_proj.fifoTx.count[3] ),
    .B(_0960_),
    .Y(_1206_));
 sg13g2_nand2_1 _1695_ (.Y(_1207_),
    .A(\uart_proj.fifoTx.REN ),
    .B(net441));
 sg13g2_mux2_1 _1696_ (.A0(_0031_),
    .A1(_1207_),
    .S(_1206_),
    .X(_1208_));
 sg13g2_nor2_2 _1697_ (.A(_1205_),
    .B(_1208_),
    .Y(_1209_));
 sg13g2_xnor2_1 _1698_ (.Y(_1210_),
    .A(_1205_),
    .B(_1208_));
 sg13g2_nor2_1 _1699_ (.A(net371),
    .B(_0961_),
    .Y(_1211_));
 sg13g2_a22oi_1 _1700_ (.Y(_1212_),
    .B1(net372),
    .B2(_1204_),
    .A2(_1210_),
    .A1(_0961_));
 sg13g2_nor2_1 _1701_ (.A(_1201_),
    .B(_1212_),
    .Y(\uart_proj.fifoTx.count_next[0] ));
 sg13g2_nor3_2 _1702_ (.A(_0033_),
    .B(_0034_),
    .C(_1204_),
    .Y(_1213_));
 sg13g2_o21ai_1 _1703_ (.B1(_0034_),
    .Y(_1214_),
    .A1(_0033_),
    .A2(_1204_));
 sg13g2_nand2b_1 _1704_ (.Y(_1215_),
    .B(_1214_),
    .A_N(_1213_));
 sg13g2_o21ai_1 _1705_ (.B1(_0961_),
    .Y(_1216_),
    .A1(_1209_),
    .A2(_1215_));
 sg13g2_a21oi_1 _1706_ (.A1(_1209_),
    .A2(_1215_),
    .Y(_1217_),
    .B1(_1216_));
 sg13g2_nand2_1 _1707_ (.Y(_0363_),
    .A(net554),
    .B(_1204_));
 sg13g2_a21oi_1 _1708_ (.A1(\uart_proj.fifoTx.REN ),
    .A2(_1204_),
    .Y(_0364_),
    .B1(net536));
 sg13g2_o21ai_1 _1709_ (.B1(\uart_proj.fifoTx.full ),
    .Y(_0365_),
    .A1(_0920_),
    .A2(_0363_));
 sg13g2_o21ai_1 _1710_ (.B1(_1202_),
    .Y(_0366_),
    .A1(_0364_),
    .A2(_0365_));
 sg13g2_nor2_1 _1711_ (.A(_1217_),
    .B(_0366_),
    .Y(\uart_proj.fifoTx.count_next[1] ));
 sg13g2_nor2_1 _1712_ (.A(_0961_),
    .B(_0363_),
    .Y(_0367_));
 sg13g2_nand2_1 _1713_ (.Y(_0368_),
    .A(\uart_proj.fifoTx.count[2] ),
    .B(_1213_));
 sg13g2_xnor2_1 _1714_ (.Y(_0369_),
    .A(\uart_proj.fifoTx.count[2] ),
    .B(_1213_));
 sg13g2_a21oi_1 _1715_ (.A1(_1209_),
    .A2(_1215_),
    .Y(_0370_),
    .B1(_0369_));
 sg13g2_nand3_1 _1716_ (.B(_1215_),
    .C(_0369_),
    .A(_1209_),
    .Y(_0371_));
 sg13g2_nand2b_1 _1717_ (.Y(_0372_),
    .B(_0371_),
    .A_N(_0370_));
 sg13g2_a21oi_1 _1718_ (.A1(_0961_),
    .A2(_0372_),
    .Y(_0373_),
    .B1(_0367_));
 sg13g2_nor2_1 _1719_ (.A(_1201_),
    .B(_0373_),
    .Y(\uart_proj.fifoTx.count_next[2] ));
 sg13g2_xor2_1 _1720_ (.B(_0368_),
    .A(\uart_proj.fifoTx.count[3] ),
    .X(_0374_));
 sg13g2_xnor2_1 _1721_ (.Y(_0375_),
    .A(_0371_),
    .B(_0374_));
 sg13g2_a221oi_1 _1722_ (.B2(_0375_),
    .C1(_0367_),
    .B1(_0961_),
    .A1(net445),
    .Y(\uart_proj.fifoTx.count_next[3] ),
    .A2(net444));
 sg13g2_nand2_1 _1723_ (.Y(_0376_),
    .A(\uart_proj.fifoRx.count[0] ),
    .B(\uart_proj.fifoRx.WEN ));
 sg13g2_xnor2_1 _1724_ (.Y(_0377_),
    .A(net532),
    .B(\uart_proj.fifoRx.WEN ));
 sg13g2_nor2b_2 _1725_ (.A(net445),
    .B_N(net444),
    .Y(_0378_));
 sg13g2_nand2b_1 _1726_ (.Y(_0379_),
    .B(net444),
    .A_N(net445));
 sg13g2_a21oi_1 _1727_ (.A1(net230),
    .A2(\uart_proj.fifoRx.empty ),
    .Y(_0380_),
    .B1(_0379_));
 sg13g2_nand2_1 _1728_ (.Y(_0381_),
    .A(net533),
    .B(_0380_));
 sg13g2_nor2_1 _1729_ (.A(_1201_),
    .B(_0377_),
    .Y(_0382_));
 sg13g2_o21ai_1 _1730_ (.B1(_0382_),
    .Y(_0383_),
    .A1(net444),
    .A2(_0963_));
 sg13g2_o21ai_1 _1731_ (.B1(_0381_),
    .Y(\uart_proj.fifoRx.count_next[0] ),
    .A1(_0380_),
    .A2(_0383_));
 sg13g2_or2_1 _1732_ (.X(_0384_),
    .B(_0376_),
    .A(_0038_));
 sg13g2_xor2_1 _1733_ (.B(_0376_),
    .A(net370),
    .X(_0385_));
 sg13g2_or2_1 _1734_ (.X(_0386_),
    .B(_0385_),
    .A(_0381_));
 sg13g2_a21oi_1 _1735_ (.A1(_0381_),
    .A2(_0385_),
    .Y(_0387_),
    .B1(\uart_proj.fifoRx.full ));
 sg13g2_nand2_1 _1736_ (.Y(_0388_),
    .A(net230),
    .B(net440));
 sg13g2_xnor2_1 _1737_ (.Y(_0389_),
    .A(net370),
    .B(_0388_));
 sg13g2_a221oi_1 _1738_ (.B2(\uart_proj.fifoRx.full ),
    .C1(_1201_),
    .B1(_0389_),
    .A1(_0386_),
    .Y(\uart_proj.fifoRx.count_next[1] ),
    .A2(_0387_));
 sg13g2_nor2_1 _1739_ (.A(net399),
    .B(_0388_),
    .Y(_0390_));
 sg13g2_or2_1 _1740_ (.X(_0391_),
    .B(_0384_),
    .A(_0919_));
 sg13g2_xnor2_1 _1741_ (.Y(_0392_),
    .A(\uart_proj.fifoRx.count[2] ),
    .B(_0384_));
 sg13g2_nor2_1 _1742_ (.A(_0386_),
    .B(_0392_),
    .Y(_0393_));
 sg13g2_xnor2_1 _1743_ (.Y(_0394_),
    .A(_0386_),
    .B(_0392_));
 sg13g2_a21oi_1 _1744_ (.A1(_0963_),
    .A2(_0394_),
    .Y(_0395_),
    .B1(_0390_));
 sg13g2_nor2_1 _1745_ (.A(_1201_),
    .B(_0395_),
    .Y(\uart_proj.fifoRx.count_next[2] ));
 sg13g2_xnor2_1 _1746_ (.Y(_0396_),
    .A(\uart_proj.fifoRx.count[3] ),
    .B(_0391_));
 sg13g2_xnor2_1 _1747_ (.Y(_0397_),
    .A(_0393_),
    .B(_0396_));
 sg13g2_a221oi_1 _1748_ (.B2(_0397_),
    .C1(_0390_),
    .B1(net399),
    .A1(net445),
    .Y(\uart_proj.fifoRx.count_next[3] ),
    .A2(net444));
 sg13g2_nand2b_1 _1749_ (.Y(_0398_),
    .B(_0030_),
    .A_N(\uart_proj.uartTx.curState[1] ));
 sg13g2_nor2_1 _1750_ (.A(\uart_proj.uartTx.curState[3] ),
    .B(_0398_),
    .Y(_0399_));
 sg13g2_nor3_1 _1751_ (.A(\uart_proj.uartTx.curState[3] ),
    .B(\uart_proj.uartTx.enterStart ),
    .C(_0398_),
    .Y(_0400_));
 sg13g2_nand3b_1 _1752_ (.B(_0953_),
    .C(_0030_),
    .Y(_0401_),
    .A_N(_0027_));
 sg13g2_a22oi_1 _1753_ (.Y(_0402_),
    .B1(_0401_),
    .B2(_0398_),
    .A2(_0400_),
    .A1(_0027_));
 sg13g2_nand2_1 _1754_ (.Y(_0403_),
    .A(_0916_),
    .B(_0953_));
 sg13g2_a221oi_1 _1755_ (.B2(\uart_proj.uartTx.curState[1] ),
    .C1(_0399_),
    .B1(_0403_),
    .A1(\uart_proj.uartTx.curState[3] ),
    .Y(_0404_),
    .A2(\uart_proj.uartTx.enterStart ));
 sg13g2_a21oi_2 _1756_ (.B1(_0404_),
    .Y(_0405_),
    .A2(_0400_),
    .A1(_0916_));
 sg13g2_nand2_1 _1757_ (.Y(_0406_),
    .A(_0402_),
    .B(_0405_));
 sg13g2_nor2_1 _1758_ (.A(_0402_),
    .B(_0405_),
    .Y(_0407_));
 sg13g2_nor3_1 _1759_ (.A(\uart_proj.uartTx.writeBuf[0] ),
    .B(_0402_),
    .C(_0405_),
    .Y(_0408_));
 sg13g2_a21oi_1 _1760_ (.A1(_0402_),
    .A2(_0405_),
    .Y(\uart_proj.tx ),
    .B1(_0408_));
 sg13g2_nor2_1 _1761_ (.A(\uart_proj.prev_ren_wen[1] ),
    .B(net297),
    .Y(_0409_));
 sg13g2_and2_1 _1762_ (.A(net5),
    .B(net298),
    .X(_0014_));
 sg13g2_and2_1 _1763_ (.A(net6),
    .B(net298),
    .X(_0015_));
 sg13g2_nor2_1 _1764_ (.A(net135),
    .B(_1190_),
    .Y(_0004_));
 sg13g2_and2_1 _1765_ (.A(net34),
    .B(net402),
    .X(_0005_));
 sg13g2_and2_1 _1766_ (.A(net68),
    .B(net402),
    .X(_0006_));
 sg13g2_and2_1 _1767_ (.A(net39),
    .B(net402),
    .X(_0007_));
 sg13g2_and2_1 _1768_ (.A(net24),
    .B(net402),
    .X(_0008_));
 sg13g2_and2_1 _1769_ (.A(net26),
    .B(net402),
    .X(_0009_));
 sg13g2_and2_1 _1770_ (.A(net28),
    .B(net402),
    .X(_0010_));
 sg13g2_and2_1 _1771_ (.A(net30),
    .B(net402),
    .X(_0011_));
 sg13g2_and2_1 _1772_ (.A(net32),
    .B(net402),
    .X(_0012_));
 sg13g2_nor3_1 _1773_ (.A(_0925_),
    .B(_0946_),
    .C(_1206_),
    .Y(_0410_));
 sg13g2_nand3b_1 _1774_ (.B(_0410_),
    .C(_0402_),
    .Y(_0411_),
    .A_N(_0405_));
 sg13g2_inv_1 _1775_ (.Y(_0013_),
    .A(_0411_));
 sg13g2_nand2b_1 _1776_ (.Y(_0412_),
    .B(net468),
    .A_N(_0046_));
 sg13g2_o21ai_1 _1777_ (.B1(_0412_),
    .Y(_0413_),
    .A1(net467),
    .A2(_0045_));
 sg13g2_nor2b_1 _1778_ (.A(net469),
    .B_N(net466),
    .Y(_0414_));
 sg13g2_and2_1 _1779_ (.A(net469),
    .B(net464),
    .X(_0415_));
 sg13g2_a221oi_1 _1780_ (.B2(_0048_),
    .C1(_0922_),
    .B1(net437),
    .A1(_0047_),
    .Y(_0416_),
    .A2(net438));
 sg13g2_o21ai_1 _1781_ (.B1(_0416_),
    .Y(_0417_),
    .A1(net465),
    .A2(_0413_));
 sg13g2_nand2b_1 _1782_ (.Y(_0418_),
    .B(net470),
    .A_N(_0042_));
 sg13g2_o21ai_1 _1783_ (.B1(_0418_),
    .Y(_0419_),
    .A1(net470),
    .A2(_0041_));
 sg13g2_a221oi_1 _1784_ (.B2(_0044_),
    .C1(\uart_proj.fifoTx.read_ptr[2] ),
    .B1(_0415_),
    .A1(net359),
    .Y(_0420_),
    .A2(net439));
 sg13g2_o21ai_1 _1785_ (.B1(net360),
    .Y(_0421_),
    .A1(net464),
    .A2(_0419_));
 sg13g2_a21oi_1 _1786_ (.A1(_0417_),
    .A2(net361),
    .Y(_0016_),
    .B1(net411));
 sg13g2_nand2b_1 _1787_ (.Y(_0422_),
    .B(net468),
    .A_N(_0054_));
 sg13g2_o21ai_1 _1788_ (.B1(_0422_),
    .Y(_0423_),
    .A1(net467),
    .A2(_0053_));
 sg13g2_a221oi_1 _1789_ (.B2(_0056_),
    .C1(_0922_),
    .B1(net437),
    .A1(_0055_),
    .Y(_0424_),
    .A2(net438));
 sg13g2_o21ai_1 _1790_ (.B1(_0424_),
    .Y(_0425_),
    .A1(net465),
    .A2(_0423_));
 sg13g2_nand2b_1 _1791_ (.Y(_0426_),
    .B(net470),
    .A_N(_0050_));
 sg13g2_o21ai_1 _1792_ (.B1(_0426_),
    .Y(_0427_),
    .A1(net470),
    .A2(_0049_));
 sg13g2_a221oi_1 _1793_ (.B2(_0052_),
    .C1(\uart_proj.fifoTx.read_ptr[2] ),
    .B1(_0415_),
    .A1(net365),
    .Y(_0428_),
    .A2(net439));
 sg13g2_o21ai_1 _1794_ (.B1(net366),
    .Y(_0429_),
    .A1(net466),
    .A2(_0427_));
 sg13g2_a21oi_1 _1795_ (.A1(_0425_),
    .A2(net367),
    .Y(_0017_),
    .B1(net411));
 sg13g2_nand2b_1 _1796_ (.Y(_0430_),
    .B(net467),
    .A_N(_0062_));
 sg13g2_o21ai_1 _1797_ (.B1(_0430_),
    .Y(_0431_),
    .A1(net467),
    .A2(_0061_));
 sg13g2_a221oi_1 _1798_ (.B2(_0064_),
    .C1(_0922_),
    .B1(net437),
    .A1(_0063_),
    .Y(_0432_),
    .A2(net438));
 sg13g2_o21ai_1 _1799_ (.B1(_0432_),
    .Y(_0433_),
    .A1(net465),
    .A2(_0431_));
 sg13g2_nand2b_1 _1800_ (.Y(_0434_),
    .B(net469),
    .A_N(_0058_));
 sg13g2_o21ai_1 _1801_ (.B1(_0434_),
    .Y(_0435_),
    .A1(net469),
    .A2(_0057_));
 sg13g2_a221oi_1 _1802_ (.B2(net387),
    .C1(net463),
    .B1(net436),
    .A1(_0059_),
    .Y(_0436_),
    .A2(net439));
 sg13g2_o21ai_1 _1803_ (.B1(net388),
    .Y(_0437_),
    .A1(net466),
    .A2(_0435_));
 sg13g2_a21oi_1 _1804_ (.A1(_0433_),
    .A2(net389),
    .Y(_0018_),
    .B1(net411));
 sg13g2_nand2b_1 _1805_ (.Y(_0438_),
    .B(net469),
    .A_N(_0066_));
 sg13g2_o21ai_1 _1806_ (.B1(_0438_),
    .Y(_0439_),
    .A1(net469),
    .A2(_0065_));
 sg13g2_a221oi_1 _1807_ (.B2(_0068_),
    .C1(net463),
    .B1(net436),
    .A1(net378),
    .Y(_0440_),
    .A2(net439));
 sg13g2_o21ai_1 _1808_ (.B1(net379),
    .Y(_0441_),
    .A1(net464),
    .A2(_0439_));
 sg13g2_nand2b_1 _1809_ (.Y(_0442_),
    .B(net467),
    .A_N(_0070_));
 sg13g2_o21ai_1 _1810_ (.B1(_0442_),
    .Y(_0443_),
    .A1(net467),
    .A2(_0069_));
 sg13g2_a221oi_1 _1811_ (.B2(_0072_),
    .C1(_0922_),
    .B1(net437),
    .A1(_0071_),
    .Y(_0444_),
    .A2(net438));
 sg13g2_o21ai_1 _1812_ (.B1(_0444_),
    .Y(_0445_),
    .A1(net465),
    .A2(_0443_));
 sg13g2_a21oi_1 _1813_ (.A1(net380),
    .A2(_0445_),
    .Y(_0019_),
    .B1(net411));
 sg13g2_nand2b_1 _1814_ (.Y(_0446_),
    .B(net469),
    .A_N(_0074_));
 sg13g2_o21ai_1 _1815_ (.B1(_0446_),
    .Y(_0447_),
    .A1(net469),
    .A2(_0073_));
 sg13g2_a221oi_1 _1816_ (.B2(_0076_),
    .C1(net463),
    .B1(net436),
    .A1(net392),
    .Y(_0448_),
    .A2(net439));
 sg13g2_o21ai_1 _1817_ (.B1(net393),
    .Y(_0449_),
    .A1(net464),
    .A2(_0447_));
 sg13g2_nand2b_1 _1818_ (.Y(_0450_),
    .B(net467),
    .A_N(_0078_));
 sg13g2_o21ai_1 _1819_ (.B1(_0450_),
    .Y(_0451_),
    .A1(net467),
    .A2(_0077_));
 sg13g2_a221oi_1 _1820_ (.B2(_0080_),
    .C1(_0922_),
    .B1(net437),
    .A1(_0079_),
    .Y(_0452_),
    .A2(net438));
 sg13g2_o21ai_1 _1821_ (.B1(_0452_),
    .Y(_0453_),
    .A1(net465),
    .A2(_0451_));
 sg13g2_a21oi_1 _1822_ (.A1(net394),
    .A2(_0453_),
    .Y(_0020_),
    .B1(net411));
 sg13g2_nand2b_1 _1823_ (.Y(_0454_),
    .B(net468),
    .A_N(_0086_));
 sg13g2_o21ai_1 _1824_ (.B1(_0454_),
    .Y(_0455_),
    .A1(net468),
    .A2(_0085_));
 sg13g2_a22oi_1 _1825_ (.Y(_0456_),
    .B1(net437),
    .B2(_0088_),
    .A2(net438),
    .A1(_0087_));
 sg13g2_o21ai_1 _1826_ (.B1(_0456_),
    .Y(_0457_),
    .A1(net465),
    .A2(_0455_));
 sg13g2_a21oi_1 _1827_ (.A1(net471),
    .A2(_0926_),
    .Y(_0458_),
    .B1(net464));
 sg13g2_o21ai_1 _1828_ (.B1(_0458_),
    .Y(_0459_),
    .A1(net471),
    .A2(net547));
 sg13g2_a22oi_1 _1829_ (.Y(_0460_),
    .B1(net436),
    .B2(_0084_),
    .A2(net439),
    .A1(_0083_));
 sg13g2_a21oi_1 _1830_ (.A1(_0459_),
    .A2(_0460_),
    .Y(_0461_),
    .B1(net463));
 sg13g2_a21oi_1 _1831_ (.A1(net463),
    .A2(_0457_),
    .Y(_0462_),
    .B1(net548));
 sg13g2_nor2b_1 _1832_ (.A(net411),
    .B_N(_0462_),
    .Y(_0021_));
 sg13g2_nand2b_1 _1833_ (.Y(_0463_),
    .B(net471),
    .A_N(_0090_));
 sg13g2_o21ai_1 _1834_ (.B1(_0463_),
    .Y(_0464_),
    .A1(net471),
    .A2(_0089_));
 sg13g2_a221oi_1 _1835_ (.B2(_0092_),
    .C1(net463),
    .B1(net436),
    .A1(net355),
    .Y(_0465_),
    .A2(net439));
 sg13g2_o21ai_1 _1836_ (.B1(net356),
    .Y(_0466_),
    .A1(net464),
    .A2(_0464_));
 sg13g2_nand2b_1 _1837_ (.Y(_0467_),
    .B(net468),
    .A_N(_0094_));
 sg13g2_o21ai_1 _1838_ (.B1(_0467_),
    .Y(_0468_),
    .A1(net468),
    .A2(_0093_));
 sg13g2_a221oi_1 _1839_ (.B2(_0096_),
    .C1(_0922_),
    .B1(net437),
    .A1(_0095_),
    .Y(_0469_),
    .A2(net438));
 sg13g2_o21ai_1 _1840_ (.B1(_0469_),
    .Y(_0470_),
    .A1(net465),
    .A2(_0468_));
 sg13g2_a21oi_1 _1841_ (.A1(net357),
    .A2(_0470_),
    .Y(_0022_),
    .B1(net411));
 sg13g2_nand2b_1 _1842_ (.Y(_0471_),
    .B(net468),
    .A_N(_0102_));
 sg13g2_o21ai_1 _1843_ (.B1(_0471_),
    .Y(_0472_),
    .A1(net468),
    .A2(_0101_));
 sg13g2_a221oi_1 _1844_ (.B2(_0104_),
    .C1(_0922_),
    .B1(net437),
    .A1(_0103_),
    .Y(_0473_),
    .A2(net438));
 sg13g2_o21ai_1 _1845_ (.B1(_0473_),
    .Y(_0474_),
    .A1(net465),
    .A2(_0472_));
 sg13g2_nand2b_1 _1846_ (.Y(_0475_),
    .B(net471),
    .A_N(_0098_));
 sg13g2_o21ai_1 _1847_ (.B1(_0475_),
    .Y(_0476_),
    .A1(net471),
    .A2(_0097_));
 sg13g2_a221oi_1 _1848_ (.B2(_0100_),
    .C1(net463),
    .B1(net436),
    .A1(net373),
    .Y(_0477_),
    .A2(net439));
 sg13g2_o21ai_1 _1849_ (.B1(net374),
    .Y(_0478_),
    .A1(net464),
    .A2(_0476_));
 sg13g2_a21oi_1 _1850_ (.A1(_0474_),
    .A2(net375),
    .Y(_0023_),
    .B1(net411));
 sg13g2_mux4_1 _1851_ (.S0(net456),
    .A0(\uart_proj.fifoRx.fifo[0] ),
    .A1(\uart_proj.fifoRx.fifo[8] ),
    .A2(\uart_proj.fifoRx.fifo[16] ),
    .A3(\uart_proj.fifoRx.fifo[24] ),
    .S1(net450),
    .X(_0479_));
 sg13g2_nor2_1 _1852_ (.A(net447),
    .B(_0479_),
    .Y(_0480_));
 sg13g2_nor2b_1 _1853_ (.A(\uart_proj.fifoRx.fifo[40] ),
    .B_N(net456),
    .Y(_0481_));
 sg13g2_nor2_1 _1854_ (.A(net456),
    .B(\uart_proj.fifoRx.fifo[32] ),
    .Y(_0482_));
 sg13g2_nor3_1 _1855_ (.A(net450),
    .B(_0481_),
    .C(_0482_),
    .Y(_0483_));
 sg13g2_nor2b_1 _1856_ (.A(\uart_proj.fifoRx.fifo[56] ),
    .B_N(net456),
    .Y(_0484_));
 sg13g2_o21ai_1 _1857_ (.B1(net450),
    .Y(_0485_),
    .A1(net456),
    .A2(\uart_proj.fifoRx.fifo[48] ));
 sg13g2_o21ai_1 _1858_ (.B1(net447),
    .Y(_0486_),
    .A1(_0484_),
    .A2(_0485_));
 sg13g2_o21ai_1 _1859_ (.B1(net440),
    .Y(_0487_),
    .A1(_0483_),
    .A2(_0486_));
 sg13g2_nor2_2 _1860_ (.A(_0480_),
    .B(_0487_),
    .Y(uio_out[0]));
 sg13g2_nand2b_1 _1861_ (.Y(_0488_),
    .B(net461),
    .A_N(\uart_proj.fifoRx.fifo[9] ));
 sg13g2_o21ai_1 _1862_ (.B1(_0488_),
    .Y(_0489_),
    .A1(net461),
    .A2(\uart_proj.fifoRx.fifo[1] ));
 sg13g2_mux2_1 _1863_ (.A0(\uart_proj.fifoRx.fifo[17] ),
    .A1(\uart_proj.fifoRx.fifo[25] ),
    .S(net456),
    .X(_0490_));
 sg13g2_a21oi_1 _1864_ (.A1(net450),
    .A2(_0490_),
    .Y(_0491_),
    .B1(net447));
 sg13g2_o21ai_1 _1865_ (.B1(_0491_),
    .Y(_0492_),
    .A1(net452),
    .A2(_0489_));
 sg13g2_nor2b_1 _1866_ (.A(\uart_proj.fifoRx.fifo[41] ),
    .B_N(net460),
    .Y(_0493_));
 sg13g2_nor2_1 _1867_ (.A(net462),
    .B(\uart_proj.fifoRx.fifo[33] ),
    .Y(_0494_));
 sg13g2_nor3_1 _1868_ (.A(net452),
    .B(_0493_),
    .C(_0494_),
    .Y(_0495_));
 sg13g2_nor2b_1 _1869_ (.A(\uart_proj.fifoRx.fifo[57] ),
    .B_N(net457),
    .Y(_0496_));
 sg13g2_o21ai_1 _1870_ (.B1(net450),
    .Y(_0497_),
    .A1(net457),
    .A2(\uart_proj.fifoRx.fifo[49] ));
 sg13g2_o21ai_1 _1871_ (.B1(net447),
    .Y(_0498_),
    .A1(_0496_),
    .A2(_0497_));
 sg13g2_o21ai_1 _1872_ (.B1(net440),
    .Y(_0499_),
    .A1(_0495_),
    .A2(_0498_));
 sg13g2_nor2b_2 _1873_ (.A(_0499_),
    .B_N(_0492_),
    .Y(uio_out[1]));
 sg13g2_nand2b_1 _1874_ (.Y(_0500_),
    .B(net460),
    .A_N(\uart_proj.fifoRx.fifo[10] ));
 sg13g2_o21ai_1 _1875_ (.B1(_0500_),
    .Y(_0501_),
    .A1(net460),
    .A2(\uart_proj.fifoRx.fifo[2] ));
 sg13g2_mux2_2 _1876_ (.A0(\uart_proj.fifoRx.fifo[18] ),
    .A1(\uart_proj.fifoRx.fifo[26] ),
    .S(net456),
    .X(_0502_));
 sg13g2_a21oi_1 _1877_ (.A1(net453),
    .A2(_0502_),
    .Y(_0503_),
    .B1(net448));
 sg13g2_o21ai_1 _1878_ (.B1(_0503_),
    .Y(_0504_),
    .A1(net452),
    .A2(_0501_));
 sg13g2_nor2b_1 _1879_ (.A(\uart_proj.fifoRx.fifo[42] ),
    .B_N(net460),
    .Y(_0505_));
 sg13g2_nor2_1 _1880_ (.A(net460),
    .B(\uart_proj.fifoRx.fifo[34] ),
    .Y(_0506_));
 sg13g2_nor3_1 _1881_ (.A(net452),
    .B(_0505_),
    .C(_0506_),
    .Y(_0507_));
 sg13g2_nor2b_1 _1882_ (.A(\uart_proj.fifoRx.fifo[58] ),
    .B_N(net460),
    .Y(_0508_));
 sg13g2_o21ai_1 _1883_ (.B1(net453),
    .Y(_0509_),
    .A1(net460),
    .A2(\uart_proj.fifoRx.fifo[50] ));
 sg13g2_o21ai_1 _1884_ (.B1(net448),
    .Y(_0510_),
    .A1(_0508_),
    .A2(_0509_));
 sg13g2_o21ai_1 _1885_ (.B1(net440),
    .Y(_0511_),
    .A1(_0507_),
    .A2(_0510_));
 sg13g2_nor2b_1 _1886_ (.A(_0511_),
    .B_N(_0504_),
    .Y(uio_out[2]));
 sg13g2_mux4_1 _1887_ (.S0(net454),
    .A0(\uart_proj.fifoRx.fifo[3] ),
    .A1(\uart_proj.fifoRx.fifo[11] ),
    .A2(\uart_proj.fifoRx.fifo[19] ),
    .A3(\uart_proj.fifoRx.fifo[27] ),
    .S1(net449),
    .X(_0512_));
 sg13g2_nor2_1 _1888_ (.A(net446),
    .B(_0512_),
    .Y(_0513_));
 sg13g2_nor2b_1 _1889_ (.A(\uart_proj.fifoRx.fifo[43] ),
    .B_N(net454),
    .Y(_0514_));
 sg13g2_nor2_1 _1890_ (.A(net455),
    .B(\uart_proj.fifoRx.fifo[35] ),
    .Y(_0515_));
 sg13g2_nor3_1 _1891_ (.A(net449),
    .B(_0514_),
    .C(_0515_),
    .Y(_0516_));
 sg13g2_nor2b_1 _1892_ (.A(\uart_proj.fifoRx.fifo[59] ),
    .B_N(net455),
    .Y(_0517_));
 sg13g2_o21ai_1 _1893_ (.B1(net449),
    .Y(_0518_),
    .A1(net455),
    .A2(\uart_proj.fifoRx.fifo[51] ));
 sg13g2_o21ai_1 _1894_ (.B1(net446),
    .Y(_0519_),
    .A1(_0517_),
    .A2(_0518_));
 sg13g2_o21ai_1 _1895_ (.B1(net440),
    .Y(_0520_),
    .A1(_0516_),
    .A2(_0519_));
 sg13g2_nor2_2 _1896_ (.A(_0513_),
    .B(_0520_),
    .Y(uio_out[3]));
 sg13g2_nand2b_1 _1897_ (.Y(_0521_),
    .B(net458),
    .A_N(\uart_proj.fifoRx.fifo[12] ));
 sg13g2_o21ai_1 _1898_ (.B1(_0521_),
    .Y(_0522_),
    .A1(net458),
    .A2(\uart_proj.fifoRx.fifo[4] ));
 sg13g2_mux2_1 _1899_ (.A0(\uart_proj.fifoRx.fifo[20] ),
    .A1(\uart_proj.fifoRx.fifo[28] ),
    .S(net456),
    .X(_0523_));
 sg13g2_a21oi_2 _1900_ (.B1(net446),
    .Y(_0524_),
    .A2(_0523_),
    .A1(net450));
 sg13g2_o21ai_1 _1901_ (.B1(_0524_),
    .Y(_0525_),
    .A1(net452),
    .A2(_0522_));
 sg13g2_nor2b_1 _1902_ (.A(\uart_proj.fifoRx.fifo[44] ),
    .B_N(net462),
    .Y(_0526_));
 sg13g2_nor2_1 _1903_ (.A(net462),
    .B(\uart_proj.fifoRx.fifo[36] ),
    .Y(_0527_));
 sg13g2_nor3_1 _1904_ (.A(net451),
    .B(_0526_),
    .C(_0527_),
    .Y(_0528_));
 sg13g2_nor2b_1 _1905_ (.A(\uart_proj.fifoRx.fifo[60] ),
    .B_N(net459),
    .Y(_0529_));
 sg13g2_o21ai_1 _1906_ (.B1(net451),
    .Y(_0530_),
    .A1(net459),
    .A2(\uart_proj.fifoRx.fifo[52] ));
 sg13g2_o21ai_1 _1907_ (.B1(net448),
    .Y(_0531_),
    .A1(_0529_),
    .A2(_0530_));
 sg13g2_o21ai_1 _1908_ (.B1(_0378_),
    .Y(_0532_),
    .A1(_0528_),
    .A2(_0531_));
 sg13g2_nor2b_2 _1909_ (.A(_0532_),
    .B_N(_0525_),
    .Y(uio_out[4]));
 sg13g2_nand2b_1 _1910_ (.Y(_0533_),
    .B(net459),
    .A_N(\uart_proj.fifoRx.fifo[13] ));
 sg13g2_o21ai_1 _1911_ (.B1(_0533_),
    .Y(_0534_),
    .A1(net459),
    .A2(\uart_proj.fifoRx.fifo[5] ));
 sg13g2_mux2_1 _1912_ (.A0(\uart_proj.fifoRx.fifo[21] ),
    .A1(\uart_proj.fifoRx.fifo[29] ),
    .S(net454),
    .X(_0535_));
 sg13g2_a21oi_1 _1913_ (.A1(net449),
    .A2(_0535_),
    .Y(_0536_),
    .B1(net446));
 sg13g2_o21ai_1 _1914_ (.B1(_0536_),
    .Y(_0537_),
    .A1(net451),
    .A2(_0534_));
 sg13g2_nor2b_1 _1915_ (.A(\uart_proj.fifoRx.fifo[45] ),
    .B_N(net459),
    .Y(_0538_));
 sg13g2_nor2_1 _1916_ (.A(net459),
    .B(\uart_proj.fifoRx.fifo[37] ),
    .Y(_0539_));
 sg13g2_nor3_1 _1917_ (.A(net451),
    .B(_0538_),
    .C(_0539_),
    .Y(_0540_));
 sg13g2_nor2b_1 _1918_ (.A(\uart_proj.fifoRx.fifo[61] ),
    .B_N(net459),
    .Y(_0541_));
 sg13g2_o21ai_1 _1919_ (.B1(net451),
    .Y(_0542_),
    .A1(net459),
    .A2(\uart_proj.fifoRx.fifo[53] ));
 sg13g2_o21ai_1 _1920_ (.B1(net446),
    .Y(_0543_),
    .A1(_0541_),
    .A2(_0542_));
 sg13g2_o21ai_1 _1921_ (.B1(_0378_),
    .Y(_0544_),
    .A1(_0540_),
    .A2(_0543_));
 sg13g2_nor2b_2 _1922_ (.A(_0544_),
    .B_N(_0537_),
    .Y(uio_out[5]));
 sg13g2_mux4_1 _1923_ (.S0(net454),
    .A0(\uart_proj.fifoRx.fifo[6] ),
    .A1(\uart_proj.fifoRx.fifo[14] ),
    .A2(\uart_proj.fifoRx.fifo[22] ),
    .A3(\uart_proj.fifoRx.fifo[30] ),
    .S1(net449),
    .X(_0545_));
 sg13g2_nor2_1 _1924_ (.A(net446),
    .B(_0545_),
    .Y(_0546_));
 sg13g2_nor2b_1 _1925_ (.A(\uart_proj.fifoRx.fifo[46] ),
    .B_N(net454),
    .Y(_0547_));
 sg13g2_nor2_1 _1926_ (.A(net454),
    .B(\uart_proj.fifoRx.fifo[38] ),
    .Y(_0548_));
 sg13g2_nor3_1 _1927_ (.A(net449),
    .B(_0547_),
    .C(_0548_),
    .Y(_0549_));
 sg13g2_nor2b_1 _1928_ (.A(\uart_proj.fifoRx.fifo[62] ),
    .B_N(net455),
    .Y(_0550_));
 sg13g2_o21ai_1 _1929_ (.B1(net449),
    .Y(_0551_),
    .A1(net454),
    .A2(\uart_proj.fifoRx.fifo[54] ));
 sg13g2_o21ai_1 _1930_ (.B1(net446),
    .Y(_0552_),
    .A1(_0550_),
    .A2(_0551_));
 sg13g2_o21ai_1 _1931_ (.B1(net440),
    .Y(_0553_),
    .A1(_0549_),
    .A2(_0552_));
 sg13g2_nor2_2 _1932_ (.A(_0546_),
    .B(_0553_),
    .Y(uio_out[6]));
 sg13g2_nand2b_1 _1933_ (.Y(_0554_),
    .B(net458),
    .A_N(\uart_proj.fifoRx.fifo[15] ));
 sg13g2_o21ai_1 _1934_ (.B1(_0554_),
    .Y(_0555_),
    .A1(net458),
    .A2(\uart_proj.fifoRx.fifo[7] ));
 sg13g2_mux2_1 _1935_ (.A0(\uart_proj.fifoRx.fifo[23] ),
    .A1(\uart_proj.fifoRx.fifo[31] ),
    .S(net454),
    .X(_0556_));
 sg13g2_a21oi_2 _1936_ (.B1(net446),
    .Y(_0557_),
    .A2(_0556_),
    .A1(net449));
 sg13g2_o21ai_1 _1937_ (.B1(_0557_),
    .Y(_0558_),
    .A1(net451),
    .A2(_0555_));
 sg13g2_nor2b_1 _1938_ (.A(\uart_proj.fifoRx.fifo[47] ),
    .B_N(net458),
    .Y(_0559_));
 sg13g2_nor2_1 _1939_ (.A(net458),
    .B(\uart_proj.fifoRx.fifo[39] ),
    .Y(_0560_));
 sg13g2_nor3_1 _1940_ (.A(net451),
    .B(_0559_),
    .C(_0560_),
    .Y(_0561_));
 sg13g2_nor2b_1 _1941_ (.A(\uart_proj.fifoRx.fifo[63] ),
    .B_N(net458),
    .Y(_0562_));
 sg13g2_o21ai_1 _1942_ (.B1(net451),
    .Y(_0563_),
    .A1(net458),
    .A2(\uart_proj.fifoRx.fifo[55] ));
 sg13g2_o21ai_1 _1943_ (.B1(net448),
    .Y(_0564_),
    .A1(_0562_),
    .A2(_0563_));
 sg13g2_o21ai_1 _1944_ (.B1(net440),
    .Y(_0565_),
    .A1(_0561_),
    .A2(_0564_));
 sg13g2_nor2b_1 _1945_ (.A(_0565_),
    .B_N(_0558_),
    .Y(uio_out[7]));
 sg13g2_a21oi_1 _1946_ (.A1(net480),
    .A2(net428),
    .Y(_0566_),
    .B1(net531));
 sg13g2_xnor2_1 _1947_ (.Y(_0137_),
    .A(_0126_),
    .B(_0566_));
 sg13g2_a21oi_1 _1948_ (.A1(\uart_proj.bg.rate[2] ),
    .A2(net428),
    .Y(_0567_),
    .B1(net541));
 sg13g2_a21oi_1 _1949_ (.A1(_0126_),
    .A2(_0566_),
    .Y(_0568_),
    .B1(_0567_));
 sg13g2_nand3_1 _1950_ (.B(_0566_),
    .C(_0567_),
    .A(_0126_),
    .Y(_0569_));
 sg13g2_nand2b_1 _1951_ (.Y(_0138_),
    .B(_0569_),
    .A_N(_0568_));
 sg13g2_nor3_2 _1952_ (.A(_0903_),
    .B(_0932_),
    .C(_0936_),
    .Y(_0570_));
 sg13g2_nor2_1 _1953_ (.A(net551),
    .B(_0570_),
    .Y(_0571_));
 sg13g2_nand2b_1 _1954_ (.Y(_0572_),
    .B(_0571_),
    .A_N(_0569_));
 sg13g2_xor2_1 _1955_ (.B(_0571_),
    .A(_0569_),
    .X(_0139_));
 sg13g2_a21oi_1 _1956_ (.A1(net480),
    .A2(net427),
    .Y(_0573_),
    .B1(net353));
 sg13g2_nand2b_1 _1957_ (.Y(_0574_),
    .B(_0573_),
    .A_N(_0572_));
 sg13g2_xor2_1 _1958_ (.B(_0573_),
    .A(_0572_),
    .X(_0140_));
 sg13g2_a21oi_1 _1959_ (.A1(\uart_proj.bg.rate[5] ),
    .A2(net428),
    .Y(_0575_),
    .B1(net385));
 sg13g2_nand2b_1 _1960_ (.Y(_0576_),
    .B(net386),
    .A_N(_0574_));
 sg13g2_xor2_1 _1961_ (.B(net386),
    .A(_0574_),
    .X(_0141_));
 sg13g2_o21ai_1 _1962_ (.B1(_0950_),
    .Y(_0577_),
    .A1(_0909_),
    .A2(net427));
 sg13g2_nand2b_1 _1963_ (.Y(_0578_),
    .B(_0577_),
    .A_N(_0576_));
 sg13g2_xor2_1 _1964_ (.B(_0577_),
    .A(_0576_),
    .X(_0142_));
 sg13g2_a21oi_1 _1965_ (.A1(\uart_proj.bg.rate[7] ),
    .A2(net427),
    .Y(_0579_),
    .B1(net537));
 sg13g2_nand2b_1 _1966_ (.Y(_0580_),
    .B(_0579_),
    .A_N(_0578_));
 sg13g2_xor2_1 _1967_ (.B(net538),
    .A(_0578_),
    .X(_0143_));
 sg13g2_a21oi_1 _1968_ (.A1(\uart_proj.bg.rate[8] ),
    .A2(net427),
    .Y(_0581_),
    .B1(net396));
 sg13g2_nand2b_1 _1969_ (.Y(_0582_),
    .B(_0581_),
    .A_N(_0580_));
 sg13g2_xor2_1 _1970_ (.B(_0581_),
    .A(_0580_),
    .X(_0144_));
 sg13g2_nor2_1 _1971_ (.A(net550),
    .B(_0570_),
    .Y(_0583_));
 sg13g2_nand2b_1 _1972_ (.Y(_0584_),
    .B(_0583_),
    .A_N(_0582_));
 sg13g2_xor2_1 _1973_ (.B(_0583_),
    .A(_0582_),
    .X(_0145_));
 sg13g2_nor2_1 _1974_ (.A(net383),
    .B(net427),
    .Y(_0585_));
 sg13g2_a21oi_1 _1975_ (.A1(\uart_proj.bg.rate[10] ),
    .A2(net427),
    .Y(_0586_),
    .B1(_0585_));
 sg13g2_nand2b_1 _1976_ (.Y(_0587_),
    .B(_0586_),
    .A_N(_0584_));
 sg13g2_xor2_1 _1977_ (.B(_0586_),
    .A(_0584_),
    .X(_0127_));
 sg13g2_nor2_1 _1978_ (.A(net549),
    .B(_0570_),
    .Y(_0588_));
 sg13g2_nand2b_2 _1979_ (.Y(_0589_),
    .B(_0588_),
    .A_N(_0587_));
 sg13g2_xor2_1 _1980_ (.B(_0588_),
    .A(_0587_),
    .X(_0128_));
 sg13g2_nor2_1 _1981_ (.A(net539),
    .B(net427),
    .Y(_0590_));
 sg13g2_a21oi_2 _1982_ (.B1(_0590_),
    .Y(_0591_),
    .A2(net427),
    .A1(_0901_));
 sg13g2_xnor2_1 _1983_ (.Y(_0129_),
    .A(_0589_),
    .B(_0591_));
 sg13g2_nor3_2 _1984_ (.A(net377),
    .B(_0589_),
    .C(_0591_),
    .Y(_0592_));
 sg13g2_o21ai_1 _1985_ (.B1(net377),
    .Y(_0593_),
    .A1(_0589_),
    .A2(_0591_));
 sg13g2_nand2b_1 _1986_ (.Y(_0130_),
    .B(_0593_),
    .A_N(_0592_));
 sg13g2_nand2b_2 _1987_ (.Y(_0594_),
    .B(_0592_),
    .A_N(net323));
 sg13g2_xor2_1 _1988_ (.B(_0592_),
    .A(net323),
    .X(_0131_));
 sg13g2_nor2_1 _1989_ (.A(\uart_proj.bg.txCount[15] ),
    .B(_0594_),
    .Y(_0595_));
 sg13g2_xnor2_1 _1990_ (.Y(_0132_),
    .A(net343),
    .B(_0594_));
 sg13g2_nor3_2 _1991_ (.A(\uart_proj.bg.txCount[16] ),
    .B(\uart_proj.bg.txCount[15] ),
    .C(_0594_),
    .Y(_0596_));
 sg13g2_xor2_1 _1992_ (.B(_0595_),
    .A(net340),
    .X(_0133_));
 sg13g2_nand2b_1 _1993_ (.Y(_0597_),
    .B(_0596_),
    .A_N(net325));
 sg13g2_xor2_1 _1994_ (.B(_0596_),
    .A(net325),
    .X(_0134_));
 sg13g2_nor2_1 _1995_ (.A(\uart_proj.bg.txCount[18] ),
    .B(_0597_),
    .Y(_0598_));
 sg13g2_xnor2_1 _1996_ (.Y(_0135_),
    .A(net338),
    .B(_0597_));
 sg13g2_xor2_1 _1997_ (.B(_0598_),
    .A(net327),
    .X(_0136_));
 sg13g2_nand2_2 _1998_ (.Y(_0599_),
    .A(_0945_),
    .B(net414));
 sg13g2_nor2_1 _1999_ (.A(_0031_),
    .B(net412),
    .Y(_0600_));
 sg13g2_nand2_2 _2000_ (.Y(_0601_),
    .A(_0406_),
    .B(_0600_));
 sg13g2_inv_1 _2001_ (.Y(_0602_),
    .A(_0601_));
 sg13g2_and2_1 _2002_ (.A(_0599_),
    .B(_0601_),
    .X(_0603_));
 sg13g2_nor2_1 _2003_ (.A(net350),
    .B(_0599_),
    .Y(_0604_));
 sg13g2_a21o_1 _2004_ (.A2(net410),
    .A1(net350),
    .B1(_0604_),
    .X(_0163_));
 sg13g2_a21oi_1 _2005_ (.A1(net280),
    .A2(_0601_),
    .Y(_0605_),
    .B1(_0604_));
 sg13g2_a21oi_1 _2006_ (.A1(net280),
    .A2(_0604_),
    .Y(_0164_),
    .B1(_0605_));
 sg13g2_nand2_1 _2007_ (.Y(_0606_),
    .A(net282),
    .B(net410));
 sg13g2_o21ai_1 _2008_ (.B1(net282),
    .Y(_0607_),
    .A1(\uart_proj.uartTx.writeCount[0] ),
    .A2(\uart_proj.uartTx.writeCount[1] ));
 sg13g2_nor2b_1 _2009_ (.A(_0952_),
    .B_N(_0607_),
    .Y(_0608_));
 sg13g2_o21ai_1 _2010_ (.B1(_0606_),
    .Y(_0165_),
    .A1(_0599_),
    .A2(_0608_));
 sg13g2_nand2_1 _2011_ (.Y(_0609_),
    .A(net118),
    .B(net410));
 sg13g2_xor2_1 _2012_ (.B(_0952_),
    .A(\uart_proj.uartTx.writeCount[3] ),
    .X(_0610_));
 sg13g2_o21ai_1 _2013_ (.B1(_0609_),
    .Y(_0166_),
    .A1(_0599_),
    .A2(_0610_));
 sg13g2_o21ai_1 _2014_ (.B1(_0962_),
    .Y(_0611_),
    .A1(\uart_proj.fifoRx.count[3] ),
    .A2(net440));
 sg13g2_nand2_2 _2015_ (.Y(_0612_),
    .A(\uart_proj.fifoRx.WEN ),
    .B(_0611_));
 sg13g2_nor2_2 _2016_ (.A(_1201_),
    .B(_0612_),
    .Y(_0613_));
 sg13g2_nand2b_1 _2017_ (.Y(_0614_),
    .B(_0613_),
    .A_N(\uart_proj.fifoRx.write_ptr[2] ));
 sg13g2_or3_2 _2018_ (.A(\uart_proj.fifoRx.write_ptr[0] ),
    .B(\uart_proj.fifoRx.write_ptr[1] ),
    .C(net419),
    .X(_0615_));
 sg13g2_mux2_1 _2019_ (.A0(\uart_proj.fifoRx.wdata[0] ),
    .A1(net303),
    .S(_0615_),
    .X(_0167_));
 sg13g2_mux2_1 _2020_ (.A0(\uart_proj.fifoRx.wdata[1] ),
    .A1(net290),
    .S(_0615_),
    .X(_0168_));
 sg13g2_mux2_1 _2021_ (.A0(\uart_proj.fifoRx.wdata[2] ),
    .A1(net307),
    .S(_0615_),
    .X(_0169_));
 sg13g2_mux2_1 _2022_ (.A0(\uart_proj.fifoRx.wdata[3] ),
    .A1(net286),
    .S(_0615_),
    .X(_0170_));
 sg13g2_mux2_1 _2023_ (.A0(\uart_proj.fifoRx.wdata[4] ),
    .A1(net305),
    .S(_0615_),
    .X(_0171_));
 sg13g2_mux2_1 _2024_ (.A0(\uart_proj.fifoRx.wdata[5] ),
    .A1(net299),
    .S(_0615_),
    .X(_0172_));
 sg13g2_mux2_1 _2025_ (.A0(\uart_proj.fifoRx.wdata[6] ),
    .A1(net295),
    .S(_0615_),
    .X(_0173_));
 sg13g2_mux2_1 _2026_ (.A0(\uart_proj.fifoRx.wdata[7] ),
    .A1(net293),
    .S(_0615_),
    .X(_0174_));
 sg13g2_nor2b_2 _2027_ (.A(\uart_proj.fifoRx.write_ptr[1] ),
    .B_N(\uart_proj.fifoRx.write_ptr[0] ),
    .Y(_0616_));
 sg13g2_nand2b_2 _2028_ (.Y(_0617_),
    .B(net435),
    .A_N(net419));
 sg13g2_nand2_1 _2029_ (.Y(_0618_),
    .A(net192),
    .B(_0617_));
 sg13g2_nand2_1 _2030_ (.Y(_0619_),
    .A(\uart_proj.fifoRx.wdata[0] ),
    .B(net435));
 sg13g2_o21ai_1 _2031_ (.B1(_0618_),
    .Y(_0175_),
    .A1(net419),
    .A2(_0619_));
 sg13g2_nand2_1 _2032_ (.Y(_0620_),
    .A(net107),
    .B(_0617_));
 sg13g2_nand2_1 _2033_ (.Y(_0621_),
    .A(\uart_proj.fifoRx.wdata[1] ),
    .B(net435));
 sg13g2_o21ai_1 _2034_ (.B1(_0620_),
    .Y(_0176_),
    .A1(net420),
    .A2(_0621_));
 sg13g2_nand2_1 _2035_ (.Y(_0622_),
    .A(net110),
    .B(_0617_));
 sg13g2_nand2_1 _2036_ (.Y(_0623_),
    .A(\uart_proj.fifoRx.wdata[2] ),
    .B(net435));
 sg13g2_o21ai_1 _2037_ (.B1(_0622_),
    .Y(_0177_),
    .A1(net420),
    .A2(_0623_));
 sg13g2_nand2_1 _2038_ (.Y(_0624_),
    .A(net158),
    .B(_0617_));
 sg13g2_nand2_1 _2039_ (.Y(_0625_),
    .A(\uart_proj.fifoRx.wdata[3] ),
    .B(net435));
 sg13g2_o21ai_1 _2040_ (.B1(_0624_),
    .Y(_0178_),
    .A1(net419),
    .A2(_0625_));
 sg13g2_nand2_1 _2041_ (.Y(_0626_),
    .A(net127),
    .B(_0617_));
 sg13g2_nand2_1 _2042_ (.Y(_0627_),
    .A(\uart_proj.fifoRx.wdata[4] ),
    .B(_0616_));
 sg13g2_o21ai_1 _2043_ (.B1(_0626_),
    .Y(_0179_),
    .A1(net420),
    .A2(_0627_));
 sg13g2_nand2_1 _2044_ (.Y(_0628_),
    .A(net137),
    .B(_0617_));
 sg13g2_nand2_1 _2045_ (.Y(_0629_),
    .A(\uart_proj.fifoRx.wdata[5] ),
    .B(_0616_));
 sg13g2_o21ai_1 _2046_ (.B1(_0628_),
    .Y(_0180_),
    .A1(net420),
    .A2(_0629_));
 sg13g2_nand2_1 _2047_ (.Y(_0630_),
    .A(net102),
    .B(_0617_));
 sg13g2_nand2_1 _2048_ (.Y(_0631_),
    .A(\uart_proj.fifoRx.wdata[6] ),
    .B(net435));
 sg13g2_o21ai_1 _2049_ (.B1(_0630_),
    .Y(_0181_),
    .A1(net419),
    .A2(_0631_));
 sg13g2_nand2_1 _2050_ (.Y(_0632_),
    .A(net149),
    .B(_0617_));
 sg13g2_nand2_1 _2051_ (.Y(_0633_),
    .A(\uart_proj.fifoRx.wdata[7] ),
    .B(_0616_));
 sg13g2_o21ai_1 _2052_ (.B1(_0632_),
    .Y(_0182_),
    .A1(net419),
    .A2(_0633_));
 sg13g2_nand2b_2 _2053_ (.Y(_0634_),
    .B(\uart_proj.fifoRx.write_ptr[1] ),
    .A_N(\uart_proj.fifoRx.write_ptr[0] ));
 sg13g2_nor2_2 _2054_ (.A(net419),
    .B(_0634_),
    .Y(_0635_));
 sg13g2_mux2_1 _2055_ (.A0(net264),
    .A1(\uart_proj.fifoRx.wdata[0] ),
    .S(_0635_),
    .X(_0183_));
 sg13g2_mux2_1 _2056_ (.A0(net167),
    .A1(\uart_proj.fifoRx.wdata[1] ),
    .S(_0635_),
    .X(_0184_));
 sg13g2_mux2_1 _2057_ (.A0(net174),
    .A1(\uart_proj.fifoRx.wdata[2] ),
    .S(_0635_),
    .X(_0185_));
 sg13g2_mux2_1 _2058_ (.A0(net259),
    .A1(\uart_proj.fifoRx.wdata[3] ),
    .S(_0635_),
    .X(_0186_));
 sg13g2_mux2_1 _2059_ (.A0(net151),
    .A1(\uart_proj.fifoRx.wdata[4] ),
    .S(_0635_),
    .X(_0187_));
 sg13g2_mux2_1 _2060_ (.A0(net169),
    .A1(\uart_proj.fifoRx.wdata[5] ),
    .S(_0635_),
    .X(_0188_));
 sg13g2_mux2_1 _2061_ (.A0(net218),
    .A1(\uart_proj.fifoRx.wdata[6] ),
    .S(_0635_),
    .X(_0189_));
 sg13g2_mux2_1 _2062_ (.A0(net139),
    .A1(\uart_proj.fifoRx.wdata[7] ),
    .S(_0635_),
    .X(_0190_));
 sg13g2_nand2_2 _2063_ (.Y(_0636_),
    .A(\uart_proj.fifoRx.write_ptr[0] ),
    .B(\uart_proj.fifoRx.write_ptr[1] ));
 sg13g2_nor2_2 _2064_ (.A(net419),
    .B(_0636_),
    .Y(_0637_));
 sg13g2_mux2_1 _2065_ (.A0(net189),
    .A1(\uart_proj.fifoRx.wdata[0] ),
    .S(_0637_),
    .X(_0191_));
 sg13g2_mux2_1 _2066_ (.A0(net204),
    .A1(\uart_proj.fifoRx.wdata[1] ),
    .S(_0637_),
    .X(_0192_));
 sg13g2_mux2_1 _2067_ (.A0(net266),
    .A1(\uart_proj.fifoRx.wdata[2] ),
    .S(_0637_),
    .X(_0193_));
 sg13g2_mux2_1 _2068_ (.A0(net284),
    .A1(\uart_proj.fifoRx.wdata[3] ),
    .S(_0637_),
    .X(_0194_));
 sg13g2_mux2_1 _2069_ (.A0(net202),
    .A1(\uart_proj.fifoRx.wdata[4] ),
    .S(_0637_),
    .X(_0195_));
 sg13g2_mux2_1 _2070_ (.A0(net223),
    .A1(\uart_proj.fifoRx.wdata[5] ),
    .S(_0637_),
    .X(_0196_));
 sg13g2_mux2_1 _2071_ (.A0(net243),
    .A1(\uart_proj.fifoRx.wdata[6] ),
    .S(_0637_),
    .X(_0197_));
 sg13g2_mux2_1 _2072_ (.A0(net220),
    .A1(\uart_proj.fifoRx.wdata[7] ),
    .S(_0637_),
    .X(_0198_));
 sg13g2_nand2_1 _2073_ (.Y(_0638_),
    .A(net36),
    .B(_0613_));
 sg13g2_o21ai_1 _2074_ (.B1(\uart_proj.fifoRx.write_ptr[2] ),
    .Y(_0639_),
    .A1(\uart_proj.fifoRx.write_ptr[0] ),
    .A2(\uart_proj.fifoRx.write_ptr[1] ));
 sg13g2_nand2b_1 _2075_ (.Y(_0640_),
    .B(_0636_),
    .A_N(\uart_proj.fifoRx.write_ptr[2] ));
 sg13g2_nand4_1 _2076_ (.B(_0613_),
    .C(_0639_),
    .A(_0040_),
    .Y(_0641_),
    .D(_0640_));
 sg13g2_nand2_2 _2077_ (.Y(_0642_),
    .A(\uart_proj.fifoRx.write_ptr[2] ),
    .B(_0613_));
 sg13g2_nor3_2 _2078_ (.A(\uart_proj.fifoRx.write_ptr[0] ),
    .B(\uart_proj.fifoRx.write_ptr[1] ),
    .C(net418),
    .Y(_0643_));
 sg13g2_a22oi_1 _2079_ (.Y(_0644_),
    .B1(_0643_),
    .B2(\uart_proj.fifoRx.wdata[0] ),
    .A2(_0641_),
    .A1(net268));
 sg13g2_inv_1 _2080_ (.Y(_0199_),
    .A(net269));
 sg13g2_a22oi_1 _2081_ (.Y(_0645_),
    .B1(_0643_),
    .B2(\uart_proj.fifoRx.wdata[1] ),
    .A2(_0641_),
    .A1(net180));
 sg13g2_inv_1 _2082_ (.Y(_0200_),
    .A(net181));
 sg13g2_a22oi_1 _2083_ (.Y(_0646_),
    .B1(_0643_),
    .B2(\uart_proj.fifoRx.wdata[2] ),
    .A2(_0641_),
    .A1(net208));
 sg13g2_inv_1 _2084_ (.Y(_0201_),
    .A(net209));
 sg13g2_a22oi_1 _2085_ (.Y(_0647_),
    .B1(_0643_),
    .B2(\uart_proj.fifoRx.wdata[3] ),
    .A2(_0641_),
    .A1(net172));
 sg13g2_inv_1 _2086_ (.Y(_0202_),
    .A(net173));
 sg13g2_a22oi_1 _2087_ (.Y(_0648_),
    .B1(_0643_),
    .B2(\uart_proj.fifoRx.wdata[4] ),
    .A2(_0641_),
    .A1(net206));
 sg13g2_inv_1 _2088_ (.Y(_0203_),
    .A(net207));
 sg13g2_a22oi_1 _2089_ (.Y(_0649_),
    .B1(_0643_),
    .B2(\uart_proj.fifoRx.wdata[5] ),
    .A2(_0641_),
    .A1(net196));
 sg13g2_inv_1 _2090_ (.Y(_0204_),
    .A(net197));
 sg13g2_a22oi_1 _2091_ (.Y(_0650_),
    .B1(_0643_),
    .B2(\uart_proj.fifoRx.wdata[6] ),
    .A2(_0641_),
    .A1(net252));
 sg13g2_inv_1 _2092_ (.Y(_0205_),
    .A(net253));
 sg13g2_a22oi_1 _2093_ (.Y(_0651_),
    .B1(_0643_),
    .B2(\uart_proj.fifoRx.wdata[7] ),
    .A2(_0641_),
    .A1(net153));
 sg13g2_inv_1 _2094_ (.Y(_0206_),
    .A(net154));
 sg13g2_nand3_1 _2095_ (.B(_0613_),
    .C(net435),
    .A(\uart_proj.fifoRx.write_ptr[2] ),
    .Y(_0652_));
 sg13g2_nand2_1 _2096_ (.Y(_0653_),
    .A(net176),
    .B(_0652_));
 sg13g2_o21ai_1 _2097_ (.B1(_0653_),
    .Y(_0207_),
    .A1(_0619_),
    .A2(net418));
 sg13g2_nand2_1 _2098_ (.Y(_0654_),
    .A(net116),
    .B(_0652_));
 sg13g2_o21ai_1 _2099_ (.B1(_0654_),
    .Y(_0208_),
    .A1(_0621_),
    .A2(net418));
 sg13g2_nand2_1 _2100_ (.Y(_0655_),
    .A(net145),
    .B(_0652_));
 sg13g2_o21ai_1 _2101_ (.B1(_0655_),
    .Y(_0209_),
    .A1(_0623_),
    .A2(net418));
 sg13g2_nand2_1 _2102_ (.Y(_0656_),
    .A(net125),
    .B(_0652_));
 sg13g2_o21ai_1 _2103_ (.B1(_0656_),
    .Y(_0210_),
    .A1(_0625_),
    .A2(net418));
 sg13g2_nand2_1 _2104_ (.Y(_0657_),
    .A(net104),
    .B(_0652_));
 sg13g2_o21ai_1 _2105_ (.B1(_0657_),
    .Y(_0211_),
    .A1(_0627_),
    .A2(_0642_));
 sg13g2_nand2_1 _2106_ (.Y(_0658_),
    .A(net163),
    .B(_0652_));
 sg13g2_o21ai_1 _2107_ (.B1(_0658_),
    .Y(_0212_),
    .A1(_0629_),
    .A2(_0642_));
 sg13g2_nand2_1 _2108_ (.Y(_0659_),
    .A(net178),
    .B(_0652_));
 sg13g2_o21ai_1 _2109_ (.B1(_0659_),
    .Y(_0213_),
    .A1(_0631_),
    .A2(net418));
 sg13g2_nand2_1 _2110_ (.Y(_0660_),
    .A(net147),
    .B(_0652_));
 sg13g2_o21ai_1 _2111_ (.B1(_0660_),
    .Y(_0214_),
    .A1(_0633_),
    .A2(_0642_));
 sg13g2_nor2_2 _2112_ (.A(_0634_),
    .B(net418),
    .Y(_0661_));
 sg13g2_mux2_1 _2113_ (.A0(net225),
    .A1(\uart_proj.fifoRx.wdata[0] ),
    .S(_0661_),
    .X(_0215_));
 sg13g2_mux2_1 _2114_ (.A0(net200),
    .A1(\uart_proj.fifoRx.wdata[1] ),
    .S(_0661_),
    .X(_0216_));
 sg13g2_mux2_1 _2115_ (.A0(net247),
    .A1(\uart_proj.fifoRx.wdata[2] ),
    .S(_0661_),
    .X(_0217_));
 sg13g2_mux2_1 _2116_ (.A0(net228),
    .A1(\uart_proj.fifoRx.wdata[3] ),
    .S(_0661_),
    .X(_0218_));
 sg13g2_mux2_1 _2117_ (.A0(net314),
    .A1(\uart_proj.fifoRx.wdata[4] ),
    .S(_0661_),
    .X(_0219_));
 sg13g2_mux2_1 _2118_ (.A0(net239),
    .A1(\uart_proj.fifoRx.wdata[5] ),
    .S(_0661_),
    .X(_0220_));
 sg13g2_mux2_1 _2119_ (.A0(net278),
    .A1(\uart_proj.fifoRx.wdata[6] ),
    .S(_0661_),
    .X(_0221_));
 sg13g2_mux2_1 _2120_ (.A0(net276),
    .A1(\uart_proj.fifoRx.wdata[7] ),
    .S(_0661_),
    .X(_0222_));
 sg13g2_nor2_1 _2121_ (.A(_0612_),
    .B(_0636_),
    .Y(_0662_));
 sg13g2_nor2_2 _2122_ (.A(_0636_),
    .B(net418),
    .Y(_0663_));
 sg13g2_mux2_1 _2123_ (.A0(net212),
    .A1(\uart_proj.fifoRx.wdata[0] ),
    .S(_0663_),
    .X(_0223_));
 sg13g2_mux2_1 _2124_ (.A0(net198),
    .A1(\uart_proj.fifoRx.wdata[1] ),
    .S(_0663_),
    .X(_0224_));
 sg13g2_mux2_1 _2125_ (.A0(net273),
    .A1(\uart_proj.fifoRx.wdata[2] ),
    .S(_0663_),
    .X(_0225_));
 sg13g2_mux2_1 _2126_ (.A0(net257),
    .A1(\uart_proj.fifoRx.wdata[3] ),
    .S(_0663_),
    .X(_0226_));
 sg13g2_mux2_1 _2127_ (.A0(net255),
    .A1(\uart_proj.fifoRx.wdata[4] ),
    .S(_0663_),
    .X(_0227_));
 sg13g2_mux2_1 _2128_ (.A0(net250),
    .A1(\uart_proj.fifoRx.wdata[5] ),
    .S(_0663_),
    .X(_0228_));
 sg13g2_mux2_1 _2129_ (.A0(net184),
    .A1(\uart_proj.fifoRx.wdata[6] ),
    .S(_0663_),
    .X(_0229_));
 sg13g2_mux2_1 _2130_ (.A0(net210),
    .A1(\uart_proj.fifoRx.wdata[7] ),
    .S(_0663_),
    .X(_0230_));
 sg13g2_o21ai_1 _2131_ (.B1(_0959_),
    .Y(_0664_),
    .A1(_0917_),
    .A2(\uart_proj.fifoTx.count[3] ));
 sg13g2_and2_2 _2132_ (.A(net442),
    .B(_0664_),
    .X(_0665_));
 sg13g2_nand2_2 _2133_ (.Y(_0666_),
    .A(net442),
    .B(_0664_));
 sg13g2_o21ai_1 _2134_ (.B1(net443),
    .Y(_0667_),
    .A1(\uart_proj.fifoTx.write_ptr[0] ),
    .A2(_0665_));
 sg13g2_a21oi_1 _2135_ (.A1(_0923_),
    .A2(_0665_),
    .Y(_0231_),
    .B1(_0667_));
 sg13g2_nor2_2 _2136_ (.A(\uart_proj.fifoTx.write_ptr[0] ),
    .B(\uart_proj.fifoTx.write_ptr[1] ),
    .Y(_0668_));
 sg13g2_nand2_1 _2137_ (.Y(_0669_),
    .A(\uart_proj.fifoTx.write_ptr[0] ),
    .B(\uart_proj.fifoTx.write_ptr[1] ));
 sg13g2_nor2b_1 _2138_ (.A(_0668_),
    .B_N(_0669_),
    .Y(_0670_));
 sg13g2_nand2b_1 _2139_ (.Y(_0671_),
    .B(_0669_),
    .A_N(_0668_));
 sg13g2_o21ai_1 _2140_ (.B1(net443),
    .Y(_0672_),
    .A1(_0666_),
    .A2(net430));
 sg13g2_a21oi_1 _2141_ (.A1(_0924_),
    .A2(_0666_),
    .Y(_0232_),
    .B1(_0672_));
 sg13g2_nor2_2 _2142_ (.A(_0666_),
    .B(_0669_),
    .Y(_0673_));
 sg13g2_nand2_1 _2143_ (.Y(_0674_),
    .A(\uart_proj.fifoTx.write_ptr[2] ),
    .B(_0673_));
 sg13g2_o21ai_1 _2144_ (.B1(net443),
    .Y(_0675_),
    .A1(net544),
    .A2(_0673_));
 sg13g2_nor2b_1 _2145_ (.A(_0675_),
    .B_N(net417),
    .Y(_0233_));
 sg13g2_a21oi_1 _2146_ (.A1(\uart_proj.fifoTx.count[3] ),
    .A2(_1204_),
    .Y(_0676_),
    .B1(_0960_));
 sg13g2_nor2b_2 _2147_ (.A(_0676_),
    .B_N(\uart_proj.fifoTx.REN ),
    .Y(_0677_));
 sg13g2_o21ai_1 _2148_ (.B1(net443),
    .Y(_0678_),
    .A1(net471),
    .A2(_0677_));
 sg13g2_a21oi_1 _2149_ (.A1(_0921_),
    .A2(_0677_),
    .Y(_0234_),
    .B1(_0678_));
 sg13g2_a21oi_1 _2150_ (.A1(net471),
    .A2(_0677_),
    .Y(_0679_),
    .B1(net464));
 sg13g2_a221oi_1 _2151_ (.B2(_0677_),
    .C1(_0679_),
    .B1(net436),
    .A1(net445),
    .Y(_0235_),
    .A2(net312));
 sg13g2_xor2_1 _2152_ (.B(net436),
    .A(net317),
    .X(_0680_));
 sg13g2_o21ai_1 _2153_ (.B1(net443),
    .Y(_0681_),
    .A1(net463),
    .A2(_0677_));
 sg13g2_a21oi_1 _2154_ (.A1(_0677_),
    .A2(_0680_),
    .Y(_0236_),
    .B1(_0681_));
 sg13g2_nor2_2 _2155_ (.A(net230),
    .B(_0963_),
    .Y(_0682_));
 sg13g2_nor2_1 _2156_ (.A(net135),
    .B(net231),
    .Y(_0683_));
 sg13g2_nor2_1 _2157_ (.A(_1201_),
    .B(_0683_),
    .Y(_0237_));
 sg13g2_nand3_1 _2158_ (.B(net443),
    .C(_0612_),
    .A(\uart_proj.fifoRx.write_ptr[0] ),
    .Y(_0684_));
 sg13g2_nand2_1 _2159_ (.Y(_0238_),
    .A(net37),
    .B(_0684_));
 sg13g2_and3_1 _2160_ (.X(_0685_),
    .A(net552),
    .B(net443),
    .C(_0612_));
 sg13g2_nand2b_1 _2161_ (.Y(_0686_),
    .B(_0634_),
    .A_N(net435));
 sg13g2_a21o_1 _2162_ (.A2(_0686_),
    .A1(_0613_),
    .B1(_0685_),
    .X(_0239_));
 sg13g2_o21ai_1 _2163_ (.B1(net443),
    .Y(_0687_),
    .A1(net345),
    .A2(_0662_));
 sg13g2_a21oi_1 _2164_ (.A1(net345),
    .A2(_0662_),
    .Y(_0240_),
    .B1(_0687_));
 sg13g2_nor3_2 _2165_ (.A(\uart_proj.fifoRx.empty ),
    .B(_0379_),
    .C(_0682_),
    .Y(_0688_));
 sg13g2_nor2_1 _2166_ (.A(_1201_),
    .B(_0688_),
    .Y(_0689_));
 sg13g2_inv_1 _2167_ (.Y(_0690_),
    .A(_0689_));
 sg13g2_nor2_1 _2168_ (.A(net461),
    .B(_0688_),
    .Y(_0691_));
 sg13g2_a21oi_1 _2169_ (.A1(net461),
    .A2(_0690_),
    .Y(_0241_),
    .B1(_0691_));
 sg13g2_a21oi_1 _2170_ (.A1(net461),
    .A2(_0690_),
    .Y(_0692_),
    .B1(net452));
 sg13g2_nand2_1 _2171_ (.Y(_0693_),
    .A(net460),
    .B(net452));
 sg13g2_nand2_1 _2172_ (.Y(_0694_),
    .A(_1202_),
    .B(_0693_));
 sg13g2_a21oi_1 _2173_ (.A1(_0690_),
    .A2(_0694_),
    .Y(_0242_),
    .B1(_0692_));
 sg13g2_xor2_1 _2174_ (.B(_0693_),
    .A(net301),
    .X(_0695_));
 sg13g2_a22oi_1 _2175_ (.Y(_0696_),
    .B1(_0695_),
    .B2(_0688_),
    .A2(_0689_),
    .A1(net448));
 sg13g2_inv_1 _2176_ (.Y(_0243_),
    .A(net302));
 sg13g2_a21o_1 _2177_ (.A2(_1150_),
    .A1(_1020_),
    .B1(net431),
    .X(_0697_));
 sg13g2_a21oi_2 _2178_ (.B1(net363),
    .Y(_0698_),
    .A2(net431),
    .A1(net481));
 sg13g2_mux2_1 _2179_ (.A0(net363),
    .A1(_0698_),
    .S(net404),
    .X(_0244_));
 sg13g2_nor2_1 _2180_ (.A(net369),
    .B(_0697_),
    .Y(_0699_));
 sg13g2_a21oi_2 _2181_ (.B1(net369),
    .Y(_0700_),
    .A2(net432),
    .A1(net479));
 sg13g2_nand2_1 _2182_ (.Y(_0701_),
    .A(_0698_),
    .B(_0700_));
 sg13g2_xor2_1 _2183_ (.B(_0700_),
    .A(_0698_),
    .X(_0702_));
 sg13g2_a21oi_1 _2184_ (.A1(net404),
    .A2(_0702_),
    .Y(_0245_),
    .B1(_0699_));
 sg13g2_nor2_1 _2185_ (.A(net333),
    .B(_0697_),
    .Y(_0703_));
 sg13g2_a21oi_1 _2186_ (.A1(\uart_proj.bg.rate[0] ),
    .A2(net432),
    .Y(_0704_),
    .B1(net333));
 sg13g2_nand3_1 _2187_ (.B(_0700_),
    .C(_0704_),
    .A(_0698_),
    .Y(_0705_));
 sg13g2_xnor2_1 _2188_ (.Y(_0706_),
    .A(_0701_),
    .B(_0704_));
 sg13g2_a21oi_1 _2189_ (.A1(net404),
    .A2(_0706_),
    .Y(_0246_),
    .B1(_0703_));
 sg13g2_nor2_1 _2190_ (.A(net318),
    .B(net404),
    .Y(_0707_));
 sg13g2_nand2_1 _2191_ (.Y(_0708_),
    .A(\uart_proj.bg.rate[7] ),
    .B(net432));
 sg13g2_nand2b_1 _2192_ (.Y(_0709_),
    .B(_0708_),
    .A_N(net318));
 sg13g2_or2_1 _2193_ (.X(_0710_),
    .B(_0709_),
    .A(_0705_));
 sg13g2_xor2_1 _2194_ (.B(_0709_),
    .A(_0705_),
    .X(_0711_));
 sg13g2_a21oi_1 _2195_ (.A1(_0697_),
    .A2(_0711_),
    .Y(_0247_),
    .B1(_0707_));
 sg13g2_a21oi_1 _2196_ (.A1(\uart_proj.bg.rate[8] ),
    .A2(net432),
    .Y(_0712_),
    .B1(net289));
 sg13g2_nand2b_1 _2197_ (.Y(_0713_),
    .B(_0712_),
    .A_N(_0710_));
 sg13g2_xnor2_1 _2198_ (.Y(_0714_),
    .A(_0710_),
    .B(_0712_));
 sg13g2_nor2_1 _2199_ (.A(net289),
    .B(net404),
    .Y(_0715_));
 sg13g2_a21oi_1 _2200_ (.A1(net404),
    .A2(_0714_),
    .Y(_0248_),
    .B1(_0715_));
 sg13g2_nor2_1 _2201_ (.A(net310),
    .B(net404),
    .Y(_0716_));
 sg13g2_a21oi_1 _2202_ (.A1(net474),
    .A2(net431),
    .Y(_0717_),
    .B1(net310));
 sg13g2_nand2b_1 _2203_ (.Y(_0718_),
    .B(_0717_),
    .A_N(_0713_));
 sg13g2_xnor2_1 _2204_ (.Y(_0719_),
    .A(_0713_),
    .B(_0717_));
 sg13g2_a21oi_1 _2205_ (.A1(net404),
    .A2(_0719_),
    .Y(_0249_),
    .B1(_0716_));
 sg13g2_nor2_1 _2206_ (.A(net316),
    .B(net431),
    .Y(_0720_));
 sg13g2_a21oi_1 _2207_ (.A1(_0902_),
    .A2(net431),
    .Y(_0721_),
    .B1(_0720_));
 sg13g2_or2_1 _2208_ (.X(_0722_),
    .B(_0721_),
    .A(_0718_));
 sg13g2_xor2_1 _2209_ (.B(_0721_),
    .A(_0718_),
    .X(_0723_));
 sg13g2_nor2_1 _2210_ (.A(net316),
    .B(net405),
    .Y(_0724_));
 sg13g2_a21oi_1 _2211_ (.A1(net405),
    .A2(_0723_),
    .Y(_0250_),
    .B1(_0724_));
 sg13g2_nor2_1 _2212_ (.A(net292),
    .B(net405),
    .Y(_0725_));
 sg13g2_a21oi_1 _2213_ (.A1(net474),
    .A2(net431),
    .Y(_0726_),
    .B1(net292));
 sg13g2_nor2b_1 _2214_ (.A(_0722_),
    .B_N(_0726_),
    .Y(_0727_));
 sg13g2_xnor2_1 _2215_ (.Y(_0728_),
    .A(_0722_),
    .B(_0726_));
 sg13g2_a21oi_1 _2216_ (.A1(net405),
    .A2(_0728_),
    .Y(_0251_),
    .B1(_0725_));
 sg13g2_a21oi_1 _2217_ (.A1(net478),
    .A2(net431),
    .Y(_0729_),
    .B1(net311));
 sg13g2_xor2_1 _2218_ (.B(_0729_),
    .A(_0727_),
    .X(_0730_));
 sg13g2_nor2_1 _2219_ (.A(net311),
    .B(net405),
    .Y(_0731_));
 sg13g2_a21oi_1 _2220_ (.A1(net405),
    .A2(_0730_),
    .Y(_0252_),
    .B1(_0731_));
 sg13g2_nand3_1 _2221_ (.B(_0727_),
    .C(_0729_),
    .A(net405),
    .Y(_0732_));
 sg13g2_xnor2_1 _2222_ (.Y(_0253_),
    .A(net342),
    .B(_0732_));
 sg13g2_nor3_2 _2223_ (.A(\uart_proj.bg.rxCount[9] ),
    .B(net320),
    .C(_0732_),
    .Y(_0733_));
 sg13g2_o21ai_1 _2224_ (.B1(net320),
    .Y(_0734_),
    .A1(\uart_proj.bg.rxCount[9] ),
    .A2(_0732_));
 sg13g2_nand2b_1 _2225_ (.Y(_0254_),
    .B(net321),
    .A_N(_0733_));
 sg13g2_nand2b_1 _2226_ (.Y(_0735_),
    .B(_0733_),
    .A_N(net143));
 sg13g2_xor2_1 _2227_ (.B(_0733_),
    .A(net143),
    .X(_0255_));
 sg13g2_or2_1 _2228_ (.X(_0736_),
    .B(_0735_),
    .A(net262));
 sg13g2_xnor2_1 _2229_ (.Y(_0256_),
    .A(net262),
    .B(_0735_));
 sg13g2_xnor2_1 _2230_ (.Y(_0257_),
    .A(net309),
    .B(_0736_));
 sg13g2_nor3_1 _2231_ (.A(net309),
    .B(net319),
    .C(_0736_),
    .Y(_0737_));
 sg13g2_o21ai_1 _2232_ (.B1(net319),
    .Y(_0738_),
    .A1(net309),
    .A2(_0736_));
 sg13g2_nand2b_1 _2233_ (.Y(_0258_),
    .B(_0738_),
    .A_N(_0737_));
 sg13g2_xor2_1 _2234_ (.B(_0737_),
    .A(net94),
    .X(_0259_));
 sg13g2_nor2b_1 _2235_ (.A(net414),
    .B_N(\uart_proj.txData[0] ),
    .Y(_0739_));
 sg13g2_a21oi_1 _2236_ (.A1(net130),
    .A2(net412),
    .Y(_0740_),
    .B1(_0739_));
 sg13g2_nand2_1 _2237_ (.Y(_0741_),
    .A(net232),
    .B(net410));
 sg13g2_o21ai_1 _2238_ (.B1(_0741_),
    .Y(_0260_),
    .A1(net410),
    .A2(_0740_));
 sg13g2_nor2b_1 _2239_ (.A(net412),
    .B_N(\uart_proj.txData[1] ),
    .Y(_0742_));
 sg13g2_a21oi_1 _2240_ (.A1(\uart_proj.uartTx.writeBuf[2] ),
    .A2(net412),
    .Y(_0743_),
    .B1(_0742_));
 sg13g2_nand2_1 _2241_ (.Y(_0744_),
    .A(net130),
    .B(net409));
 sg13g2_o21ai_1 _2242_ (.B1(_0744_),
    .Y(_0261_),
    .A1(net409),
    .A2(_0743_));
 sg13g2_nor2b_1 _2243_ (.A(net413),
    .B_N(\uart_proj.txData[2] ),
    .Y(_0745_));
 sg13g2_a21oi_1 _2244_ (.A1(\uart_proj.uartTx.writeBuf[3] ),
    .A2(net413),
    .Y(_0746_),
    .B1(_0745_));
 sg13g2_nand2_1 _2245_ (.Y(_0747_),
    .A(net155),
    .B(net408));
 sg13g2_o21ai_1 _2246_ (.B1(_0747_),
    .Y(_0262_),
    .A1(net408),
    .A2(_0746_));
 sg13g2_nor2b_1 _2247_ (.A(net413),
    .B_N(\uart_proj.txData[3] ),
    .Y(_0748_));
 sg13g2_a21oi_1 _2248_ (.A1(net186),
    .A2(net413),
    .Y(_0749_),
    .B1(_0748_));
 sg13g2_nand2_1 _2249_ (.Y(_0750_),
    .A(net234),
    .B(net408));
 sg13g2_o21ai_1 _2250_ (.B1(_0750_),
    .Y(_0263_),
    .A1(net408),
    .A2(_0749_));
 sg13g2_nor2b_1 _2251_ (.A(net413),
    .B_N(\uart_proj.txData[4] ),
    .Y(_0751_));
 sg13g2_a21oi_1 _2252_ (.A1(net182),
    .A2(net413),
    .Y(_0752_),
    .B1(_0751_));
 sg13g2_nand2_1 _2253_ (.Y(_0753_),
    .A(net186),
    .B(net408));
 sg13g2_o21ai_1 _2254_ (.B1(_0753_),
    .Y(_0264_),
    .A1(net408),
    .A2(_0752_));
 sg13g2_nor2b_1 _2255_ (.A(net412),
    .B_N(\uart_proj.txData[5] ),
    .Y(_0754_));
 sg13g2_a21oi_1 _2256_ (.A1(net96),
    .A2(net412),
    .Y(_0755_),
    .B1(_0754_));
 sg13g2_nand2_1 _2257_ (.Y(_0756_),
    .A(net182),
    .B(net409));
 sg13g2_o21ai_1 _2258_ (.B1(_0756_),
    .Y(_0265_),
    .A1(net408),
    .A2(_0755_));
 sg13g2_nor2b_1 _2259_ (.A(net412),
    .B_N(\uart_proj.txData[6] ),
    .Y(_0757_));
 sg13g2_a21oi_1 _2260_ (.A1(\uart_proj.uartTx.writeBuf[7] ),
    .A2(net412),
    .Y(_0758_),
    .B1(_0757_));
 sg13g2_nand2_1 _2261_ (.Y(_0759_),
    .A(net96),
    .B(net408));
 sg13g2_o21ai_1 _2262_ (.B1(_0759_),
    .Y(_0266_),
    .A1(net409),
    .A2(_0758_));
 sg13g2_a22oi_1 _2263_ (.Y(_0760_),
    .B1(net410),
    .B2(\uart_proj.uartTx.writeBuf[7] ),
    .A2(_0602_),
    .A1(net120));
 sg13g2_inv_1 _2264_ (.Y(_0267_),
    .A(net121));
 sg13g2_nor2_1 _2265_ (.A(net124),
    .B(net407),
    .Y(_0761_));
 sg13g2_a21oi_1 _2266_ (.A1(net1),
    .A2(net407),
    .Y(_0268_),
    .B1(_0761_));
 sg13g2_nor2_1 _2267_ (.A(_0946_),
    .B(_0406_),
    .Y(_0762_));
 sg13g2_a21oi_1 _2268_ (.A1(_0918_),
    .A2(_0601_),
    .Y(_0269_),
    .B1(_0762_));
 sg13g2_o21ai_1 _2269_ (.B1(_0945_),
    .Y(_0763_),
    .A1(\uart_proj.fifoTx.REN ),
    .A2(net236));
 sg13g2_nor2_1 _2270_ (.A(net414),
    .B(_0763_),
    .Y(_0764_));
 sg13g2_nor2_1 _2271_ (.A(net329),
    .B(_0764_),
    .Y(_0765_));
 sg13g2_nor2_1 _2272_ (.A(_0762_),
    .B(net330),
    .Y(_0270_));
 sg13g2_xor2_1 _2273_ (.B(_1187_),
    .A(\uart_proj.uartRx.curState[0] ),
    .X(_0766_));
 sg13g2_nand2b_1 _2274_ (.Y(_0767_),
    .B(_0915_),
    .A_N(_1197_));
 sg13g2_o21ai_1 _2275_ (.B1(\uart_proj.uartRx.curState[2] ),
    .Y(_0768_),
    .A1(_1197_),
    .A2(_1198_));
 sg13g2_xnor2_1 _2276_ (.Y(_0769_),
    .A(\uart_proj.uartRx.curState[1] ),
    .B(_1194_));
 sg13g2_a21oi_2 _2277_ (.B1(_0769_),
    .Y(_0770_),
    .A2(_0768_),
    .A1(_0767_));
 sg13g2_nand2_2 _2278_ (.Y(_0771_),
    .A(_0766_),
    .B(_0770_));
 sg13g2_a21oi_1 _2279_ (.A1(_0766_),
    .A2(_0770_),
    .Y(_0772_),
    .B1(_1159_));
 sg13g2_o21ai_1 _2280_ (.B1(_1163_),
    .Y(_0271_),
    .A1(_0914_),
    .A2(_0772_));
 sg13g2_nor3_2 _2281_ (.A(\uart_proj.fifoTx.write_ptr[0] ),
    .B(\uart_proj.fifoTx.write_ptr[1] ),
    .C(\uart_proj.fifoTx.write_ptr[2] ),
    .Y(_0773_));
 sg13g2_nand2_2 _2282_ (.Y(_0774_),
    .A(_0665_),
    .B(net433));
 sg13g2_mux2_1 _2283_ (.A0(net7),
    .A1(net195),
    .S(_0774_),
    .X(_0272_));
 sg13g2_mux2_1 _2284_ (.A0(net8),
    .A1(net288),
    .S(_0774_),
    .X(_0273_));
 sg13g2_mux2_1 _2285_ (.A0(net9),
    .A1(net238),
    .S(_0774_),
    .X(_0274_));
 sg13g2_mux2_1 _2286_ (.A0(net10),
    .A1(net245),
    .S(_0774_),
    .X(_0275_));
 sg13g2_mux2_1 _2287_ (.A0(net11),
    .A1(net246),
    .S(_0774_),
    .X(_0276_));
 sg13g2_mux2_1 _2288_ (.A0(net12),
    .A1(net249),
    .S(_0774_),
    .X(_0277_));
 sg13g2_mux2_1 _2289_ (.A0(net13),
    .A1(net254),
    .S(_0774_),
    .X(_0278_));
 sg13g2_mux2_1 _2290_ (.A0(net14),
    .A1(net261),
    .S(_0774_),
    .X(_0279_));
 sg13g2_or4_2 _2291_ (.A(\uart_proj.fifoTx.write_ptr[1] ),
    .B(\uart_proj.fifoTx.write_ptr[2] ),
    .C(_0666_),
    .D(net433),
    .X(_0775_));
 sg13g2_nand2_1 _2292_ (.Y(_0776_),
    .A(net70),
    .B(_0775_));
 sg13g2_nand2_2 _2293_ (.Y(_0777_),
    .A(net7),
    .B(net442));
 sg13g2_nor3_1 _2294_ (.A(_0037_),
    .B(net433),
    .C(_0777_),
    .Y(_0778_));
 sg13g2_nand2_1 _2295_ (.Y(_0779_),
    .A(_0670_),
    .B(_0778_));
 sg13g2_xnor2_1 _2296_ (.Y(_0780_),
    .A(\uart_proj.fifoTx.write_ptr[2] ),
    .B(_0668_));
 sg13g2_nand2_1 _2297_ (.Y(_0781_),
    .A(_0665_),
    .B(_0780_));
 sg13g2_o21ai_1 _2298_ (.B1(_0776_),
    .Y(_0280_),
    .A1(_0779_),
    .A2(net425));
 sg13g2_nand2_1 _2299_ (.Y(_0782_),
    .A(net91),
    .B(_0775_));
 sg13g2_nand2_2 _2300_ (.Y(_0783_),
    .A(net8),
    .B(net441));
 sg13g2_nor3_1 _2301_ (.A(_0037_),
    .B(net433),
    .C(_0783_),
    .Y(_0784_));
 sg13g2_nand2_2 _2302_ (.Y(_0785_),
    .A(net430),
    .B(_0784_));
 sg13g2_o21ai_1 _2303_ (.B1(_0782_),
    .Y(_0281_),
    .A1(net426),
    .A2(_0785_));
 sg13g2_nand2_1 _2304_ (.Y(_0786_),
    .A(net72),
    .B(_0775_));
 sg13g2_nand2_2 _2305_ (.Y(_0787_),
    .A(net9),
    .B(net441));
 sg13g2_nor3_2 _2306_ (.A(net473),
    .B(net433),
    .C(_0787_),
    .Y(_0788_));
 sg13g2_nand2_2 _2307_ (.Y(_0789_),
    .A(net430),
    .B(_0788_));
 sg13g2_o21ai_1 _2308_ (.B1(_0786_),
    .Y(_0282_),
    .A1(_0781_),
    .A2(_0789_));
 sg13g2_nand2_1 _2309_ (.Y(_0790_),
    .A(net57),
    .B(_0775_));
 sg13g2_nand2_2 _2310_ (.Y(_0791_),
    .A(net10),
    .B(net441));
 sg13g2_nor3_2 _2311_ (.A(net473),
    .B(_0773_),
    .C(_0791_),
    .Y(_0792_));
 sg13g2_nand2_2 _2312_ (.Y(_0793_),
    .A(net430),
    .B(_0792_));
 sg13g2_o21ai_1 _2313_ (.B1(_0790_),
    .Y(_0283_),
    .A1(net425),
    .A2(_0793_));
 sg13g2_nand2_1 _2314_ (.Y(_0794_),
    .A(net54),
    .B(_0775_));
 sg13g2_nand2_2 _2315_ (.Y(_0795_),
    .A(net11),
    .B(net441));
 sg13g2_nor3_2 _2316_ (.A(net473),
    .B(_0773_),
    .C(_0795_),
    .Y(_0796_));
 sg13g2_nand2_2 _2317_ (.Y(_0797_),
    .A(net430),
    .B(_0796_));
 sg13g2_o21ai_1 _2318_ (.B1(_0794_),
    .Y(_0284_),
    .A1(net425),
    .A2(_0797_));
 sg13g2_nand2_1 _2319_ (.Y(_0798_),
    .A(net62),
    .B(_0775_));
 sg13g2_nand2_2 _2320_ (.Y(_0799_),
    .A(net12),
    .B(net441));
 sg13g2_nor3_1 _2321_ (.A(net473),
    .B(net433),
    .C(_0799_),
    .Y(_0800_));
 sg13g2_nand2_2 _2322_ (.Y(_0801_),
    .A(net430),
    .B(_0800_));
 sg13g2_o21ai_1 _2323_ (.B1(_0798_),
    .Y(_0285_),
    .A1(net426),
    .A2(_0801_));
 sg13g2_nand2_1 _2324_ (.Y(_0802_),
    .A(net61),
    .B(_0775_));
 sg13g2_nand2_2 _2325_ (.Y(_0803_),
    .A(net13),
    .B(net441));
 sg13g2_nor3_2 _2326_ (.A(net473),
    .B(net433),
    .C(_0803_),
    .Y(_0804_));
 sg13g2_nand2_2 _2327_ (.Y(_0805_),
    .A(net430),
    .B(_0804_));
 sg13g2_o21ai_1 _2328_ (.B1(_0802_),
    .Y(_0286_),
    .A1(net426),
    .A2(_0805_));
 sg13g2_nand2_1 _2329_ (.Y(_0806_),
    .A(net79),
    .B(_0775_));
 sg13g2_nand2_2 _2330_ (.Y(_0807_),
    .A(net14),
    .B(net442));
 sg13g2_nor3_1 _2331_ (.A(net473),
    .B(net433),
    .C(_0807_),
    .Y(_0808_));
 sg13g2_nand2_2 _2332_ (.Y(_0809_),
    .A(net430),
    .B(_0808_));
 sg13g2_o21ai_1 _2333_ (.B1(_0806_),
    .Y(_0287_),
    .A1(net426),
    .A2(_0809_));
 sg13g2_nor4_2 _2334_ (.A(\uart_proj.fifoTx.write_ptr[0] ),
    .B(_0924_),
    .C(\uart_proj.fifoTx.write_ptr[2] ),
    .Y(_0810_),
    .D(_0666_));
 sg13g2_nor2_1 _2335_ (.A(net129),
    .B(net423),
    .Y(_0811_));
 sg13g2_a21oi_1 _2336_ (.A1(_0777_),
    .A2(net423),
    .Y(_0288_),
    .B1(_0811_));
 sg13g2_nor2_1 _2337_ (.A(net114),
    .B(net423),
    .Y(_0812_));
 sg13g2_a21oi_1 _2338_ (.A1(_0783_),
    .A2(net423),
    .Y(_0289_),
    .B1(_0812_));
 sg13g2_nor2_1 _2339_ (.A(net141),
    .B(net423),
    .Y(_0813_));
 sg13g2_a21oi_1 _2340_ (.A1(_0787_),
    .A2(net423),
    .Y(_0290_),
    .B1(_0813_));
 sg13g2_nor2_1 _2341_ (.A(net112),
    .B(net423),
    .Y(_0814_));
 sg13g2_a21oi_1 _2342_ (.A1(_0791_),
    .A2(_0810_),
    .Y(_0291_),
    .B1(_0814_));
 sg13g2_nor2_1 _2343_ (.A(net171),
    .B(net423),
    .Y(_0815_));
 sg13g2_a21oi_1 _2344_ (.A1(_0795_),
    .A2(net424),
    .Y(_0292_),
    .B1(_0815_));
 sg13g2_nor2_1 _2345_ (.A(net106),
    .B(net424),
    .Y(_0816_));
 sg13g2_a21oi_1 _2346_ (.A1(_0799_),
    .A2(net424),
    .Y(_0293_),
    .B1(_0816_));
 sg13g2_nor2_1 _2347_ (.A(net134),
    .B(net424),
    .Y(_0817_));
 sg13g2_a21oi_1 _2348_ (.A1(_0803_),
    .A2(net424),
    .Y(_0294_),
    .B1(_0817_));
 sg13g2_nor2_1 _2349_ (.A(net142),
    .B(net424),
    .Y(_0818_));
 sg13g2_a21oi_1 _2350_ (.A1(_0807_),
    .A2(net424),
    .Y(_0295_),
    .B1(_0818_));
 sg13g2_nand2b_2 _2351_ (.Y(_0819_),
    .B(_0673_),
    .A_N(\uart_proj.fifoTx.write_ptr[2] ));
 sg13g2_nand2_1 _2352_ (.Y(_0820_),
    .A(net84),
    .B(_0819_));
 sg13g2_nand2_1 _2353_ (.Y(_0821_),
    .A(_0671_),
    .B(_0778_));
 sg13g2_o21ai_1 _2354_ (.B1(_0820_),
    .Y(_0296_),
    .A1(net425),
    .A2(_0821_));
 sg13g2_nand2_1 _2355_ (.Y(_0822_),
    .A(net52),
    .B(_0819_));
 sg13g2_nand2_1 _2356_ (.Y(_0823_),
    .A(net429),
    .B(_0784_));
 sg13g2_o21ai_1 _2357_ (.B1(_0822_),
    .Y(_0297_),
    .A1(net425),
    .A2(_0823_));
 sg13g2_nand2_1 _2358_ (.Y(_0824_),
    .A(net74),
    .B(_0819_));
 sg13g2_nand2_2 _2359_ (.Y(_0825_),
    .A(net429),
    .B(_0788_));
 sg13g2_o21ai_1 _2360_ (.B1(_0824_),
    .Y(_0298_),
    .A1(net425),
    .A2(_0825_));
 sg13g2_nand2_1 _2361_ (.Y(_0826_),
    .A(net76),
    .B(_0819_));
 sg13g2_nand2_2 _2362_ (.Y(_0827_),
    .A(net429),
    .B(_0792_));
 sg13g2_o21ai_1 _2363_ (.B1(_0826_),
    .Y(_0299_),
    .A1(net425),
    .A2(_0827_));
 sg13g2_nand2_1 _2364_ (.Y(_0828_),
    .A(net83),
    .B(_0819_));
 sg13g2_nand2_2 _2365_ (.Y(_0829_),
    .A(net429),
    .B(_0796_));
 sg13g2_o21ai_1 _2366_ (.B1(_0828_),
    .Y(_0300_),
    .A1(net425),
    .A2(_0829_));
 sg13g2_nand2_1 _2367_ (.Y(_0830_),
    .A(net51),
    .B(_0819_));
 sg13g2_nand2_1 _2368_ (.Y(_0831_),
    .A(net429),
    .B(_0800_));
 sg13g2_o21ai_1 _2369_ (.B1(_0830_),
    .Y(_0301_),
    .A1(net426),
    .A2(_0831_));
 sg13g2_nand2_1 _2370_ (.Y(_0832_),
    .A(net73),
    .B(_0819_));
 sg13g2_nand2_2 _2371_ (.Y(_0833_),
    .A(net429),
    .B(_0804_));
 sg13g2_o21ai_1 _2372_ (.B1(_0832_),
    .Y(_0302_),
    .A1(net426),
    .A2(_0833_));
 sg13g2_nand2_1 _2373_ (.Y(_0834_),
    .A(net78),
    .B(_0819_));
 sg13g2_nand2_1 _2374_ (.Y(_0835_),
    .A(net429),
    .B(_0808_));
 sg13g2_o21ai_1 _2375_ (.B1(_0834_),
    .Y(_0303_),
    .A1(net426),
    .A2(_0835_));
 sg13g2_nand4_1 _2376_ (.B(_0665_),
    .C(net429),
    .A(net473),
    .Y(_0836_),
    .D(_0780_));
 sg13g2_nand2_2 _2377_ (.Y(_0837_),
    .A(_0664_),
    .B(_0668_));
 sg13g2_nor3_1 _2378_ (.A(net434),
    .B(_0777_),
    .C(_0837_),
    .Y(_0838_));
 sg13g2_a21o_1 _2379_ (.A2(_0836_),
    .A1(net166),
    .B1(_0838_),
    .X(_0304_));
 sg13g2_nor3_1 _2380_ (.A(net434),
    .B(_0783_),
    .C(_0837_),
    .Y(_0839_));
 sg13g2_a21o_1 _2381_ (.A2(_0836_),
    .A1(net157),
    .B1(_0839_),
    .X(_0305_));
 sg13g2_nor3_1 _2382_ (.A(net434),
    .B(_0787_),
    .C(_0837_),
    .Y(_0840_));
 sg13g2_a21o_1 _2383_ (.A2(_0836_),
    .A1(net160),
    .B1(_0840_),
    .X(_0306_));
 sg13g2_nor3_1 _2384_ (.A(net434),
    .B(_0791_),
    .C(_0837_),
    .Y(_0841_));
 sg13g2_a21o_1 _2385_ (.A2(_0836_),
    .A1(net162),
    .B1(_0841_),
    .X(_0307_));
 sg13g2_nor3_1 _2386_ (.A(net434),
    .B(_0795_),
    .C(_0837_),
    .Y(_0842_));
 sg13g2_a21o_1 _2387_ (.A2(_0836_),
    .A1(net161),
    .B1(_0842_),
    .X(_0308_));
 sg13g2_nor3_1 _2388_ (.A(net434),
    .B(_0799_),
    .C(_0837_),
    .Y(_0843_));
 sg13g2_a21o_1 _2389_ (.A2(_0836_),
    .A1(net194),
    .B1(_0843_),
    .X(_0309_));
 sg13g2_nor3_1 _2390_ (.A(net434),
    .B(_0803_),
    .C(_0837_),
    .Y(_0844_));
 sg13g2_a21o_1 _2391_ (.A2(_0836_),
    .A1(net165),
    .B1(_0844_),
    .X(_0310_));
 sg13g2_nor3_1 _2392_ (.A(net434),
    .B(_0807_),
    .C(_0837_),
    .Y(_0845_));
 sg13g2_a21o_1 _2393_ (.A2(_0836_),
    .A1(net188),
    .B1(_0845_),
    .X(_0311_));
 sg13g2_nand2b_1 _2394_ (.Y(_0846_),
    .B(_0665_),
    .A_N(_0780_));
 sg13g2_nand4_1 _2395_ (.B(_0924_),
    .C(\uart_proj.fifoTx.write_ptr[2] ),
    .A(\uart_proj.fifoTx.write_ptr[0] ),
    .Y(_0847_),
    .D(_0665_));
 sg13g2_nand2_1 _2396_ (.Y(_0848_),
    .A(net132),
    .B(_0847_));
 sg13g2_o21ai_1 _2397_ (.B1(_0848_),
    .Y(_0312_),
    .A1(_0779_),
    .A2(_0846_));
 sg13g2_nand2_1 _2398_ (.Y(_0849_),
    .A(net86),
    .B(_0847_));
 sg13g2_o21ai_1 _2399_ (.B1(_0849_),
    .Y(_0313_),
    .A1(_0785_),
    .A2(net421));
 sg13g2_nand2_1 _2400_ (.Y(_0850_),
    .A(net43),
    .B(_0847_));
 sg13g2_o21ai_1 _2401_ (.B1(_0850_),
    .Y(_0314_),
    .A1(_0789_),
    .A2(net421));
 sg13g2_nand2_1 _2402_ (.Y(_0851_),
    .A(net113),
    .B(_0847_));
 sg13g2_o21ai_1 _2403_ (.B1(_0851_),
    .Y(_0315_),
    .A1(_0793_),
    .A2(net421));
 sg13g2_nand2_1 _2404_ (.Y(_0852_),
    .A(net77),
    .B(_0847_));
 sg13g2_o21ai_1 _2405_ (.B1(_0852_),
    .Y(_0316_),
    .A1(_0797_),
    .A2(net421));
 sg13g2_nand2_1 _2406_ (.Y(_0853_),
    .A(net60),
    .B(_0847_));
 sg13g2_o21ai_1 _2407_ (.B1(_0853_),
    .Y(_0317_),
    .A1(_0801_),
    .A2(net422));
 sg13g2_nand2_1 _2408_ (.Y(_0854_),
    .A(net64),
    .B(_0847_));
 sg13g2_o21ai_1 _2409_ (.B1(_0854_),
    .Y(_0318_),
    .A1(_0805_),
    .A2(net422));
 sg13g2_nand2_1 _2410_ (.Y(_0855_),
    .A(net109),
    .B(_0847_));
 sg13g2_o21ai_1 _2411_ (.B1(_0855_),
    .Y(_0319_),
    .A1(_0809_),
    .A2(net422));
 sg13g2_or3_1 _2412_ (.A(\uart_proj.fifoTx.write_ptr[0] ),
    .B(_0924_),
    .C(net422),
    .X(_0856_));
 sg13g2_nand2_1 _2413_ (.Y(_0857_),
    .A(net59),
    .B(net416));
 sg13g2_o21ai_1 _2414_ (.B1(_0857_),
    .Y(_0320_),
    .A1(_0777_),
    .A2(net416));
 sg13g2_nand2_1 _2415_ (.Y(_0858_),
    .A(net115),
    .B(net416));
 sg13g2_o21ai_1 _2416_ (.B1(_0858_),
    .Y(_0321_),
    .A1(_0783_),
    .A2(net416));
 sg13g2_nand2_1 _2417_ (.Y(_0859_),
    .A(net75),
    .B(net416));
 sg13g2_o21ai_1 _2418_ (.B1(_0859_),
    .Y(_0322_),
    .A1(_0787_),
    .A2(net416));
 sg13g2_nand2_1 _2419_ (.Y(_0860_),
    .A(net50),
    .B(net416));
 sg13g2_o21ai_1 _2420_ (.B1(_0860_),
    .Y(_0323_),
    .A1(_0791_),
    .A2(net416));
 sg13g2_nand2_1 _2421_ (.Y(_0861_),
    .A(net55),
    .B(net415));
 sg13g2_o21ai_1 _2422_ (.B1(_0861_),
    .Y(_0324_),
    .A1(_0795_),
    .A2(net415));
 sg13g2_nand2_1 _2423_ (.Y(_0862_),
    .A(net98),
    .B(net415));
 sg13g2_o21ai_1 _2424_ (.B1(_0862_),
    .Y(_0325_),
    .A1(_0799_),
    .A2(net415));
 sg13g2_nand2_1 _2425_ (.Y(_0863_),
    .A(net63),
    .B(net415));
 sg13g2_o21ai_1 _2426_ (.B1(_0863_),
    .Y(_0326_),
    .A1(_0803_),
    .A2(net415));
 sg13g2_nand2_1 _2427_ (.Y(_0864_),
    .A(net58),
    .B(net415));
 sg13g2_o21ai_1 _2428_ (.B1(_0864_),
    .Y(_0327_),
    .A1(_0807_),
    .A2(net415));
 sg13g2_nand2_1 _2429_ (.Y(_0865_),
    .A(net47),
    .B(_0674_));
 sg13g2_o21ai_1 _2430_ (.B1(net48),
    .Y(_0328_),
    .A1(_0821_),
    .A2(net421));
 sg13g2_nand2_1 _2431_ (.Y(_0866_),
    .A(net81),
    .B(net417));
 sg13g2_o21ai_1 _2432_ (.B1(_0866_),
    .Y(_0329_),
    .A1(_0823_),
    .A2(_0846_));
 sg13g2_nand2_1 _2433_ (.Y(_0867_),
    .A(net56),
    .B(net417));
 sg13g2_o21ai_1 _2434_ (.B1(_0867_),
    .Y(_0330_),
    .A1(_0825_),
    .A2(net421));
 sg13g2_nand2_1 _2435_ (.Y(_0868_),
    .A(net80),
    .B(net417));
 sg13g2_o21ai_1 _2436_ (.B1(_0868_),
    .Y(_0331_),
    .A1(_0827_),
    .A2(net421));
 sg13g2_nand2_1 _2437_ (.Y(_0869_),
    .A(net99),
    .B(net417));
 sg13g2_o21ai_1 _2438_ (.B1(_0869_),
    .Y(_0332_),
    .A1(_0829_),
    .A2(net421));
 sg13g2_nand2_1 _2439_ (.Y(_0870_),
    .A(net67),
    .B(net417));
 sg13g2_o21ai_1 _2440_ (.B1(_0870_),
    .Y(_0333_),
    .A1(_0831_),
    .A2(net422));
 sg13g2_nand2_1 _2441_ (.Y(_0871_),
    .A(net93),
    .B(net417));
 sg13g2_o21ai_1 _2442_ (.B1(_0871_),
    .Y(_0334_),
    .A1(_0833_),
    .A2(net422));
 sg13g2_nand2_1 _2443_ (.Y(_0872_),
    .A(net46),
    .B(net417));
 sg13g2_o21ai_1 _2444_ (.B1(_0872_),
    .Y(_0335_),
    .A1(_0835_),
    .A2(net422));
 sg13g2_nor2_1 _2445_ (.A(net391),
    .B(net407),
    .Y(_0873_));
 sg13g2_a21oi_1 _2446_ (.A1(net407),
    .A2(_1187_),
    .Y(_0336_),
    .B1(_0873_));
 sg13g2_nor2_1 _2447_ (.A(net382),
    .B(net406),
    .Y(_0874_));
 sg13g2_a21oi_1 _2448_ (.A1(net406),
    .A2(_1194_),
    .Y(_0337_),
    .B1(_0874_));
 sg13g2_nor2_1 _2449_ (.A(_1159_),
    .B(_1199_),
    .Y(_0875_));
 sg13g2_a21oi_1 _2450_ (.A1(_0915_),
    .A2(_1159_),
    .Y(_0338_),
    .B1(_0875_));
 sg13g2_mux2_1 _2451_ (.A0(net34),
    .A1(net191),
    .S(net403),
    .X(_0339_));
 sg13g2_mux2_1 _2452_ (.A0(net68),
    .A1(net271),
    .S(_1189_),
    .X(_0340_));
 sg13g2_mux2_1 _2453_ (.A0(net39),
    .A1(net217),
    .S(net403),
    .X(_0341_));
 sg13g2_mux2_1 _2454_ (.A0(net24),
    .A1(net270),
    .S(net403),
    .X(_0342_));
 sg13g2_mux2_1 _2455_ (.A0(net26),
    .A1(net214),
    .S(net403),
    .X(_0343_));
 sg13g2_mux2_1 _2456_ (.A0(net28),
    .A1(net275),
    .S(net403),
    .X(_0344_));
 sg13g2_mux2_1 _2457_ (.A0(net30),
    .A1(net227),
    .S(net403),
    .X(_0345_));
 sg13g2_mux2_1 _2458_ (.A0(net32),
    .A1(net222),
    .S(net403),
    .X(_0346_));
 sg13g2_nor3_2 _2459_ (.A(_1194_),
    .B(_1197_),
    .C(_1198_),
    .Y(_0876_));
 sg13g2_a21o_1 _2460_ (.A2(_0876_),
    .A1(_1175_),
    .B1(_1159_),
    .X(_0877_));
 sg13g2_nand2_1 _2461_ (.Y(_0878_),
    .A(net21),
    .B(_0877_));
 sg13g2_nor2b_1 _2462_ (.A(_1176_),
    .B_N(_0876_),
    .Y(_0879_));
 sg13g2_nand2b_2 _2463_ (.Y(_0880_),
    .B(_0876_),
    .A_N(_1176_));
 sg13g2_o21ai_1 _2464_ (.B1(_0878_),
    .Y(_0347_),
    .A1(net21),
    .A2(_0880_));
 sg13g2_nand2_1 _2465_ (.Y(_0881_),
    .A(\uart_proj.uartRx.readCount[1] ),
    .B(_0877_));
 sg13g2_xor2_1 _2466_ (.B(net21),
    .A(\uart_proj.uartRx.readCount[1] ),
    .X(_0882_));
 sg13g2_o21ai_1 _2467_ (.B1(_0881_),
    .Y(_0348_),
    .A1(_0880_),
    .A2(net22));
 sg13g2_nand2_1 _2468_ (.Y(_0883_),
    .A(net241),
    .B(_0877_));
 sg13g2_o21ai_1 _2469_ (.B1(net241),
    .Y(_0884_),
    .A1(\uart_proj.uartRx.readCount[1] ),
    .A2(net21));
 sg13g2_nor2b_1 _2470_ (.A(_1180_),
    .B_N(_0884_),
    .Y(_0885_));
 sg13g2_o21ai_1 _2471_ (.B1(_0883_),
    .Y(_0349_),
    .A1(_0880_),
    .A2(_0885_));
 sg13g2_nand2_1 _2472_ (.Y(_0886_),
    .A(net44),
    .B(_0877_));
 sg13g2_xor2_1 _2473_ (.B(_1180_),
    .A(\uart_proj.uartRx.readCount[3] ),
    .X(_0887_));
 sg13g2_o21ai_1 _2474_ (.B1(_0886_),
    .Y(_0350_),
    .A1(_0880_),
    .A2(_0887_));
 sg13g2_nand2_1 _2475_ (.Y(_0888_),
    .A(net122),
    .B(_1159_));
 sg13g2_nand2_1 _2476_ (.Y(_0889_),
    .A(\uart_proj.uartRx.sampleCount[0] ),
    .B(_1158_));
 sg13g2_o21ai_1 _2477_ (.B1(_0888_),
    .Y(_0351_),
    .A1(_0771_),
    .A2(_0889_));
 sg13g2_nand2_1 _2478_ (.Y(_0890_),
    .A(net89),
    .B(_1159_));
 sg13g2_nand2_1 _2479_ (.Y(_0891_),
    .A(\uart_proj.uartRx.sampleCount[0] ),
    .B(\uart_proj.uartRx.sampleCount[1] ));
 sg13g2_nand3b_1 _2480_ (.B(_0891_),
    .C(_1158_),
    .Y(_0892_),
    .A_N(_1165_));
 sg13g2_o21ai_1 _2481_ (.B1(_0890_),
    .Y(_0352_),
    .A1(_0771_),
    .A2(_0892_));
 sg13g2_nand2_1 _2482_ (.Y(_0893_),
    .A(net100),
    .B(_1159_));
 sg13g2_o21ai_1 _2483_ (.B1(\uart_proj.uartRx.sampleCount[2] ),
    .Y(_0894_),
    .A1(\uart_proj.uartRx.sampleCount[0] ),
    .A2(\uart_proj.uartRx.sampleCount[1] ));
 sg13g2_nand3_1 _2484_ (.B(_1167_),
    .C(_0894_),
    .A(net407),
    .Y(_0895_));
 sg13g2_o21ai_1 _2485_ (.B1(_0893_),
    .Y(_0353_),
    .A1(_0771_),
    .A2(_0895_));
 sg13g2_nand2_1 _2486_ (.Y(_0896_),
    .A(net65),
    .B(_1159_));
 sg13g2_nand3b_1 _2487_ (.B(net407),
    .C(_1167_),
    .Y(_0897_),
    .A_N(\uart_proj.uartRx.sampleCount[3] ));
 sg13g2_and2_1 _2488_ (.A(_1176_),
    .B(_0897_),
    .X(_0898_));
 sg13g2_o21ai_1 _2489_ (.B1(_0896_),
    .Y(_0354_),
    .A1(_0771_),
    .A2(_0898_));
 sg13g2_mux2_1 _2490_ (.A0(net191),
    .A1(net271),
    .S(net401),
    .X(_0355_));
 sg13g2_mux2_1 _2491_ (.A0(net271),
    .A1(net217),
    .S(_0879_),
    .X(_0356_));
 sg13g2_mux2_1 _2492_ (.A0(net217),
    .A1(net270),
    .S(net401),
    .X(_0357_));
 sg13g2_mux2_1 _2493_ (.A0(net270),
    .A1(net214),
    .S(net401),
    .X(_0358_));
 sg13g2_mux2_1 _2494_ (.A0(net214),
    .A1(net275),
    .S(net401),
    .X(_0359_));
 sg13g2_mux2_1 _2495_ (.A0(net275),
    .A1(net227),
    .S(net401),
    .X(_0360_));
 sg13g2_mux2_1 _2496_ (.A0(net227),
    .A1(net222),
    .S(net401),
    .X(_0361_));
 sg13g2_nor2_1 _2497_ (.A(net222),
    .B(net401),
    .Y(_0899_));
 sg13g2_a21oi_1 _2498_ (.A1(_0900_),
    .A2(net401),
    .Y(_0362_),
    .B1(_0899_));
 sg13g2_buf_1 _2499_ (.A(net3),
    .X(_0162_));
 sg13g2_nor2b_1 _2500_ (.A(net4),
    .B_N(net3),
    .Y(\uart_proj.new_rate[11] ));
 sg13g2_and2_1 _2501_ (.A(net4),
    .B(net3),
    .X(\uart_proj.new_rate[7] ));
 sg13g2_buf_1 _2502_ (.A(net3),
    .X(\uart_proj.new_rate[5] ));
 sg13g2_buf_1 _2503_ (.A(net4),
    .X(\uart_proj.new_rate[8] ));
 sg13g2_dfrbp_1 _2504_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net517),
    .D(_0163_),
    .Q_N(_1341_),
    .Q(\uart_proj.uartTx.writeCount[0] ));
 sg13g2_dfrbp_1 _2505_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net517),
    .D(net281),
    .Q_N(_1340_),
    .Q(\uart_proj.uartTx.writeCount[1] ));
 sg13g2_dfrbp_1 _2506_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net517),
    .D(net283),
    .Q_N(_1339_),
    .Q(\uart_proj.uartTx.writeCount[2] ));
 sg13g2_dfrbp_1 _2507_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net518),
    .D(net119),
    .Q_N(\uart_proj.uartTx.writeCount[3] ),
    .Q(_0146_));
 sg13g2_dfrbp_1 _2508_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net496),
    .D(net19),
    .Q_N(\uart_proj.uartTx.curState[0] ),
    .Q(_0147_));
 sg13g2_dfrbp_1 _2509_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net518),
    .D(net337),
    .Q_N(_1342_),
    .Q(\uart_proj.uartTx.curState[1] ));
 sg13g2_dfrbp_1 _2510_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net518),
    .D(net42),
    .Q_N(_0030_),
    .Q(\uart_proj.uartTx.curState[2] ));
 sg13g2_dfrbp_1 _2511_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net516),
    .D(net352),
    .Q_N(_1338_),
    .Q(\uart_proj.uartTx.curState[3] ));
 sg13g2_dfrbp_1 _2512_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net502),
    .D(net304),
    .Q_N(_1337_),
    .Q(\uart_proj.fifoRx.fifo[0] ));
 sg13g2_dfrbp_1 _2513_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net509),
    .D(net291),
    .Q_N(_1336_),
    .Q(\uart_proj.fifoRx.fifo[1] ));
 sg13g2_dfrbp_1 _2514_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net509),
    .D(net308),
    .Q_N(_1335_),
    .Q(\uart_proj.fifoRx.fifo[2] ));
 sg13g2_dfrbp_1 _2515_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net498),
    .D(net287),
    .Q_N(_1334_),
    .Q(\uart_proj.fifoRx.fifo[3] ));
 sg13g2_dfrbp_1 _2516_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net507),
    .D(net306),
    .Q_N(_1333_),
    .Q(\uart_proj.fifoRx.fifo[4] ));
 sg13g2_dfrbp_1 _2517_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net505),
    .D(net300),
    .Q_N(_1332_),
    .Q(\uart_proj.fifoRx.fifo[5] ));
 sg13g2_dfrbp_1 _2518_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net499),
    .D(net296),
    .Q_N(_1331_),
    .Q(\uart_proj.fifoRx.fifo[6] ));
 sg13g2_dfrbp_1 _2519_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net506),
    .D(net294),
    .Q_N(_1330_),
    .Q(\uart_proj.fifoRx.fifo[7] ));
 sg13g2_dfrbp_1 _2520_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net497),
    .D(net193),
    .Q_N(_1329_),
    .Q(\uart_proj.fifoRx.fifo[8] ));
 sg13g2_dfrbp_1 _2521_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net509),
    .D(net108),
    .Q_N(_1328_),
    .Q(\uart_proj.fifoRx.fifo[9] ));
 sg13g2_dfrbp_1 _2522_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net507),
    .D(net111),
    .Q_N(_1327_),
    .Q(\uart_proj.fifoRx.fifo[10] ));
 sg13g2_dfrbp_1 _2523_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net498),
    .D(net159),
    .Q_N(_1326_),
    .Q(\uart_proj.fifoRx.fifo[11] ));
 sg13g2_dfrbp_1 _2524_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net507),
    .D(net128),
    .Q_N(_1325_),
    .Q(\uart_proj.fifoRx.fifo[12] ));
 sg13g2_dfrbp_1 _2525_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net505),
    .D(net138),
    .Q_N(_1324_),
    .Q(\uart_proj.fifoRx.fifo[13] ));
 sg13g2_dfrbp_1 _2526_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net499),
    .D(net103),
    .Q_N(_1323_),
    .Q(\uart_proj.fifoRx.fifo[14] ));
 sg13g2_dfrbp_1 _2527_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net506),
    .D(net150),
    .Q_N(_1322_),
    .Q(\uart_proj.fifoRx.fifo[15] ));
 sg13g2_dfrbp_1 _2528_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net502),
    .D(net265),
    .Q_N(_1321_),
    .Q(\uart_proj.fifoRx.fifo[16] ));
 sg13g2_dfrbp_1 _2529_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net502),
    .D(net168),
    .Q_N(_1320_),
    .Q(\uart_proj.fifoRx.fifo[17] ));
 sg13g2_dfrbp_1 _2530_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net502),
    .D(net175),
    .Q_N(_1319_),
    .Q(\uart_proj.fifoRx.fifo[18] ));
 sg13g2_dfrbp_1 _2531_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net498),
    .D(net260),
    .Q_N(_1318_),
    .Q(\uart_proj.fifoRx.fifo[19] ));
 sg13g2_dfrbp_1 _2532_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net497),
    .D(net152),
    .Q_N(_1317_),
    .Q(\uart_proj.fifoRx.fifo[20] ));
 sg13g2_dfrbp_1 _2533_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net497),
    .D(net170),
    .Q_N(_1316_),
    .Q(\uart_proj.fifoRx.fifo[21] ));
 sg13g2_dfrbp_1 _2534_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net499),
    .D(net219),
    .Q_N(_1315_),
    .Q(\uart_proj.fifoRx.fifo[22] ));
 sg13g2_dfrbp_1 _2535_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net497),
    .D(net140),
    .Q_N(_1314_),
    .Q(\uart_proj.fifoRx.fifo[23] ));
 sg13g2_dfrbp_1 _2536_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net502),
    .D(net190),
    .Q_N(_1313_),
    .Q(\uart_proj.fifoRx.fifo[24] ));
 sg13g2_dfrbp_1 _2537_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net502),
    .D(net205),
    .Q_N(_1312_),
    .Q(\uart_proj.fifoRx.fifo[25] ));
 sg13g2_dfrbp_1 _2538_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net502),
    .D(net267),
    .Q_N(_1311_),
    .Q(\uart_proj.fifoRx.fifo[26] ));
 sg13g2_dfrbp_1 _2539_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net497),
    .D(net285),
    .Q_N(_1310_),
    .Q(\uart_proj.fifoRx.fifo[27] ));
 sg13g2_dfrbp_1 _2540_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net498),
    .D(net203),
    .Q_N(_1309_),
    .Q(\uart_proj.fifoRx.fifo[28] ));
 sg13g2_dfrbp_1 _2541_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net497),
    .D(net224),
    .Q_N(_1308_),
    .Q(\uart_proj.fifoRx.fifo[29] ));
 sg13g2_dfrbp_1 _2542_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net497),
    .D(net244),
    .Q_N(_1307_),
    .Q(\uart_proj.fifoRx.fifo[30] ));
 sg13g2_dfrbp_1 _2543_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net497),
    .D(net221),
    .Q_N(_1306_),
    .Q(\uart_proj.fifoRx.fifo[31] ));
 sg13g2_dfrbp_1 _2544_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net500),
    .D(_0199_),
    .Q_N(_1305_),
    .Q(\uart_proj.fifoRx.fifo[32] ));
 sg13g2_dfrbp_1 _2545_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net510),
    .D(_0200_),
    .Q_N(_1304_),
    .Q(\uart_proj.fifoRx.fifo[33] ));
 sg13g2_dfrbp_1 _2546_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net506),
    .D(_0201_),
    .Q_N(_1303_),
    .Q(\uart_proj.fifoRx.fifo[34] ));
 sg13g2_dfrbp_1 _2547_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net500),
    .D(_0202_),
    .Q_N(_1302_),
    .Q(\uart_proj.fifoRx.fifo[35] ));
 sg13g2_dfrbp_1 _2548_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net505),
    .D(_0203_),
    .Q_N(_1301_),
    .Q(\uart_proj.fifoRx.fifo[36] ));
 sg13g2_dfrbp_1 _2549_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net505),
    .D(_0204_),
    .Q_N(_1300_),
    .Q(\uart_proj.fifoRx.fifo[37] ));
 sg13g2_dfrbp_1 _2550_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net499),
    .D(_0205_),
    .Q_N(_1299_),
    .Q(\uart_proj.fifoRx.fifo[38] ));
 sg13g2_dfrbp_1 _2551_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net506),
    .D(_0206_),
    .Q_N(_1298_),
    .Q(\uart_proj.fifoRx.fifo[39] ));
 sg13g2_dfrbp_1 _2552_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net500),
    .D(net177),
    .Q_N(_1297_),
    .Q(\uart_proj.fifoRx.fifo[40] ));
 sg13g2_dfrbp_1 _2553_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net510),
    .D(net117),
    .Q_N(_1296_),
    .Q(\uart_proj.fifoRx.fifo[41] ));
 sg13g2_dfrbp_1 _2554_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net506),
    .D(net146),
    .Q_N(_1295_),
    .Q(\uart_proj.fifoRx.fifo[42] ));
 sg13g2_dfrbp_1 _2555_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net499),
    .D(net126),
    .Q_N(_1294_),
    .Q(\uart_proj.fifoRx.fifo[43] ));
 sg13g2_dfrbp_1 _2556_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net507),
    .D(net105),
    .Q_N(_1293_),
    .Q(\uart_proj.fifoRx.fifo[44] ));
 sg13g2_dfrbp_1 _2557_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net505),
    .D(net164),
    .Q_N(_1292_),
    .Q(\uart_proj.fifoRx.fifo[45] ));
 sg13g2_dfrbp_1 _2558_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net499),
    .D(net179),
    .Q_N(_1291_),
    .Q(\uart_proj.fifoRx.fifo[46] ));
 sg13g2_dfrbp_1 _2559_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net506),
    .D(net148),
    .Q_N(_1290_),
    .Q(\uart_proj.fifoRx.fifo[47] ));
 sg13g2_dfrbp_1 _2560_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net503),
    .D(net226),
    .Q_N(_1289_),
    .Q(\uart_proj.fifoRx.fifo[48] ));
 sg13g2_dfrbp_1 _2561_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net503),
    .D(net201),
    .Q_N(_1288_),
    .Q(\uart_proj.fifoRx.fifo[49] ));
 sg13g2_dfrbp_1 _2562_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net509),
    .D(net248),
    .Q_N(_1287_),
    .Q(\uart_proj.fifoRx.fifo[50] ));
 sg13g2_dfrbp_1 _2563_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net500),
    .D(net229),
    .Q_N(_1286_),
    .Q(\uart_proj.fifoRx.fifo[51] ));
 sg13g2_dfrbp_1 _2564_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net508),
    .D(net315),
    .Q_N(_1285_),
    .Q(\uart_proj.fifoRx.fifo[52] ));
 sg13g2_dfrbp_1 _2565_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net505),
    .D(net240),
    .Q_N(_1284_),
    .Q(\uart_proj.fifoRx.fifo[53] ));
 sg13g2_dfrbp_1 _2566_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net499),
    .D(net279),
    .Q_N(_1283_),
    .Q(\uart_proj.fifoRx.fifo[54] ));
 sg13g2_dfrbp_1 _2567_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net506),
    .D(net277),
    .Q_N(_1282_),
    .Q(\uart_proj.fifoRx.fifo[55] ));
 sg13g2_dfrbp_1 _2568_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net503),
    .D(net213),
    .Q_N(_1281_),
    .Q(\uart_proj.fifoRx.fifo[56] ));
 sg13g2_dfrbp_1 _2569_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net503),
    .D(net199),
    .Q_N(_1280_),
    .Q(\uart_proj.fifoRx.fifo[57] ));
 sg13g2_dfrbp_1 _2570_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net509),
    .D(net274),
    .Q_N(_1279_),
    .Q(\uart_proj.fifoRx.fifo[58] ));
 sg13g2_dfrbp_1 _2571_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net500),
    .D(net258),
    .Q_N(_1278_),
    .Q(\uart_proj.fifoRx.fifo[59] ));
 sg13g2_dfrbp_1 _2572_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net505),
    .D(net256),
    .Q_N(_1277_),
    .Q(\uart_proj.fifoRx.fifo[60] ));
 sg13g2_dfrbp_1 _2573_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net505),
    .D(net251),
    .Q_N(_1276_),
    .Q(\uart_proj.fifoRx.fifo[61] ));
 sg13g2_dfrbp_1 _2574_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net499),
    .D(net185),
    .Q_N(_1275_),
    .Q(\uart_proj.fifoRx.fifo[62] ));
 sg13g2_dfrbp_1 _2575_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net506),
    .D(net211),
    .Q_N(_1274_),
    .Q(\uart_proj.fifoRx.fifo[63] ));
 sg13g2_dfrbp_1 _2576_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net495),
    .D(_0159_),
    .Q_N(\uart_proj.bg.rate[2] ),
    .Q(_0148_));
 sg13g2_dfrbp_1 _2577_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net495),
    .D(_0160_),
    .Q_N(\uart_proj.bg.rate[1] ),
    .Q(_0149_));
 sg13g2_dfrbp_1 _2578_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net495),
    .D(\uart_proj.new_rate[5] ),
    .Q_N(_0118_),
    .Q(\uart_proj.bg.rate[5] ));
 sg13g2_dfrbp_1 _2579_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net495),
    .D(_0161_),
    .Q_N(\uart_proj.bg.rate[0] ),
    .Q(_0150_));
 sg13g2_dfrbp_1 _2580_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net495),
    .D(\uart_proj.new_rate[7] ),
    .Q_N(_0116_),
    .Q(\uart_proj.bg.rate[7] ));
 sg13g2_dfrbp_1 _2581_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net493),
    .D(\uart_proj.new_rate[8] ),
    .Q_N(_0115_),
    .Q(\uart_proj.bg.rate[8] ));
 sg13g2_dfrbp_1 _2582_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net493),
    .D(_0162_),
    .Q_N(\uart_proj.bg.rate[10] ),
    .Q(_0151_));
 sg13g2_dfrbp_1 _2583_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net495),
    .D(\uart_proj.new_rate[11] ),
    .Q_N(_0121_),
    .Q(\uart_proj.bg.rate[11] ));
 sg13g2_dfrbp_1 _2584_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net513),
    .D(net530),
    .Q_N(_0037_),
    .Q(\uart_proj.fifoTx.write_ptr[0] ));
 sg13g2_dfrbp_1 _2585_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net503),
    .D(_0232_),
    .Q_N(_1273_),
    .Q(\uart_proj.fifoTx.write_ptr[1] ));
 sg13g2_dfrbp_1 _2586_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net502),
    .D(_0233_),
    .Q_N(_1272_),
    .Q(\uart_proj.fifoTx.write_ptr[2] ));
 sg13g2_dfrbp_1 _2587_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net519),
    .D(_0234_),
    .Q_N(_0035_),
    .Q(\uart_proj.fifoTx.read_ptr[0] ));
 sg13g2_dfrbp_1 _2588_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net520),
    .D(net313),
    .Q_N(_1271_),
    .Q(\uart_proj.fifoTx.read_ptr[1] ));
 sg13g2_dfrbp_1 _2589_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net519),
    .D(_0236_),
    .Q_N(_0036_),
    .Q(\uart_proj.fifoTx.read_ptr[2] ));
 sg13g2_dfrbp_1 _2590_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net511),
    .D(\uart_proj.fifoTx.count_next[0] ),
    .Q_N(_0033_),
    .Q(\uart_proj.fifoTx.count[0] ));
 sg13g2_dfrbp_1 _2591_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net511),
    .D(\uart_proj.fifoTx.count_next[1] ),
    .Q_N(_0034_),
    .Q(\uart_proj.fifoTx.count[1] ));
 sg13g2_dfrbp_1 _2592_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net510),
    .D(\uart_proj.fifoTx.count_next[2] ),
    .Q_N(_1343_),
    .Q(\uart_proj.fifoTx.count[2] ));
 sg13g2_dfrbp_1 _2593_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net520),
    .D(net543),
    .Q_N(_1270_),
    .Q(\uart_proj.fifoTx.count[3] ));
 sg13g2_dfrbp_1 _2594_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net504),
    .D(_0237_),
    .Q_N(_1269_),
    .Q(\uart_proj.fifoRx.overrun ));
 sg13g2_dfrbp_1 _2595_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net503),
    .D(net38),
    .Q_N(_0040_),
    .Q(\uart_proj.fifoRx.write_ptr[0] ));
 sg13g2_dfrbp_1 _2596_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net503),
    .D(net553),
    .Q_N(_1268_),
    .Q(\uart_proj.fifoRx.write_ptr[1] ));
 sg13g2_dfrbp_1 _2597_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net503),
    .D(net346),
    .Q_N(_1267_),
    .Q(\uart_proj.fifoRx.write_ptr[2] ));
 sg13g2_dfrbp_1 _2598_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net509),
    .D(_0241_),
    .Q_N(_1266_),
    .Q(\uart_proj.fifoRx.read_ptr[0] ));
 sg13g2_dfrbp_1 _2599_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net509),
    .D(_0242_),
    .Q_N(_1265_),
    .Q(\uart_proj.fifoRx.read_ptr[1] ));
 sg13g2_dfrbp_1 _2600_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net509),
    .D(_0243_),
    .Q_N(_0039_),
    .Q(\uart_proj.fifoRx.read_ptr[2] ));
 sg13g2_dfrbp_1 _2601_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net493),
    .D(net364),
    .Q_N(_1264_),
    .Q(\uart_proj.bg.rxCount[0] ));
 sg13g2_dfrbp_1 _2602_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net489),
    .D(_0245_),
    .Q_N(_1263_),
    .Q(\uart_proj.bg.rxCount[1] ));
 sg13g2_dfrbp_1 _2603_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net489),
    .D(net334),
    .Q_N(_1262_),
    .Q(\uart_proj.bg.rxCount[2] ));
 sg13g2_dfrbp_1 _2604_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net489),
    .D(_0247_),
    .Q_N(_1261_),
    .Q(\uart_proj.bg.rxCount[3] ));
 sg13g2_dfrbp_1 _2605_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net489),
    .D(_0248_),
    .Q_N(_1260_),
    .Q(\uart_proj.bg.rxCount[4] ));
 sg13g2_dfrbp_1 _2606_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net489),
    .D(_0249_),
    .Q_N(_1259_),
    .Q(\uart_proj.bg.rxCount[5] ));
 sg13g2_dfrbp_1 _2607_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net488),
    .D(_0250_),
    .Q_N(_1258_),
    .Q(\uart_proj.bg.rxCount[6] ));
 sg13g2_dfrbp_1 _2608_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net488),
    .D(_0251_),
    .Q_N(_1257_),
    .Q(\uart_proj.bg.rxCount[7] ));
 sg13g2_dfrbp_1 _2609_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net488),
    .D(_0252_),
    .Q_N(_1256_),
    .Q(\uart_proj.bg.rxCount[8] ));
 sg13g2_dfrbp_1 _2610_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net488),
    .D(_0253_),
    .Q_N(_1255_),
    .Q(\uart_proj.bg.rxCount[9] ));
 sg13g2_dfrbp_1 _2611_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net488),
    .D(net322),
    .Q_N(_1254_),
    .Q(\uart_proj.bg.rxCount[10] ));
 sg13g2_dfrbp_1 _2612_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net487),
    .D(net144),
    .Q_N(_1253_),
    .Q(\uart_proj.bg.rxCount[11] ));
 sg13g2_dfrbp_1 _2613_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net487),
    .D(net263),
    .Q_N(_1252_),
    .Q(\uart_proj.bg.rxCount[12] ));
 sg13g2_dfrbp_1 _2614_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net487),
    .D(_0257_),
    .Q_N(_1251_),
    .Q(\uart_proj.bg.rxCount[13] ));
 sg13g2_dfrbp_1 _2615_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net487),
    .D(_0258_),
    .Q_N(_1250_),
    .Q(\uart_proj.bg.rxCount[14] ));
 sg13g2_dfrbp_1 _2616_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net487),
    .D(net95),
    .Q_N(_1344_),
    .Q(\uart_proj.bg.rxCount[15] ));
 sg13g2_dfrbp_1 _2617_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net510),
    .D(net534),
    .Q_N(_1345_),
    .Q(\uart_proj.fifoRx.count[0] ));
 sg13g2_dfrbp_1 _2618_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net510),
    .D(\uart_proj.fifoRx.count_next[1] ),
    .Q_N(_0038_),
    .Q(\uart_proj.fifoRx.count[1] ));
 sg13g2_dfrbp_1 _2619_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net510),
    .D(\uart_proj.fifoRx.count_next[2] ),
    .Q_N(_1346_),
    .Q(\uart_proj.fifoRx.count[2] ));
 sg13g2_dfrbp_1 _2620_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net510),
    .D(net400),
    .Q_N(_1347_),
    .Q(\uart_proj.fifoRx.count[3] ));
 sg13g2_dfrbp_1 _2621_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net516),
    .D(net348),
    .Q_N(_1348_),
    .Q(_0026_));
 sg13g2_dfrbp_1 _2622_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net516),
    .D(_0025_),
    .Q_N(_1249_),
    .Q(_0027_));
 sg13g2_dfrbp_1 _2623_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net522),
    .D(net233),
    .Q_N(_1248_),
    .Q(\uart_proj.uartTx.writeBuf[0] ));
 sg13g2_dfrbp_1 _2624_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net522),
    .D(net131),
    .Q_N(_1247_),
    .Q(\uart_proj.uartTx.writeBuf[1] ));
 sg13g2_dfrbp_1 _2625_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net524),
    .D(net156),
    .Q_N(_1246_),
    .Q(\uart_proj.uartTx.writeBuf[2] ));
 sg13g2_dfrbp_1 _2626_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net524),
    .D(net235),
    .Q_N(_1245_),
    .Q(\uart_proj.uartTx.writeBuf[3] ));
 sg13g2_dfrbp_1 _2627_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net524),
    .D(net187),
    .Q_N(_1244_),
    .Q(\uart_proj.uartTx.writeBuf[4] ));
 sg13g2_dfrbp_1 _2628_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net524),
    .D(net183),
    .Q_N(_1243_),
    .Q(\uart_proj.uartTx.writeBuf[5] ));
 sg13g2_dfrbp_1 _2629_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net524),
    .D(net97),
    .Q_N(_1242_),
    .Q(\uart_proj.uartTx.writeBuf[6] ));
 sg13g2_dfrbp_1 _2630_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net521),
    .D(_0267_),
    .Q_N(_1241_),
    .Q(\uart_proj.uartTx.writeBuf[7] ));
 sg13g2_dfrbp_1 _2631_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net494),
    .D(_0268_),
    .Q_N(\uart_proj.uartRx.cmp ),
    .Q(_0152_));
 sg13g2_dfrbp_1 _2632_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net518),
    .D(net237),
    .Q_N(_1240_),
    .Q(\uart_proj.uartTx.hasData ));
 sg13g2_dfrbp_1 _2633_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net516),
    .D(_0270_),
    .Q_N(_1239_),
    .Q(\uart_proj.uartTx.enterStart ));
 sg13g2_dfrbp_1 _2634_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net493),
    .D(net216),
    .Q_N(_1238_),
    .Q(\uart_proj.uartRx.edgeCmp ));
 sg13g2_dfrbp_1 _2635_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net523),
    .D(_0272_),
    .Q_N(_0041_),
    .Q(\uart_proj.fifoTx.fifo[0] ));
 sg13g2_dfrbp_1 _2636_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net523),
    .D(_0273_),
    .Q_N(_0049_),
    .Q(\uart_proj.fifoTx.fifo[1] ));
 sg13g2_dfrbp_1 _2637_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net523),
    .D(_0274_),
    .Q_N(_0057_),
    .Q(\uart_proj.fifoTx.fifo[2] ));
 sg13g2_dfrbp_1 _2638_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net520),
    .D(_0275_),
    .Q_N(_0065_),
    .Q(\uart_proj.fifoTx.fifo[3] ));
 sg13g2_dfrbp_1 _2639_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net520),
    .D(_0276_),
    .Q_N(_0073_),
    .Q(\uart_proj.fifoTx.fifo[4] ));
 sg13g2_dfrbp_1 _2640_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net520),
    .D(_0277_),
    .Q_N(_0081_),
    .Q(\uart_proj.fifoTx.fifo[5] ));
 sg13g2_dfrbp_1 _2641_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net520),
    .D(_0278_),
    .Q_N(_0089_),
    .Q(\uart_proj.fifoTx.fifo[6] ));
 sg13g2_dfrbp_1 _2642_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net519),
    .D(_0279_),
    .Q_N(_0097_),
    .Q(\uart_proj.fifoTx.fifo[7] ));
 sg13g2_dfrbp_1 _2643_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net517),
    .D(net71),
    .Q_N(_0042_),
    .Q(\uart_proj.fifoTx.fifo[8] ));
 sg13g2_dfrbp_1 _2644_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net517),
    .D(net92),
    .Q_N(_0050_),
    .Q(\uart_proj.fifoTx.fifo[9] ));
 sg13g2_dfrbp_1 _2645_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net517),
    .D(_0282_),
    .Q_N(_0058_),
    .Q(\uart_proj.fifoTx.fifo[10] ));
 sg13g2_dfrbp_1 _2646_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net514),
    .D(_0283_),
    .Q_N(_0066_),
    .Q(\uart_proj.fifoTx.fifo[11] ));
 sg13g2_dfrbp_1 _2647_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net513),
    .D(_0284_),
    .Q_N(_0074_),
    .Q(\uart_proj.fifoTx.fifo[12] ));
 sg13g2_dfrbp_1 _2648_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net513),
    .D(_0285_),
    .Q_N(_0082_),
    .Q(\uart_proj.fifoTx.fifo[13] ));
 sg13g2_dfrbp_1 _2649_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net513),
    .D(_0286_),
    .Q_N(_0090_),
    .Q(\uart_proj.fifoTx.fifo[14] ));
 sg13g2_dfrbp_1 _2650_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net513),
    .D(_0287_),
    .Q_N(_0098_),
    .Q(\uart_proj.fifoTx.fifo[15] ));
 sg13g2_dfrbp_1 _2651_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net521),
    .D(_0288_),
    .Q_N(_0043_),
    .Q(\uart_proj.fifoTx.fifo[16] ));
 sg13g2_dfrbp_1 _2652_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net521),
    .D(_0289_),
    .Q_N(_0051_),
    .Q(\uart_proj.fifoTx.fifo[17] ));
 sg13g2_dfrbp_1 _2653_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net523),
    .D(_0290_),
    .Q_N(_0059_),
    .Q(\uart_proj.fifoTx.fifo[18] ));
 sg13g2_dfrbp_1 _2654_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net521),
    .D(_0291_),
    .Q_N(_0067_),
    .Q(\uart_proj.fifoTx.fifo[19] ));
 sg13g2_dfrbp_1 _2655_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net519),
    .D(_0292_),
    .Q_N(_0075_),
    .Q(\uart_proj.fifoTx.fifo[20] ));
 sg13g2_dfrbp_1 _2656_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net519),
    .D(_0293_),
    .Q_N(_0083_),
    .Q(\uart_proj.fifoTx.fifo[21] ));
 sg13g2_dfrbp_1 _2657_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net519),
    .D(_0294_),
    .Q_N(_0091_),
    .Q(\uart_proj.fifoTx.fifo[22] ));
 sg13g2_dfrbp_1 _2658_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net519),
    .D(_0295_),
    .Q_N(_0099_),
    .Q(\uart_proj.fifoTx.fifo[23] ));
 sg13g2_dfrbp_1 _2659_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net517),
    .D(net85),
    .Q_N(_0044_),
    .Q(\uart_proj.fifoTx.fifo[24] ));
 sg13g2_dfrbp_1 _2660_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net517),
    .D(net53),
    .Q_N(_0052_),
    .Q(\uart_proj.fifoTx.fifo[25] ));
 sg13g2_dfrbp_1 _2661_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net521),
    .D(_0298_),
    .Q_N(_0060_),
    .Q(\uart_proj.fifoTx.fifo[26] ));
 sg13g2_dfrbp_1 _2662_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net521),
    .D(_0299_),
    .Q_N(_0068_),
    .Q(\uart_proj.fifoTx.fifo[27] ));
 sg13g2_dfrbp_1 _2663_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net519),
    .D(_0300_),
    .Q_N(_0076_),
    .Q(\uart_proj.fifoTx.fifo[28] ));
 sg13g2_dfrbp_1 _2664_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net513),
    .D(_0301_),
    .Q_N(_0084_),
    .Q(\uart_proj.fifoTx.fifo[29] ));
 sg13g2_dfrbp_1 _2665_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net513),
    .D(_0302_),
    .Q_N(_0092_),
    .Q(\uart_proj.fifoTx.fifo[30] ));
 sg13g2_dfrbp_1 _2666_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net513),
    .D(_0303_),
    .Q_N(_0100_),
    .Q(\uart_proj.fifoTx.fifo[31] ));
 sg13g2_dfrbp_1 _2667_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net515),
    .D(_0304_),
    .Q_N(_0045_),
    .Q(\uart_proj.fifoTx.fifo[32] ));
 sg13g2_dfrbp_1 _2668_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net495),
    .D(_0305_),
    .Q_N(_0053_),
    .Q(\uart_proj.fifoTx.fifo[33] ));
 sg13g2_dfrbp_1 _2669_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net495),
    .D(_0306_),
    .Q_N(_0061_),
    .Q(\uart_proj.fifoTx.fifo[34] ));
 sg13g2_dfrbp_1 _2670_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net494),
    .D(_0307_),
    .Q_N(_0069_),
    .Q(\uart_proj.fifoTx.fifo[35] ));
 sg13g2_dfrbp_1 _2671_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net494),
    .D(_0308_),
    .Q_N(_0077_),
    .Q(\uart_proj.fifoTx.fifo[36] ));
 sg13g2_dfrbp_1 _2672_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net512),
    .D(_0309_),
    .Q_N(_0085_),
    .Q(\uart_proj.fifoTx.fifo[37] ));
 sg13g2_dfrbp_1 _2673_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net493),
    .D(_0310_),
    .Q_N(_0093_),
    .Q(\uart_proj.fifoTx.fifo[38] ));
 sg13g2_dfrbp_1 _2674_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net493),
    .D(_0311_),
    .Q_N(_0101_),
    .Q(\uart_proj.fifoTx.fifo[39] ));
 sg13g2_dfrbp_1 _2675_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net516),
    .D(net133),
    .Q_N(_0046_),
    .Q(\uart_proj.fifoTx.fifo[40] ));
 sg13g2_dfrbp_1 _2676_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net515),
    .D(net87),
    .Q_N(_0054_),
    .Q(\uart_proj.fifoTx.fifo[41] ));
 sg13g2_dfrbp_1 _2677_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net496),
    .D(_0314_),
    .Q_N(_0062_),
    .Q(\uart_proj.fifoTx.fifo[42] ));
 sg13g2_dfrbp_1 _2678_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net494),
    .D(_0315_),
    .Q_N(_0070_),
    .Q(\uart_proj.fifoTx.fifo[43] ));
 sg13g2_dfrbp_1 _2679_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net494),
    .D(_0316_),
    .Q_N(_0078_),
    .Q(\uart_proj.fifoTx.fifo[44] ));
 sg13g2_dfrbp_1 _2680_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net512),
    .D(_0317_),
    .Q_N(_0086_),
    .Q(\uart_proj.fifoTx.fifo[45] ));
 sg13g2_dfrbp_1 _2681_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net512),
    .D(_0318_),
    .Q_N(_0094_),
    .Q(\uart_proj.fifoTx.fifo[46] ));
 sg13g2_dfrbp_1 _2682_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net493),
    .D(_0319_),
    .Q_N(_0102_),
    .Q(\uart_proj.fifoTx.fifo[47] ));
 sg13g2_dfrbp_1 _2683_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net516),
    .D(_0320_),
    .Q_N(_0047_),
    .Q(\uart_proj.fifoTx.fifo[48] ));
 sg13g2_dfrbp_1 _2684_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net516),
    .D(_0321_),
    .Q_N(_0055_),
    .Q(\uart_proj.fifoTx.fifo[49] ));
 sg13g2_dfrbp_1 _2685_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net515),
    .D(_0322_),
    .Q_N(_0063_),
    .Q(\uart_proj.fifoTx.fifo[50] ));
 sg13g2_dfrbp_1 _2686_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net515),
    .D(_0323_),
    .Q_N(_0071_),
    .Q(\uart_proj.fifoTx.fifo[51] ));
 sg13g2_dfrbp_1 _2687_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net512),
    .D(_0324_),
    .Q_N(_0079_),
    .Q(\uart_proj.fifoTx.fifo[52] ));
 sg13g2_dfrbp_1 _2688_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net512),
    .D(_0325_),
    .Q_N(_0087_),
    .Q(\uart_proj.fifoTx.fifo[53] ));
 sg13g2_dfrbp_1 _2689_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net512),
    .D(_0326_),
    .Q_N(_0095_),
    .Q(\uart_proj.fifoTx.fifo[54] ));
 sg13g2_dfrbp_1 _2690_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net514),
    .D(_0327_),
    .Q_N(_0103_),
    .Q(\uart_proj.fifoTx.fifo[55] ));
 sg13g2_dfrbp_1 _2691_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net515),
    .D(net49),
    .Q_N(_0048_),
    .Q(\uart_proj.fifoTx.fifo[56] ));
 sg13g2_dfrbp_1 _2692_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net515),
    .D(net82),
    .Q_N(_0056_),
    .Q(\uart_proj.fifoTx.fifo[57] ));
 sg13g2_dfrbp_1 _2693_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net515),
    .D(_0330_),
    .Q_N(_0064_),
    .Q(\uart_proj.fifoTx.fifo[58] ));
 sg13g2_dfrbp_1 _2694_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net515),
    .D(_0331_),
    .Q_N(_0072_),
    .Q(\uart_proj.fifoTx.fifo[59] ));
 sg13g2_dfrbp_1 _2695_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net512),
    .D(_0332_),
    .Q_N(_0080_),
    .Q(\uart_proj.fifoTx.fifo[60] ));
 sg13g2_dfrbp_1 _2696_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net512),
    .D(_0333_),
    .Q_N(_0088_),
    .Q(\uart_proj.fifoTx.fifo[61] ));
 sg13g2_dfrbp_1 _2697_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net514),
    .D(_0334_),
    .Q_N(_0096_),
    .Q(\uart_proj.fifoTx.fifo[62] ));
 sg13g2_dfrbp_1 _2698_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net514),
    .D(_0335_),
    .Q_N(_0104_),
    .Q(\uart_proj.fifoTx.fifo[63] ));
 sg13g2_dfrbp_1 _2699_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net493),
    .D(_0336_),
    .Q_N(_1237_),
    .Q(\uart_proj.uartRx.curState[0] ));
 sg13g2_dfrbp_1 _2700_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net484),
    .D(_0337_),
    .Q_N(_0028_),
    .Q(\uart_proj.uartRx.curState[1] ));
 sg13g2_dfrbp_1 _2701_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net484),
    .D(_0338_),
    .Q_N(_0029_),
    .Q(\uart_proj.uartRx.curState[2] ));
 sg13g2_dfrbp_1 _2702_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net485),
    .D(_0339_),
    .Q_N(_1236_),
    .Q(\uart_proj.rxData[0] ));
 sg13g2_dfrbp_1 _2703_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net485),
    .D(net272),
    .Q_N(_1235_),
    .Q(\uart_proj.rxData[1] ));
 sg13g2_dfrbp_1 _2704_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net483),
    .D(_0341_),
    .Q_N(_1234_),
    .Q(\uart_proj.rxData[2] ));
 sg13g2_dfrbp_1 _2705_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net483),
    .D(_0342_),
    .Q_N(_1233_),
    .Q(\uart_proj.rxData[3] ));
 sg13g2_dfrbp_1 _2706_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net483),
    .D(_0343_),
    .Q_N(_1232_),
    .Q(\uart_proj.rxData[4] ));
 sg13g2_dfrbp_1 _2707_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net482),
    .D(_0344_),
    .Q_N(_1231_),
    .Q(\uart_proj.rxData[5] ));
 sg13g2_dfrbp_1 _2708_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net482),
    .D(_0345_),
    .Q_N(_1230_),
    .Q(\uart_proj.rxData[6] ));
 sg13g2_dfrbp_1 _2709_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net482),
    .D(_0346_),
    .Q_N(_1229_),
    .Q(\uart_proj.rxData[7] ));
 sg13g2_dfrbp_1 _2710_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net487),
    .D(_0347_),
    .Q_N(_1228_),
    .Q(\uart_proj.uartRx.readCount[0] ));
 sg13g2_dfrbp_1 _2711_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net487),
    .D(net23),
    .Q_N(_1227_),
    .Q(\uart_proj.uartRx.readCount[1] ));
 sg13g2_dfrbp_1 _2712_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net484),
    .D(net242),
    .Q_N(_1226_),
    .Q(\uart_proj.uartRx.readCount[2] ));
 sg13g2_dfrbp_1 _2713_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net484),
    .D(net45),
    .Q_N(\uart_proj.uartRx.readCount[3] ),
    .Q(_0153_));
 sg13g2_dfrbp_1 _2714_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net485),
    .D(net123),
    .Q_N(\uart_proj.uartRx.sampleCount[0] ),
    .Q(_0154_));
 sg13g2_dfrbp_1 _2715_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net485),
    .D(net90),
    .Q_N(\uart_proj.uartRx.sampleCount[1] ),
    .Q(_0155_));
 sg13g2_dfrbp_1 _2716_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net485),
    .D(net101),
    .Q_N(\uart_proj.uartRx.sampleCount[2] ),
    .Q(_0156_));
 sg13g2_dfrbp_1 _2717_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net484),
    .D(net66),
    .Q_N(\uart_proj.uartRx.sampleCount[3] ),
    .Q(_0157_));
 sg13g2_dfrbp_1 _2718_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net484),
    .D(_0355_),
    .Q_N(_1225_),
    .Q(\uart_proj.uartRx.readBuf[0] ));
 sg13g2_dfrbp_1 _2719_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net484),
    .D(_0356_),
    .Q_N(_1224_),
    .Q(\uart_proj.uartRx.readBuf[1] ));
 sg13g2_dfrbp_1 _2720_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net482),
    .D(_0357_),
    .Q_N(_1223_),
    .Q(\uart_proj.uartRx.readBuf[2] ));
 sg13g2_dfrbp_1 _2721_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net482),
    .D(_0358_),
    .Q_N(_1222_),
    .Q(\uart_proj.uartRx.readBuf[3] ));
 sg13g2_dfrbp_1 _2722_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net482),
    .D(_0359_),
    .Q_N(_1221_),
    .Q(\uart_proj.uartRx.readBuf[4] ));
 sg13g2_dfrbp_1 _2723_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net482),
    .D(_0360_),
    .Q_N(_1220_),
    .Q(\uart_proj.uartRx.readBuf[5] ));
 sg13g2_dfrbp_1 _2724_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net482),
    .D(_0361_),
    .Q_N(_1219_),
    .Q(\uart_proj.uartRx.readBuf[6] ));
 sg13g2_dfrbp_1 _2725_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net484),
    .D(_0362_),
    .Q_N(_1349_),
    .Q(\uart_proj.uartRx.readBuf[7] ));
 sg13g2_dfrbp_1 _2726_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net492),
    .D(_0126_),
    .Q_N(_0123_),
    .Q(\uart_proj.bg.txCount[0] ));
 sg13g2_dfrbp_1 _2727_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net491),
    .D(_0137_),
    .Q_N(_1350_),
    .Q(\uart_proj.bg.txCount[1] ));
 sg13g2_dfrbp_1 _2728_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net491),
    .D(_0138_),
    .Q_N(_0122_),
    .Q(\uart_proj.bg.txCount[2] ));
 sg13g2_dfrbp_1 _2729_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net492),
    .D(_0139_),
    .Q_N(_1351_),
    .Q(\uart_proj.bg.txCount[3] ));
 sg13g2_dfrbp_1 _2730_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net491),
    .D(net354),
    .Q_N(_0120_),
    .Q(\uart_proj.bg.txCount[4] ));
 sg13g2_dfrbp_1 _2731_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net491),
    .D(_0141_),
    .Q_N(_0119_),
    .Q(\uart_proj.bg.txCount[5] ));
 sg13g2_dfrbp_1 _2732_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net491),
    .D(_0142_),
    .Q_N(_0117_),
    .Q(\uart_proj.bg.txCount[6] ));
 sg13g2_dfrbp_1 _2733_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net491),
    .D(_0143_),
    .Q_N(_1352_),
    .Q(\uart_proj.bg.txCount[7] ));
 sg13g2_dfrbp_1 _2734_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net491),
    .D(net397),
    .Q_N(_0114_),
    .Q(\uart_proj.bg.txCount[8] ));
 sg13g2_dfrbp_1 _2735_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net491),
    .D(_0145_),
    .Q_N(_0113_),
    .Q(\uart_proj.bg.txCount[9] ));
 sg13g2_dfrbp_1 _2736_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net490),
    .D(net384),
    .Q_N(_0112_),
    .Q(\uart_proj.bg.txCount[10] ));
 sg13g2_dfrbp_1 _2737_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net490),
    .D(_0128_),
    .Q_N(_0111_),
    .Q(\uart_proj.bg.txCount[11] ));
 sg13g2_dfrbp_1 _2738_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net490),
    .D(net540),
    .Q_N(_0125_),
    .Q(\uart_proj.bg.txCount[12] ));
 sg13g2_dfrbp_1 _2739_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net488),
    .D(_0130_),
    .Q_N(_0110_),
    .Q(\uart_proj.bg.txCount[13] ));
 sg13g2_dfrbp_1 _2740_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net488),
    .D(net324),
    .Q_N(_0109_),
    .Q(\uart_proj.bg.txCount[14] ));
 sg13g2_dfrbp_1 _2741_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net488),
    .D(net344),
    .Q_N(_0108_),
    .Q(\uart_proj.bg.txCount[15] ));
 sg13g2_dfrbp_1 _2742_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net490),
    .D(net341),
    .Q_N(_0124_),
    .Q(\uart_proj.bg.txCount[16] ));
 sg13g2_dfrbp_1 _2743_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net489),
    .D(net326),
    .Q_N(_0107_),
    .Q(\uart_proj.bg.txCount[17] ));
 sg13g2_dfrbp_1 _2744_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net489),
    .D(net339),
    .Q_N(_0106_),
    .Q(\uart_proj.bg.txCount[18] ));
 sg13g2_dfrbp_1 _2745_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net489),
    .D(net328),
    .Q_N(_0105_),
    .Q(\uart_proj.bg.txCount[19] ));
 sg13g2_dfrbp_1 _2746_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net485),
    .D(net35),
    .Q_N(_1353_),
    .Q(\uart_proj.fifoRx.wdata[0] ));
 sg13g2_dfrbp_1 _2747_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net485),
    .D(net69),
    .Q_N(_1354_),
    .Q(\uart_proj.fifoRx.wdata[1] ));
 sg13g2_dfrbp_1 _2748_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net485),
    .D(net40),
    .Q_N(_1355_),
    .Q(\uart_proj.fifoRx.wdata[2] ));
 sg13g2_dfrbp_1 _2749_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net483),
    .D(net25),
    .Q_N(_1356_),
    .Q(\uart_proj.fifoRx.wdata[3] ));
 sg13g2_dfrbp_1 _2750_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net483),
    .D(net27),
    .Q_N(_1357_),
    .Q(\uart_proj.fifoRx.wdata[4] ));
 sg13g2_dfrbp_1 _2751_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net483),
    .D(net29),
    .Q_N(_1358_),
    .Q(\uart_proj.fifoRx.wdata[5] ));
 sg13g2_dfrbp_1 _2752_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net483),
    .D(net31),
    .Q_N(_1359_),
    .Q(\uart_proj.fifoRx.wdata[6] ));
 sg13g2_dfrbp_1 _2753_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net483),
    .D(net33),
    .Q_N(_1360_),
    .Q(\uart_proj.fifoRx.wdata[7] ));
 sg13g2_dfrbp_1 _2754_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net504),
    .D(net136),
    .Q_N(_0032_),
    .Q(\uart_proj.fifoRx.WEN ));
 sg13g2_dfrbp_1 _2755_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net520),
    .D(_0014_),
    .Q_N(_1361_),
    .Q(\uart_proj.ren_wen_nidle[0] ));
 sg13g2_dfrbp_1 _2756_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net520),
    .D(_0015_),
    .Q_N(_1362_),
    .Q(\uart_proj.ren_wen_nidle[1] ));
 sg13g2_dfrbp_1 _2757_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net523),
    .D(_0013_),
    .Q_N(_0031_),
    .Q(\uart_proj.fifoTx.REN ));
 sg13g2_dfrbp_1 _2758_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net522),
    .D(net362),
    .Q_N(_1363_),
    .Q(\uart_proj.txData[0] ));
 sg13g2_dfrbp_1 _2759_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net522),
    .D(net368),
    .Q_N(_1364_),
    .Q(\uart_proj.txData[1] ));
 sg13g2_dfrbp_1 _2760_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net524),
    .D(net390),
    .Q_N(_1365_),
    .Q(\uart_proj.txData[2] ));
 sg13g2_dfrbp_1 _2761_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net524),
    .D(net381),
    .Q_N(_1366_),
    .Q(\uart_proj.txData[3] ));
 sg13g2_dfrbp_1 _2762_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net523),
    .D(net395),
    .Q_N(_1367_),
    .Q(\uart_proj.txData[4] ));
 sg13g2_dfrbp_1 _2763_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net524),
    .D(_0021_),
    .Q_N(_1368_),
    .Q(\uart_proj.txData[5] ));
 sg13g2_dfrbp_1 _2764_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net521),
    .D(net358),
    .Q_N(_1369_),
    .Q(\uart_proj.txData[6] ));
 sg13g2_dfrbp_1 _2765_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net521),
    .D(net376),
    .Q_N(_1370_),
    .Q(\uart_proj.txData[7] ));
 sg13g2_dfrbp_1 _2766_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net504),
    .D(_0003_),
    .Q_N(_1371_),
    .Q(\uart_proj.err ));
 sg13g2_dfrbp_1 _2767_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net523),
    .D(net5),
    .Q_N(_1372_),
    .Q(\uart_proj.prev_ren_wen[0] ));
 sg13g2_dfrbp_1 _2768_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net523),
    .D(net6),
    .Q_N(_1218_),
    .Q(\uart_proj.prev_ren_wen[1] ));
 sg13g2_tielo tt_um_purdue_socet_uart_16 (.L_LO(net16));
 sg13g2_tielo tt_um_purdue_socet_uart_17 (.L_LO(net17));
 sg13g2_buf_2 clkbuf_leaf_0_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_buf_1 _2772_ (.A(uio_oe[7]),
    .X(uio_oe[0]));
 sg13g2_buf_1 _2773_ (.A(uio_oe[7]),
    .X(uio_oe[1]));
 sg13g2_buf_1 _2774_ (.A(uio_oe[7]),
    .X(uio_oe[2]));
 sg13g2_buf_1 _2775_ (.A(uio_oe[7]),
    .X(uio_oe[3]));
 sg13g2_buf_1 _2776_ (.A(uio_oe[7]),
    .X(uio_oe[4]));
 sg13g2_buf_1 _2777_ (.A(uio_oe[7]),
    .X(uio_oe[5]));
 sg13g2_buf_1 _2778_ (.A(uio_oe[7]),
    .X(uio_oe[6]));
 sg13g2_buf_2 _2779_ (.A(\uart_proj.tx ),
    .X(uo_out[0]));
 sg13g2_buf_2 _2780_ (.A(\uart_proj.fifoRx.full ),
    .X(uo_out[1]));
 sg13g2_buf_2 _2781_ (.A(\uart_proj.err ),
    .X(uo_out[2]));
 sg13g2_buf_1 _2782_ (.A(\uart_proj.fifoTx.full ),
    .X(uo_out[3]));
 sg13g2_buf_2 _2783_ (.A(\uart_proj.fifoRx.empty ),
    .X(uo_out[4]));
 sg13g2_buf_4 fanout401 (.X(net401),
    .A(_0879_));
 sg13g2_buf_2 fanout402 (.A(_0004_),
    .X(net402));
 sg13g2_buf_4 fanout403 (.X(net403),
    .A(_1189_));
 sg13g2_buf_2 fanout404 (.A(net405),
    .X(net404));
 sg13g2_buf_2 fanout405 (.A(_0697_),
    .X(net405));
 sg13g2_buf_2 fanout406 (.A(net407),
    .X(net406));
 sg13g2_buf_2 fanout407 (.A(_1158_),
    .X(net407));
 sg13g2_buf_2 fanout408 (.A(net409),
    .X(net408));
 sg13g2_buf_1 fanout409 (.A(net410),
    .X(net409));
 sg13g2_buf_2 fanout410 (.A(_0603_),
    .X(net410));
 sg13g2_buf_2 fanout411 (.A(_0411_),
    .X(net411));
 sg13g2_buf_2 fanout412 (.A(net414),
    .X(net412));
 sg13g2_buf_1 fanout413 (.A(net414),
    .X(net413));
 sg13g2_buf_2 fanout414 (.A(_0407_),
    .X(net414));
 sg13g2_buf_2 fanout415 (.A(_0856_),
    .X(net415));
 sg13g2_buf_2 fanout416 (.A(_0856_),
    .X(net416));
 sg13g2_buf_2 fanout417 (.A(_0674_),
    .X(net417));
 sg13g2_buf_4 fanout418 (.X(net418),
    .A(_0642_));
 sg13g2_buf_4 fanout419 (.X(net419),
    .A(_0614_));
 sg13g2_buf_2 fanout420 (.A(_0614_),
    .X(net420));
 sg13g2_buf_4 fanout421 (.X(net421),
    .A(net422));
 sg13g2_buf_4 fanout422 (.X(net422),
    .A(_0846_));
 sg13g2_buf_2 fanout423 (.A(net424),
    .X(net423));
 sg13g2_buf_2 fanout424 (.A(_0810_),
    .X(net424));
 sg13g2_buf_2 fanout425 (.A(net426),
    .X(net425));
 sg13g2_buf_2 fanout426 (.A(_0781_),
    .X(net426));
 sg13g2_buf_2 fanout427 (.A(net428),
    .X(net427));
 sg13g2_buf_4 fanout428 (.X(net428),
    .A(_0937_));
 sg13g2_buf_2 fanout429 (.A(_0671_),
    .X(net429));
 sg13g2_buf_4 fanout430 (.X(net430),
    .A(_0670_));
 sg13g2_buf_2 fanout431 (.A(_1155_),
    .X(net431));
 sg13g2_buf_2 fanout432 (.A(_1155_),
    .X(net432));
 sg13g2_buf_2 fanout433 (.A(_0773_),
    .X(net433));
 sg13g2_buf_2 fanout434 (.A(_0773_),
    .X(net434));
 sg13g2_buf_4 fanout435 (.X(net435),
    .A(_0616_));
 sg13g2_buf_2 fanout436 (.A(_0415_),
    .X(net436));
 sg13g2_buf_2 fanout437 (.A(_0415_),
    .X(net437));
 sg13g2_buf_4 fanout438 (.X(net438),
    .A(_0414_));
 sg13g2_buf_2 fanout439 (.A(_0414_),
    .X(net439));
 sg13g2_buf_4 fanout440 (.X(net440),
    .A(_0378_));
 sg13g2_buf_4 fanout441 (.X(net441),
    .A(net442));
 sg13g2_buf_2 fanout442 (.A(_1203_),
    .X(net442));
 sg13g2_buf_4 fanout443 (.X(net443),
    .A(_1202_));
 sg13g2_buf_4 fanout444 (.X(net444),
    .A(net312));
 sg13g2_buf_4 fanout445 (.X(net445),
    .A(net542));
 sg13g2_buf_4 fanout446 (.X(net446),
    .A(net448));
 sg13g2_buf_1 fanout447 (.A(net448),
    .X(net447));
 sg13g2_buf_4 fanout448 (.X(net448),
    .A(\uart_proj.fifoRx.read_ptr[2] ));
 sg13g2_buf_4 fanout449 (.X(net449),
    .A(net453));
 sg13g2_buf_2 fanout450 (.A(net453),
    .X(net450));
 sg13g2_buf_2 fanout451 (.A(net452),
    .X(net451));
 sg13g2_buf_2 fanout452 (.A(net453),
    .X(net452));
 sg13g2_buf_2 fanout453 (.A(\uart_proj.fifoRx.read_ptr[1] ),
    .X(net453));
 sg13g2_buf_4 fanout454 (.X(net454),
    .A(net457));
 sg13g2_buf_1 fanout455 (.A(net457),
    .X(net455));
 sg13g2_buf_4 fanout456 (.X(net456),
    .A(net457));
 sg13g2_buf_2 fanout457 (.A(\uart_proj.fifoRx.read_ptr[0] ),
    .X(net457));
 sg13g2_buf_2 fanout458 (.A(net462),
    .X(net458));
 sg13g2_buf_2 fanout459 (.A(net462),
    .X(net459));
 sg13g2_buf_2 fanout460 (.A(net462),
    .X(net460));
 sg13g2_buf_1 fanout461 (.A(net462),
    .X(net461));
 sg13g2_buf_2 fanout462 (.A(\uart_proj.fifoRx.read_ptr[0] ),
    .X(net462));
 sg13g2_buf_2 fanout463 (.A(\uart_proj.fifoTx.read_ptr[2] ),
    .X(net463));
 sg13g2_buf_2 fanout464 (.A(net466),
    .X(net464));
 sg13g2_buf_4 fanout465 (.X(net465),
    .A(\uart_proj.fifoTx.read_ptr[1] ));
 sg13g2_buf_1 fanout466 (.A(\uart_proj.fifoTx.read_ptr[1] ),
    .X(net466));
 sg13g2_buf_4 fanout467 (.X(net467),
    .A(net472));
 sg13g2_buf_4 fanout468 (.X(net468),
    .A(net472));
 sg13g2_buf_2 fanout469 (.A(net470),
    .X(net469));
 sg13g2_buf_2 fanout470 (.A(net472),
    .X(net470));
 sg13g2_buf_2 fanout471 (.A(net472),
    .X(net471));
 sg13g2_buf_2 fanout472 (.A(\uart_proj.fifoTx.read_ptr[0] ),
    .X(net472));
 sg13g2_buf_4 fanout473 (.X(net473),
    .A(net529));
 sg13g2_buf_4 fanout474 (.X(net474),
    .A(\uart_proj.bg.rate[11] ));
 sg13g2_buf_2 fanout475 (.A(\uart_proj.bg.rate[11] ),
    .X(net475));
 sg13g2_buf_2 fanout476 (.A(net477),
    .X(net476));
 sg13g2_buf_1 fanout477 (.A(net478),
    .X(net477));
 sg13g2_buf_4 fanout478 (.X(net478),
    .A(\uart_proj.bg.rate[0] ));
 sg13g2_buf_2 fanout479 (.A(\uart_proj.bg.rate[5] ),
    .X(net479));
 sg13g2_buf_4 fanout480 (.X(net480),
    .A(net481));
 sg13g2_buf_2 fanout481 (.A(\uart_proj.bg.rate[1] ),
    .X(net481));
 sg13g2_buf_4 fanout482 (.X(net482),
    .A(net486));
 sg13g2_buf_4 fanout483 (.X(net483),
    .A(net486));
 sg13g2_buf_4 fanout484 (.X(net484),
    .A(net486));
 sg13g2_buf_4 fanout485 (.X(net485),
    .A(net486));
 sg13g2_buf_2 fanout486 (.A(net487),
    .X(net486));
 sg13g2_buf_4 fanout487 (.X(net487),
    .A(net528));
 sg13g2_buf_4 fanout488 (.X(net488),
    .A(net490));
 sg13g2_buf_4 fanout489 (.X(net489),
    .A(net490));
 sg13g2_buf_4 fanout490 (.X(net490),
    .A(net492));
 sg13g2_buf_4 fanout491 (.X(net491),
    .A(net492));
 sg13g2_buf_2 fanout492 (.A(net528),
    .X(net492));
 sg13g2_buf_4 fanout493 (.X(net493),
    .A(net496));
 sg13g2_buf_2 fanout494 (.A(net496),
    .X(net494));
 sg13g2_buf_4 fanout495 (.X(net495),
    .A(net496));
 sg13g2_buf_2 fanout496 (.A(net528),
    .X(net496));
 sg13g2_buf_4 fanout497 (.X(net497),
    .A(net501));
 sg13g2_buf_2 fanout498 (.A(net501),
    .X(net498));
 sg13g2_buf_4 fanout499 (.X(net499),
    .A(net501));
 sg13g2_buf_2 fanout500 (.A(net501),
    .X(net500));
 sg13g2_buf_1 fanout501 (.A(net527),
    .X(net501));
 sg13g2_buf_4 fanout502 (.X(net502),
    .A(net504));
 sg13g2_buf_4 fanout503 (.X(net503),
    .A(net504));
 sg13g2_buf_2 fanout504 (.A(net527),
    .X(net504));
 sg13g2_buf_4 fanout505 (.X(net505),
    .A(net508));
 sg13g2_buf_4 fanout506 (.X(net506),
    .A(net508));
 sg13g2_buf_2 fanout507 (.A(net508),
    .X(net507));
 sg13g2_buf_2 fanout508 (.A(net511),
    .X(net508));
 sg13g2_buf_4 fanout509 (.X(net509),
    .A(net510));
 sg13g2_buf_4 fanout510 (.X(net510),
    .A(net511));
 sg13g2_buf_2 fanout511 (.A(net527),
    .X(net511));
 sg13g2_buf_4 fanout512 (.X(net512),
    .A(net514));
 sg13g2_buf_4 fanout513 (.X(net513),
    .A(net514));
 sg13g2_buf_4 fanout514 (.X(net514),
    .A(net526));
 sg13g2_buf_4 fanout515 (.X(net515),
    .A(net516));
 sg13g2_buf_4 fanout516 (.X(net516),
    .A(net518));
 sg13g2_buf_4 fanout517 (.X(net517),
    .A(net518));
 sg13g2_buf_4 fanout518 (.X(net518),
    .A(net526));
 sg13g2_buf_4 fanout519 (.X(net519),
    .A(net526));
 sg13g2_buf_4 fanout520 (.X(net520),
    .A(net526));
 sg13g2_buf_4 fanout521 (.X(net521),
    .A(net525));
 sg13g2_buf_2 fanout522 (.A(net525),
    .X(net522));
 sg13g2_buf_4 fanout523 (.X(net523),
    .A(net525));
 sg13g2_buf_4 fanout524 (.X(net524),
    .A(net525));
 sg13g2_buf_2 fanout525 (.A(net526),
    .X(net525));
 sg13g2_buf_2 fanout526 (.A(net527),
    .X(net526));
 sg13g2_buf_2 fanout527 (.A(net528),
    .X(net527));
 sg13g2_buf_2 fanout528 (.A(rst_n),
    .X(net528));
 sg13g2_buf_4 input1 (.X(net1),
    .A(ui_in[0]));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_4 input3 (.X(net3),
    .A(ui_in[2]));
 sg13g2_buf_4 input4 (.X(net4),
    .A(ui_in[3]));
 sg13g2_buf_1 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[5]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(uio_in[0]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(uio_in[1]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(uio_in[2]),
    .X(net9));
 sg13g2_buf_1 input10 (.A(uio_in[3]),
    .X(net10));
 sg13g2_buf_1 input11 (.A(uio_in[4]),
    .X(net11));
 sg13g2_buf_1 input12 (.A(uio_in[5]),
    .X(net12));
 sg13g2_buf_1 input13 (.A(uio_in[6]),
    .X(net13));
 sg13g2_buf_1 input14 (.A(uio_in[7]),
    .X(net14));
 sg13g2_tielo tt_um_purdue_socet_uart_15 (.L_LO(net15));
 sg13g2_buf_2 clkbuf_leaf_1_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_2 clkbuf_leaf_2_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_2 clkbuf_leaf_3_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_2 clkbuf_leaf_4_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_2 clkbuf_leaf_5_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_2 clkbuf_leaf_6_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_2 clkbuf_leaf_7_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_2 clkbuf_leaf_8_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_2 clkbuf_leaf_9_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_2 clkbuf_leaf_10_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_2 clkbuf_leaf_11_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_2 clkbuf_leaf_12_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_2 clkbuf_leaf_13_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_2 clkbuf_leaf_14_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_2 clkbuf_leaf_15_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_2 clkbuf_leaf_16_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_2 clkbuf_leaf_17_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_2 clkbuf_leaf_18_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_2 clkbuf_leaf_19_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_2 clkbuf_leaf_20_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_2 clkbuf_leaf_21_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_2 clkbuf_leaf_22_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_2 clkbuf_leaf_23_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_2 clkbuf_leaf_24_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_2 clkbuf_leaf_25_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_2 clkbuf_leaf_26_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_2 clkbuf_leaf_27_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_2 clkbuf_leaf_28_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_2 clkbuf_leaf_29_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_2 clkbuf_leaf_30_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_2 clkbuf_leaf_31_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_31_clk));
 sg13g2_buf_2 clkbuf_leaf_32_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_32_clk));
 sg13g2_buf_2 clkbuf_leaf_34_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_34_clk));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_2 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sg13g2_buf_2 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sg13g2_buf_2 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sg13g2_buf_2 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sg13g2_buf_2 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sg13g2_buf_2 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sg13g2_buf_2 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sg13g2_buf_2 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_3_1__leaf_clk));
 sg13g2_buf_1 clkload1 (.A(clknet_3_2__leaf_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_3_3__leaf_clk));
 sg13g2_buf_1 clkload3 (.A(clknet_3_4__leaf_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_3_5__leaf_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_3_6__leaf_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_3_7__leaf_clk));
 sg13g2_inv_1 clkload7 (.A(clknet_leaf_34_clk));
 sg13g2_inv_8 clkload8 (.A(clknet_leaf_26_clk));
 sg13g2_inv_1 clkload9 (.A(clknet_leaf_31_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\uart_proj.uartTx.curState[0] ),
    .X(net18));
 sg13g2_dlygate4sd3_1 hold2 (.A(_0158_),
    .X(net19));
 sg13g2_dlygate4sd3_1 hold3 (.A(_0035_),
    .X(net20));
 sg13g2_dlygate4sd3_1 hold4 (.A(\uart_proj.uartRx.readCount[0] ),
    .X(net21));
 sg13g2_dlygate4sd3_1 hold5 (.A(_0882_),
    .X(net22));
 sg13g2_dlygate4sd3_1 hold6 (.A(_0348_),
    .X(net23));
 sg13g2_dlygate4sd3_1 hold7 (.A(\uart_proj.rxData[3] ),
    .X(net24));
 sg13g2_dlygate4sd3_1 hold8 (.A(_0008_),
    .X(net25));
 sg13g2_dlygate4sd3_1 hold9 (.A(\uart_proj.rxData[4] ),
    .X(net26));
 sg13g2_dlygate4sd3_1 hold10 (.A(_0009_),
    .X(net27));
 sg13g2_dlygate4sd3_1 hold11 (.A(\uart_proj.rxData[5] ),
    .X(net28));
 sg13g2_dlygate4sd3_1 hold12 (.A(_0010_),
    .X(net29));
 sg13g2_dlygate4sd3_1 hold13 (.A(\uart_proj.rxData[6] ),
    .X(net30));
 sg13g2_dlygate4sd3_1 hold14 (.A(_0011_),
    .X(net31));
 sg13g2_dlygate4sd3_1 hold15 (.A(\uart_proj.rxData[7] ),
    .X(net32));
 sg13g2_dlygate4sd3_1 hold16 (.A(_0012_),
    .X(net33));
 sg13g2_dlygate4sd3_1 hold17 (.A(\uart_proj.rxData[0] ),
    .X(net34));
 sg13g2_dlygate4sd3_1 hold18 (.A(_0005_),
    .X(net35));
 sg13g2_dlygate4sd3_1 hold19 (.A(_0040_),
    .X(net36));
 sg13g2_dlygate4sd3_1 hold20 (.A(_0638_),
    .X(net37));
 sg13g2_dlygate4sd3_1 hold21 (.A(_0238_),
    .X(net38));
 sg13g2_dlygate4sd3_1 hold22 (.A(\uart_proj.rxData[2] ),
    .X(net39));
 sg13g2_dlygate4sd3_1 hold23 (.A(_0007_),
    .X(net40));
 sg13g2_dlygate4sd3_1 hold24 (.A(_0030_),
    .X(net41));
 sg13g2_dlygate4sd3_1 hold25 (.A(_0001_),
    .X(net42));
 sg13g2_dlygate4sd3_1 hold26 (.A(\uart_proj.fifoTx.fifo[42] ),
    .X(net43));
 sg13g2_dlygate4sd3_1 hold27 (.A(_0153_),
    .X(net44));
 sg13g2_dlygate4sd3_1 hold28 (.A(_0350_),
    .X(net45));
 sg13g2_dlygate4sd3_1 hold29 (.A(\uart_proj.fifoTx.fifo[63] ),
    .X(net46));
 sg13g2_dlygate4sd3_1 hold30 (.A(\uart_proj.fifoTx.fifo[56] ),
    .X(net47));
 sg13g2_dlygate4sd3_1 hold31 (.A(_0865_),
    .X(net48));
 sg13g2_dlygate4sd3_1 hold32 (.A(_0328_),
    .X(net49));
 sg13g2_dlygate4sd3_1 hold33 (.A(\uart_proj.fifoTx.fifo[51] ),
    .X(net50));
 sg13g2_dlygate4sd3_1 hold34 (.A(\uart_proj.fifoTx.fifo[29] ),
    .X(net51));
 sg13g2_dlygate4sd3_1 hold35 (.A(\uart_proj.fifoTx.fifo[25] ),
    .X(net52));
 sg13g2_dlygate4sd3_1 hold36 (.A(_0297_),
    .X(net53));
 sg13g2_dlygate4sd3_1 hold37 (.A(\uart_proj.fifoTx.fifo[12] ),
    .X(net54));
 sg13g2_dlygate4sd3_1 hold38 (.A(\uart_proj.fifoTx.fifo[52] ),
    .X(net55));
 sg13g2_dlygate4sd3_1 hold39 (.A(\uart_proj.fifoTx.fifo[58] ),
    .X(net56));
 sg13g2_dlygate4sd3_1 hold40 (.A(\uart_proj.fifoTx.fifo[11] ),
    .X(net57));
 sg13g2_dlygate4sd3_1 hold41 (.A(\uart_proj.fifoTx.fifo[55] ),
    .X(net58));
 sg13g2_dlygate4sd3_1 hold42 (.A(\uart_proj.fifoTx.fifo[48] ),
    .X(net59));
 sg13g2_dlygate4sd3_1 hold43 (.A(\uart_proj.fifoTx.fifo[45] ),
    .X(net60));
 sg13g2_dlygate4sd3_1 hold44 (.A(\uart_proj.fifoTx.fifo[14] ),
    .X(net61));
 sg13g2_dlygate4sd3_1 hold45 (.A(\uart_proj.fifoTx.fifo[13] ),
    .X(net62));
 sg13g2_dlygate4sd3_1 hold46 (.A(\uart_proj.fifoTx.fifo[54] ),
    .X(net63));
 sg13g2_dlygate4sd3_1 hold47 (.A(\uart_proj.fifoTx.fifo[46] ),
    .X(net64));
 sg13g2_dlygate4sd3_1 hold48 (.A(_0157_),
    .X(net65));
 sg13g2_dlygate4sd3_1 hold49 (.A(_0354_),
    .X(net66));
 sg13g2_dlygate4sd3_1 hold50 (.A(\uart_proj.fifoTx.fifo[61] ),
    .X(net67));
 sg13g2_dlygate4sd3_1 hold51 (.A(\uart_proj.rxData[1] ),
    .X(net68));
 sg13g2_dlygate4sd3_1 hold52 (.A(_0006_),
    .X(net69));
 sg13g2_dlygate4sd3_1 hold53 (.A(\uart_proj.fifoTx.fifo[8] ),
    .X(net70));
 sg13g2_dlygate4sd3_1 hold54 (.A(_0280_),
    .X(net71));
 sg13g2_dlygate4sd3_1 hold55 (.A(\uart_proj.fifoTx.fifo[10] ),
    .X(net72));
 sg13g2_dlygate4sd3_1 hold56 (.A(\uart_proj.fifoTx.fifo[30] ),
    .X(net73));
 sg13g2_dlygate4sd3_1 hold57 (.A(\uart_proj.fifoTx.fifo[26] ),
    .X(net74));
 sg13g2_dlygate4sd3_1 hold58 (.A(\uart_proj.fifoTx.fifo[50] ),
    .X(net75));
 sg13g2_dlygate4sd3_1 hold59 (.A(\uart_proj.fifoTx.fifo[27] ),
    .X(net76));
 sg13g2_dlygate4sd3_1 hold60 (.A(\uart_proj.fifoTx.fifo[44] ),
    .X(net77));
 sg13g2_dlygate4sd3_1 hold61 (.A(\uart_proj.fifoTx.fifo[31] ),
    .X(net78));
 sg13g2_dlygate4sd3_1 hold62 (.A(\uart_proj.fifoTx.fifo[15] ),
    .X(net79));
 sg13g2_dlygate4sd3_1 hold63 (.A(\uart_proj.fifoTx.fifo[59] ),
    .X(net80));
 sg13g2_dlygate4sd3_1 hold64 (.A(\uart_proj.fifoTx.fifo[57] ),
    .X(net81));
 sg13g2_dlygate4sd3_1 hold65 (.A(_0329_),
    .X(net82));
 sg13g2_dlygate4sd3_1 hold66 (.A(\uart_proj.fifoTx.fifo[28] ),
    .X(net83));
 sg13g2_dlygate4sd3_1 hold67 (.A(\uart_proj.fifoTx.fifo[24] ),
    .X(net84));
 sg13g2_dlygate4sd3_1 hold68 (.A(_0296_),
    .X(net85));
 sg13g2_dlygate4sd3_1 hold69 (.A(\uart_proj.fifoTx.fifo[41] ),
    .X(net86));
 sg13g2_dlygate4sd3_1 hold70 (.A(_0313_),
    .X(net87));
 sg13g2_dlygate4sd3_1 hold71 (.A(\uart_proj.err ),
    .X(net88));
 sg13g2_dlygate4sd3_1 hold72 (.A(_0155_),
    .X(net89));
 sg13g2_dlygate4sd3_1 hold73 (.A(_0352_),
    .X(net90));
 sg13g2_dlygate4sd3_1 hold74 (.A(\uart_proj.fifoTx.fifo[9] ),
    .X(net91));
 sg13g2_dlygate4sd3_1 hold75 (.A(_0281_),
    .X(net92));
 sg13g2_dlygate4sd3_1 hold76 (.A(\uart_proj.fifoTx.fifo[62] ),
    .X(net93));
 sg13g2_dlygate4sd3_1 hold77 (.A(\uart_proj.bg.rxCount[15] ),
    .X(net94));
 sg13g2_dlygate4sd3_1 hold78 (.A(_0259_),
    .X(net95));
 sg13g2_dlygate4sd3_1 hold79 (.A(\uart_proj.uartTx.writeBuf[6] ),
    .X(net96));
 sg13g2_dlygate4sd3_1 hold80 (.A(_0266_),
    .X(net97));
 sg13g2_dlygate4sd3_1 hold81 (.A(\uart_proj.fifoTx.fifo[53] ),
    .X(net98));
 sg13g2_dlygate4sd3_1 hold82 (.A(\uart_proj.fifoTx.fifo[60] ),
    .X(net99));
 sg13g2_dlygate4sd3_1 hold83 (.A(_0156_),
    .X(net100));
 sg13g2_dlygate4sd3_1 hold84 (.A(_0353_),
    .X(net101));
 sg13g2_dlygate4sd3_1 hold85 (.A(\uart_proj.fifoRx.fifo[14] ),
    .X(net102));
 sg13g2_dlygate4sd3_1 hold86 (.A(_0181_),
    .X(net103));
 sg13g2_dlygate4sd3_1 hold87 (.A(\uart_proj.fifoRx.fifo[44] ),
    .X(net104));
 sg13g2_dlygate4sd3_1 hold88 (.A(_0211_),
    .X(net105));
 sg13g2_dlygate4sd3_1 hold89 (.A(\uart_proj.fifoTx.fifo[21] ),
    .X(net106));
 sg13g2_dlygate4sd3_1 hold90 (.A(\uart_proj.fifoRx.fifo[9] ),
    .X(net107));
 sg13g2_dlygate4sd3_1 hold91 (.A(_0176_),
    .X(net108));
 sg13g2_dlygate4sd3_1 hold92 (.A(\uart_proj.fifoTx.fifo[47] ),
    .X(net109));
 sg13g2_dlygate4sd3_1 hold93 (.A(\uart_proj.fifoRx.fifo[10] ),
    .X(net110));
 sg13g2_dlygate4sd3_1 hold94 (.A(_0177_),
    .X(net111));
 sg13g2_dlygate4sd3_1 hold95 (.A(\uart_proj.fifoTx.fifo[19] ),
    .X(net112));
 sg13g2_dlygate4sd3_1 hold96 (.A(\uart_proj.fifoTx.fifo[43] ),
    .X(net113));
 sg13g2_dlygate4sd3_1 hold97 (.A(\uart_proj.fifoTx.fifo[17] ),
    .X(net114));
 sg13g2_dlygate4sd3_1 hold98 (.A(\uart_proj.fifoTx.fifo[49] ),
    .X(net115));
 sg13g2_dlygate4sd3_1 hold99 (.A(\uart_proj.fifoRx.fifo[41] ),
    .X(net116));
 sg13g2_dlygate4sd3_1 hold100 (.A(_0208_),
    .X(net117));
 sg13g2_dlygate4sd3_1 hold101 (.A(_0146_),
    .X(net118));
 sg13g2_dlygate4sd3_1 hold102 (.A(_0166_),
    .X(net119));
 sg13g2_dlygate4sd3_1 hold103 (.A(\uart_proj.txData[7] ),
    .X(net120));
 sg13g2_dlygate4sd3_1 hold104 (.A(_0760_),
    .X(net121));
 sg13g2_dlygate4sd3_1 hold105 (.A(_0154_),
    .X(net122));
 sg13g2_dlygate4sd3_1 hold106 (.A(_0351_),
    .X(net123));
 sg13g2_dlygate4sd3_1 hold107 (.A(_0152_),
    .X(net124));
 sg13g2_dlygate4sd3_1 hold108 (.A(\uart_proj.fifoRx.fifo[43] ),
    .X(net125));
 sg13g2_dlygate4sd3_1 hold109 (.A(_0210_),
    .X(net126));
 sg13g2_dlygate4sd3_1 hold110 (.A(\uart_proj.fifoRx.fifo[12] ),
    .X(net127));
 sg13g2_dlygate4sd3_1 hold111 (.A(_0179_),
    .X(net128));
 sg13g2_dlygate4sd3_1 hold112 (.A(\uart_proj.fifoTx.fifo[16] ),
    .X(net129));
 sg13g2_dlygate4sd3_1 hold113 (.A(\uart_proj.uartTx.writeBuf[1] ),
    .X(net130));
 sg13g2_dlygate4sd3_1 hold114 (.A(_0261_),
    .X(net131));
 sg13g2_dlygate4sd3_1 hold115 (.A(\uart_proj.fifoTx.fifo[40] ),
    .X(net132));
 sg13g2_dlygate4sd3_1 hold116 (.A(_0312_),
    .X(net133));
 sg13g2_dlygate4sd3_1 hold117 (.A(\uart_proj.fifoTx.fifo[22] ),
    .X(net134));
 sg13g2_dlygate4sd3_1 hold118 (.A(\uart_proj.fifoRx.overrun ),
    .X(net135));
 sg13g2_dlygate4sd3_1 hold119 (.A(_0004_),
    .X(net136));
 sg13g2_dlygate4sd3_1 hold120 (.A(\uart_proj.fifoRx.fifo[13] ),
    .X(net137));
 sg13g2_dlygate4sd3_1 hold121 (.A(_0180_),
    .X(net138));
 sg13g2_dlygate4sd3_1 hold122 (.A(\uart_proj.fifoRx.fifo[23] ),
    .X(net139));
 sg13g2_dlygate4sd3_1 hold123 (.A(_0190_),
    .X(net140));
 sg13g2_dlygate4sd3_1 hold124 (.A(\uart_proj.fifoTx.fifo[18] ),
    .X(net141));
 sg13g2_dlygate4sd3_1 hold125 (.A(\uart_proj.fifoTx.fifo[23] ),
    .X(net142));
 sg13g2_dlygate4sd3_1 hold126 (.A(\uart_proj.bg.rxCount[11] ),
    .X(net143));
 sg13g2_dlygate4sd3_1 hold127 (.A(_0255_),
    .X(net144));
 sg13g2_dlygate4sd3_1 hold128 (.A(\uart_proj.fifoRx.fifo[42] ),
    .X(net145));
 sg13g2_dlygate4sd3_1 hold129 (.A(_0209_),
    .X(net146));
 sg13g2_dlygate4sd3_1 hold130 (.A(\uart_proj.fifoRx.fifo[47] ),
    .X(net147));
 sg13g2_dlygate4sd3_1 hold131 (.A(_0214_),
    .X(net148));
 sg13g2_dlygate4sd3_1 hold132 (.A(\uart_proj.fifoRx.fifo[15] ),
    .X(net149));
 sg13g2_dlygate4sd3_1 hold133 (.A(_0182_),
    .X(net150));
 sg13g2_dlygate4sd3_1 hold134 (.A(\uart_proj.fifoRx.fifo[20] ),
    .X(net151));
 sg13g2_dlygate4sd3_1 hold135 (.A(_0187_),
    .X(net152));
 sg13g2_dlygate4sd3_1 hold136 (.A(\uart_proj.fifoRx.fifo[39] ),
    .X(net153));
 sg13g2_dlygate4sd3_1 hold137 (.A(_0651_),
    .X(net154));
 sg13g2_dlygate4sd3_1 hold138 (.A(\uart_proj.uartTx.writeBuf[2] ),
    .X(net155));
 sg13g2_dlygate4sd3_1 hold139 (.A(_0262_),
    .X(net156));
 sg13g2_dlygate4sd3_1 hold140 (.A(\uart_proj.fifoTx.fifo[33] ),
    .X(net157));
 sg13g2_dlygate4sd3_1 hold141 (.A(\uart_proj.fifoRx.fifo[11] ),
    .X(net158));
 sg13g2_dlygate4sd3_1 hold142 (.A(_0178_),
    .X(net159));
 sg13g2_dlygate4sd3_1 hold143 (.A(\uart_proj.fifoTx.fifo[34] ),
    .X(net160));
 sg13g2_dlygate4sd3_1 hold144 (.A(\uart_proj.fifoTx.fifo[36] ),
    .X(net161));
 sg13g2_dlygate4sd3_1 hold145 (.A(\uart_proj.fifoTx.fifo[35] ),
    .X(net162));
 sg13g2_dlygate4sd3_1 hold146 (.A(\uart_proj.fifoRx.fifo[45] ),
    .X(net163));
 sg13g2_dlygate4sd3_1 hold147 (.A(_0212_),
    .X(net164));
 sg13g2_dlygate4sd3_1 hold148 (.A(\uart_proj.fifoTx.fifo[38] ),
    .X(net165));
 sg13g2_dlygate4sd3_1 hold149 (.A(\uart_proj.fifoTx.fifo[32] ),
    .X(net166));
 sg13g2_dlygate4sd3_1 hold150 (.A(\uart_proj.fifoRx.fifo[17] ),
    .X(net167));
 sg13g2_dlygate4sd3_1 hold151 (.A(_0184_),
    .X(net168));
 sg13g2_dlygate4sd3_1 hold152 (.A(\uart_proj.fifoRx.fifo[21] ),
    .X(net169));
 sg13g2_dlygate4sd3_1 hold153 (.A(_0188_),
    .X(net170));
 sg13g2_dlygate4sd3_1 hold154 (.A(\uart_proj.fifoTx.fifo[20] ),
    .X(net171));
 sg13g2_dlygate4sd3_1 hold155 (.A(\uart_proj.fifoRx.fifo[35] ),
    .X(net172));
 sg13g2_dlygate4sd3_1 hold156 (.A(_0647_),
    .X(net173));
 sg13g2_dlygate4sd3_1 hold157 (.A(\uart_proj.fifoRx.fifo[18] ),
    .X(net174));
 sg13g2_dlygate4sd3_1 hold158 (.A(_0185_),
    .X(net175));
 sg13g2_dlygate4sd3_1 hold159 (.A(\uart_proj.fifoRx.fifo[40] ),
    .X(net176));
 sg13g2_dlygate4sd3_1 hold160 (.A(_0207_),
    .X(net177));
 sg13g2_dlygate4sd3_1 hold161 (.A(\uart_proj.fifoRx.fifo[46] ),
    .X(net178));
 sg13g2_dlygate4sd3_1 hold162 (.A(_0213_),
    .X(net179));
 sg13g2_dlygate4sd3_1 hold163 (.A(\uart_proj.fifoRx.fifo[33] ),
    .X(net180));
 sg13g2_dlygate4sd3_1 hold164 (.A(_0645_),
    .X(net181));
 sg13g2_dlygate4sd3_1 hold165 (.A(\uart_proj.uartTx.writeBuf[5] ),
    .X(net182));
 sg13g2_dlygate4sd3_1 hold166 (.A(_0265_),
    .X(net183));
 sg13g2_dlygate4sd3_1 hold167 (.A(\uart_proj.fifoRx.fifo[62] ),
    .X(net184));
 sg13g2_dlygate4sd3_1 hold168 (.A(_0229_),
    .X(net185));
 sg13g2_dlygate4sd3_1 hold169 (.A(\uart_proj.uartTx.writeBuf[4] ),
    .X(net186));
 sg13g2_dlygate4sd3_1 hold170 (.A(_0264_),
    .X(net187));
 sg13g2_dlygate4sd3_1 hold171 (.A(\uart_proj.fifoTx.fifo[39] ),
    .X(net188));
 sg13g2_dlygate4sd3_1 hold172 (.A(\uart_proj.fifoRx.fifo[24] ),
    .X(net189));
 sg13g2_dlygate4sd3_1 hold173 (.A(_0191_),
    .X(net190));
 sg13g2_dlygate4sd3_1 hold174 (.A(\uart_proj.uartRx.readBuf[0] ),
    .X(net191));
 sg13g2_dlygate4sd3_1 hold175 (.A(\uart_proj.fifoRx.fifo[8] ),
    .X(net192));
 sg13g2_dlygate4sd3_1 hold176 (.A(_0175_),
    .X(net193));
 sg13g2_dlygate4sd3_1 hold177 (.A(\uart_proj.fifoTx.fifo[37] ),
    .X(net194));
 sg13g2_dlygate4sd3_1 hold178 (.A(\uart_proj.fifoTx.fifo[0] ),
    .X(net195));
 sg13g2_dlygate4sd3_1 hold179 (.A(\uart_proj.fifoRx.fifo[37] ),
    .X(net196));
 sg13g2_dlygate4sd3_1 hold180 (.A(_0649_),
    .X(net197));
 sg13g2_dlygate4sd3_1 hold181 (.A(\uart_proj.fifoRx.fifo[57] ),
    .X(net198));
 sg13g2_dlygate4sd3_1 hold182 (.A(_0224_),
    .X(net199));
 sg13g2_dlygate4sd3_1 hold183 (.A(\uart_proj.fifoRx.fifo[49] ),
    .X(net200));
 sg13g2_dlygate4sd3_1 hold184 (.A(_0216_),
    .X(net201));
 sg13g2_dlygate4sd3_1 hold185 (.A(\uart_proj.fifoRx.fifo[28] ),
    .X(net202));
 sg13g2_dlygate4sd3_1 hold186 (.A(_0195_),
    .X(net203));
 sg13g2_dlygate4sd3_1 hold187 (.A(\uart_proj.fifoRx.fifo[25] ),
    .X(net204));
 sg13g2_dlygate4sd3_1 hold188 (.A(_0192_),
    .X(net205));
 sg13g2_dlygate4sd3_1 hold189 (.A(\uart_proj.fifoRx.fifo[36] ),
    .X(net206));
 sg13g2_dlygate4sd3_1 hold190 (.A(_0648_),
    .X(net207));
 sg13g2_dlygate4sd3_1 hold191 (.A(\uart_proj.fifoRx.fifo[34] ),
    .X(net208));
 sg13g2_dlygate4sd3_1 hold192 (.A(_0646_),
    .X(net209));
 sg13g2_dlygate4sd3_1 hold193 (.A(\uart_proj.fifoRx.fifo[63] ),
    .X(net210));
 sg13g2_dlygate4sd3_1 hold194 (.A(_0230_),
    .X(net211));
 sg13g2_dlygate4sd3_1 hold195 (.A(\uart_proj.fifoRx.fifo[56] ),
    .X(net212));
 sg13g2_dlygate4sd3_1 hold196 (.A(_0223_),
    .X(net213));
 sg13g2_dlygate4sd3_1 hold197 (.A(\uart_proj.uartRx.readBuf[4] ),
    .X(net214));
 sg13g2_dlygate4sd3_1 hold198 (.A(\uart_proj.uartRx.edgeCmp ),
    .X(net215));
 sg13g2_dlygate4sd3_1 hold199 (.A(_0271_),
    .X(net216));
 sg13g2_dlygate4sd3_1 hold200 (.A(\uart_proj.uartRx.readBuf[2] ),
    .X(net217));
 sg13g2_dlygate4sd3_1 hold201 (.A(\uart_proj.fifoRx.fifo[22] ),
    .X(net218));
 sg13g2_dlygate4sd3_1 hold202 (.A(_0189_),
    .X(net219));
 sg13g2_dlygate4sd3_1 hold203 (.A(\uart_proj.fifoRx.fifo[31] ),
    .X(net220));
 sg13g2_dlygate4sd3_1 hold204 (.A(_0198_),
    .X(net221));
 sg13g2_dlygate4sd3_1 hold205 (.A(\uart_proj.uartRx.readBuf[7] ),
    .X(net222));
 sg13g2_dlygate4sd3_1 hold206 (.A(\uart_proj.fifoRx.fifo[29] ),
    .X(net223));
 sg13g2_dlygate4sd3_1 hold207 (.A(_0196_),
    .X(net224));
 sg13g2_dlygate4sd3_1 hold208 (.A(\uart_proj.fifoRx.fifo[48] ),
    .X(net225));
 sg13g2_dlygate4sd3_1 hold209 (.A(_0215_),
    .X(net226));
 sg13g2_dlygate4sd3_1 hold210 (.A(\uart_proj.uartRx.readBuf[6] ),
    .X(net227));
 sg13g2_dlygate4sd3_1 hold211 (.A(\uart_proj.fifoRx.fifo[51] ),
    .X(net228));
 sg13g2_dlygate4sd3_1 hold212 (.A(_0218_),
    .X(net229));
 sg13g2_dlygate4sd3_1 hold213 (.A(_0032_),
    .X(net230));
 sg13g2_dlygate4sd3_1 hold214 (.A(_0682_),
    .X(net231));
 sg13g2_dlygate4sd3_1 hold215 (.A(\uart_proj.uartTx.writeBuf[0] ),
    .X(net232));
 sg13g2_dlygate4sd3_1 hold216 (.A(_0260_),
    .X(net233));
 sg13g2_dlygate4sd3_1 hold217 (.A(\uart_proj.uartTx.writeBuf[3] ),
    .X(net234));
 sg13g2_dlygate4sd3_1 hold218 (.A(_0263_),
    .X(net235));
 sg13g2_dlygate4sd3_1 hold219 (.A(\uart_proj.uartTx.hasData ),
    .X(net236));
 sg13g2_dlygate4sd3_1 hold220 (.A(_0269_),
    .X(net237));
 sg13g2_dlygate4sd3_1 hold221 (.A(\uart_proj.fifoTx.fifo[2] ),
    .X(net238));
 sg13g2_dlygate4sd3_1 hold222 (.A(\uart_proj.fifoRx.fifo[53] ),
    .X(net239));
 sg13g2_dlygate4sd3_1 hold223 (.A(_0220_),
    .X(net240));
 sg13g2_dlygate4sd3_1 hold224 (.A(\uart_proj.uartRx.readCount[2] ),
    .X(net241));
 sg13g2_dlygate4sd3_1 hold225 (.A(_0349_),
    .X(net242));
 sg13g2_dlygate4sd3_1 hold226 (.A(\uart_proj.fifoRx.fifo[30] ),
    .X(net243));
 sg13g2_dlygate4sd3_1 hold227 (.A(_0197_),
    .X(net244));
 sg13g2_dlygate4sd3_1 hold228 (.A(\uart_proj.fifoTx.fifo[3] ),
    .X(net245));
 sg13g2_dlygate4sd3_1 hold229 (.A(\uart_proj.fifoTx.fifo[4] ),
    .X(net246));
 sg13g2_dlygate4sd3_1 hold230 (.A(\uart_proj.fifoRx.fifo[50] ),
    .X(net247));
 sg13g2_dlygate4sd3_1 hold231 (.A(_0217_),
    .X(net248));
 sg13g2_dlygate4sd3_1 hold232 (.A(\uart_proj.fifoTx.fifo[5] ),
    .X(net249));
 sg13g2_dlygate4sd3_1 hold233 (.A(\uart_proj.fifoRx.fifo[61] ),
    .X(net250));
 sg13g2_dlygate4sd3_1 hold234 (.A(_0228_),
    .X(net251));
 sg13g2_dlygate4sd3_1 hold235 (.A(\uart_proj.fifoRx.fifo[38] ),
    .X(net252));
 sg13g2_dlygate4sd3_1 hold236 (.A(_0650_),
    .X(net253));
 sg13g2_dlygate4sd3_1 hold237 (.A(\uart_proj.fifoTx.fifo[6] ),
    .X(net254));
 sg13g2_dlygate4sd3_1 hold238 (.A(\uart_proj.fifoRx.fifo[60] ),
    .X(net255));
 sg13g2_dlygate4sd3_1 hold239 (.A(_0227_),
    .X(net256));
 sg13g2_dlygate4sd3_1 hold240 (.A(\uart_proj.fifoRx.fifo[59] ),
    .X(net257));
 sg13g2_dlygate4sd3_1 hold241 (.A(_0226_),
    .X(net258));
 sg13g2_dlygate4sd3_1 hold242 (.A(\uart_proj.fifoRx.fifo[19] ),
    .X(net259));
 sg13g2_dlygate4sd3_1 hold243 (.A(_0186_),
    .X(net260));
 sg13g2_dlygate4sd3_1 hold244 (.A(\uart_proj.fifoTx.fifo[7] ),
    .X(net261));
 sg13g2_dlygate4sd3_1 hold245 (.A(\uart_proj.bg.rxCount[12] ),
    .X(net262));
 sg13g2_dlygate4sd3_1 hold246 (.A(_0256_),
    .X(net263));
 sg13g2_dlygate4sd3_1 hold247 (.A(\uart_proj.fifoRx.fifo[16] ),
    .X(net264));
 sg13g2_dlygate4sd3_1 hold248 (.A(_0183_),
    .X(net265));
 sg13g2_dlygate4sd3_1 hold249 (.A(\uart_proj.fifoRx.fifo[26] ),
    .X(net266));
 sg13g2_dlygate4sd3_1 hold250 (.A(_0193_),
    .X(net267));
 sg13g2_dlygate4sd3_1 hold251 (.A(\uart_proj.fifoRx.fifo[32] ),
    .X(net268));
 sg13g2_dlygate4sd3_1 hold252 (.A(_0644_),
    .X(net269));
 sg13g2_dlygate4sd3_1 hold253 (.A(\uart_proj.uartRx.readBuf[3] ),
    .X(net270));
 sg13g2_dlygate4sd3_1 hold254 (.A(\uart_proj.uartRx.readBuf[1] ),
    .X(net271));
 sg13g2_dlygate4sd3_1 hold255 (.A(_0340_),
    .X(net272));
 sg13g2_dlygate4sd3_1 hold256 (.A(\uart_proj.fifoRx.fifo[58] ),
    .X(net273));
 sg13g2_dlygate4sd3_1 hold257 (.A(_0225_),
    .X(net274));
 sg13g2_dlygate4sd3_1 hold258 (.A(\uart_proj.uartRx.readBuf[5] ),
    .X(net275));
 sg13g2_dlygate4sd3_1 hold259 (.A(\uart_proj.fifoRx.fifo[55] ),
    .X(net276));
 sg13g2_dlygate4sd3_1 hold260 (.A(_0222_),
    .X(net277));
 sg13g2_dlygate4sd3_1 hold261 (.A(\uart_proj.fifoRx.fifo[54] ),
    .X(net278));
 sg13g2_dlygate4sd3_1 hold262 (.A(_0221_),
    .X(net279));
 sg13g2_dlygate4sd3_1 hold263 (.A(\uart_proj.uartTx.writeCount[1] ),
    .X(net280));
 sg13g2_dlygate4sd3_1 hold264 (.A(_0164_),
    .X(net281));
 sg13g2_dlygate4sd3_1 hold265 (.A(\uart_proj.uartTx.writeCount[2] ),
    .X(net282));
 sg13g2_dlygate4sd3_1 hold266 (.A(_0165_),
    .X(net283));
 sg13g2_dlygate4sd3_1 hold267 (.A(\uart_proj.fifoRx.fifo[27] ),
    .X(net284));
 sg13g2_dlygate4sd3_1 hold268 (.A(_0194_),
    .X(net285));
 sg13g2_dlygate4sd3_1 hold269 (.A(\uart_proj.fifoRx.fifo[3] ),
    .X(net286));
 sg13g2_dlygate4sd3_1 hold270 (.A(_0170_),
    .X(net287));
 sg13g2_dlygate4sd3_1 hold271 (.A(\uart_proj.fifoTx.fifo[1] ),
    .X(net288));
 sg13g2_dlygate4sd3_1 hold272 (.A(\uart_proj.bg.rxCount[4] ),
    .X(net289));
 sg13g2_dlygate4sd3_1 hold273 (.A(\uart_proj.fifoRx.fifo[1] ),
    .X(net290));
 sg13g2_dlygate4sd3_1 hold274 (.A(_0168_),
    .X(net291));
 sg13g2_dlygate4sd3_1 hold275 (.A(\uart_proj.bg.rxCount[7] ),
    .X(net292));
 sg13g2_dlygate4sd3_1 hold276 (.A(\uart_proj.fifoRx.fifo[7] ),
    .X(net293));
 sg13g2_dlygate4sd3_1 hold277 (.A(_0174_),
    .X(net294));
 sg13g2_dlygate4sd3_1 hold278 (.A(\uart_proj.fifoRx.fifo[6] ),
    .X(net295));
 sg13g2_dlygate4sd3_1 hold279 (.A(_0173_),
    .X(net296));
 sg13g2_dlygate4sd3_1 hold280 (.A(\uart_proj.prev_ren_wen[0] ),
    .X(net297));
 sg13g2_dlygate4sd3_1 hold281 (.A(_0409_),
    .X(net298));
 sg13g2_dlygate4sd3_1 hold282 (.A(\uart_proj.fifoRx.fifo[5] ),
    .X(net299));
 sg13g2_dlygate4sd3_1 hold283 (.A(_0172_),
    .X(net300));
 sg13g2_dlygate4sd3_1 hold284 (.A(_0039_),
    .X(net301));
 sg13g2_dlygate4sd3_1 hold285 (.A(_0696_),
    .X(net302));
 sg13g2_dlygate4sd3_1 hold286 (.A(\uart_proj.fifoRx.fifo[0] ),
    .X(net303));
 sg13g2_dlygate4sd3_1 hold287 (.A(_0167_),
    .X(net304));
 sg13g2_dlygate4sd3_1 hold288 (.A(\uart_proj.fifoRx.fifo[4] ),
    .X(net305));
 sg13g2_dlygate4sd3_1 hold289 (.A(_0171_),
    .X(net306));
 sg13g2_dlygate4sd3_1 hold290 (.A(\uart_proj.fifoRx.fifo[2] ),
    .X(net307));
 sg13g2_dlygate4sd3_1 hold291 (.A(_0169_),
    .X(net308));
 sg13g2_dlygate4sd3_1 hold292 (.A(\uart_proj.bg.rxCount[13] ),
    .X(net309));
 sg13g2_dlygate4sd3_1 hold293 (.A(\uart_proj.bg.rxCount[5] ),
    .X(net310));
 sg13g2_dlygate4sd3_1 hold294 (.A(\uart_proj.bg.rxCount[8] ),
    .X(net311));
 sg13g2_dlygate4sd3_1 hold295 (.A(\uart_proj.ren_wen_nidle[1] ),
    .X(net312));
 sg13g2_dlygate4sd3_1 hold296 (.A(_0235_),
    .X(net313));
 sg13g2_dlygate4sd3_1 hold297 (.A(\uart_proj.fifoRx.fifo[52] ),
    .X(net314));
 sg13g2_dlygate4sd3_1 hold298 (.A(_0219_),
    .X(net315));
 sg13g2_dlygate4sd3_1 hold299 (.A(\uart_proj.bg.rxCount[6] ),
    .X(net316));
 sg13g2_dlygate4sd3_1 hold300 (.A(_0036_),
    .X(net317));
 sg13g2_dlygate4sd3_1 hold301 (.A(\uart_proj.bg.rxCount[3] ),
    .X(net318));
 sg13g2_dlygate4sd3_1 hold302 (.A(\uart_proj.bg.rxCount[14] ),
    .X(net319));
 sg13g2_dlygate4sd3_1 hold303 (.A(\uart_proj.bg.rxCount[10] ),
    .X(net320));
 sg13g2_dlygate4sd3_1 hold304 (.A(_0734_),
    .X(net321));
 sg13g2_dlygate4sd3_1 hold305 (.A(_0254_),
    .X(net322));
 sg13g2_dlygate4sd3_1 hold306 (.A(\uart_proj.bg.txCount[14] ),
    .X(net323));
 sg13g2_dlygate4sd3_1 hold307 (.A(_0131_),
    .X(net324));
 sg13g2_dlygate4sd3_1 hold308 (.A(\uart_proj.bg.txCount[17] ),
    .X(net325));
 sg13g2_dlygate4sd3_1 hold309 (.A(_0134_),
    .X(net326));
 sg13g2_dlygate4sd3_1 hold310 (.A(\uart_proj.bg.txCount[19] ),
    .X(net327));
 sg13g2_dlygate4sd3_1 hold311 (.A(_0136_),
    .X(net328));
 sg13g2_dlygate4sd3_1 hold312 (.A(\uart_proj.uartTx.enterStart ),
    .X(net329));
 sg13g2_dlygate4sd3_1 hold313 (.A(_0765_),
    .X(net330));
 sg13g2_dlygate4sd3_1 hold314 (.A(_0028_),
    .X(net331));
 sg13g2_dlygate4sd3_1 hold315 (.A(_1193_),
    .X(net332));
 sg13g2_dlygate4sd3_1 hold316 (.A(\uart_proj.bg.rxCount[2] ),
    .X(net333));
 sg13g2_dlygate4sd3_1 hold317 (.A(_0246_),
    .X(net334));
 sg13g2_dlygate4sd3_1 hold318 (.A(\uart_proj.uartTx.curState[1] ),
    .X(net335));
 sg13g2_dlygate4sd3_1 hold319 (.A(_0956_),
    .X(net336));
 sg13g2_dlygate4sd3_1 hold320 (.A(_0000_),
    .X(net337));
 sg13g2_dlygate4sd3_1 hold321 (.A(\uart_proj.bg.txCount[18] ),
    .X(net338));
 sg13g2_dlygate4sd3_1 hold322 (.A(_0135_),
    .X(net339));
 sg13g2_dlygate4sd3_1 hold323 (.A(\uart_proj.bg.txCount[16] ),
    .X(net340));
 sg13g2_dlygate4sd3_1 hold324 (.A(_0133_),
    .X(net341));
 sg13g2_dlygate4sd3_1 hold325 (.A(\uart_proj.bg.rxCount[9] ),
    .X(net342));
 sg13g2_dlygate4sd3_1 hold326 (.A(\uart_proj.bg.txCount[15] ),
    .X(net343));
 sg13g2_dlygate4sd3_1 hold327 (.A(_0132_),
    .X(net344));
 sg13g2_dlygate4sd3_1 hold328 (.A(\uart_proj.fifoRx.write_ptr[2] ),
    .X(net345));
 sg13g2_dlygate4sd3_1 hold329 (.A(_0240_),
    .X(net346));
 sg13g2_dlygate4sd3_1 hold330 (.A(\uart_proj.uartTx.curState[2] ),
    .X(net347));
 sg13g2_dlygate4sd3_1 hold331 (.A(_0024_),
    .X(net348));
 sg13g2_dlygate4sd3_1 hold332 (.A(\uart_proj.uartRx.curState[2] ),
    .X(net349));
 sg13g2_dlygate4sd3_1 hold333 (.A(\uart_proj.uartTx.writeCount[0] ),
    .X(net350));
 sg13g2_dlygate4sd3_1 hold334 (.A(\uart_proj.uartTx.curState[3] ),
    .X(net351));
 sg13g2_dlygate4sd3_1 hold335 (.A(_0002_),
    .X(net352));
 sg13g2_dlygate4sd3_1 hold336 (.A(\uart_proj.bg.txCount[4] ),
    .X(net353));
 sg13g2_dlygate4sd3_1 hold337 (.A(_0140_),
    .X(net354));
 sg13g2_dlygate4sd3_1 hold338 (.A(_0091_),
    .X(net355));
 sg13g2_dlygate4sd3_1 hold339 (.A(_0465_),
    .X(net356));
 sg13g2_dlygate4sd3_1 hold340 (.A(_0466_),
    .X(net357));
 sg13g2_dlygate4sd3_1 hold341 (.A(_0022_),
    .X(net358));
 sg13g2_dlygate4sd3_1 hold342 (.A(_0043_),
    .X(net359));
 sg13g2_dlygate4sd3_1 hold343 (.A(_0420_),
    .X(net360));
 sg13g2_dlygate4sd3_1 hold344 (.A(_0421_),
    .X(net361));
 sg13g2_dlygate4sd3_1 hold345 (.A(_0016_),
    .X(net362));
 sg13g2_dlygate4sd3_1 hold346 (.A(\uart_proj.bg.rxCount[0] ),
    .X(net363));
 sg13g2_dlygate4sd3_1 hold347 (.A(_0244_),
    .X(net364));
 sg13g2_dlygate4sd3_1 hold348 (.A(_0051_),
    .X(net365));
 sg13g2_dlygate4sd3_1 hold349 (.A(_0428_),
    .X(net366));
 sg13g2_dlygate4sd3_1 hold350 (.A(_0429_),
    .X(net367));
 sg13g2_dlygate4sd3_1 hold351 (.A(_0017_),
    .X(net368));
 sg13g2_dlygate4sd3_1 hold352 (.A(\uart_proj.bg.rxCount[1] ),
    .X(net369));
 sg13g2_dlygate4sd3_1 hold353 (.A(_0038_),
    .X(net370));
 sg13g2_dlygate4sd3_1 hold354 (.A(_0031_),
    .X(net371));
 sg13g2_dlygate4sd3_1 hold355 (.A(_1211_),
    .X(net372));
 sg13g2_dlygate4sd3_1 hold356 (.A(_0099_),
    .X(net373));
 sg13g2_dlygate4sd3_1 hold357 (.A(_0477_),
    .X(net374));
 sg13g2_dlygate4sd3_1 hold358 (.A(_0478_),
    .X(net375));
 sg13g2_dlygate4sd3_1 hold359 (.A(_0023_),
    .X(net376));
 sg13g2_dlygate4sd3_1 hold360 (.A(\uart_proj.bg.txCount[13] ),
    .X(net377));
 sg13g2_dlygate4sd3_1 hold361 (.A(_0067_),
    .X(net378));
 sg13g2_dlygate4sd3_1 hold362 (.A(_0440_),
    .X(net379));
 sg13g2_dlygate4sd3_1 hold363 (.A(_0441_),
    .X(net380));
 sg13g2_dlygate4sd3_1 hold364 (.A(_0019_),
    .X(net381));
 sg13g2_dlygate4sd3_1 hold365 (.A(\uart_proj.uartRx.curState[1] ),
    .X(net382));
 sg13g2_dlygate4sd3_1 hold366 (.A(_0112_),
    .X(net383));
 sg13g2_dlygate4sd3_1 hold367 (.A(_0127_),
    .X(net384));
 sg13g2_dlygate4sd3_1 hold368 (.A(\uart_proj.bg.txCount[5] ),
    .X(net385));
 sg13g2_dlygate4sd3_1 hold369 (.A(_0575_),
    .X(net386));
 sg13g2_dlygate4sd3_1 hold370 (.A(_0060_),
    .X(net387));
 sg13g2_dlygate4sd3_1 hold371 (.A(_0436_),
    .X(net388));
 sg13g2_dlygate4sd3_1 hold372 (.A(_0437_),
    .X(net389));
 sg13g2_dlygate4sd3_1 hold373 (.A(_0018_),
    .X(net390));
 sg13g2_dlygate4sd3_1 hold374 (.A(\uart_proj.uartRx.curState[0] ),
    .X(net391));
 sg13g2_dlygate4sd3_1 hold375 (.A(_0075_),
    .X(net392));
 sg13g2_dlygate4sd3_1 hold376 (.A(_0448_),
    .X(net393));
 sg13g2_dlygate4sd3_1 hold377 (.A(_0449_),
    .X(net394));
 sg13g2_dlygate4sd3_1 hold378 (.A(_0020_),
    .X(net395));
 sg13g2_dlygate4sd3_1 hold379 (.A(\uart_proj.bg.txCount[8] ),
    .X(net396));
 sg13g2_dlygate4sd3_1 hold380 (.A(_0144_),
    .X(net397));
 sg13g2_dlygate4sd3_1 hold381 (.A(\uart_proj.fifoRx.count[3] ),
    .X(net398));
 sg13g2_dlygate4sd3_1 hold382 (.A(_0963_),
    .X(net399));
 sg13g2_dlygate4sd3_1 hold383 (.A(\uart_proj.fifoRx.count_next[3] ),
    .X(net400));
 sg13g2_dlygate4sd3_1 hold384 (.A(_0037_),
    .X(net529));
 sg13g2_dlygate4sd3_1 hold385 (.A(_0231_),
    .X(net530));
 sg13g2_dlygate4sd3_1 hold386 (.A(\uart_proj.bg.txCount[1] ),
    .X(net531));
 sg13g2_dlygate4sd3_1 hold387 (.A(\uart_proj.fifoRx.count[0] ),
    .X(net532));
 sg13g2_dlygate4sd3_1 hold388 (.A(_0377_),
    .X(net533));
 sg13g2_dlygate4sd3_1 hold389 (.A(\uart_proj.fifoRx.count_next[0] ),
    .X(net534));
 sg13g2_dlygate4sd3_1 hold390 (.A(_0123_),
    .X(net535));
 sg13g2_dlygate4sd3_1 hold391 (.A(_0034_),
    .X(net536));
 sg13g2_dlygate4sd3_1 hold392 (.A(\uart_proj.bg.txCount[7] ),
    .X(net537));
 sg13g2_dlygate4sd3_1 hold393 (.A(_0579_),
    .X(net538));
 sg13g2_dlygate4sd3_1 hold394 (.A(\uart_proj.bg.txCount[12] ),
    .X(net539));
 sg13g2_dlygate4sd3_1 hold395 (.A(_0129_),
    .X(net540));
 sg13g2_dlygate4sd3_1 hold396 (.A(\uart_proj.bg.txCount[2] ),
    .X(net541));
 sg13g2_dlygate4sd3_1 hold397 (.A(\uart_proj.ren_wen_nidle[0] ),
    .X(net542));
 sg13g2_dlygate4sd3_1 hold398 (.A(\uart_proj.fifoTx.count_next[3] ),
    .X(net543));
 sg13g2_dlygate4sd3_1 hold399 (.A(\uart_proj.fifoTx.write_ptr[2] ),
    .X(net544));
 sg13g2_dlygate4sd3_1 hold400 (.A(\uart_proj.fifoTx.write_ptr[1] ),
    .X(net545));
 sg13g2_dlygate4sd3_1 hold401 (.A(_0117_),
    .X(net546));
 sg13g2_dlygate4sd3_1 hold402 (.A(_0081_),
    .X(net547));
 sg13g2_dlygate4sd3_1 hold403 (.A(_0461_),
    .X(net548));
 sg13g2_dlygate4sd3_1 hold404 (.A(\uart_proj.bg.txCount[11] ),
    .X(net549));
 sg13g2_dlygate4sd3_1 hold405 (.A(\uart_proj.bg.txCount[9] ),
    .X(net550));
 sg13g2_dlygate4sd3_1 hold406 (.A(\uart_proj.bg.txCount[3] ),
    .X(net551));
 sg13g2_dlygate4sd3_1 hold407 (.A(\uart_proj.fifoRx.write_ptr[1] ),
    .X(net552));
 sg13g2_dlygate4sd3_1 hold408 (.A(_0239_),
    .X(net553));
 sg13g2_dlygate4sd3_1 hold409 (.A(\uart_proj.fifoTx.REN ),
    .X(net554));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_fill_2 FILLER_10_301 ();
 sg13g2_fill_1 FILLER_10_303 ();
 sg13g2_decap_8 FILLER_10_309 ();
 sg13g2_decap_8 FILLER_10_316 ();
 sg13g2_decap_8 FILLER_10_332 ();
 sg13g2_decap_8 FILLER_10_339 ();
 sg13g2_decap_8 FILLER_10_346 ();
 sg13g2_decap_8 FILLER_10_353 ();
 sg13g2_decap_8 FILLER_10_360 ();
 sg13g2_decap_8 FILLER_10_367 ();
 sg13g2_decap_8 FILLER_10_374 ();
 sg13g2_decap_8 FILLER_10_381 ();
 sg13g2_decap_8 FILLER_10_388 ();
 sg13g2_decap_8 FILLER_10_395 ();
 sg13g2_decap_8 FILLER_10_402 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_4 FILLER_11_294 ();
 sg13g2_fill_2 FILLER_11_298 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_4 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_377 ();
 sg13g2_decap_8 FILLER_12_384 ();
 sg13g2_decap_8 FILLER_12_391 ();
 sg13g2_decap_8 FILLER_12_398 ();
 sg13g2_decap_4 FILLER_12_405 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_fill_2 FILLER_13_259 ();
 sg13g2_fill_1 FILLER_13_261 ();
 sg13g2_decap_4 FILLER_13_288 ();
 sg13g2_fill_1 FILLER_13_292 ();
 sg13g2_fill_1 FILLER_13_301 ();
 sg13g2_fill_2 FILLER_13_354 ();
 sg13g2_fill_1 FILLER_13_356 ();
 sg13g2_decap_8 FILLER_13_379 ();
 sg13g2_decap_8 FILLER_13_386 ();
 sg13g2_decap_8 FILLER_13_393 ();
 sg13g2_decap_8 FILLER_13_400 ();
 sg13g2_fill_2 FILLER_13_407 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_4 FILLER_14_252 ();
 sg13g2_fill_1 FILLER_14_295 ();
 sg13g2_fill_2 FILLER_14_317 ();
 sg13g2_fill_2 FILLER_14_359 ();
 sg13g2_fill_1 FILLER_14_370 ();
 sg13g2_decap_8 FILLER_14_379 ();
 sg13g2_decap_8 FILLER_14_386 ();
 sg13g2_decap_8 FILLER_14_393 ();
 sg13g2_decap_8 FILLER_14_400 ();
 sg13g2_fill_2 FILLER_14_407 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_4 FILLER_15_238 ();
 sg13g2_fill_1 FILLER_15_242 ();
 sg13g2_fill_2 FILLER_15_279 ();
 sg13g2_fill_1 FILLER_15_320 ();
 sg13g2_fill_1 FILLER_15_346 ();
 sg13g2_decap_4 FILLER_15_357 ();
 sg13g2_decap_8 FILLER_15_397 ();
 sg13g2_decap_4 FILLER_15_404 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_decap_8 FILLER_16_217 ();
 sg13g2_decap_8 FILLER_16_224 ();
 sg13g2_decap_8 FILLER_16_231 ();
 sg13g2_decap_4 FILLER_16_238 ();
 sg13g2_fill_1 FILLER_16_242 ();
 sg13g2_fill_2 FILLER_16_334 ();
 sg13g2_fill_2 FILLER_16_348 ();
 sg13g2_fill_2 FILLER_16_358 ();
 sg13g2_fill_1 FILLER_16_360 ();
 sg13g2_decap_8 FILLER_16_401 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_decap_8 FILLER_17_168 ();
 sg13g2_decap_8 FILLER_17_175 ();
 sg13g2_decap_8 FILLER_17_182 ();
 sg13g2_decap_8 FILLER_17_189 ();
 sg13g2_decap_8 FILLER_17_196 ();
 sg13g2_decap_8 FILLER_17_203 ();
 sg13g2_decap_8 FILLER_17_210 ();
 sg13g2_decap_8 FILLER_17_217 ();
 sg13g2_decap_8 FILLER_17_224 ();
 sg13g2_decap_4 FILLER_17_231 ();
 sg13g2_fill_2 FILLER_17_282 ();
 sg13g2_fill_1 FILLER_17_294 ();
 sg13g2_fill_1 FILLER_17_304 ();
 sg13g2_fill_2 FILLER_17_331 ();
 sg13g2_decap_4 FILLER_17_370 ();
 sg13g2_decap_8 FILLER_17_400 ();
 sg13g2_fill_2 FILLER_17_407 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_decap_8 FILLER_18_147 ();
 sg13g2_decap_8 FILLER_18_154 ();
 sg13g2_decap_8 FILLER_18_161 ();
 sg13g2_decap_8 FILLER_18_168 ();
 sg13g2_decap_8 FILLER_18_175 ();
 sg13g2_decap_8 FILLER_18_182 ();
 sg13g2_decap_8 FILLER_18_189 ();
 sg13g2_decap_8 FILLER_18_196 ();
 sg13g2_decap_8 FILLER_18_203 ();
 sg13g2_decap_8 FILLER_18_210 ();
 sg13g2_decap_8 FILLER_18_217 ();
 sg13g2_decap_8 FILLER_18_224 ();
 sg13g2_fill_2 FILLER_18_231 ();
 sg13g2_fill_2 FILLER_18_267 ();
 sg13g2_fill_1 FILLER_18_269 ();
 sg13g2_fill_2 FILLER_18_288 ();
 sg13g2_fill_1 FILLER_18_290 ();
 sg13g2_fill_1 FILLER_18_309 ();
 sg13g2_fill_1 FILLER_18_388 ();
 sg13g2_decap_8 FILLER_18_398 ();
 sg13g2_decap_4 FILLER_18_405 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_decap_8 FILLER_19_140 ();
 sg13g2_decap_8 FILLER_19_147 ();
 sg13g2_decap_8 FILLER_19_154 ();
 sg13g2_decap_8 FILLER_19_161 ();
 sg13g2_decap_8 FILLER_19_168 ();
 sg13g2_decap_8 FILLER_19_175 ();
 sg13g2_decap_8 FILLER_19_182 ();
 sg13g2_decap_8 FILLER_19_189 ();
 sg13g2_decap_8 FILLER_19_196 ();
 sg13g2_decap_8 FILLER_19_203 ();
 sg13g2_decap_4 FILLER_19_210 ();
 sg13g2_fill_1 FILLER_19_214 ();
 sg13g2_fill_2 FILLER_19_274 ();
 sg13g2_fill_1 FILLER_19_276 ();
 sg13g2_fill_2 FILLER_19_358 ();
 sg13g2_decap_4 FILLER_19_368 ();
 sg13g2_fill_2 FILLER_19_372 ();
 sg13g2_decap_8 FILLER_19_387 ();
 sg13g2_decap_8 FILLER_19_394 ();
 sg13g2_decap_8 FILLER_19_401 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_decap_8 FILLER_20_126 ();
 sg13g2_decap_8 FILLER_20_133 ();
 sg13g2_decap_8 FILLER_20_140 ();
 sg13g2_decap_8 FILLER_20_147 ();
 sg13g2_decap_8 FILLER_20_154 ();
 sg13g2_decap_8 FILLER_20_161 ();
 sg13g2_decap_8 FILLER_20_168 ();
 sg13g2_decap_8 FILLER_20_175 ();
 sg13g2_decap_8 FILLER_20_182 ();
 sg13g2_decap_8 FILLER_20_189 ();
 sg13g2_decap_8 FILLER_20_196 ();
 sg13g2_fill_2 FILLER_20_203 ();
 sg13g2_fill_2 FILLER_20_236 ();
 sg13g2_fill_1 FILLER_20_333 ();
 sg13g2_decap_4 FILLER_20_351 ();
 sg13g2_fill_2 FILLER_20_355 ();
 sg13g2_decap_4 FILLER_20_403 ();
 sg13g2_fill_2 FILLER_20_407 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_decap_8 FILLER_21_119 ();
 sg13g2_decap_8 FILLER_21_126 ();
 sg13g2_decap_8 FILLER_21_133 ();
 sg13g2_decap_8 FILLER_21_140 ();
 sg13g2_decap_8 FILLER_21_147 ();
 sg13g2_decap_8 FILLER_21_154 ();
 sg13g2_decap_8 FILLER_21_161 ();
 sg13g2_decap_8 FILLER_21_168 ();
 sg13g2_decap_8 FILLER_21_175 ();
 sg13g2_decap_4 FILLER_21_182 ();
 sg13g2_decap_4 FILLER_21_279 ();
 sg13g2_fill_1 FILLER_21_283 ();
 sg13g2_fill_1 FILLER_21_330 ();
 sg13g2_fill_2 FILLER_21_343 ();
 sg13g2_fill_1 FILLER_21_345 ();
 sg13g2_decap_4 FILLER_21_404 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_8 FILLER_22_105 ();
 sg13g2_decap_8 FILLER_22_112 ();
 sg13g2_decap_8 FILLER_22_119 ();
 sg13g2_decap_8 FILLER_22_126 ();
 sg13g2_decap_8 FILLER_22_133 ();
 sg13g2_decap_8 FILLER_22_140 ();
 sg13g2_decap_8 FILLER_22_147 ();
 sg13g2_decap_8 FILLER_22_154 ();
 sg13g2_decap_8 FILLER_22_161 ();
 sg13g2_decap_8 FILLER_22_168 ();
 sg13g2_decap_8 FILLER_22_175 ();
 sg13g2_decap_4 FILLER_22_182 ();
 sg13g2_fill_1 FILLER_22_212 ();
 sg13g2_fill_2 FILLER_22_266 ();
 sg13g2_fill_2 FILLER_22_292 ();
 sg13g2_fill_1 FILLER_22_294 ();
 sg13g2_fill_2 FILLER_22_315 ();
 sg13g2_fill_1 FILLER_22_317 ();
 sg13g2_fill_2 FILLER_22_343 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_98 ();
 sg13g2_decap_8 FILLER_23_105 ();
 sg13g2_decap_8 FILLER_23_112 ();
 sg13g2_decap_8 FILLER_23_119 ();
 sg13g2_decap_8 FILLER_23_126 ();
 sg13g2_decap_8 FILLER_23_133 ();
 sg13g2_decap_8 FILLER_23_140 ();
 sg13g2_decap_8 FILLER_23_147 ();
 sg13g2_decap_8 FILLER_23_154 ();
 sg13g2_decap_8 FILLER_23_161 ();
 sg13g2_decap_8 FILLER_23_168 ();
 sg13g2_decap_4 FILLER_23_175 ();
 sg13g2_fill_1 FILLER_23_179 ();
 sg13g2_fill_2 FILLER_23_274 ();
 sg13g2_fill_1 FILLER_23_276 ();
 sg13g2_fill_1 FILLER_23_309 ();
 sg13g2_decap_8 FILLER_23_326 ();
 sg13g2_decap_8 FILLER_23_333 ();
 sg13g2_fill_1 FILLER_23_340 ();
 sg13g2_decap_8 FILLER_23_345 ();
 sg13g2_fill_2 FILLER_23_352 ();
 sg13g2_decap_8 FILLER_23_361 ();
 sg13g2_fill_2 FILLER_23_368 ();
 sg13g2_fill_1 FILLER_23_370 ();
 sg13g2_decap_8 FILLER_23_375 ();
 sg13g2_fill_2 FILLER_23_382 ();
 sg13g2_decap_8 FILLER_23_402 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_decap_8 FILLER_24_98 ();
 sg13g2_decap_8 FILLER_24_105 ();
 sg13g2_decap_8 FILLER_24_112 ();
 sg13g2_decap_8 FILLER_24_119 ();
 sg13g2_decap_8 FILLER_24_126 ();
 sg13g2_decap_8 FILLER_24_133 ();
 sg13g2_decap_8 FILLER_24_140 ();
 sg13g2_decap_8 FILLER_24_147 ();
 sg13g2_decap_8 FILLER_24_154 ();
 sg13g2_decap_8 FILLER_24_161 ();
 sg13g2_decap_8 FILLER_24_168 ();
 sg13g2_decap_4 FILLER_24_175 ();
 sg13g2_fill_1 FILLER_24_179 ();
 sg13g2_fill_1 FILLER_24_199 ();
 sg13g2_fill_2 FILLER_24_214 ();
 sg13g2_fill_1 FILLER_24_216 ();
 sg13g2_fill_1 FILLER_24_231 ();
 sg13g2_fill_2 FILLER_24_236 ();
 sg13g2_fill_1 FILLER_24_238 ();
 sg13g2_fill_2 FILLER_24_248 ();
 sg13g2_fill_1 FILLER_24_250 ();
 sg13g2_fill_1 FILLER_24_277 ();
 sg13g2_decap_8 FILLER_24_321 ();
 sg13g2_fill_1 FILLER_24_328 ();
 sg13g2_decap_8 FILLER_24_338 ();
 sg13g2_fill_1 FILLER_24_345 ();
 sg13g2_fill_1 FILLER_24_361 ();
 sg13g2_fill_2 FILLER_24_366 ();
 sg13g2_fill_2 FILLER_24_377 ();
 sg13g2_fill_1 FILLER_24_382 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_8 FILLER_25_91 ();
 sg13g2_decap_8 FILLER_25_98 ();
 sg13g2_decap_8 FILLER_25_105 ();
 sg13g2_decap_8 FILLER_25_112 ();
 sg13g2_decap_8 FILLER_25_119 ();
 sg13g2_decap_8 FILLER_25_126 ();
 sg13g2_decap_8 FILLER_25_133 ();
 sg13g2_decap_8 FILLER_25_140 ();
 sg13g2_decap_8 FILLER_25_147 ();
 sg13g2_decap_8 FILLER_25_154 ();
 sg13g2_decap_8 FILLER_25_161 ();
 sg13g2_decap_8 FILLER_25_168 ();
 sg13g2_decap_8 FILLER_25_175 ();
 sg13g2_decap_4 FILLER_25_182 ();
 sg13g2_fill_2 FILLER_25_186 ();
 sg13g2_fill_2 FILLER_25_240 ();
 sg13g2_fill_1 FILLER_25_242 ();
 sg13g2_fill_1 FILLER_25_251 ();
 sg13g2_fill_2 FILLER_25_300 ();
 sg13g2_fill_1 FILLER_25_302 ();
 sg13g2_fill_1 FILLER_25_323 ();
 sg13g2_fill_2 FILLER_25_365 ();
 sg13g2_fill_1 FILLER_25_367 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_decap_8 FILLER_26_91 ();
 sg13g2_decap_8 FILLER_26_98 ();
 sg13g2_decap_8 FILLER_26_105 ();
 sg13g2_decap_8 FILLER_26_112 ();
 sg13g2_decap_8 FILLER_26_119 ();
 sg13g2_decap_8 FILLER_26_126 ();
 sg13g2_decap_8 FILLER_26_133 ();
 sg13g2_decap_8 FILLER_26_140 ();
 sg13g2_decap_8 FILLER_26_147 ();
 sg13g2_decap_8 FILLER_26_154 ();
 sg13g2_decap_8 FILLER_26_161 ();
 sg13g2_decap_8 FILLER_26_168 ();
 sg13g2_decap_8 FILLER_26_175 ();
 sg13g2_fill_2 FILLER_26_182 ();
 sg13g2_fill_2 FILLER_26_189 ();
 sg13g2_fill_1 FILLER_26_191 ();
 sg13g2_decap_8 FILLER_26_196 ();
 sg13g2_fill_1 FILLER_26_203 ();
 sg13g2_fill_2 FILLER_26_257 ();
 sg13g2_fill_1 FILLER_26_303 ();
 sg13g2_fill_1 FILLER_26_341 ();
 sg13g2_fill_2 FILLER_26_348 ();
 sg13g2_fill_1 FILLER_26_350 ();
 sg13g2_fill_2 FILLER_26_357 ();
 sg13g2_fill_2 FILLER_26_364 ();
 sg13g2_fill_1 FILLER_26_374 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_decap_8 FILLER_27_84 ();
 sg13g2_decap_8 FILLER_27_91 ();
 sg13g2_decap_8 FILLER_27_98 ();
 sg13g2_decap_8 FILLER_27_105 ();
 sg13g2_decap_4 FILLER_27_112 ();
 sg13g2_fill_2 FILLER_27_116 ();
 sg13g2_decap_8 FILLER_27_136 ();
 sg13g2_decap_8 FILLER_27_143 ();
 sg13g2_decap_8 FILLER_27_150 ();
 sg13g2_decap_8 FILLER_27_157 ();
 sg13g2_decap_8 FILLER_27_164 ();
 sg13g2_fill_2 FILLER_27_171 ();
 sg13g2_fill_1 FILLER_27_173 ();
 sg13g2_decap_4 FILLER_27_182 ();
 sg13g2_fill_2 FILLER_27_186 ();
 sg13g2_fill_2 FILLER_27_205 ();
 sg13g2_fill_2 FILLER_27_214 ();
 sg13g2_fill_2 FILLER_27_221 ();
 sg13g2_fill_1 FILLER_27_228 ();
 sg13g2_fill_2 FILLER_27_244 ();
 sg13g2_fill_1 FILLER_27_273 ();
 sg13g2_fill_1 FILLER_27_287 ();
 sg13g2_fill_2 FILLER_27_326 ();
 sg13g2_fill_1 FILLER_27_328 ();
 sg13g2_fill_2 FILLER_27_374 ();
 sg13g2_fill_2 FILLER_27_392 ();
 sg13g2_fill_1 FILLER_27_394 ();
 sg13g2_decap_4 FILLER_27_404 ();
 sg13g2_fill_1 FILLER_27_408 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_decap_8 FILLER_28_84 ();
 sg13g2_decap_8 FILLER_28_91 ();
 sg13g2_decap_4 FILLER_28_98 ();
 sg13g2_fill_2 FILLER_28_172 ();
 sg13g2_fill_1 FILLER_28_174 ();
 sg13g2_fill_1 FILLER_28_180 ();
 sg13g2_fill_1 FILLER_28_238 ();
 sg13g2_fill_2 FILLER_28_246 ();
 sg13g2_fill_1 FILLER_28_248 ();
 sg13g2_fill_1 FILLER_28_262 ();
 sg13g2_fill_1 FILLER_28_287 ();
 sg13g2_fill_2 FILLER_28_308 ();
 sg13g2_fill_1 FILLER_28_310 ();
 sg13g2_fill_2 FILLER_28_332 ();
 sg13g2_fill_1 FILLER_28_357 ();
 sg13g2_fill_2 FILLER_28_363 ();
 sg13g2_fill_2 FILLER_28_373 ();
 sg13g2_fill_1 FILLER_28_375 ();
 sg13g2_fill_2 FILLER_28_379 ();
 sg13g2_fill_1 FILLER_28_381 ();
 sg13g2_decap_8 FILLER_28_387 ();
 sg13g2_decap_4 FILLER_28_394 ();
 sg13g2_fill_2 FILLER_28_407 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_decap_8 FILLER_29_84 ();
 sg13g2_fill_2 FILLER_29_91 ();
 sg13g2_decap_4 FILLER_29_191 ();
 sg13g2_fill_2 FILLER_29_208 ();
 sg13g2_fill_1 FILLER_29_210 ();
 sg13g2_fill_1 FILLER_29_233 ();
 sg13g2_fill_1 FILLER_29_258 ();
 sg13g2_fill_2 FILLER_29_300 ();
 sg13g2_fill_2 FILLER_29_312 ();
 sg13g2_fill_1 FILLER_29_314 ();
 sg13g2_fill_2 FILLER_29_320 ();
 sg13g2_fill_1 FILLER_29_348 ();
 sg13g2_fill_1 FILLER_29_361 ();
 sg13g2_fill_2 FILLER_29_376 ();
 sg13g2_decap_4 FILLER_29_391 ();
 sg13g2_fill_2 FILLER_29_395 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_77 ();
 sg13g2_decap_4 FILLER_30_84 ();
 sg13g2_fill_2 FILLER_30_114 ();
 sg13g2_fill_1 FILLER_30_141 ();
 sg13g2_decap_8 FILLER_30_183 ();
 sg13g2_decap_8 FILLER_30_190 ();
 sg13g2_decap_8 FILLER_30_197 ();
 sg13g2_fill_1 FILLER_30_204 ();
 sg13g2_fill_1 FILLER_30_240 ();
 sg13g2_fill_2 FILLER_30_280 ();
 sg13g2_fill_1 FILLER_30_282 ();
 sg13g2_fill_2 FILLER_30_300 ();
 sg13g2_fill_2 FILLER_30_307 ();
 sg13g2_fill_2 FILLER_30_350 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_decap_4 FILLER_31_84 ();
 sg13g2_fill_2 FILLER_31_88 ();
 sg13g2_fill_1 FILLER_31_126 ();
 sg13g2_fill_2 FILLER_31_137 ();
 sg13g2_fill_2 FILLER_31_227 ();
 sg13g2_fill_2 FILLER_31_253 ();
 sg13g2_fill_1 FILLER_31_255 ();
 sg13g2_fill_1 FILLER_31_268 ();
 sg13g2_fill_2 FILLER_31_278 ();
 sg13g2_fill_2 FILLER_31_324 ();
 sg13g2_decap_8 FILLER_31_340 ();
 sg13g2_fill_2 FILLER_31_347 ();
 sg13g2_decap_8 FILLER_31_353 ();
 sg13g2_fill_2 FILLER_31_360 ();
 sg13g2_fill_1 FILLER_31_362 ();
 sg13g2_fill_1 FILLER_31_377 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_8 FILLER_32_84 ();
 sg13g2_decap_8 FILLER_32_91 ();
 sg13g2_decap_4 FILLER_32_98 ();
 sg13g2_fill_1 FILLER_32_102 ();
 sg13g2_fill_2 FILLER_32_148 ();
 sg13g2_fill_2 FILLER_32_221 ();
 sg13g2_fill_2 FILLER_32_229 ();
 sg13g2_fill_1 FILLER_32_231 ();
 sg13g2_decap_4 FILLER_32_252 ();
 sg13g2_fill_2 FILLER_32_256 ();
 sg13g2_decap_8 FILLER_32_267 ();
 sg13g2_decap_4 FILLER_32_274 ();
 sg13g2_fill_2 FILLER_32_281 ();
 sg13g2_decap_8 FILLER_32_331 ();
 sg13g2_decap_4 FILLER_32_338 ();
 sg13g2_fill_2 FILLER_32_342 ();
 sg13g2_decap_8 FILLER_32_365 ();
 sg13g2_decap_8 FILLER_32_372 ();
 sg13g2_fill_2 FILLER_32_379 ();
 sg13g2_decap_4 FILLER_32_386 ();
 sg13g2_fill_1 FILLER_32_390 ();
 sg13g2_fill_1 FILLER_32_396 ();
 sg13g2_decap_4 FILLER_32_403 ();
 sg13g2_fill_2 FILLER_32_407 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_4 FILLER_33_84 ();
 sg13g2_fill_1 FILLER_33_88 ();
 sg13g2_fill_2 FILLER_33_173 ();
 sg13g2_fill_2 FILLER_33_192 ();
 sg13g2_fill_2 FILLER_33_241 ();
 sg13g2_fill_1 FILLER_33_243 ();
 sg13g2_fill_2 FILLER_33_291 ();
 sg13g2_fill_2 FILLER_33_324 ();
 sg13g2_fill_1 FILLER_33_326 ();
 sg13g2_decap_4 FILLER_33_375 ();
 sg13g2_fill_2 FILLER_33_379 ();
 sg13g2_decap_4 FILLER_33_404 ();
 sg13g2_fill_1 FILLER_33_408 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_fill_2 FILLER_34_77 ();
 sg13g2_fill_1 FILLER_34_79 ();
 sg13g2_fill_2 FILLER_34_125 ();
 sg13g2_fill_1 FILLER_34_221 ();
 sg13g2_fill_2 FILLER_34_317 ();
 sg13g2_fill_2 FILLER_34_355 ();
 sg13g2_fill_1 FILLER_34_408 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_fill_2 FILLER_35_84 ();
 sg13g2_fill_2 FILLER_35_124 ();
 sg13g2_fill_1 FILLER_35_126 ();
 sg13g2_fill_1 FILLER_35_167 ();
 sg13g2_fill_2 FILLER_35_216 ();
 sg13g2_fill_1 FILLER_35_218 ();
 sg13g2_fill_2 FILLER_35_224 ();
 sg13g2_fill_1 FILLER_35_264 ();
 sg13g2_decap_4 FILLER_35_346 ();
 sg13g2_fill_2 FILLER_35_375 ();
 sg13g2_fill_2 FILLER_35_394 ();
 sg13g2_fill_1 FILLER_35_396 ();
 sg13g2_fill_2 FILLER_35_407 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_fill_1 FILLER_36_91 ();
 sg13g2_fill_2 FILLER_36_158 ();
 sg13g2_fill_1 FILLER_36_160 ();
 sg13g2_fill_1 FILLER_36_190 ();
 sg13g2_fill_2 FILLER_36_242 ();
 sg13g2_fill_2 FILLER_36_258 ();
 sg13g2_fill_2 FILLER_36_269 ();
 sg13g2_fill_1 FILLER_36_271 ();
 sg13g2_fill_2 FILLER_36_282 ();
 sg13g2_fill_1 FILLER_36_301 ();
 sg13g2_decap_8 FILLER_36_328 ();
 sg13g2_decap_8 FILLER_36_335 ();
 sg13g2_decap_8 FILLER_36_342 ();
 sg13g2_decap_8 FILLER_36_349 ();
 sg13g2_decap_8 FILLER_36_361 ();
 sg13g2_fill_2 FILLER_36_368 ();
 sg13g2_decap_8 FILLER_36_375 ();
 sg13g2_decap_8 FILLER_36_382 ();
 sg13g2_fill_1 FILLER_36_408 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_4 FILLER_37_91 ();
 sg13g2_fill_1 FILLER_37_135 ();
 sg13g2_fill_2 FILLER_37_193 ();
 sg13g2_fill_1 FILLER_37_195 ();
 sg13g2_fill_1 FILLER_37_236 ();
 sg13g2_fill_1 FILLER_37_266 ();
 sg13g2_decap_4 FILLER_37_272 ();
 sg13g2_fill_1 FILLER_37_276 ();
 sg13g2_decap_4 FILLER_37_303 ();
 sg13g2_fill_2 FILLER_37_311 ();
 sg13g2_decap_4 FILLER_37_370 ();
 sg13g2_fill_1 FILLER_37_374 ();
 sg13g2_decap_4 FILLER_37_380 ();
 sg13g2_fill_2 FILLER_37_389 ();
 sg13g2_fill_1 FILLER_37_391 ();
 sg13g2_fill_2 FILLER_37_407 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_8 FILLER_38_56 ();
 sg13g2_decap_8 FILLER_38_63 ();
 sg13g2_decap_8 FILLER_38_70 ();
 sg13g2_decap_8 FILLER_38_77 ();
 sg13g2_decap_8 FILLER_38_84 ();
 sg13g2_decap_8 FILLER_38_91 ();
 sg13g2_fill_2 FILLER_38_98 ();
 sg13g2_decap_4 FILLER_38_135 ();
 sg13g2_decap_8 FILLER_38_184 ();
 sg13g2_fill_1 FILLER_38_191 ();
 sg13g2_fill_2 FILLER_38_197 ();
 sg13g2_decap_8 FILLER_38_272 ();
 sg13g2_fill_1 FILLER_38_279 ();
 sg13g2_decap_4 FILLER_38_289 ();
 sg13g2_fill_2 FILLER_38_293 ();
 sg13g2_decap_8 FILLER_38_300 ();
 sg13g2_decap_8 FILLER_38_307 ();
 sg13g2_decap_8 FILLER_38_314 ();
 sg13g2_fill_1 FILLER_38_321 ();
 sg13g2_fill_2 FILLER_38_327 ();
 sg13g2_fill_2 FILLER_38_406 ();
 sg13g2_fill_1 FILLER_38_408 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_14 ();
 sg13g2_decap_8 FILLER_39_21 ();
 sg13g2_decap_8 FILLER_39_28 ();
 sg13g2_decap_8 FILLER_39_35 ();
 sg13g2_decap_8 FILLER_39_42 ();
 sg13g2_decap_8 FILLER_39_49 ();
 sg13g2_decap_8 FILLER_39_56 ();
 sg13g2_decap_8 FILLER_39_63 ();
 sg13g2_decap_8 FILLER_39_70 ();
 sg13g2_decap_8 FILLER_39_77 ();
 sg13g2_decap_8 FILLER_39_84 ();
 sg13g2_decap_8 FILLER_39_91 ();
 sg13g2_decap_4 FILLER_39_98 ();
 sg13g2_fill_1 FILLER_39_102 ();
 sg13g2_decap_8 FILLER_39_108 ();
 sg13g2_decap_4 FILLER_39_115 ();
 sg13g2_fill_2 FILLER_39_119 ();
 sg13g2_fill_2 FILLER_39_163 ();
 sg13g2_fill_1 FILLER_39_165 ();
 sg13g2_fill_1 FILLER_39_175 ();
 sg13g2_decap_8 FILLER_39_194 ();
 sg13g2_fill_1 FILLER_39_201 ();
 sg13g2_fill_2 FILLER_39_215 ();
 sg13g2_fill_2 FILLER_39_231 ();
 sg13g2_fill_1 FILLER_39_259 ();
 sg13g2_decap_8 FILLER_39_274 ();
 sg13g2_decap_8 FILLER_39_281 ();
 sg13g2_fill_2 FILLER_39_288 ();
 sg13g2_fill_1 FILLER_39_290 ();
 sg13g2_decap_4 FILLER_39_322 ();
 sg13g2_fill_2 FILLER_39_326 ();
 sg13g2_decap_4 FILLER_39_359 ();
 sg13g2_fill_2 FILLER_39_407 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_14 ();
 sg13g2_decap_8 FILLER_40_21 ();
 sg13g2_decap_8 FILLER_40_28 ();
 sg13g2_decap_8 FILLER_40_35 ();
 sg13g2_decap_8 FILLER_40_42 ();
 sg13g2_decap_8 FILLER_40_49 ();
 sg13g2_decap_8 FILLER_40_56 ();
 sg13g2_decap_8 FILLER_40_63 ();
 sg13g2_decap_8 FILLER_40_70 ();
 sg13g2_decap_8 FILLER_40_77 ();
 sg13g2_decap_8 FILLER_40_84 ();
 sg13g2_decap_8 FILLER_40_91 ();
 sg13g2_decap_4 FILLER_40_134 ();
 sg13g2_decap_8 FILLER_40_204 ();
 sg13g2_fill_1 FILLER_40_211 ();
 sg13g2_decap_8 FILLER_40_237 ();
 sg13g2_decap_8 FILLER_40_244 ();
 sg13g2_decap_8 FILLER_40_251 ();
 sg13g2_fill_2 FILLER_40_258 ();
 sg13g2_fill_1 FILLER_40_260 ();
 sg13g2_decap_8 FILLER_40_326 ();
 sg13g2_decap_8 FILLER_40_333 ();
 sg13g2_decap_8 FILLER_40_340 ();
 sg13g2_decap_8 FILLER_40_347 ();
 sg13g2_decap_8 FILLER_40_354 ();
 sg13g2_decap_4 FILLER_40_361 ();
 sg13g2_fill_1 FILLER_40_365 ();
 sg13g2_fill_2 FILLER_40_370 ();
 sg13g2_fill_2 FILLER_40_389 ();
 sg13g2_fill_1 FILLER_40_391 ();
 sg13g2_decap_8 FILLER_40_402 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_8 FILLER_41_14 ();
 sg13g2_decap_8 FILLER_41_21 ();
 sg13g2_decap_8 FILLER_41_28 ();
 sg13g2_decap_8 FILLER_41_35 ();
 sg13g2_decap_8 FILLER_41_42 ();
 sg13g2_decap_8 FILLER_41_49 ();
 sg13g2_decap_8 FILLER_41_56 ();
 sg13g2_decap_8 FILLER_41_63 ();
 sg13g2_decap_8 FILLER_41_70 ();
 sg13g2_decap_8 FILLER_41_77 ();
 sg13g2_decap_8 FILLER_41_84 ();
 sg13g2_decap_8 FILLER_41_91 ();
 sg13g2_decap_4 FILLER_41_98 ();
 sg13g2_fill_2 FILLER_41_199 ();
 sg13g2_fill_2 FILLER_41_210 ();
 sg13g2_fill_1 FILLER_41_221 ();
 sg13g2_fill_2 FILLER_41_226 ();
 sg13g2_fill_1 FILLER_41_228 ();
 sg13g2_fill_1 FILLER_41_234 ();
 sg13g2_decap_4 FILLER_41_254 ();
 sg13g2_fill_1 FILLER_41_258 ();
 sg13g2_decap_8 FILLER_41_336 ();
 sg13g2_decap_4 FILLER_41_343 ();
 sg13g2_fill_1 FILLER_41_347 ();
 sg13g2_fill_2 FILLER_41_358 ();
 sg13g2_decap_8 FILLER_41_377 ();
 sg13g2_decap_8 FILLER_41_384 ();
 sg13g2_decap_8 FILLER_41_391 ();
 sg13g2_decap_8 FILLER_41_398 ();
 sg13g2_decap_4 FILLER_41_405 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_decap_8 FILLER_42_14 ();
 sg13g2_decap_8 FILLER_42_21 ();
 sg13g2_decap_8 FILLER_42_28 ();
 sg13g2_decap_8 FILLER_42_35 ();
 sg13g2_decap_8 FILLER_42_42 ();
 sg13g2_decap_8 FILLER_42_49 ();
 sg13g2_decap_8 FILLER_42_56 ();
 sg13g2_decap_8 FILLER_42_63 ();
 sg13g2_decap_8 FILLER_42_70 ();
 sg13g2_decap_8 FILLER_42_77 ();
 sg13g2_decap_8 FILLER_42_84 ();
 sg13g2_decap_8 FILLER_42_91 ();
 sg13g2_fill_2 FILLER_42_98 ();
 sg13g2_fill_1 FILLER_42_100 ();
 sg13g2_fill_2 FILLER_42_165 ();
 sg13g2_fill_1 FILLER_42_167 ();
 sg13g2_fill_2 FILLER_42_219 ();
 sg13g2_fill_1 FILLER_42_221 ();
 sg13g2_fill_2 FILLER_42_310 ();
 sg13g2_decap_8 FILLER_42_365 ();
 sg13g2_fill_1 FILLER_42_372 ();
 sg13g2_decap_8 FILLER_42_381 ();
 sg13g2_decap_8 FILLER_42_388 ();
 sg13g2_decap_8 FILLER_42_395 ();
 sg13g2_decap_8 FILLER_42_402 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_decap_8 FILLER_43_14 ();
 sg13g2_decap_8 FILLER_43_21 ();
 sg13g2_decap_8 FILLER_43_28 ();
 sg13g2_decap_8 FILLER_43_35 ();
 sg13g2_decap_8 FILLER_43_42 ();
 sg13g2_decap_8 FILLER_43_49 ();
 sg13g2_decap_8 FILLER_43_56 ();
 sg13g2_decap_8 FILLER_43_63 ();
 sg13g2_decap_8 FILLER_43_70 ();
 sg13g2_decap_8 FILLER_43_77 ();
 sg13g2_decap_8 FILLER_43_84 ();
 sg13g2_fill_1 FILLER_43_91 ();
 sg13g2_decap_4 FILLER_43_118 ();
 sg13g2_fill_1 FILLER_43_122 ();
 sg13g2_fill_2 FILLER_43_168 ();
 sg13g2_fill_2 FILLER_43_242 ();
 sg13g2_fill_1 FILLER_43_244 ();
 sg13g2_fill_2 FILLER_43_271 ();
 sg13g2_fill_1 FILLER_43_273 ();
 sg13g2_fill_2 FILLER_43_288 ();
 sg13g2_fill_1 FILLER_43_290 ();
 sg13g2_fill_2 FILLER_43_360 ();
 sg13g2_decap_8 FILLER_43_377 ();
 sg13g2_decap_8 FILLER_43_384 ();
 sg13g2_decap_8 FILLER_43_391 ();
 sg13g2_decap_8 FILLER_43_398 ();
 sg13g2_decap_4 FILLER_43_405 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_decap_8 FILLER_44_14 ();
 sg13g2_decap_8 FILLER_44_21 ();
 sg13g2_decap_8 FILLER_44_28 ();
 sg13g2_decap_8 FILLER_44_35 ();
 sg13g2_decap_8 FILLER_44_42 ();
 sg13g2_decap_8 FILLER_44_49 ();
 sg13g2_decap_8 FILLER_44_56 ();
 sg13g2_decap_8 FILLER_44_63 ();
 sg13g2_decap_8 FILLER_44_70 ();
 sg13g2_decap_8 FILLER_44_77 ();
 sg13g2_decap_8 FILLER_44_84 ();
 sg13g2_decap_4 FILLER_44_91 ();
 sg13g2_decap_4 FILLER_44_131 ();
 sg13g2_fill_1 FILLER_44_163 ();
 sg13g2_fill_2 FILLER_44_193 ();
 sg13g2_fill_2 FILLER_44_205 ();
 sg13g2_fill_2 FILLER_44_265 ();
 sg13g2_fill_2 FILLER_44_296 ();
 sg13g2_fill_1 FILLER_44_298 ();
 sg13g2_fill_2 FILLER_44_334 ();
 sg13g2_decap_4 FILLER_44_397 ();
 sg13g2_fill_1 FILLER_44_401 ();
 sg13g2_fill_2 FILLER_44_406 ();
 sg13g2_fill_1 FILLER_44_408 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_7 ();
 sg13g2_decap_8 FILLER_45_14 ();
 sg13g2_decap_8 FILLER_45_21 ();
 sg13g2_decap_8 FILLER_45_28 ();
 sg13g2_decap_8 FILLER_45_35 ();
 sg13g2_decap_8 FILLER_45_42 ();
 sg13g2_decap_8 FILLER_45_49 ();
 sg13g2_decap_8 FILLER_45_56 ();
 sg13g2_decap_8 FILLER_45_63 ();
 sg13g2_decap_8 FILLER_45_70 ();
 sg13g2_decap_8 FILLER_45_77 ();
 sg13g2_decap_4 FILLER_45_122 ();
 sg13g2_decap_4 FILLER_45_152 ();
 sg13g2_fill_2 FILLER_45_186 ();
 sg13g2_fill_1 FILLER_45_188 ();
 sg13g2_fill_2 FILLER_45_198 ();
 sg13g2_decap_4 FILLER_45_225 ();
 sg13g2_fill_1 FILLER_45_229 ();
 sg13g2_decap_8 FILLER_45_238 ();
 sg13g2_fill_1 FILLER_45_317 ();
 sg13g2_fill_2 FILLER_45_327 ();
 sg13g2_fill_1 FILLER_45_336 ();
 sg13g2_fill_1 FILLER_45_367 ();
 sg13g2_fill_2 FILLER_45_399 ();
 sg13g2_fill_1 FILLER_45_401 ();
 sg13g2_fill_2 FILLER_45_406 ();
 sg13g2_fill_1 FILLER_45_408 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_7 ();
 sg13g2_decap_8 FILLER_46_14 ();
 sg13g2_decap_8 FILLER_46_21 ();
 sg13g2_decap_8 FILLER_46_28 ();
 sg13g2_decap_8 FILLER_46_35 ();
 sg13g2_decap_8 FILLER_46_42 ();
 sg13g2_decap_8 FILLER_46_49 ();
 sg13g2_decap_8 FILLER_46_56 ();
 sg13g2_decap_8 FILLER_46_63 ();
 sg13g2_decap_8 FILLER_46_70 ();
 sg13g2_decap_8 FILLER_46_77 ();
 sg13g2_decap_8 FILLER_46_84 ();
 sg13g2_fill_2 FILLER_46_91 ();
 sg13g2_fill_1 FILLER_46_172 ();
 sg13g2_decap_8 FILLER_46_222 ();
 sg13g2_decap_8 FILLER_46_229 ();
 sg13g2_fill_1 FILLER_46_236 ();
 sg13g2_fill_2 FILLER_46_268 ();
 sg13g2_fill_1 FILLER_46_270 ();
 sg13g2_fill_2 FILLER_46_311 ();
 sg13g2_fill_1 FILLER_46_313 ();
 sg13g2_fill_2 FILLER_46_334 ();
 sg13g2_fill_1 FILLER_46_336 ();
 sg13g2_fill_2 FILLER_46_407 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_7 ();
 sg13g2_decap_8 FILLER_47_14 ();
 sg13g2_decap_8 FILLER_47_21 ();
 sg13g2_decap_8 FILLER_47_28 ();
 sg13g2_decap_8 FILLER_47_35 ();
 sg13g2_decap_8 FILLER_47_42 ();
 sg13g2_decap_8 FILLER_47_49 ();
 sg13g2_decap_8 FILLER_47_56 ();
 sg13g2_decap_8 FILLER_47_63 ();
 sg13g2_decap_8 FILLER_47_70 ();
 sg13g2_decap_4 FILLER_47_77 ();
 sg13g2_fill_2 FILLER_47_81 ();
 sg13g2_fill_1 FILLER_47_161 ();
 sg13g2_fill_1 FILLER_47_186 ();
 sg13g2_fill_1 FILLER_47_222 ();
 sg13g2_decap_4 FILLER_47_245 ();
 sg13g2_fill_2 FILLER_47_249 ();
 sg13g2_fill_2 FILLER_47_256 ();
 sg13g2_fill_1 FILLER_47_258 ();
 sg13g2_fill_2 FILLER_47_287 ();
 sg13g2_fill_2 FILLER_47_367 ();
 sg13g2_fill_2 FILLER_47_395 ();
 sg13g2_fill_1 FILLER_47_397 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_decap_8 FILLER_48_14 ();
 sg13g2_decap_8 FILLER_48_21 ();
 sg13g2_decap_8 FILLER_48_28 ();
 sg13g2_decap_8 FILLER_48_35 ();
 sg13g2_decap_8 FILLER_48_42 ();
 sg13g2_decap_8 FILLER_48_49 ();
 sg13g2_decap_8 FILLER_48_56 ();
 sg13g2_decap_8 FILLER_48_63 ();
 sg13g2_decap_4 FILLER_48_70 ();
 sg13g2_fill_2 FILLER_48_74 ();
 sg13g2_fill_2 FILLER_48_130 ();
 sg13g2_fill_1 FILLER_48_132 ();
 sg13g2_decap_4 FILLER_48_254 ();
 sg13g2_fill_2 FILLER_48_262 ();
 sg13g2_fill_1 FILLER_48_285 ();
 sg13g2_fill_1 FILLER_48_306 ();
 sg13g2_fill_1 FILLER_48_321 ();
 sg13g2_fill_2 FILLER_48_341 ();
 sg13g2_fill_1 FILLER_48_408 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_7 ();
 sg13g2_decap_8 FILLER_49_14 ();
 sg13g2_decap_8 FILLER_49_21 ();
 sg13g2_decap_8 FILLER_49_28 ();
 sg13g2_decap_8 FILLER_49_35 ();
 sg13g2_decap_8 FILLER_49_42 ();
 sg13g2_decap_8 FILLER_49_49 ();
 sg13g2_decap_8 FILLER_49_56 ();
 sg13g2_decap_8 FILLER_49_63 ();
 sg13g2_decap_8 FILLER_49_70 ();
 sg13g2_decap_8 FILLER_49_77 ();
 sg13g2_fill_2 FILLER_49_84 ();
 sg13g2_fill_2 FILLER_49_133 ();
 sg13g2_fill_2 FILLER_49_201 ();
 sg13g2_fill_2 FILLER_49_273 ();
 sg13g2_fill_2 FILLER_49_285 ();
 sg13g2_fill_2 FILLER_49_301 ();
 sg13g2_fill_1 FILLER_49_372 ();
 sg13g2_fill_1 FILLER_49_408 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_8 FILLER_50_7 ();
 sg13g2_decap_8 FILLER_50_14 ();
 sg13g2_decap_8 FILLER_50_21 ();
 sg13g2_decap_8 FILLER_50_28 ();
 sg13g2_decap_8 FILLER_50_35 ();
 sg13g2_decap_8 FILLER_50_42 ();
 sg13g2_decap_8 FILLER_50_49 ();
 sg13g2_decap_8 FILLER_50_56 ();
 sg13g2_decap_8 FILLER_50_63 ();
 sg13g2_decap_8 FILLER_50_70 ();
 sg13g2_decap_8 FILLER_50_77 ();
 sg13g2_decap_8 FILLER_50_84 ();
 sg13g2_fill_1 FILLER_50_91 ();
 sg13g2_fill_1 FILLER_50_123 ();
 sg13g2_fill_1 FILLER_50_139 ();
 sg13g2_fill_2 FILLER_50_193 ();
 sg13g2_fill_2 FILLER_50_213 ();
 sg13g2_fill_1 FILLER_50_233 ();
 sg13g2_fill_2 FILLER_50_243 ();
 sg13g2_fill_1 FILLER_50_315 ();
 sg13g2_fill_2 FILLER_50_334 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_decap_8 FILLER_51_7 ();
 sg13g2_decap_8 FILLER_51_14 ();
 sg13g2_decap_8 FILLER_51_21 ();
 sg13g2_decap_8 FILLER_51_28 ();
 sg13g2_decap_8 FILLER_51_35 ();
 sg13g2_decap_8 FILLER_51_42 ();
 sg13g2_decap_8 FILLER_51_49 ();
 sg13g2_decap_8 FILLER_51_56 ();
 sg13g2_decap_8 FILLER_51_63 ();
 sg13g2_decap_8 FILLER_51_70 ();
 sg13g2_decap_4 FILLER_51_77 ();
 sg13g2_fill_1 FILLER_51_81 ();
 sg13g2_fill_1 FILLER_51_154 ();
 sg13g2_fill_2 FILLER_51_234 ();
 sg13g2_fill_2 FILLER_51_250 ();
 sg13g2_fill_1 FILLER_51_252 ();
 sg13g2_fill_2 FILLER_51_305 ();
 sg13g2_fill_1 FILLER_51_307 ();
 sg13g2_fill_1 FILLER_51_338 ();
 sg13g2_fill_1 FILLER_51_365 ();
 sg13g2_fill_1 FILLER_51_408 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_decap_8 FILLER_52_7 ();
 sg13g2_decap_8 FILLER_52_14 ();
 sg13g2_decap_8 FILLER_52_21 ();
 sg13g2_decap_8 FILLER_52_28 ();
 sg13g2_decap_8 FILLER_52_35 ();
 sg13g2_decap_8 FILLER_52_42 ();
 sg13g2_decap_8 FILLER_52_49 ();
 sg13g2_decap_8 FILLER_52_56 ();
 sg13g2_decap_8 FILLER_52_63 ();
 sg13g2_decap_8 FILLER_52_70 ();
 sg13g2_decap_4 FILLER_52_77 ();
 sg13g2_fill_1 FILLER_52_122 ();
 sg13g2_fill_2 FILLER_52_132 ();
 sg13g2_fill_2 FILLER_52_142 ();
 sg13g2_fill_1 FILLER_52_212 ();
 sg13g2_decap_8 FILLER_52_236 ();
 sg13g2_decap_4 FILLER_52_243 ();
 sg13g2_fill_2 FILLER_52_247 ();
 sg13g2_fill_2 FILLER_52_254 ();
 sg13g2_fill_1 FILLER_52_256 ();
 sg13g2_fill_1 FILLER_52_310 ();
 sg13g2_fill_1 FILLER_52_324 ();
 sg13g2_fill_1 FILLER_52_342 ();
 sg13g2_fill_2 FILLER_52_367 ();
 sg13g2_fill_1 FILLER_52_408 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_decap_8 FILLER_53_7 ();
 sg13g2_decap_8 FILLER_53_14 ();
 sg13g2_decap_8 FILLER_53_21 ();
 sg13g2_decap_8 FILLER_53_28 ();
 sg13g2_decap_8 FILLER_53_35 ();
 sg13g2_decap_8 FILLER_53_42 ();
 sg13g2_decap_8 FILLER_53_49 ();
 sg13g2_decap_8 FILLER_53_56 ();
 sg13g2_decap_8 FILLER_53_63 ();
 sg13g2_decap_8 FILLER_53_70 ();
 sg13g2_fill_1 FILLER_53_77 ();
 sg13g2_fill_1 FILLER_53_142 ();
 sg13g2_fill_1 FILLER_53_157 ();
 sg13g2_fill_2 FILLER_53_184 ();
 sg13g2_fill_2 FILLER_53_231 ();
 sg13g2_fill_1 FILLER_53_233 ();
 sg13g2_fill_2 FILLER_53_250 ();
 sg13g2_fill_1 FILLER_53_252 ();
 sg13g2_decap_4 FILLER_53_257 ();
 sg13g2_fill_1 FILLER_53_261 ();
 sg13g2_fill_1 FILLER_53_276 ();
 sg13g2_decap_8 FILLER_53_286 ();
 sg13g2_fill_1 FILLER_53_293 ();
 sg13g2_fill_2 FILLER_53_299 ();
 sg13g2_fill_1 FILLER_53_314 ();
 sg13g2_fill_2 FILLER_53_337 ();
 sg13g2_fill_1 FILLER_53_365 ();
 sg13g2_fill_2 FILLER_53_393 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_decap_8 FILLER_54_7 ();
 sg13g2_decap_8 FILLER_54_14 ();
 sg13g2_decap_8 FILLER_54_21 ();
 sg13g2_decap_8 FILLER_54_28 ();
 sg13g2_decap_8 FILLER_54_35 ();
 sg13g2_decap_8 FILLER_54_42 ();
 sg13g2_decap_8 FILLER_54_49 ();
 sg13g2_decap_8 FILLER_54_56 ();
 sg13g2_decap_8 FILLER_54_63 ();
 sg13g2_decap_8 FILLER_54_70 ();
 sg13g2_decap_8 FILLER_54_77 ();
 sg13g2_fill_2 FILLER_54_157 ();
 sg13g2_fill_1 FILLER_54_159 ();
 sg13g2_fill_1 FILLER_54_186 ();
 sg13g2_fill_1 FILLER_54_282 ();
 sg13g2_fill_1 FILLER_54_289 ();
 sg13g2_fill_2 FILLER_54_301 ();
 sg13g2_fill_1 FILLER_54_303 ();
 sg13g2_fill_2 FILLER_54_322 ();
 sg13g2_fill_1 FILLER_54_324 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_decap_8 FILLER_55_7 ();
 sg13g2_decap_8 FILLER_55_14 ();
 sg13g2_decap_8 FILLER_55_21 ();
 sg13g2_decap_8 FILLER_55_28 ();
 sg13g2_decap_8 FILLER_55_35 ();
 sg13g2_decap_8 FILLER_55_42 ();
 sg13g2_decap_8 FILLER_55_49 ();
 sg13g2_decap_8 FILLER_55_56 ();
 sg13g2_decap_8 FILLER_55_63 ();
 sg13g2_decap_8 FILLER_55_70 ();
 sg13g2_decap_8 FILLER_55_77 ();
 sg13g2_fill_2 FILLER_55_84 ();
 sg13g2_fill_1 FILLER_55_86 ();
 sg13g2_fill_1 FILLER_55_165 ();
 sg13g2_fill_2 FILLER_55_184 ();
 sg13g2_fill_1 FILLER_55_186 ();
 sg13g2_fill_2 FILLER_55_213 ();
 sg13g2_fill_1 FILLER_55_229 ();
 sg13g2_decap_8 FILLER_55_251 ();
 sg13g2_decap_4 FILLER_55_258 ();
 sg13g2_fill_1 FILLER_55_262 ();
 sg13g2_fill_1 FILLER_55_286 ();
 sg13g2_fill_2 FILLER_55_302 ();
 sg13g2_fill_1 FILLER_55_304 ();
 sg13g2_fill_2 FILLER_55_310 ();
 sg13g2_fill_1 FILLER_55_312 ();
 sg13g2_fill_2 FILLER_55_380 ();
 sg13g2_fill_1 FILLER_55_382 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_decap_8 FILLER_56_7 ();
 sg13g2_decap_8 FILLER_56_14 ();
 sg13g2_decap_8 FILLER_56_21 ();
 sg13g2_decap_8 FILLER_56_28 ();
 sg13g2_decap_8 FILLER_56_35 ();
 sg13g2_decap_8 FILLER_56_42 ();
 sg13g2_decap_8 FILLER_56_49 ();
 sg13g2_decap_8 FILLER_56_56 ();
 sg13g2_decap_8 FILLER_56_63 ();
 sg13g2_decap_8 FILLER_56_70 ();
 sg13g2_decap_8 FILLER_56_77 ();
 sg13g2_decap_4 FILLER_56_84 ();
 sg13g2_fill_2 FILLER_56_111 ();
 sg13g2_fill_1 FILLER_56_113 ();
 sg13g2_fill_2 FILLER_56_177 ();
 sg13g2_fill_1 FILLER_56_211 ();
 sg13g2_fill_1 FILLER_56_236 ();
 sg13g2_fill_1 FILLER_56_263 ();
 sg13g2_fill_2 FILLER_56_320 ();
 sg13g2_fill_2 FILLER_56_406 ();
 sg13g2_fill_1 FILLER_56_408 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_decap_8 FILLER_57_7 ();
 sg13g2_decap_8 FILLER_57_14 ();
 sg13g2_decap_8 FILLER_57_21 ();
 sg13g2_decap_8 FILLER_57_28 ();
 sg13g2_decap_8 FILLER_57_35 ();
 sg13g2_decap_8 FILLER_57_42 ();
 sg13g2_decap_8 FILLER_57_49 ();
 sg13g2_decap_8 FILLER_57_56 ();
 sg13g2_decap_8 FILLER_57_63 ();
 sg13g2_decap_8 FILLER_57_70 ();
 sg13g2_decap_8 FILLER_57_77 ();
 sg13g2_decap_8 FILLER_57_84 ();
 sg13g2_fill_1 FILLER_57_91 ();
 sg13g2_fill_2 FILLER_57_119 ();
 sg13g2_fill_1 FILLER_57_121 ();
 sg13g2_fill_1 FILLER_57_161 ();
 sg13g2_fill_2 FILLER_57_184 ();
 sg13g2_fill_2 FILLER_57_201 ();
 sg13g2_fill_1 FILLER_57_259 ();
 sg13g2_fill_1 FILLER_57_282 ();
 sg13g2_fill_1 FILLER_57_312 ();
 sg13g2_fill_2 FILLER_57_363 ();
 sg13g2_fill_1 FILLER_57_365 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_decap_8 FILLER_58_7 ();
 sg13g2_decap_8 FILLER_58_14 ();
 sg13g2_decap_8 FILLER_58_21 ();
 sg13g2_decap_8 FILLER_58_28 ();
 sg13g2_decap_8 FILLER_58_35 ();
 sg13g2_decap_8 FILLER_58_42 ();
 sg13g2_decap_8 FILLER_58_49 ();
 sg13g2_decap_8 FILLER_58_56 ();
 sg13g2_decap_8 FILLER_58_63 ();
 sg13g2_decap_8 FILLER_58_70 ();
 sg13g2_decap_8 FILLER_58_77 ();
 sg13g2_decap_8 FILLER_58_84 ();
 sg13g2_fill_2 FILLER_58_91 ();
 sg13g2_fill_1 FILLER_58_128 ();
 sg13g2_fill_1 FILLER_58_142 ();
 sg13g2_fill_2 FILLER_58_160 ();
 sg13g2_fill_1 FILLER_58_162 ();
 sg13g2_decap_4 FILLER_58_241 ();
 sg13g2_fill_2 FILLER_58_249 ();
 sg13g2_fill_2 FILLER_58_290 ();
 sg13g2_fill_1 FILLER_58_292 ();
 sg13g2_fill_1 FILLER_58_339 ();
 sg13g2_fill_2 FILLER_58_345 ();
 sg13g2_fill_1 FILLER_58_368 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_decap_8 FILLER_59_7 ();
 sg13g2_decap_8 FILLER_59_14 ();
 sg13g2_decap_8 FILLER_59_21 ();
 sg13g2_decap_8 FILLER_59_28 ();
 sg13g2_decap_8 FILLER_59_35 ();
 sg13g2_decap_8 FILLER_59_42 ();
 sg13g2_decap_8 FILLER_59_49 ();
 sg13g2_decap_8 FILLER_59_56 ();
 sg13g2_decap_8 FILLER_59_63 ();
 sg13g2_decap_8 FILLER_59_70 ();
 sg13g2_decap_8 FILLER_59_77 ();
 sg13g2_decap_4 FILLER_59_84 ();
 sg13g2_fill_2 FILLER_59_88 ();
 sg13g2_fill_1 FILLER_59_143 ();
 sg13g2_fill_2 FILLER_59_203 ();
 sg13g2_fill_2 FILLER_59_223 ();
 sg13g2_fill_1 FILLER_59_225 ();
 sg13g2_decap_8 FILLER_59_231 ();
 sg13g2_decap_4 FILLER_59_238 ();
 sg13g2_fill_2 FILLER_59_242 ();
 sg13g2_fill_2 FILLER_59_257 ();
 sg13g2_fill_1 FILLER_59_259 ();
 sg13g2_fill_2 FILLER_59_284 ();
 sg13g2_fill_1 FILLER_59_292 ();
 sg13g2_fill_1 FILLER_59_392 ();
 sg13g2_fill_2 FILLER_59_398 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_decap_8 FILLER_60_7 ();
 sg13g2_decap_8 FILLER_60_14 ();
 sg13g2_decap_8 FILLER_60_21 ();
 sg13g2_decap_8 FILLER_60_28 ();
 sg13g2_decap_8 FILLER_60_35 ();
 sg13g2_decap_8 FILLER_60_42 ();
 sg13g2_decap_8 FILLER_60_49 ();
 sg13g2_decap_8 FILLER_60_56 ();
 sg13g2_decap_8 FILLER_60_63 ();
 sg13g2_decap_8 FILLER_60_70 ();
 sg13g2_decap_8 FILLER_60_77 ();
 sg13g2_decap_8 FILLER_60_84 ();
 sg13g2_fill_2 FILLER_60_91 ();
 sg13g2_fill_1 FILLER_60_93 ();
 sg13g2_fill_1 FILLER_60_114 ();
 sg13g2_fill_2 FILLER_60_157 ();
 sg13g2_fill_1 FILLER_60_199 ();
 sg13g2_decap_4 FILLER_60_226 ();
 sg13g2_fill_2 FILLER_60_230 ();
 sg13g2_fill_2 FILLER_60_319 ();
 sg13g2_fill_1 FILLER_60_321 ();
 sg13g2_fill_1 FILLER_60_357 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_decap_8 FILLER_61_7 ();
 sg13g2_decap_8 FILLER_61_14 ();
 sg13g2_decap_8 FILLER_61_21 ();
 sg13g2_decap_8 FILLER_61_28 ();
 sg13g2_decap_8 FILLER_61_35 ();
 sg13g2_decap_8 FILLER_61_42 ();
 sg13g2_decap_8 FILLER_61_49 ();
 sg13g2_decap_8 FILLER_61_56 ();
 sg13g2_decap_8 FILLER_61_63 ();
 sg13g2_decap_8 FILLER_61_70 ();
 sg13g2_decap_8 FILLER_61_77 ();
 sg13g2_fill_1 FILLER_61_84 ();
 sg13g2_fill_1 FILLER_61_113 ();
 sg13g2_fill_2 FILLER_61_123 ();
 sg13g2_fill_1 FILLER_61_125 ();
 sg13g2_fill_1 FILLER_61_156 ();
 sg13g2_fill_1 FILLER_61_163 ();
 sg13g2_fill_2 FILLER_61_213 ();
 sg13g2_fill_1 FILLER_61_224 ();
 sg13g2_fill_1 FILLER_61_280 ();
 sg13g2_fill_2 FILLER_61_295 ();
 sg13g2_fill_2 FILLER_61_307 ();
 sg13g2_fill_1 FILLER_61_309 ();
 sg13g2_fill_1 FILLER_61_320 ();
 sg13g2_fill_2 FILLER_61_326 ();
 sg13g2_fill_1 FILLER_61_328 ();
 sg13g2_fill_2 FILLER_61_407 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_decap_8 FILLER_62_7 ();
 sg13g2_decap_8 FILLER_62_14 ();
 sg13g2_decap_8 FILLER_62_21 ();
 sg13g2_decap_8 FILLER_62_28 ();
 sg13g2_decap_8 FILLER_62_35 ();
 sg13g2_decap_8 FILLER_62_42 ();
 sg13g2_decap_8 FILLER_62_49 ();
 sg13g2_decap_8 FILLER_62_56 ();
 sg13g2_decap_8 FILLER_62_63 ();
 sg13g2_decap_8 FILLER_62_70 ();
 sg13g2_decap_8 FILLER_62_77 ();
 sg13g2_fill_2 FILLER_62_84 ();
 sg13g2_fill_1 FILLER_62_86 ();
 sg13g2_fill_2 FILLER_62_117 ();
 sg13g2_fill_1 FILLER_62_119 ();
 sg13g2_fill_1 FILLER_62_241 ();
 sg13g2_fill_2 FILLER_62_287 ();
 sg13g2_fill_1 FILLER_62_324 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_decap_8 FILLER_63_7 ();
 sg13g2_decap_8 FILLER_63_14 ();
 sg13g2_decap_8 FILLER_63_21 ();
 sg13g2_decap_8 FILLER_63_28 ();
 sg13g2_decap_8 FILLER_63_35 ();
 sg13g2_decap_8 FILLER_63_42 ();
 sg13g2_decap_8 FILLER_63_49 ();
 sg13g2_decap_8 FILLER_63_56 ();
 sg13g2_decap_8 FILLER_63_63 ();
 sg13g2_decap_8 FILLER_63_70 ();
 sg13g2_decap_8 FILLER_63_77 ();
 sg13g2_decap_8 FILLER_63_84 ();
 sg13g2_fill_1 FILLER_63_91 ();
 sg13g2_fill_2 FILLER_63_146 ();
 sg13g2_fill_1 FILLER_63_148 ();
 sg13g2_fill_1 FILLER_63_162 ();
 sg13g2_fill_1 FILLER_63_261 ();
 sg13g2_fill_1 FILLER_63_297 ();
 sg13g2_fill_1 FILLER_63_357 ();
 sg13g2_fill_2 FILLER_63_407 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_8 FILLER_64_7 ();
 sg13g2_decap_8 FILLER_64_14 ();
 sg13g2_decap_8 FILLER_64_21 ();
 sg13g2_decap_8 FILLER_64_28 ();
 sg13g2_decap_8 FILLER_64_35 ();
 sg13g2_decap_8 FILLER_64_42 ();
 sg13g2_decap_8 FILLER_64_49 ();
 sg13g2_decap_8 FILLER_64_56 ();
 sg13g2_decap_8 FILLER_64_63 ();
 sg13g2_decap_8 FILLER_64_70 ();
 sg13g2_decap_8 FILLER_64_77 ();
 sg13g2_decap_8 FILLER_64_84 ();
 sg13g2_fill_1 FILLER_64_91 ();
 sg13g2_fill_2 FILLER_64_118 ();
 sg13g2_fill_2 FILLER_64_138 ();
 sg13g2_fill_1 FILLER_64_140 ();
 sg13g2_fill_2 FILLER_64_146 ();
 sg13g2_fill_1 FILLER_64_148 ();
 sg13g2_fill_1 FILLER_64_187 ();
 sg13g2_fill_2 FILLER_64_193 ();
 sg13g2_fill_1 FILLER_64_210 ();
 sg13g2_fill_1 FILLER_64_237 ();
 sg13g2_fill_1 FILLER_64_285 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_8 FILLER_65_7 ();
 sg13g2_decap_8 FILLER_65_14 ();
 sg13g2_decap_8 FILLER_65_21 ();
 sg13g2_decap_8 FILLER_65_28 ();
 sg13g2_decap_8 FILLER_65_35 ();
 sg13g2_decap_8 FILLER_65_42 ();
 sg13g2_decap_8 FILLER_65_49 ();
 sg13g2_decap_8 FILLER_65_56 ();
 sg13g2_decap_8 FILLER_65_63 ();
 sg13g2_decap_8 FILLER_65_70 ();
 sg13g2_decap_8 FILLER_65_77 ();
 sg13g2_decap_8 FILLER_65_84 ();
 sg13g2_decap_4 FILLER_65_91 ();
 sg13g2_fill_1 FILLER_65_104 ();
 sg13g2_fill_2 FILLER_65_118 ();
 sg13g2_fill_1 FILLER_65_120 ();
 sg13g2_fill_2 FILLER_65_239 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_8 FILLER_66_7 ();
 sg13g2_decap_8 FILLER_66_14 ();
 sg13g2_decap_8 FILLER_66_21 ();
 sg13g2_decap_8 FILLER_66_28 ();
 sg13g2_decap_8 FILLER_66_35 ();
 sg13g2_decap_8 FILLER_66_42 ();
 sg13g2_decap_8 FILLER_66_49 ();
 sg13g2_decap_8 FILLER_66_56 ();
 sg13g2_decap_8 FILLER_66_63 ();
 sg13g2_decap_8 FILLER_66_70 ();
 sg13g2_decap_8 FILLER_66_77 ();
 sg13g2_decap_8 FILLER_66_84 ();
 sg13g2_decap_8 FILLER_66_91 ();
 sg13g2_fill_2 FILLER_66_98 ();
 sg13g2_fill_1 FILLER_66_100 ();
 sg13g2_fill_1 FILLER_66_160 ();
 sg13g2_fill_2 FILLER_66_254 ();
 sg13g2_fill_1 FILLER_66_271 ();
 sg13g2_fill_2 FILLER_66_287 ();
 sg13g2_fill_2 FILLER_66_298 ();
 sg13g2_fill_1 FILLER_66_300 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_8 FILLER_67_7 ();
 sg13g2_decap_8 FILLER_67_14 ();
 sg13g2_decap_8 FILLER_67_21 ();
 sg13g2_decap_8 FILLER_67_28 ();
 sg13g2_decap_8 FILLER_67_35 ();
 sg13g2_decap_8 FILLER_67_42 ();
 sg13g2_decap_8 FILLER_67_49 ();
 sg13g2_decap_8 FILLER_67_56 ();
 sg13g2_decap_8 FILLER_67_63 ();
 sg13g2_decap_8 FILLER_67_70 ();
 sg13g2_decap_8 FILLER_67_77 ();
 sg13g2_decap_8 FILLER_67_84 ();
 sg13g2_decap_8 FILLER_67_91 ();
 sg13g2_fill_2 FILLER_67_149 ();
 sg13g2_fill_1 FILLER_67_151 ();
 sg13g2_fill_1 FILLER_67_220 ();
 sg13g2_fill_2 FILLER_67_244 ();
 sg13g2_fill_1 FILLER_67_331 ();
 sg13g2_fill_2 FILLER_67_340 ();
 sg13g2_fill_1 FILLER_67_342 ();
 sg13g2_fill_2 FILLER_67_386 ();
 sg13g2_fill_2 FILLER_67_393 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_8 FILLER_68_7 ();
 sg13g2_decap_8 FILLER_68_14 ();
 sg13g2_decap_8 FILLER_68_21 ();
 sg13g2_decap_8 FILLER_68_28 ();
 sg13g2_decap_8 FILLER_68_35 ();
 sg13g2_decap_8 FILLER_68_42 ();
 sg13g2_decap_8 FILLER_68_49 ();
 sg13g2_decap_8 FILLER_68_56 ();
 sg13g2_decap_8 FILLER_68_63 ();
 sg13g2_decap_8 FILLER_68_70 ();
 sg13g2_decap_8 FILLER_68_77 ();
 sg13g2_decap_8 FILLER_68_84 ();
 sg13g2_decap_8 FILLER_68_91 ();
 sg13g2_fill_2 FILLER_68_98 ();
 sg13g2_fill_1 FILLER_68_100 ();
 sg13g2_fill_2 FILLER_68_155 ();
 sg13g2_fill_1 FILLER_68_157 ();
 sg13g2_fill_1 FILLER_68_212 ();
 sg13g2_fill_1 FILLER_68_232 ();
 sg13g2_fill_2 FILLER_68_314 ();
 sg13g2_fill_1 FILLER_68_316 ();
 sg13g2_fill_2 FILLER_68_327 ();
 sg13g2_fill_1 FILLER_68_349 ();
 sg13g2_fill_2 FILLER_68_359 ();
 sg13g2_fill_2 FILLER_68_387 ();
 sg13g2_fill_2 FILLER_68_398 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_8 FILLER_69_7 ();
 sg13g2_decap_8 FILLER_69_14 ();
 sg13g2_decap_8 FILLER_69_21 ();
 sg13g2_decap_8 FILLER_69_28 ();
 sg13g2_decap_8 FILLER_69_35 ();
 sg13g2_decap_8 FILLER_69_42 ();
 sg13g2_decap_8 FILLER_69_49 ();
 sg13g2_decap_8 FILLER_69_56 ();
 sg13g2_decap_8 FILLER_69_63 ();
 sg13g2_decap_8 FILLER_69_70 ();
 sg13g2_decap_8 FILLER_69_77 ();
 sg13g2_decap_8 FILLER_69_84 ();
 sg13g2_decap_4 FILLER_69_91 ();
 sg13g2_fill_1 FILLER_69_181 ();
 sg13g2_fill_2 FILLER_69_340 ();
 sg13g2_fill_1 FILLER_69_382 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_decap_8 FILLER_70_14 ();
 sg13g2_decap_8 FILLER_70_21 ();
 sg13g2_decap_8 FILLER_70_28 ();
 sg13g2_decap_8 FILLER_70_35 ();
 sg13g2_decap_8 FILLER_70_42 ();
 sg13g2_decap_8 FILLER_70_49 ();
 sg13g2_decap_8 FILLER_70_56 ();
 sg13g2_decap_8 FILLER_70_63 ();
 sg13g2_decap_8 FILLER_70_70 ();
 sg13g2_decap_8 FILLER_70_77 ();
 sg13g2_decap_8 FILLER_70_84 ();
 sg13g2_fill_2 FILLER_70_91 ();
 sg13g2_fill_1 FILLER_70_93 ();
 sg13g2_fill_1 FILLER_70_128 ();
 sg13g2_fill_2 FILLER_70_170 ();
 sg13g2_fill_1 FILLER_70_190 ();
 sg13g2_fill_1 FILLER_70_236 ();
 sg13g2_fill_2 FILLER_70_253 ();
 sg13g2_fill_2 FILLER_70_275 ();
 sg13g2_fill_2 FILLER_70_323 ();
 sg13g2_fill_1 FILLER_70_334 ();
 sg13g2_fill_2 FILLER_70_353 ();
 sg13g2_fill_1 FILLER_70_388 ();
 sg13g2_fill_2 FILLER_70_398 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_decap_8 FILLER_71_7 ();
 sg13g2_decap_8 FILLER_71_14 ();
 sg13g2_decap_8 FILLER_71_21 ();
 sg13g2_decap_8 FILLER_71_28 ();
 sg13g2_decap_8 FILLER_71_35 ();
 sg13g2_decap_8 FILLER_71_42 ();
 sg13g2_decap_8 FILLER_71_49 ();
 sg13g2_decap_8 FILLER_71_56 ();
 sg13g2_decap_8 FILLER_71_63 ();
 sg13g2_decap_8 FILLER_71_70 ();
 sg13g2_decap_8 FILLER_71_77 ();
 sg13g2_decap_8 FILLER_71_84 ();
 sg13g2_decap_8 FILLER_71_91 ();
 sg13g2_fill_2 FILLER_71_98 ();
 sg13g2_fill_2 FILLER_71_140 ();
 sg13g2_fill_2 FILLER_71_191 ();
 sg13g2_fill_2 FILLER_71_204 ();
 sg13g2_fill_1 FILLER_71_214 ();
 sg13g2_fill_1 FILLER_71_245 ();
 sg13g2_fill_2 FILLER_71_269 ();
 sg13g2_fill_2 FILLER_71_350 ();
 sg13g2_fill_1 FILLER_71_408 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_decap_8 FILLER_72_14 ();
 sg13g2_decap_8 FILLER_72_21 ();
 sg13g2_decap_8 FILLER_72_28 ();
 sg13g2_decap_8 FILLER_72_35 ();
 sg13g2_decap_8 FILLER_72_42 ();
 sg13g2_decap_8 FILLER_72_49 ();
 sg13g2_decap_8 FILLER_72_56 ();
 sg13g2_decap_8 FILLER_72_63 ();
 sg13g2_decap_8 FILLER_72_70 ();
 sg13g2_decap_8 FILLER_72_77 ();
 sg13g2_decap_8 FILLER_72_84 ();
 sg13g2_decap_8 FILLER_72_91 ();
 sg13g2_decap_4 FILLER_72_98 ();
 sg13g2_fill_2 FILLER_72_102 ();
 sg13g2_fill_1 FILLER_72_222 ();
 sg13g2_fill_1 FILLER_72_244 ();
 sg13g2_fill_2 FILLER_72_299 ();
 sg13g2_fill_2 FILLER_72_345 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_decap_8 FILLER_73_14 ();
 sg13g2_decap_8 FILLER_73_21 ();
 sg13g2_decap_8 FILLER_73_28 ();
 sg13g2_decap_8 FILLER_73_35 ();
 sg13g2_decap_8 FILLER_73_42 ();
 sg13g2_decap_8 FILLER_73_49 ();
 sg13g2_decap_8 FILLER_73_56 ();
 sg13g2_decap_8 FILLER_73_63 ();
 sg13g2_decap_8 FILLER_73_70 ();
 sg13g2_decap_8 FILLER_73_77 ();
 sg13g2_decap_8 FILLER_73_84 ();
 sg13g2_decap_8 FILLER_73_91 ();
 sg13g2_fill_2 FILLER_73_98 ();
 sg13g2_fill_1 FILLER_73_100 ();
 sg13g2_fill_2 FILLER_73_134 ();
 sg13g2_fill_1 FILLER_73_136 ();
 sg13g2_fill_1 FILLER_73_156 ();
 sg13g2_fill_1 FILLER_73_221 ();
 sg13g2_fill_2 FILLER_73_307 ();
 sg13g2_fill_2 FILLER_73_314 ();
 sg13g2_fill_2 FILLER_73_381 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_decap_8 FILLER_74_14 ();
 sg13g2_decap_8 FILLER_74_21 ();
 sg13g2_decap_8 FILLER_74_28 ();
 sg13g2_decap_8 FILLER_74_35 ();
 sg13g2_decap_8 FILLER_74_42 ();
 sg13g2_decap_8 FILLER_74_49 ();
 sg13g2_decap_8 FILLER_74_56 ();
 sg13g2_decap_8 FILLER_74_63 ();
 sg13g2_decap_8 FILLER_74_70 ();
 sg13g2_decap_8 FILLER_74_77 ();
 sg13g2_decap_8 FILLER_74_84 ();
 sg13g2_decap_8 FILLER_74_91 ();
 sg13g2_fill_1 FILLER_74_98 ();
 sg13g2_fill_2 FILLER_74_139 ();
 sg13g2_fill_1 FILLER_74_141 ();
 sg13g2_fill_1 FILLER_74_173 ();
 sg13g2_fill_1 FILLER_74_194 ();
 sg13g2_fill_2 FILLER_74_259 ();
 sg13g2_fill_1 FILLER_74_261 ();
 sg13g2_fill_2 FILLER_74_271 ();
 sg13g2_fill_1 FILLER_74_273 ();
 sg13g2_fill_1 FILLER_74_303 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_14 ();
 sg13g2_decap_8 FILLER_75_21 ();
 sg13g2_decap_8 FILLER_75_28 ();
 sg13g2_decap_8 FILLER_75_35 ();
 sg13g2_decap_8 FILLER_75_42 ();
 sg13g2_decap_8 FILLER_75_49 ();
 sg13g2_decap_8 FILLER_75_56 ();
 sg13g2_decap_8 FILLER_75_63 ();
 sg13g2_decap_8 FILLER_75_70 ();
 sg13g2_decap_8 FILLER_75_77 ();
 sg13g2_decap_4 FILLER_75_84 ();
 sg13g2_fill_2 FILLER_75_88 ();
 sg13g2_fill_2 FILLER_75_117 ();
 sg13g2_fill_2 FILLER_75_156 ();
 sg13g2_fill_1 FILLER_75_167 ();
 sg13g2_fill_1 FILLER_75_191 ();
 sg13g2_fill_2 FILLER_75_212 ();
 sg13g2_fill_1 FILLER_75_214 ();
 sg13g2_fill_1 FILLER_75_267 ();
 sg13g2_fill_2 FILLER_75_320 ();
 sg13g2_fill_1 FILLER_75_322 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_8 FILLER_76_21 ();
 sg13g2_decap_8 FILLER_76_28 ();
 sg13g2_decap_8 FILLER_76_35 ();
 sg13g2_decap_8 FILLER_76_42 ();
 sg13g2_decap_8 FILLER_76_49 ();
 sg13g2_decap_8 FILLER_76_56 ();
 sg13g2_decap_8 FILLER_76_63 ();
 sg13g2_decap_8 FILLER_76_70 ();
 sg13g2_decap_8 FILLER_76_77 ();
 sg13g2_decap_8 FILLER_76_84 ();
 sg13g2_fill_2 FILLER_76_91 ();
 sg13g2_fill_1 FILLER_76_93 ();
 sg13g2_fill_2 FILLER_76_133 ();
 sg13g2_fill_1 FILLER_76_218 ();
 sg13g2_fill_2 FILLER_76_260 ();
 sg13g2_fill_2 FILLER_76_288 ();
 sg13g2_fill_1 FILLER_76_290 ();
 sg13g2_fill_1 FILLER_76_306 ();
 sg13g2_fill_2 FILLER_76_332 ();
 sg13g2_fill_2 FILLER_76_366 ();
 sg13g2_fill_2 FILLER_76_381 ();
 sg13g2_fill_1 FILLER_76_383 ();
 sg13g2_fill_2 FILLER_76_398 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_decap_8 FILLER_77_28 ();
 sg13g2_decap_8 FILLER_77_35 ();
 sg13g2_decap_8 FILLER_77_42 ();
 sg13g2_decap_8 FILLER_77_49 ();
 sg13g2_decap_8 FILLER_77_56 ();
 sg13g2_decap_8 FILLER_77_63 ();
 sg13g2_decap_8 FILLER_77_70 ();
 sg13g2_decap_8 FILLER_77_77 ();
 sg13g2_decap_8 FILLER_77_84 ();
 sg13g2_decap_8 FILLER_77_91 ();
 sg13g2_fill_2 FILLER_77_98 ();
 sg13g2_fill_1 FILLER_77_100 ();
 sg13g2_fill_1 FILLER_77_158 ();
 sg13g2_fill_1 FILLER_77_225 ();
 sg13g2_fill_2 FILLER_77_252 ();
 sg13g2_fill_1 FILLER_77_254 ();
 sg13g2_fill_1 FILLER_77_290 ();
 sg13g2_fill_2 FILLER_77_300 ();
 sg13g2_fill_2 FILLER_77_380 ();
 sg13g2_fill_1 FILLER_77_382 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_decap_8 FILLER_78_28 ();
 sg13g2_decap_8 FILLER_78_35 ();
 sg13g2_decap_8 FILLER_78_42 ();
 sg13g2_decap_8 FILLER_78_49 ();
 sg13g2_decap_8 FILLER_78_56 ();
 sg13g2_decap_8 FILLER_78_63 ();
 sg13g2_decap_8 FILLER_78_70 ();
 sg13g2_decap_8 FILLER_78_77 ();
 sg13g2_decap_8 FILLER_78_84 ();
 sg13g2_decap_8 FILLER_78_91 ();
 sg13g2_fill_1 FILLER_78_98 ();
 sg13g2_fill_2 FILLER_78_131 ();
 sg13g2_fill_1 FILLER_78_133 ();
 sg13g2_fill_2 FILLER_78_210 ();
 sg13g2_fill_2 FILLER_78_243 ();
 sg13g2_fill_1 FILLER_78_245 ();
 sg13g2_fill_2 FILLER_78_286 ();
 sg13g2_fill_1 FILLER_78_288 ();
 sg13g2_fill_2 FILLER_78_315 ();
 sg13g2_fill_1 FILLER_78_317 ();
 sg13g2_fill_2 FILLER_78_344 ();
 sg13g2_fill_2 FILLER_78_372 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_decap_8 FILLER_79_35 ();
 sg13g2_decap_8 FILLER_79_42 ();
 sg13g2_decap_8 FILLER_79_49 ();
 sg13g2_decap_8 FILLER_79_56 ();
 sg13g2_decap_8 FILLER_79_63 ();
 sg13g2_decap_8 FILLER_79_70 ();
 sg13g2_decap_8 FILLER_79_77 ();
 sg13g2_decap_4 FILLER_79_84 ();
 sg13g2_fill_1 FILLER_79_88 ();
 sg13g2_fill_1 FILLER_79_153 ();
 sg13g2_fill_1 FILLER_79_190 ();
 sg13g2_fill_2 FILLER_79_204 ();
 sg13g2_fill_1 FILLER_79_206 ();
 sg13g2_fill_1 FILLER_79_245 ();
 sg13g2_fill_2 FILLER_79_283 ();
 sg13g2_fill_2 FILLER_79_327 ();
 sg13g2_fill_2 FILLER_79_381 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_42 ();
 sg13g2_decap_8 FILLER_80_49 ();
 sg13g2_decap_8 FILLER_80_56 ();
 sg13g2_decap_8 FILLER_80_63 ();
 sg13g2_decap_8 FILLER_80_70 ();
 sg13g2_decap_4 FILLER_80_77 ();
 sg13g2_fill_1 FILLER_80_81 ();
 sg13g2_fill_1 FILLER_80_153 ();
 sg13g2_fill_1 FILLER_80_193 ();
 sg13g2_fill_2 FILLER_80_203 ();
 sg13g2_fill_2 FILLER_80_239 ();
 sg13g2_fill_2 FILLER_80_250 ();
 sg13g2_fill_2 FILLER_80_286 ();
 sg13g2_fill_2 FILLER_80_335 ();
 sg13g2_fill_1 FILLER_80_337 ();
 sg13g2_fill_2 FILLER_80_377 ();
 sg13g2_fill_2 FILLER_80_397 ();
 sg13g2_fill_1 FILLER_80_399 ();
 assign uo_out[5] = net15;
 assign uo_out[6] = net16;
 assign uo_out[7] = net17;
endmodule

module tt_um_NicklausThompson_SkyKing (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire \BNC1_out[0] ;
 wire \BNC1_out[1] ;
 wire \BNC1_out[2] ;
 wire \BNC1_out[3] ;
 wire \BNC1_out[4] ;
 wire \BNC1_out[5] ;
 wire \BNC1_out[6] ;
 wire \BNC1_out[7] ;
 wire \BNC2X_out[0] ;
 wire \BNC2X_out[1] ;
 wire \BNC2X_out[4] ;
 wire \BNC2X_out[5] ;
 wire \BNC2Y_out[0] ;
 wire \BNC2Y_out[1] ;
 wire \BNC2Y_out[4] ;
 wire \BNC2Y_out[5] ;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire \bnc_image_generator.counter[0] ;
 wire \bnc_image_generator.counter[1] ;
 wire \bnc_image_generator.counter[2] ;
 wire \bnc_image_generator.counter[4] ;
 wire hsync;
 wire \hvsync_gen.hpos[0] ;
 wire \hvsync_gen.hpos[1] ;
 wire \hvsync_gen.hpos[2] ;
 wire \hvsync_gen.hpos[3] ;
 wire \hvsync_gen.hpos[4] ;
 wire \hvsync_gen.hpos[5] ;
 wire \hvsync_gen.hpos[6] ;
 wire \hvsync_gen.hpos[7] ;
 wire \hvsync_gen.hpos[8] ;
 wire \hvsync_gen.hpos[9] ;
 wire \hvsync_gen.vpos[0] ;
 wire \hvsync_gen.vpos[1] ;
 wire \hvsync_gen.vpos[2] ;
 wire \hvsync_gen.vpos[3] ;
 wire \hvsync_gen.vpos[4] ;
 wire \hvsync_gen.vpos[5] ;
 wire \hvsync_gen.vpos[6] ;
 wire \hvsync_gen.vpos[7] ;
 wire \hvsync_gen.vpos[8] ;
 wire \hvsync_gen.vpos[9] ;
 wire \hvsync_gen.vsync ;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire clknet_0_clk;
 wire \vga_image_generator.character_hold[0] ;
 wire \vga_image_generator.character_hold[10] ;
 wire \vga_image_generator.character_hold[11] ;
 wire \vga_image_generator.character_hold[12] ;
 wire \vga_image_generator.character_hold[13] ;
 wire \vga_image_generator.character_hold[14] ;
 wire \vga_image_generator.character_hold[15] ;
 wire \vga_image_generator.character_hold[16] ;
 wire \vga_image_generator.character_hold[17] ;
 wire \vga_image_generator.character_hold[1] ;
 wire \vga_image_generator.character_hold[2] ;
 wire \vga_image_generator.character_hold[3] ;
 wire \vga_image_generator.character_hold[4] ;
 wire \vga_image_generator.character_hold[5] ;
 wire \vga_image_generator.character_hold[6] ;
 wire \vga_image_generator.character_hold[7] ;
 wire \vga_image_generator.character_hold[8] ;
 wire \vga_image_generator.character_hold[9] ;
 wire \vga_image_generator.counter[0] ;
 wire \vga_image_generator.counter[10] ;
 wire \vga_image_generator.counter[11] ;
 wire \vga_image_generator.counter[12] ;
 wire \vga_image_generator.counter[13] ;
 wire \vga_image_generator.counter[14] ;
 wire \vga_image_generator.counter[15] ;
 wire \vga_image_generator.counter[16] ;
 wire \vga_image_generator.counter[17] ;
 wire \vga_image_generator.counter[18] ;
 wire \vga_image_generator.counter[19] ;
 wire \vga_image_generator.counter[1] ;
 wire \vga_image_generator.counter[20] ;
 wire \vga_image_generator.counter[21] ;
 wire \vga_image_generator.counter[22] ;
 wire \vga_image_generator.counter[23] ;
 wire \vga_image_generator.counter[24] ;
 wire \vga_image_generator.counter[2] ;
 wire \vga_image_generator.counter[3] ;
 wire \vga_image_generator.counter[4] ;
 wire \vga_image_generator.counter[5] ;
 wire \vga_image_generator.counter[6] ;
 wire \vga_image_generator.counter[7] ;
 wire \vga_image_generator.counter[8] ;
 wire \vga_image_generator.counter[9] ;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net282;
 wire net283;
 wire net284;

 sg13g2_inv_1 _0837_ (.Y(_0096_),
    .A(net101));
 sg13g2_inv_2 _0838_ (.Y(_0097_),
    .A(\hvsync_gen.vpos[8] ));
 sg13g2_inv_1 _0839_ (.Y(_0098_),
    .A(net251));
 sg13g2_inv_1 _0840_ (.Y(_0099_),
    .A(\hvsync_gen.vpos[9] ));
 sg13g2_inv_1 _0841_ (.Y(_0100_),
    .A(net190));
 sg13g2_inv_1 _0842_ (.Y(_0101_),
    .A(net256));
 sg13g2_inv_2 _0843_ (.Y(_0102_),
    .A(net227));
 sg13g2_inv_2 _0844_ (.Y(_0103_),
    .A(net228));
 sg13g2_inv_1 _0845_ (.Y(_0104_),
    .A(\hvsync_gen.hpos[1] ));
 sg13g2_inv_1 _0846_ (.Y(_0105_),
    .A(\hvsync_gen.hpos[0] ));
 sg13g2_inv_1 _0847_ (.Y(_0106_),
    .A(net240));
 sg13g2_inv_1 _0848_ (.Y(_0107_),
    .A(net237));
 sg13g2_inv_2 _0849_ (.Y(_0108_),
    .A(net262));
 sg13g2_inv_2 _0850_ (.Y(_0109_),
    .A(net275));
 sg13g2_inv_1 _0851_ (.Y(_0110_),
    .A(_0022_));
 sg13g2_inv_1 _0852_ (.Y(_0111_),
    .A(net4));
 sg13g2_inv_1 _0853_ (.Y(_0112_),
    .A(_0018_));
 sg13g2_inv_1 _0854_ (.Y(_0113_),
    .A(net201));
 sg13g2_inv_1 _0855_ (.Y(_0114_),
    .A(net264));
 sg13g2_inv_1 _0856_ (.Y(_0115_),
    .A(net257));
 sg13g2_inv_1 _0857_ (.Y(_0116_),
    .A(net200));
 sg13g2_inv_1 _0858_ (.Y(_0117_),
    .A(net164));
 sg13g2_inv_1 _0859_ (.Y(_0118_),
    .A(net196));
 sg13g2_inv_2 _0860_ (.Y(_0119_),
    .A(net280));
 sg13g2_nor2_1 _0861_ (.A(net248),
    .B(\hvsync_gen.vpos[6] ),
    .Y(_0120_));
 sg13g2_nand2b_1 _0862_ (.Y(_0121_),
    .B(\hvsync_gen.vpos[8] ),
    .A_N(net186));
 sg13g2_nor2b_2 _0863_ (.A(net251),
    .B_N(net250),
    .Y(_0122_));
 sg13g2_nand2b_2 _0864_ (.Y(_0123_),
    .B(net250),
    .A_N(net251));
 sg13g2_nor4_2 _0865_ (.A(net248),
    .B(net249),
    .C(_0121_),
    .Y(_0124_),
    .D(_0123_));
 sg13g2_nor2_1 _0866_ (.A(\hvsync_gen.vpos[1] ),
    .B(\hvsync_gen.vpos[0] ),
    .Y(_0125_));
 sg13g2_or2_1 _0867_ (.X(_0126_),
    .B(\hvsync_gen.vpos[0] ),
    .A(\hvsync_gen.vpos[1] ));
 sg13g2_and2_1 _0868_ (.A(net254),
    .B(net256),
    .X(_0127_));
 sg13g2_nand2_1 _0869_ (.Y(_0128_),
    .A(_0126_),
    .B(_0127_));
 sg13g2_nand2_1 _0870_ (.Y(_0129_),
    .A(_0124_),
    .B(_0128_));
 sg13g2_nor3_2 _0871_ (.A(net248),
    .B(net249),
    .C(net250),
    .Y(_0130_));
 sg13g2_nor2_1 _0872_ (.A(_0097_),
    .B(_0130_),
    .Y(_0131_));
 sg13g2_o21ai_1 _0873_ (.B1(_0099_),
    .Y(_0132_),
    .A1(_0097_),
    .A2(_0130_));
 sg13g2_and2_1 _0874_ (.A(_0129_),
    .B(_0132_),
    .X(_0133_));
 sg13g2_nand3_1 _0875_ (.B(\hvsync_gen.vpos[5] ),
    .C(net252),
    .A(net248),
    .Y(_0134_));
 sg13g2_nor2_1 _0876_ (.A(\hvsync_gen.vpos[8] ),
    .B(\hvsync_gen.vpos[9] ),
    .Y(_0135_));
 sg13g2_and2_2 _0877_ (.A(net248),
    .B(net249),
    .X(_0136_));
 sg13g2_nor2b_1 _0878_ (.A(_0136_),
    .B_N(_0135_),
    .Y(_0137_));
 sg13g2_nor2b_1 _0879_ (.A(net253),
    .B_N(net255),
    .Y(_0138_));
 sg13g2_nand2b_1 _0880_ (.Y(_0139_),
    .B(net256),
    .A_N(net254));
 sg13g2_a21oi_1 _0881_ (.A1(net256),
    .A2(_0126_),
    .Y(_0140_),
    .B1(net254));
 sg13g2_nor4_1 _0882_ (.A(\hvsync_gen.vpos[8] ),
    .B(\hvsync_gen.vpos[6] ),
    .C(\hvsync_gen.vpos[9] ),
    .D(_0134_),
    .Y(_0141_));
 sg13g2_a22oi_1 _0883_ (.Y(_0142_),
    .B1(_0140_),
    .B2(_0141_),
    .A2(_0137_),
    .A1(_0134_));
 sg13g2_nor4_1 _0884_ (.A(\hvsync_gen.vpos[6] ),
    .B(_0126_),
    .C(_0134_),
    .D(_0139_),
    .Y(_0143_));
 sg13g2_nor2_2 _0885_ (.A(\hvsync_gen.hpos[7] ),
    .B(net231),
    .Y(_0144_));
 sg13g2_or2_2 _0886_ (.X(_0145_),
    .B(net231),
    .A(net228));
 sg13g2_nor2b_2 _0887_ (.A(net224),
    .B_N(\hvsync_gen.hpos[8] ),
    .Y(_0146_));
 sg13g2_nand2b_2 _0888_ (.Y(_0147_),
    .B(\hvsync_gen.hpos[8] ),
    .A_N(net224));
 sg13g2_nor2_1 _0889_ (.A(_0145_),
    .B(_0147_),
    .Y(_0148_));
 sg13g2_nor2_2 _0890_ (.A(net238),
    .B(net243),
    .Y(_0149_));
 sg13g2_or2_1 _0891_ (.X(_0150_),
    .B(net242),
    .A(net241));
 sg13g2_a21o_1 _0892_ (.A2(net242),
    .A1(net244),
    .B1(net240),
    .X(_0151_));
 sg13g2_and2_1 _0893_ (.A(net233),
    .B(net236),
    .X(_0152_));
 sg13g2_nand4_1 _0894_ (.B(_0146_),
    .C(_0151_),
    .A(_0144_),
    .Y(_0153_),
    .D(net219));
 sg13g2_nor2_2 _0895_ (.A(_0104_),
    .B(_0105_),
    .Y(_0154_));
 sg13g2_a21oi_1 _0896_ (.A1(net244),
    .A2(net204),
    .Y(_0155_),
    .B1(net242));
 sg13g2_nor2_1 _0897_ (.A(_0106_),
    .B(_0155_),
    .Y(_0156_));
 sg13g2_nor2b_1 _0898_ (.A(net234),
    .B_N(net230),
    .Y(_0157_));
 sg13g2_nand2b_2 _0899_ (.Y(_0158_),
    .B(net231),
    .A_N(net228));
 sg13g2_nor2_1 _0900_ (.A(net233),
    .B(_0158_),
    .Y(_0159_));
 sg13g2_nor2_2 _0901_ (.A(net234),
    .B(net237),
    .Y(_0160_));
 sg13g2_nor2b_1 _0902_ (.A(_0158_),
    .B_N(_0160_),
    .Y(_0161_));
 sg13g2_nand4_1 _0903_ (.B(net232),
    .C(_0146_),
    .A(_0103_),
    .Y(_0162_),
    .D(_0160_));
 sg13g2_o21ai_1 _0904_ (.B1(_0153_),
    .Y(_0163_),
    .A1(_0156_),
    .A2(_0162_));
 sg13g2_o21ai_1 _0905_ (.B1(_0163_),
    .Y(_0164_),
    .A1(_0142_),
    .A2(_0143_));
 sg13g2_nand2_1 _0906_ (.Y(_0165_),
    .A(net203),
    .B(\hvsync_gen.vpos[0] ));
 sg13g2_nor2_1 _0907_ (.A(_0139_),
    .B(_0165_),
    .Y(_0166_));
 sg13g2_or2_1 _0908_ (.X(_0167_),
    .B(_0165_),
    .A(_0139_));
 sg13g2_nor2_1 _0909_ (.A(net254),
    .B(net252),
    .Y(_0168_));
 sg13g2_nand2_1 _0910_ (.Y(_0169_),
    .A(_0120_),
    .B(_0168_));
 sg13g2_and2_1 _0911_ (.A(_0131_),
    .B(_0169_),
    .X(_0170_));
 sg13g2_a221oi_1 _0912_ (.B2(_0131_),
    .C1(\hvsync_gen.vpos[9] ),
    .B1(_0169_),
    .A1(_0124_),
    .Y(_0171_),
    .A2(_0166_));
 sg13g2_nor3_2 _0913_ (.A(\hvsync_gen.hpos[5] ),
    .B(_0147_),
    .C(_0158_),
    .Y(_0172_));
 sg13g2_and2_1 _0914_ (.A(net243),
    .B(_0154_),
    .X(_0173_));
 sg13g2_and2_2 _0915_ (.A(net240),
    .B(net242),
    .X(_0174_));
 sg13g2_and4_2 _0916_ (.A(net213),
    .B(\hvsync_gen.hpos[0] ),
    .C(net240),
    .D(net242),
    .X(_0175_));
 sg13g2_and2_1 _0917_ (.A(net236),
    .B(_0175_),
    .X(_0176_));
 sg13g2_nand2_1 _0918_ (.Y(_0177_),
    .A(net235),
    .B(_0175_));
 sg13g2_a21oi_1 _0919_ (.A1(_0172_),
    .A2(_0177_),
    .Y(_0178_),
    .B1(_0148_));
 sg13g2_nor3_2 _0920_ (.A(net228),
    .B(net231),
    .C(net233),
    .Y(_0179_));
 sg13g2_nand2b_2 _0921_ (.Y(_0180_),
    .B(_0144_),
    .A_N(\hvsync_gen.hpos[5] ));
 sg13g2_nor2b_2 _0922_ (.A(net236),
    .B_N(net233),
    .Y(_0181_));
 sg13g2_nand2b_2 _0923_ (.Y(_0182_),
    .B(net234),
    .A_N(net237));
 sg13g2_nor2_2 _0924_ (.A(_0145_),
    .B(_0182_),
    .Y(_0183_));
 sg13g2_nand4_1 _0925_ (.B(_0144_),
    .C(_0155_),
    .A(_0106_),
    .Y(_0184_),
    .D(_0181_));
 sg13g2_nor2_1 _0926_ (.A(net239),
    .B(_0182_),
    .Y(_0185_));
 sg13g2_nand2_1 _0927_ (.Y(_0186_),
    .A(_0149_),
    .B(_0181_));
 sg13g2_nor3_1 _0928_ (.A(_0104_),
    .B(\hvsync_gen.hpos[0] ),
    .C(_0150_),
    .Y(_0187_));
 sg13g2_a22oi_1 _0929_ (.Y(_0188_),
    .B1(_0187_),
    .B2(_0183_),
    .A2(_0184_),
    .A1(_0180_));
 sg13g2_or3_1 _0930_ (.A(_0171_),
    .B(_0178_),
    .C(_0188_),
    .X(_0189_));
 sg13g2_a21o_1 _0931_ (.A2(_0189_),
    .A1(_0164_),
    .B1(_0133_),
    .X(_0190_));
 sg13g2_nor3_1 _0932_ (.A(net244),
    .B(_0105_),
    .C(_0147_),
    .Y(_0191_));
 sg13g2_nor2b_2 _0933_ (.A(net240),
    .B_N(net242),
    .Y(_0192_));
 sg13g2_nand2b_1 _0934_ (.Y(_0193_),
    .B(net243),
    .A_N(net238));
 sg13g2_nor4_1 _0935_ (.A(net244),
    .B(_0105_),
    .C(_0147_),
    .D(_0193_),
    .Y(_0194_));
 sg13g2_o21ai_1 _0936_ (.B1(net226),
    .Y(_0195_),
    .A1(net229),
    .A2(net232));
 sg13g2_nor2_2 _0937_ (.A(net238),
    .B(net237),
    .Y(_0196_));
 sg13g2_nor4_1 _0938_ (.A(net233),
    .B(net235),
    .C(_0151_),
    .D(_0158_),
    .Y(_0197_));
 sg13g2_or2_1 _0939_ (.X(_0198_),
    .B(_0197_),
    .A(_0195_));
 sg13g2_a22oi_1 _0940_ (.Y(_0199_),
    .B1(_0198_),
    .B2(net223),
    .A2(_0194_),
    .A1(_0161_));
 sg13g2_nor2_2 _0941_ (.A(net226),
    .B(net224),
    .Y(_0200_));
 sg13g2_or2_1 _0942_ (.X(_0201_),
    .B(\hvsync_gen.hpos[9] ),
    .A(net226));
 sg13g2_nand2_1 _0943_ (.Y(_0202_),
    .A(net235),
    .B(_0174_));
 sg13g2_nand2_1 _0944_ (.Y(_0203_),
    .A(net219),
    .B(_0174_));
 sg13g2_a21oi_1 _0945_ (.A1(_0148_),
    .A2(_0203_),
    .Y(_0204_),
    .B1(_0200_));
 sg13g2_nor2b_2 _0946_ (.A(net242),
    .B_N(net240),
    .Y(_0205_));
 sg13g2_nand4_1 _0947_ (.B(net219),
    .C(_0154_),
    .A(_0148_),
    .Y(_0206_),
    .D(_0205_));
 sg13g2_nor2b_1 _0948_ (.A(_0204_),
    .B_N(_0206_),
    .Y(_0207_));
 sg13g2_and3_1 _0949_ (.X(_0208_),
    .A(\hvsync_gen.vpos[1] ),
    .B(\hvsync_gen.vpos[0] ),
    .C(_0127_));
 sg13g2_nor2b_2 _0950_ (.A(net249),
    .B_N(\hvsync_gen.vpos[7] ),
    .Y(_0209_));
 sg13g2_nand2b_2 _0951_ (.Y(_0210_),
    .B(net248),
    .A_N(net249));
 sg13g2_nand3_1 _0952_ (.B(_0208_),
    .C(_0209_),
    .A(_0122_),
    .Y(_0211_));
 sg13g2_and3_1 _0953_ (.X(_0212_),
    .A(_0134_),
    .B(_0137_),
    .C(_0211_));
 sg13g2_or4_1 _0954_ (.A(_0142_),
    .B(_0199_),
    .C(_0207_),
    .D(_0212_),
    .X(_0213_));
 sg13g2_nor2_2 _0955_ (.A(net244),
    .B(net204),
    .Y(_0214_));
 sg13g2_or2_2 _0956_ (.X(_0215_),
    .B(\hvsync_gen.hpos[0] ),
    .A(net244));
 sg13g2_nand2_1 _0957_ (.Y(_0216_),
    .A(_0174_),
    .B(_0215_));
 sg13g2_a21o_1 _0958_ (.A2(_0216_),
    .A1(_0183_),
    .B1(_0179_),
    .X(_0217_));
 sg13g2_nand3_1 _0959_ (.B(_0183_),
    .C(_0214_),
    .A(_0174_),
    .Y(_0218_));
 sg13g2_o21ai_1 _0960_ (.B1(_0218_),
    .Y(_0219_),
    .A1(_0200_),
    .A2(_0217_));
 sg13g2_o21ai_1 _0961_ (.B1(_0168_),
    .Y(_0220_),
    .A1(_0100_),
    .A2(_0101_));
 sg13g2_nand2_1 _0962_ (.Y(_0221_),
    .A(\hvsync_gen.vpos[5] ),
    .B(_0220_));
 sg13g2_nand4_1 _0963_ (.B(\hvsync_gen.vpos[0] ),
    .C(_0122_),
    .A(_0100_),
    .Y(_0222_),
    .D(_0138_));
 sg13g2_nand3_1 _0964_ (.B(_0221_),
    .C(_0222_),
    .A(_0120_),
    .Y(_0223_));
 sg13g2_o21ai_1 _0965_ (.B1(net235),
    .Y(_0224_),
    .A1(net240),
    .A2(net242));
 sg13g2_a21o_1 _0966_ (.A2(_0214_),
    .A1(_0192_),
    .B1(_0224_),
    .X(_0225_));
 sg13g2_a21oi_2 _0967_ (.B1(_0144_),
    .Y(_0226_),
    .A2(_0225_),
    .A1(_0159_));
 sg13g2_nor4_1 _0968_ (.A(_0121_),
    .B(_0147_),
    .C(_0170_),
    .D(_0226_),
    .Y(_0227_));
 sg13g2_nand3_1 _0969_ (.B(_0223_),
    .C(_0227_),
    .A(_0219_),
    .Y(_0228_));
 sg13g2_and2_2 _0970_ (.A(\hvsync_gen.vpos[5] ),
    .B(_0136_),
    .X(_0229_));
 sg13g2_nand2_1 _0971_ (.Y(_0230_),
    .A(net250),
    .B(_0136_));
 sg13g2_nor2_2 _0972_ (.A(net226),
    .B(net229),
    .Y(_0231_));
 sg13g2_nor2_1 _0973_ (.A(\hvsync_gen.vpos[9] ),
    .B(net2),
    .Y(_0232_));
 sg13g2_o21ai_1 _0974_ (.B1(_0232_),
    .Y(_0233_),
    .A1(net223),
    .A2(_0231_));
 sg13g2_a21oi_1 _0975_ (.A1(\hvsync_gen.vpos[8] ),
    .A2(_0229_),
    .Y(_0234_),
    .B1(_0233_));
 sg13g2_nand4_1 _0976_ (.B(_0213_),
    .C(_0228_),
    .A(_0190_),
    .Y(_0235_),
    .D(_0234_));
 sg13g2_nor2b_1 _0977_ (.A(net224),
    .B_N(_0195_),
    .Y(_0236_));
 sg13g2_a21o_1 _0978_ (.A2(_0202_),
    .A1(_0172_),
    .B1(_0236_),
    .X(_0237_));
 sg13g2_nand4_1 _0979_ (.B(_0154_),
    .C(_0172_),
    .A(net235),
    .Y(_0238_),
    .D(_0205_));
 sg13g2_nor2_1 _0980_ (.A(_0158_),
    .B(_0182_),
    .Y(_0239_));
 sg13g2_nand3_1 _0981_ (.B(_0191_),
    .C(_0239_),
    .A(_0149_),
    .Y(_0240_));
 sg13g2_nor3_1 _0982_ (.A(net228),
    .B(net244),
    .C(net243),
    .Y(_0241_));
 sg13g2_nand2_2 _0983_ (.Y(_0242_),
    .A(net231),
    .B(net234));
 sg13g2_a221oi_1 _0984_ (.B2(_0103_),
    .C1(_0102_),
    .B1(_0242_),
    .A1(_0196_),
    .Y(_0243_),
    .A2(_0241_));
 sg13g2_nand2b_1 _0985_ (.Y(_0244_),
    .B(net223),
    .A_N(_0243_));
 sg13g2_a22oi_1 _0986_ (.Y(_0245_),
    .B1(_0240_),
    .B2(_0244_),
    .A2(_0238_),
    .A1(_0237_));
 sg13g2_and2_1 _0987_ (.A(net226),
    .B(net233),
    .X(_0246_));
 sg13g2_o21ai_1 _0988_ (.B1(_0246_),
    .Y(_0247_),
    .A1(net235),
    .A2(_0151_));
 sg13g2_and2_1 _0989_ (.A(net223),
    .B(_0195_),
    .X(_0248_));
 sg13g2_a22oi_1 _0990_ (.Y(_0249_),
    .B1(_0247_),
    .B2(_0248_),
    .A2(_0194_),
    .A1(_0183_));
 sg13g2_nor3_1 _0991_ (.A(net224),
    .B(_0176_),
    .C(_0180_),
    .Y(_0250_));
 sg13g2_nor3_1 _0992_ (.A(_0200_),
    .B(_0249_),
    .C(_0250_),
    .Y(_0251_));
 sg13g2_nand2_1 _0993_ (.Y(_0252_),
    .A(net252),
    .B(_0136_));
 sg13g2_nor2_1 _0994_ (.A(net250),
    .B(_0252_),
    .Y(_0253_));
 sg13g2_nor3_1 _0995_ (.A(net254),
    .B(\hvsync_gen.vpos[1] ),
    .C(net255),
    .Y(_0254_));
 sg13g2_a22oi_1 _0996_ (.Y(_0255_),
    .B1(_0253_),
    .B2(_0254_),
    .A2(_0252_),
    .A1(_0230_));
 sg13g2_o21ai_1 _0997_ (.B1(_0255_),
    .Y(_0256_),
    .A1(_0245_),
    .A2(_0251_));
 sg13g2_nand3_1 _0998_ (.B(_0105_),
    .C(_0174_),
    .A(net244),
    .Y(_0257_));
 sg13g2_nand2b_1 _0999_ (.Y(_0258_),
    .B(_0160_),
    .A_N(net232));
 sg13g2_nor3_1 _1000_ (.A(net236),
    .B(_0175_),
    .C(_0180_),
    .Y(_0259_));
 sg13g2_o21ai_1 _1001_ (.B1(_0257_),
    .Y(_0260_),
    .A1(_0200_),
    .A2(_0259_));
 sg13g2_and3_2 _1002_ (.X(_0261_),
    .A(net231),
    .B(net233),
    .C(net236));
 sg13g2_o21ai_1 _1003_ (.B1(_0261_),
    .Y(_0262_),
    .A1(_0150_),
    .A2(_0154_));
 sg13g2_and3_1 _1004_ (.X(_0263_),
    .A(net252),
    .B(_0140_),
    .C(_0262_));
 sg13g2_nor3_1 _1005_ (.A(net235),
    .B(_0150_),
    .C(_0180_),
    .Y(_0264_));
 sg13g2_nand4_1 _1006_ (.B(_0179_),
    .C(_0192_),
    .A(_0107_),
    .Y(_0265_),
    .D(_0214_));
 sg13g2_o21ai_1 _1007_ (.B1(_0265_),
    .Y(_0266_),
    .A1(_0200_),
    .A2(_0264_));
 sg13g2_nor2_1 _1008_ (.A(_0202_),
    .B(_0242_),
    .Y(_0267_));
 sg13g2_nor3_1 _1009_ (.A(net254),
    .B(net256),
    .C(_0126_),
    .Y(_0268_));
 sg13g2_o21ai_1 _1010_ (.B1(_0220_),
    .Y(_0269_),
    .A1(_0098_),
    .A2(_0268_));
 sg13g2_a21oi_1 _1011_ (.A1(_0215_),
    .A2(_0267_),
    .Y(_0270_),
    .B1(_0269_));
 sg13g2_a22oi_1 _1012_ (.Y(_0271_),
    .B1(_0266_),
    .B2(_0270_),
    .A2(_0263_),
    .A1(_0260_));
 sg13g2_nand3_1 _1013_ (.B(_0146_),
    .C(_0229_),
    .A(_0103_),
    .Y(_0272_));
 sg13g2_o21ai_1 _1014_ (.B1(_0256_),
    .Y(_0273_),
    .A1(_0271_),
    .A2(_0272_));
 sg13g2_o21ai_1 _1015_ (.B1(net241),
    .Y(_0274_),
    .A1(net243),
    .A2(_0215_));
 sg13g2_a22oi_1 _1016_ (.Y(_0275_),
    .B1(_0274_),
    .B2(_0239_),
    .A2(_0242_),
    .A1(_0103_));
 sg13g2_nor2b_1 _1017_ (.A(net234),
    .B_N(net237),
    .Y(_0276_));
 sg13g2_and2_2 _1018_ (.A(_0192_),
    .B(_0276_),
    .X(_0277_));
 sg13g2_nor2_1 _1019_ (.A(_0158_),
    .B(_0215_),
    .Y(_0278_));
 sg13g2_a22oi_1 _1020_ (.Y(_0279_),
    .B1(_0277_),
    .B2(_0278_),
    .A2(_0226_),
    .A1(_0201_));
 sg13g2_a21oi_1 _1021_ (.A1(net241),
    .A2(net235),
    .Y(_0280_),
    .B1(_0180_));
 sg13g2_nand4_1 _1022_ (.B(_0179_),
    .C(_0205_),
    .A(net236),
    .Y(_0281_),
    .D(_0214_));
 sg13g2_o21ai_1 _1023_ (.B1(_0281_),
    .Y(_0282_),
    .A1(_0200_),
    .A2(_0280_));
 sg13g2_nand2_1 _1024_ (.Y(_0283_),
    .A(_0217_),
    .B(_0282_));
 sg13g2_o21ai_1 _1025_ (.B1(_0283_),
    .Y(_0284_),
    .A1(_0275_),
    .A2(_0279_));
 sg13g2_nand3_1 _1026_ (.B(net252),
    .C(_0136_),
    .A(net254),
    .Y(_0285_));
 sg13g2_and3_1 _1027_ (.X(_0286_),
    .A(_0167_),
    .B(_0230_),
    .C(_0285_));
 sg13g2_nor2b_2 _1028_ (.A(net255),
    .B_N(net253),
    .Y(_0287_));
 sg13g2_a22oi_1 _1029_ (.Y(_0288_),
    .B1(_0287_),
    .B2(_0125_),
    .A2(_0285_),
    .A1(_0230_));
 sg13g2_nand2_1 _1030_ (.Y(_0289_),
    .A(_0135_),
    .B(_0253_));
 sg13g2_nor4_1 _1031_ (.A(_0147_),
    .B(_0286_),
    .C(_0288_),
    .D(_0289_),
    .Y(_0290_));
 sg13g2_a221oi_1 _1032_ (.B2(_0290_),
    .C1(_0235_),
    .B1(_0284_),
    .A1(_0135_),
    .Y(_0291_),
    .A2(_0273_));
 sg13g2_o21ai_1 _1033_ (.B1(net277),
    .Y(_0292_),
    .A1(\BNC2Y_out[0] ),
    .A2(_0109_));
 sg13g2_a21o_1 _1034_ (.A2(_0109_),
    .A1(_0108_),
    .B1(_0292_),
    .X(_0293_));
 sg13g2_nand2b_1 _1035_ (.Y(uo_out[0]),
    .B(_0293_),
    .A_N(_0291_));
 sg13g2_nand2_1 _1036_ (.Y(_0294_),
    .A(_0097_),
    .B(_0291_));
 sg13g2_nor2_1 _1037_ (.A(net275),
    .B(\BNC1_out[1] ),
    .Y(_0295_));
 sg13g2_o21ai_1 _1038_ (.B1(net277),
    .Y(_0296_),
    .A1(_0109_),
    .A2(\BNC2Y_out[1] ));
 sg13g2_or2_1 _1039_ (.X(_0297_),
    .B(_0296_),
    .A(_0295_));
 sg13g2_or3_1 _1040_ (.A(net253),
    .B(net255),
    .C(_0022_),
    .X(_0298_));
 sg13g2_nand3b_1 _1041_ (.B(net250),
    .C(\hvsync_gen.vpos[7] ),
    .Y(_0299_),
    .A_N(net249));
 sg13g2_nor2_1 _1042_ (.A(_0298_),
    .B(_0299_),
    .Y(_0300_));
 sg13g2_or2_2 _1043_ (.X(_0301_),
    .B(_0299_),
    .A(_0298_));
 sg13g2_nor3_2 _1044_ (.A(_0098_),
    .B(_0298_),
    .C(_0299_),
    .Y(_0302_));
 sg13g2_or3_1 _1045_ (.A(_0098_),
    .B(_0298_),
    .C(_0299_),
    .X(_0303_));
 sg13g2_nor3_2 _1046_ (.A(_0022_),
    .B(_0123_),
    .C(_0210_),
    .Y(_0304_));
 sg13g2_nand3_1 _1047_ (.B(_0122_),
    .C(_0209_),
    .A(_0110_),
    .Y(_0305_));
 sg13g2_nor3_1 _1048_ (.A(net253),
    .B(net255),
    .C(net225),
    .Y(_0306_));
 sg13g2_a22oi_1 _1049_ (.Y(_0307_),
    .B1(_0304_),
    .B2(_0306_),
    .A2(_0302_),
    .A1(net222));
 sg13g2_and4_1 _1050_ (.A(_0110_),
    .B(_0122_),
    .C(_0209_),
    .D(_0287_),
    .X(_0308_));
 sg13g2_nand2_1 _1051_ (.Y(_0309_),
    .A(_0287_),
    .B(_0304_));
 sg13g2_and2_1 _1052_ (.A(net222),
    .B(_0308_),
    .X(_0310_));
 sg13g2_nand2b_1 _1053_ (.Y(_0311_),
    .B(_0307_),
    .A_N(_0310_));
 sg13g2_nor2_2 _1054_ (.A(net227),
    .B(_0145_),
    .Y(_0312_));
 sg13g2_and2_1 _1055_ (.A(net218),
    .B(_0312_),
    .X(_0313_));
 sg13g2_nand2_1 _1056_ (.Y(_0314_),
    .A(_0149_),
    .B(net218));
 sg13g2_nand2_1 _1057_ (.Y(_0315_),
    .A(net222),
    .B(_0231_));
 sg13g2_nand3_1 _1058_ (.B(_0304_),
    .C(_0312_),
    .A(net222),
    .Y(_0316_));
 sg13g2_o21ai_1 _1059_ (.B1(net4),
    .Y(_0317_),
    .A1(_0314_),
    .A2(_0316_));
 sg13g2_a21oi_1 _1060_ (.A1(_0311_),
    .A2(_0313_),
    .Y(_0318_),
    .B1(_0317_));
 sg13g2_nand2_2 _1061_ (.Y(_0319_),
    .A(net232),
    .B(_0231_));
 sg13g2_nand2_1 _1062_ (.Y(_0320_),
    .A(_0149_),
    .B(_0160_));
 sg13g2_nor4_1 _1063_ (.A(net225),
    .B(_0305_),
    .C(_0319_),
    .D(_0320_),
    .Y(_0321_));
 sg13g2_nand4_1 _1064_ (.B(_0018_),
    .C(_0161_),
    .A(net222),
    .Y(_0322_),
    .D(_0302_));
 sg13g2_nand2_1 _1065_ (.Y(_0323_),
    .A(_0111_),
    .B(_0322_));
 sg13g2_o21ai_1 _1066_ (.B1(\vga_image_generator.character_hold[2] ),
    .Y(_0324_),
    .A1(_0321_),
    .A2(_0323_));
 sg13g2_or2_1 _1067_ (.X(_0325_),
    .B(_0324_),
    .A(_0318_));
 sg13g2_nand2_1 _1068_ (.Y(_0326_),
    .A(net239),
    .B(_0276_));
 sg13g2_nor2b_2 _1069_ (.A(net231),
    .B_N(net238),
    .Y(_0327_));
 sg13g2_nor2b_1 _1070_ (.A(net230),
    .B_N(net234),
    .Y(_0328_));
 sg13g2_a22oi_1 _1071_ (.Y(_0329_),
    .B1(_0328_),
    .B2(_0196_),
    .A2(_0327_),
    .A1(net216));
 sg13g2_nor2_1 _1072_ (.A(_0103_),
    .B(net230),
    .Y(_0330_));
 sg13g2_nand2_1 _1073_ (.Y(_0331_),
    .A(_0112_),
    .B(_0330_));
 sg13g2_nand2_1 _1074_ (.Y(_0332_),
    .A(net217),
    .B(net216));
 sg13g2_nor2_1 _1075_ (.A(_0182_),
    .B(_0193_),
    .Y(_0333_));
 sg13g2_a22oi_1 _1076_ (.Y(_0334_),
    .B1(net217),
    .B2(net216),
    .A2(_0192_),
    .A1(_0181_));
 sg13g2_nor4_2 _1077_ (.A(net255),
    .B(_0022_),
    .C(_0123_),
    .Y(_0335_),
    .D(_0210_));
 sg13g2_nor2_1 _1078_ (.A(_0302_),
    .B(_0335_),
    .Y(_0336_));
 sg13g2_nor4_2 _1079_ (.A(_0097_),
    .B(net253),
    .C(_0123_),
    .Y(_0337_),
    .D(_0210_));
 sg13g2_and4_2 _1080_ (.A(\hvsync_gen.vpos[8] ),
    .B(net253),
    .C(_0122_),
    .D(_0209_),
    .X(_0338_));
 sg13g2_nand4_1 _1081_ (.B(net253),
    .C(_0122_),
    .A(\hvsync_gen.vpos[8] ),
    .Y(_0339_),
    .D(_0209_));
 sg13g2_a22oi_1 _1082_ (.Y(_0340_),
    .B1(_0338_),
    .B2(_0174_),
    .A2(_0337_),
    .A1(_0149_));
 sg13g2_nand2b_1 _1083_ (.Y(_0341_),
    .B(net229),
    .A_N(net227));
 sg13g2_nor2_1 _1084_ (.A(net230),
    .B(_0341_),
    .Y(_0342_));
 sg13g2_nand3_1 _1085_ (.B(net218),
    .C(_0342_),
    .A(\vga_image_generator.character_hold[6] ),
    .Y(_0343_));
 sg13g2_a21oi_1 _1086_ (.A1(_0336_),
    .A2(_0340_),
    .Y(_0344_),
    .B1(_0343_));
 sg13g2_nand2_1 _1087_ (.Y(_0345_),
    .A(net238),
    .B(_0261_));
 sg13g2_nand3_1 _1088_ (.B(_0179_),
    .C(_0196_),
    .A(net227),
    .Y(_0346_));
 sg13g2_o21ai_1 _1089_ (.B1(_0346_),
    .Y(_0347_),
    .A1(_0341_),
    .A2(_0345_));
 sg13g2_nand2_1 _1090_ (.Y(_0348_),
    .A(\vga_image_generator.character_hold[9] ),
    .B(_0347_));
 sg13g2_nand4_1 _1091_ (.B(net227),
    .C(net237),
    .A(\vga_image_generator.character_hold[10] ),
    .Y(_0349_),
    .D(_0179_));
 sg13g2_a22oi_1 _1092_ (.Y(_0350_),
    .B1(_0327_),
    .B2(net218),
    .A2(_0196_),
    .A1(_0157_));
 sg13g2_nor2b_1 _1093_ (.A(_0350_),
    .B_N(\vga_image_generator.character_hold[11] ),
    .Y(_0351_));
 sg13g2_nand3_1 _1094_ (.B(_0103_),
    .C(_0351_),
    .A(net227),
    .Y(_0352_));
 sg13g2_nand2_1 _1095_ (.Y(_0353_),
    .A(net225),
    .B(_0111_));
 sg13g2_xnor2_1 _1096_ (.Y(_0354_),
    .A(net238),
    .B(net237));
 sg13g2_nor2_2 _1097_ (.A(net234),
    .B(_0354_),
    .Y(_0355_));
 sg13g2_nand2_1 _1098_ (.Y(_0356_),
    .A(_0302_),
    .B(_0355_));
 sg13g2_a22oi_1 _1099_ (.Y(_0357_),
    .B1(_0277_),
    .B2(net4),
    .A2(net217),
    .A1(_0160_));
 sg13g2_o21ai_1 _1100_ (.B1(_0356_),
    .Y(_0358_),
    .A1(_0305_),
    .A2(_0357_));
 sg13g2_nor2b_1 _1101_ (.A(net4),
    .B_N(net222),
    .Y(_0359_));
 sg13g2_o21ai_1 _1102_ (.B1(net253),
    .Y(_0360_),
    .A1(net238),
    .A2(_0107_));
 sg13g2_nand3_1 _1103_ (.B(_0355_),
    .C(_0360_),
    .A(_0335_),
    .Y(_0361_));
 sg13g2_nand2_1 _1104_ (.Y(_0362_),
    .A(_0277_),
    .B(_0338_));
 sg13g2_nand2_1 _1105_ (.Y(_0363_),
    .A(_0361_),
    .B(_0362_));
 sg13g2_a22oi_1 _1106_ (.Y(_0364_),
    .B1(_0359_),
    .B2(_0363_),
    .A2(_0358_),
    .A1(_0353_));
 sg13g2_nand3b_1 _1107_ (.B(_0342_),
    .C(\vga_image_generator.character_hold[5] ),
    .Y(_0365_),
    .A_N(_0364_));
 sg13g2_nand2_1 _1108_ (.Y(_0366_),
    .A(_0301_),
    .B(_0305_));
 sg13g2_nand3_1 _1109_ (.B(_0160_),
    .C(net217),
    .A(\vga_image_generator.character_hold[7] ),
    .Y(_0367_));
 sg13g2_xnor2_1 _1110_ (.Y(_0368_),
    .A(net238),
    .B(net243));
 sg13g2_and2_1 _1111_ (.A(\vga_image_generator.character_hold[8] ),
    .B(_0181_),
    .X(_0369_));
 sg13g2_o21ai_1 _1112_ (.B1(_0369_),
    .Y(_0370_),
    .A1(_0335_),
    .A2(_0368_));
 sg13g2_a22oi_1 _1113_ (.Y(_0371_),
    .B1(_0367_),
    .B2(_0370_),
    .A2(_0305_),
    .A1(_0301_));
 sg13g2_nand4_1 _1114_ (.B(net218),
    .C(net217),
    .A(\vga_image_generator.character_hold[9] ),
    .Y(_0372_),
    .D(_0304_));
 sg13g2_a22oi_1 _1115_ (.Y(_0373_),
    .B1(_0355_),
    .B2(_0335_),
    .A2(_0337_),
    .A1(_0277_));
 sg13g2_nand2b_1 _1116_ (.Y(_0374_),
    .B(\vga_image_generator.character_hold[7] ),
    .A_N(_0373_));
 sg13g2_nand3b_1 _1117_ (.B(_0372_),
    .C(_0374_),
    .Y(_0375_),
    .A_N(_0371_));
 sg13g2_nand4_1 _1118_ (.B(net229),
    .C(net230),
    .A(_0102_),
    .Y(_0376_),
    .D(_0375_));
 sg13g2_a21o_1 _1119_ (.A2(_0327_),
    .A1(net216),
    .B1(net251),
    .X(_0377_));
 sg13g2_a22oi_1 _1120_ (.Y(_0378_),
    .B1(_0333_),
    .B2(_0111_),
    .A2(net216),
    .A1(net217));
 sg13g2_nor2b_1 _1121_ (.A(_0340_),
    .B_N(net222),
    .Y(_0379_));
 sg13g2_and3_1 _1122_ (.X(_0380_),
    .A(\vga_image_generator.character_hold[0] ),
    .B(_0160_),
    .C(_0312_));
 sg13g2_o21ai_1 _1123_ (.B1(_0380_),
    .Y(_0381_),
    .A1(_0311_),
    .A2(_0379_));
 sg13g2_nor4_1 _1124_ (.A(_0102_),
    .B(_0103_),
    .C(net230),
    .D(_0309_),
    .Y(_0382_));
 sg13g2_nor3_1 _1125_ (.A(_0302_),
    .B(_0338_),
    .C(_0368_),
    .Y(_0383_));
 sg13g2_nor2b_1 _1126_ (.A(_0337_),
    .B_N(_0368_),
    .Y(_0384_));
 sg13g2_nor3_1 _1127_ (.A(_0331_),
    .B(_0383_),
    .C(_0384_),
    .Y(_0385_));
 sg13g2_and2_1 _1128_ (.A(\vga_image_generator.character_hold[16] ),
    .B(net218),
    .X(_0386_));
 sg13g2_o21ai_1 _1129_ (.B1(_0386_),
    .Y(_0387_),
    .A1(_0382_),
    .A2(_0385_));
 sg13g2_and4_1 _1130_ (.A(\vga_image_generator.character_hold[17] ),
    .B(net227),
    .C(net229),
    .D(net247),
    .X(_0388_));
 sg13g2_nor2_1 _1131_ (.A(_0018_),
    .B(_0158_),
    .Y(_0389_));
 sg13g2_nand3_1 _1132_ (.B(net216),
    .C(_0389_),
    .A(\vga_image_generator.character_hold[12] ),
    .Y(_0390_));
 sg13g2_nand2_1 _1133_ (.Y(_0391_),
    .A(_0304_),
    .B(_0368_));
 sg13g2_nand3_1 _1134_ (.B(net218),
    .C(net217),
    .A(\vga_image_generator.character_hold[11] ),
    .Y(_0392_));
 sg13g2_nand3_1 _1135_ (.B(_0149_),
    .C(net216),
    .A(\vga_image_generator.character_hold[10] ),
    .Y(_0393_));
 sg13g2_and2_1 _1136_ (.A(_0392_),
    .B(_0393_),
    .X(_0394_));
 sg13g2_nor4_1 _1137_ (.A(_0018_),
    .B(_0145_),
    .C(_0305_),
    .D(_0394_),
    .Y(_0395_));
 sg13g2_nand4_1 _1138_ (.B(_0112_),
    .C(_0160_),
    .A(\vga_image_generator.character_hold[14] ),
    .Y(_0396_),
    .D(_0330_));
 sg13g2_a21oi_1 _1139_ (.A1(_0336_),
    .A2(_0391_),
    .Y(_0397_),
    .B1(_0396_));
 sg13g2_a22oi_1 _1140_ (.Y(_0398_),
    .B1(net217),
    .B2(_0181_),
    .A2(_0192_),
    .A1(net218));
 sg13g2_nor2b_1 _1141_ (.A(_0398_),
    .B_N(_0389_),
    .Y(_0399_));
 sg13g2_nor4_1 _1142_ (.A(_0102_),
    .B(net228),
    .C(_0242_),
    .D(_0354_),
    .Y(_0400_));
 sg13g2_a22oi_1 _1143_ (.Y(_0401_),
    .B1(_0400_),
    .B2(_0338_),
    .A2(_0399_),
    .A1(_0366_));
 sg13g2_nor2b_1 _1144_ (.A(_0401_),
    .B_N(\vga_image_generator.character_hold[13] ),
    .Y(_0402_));
 sg13g2_a21o_1 _1145_ (.A2(_0368_),
    .A1(net251),
    .B1(net4),
    .X(_0403_));
 sg13g2_a22oi_1 _1146_ (.Y(_0404_),
    .B1(_0403_),
    .B2(_0300_),
    .A2(_0308_),
    .A1(_0111_));
 sg13g2_nand2b_1 _1147_ (.Y(_0405_),
    .B(_0261_),
    .A_N(_0404_));
 sg13g2_nand3b_1 _1148_ (.B(_0138_),
    .C(_0261_),
    .Y(_0406_),
    .A_N(net239));
 sg13g2_nand3_1 _1149_ (.B(_0127_),
    .C(_0261_),
    .A(net239),
    .Y(_0407_));
 sg13g2_a21oi_1 _1150_ (.A1(_0406_),
    .A2(_0407_),
    .Y(_0408_),
    .B1(net4));
 sg13g2_o21ai_1 _1151_ (.B1(_0304_),
    .Y(_0409_),
    .A1(_0267_),
    .A2(_0408_));
 sg13g2_a21oi_1 _1152_ (.A1(_0405_),
    .A2(_0409_),
    .Y(_0410_),
    .B1(_0315_));
 sg13g2_nor4_1 _1153_ (.A(net225),
    .B(_0305_),
    .C(_0314_),
    .D(_0319_),
    .Y(_0411_));
 sg13g2_o21ai_1 _1154_ (.B1(\vga_image_generator.character_hold[4] ),
    .Y(_0412_),
    .A1(_0410_),
    .A2(_0411_));
 sg13g2_nand2_1 _1155_ (.Y(_0413_),
    .A(_0174_),
    .B(net216));
 sg13g2_nor3_1 _1156_ (.A(_0305_),
    .B(_0331_),
    .C(_0334_),
    .Y(_0414_));
 sg13g2_nand4_1 _1157_ (.B(net234),
    .C(_0196_),
    .A(net232),
    .Y(_0415_),
    .D(_0231_));
 sg13g2_o21ai_1 _1158_ (.B1(_0415_),
    .Y(_0416_),
    .A1(_0319_),
    .A2(_0326_));
 sg13g2_nand3_1 _1159_ (.B(net223),
    .C(_0231_),
    .A(net230),
    .Y(_0417_));
 sg13g2_a221oi_1 _1160_ (.B2(_0186_),
    .C1(_0417_),
    .B1(_0413_),
    .A1(_0303_),
    .Y(_0418_),
    .A2(_0339_));
 sg13g2_nand3_1 _1161_ (.B(_0181_),
    .C(_0192_),
    .A(net223),
    .Y(_0419_));
 sg13g2_o21ai_1 _1162_ (.B1(_0419_),
    .Y(_0420_),
    .A1(net225),
    .A2(_0332_));
 sg13g2_nor4_1 _1163_ (.A(net4),
    .B(_0307_),
    .C(_0319_),
    .D(_0326_),
    .Y(_0421_));
 sg13g2_nor2_1 _1164_ (.A(_0301_),
    .B(_0415_),
    .Y(_0422_));
 sg13g2_nor3_1 _1165_ (.A(_0305_),
    .B(_0319_),
    .C(_0334_),
    .Y(_0423_));
 sg13g2_o21ai_1 _1166_ (.B1(_0359_),
    .Y(_0424_),
    .A1(_0422_),
    .A2(_0423_));
 sg13g2_a22oi_1 _1167_ (.Y(_0425_),
    .B1(_0377_),
    .B2(_0300_),
    .A2(_0308_),
    .A1(net4));
 sg13g2_nor3_1 _1168_ (.A(_0315_),
    .B(_0329_),
    .C(_0425_),
    .Y(_0426_));
 sg13g2_nand4_1 _1169_ (.B(_0304_),
    .C(_0306_),
    .A(_0185_),
    .Y(_0427_),
    .D(_0312_));
 sg13g2_o21ai_1 _1170_ (.B1(_0427_),
    .Y(_0428_),
    .A1(_0316_),
    .A2(_0378_));
 sg13g2_o21ai_1 _1171_ (.B1(\vga_image_generator.character_hold[1] ),
    .Y(_0429_),
    .A1(_0426_),
    .A2(_0428_));
 sg13g2_nand4_1 _1172_ (.B(_0302_),
    .C(_0355_),
    .A(net230),
    .Y(_0430_),
    .D(_0388_));
 sg13g2_o21ai_1 _1173_ (.B1(_0430_),
    .Y(_0431_),
    .A1(_0309_),
    .A2(_0349_));
 sg13g2_nor4_1 _1174_ (.A(_0344_),
    .B(_0395_),
    .C(_0397_),
    .D(_0431_),
    .Y(_0432_));
 sg13g2_and2_1 _1175_ (.A(_0429_),
    .B(_0432_),
    .X(_0433_));
 sg13g2_nand4_1 _1176_ (.B(_0365_),
    .C(_0376_),
    .A(_0325_),
    .Y(_0434_),
    .D(_0433_));
 sg13g2_o21ai_1 _1177_ (.B1(_0301_),
    .Y(_0435_),
    .A1(_0390_),
    .A2(_0391_));
 sg13g2_nand4_1 _1178_ (.B(_0349_),
    .C(_0352_),
    .A(_0348_),
    .Y(_0436_),
    .D(_0390_));
 sg13g2_nor4_1 _1179_ (.A(_0102_),
    .B(_0103_),
    .C(_0301_),
    .D(_0329_),
    .Y(_0437_));
 sg13g2_or2_1 _1180_ (.X(_0438_),
    .B(_0437_),
    .A(_0414_));
 sg13g2_a221oi_1 _1181_ (.B2(\vga_image_generator.character_hold[15] ),
    .C1(_0402_),
    .B1(_0438_),
    .A1(_0435_),
    .Y(_0439_),
    .A2(_0436_));
 sg13g2_and2_1 _1182_ (.A(_0381_),
    .B(_0387_),
    .X(_0440_));
 sg13g2_nor2b_1 _1183_ (.A(_0319_),
    .B_N(_0337_),
    .Y(_0441_));
 sg13g2_a221oi_1 _1184_ (.B2(_0441_),
    .C1(_0418_),
    .B1(_0420_),
    .A1(_0310_),
    .Y(_0442_),
    .A2(_0416_));
 sg13g2_o21ai_1 _1185_ (.B1(_0424_),
    .Y(_0443_),
    .A1(_0111_),
    .A2(_0442_));
 sg13g2_o21ai_1 _1186_ (.B1(\vga_image_generator.character_hold[3] ),
    .Y(_0444_),
    .A1(_0421_),
    .A2(_0443_));
 sg13g2_nand4_1 _1187_ (.B(_0439_),
    .C(_0440_),
    .A(_0412_),
    .Y(_0445_),
    .D(_0444_));
 sg13g2_o21ai_1 _1188_ (.B1(_0291_),
    .Y(_0446_),
    .A1(_0434_),
    .A2(_0445_));
 sg13g2_nand3_1 _1189_ (.B(_0297_),
    .C(_0446_),
    .A(_0294_),
    .Y(uo_out[1]));
 sg13g2_nor2_1 _1190_ (.A(_0109_),
    .B(\BNC1_out[5] ),
    .Y(_0447_));
 sg13g2_o21ai_1 _1191_ (.B1(net277),
    .Y(_0448_),
    .A1(net275),
    .A2(\BNC1_out[2] ));
 sg13g2_o21ai_1 _1192_ (.B1(_0446_),
    .Y(uo_out[2]),
    .A1(_0447_),
    .A2(_0448_));
 sg13g2_nand2b_1 _1193_ (.Y(_0449_),
    .B(\hvsync_gen.vsync ),
    .A_N(net2));
 sg13g2_nor2_1 _1194_ (.A(net3),
    .B(\BNC1_out[3] ),
    .Y(_0450_));
 sg13g2_o21ai_1 _1195_ (.B1(net277),
    .Y(_0451_),
    .A1(_0109_),
    .A2(\BNC1_out[4] ));
 sg13g2_o21ai_1 _1196_ (.B1(_0449_),
    .Y(uo_out[3]),
    .A1(_0450_),
    .A2(_0451_));
 sg13g2_nor2_1 _1197_ (.A(net275),
    .B(\BNC1_out[4] ),
    .Y(_0452_));
 sg13g2_o21ai_1 _1198_ (.B1(net277),
    .Y(_0453_),
    .A1(_0109_),
    .A2(\BNC2Y_out[4] ));
 sg13g2_or2_1 _1199_ (.X(_0454_),
    .B(_0453_),
    .A(_0452_));
 sg13g2_nand2b_1 _1200_ (.Y(_0455_),
    .B(_0291_),
    .A_N(net248));
 sg13g2_nand4_1 _1201_ (.B(_0446_),
    .C(_0454_),
    .A(_0294_),
    .Y(uo_out[4]),
    .D(_0455_));
 sg13g2_nor2_1 _1202_ (.A(net275),
    .B(\BNC1_out[5] ),
    .Y(_0456_));
 sg13g2_o21ai_1 _1203_ (.B1(net277),
    .Y(_0457_),
    .A1(_0109_),
    .A2(\BNC2Y_out[5] ));
 sg13g2_or2_1 _1204_ (.X(_0458_),
    .B(_0457_),
    .A(_0456_));
 sg13g2_nand3_1 _1205_ (.B(_0455_),
    .C(_0458_),
    .A(_0446_),
    .Y(uo_out[5]));
 sg13g2_nor2_1 _1206_ (.A(net275),
    .B(\BNC1_out[6] ),
    .Y(_0459_));
 sg13g2_o21ai_1 _1207_ (.B1(net277),
    .Y(_0460_),
    .A1(_0109_),
    .A2(\BNC1_out[1] ));
 sg13g2_o21ai_1 _1208_ (.B1(_0446_),
    .Y(uo_out[6]),
    .A1(_0459_),
    .A2(_0460_));
 sg13g2_nor2_1 _1209_ (.A(net275),
    .B(\BNC1_out[7] ),
    .Y(_0461_));
 sg13g2_a21oi_1 _1210_ (.A1(_0108_),
    .A2(net275),
    .Y(_0462_),
    .B1(_0461_));
 sg13g2_mux2_1 _1211_ (.A0(hsync),
    .A1(_0462_),
    .S(net277),
    .X(uo_out[7]));
 sg13g2_and2_1 _1212_ (.A(net276),
    .B(\BNC2X_out[0] ),
    .X(uio_out[0]));
 sg13g2_and2_1 _1213_ (.A(net276),
    .B(\BNC2X_out[1] ),
    .X(uio_out[1]));
 sg13g2_and2_1 _1214_ (.A(net276),
    .B(\BNC1_out[7] ),
    .X(uio_out[2]));
 sg13g2_and2_1 _1215_ (.A(net276),
    .B(\BNC1_out[6] ),
    .X(uio_out[3]));
 sg13g2_and2_1 _1216_ (.A(net276),
    .B(\BNC2X_out[4] ),
    .X(uio_out[4]));
 sg13g2_and2_1 _1217_ (.A(net276),
    .B(\BNC2X_out[5] ),
    .X(uio_out[5]));
 sg13g2_and2_1 _1218_ (.A(net276),
    .B(\BNC1_out[3] ),
    .X(uio_out[6]));
 sg13g2_and2_1 _1219_ (.A(net276),
    .B(\BNC1_out[2] ),
    .X(uio_out[7]));
 sg13g2_nand2_1 _1220_ (.Y(_0463_),
    .A(net270),
    .B(_0114_));
 sg13g2_nor2_1 _1221_ (.A(_0113_),
    .B(net268),
    .Y(_0464_));
 sg13g2_nor2_2 _1222_ (.A(net268),
    .B(_0463_),
    .Y(_0465_));
 sg13g2_nand2_1 _1223_ (.Y(_0466_),
    .A(net282),
    .B(net264));
 sg13g2_nor2b_1 _1224_ (.A(_0465_),
    .B_N(_0466_),
    .Y(_0467_));
 sg13g2_inv_1 _1225_ (.Y(_0468_),
    .A(_0467_));
 sg13g2_nor2_2 _1226_ (.A(net201),
    .B(net268),
    .Y(_0469_));
 sg13g2_or2_2 _1227_ (.X(_0470_),
    .B(net268),
    .A(net270));
 sg13g2_nand3_1 _1228_ (.B(net265),
    .C(_0469_),
    .A(net263),
    .Y(_0471_));
 sg13g2_nor2_1 _1229_ (.A(_0108_),
    .B(net266),
    .Y(_0472_));
 sg13g2_a21oi_1 _1230_ (.A1(net269),
    .A2(_0472_),
    .Y(_0473_),
    .B1(net181));
 sg13g2_o21ai_1 _1231_ (.B1(_0473_),
    .Y(_0474_),
    .A1(net262),
    .A2(_0467_));
 sg13g2_inv_1 _1232_ (.Y(_0475_),
    .A(_0474_));
 sg13g2_nor2b_2 _1233_ (.A(net270),
    .B_N(net268),
    .Y(_0476_));
 sg13g2_nor2_2 _1234_ (.A(net265),
    .B(_0476_),
    .Y(_0477_));
 sg13g2_nand2_2 _1235_ (.Y(_0478_),
    .A(net269),
    .B(net265));
 sg13g2_o21ai_1 _1236_ (.B1(net257),
    .Y(_0479_),
    .A1(net263),
    .A2(_0478_));
 sg13g2_nor2_1 _1237_ (.A(_0477_),
    .B(_0479_),
    .Y(_0480_));
 sg13g2_a21oi_1 _1238_ (.A1(_0471_),
    .A2(_0475_),
    .Y(_0008_),
    .B1(_0480_));
 sg13g2_and2_2 _1239_ (.A(net270),
    .B(net268),
    .X(_0481_));
 sg13g2_nand2_2 _1240_ (.Y(_0482_),
    .A(net270),
    .B(net268));
 sg13g2_nand2_1 _1241_ (.Y(_0483_),
    .A(_0470_),
    .B(_0482_));
 sg13g2_nand3_1 _1242_ (.B(_0470_),
    .C(_0482_),
    .A(net264),
    .Y(_0484_));
 sg13g2_nor2_1 _1243_ (.A(net270),
    .B(net266),
    .Y(_0485_));
 sg13g2_nand2_1 _1244_ (.Y(_0486_),
    .A(net267),
    .B(_0483_));
 sg13g2_and2_1 _1245_ (.A(_0463_),
    .B(_0484_),
    .X(_0487_));
 sg13g2_or2_1 _1246_ (.X(_0488_),
    .B(_0487_),
    .A(net260));
 sg13g2_nor2_2 _1247_ (.A(net263),
    .B(net265),
    .Y(_0489_));
 sg13g2_mux2_1 _1248_ (.A0(net261),
    .A1(_0489_),
    .S(_0487_),
    .X(_0490_));
 sg13g2_inv_1 _1249_ (.Y(_0491_),
    .A(_0490_));
 sg13g2_nand2_1 _1250_ (.Y(_0492_),
    .A(_0113_),
    .B(_0478_));
 sg13g2_a21oi_1 _1251_ (.A1(net263),
    .A2(_0492_),
    .Y(_0493_),
    .B1(_0489_));
 sg13g2_o21ai_1 _1252_ (.B1(net220),
    .Y(_0494_),
    .A1(_0481_),
    .A2(_0493_));
 sg13g2_o21ai_1 _1253_ (.B1(_0494_),
    .Y(_0009_),
    .A1(net220),
    .A2(_0491_));
 sg13g2_nor2_1 _1254_ (.A(net265),
    .B(_0481_),
    .Y(_0495_));
 sg13g2_nand2_1 _1255_ (.Y(_0496_),
    .A(net264),
    .B(_0027_));
 sg13g2_o21ai_1 _1256_ (.B1(_0496_),
    .Y(_0497_),
    .A1(net264),
    .A2(_0481_));
 sg13g2_nand2_1 _1257_ (.Y(_0498_),
    .A(_0472_),
    .B(_0476_));
 sg13g2_o21ai_1 _1258_ (.B1(_0498_),
    .Y(_0499_),
    .A1(net262),
    .A2(_0497_));
 sg13g2_o21ai_1 _1259_ (.B1(net270),
    .Y(_0500_),
    .A1(net269),
    .A2(net266));
 sg13g2_or2_1 _1260_ (.X(_0501_),
    .B(_0500_),
    .A(net261));
 sg13g2_a22oi_1 _1261_ (.Y(_0010_),
    .B1(_0501_),
    .B2(_0473_),
    .A2(_0499_),
    .A1(net257));
 sg13g2_o21ai_1 _1262_ (.B1(net261),
    .Y(_0502_),
    .A1(net266),
    .A2(_0469_));
 sg13g2_o21ai_1 _1263_ (.B1(_0502_),
    .Y(_0503_),
    .A1(net261),
    .A2(_0467_));
 sg13g2_o21ai_1 _1264_ (.B1(_0108_),
    .Y(_0504_),
    .A1(net269),
    .A2(_0485_));
 sg13g2_nand2_1 _1265_ (.Y(_0505_),
    .A(net260),
    .B(_0482_));
 sg13g2_nand2_1 _1266_ (.Y(_0506_),
    .A(_0504_),
    .B(_0505_));
 sg13g2_and2_1 _1267_ (.A(net220),
    .B(_0502_),
    .X(_0507_));
 sg13g2_a22oi_1 _1268_ (.Y(_0508_),
    .B1(_0506_),
    .B2(_0507_),
    .A2(_0503_),
    .A1(net257));
 sg13g2_inv_1 _1269_ (.Y(_0011_),
    .A(_0508_));
 sg13g2_xnor2_1 _1270_ (.Y(_0509_),
    .A(net270),
    .B(net264));
 sg13g2_a21oi_1 _1271_ (.A1(_0470_),
    .A2(_0509_),
    .Y(_0510_),
    .B1(net259));
 sg13g2_nand2_1 _1272_ (.Y(_0511_),
    .A(net259),
    .B(_0465_));
 sg13g2_nand2_1 _1273_ (.Y(_0512_),
    .A(net258),
    .B(_0511_));
 sg13g2_nor2b_1 _1274_ (.A(_0477_),
    .B_N(_0496_),
    .Y(_0513_));
 sg13g2_o21ai_1 _1275_ (.B1(_0511_),
    .Y(_0514_),
    .A1(net259),
    .A2(_0513_));
 sg13g2_nand2_1 _1276_ (.Y(_0515_),
    .A(net221),
    .B(_0514_));
 sg13g2_o21ai_1 _1277_ (.B1(_0515_),
    .Y(_0012_),
    .A1(_0510_),
    .A2(_0512_));
 sg13g2_o21ai_1 _1278_ (.B1(net261),
    .Y(_0516_),
    .A1(net266),
    .A2(_0470_));
 sg13g2_a21oi_1 _1279_ (.A1(net269),
    .A2(net265),
    .Y(_0517_),
    .B1(net263));
 sg13g2_o21ai_1 _1280_ (.B1(_0517_),
    .Y(_0518_),
    .A1(net265),
    .A2(_0481_));
 sg13g2_nand2_1 _1281_ (.Y(_0519_),
    .A(_0516_),
    .B(_0518_));
 sg13g2_o21ai_1 _1282_ (.B1(_0466_),
    .Y(_0520_),
    .A1(net264),
    .A2(_0482_));
 sg13g2_a21oi_1 _1283_ (.A1(_0108_),
    .A2(_0520_),
    .Y(_0521_),
    .B1(net220));
 sg13g2_a22oi_1 _1284_ (.Y(_0013_),
    .B1(_0521_),
    .B2(_0516_),
    .A2(_0519_),
    .A1(net220));
 sg13g2_a21oi_1 _1285_ (.A1(net119),
    .A2(_0478_),
    .Y(_0522_),
    .B1(net257));
 sg13g2_a21oi_1 _1286_ (.A1(net257),
    .A2(_0517_),
    .Y(_0014_),
    .B1(_0522_));
 sg13g2_a21oi_2 _1287_ (.B1(net259),
    .Y(_0523_),
    .A2(_0470_),
    .A1(_0114_));
 sg13g2_nor3_1 _1288_ (.A(net258),
    .B(_0464_),
    .C(_0477_),
    .Y(_0524_));
 sg13g2_nand2_1 _1289_ (.Y(_0525_),
    .A(net268),
    .B(net258));
 sg13g2_o21ai_1 _1290_ (.B1(net259),
    .Y(_0526_),
    .A1(_0509_),
    .A2(_0525_));
 sg13g2_nor2_1 _1291_ (.A(_0524_),
    .B(_0526_),
    .Y(_0527_));
 sg13g2_a21oi_1 _1292_ (.A1(_0486_),
    .A2(_0523_),
    .Y(_0000_),
    .B1(_0527_));
 sg13g2_a21o_1 _1293_ (.A2(_0505_),
    .A1(_0463_),
    .B1(_0512_),
    .X(_0528_));
 sg13g2_nor2_1 _1294_ (.A(net259),
    .B(_0477_),
    .Y(_0529_));
 sg13g2_nand2_1 _1295_ (.Y(_0530_),
    .A(_0484_),
    .B(_0529_));
 sg13g2_nand2_1 _1296_ (.Y(_0531_),
    .A(net263),
    .B(_0478_));
 sg13g2_o21ai_1 _1297_ (.B1(_0530_),
    .Y(_0532_),
    .A1(_0465_),
    .A2(_0531_));
 sg13g2_o21ai_1 _1298_ (.B1(_0528_),
    .Y(_0001_),
    .A1(net258),
    .A2(_0532_));
 sg13g2_xnor2_1 _1299_ (.Y(_0533_),
    .A(net264),
    .B(_0481_));
 sg13g2_a21oi_1 _1300_ (.A1(net261),
    .A2(_0520_),
    .Y(_0534_),
    .B1(net258));
 sg13g2_o21ai_1 _1301_ (.B1(_0108_),
    .Y(_0535_),
    .A1(net175),
    .A2(_0483_));
 sg13g2_a21oi_1 _1302_ (.A1(net260),
    .A2(_0533_),
    .Y(_0536_),
    .B1(net221));
 sg13g2_a22oi_1 _1303_ (.Y(_0002_),
    .B1(_0535_),
    .B2(_0536_),
    .A2(net182),
    .A1(_0488_));
 sg13g2_nor2_1 _1304_ (.A(_0108_),
    .B(_0497_),
    .Y(_0537_));
 sg13g2_nor3_1 _1305_ (.A(net221),
    .B(_0523_),
    .C(_0537_),
    .Y(_0538_));
 sg13g2_a22oi_1 _1306_ (.Y(_0539_),
    .B1(_0500_),
    .B2(net261),
    .A2(_0489_),
    .A1(_0476_));
 sg13g2_a21o_1 _1307_ (.A2(_0539_),
    .A1(net221),
    .B1(_0538_),
    .X(_0003_));
 sg13g2_a22oi_1 _1308_ (.Y(_0540_),
    .B1(_0476_),
    .B2(_0489_),
    .A2(_0468_),
    .A1(net262));
 sg13g2_o21ai_1 _1309_ (.B1(net262),
    .Y(_0541_),
    .A1(net269),
    .A2(_0485_));
 sg13g2_nor2_1 _1310_ (.A(net258),
    .B(_0523_),
    .Y(_0542_));
 sg13g2_a22oi_1 _1311_ (.Y(_0004_),
    .B1(_0541_),
    .B2(_0542_),
    .A2(_0540_),
    .A1(net258));
 sg13g2_nand3_1 _1312_ (.B(_0470_),
    .C(_0509_),
    .A(net259),
    .Y(_0543_));
 sg13g2_mux2_1 _1313_ (.A0(_0465_),
    .A1(_0513_),
    .S(net259),
    .X(_0544_));
 sg13g2_a21oi_1 _1314_ (.A1(_0464_),
    .A2(_0489_),
    .Y(_0545_),
    .B1(net221));
 sg13g2_a22oi_1 _1315_ (.Y(_0005_),
    .B1(_0545_),
    .B2(_0543_),
    .A2(_0544_),
    .A1(net221));
 sg13g2_nand2_1 _1316_ (.Y(_0546_),
    .A(_0469_),
    .B(_0489_));
 sg13g2_o21ai_1 _1317_ (.B1(_0546_),
    .Y(_0547_),
    .A1(_0495_),
    .A2(_0531_));
 sg13g2_a221oi_1 _1318_ (.B2(net261),
    .C1(net221),
    .B1(_0520_),
    .A1(_0469_),
    .Y(_0548_),
    .A2(_0489_));
 sg13g2_a21oi_1 _1319_ (.A1(net220),
    .A2(_0547_),
    .Y(_0006_),
    .B1(_0548_));
 sg13g2_nand3_1 _1320_ (.B(net269),
    .C(net265),
    .A(net263),
    .Y(_0549_));
 sg13g2_nor3_1 _1321_ (.A(net220),
    .B(net119),
    .C(_0478_),
    .Y(_0550_));
 sg13g2_a21oi_1 _1322_ (.A1(net220),
    .A2(_0549_),
    .Y(_0551_),
    .B1(_0550_));
 sg13g2_inv_1 _1323_ (.Y(_0007_),
    .A(_0551_));
 sg13g2_nand3_1 _1324_ (.B(_0136_),
    .C(_0287_),
    .A(net190),
    .Y(_0552_));
 sg13g2_nor3_1 _1325_ (.A(_0121_),
    .B(_0123_),
    .C(_0552_),
    .Y(_0016_));
 sg13g2_nand2_1 _1326_ (.Y(_0553_),
    .A(net227),
    .B(net225));
 sg13g2_nand3_1 _1327_ (.B(net225),
    .C(_0258_),
    .A(net229),
    .Y(_0554_));
 sg13g2_nand2_1 _1328_ (.Y(_0555_),
    .A(_0102_),
    .B(net225));
 sg13g2_a21oi_1 _1329_ (.A1(net229),
    .A2(_0261_),
    .Y(_0556_),
    .B1(_0555_));
 sg13g2_nor2_1 _1330_ (.A(net222),
    .B(_0556_),
    .Y(_0557_));
 sg13g2_a21oi_1 _1331_ (.A1(_0553_),
    .A2(_0554_),
    .Y(_0015_),
    .B1(_0557_));
 sg13g2_and2_1 _1332_ (.A(net100),
    .B(net280),
    .X(_0028_));
 sg13g2_nor3_1 _1333_ (.A(net273),
    .B(_0469_),
    .C(_0481_),
    .Y(_0029_));
 sg13g2_nor2_1 _1334_ (.A(net273),
    .B(_0533_),
    .Y(_0030_));
 sg13g2_nor2_1 _1335_ (.A(net175),
    .B(_0482_),
    .Y(_0558_));
 sg13g2_o21ai_1 _1336_ (.B1(net280),
    .Y(_0559_),
    .A1(net260),
    .A2(_0558_));
 sg13g2_a21oi_1 _1337_ (.A1(net260),
    .A2(_0558_),
    .Y(_0031_),
    .B1(_0559_));
 sg13g2_nor2_1 _1338_ (.A(_0113_),
    .B(_0549_),
    .Y(_0560_));
 sg13g2_o21ai_1 _1339_ (.B1(net280),
    .Y(_0561_),
    .A1(net257),
    .A2(_0560_));
 sg13g2_a21oi_1 _1340_ (.A1(net257),
    .A2(_0560_),
    .Y(_0032_),
    .B1(_0561_));
 sg13g2_nand4_1 _1341_ (.B(net224),
    .C(_0176_),
    .A(net226),
    .Y(_0562_),
    .D(_0179_));
 sg13g2_and2_2 _1342_ (.A(net281),
    .B(_0562_),
    .X(_0563_));
 sg13g2_nand2_2 _1343_ (.Y(_0564_),
    .A(net281),
    .B(_0562_));
 sg13g2_nand2_1 _1344_ (.Y(_0565_),
    .A(\hvsync_gen.vpos[0] ),
    .B(_0563_));
 sg13g2_nand2_1 _1345_ (.Y(_0566_),
    .A(_0125_),
    .B(_0127_));
 sg13g2_nor4_1 _1346_ (.A(\hvsync_gen.vpos[8] ),
    .B(net252),
    .C(_0099_),
    .D(_0566_),
    .Y(_0567_));
 sg13g2_a21oi_1 _1347_ (.A1(_0130_),
    .A2(_0567_),
    .Y(_0568_),
    .B1(net274));
 sg13g2_nand2b_1 _1348_ (.Y(_0569_),
    .B(_0568_),
    .A_N(_0562_));
 sg13g2_o21ai_1 _1349_ (.B1(_0565_),
    .Y(_0033_),
    .A1(_0096_),
    .A2(_0569_));
 sg13g2_nand3b_1 _1350_ (.B(_0165_),
    .C(_0126_),
    .Y(_0570_),
    .A_N(_0569_));
 sg13g2_o21ai_1 _1351_ (.B1(_0570_),
    .Y(_0034_),
    .A1(_0100_),
    .A2(_0564_));
 sg13g2_nor2_1 _1352_ (.A(_0165_),
    .B(_0563_),
    .Y(_0571_));
 sg13g2_and2_1 _1353_ (.A(net255),
    .B(_0571_),
    .X(_0572_));
 sg13g2_nor2_2 _1354_ (.A(_0563_),
    .B(_0568_),
    .Y(_0573_));
 sg13g2_nor2_1 _1355_ (.A(net255),
    .B(_0571_),
    .Y(_0574_));
 sg13g2_nor3_1 _1356_ (.A(_0572_),
    .B(_0573_),
    .C(_0574_),
    .Y(_0035_));
 sg13g2_nor2_1 _1357_ (.A(net254),
    .B(_0572_),
    .Y(_0575_));
 sg13g2_and2_1 _1358_ (.A(_0208_),
    .B(_0564_),
    .X(_0576_));
 sg13g2_nor3_1 _1359_ (.A(_0573_),
    .B(_0575_),
    .C(_0576_),
    .Y(_0036_));
 sg13g2_and2_1 _1360_ (.A(net251),
    .B(_0576_),
    .X(_0577_));
 sg13g2_nor2_1 _1361_ (.A(net251),
    .B(_0576_),
    .Y(_0578_));
 sg13g2_nor3_1 _1362_ (.A(_0573_),
    .B(_0577_),
    .C(_0578_),
    .Y(_0037_));
 sg13g2_nor2_1 _1363_ (.A(net250),
    .B(_0577_),
    .Y(_0579_));
 sg13g2_and2_1 _1364_ (.A(net250),
    .B(_0577_),
    .X(_0580_));
 sg13g2_nor3_1 _1365_ (.A(_0573_),
    .B(_0579_),
    .C(_0580_),
    .Y(_0038_));
 sg13g2_xnor2_1 _1366_ (.Y(_0581_),
    .A(net249),
    .B(_0580_));
 sg13g2_nor2_1 _1367_ (.A(_0573_),
    .B(_0581_),
    .Y(_0039_));
 sg13g2_a21oi_1 _1368_ (.A1(net249),
    .A2(_0580_),
    .Y(_0582_),
    .B1(net248));
 sg13g2_nand2_1 _1369_ (.Y(_0583_),
    .A(_0229_),
    .B(_0577_));
 sg13g2_a21oi_1 _1370_ (.A1(_0229_),
    .A2(_0577_),
    .Y(_0584_),
    .B1(_0573_));
 sg13g2_nor2b_1 _1371_ (.A(net199),
    .B_N(_0584_),
    .Y(_0040_));
 sg13g2_xnor2_1 _1372_ (.Y(_0585_),
    .A(_0097_),
    .B(_0583_));
 sg13g2_nor2_1 _1373_ (.A(_0573_),
    .B(_0585_),
    .Y(_0041_));
 sg13g2_nand2_1 _1374_ (.Y(_0586_),
    .A(net186),
    .B(_0563_));
 sg13g2_nand4_1 _1375_ (.B(_0110_),
    .C(_0208_),
    .A(net251),
    .Y(_0587_),
    .D(_0229_));
 sg13g2_xnor2_1 _1376_ (.Y(_0588_),
    .A(_0099_),
    .B(_0587_));
 sg13g2_o21ai_1 _1377_ (.B1(_0586_),
    .Y(_0042_),
    .A1(_0569_),
    .A2(_0588_));
 sg13g2_and3_1 _1378_ (.X(_0589_),
    .A(net246),
    .B(net245),
    .C(_0118_));
 sg13g2_and2_1 _1379_ (.A(\vga_image_generator.counter[20] ),
    .B(\vga_image_generator.counter[21] ),
    .X(_0590_));
 sg13g2_a21oi_1 _1380_ (.A1(_0589_),
    .A2(_0590_),
    .Y(_0591_),
    .B1(net154));
 sg13g2_nor2_1 _1381_ (.A(net272),
    .B(_0591_),
    .Y(_0043_));
 sg13g2_nand2b_2 _1382_ (.Y(_0592_),
    .B(\vga_image_generator.counter[21] ),
    .A_N(\vga_image_generator.counter[20] ));
 sg13g2_inv_1 _1383_ (.Y(_0593_),
    .A(_0592_));
 sg13g2_a21oi_1 _1384_ (.A1(_0589_),
    .A2(_0593_),
    .Y(_0594_),
    .B1(net113));
 sg13g2_nor2_1 _1385_ (.A(net274),
    .B(net114),
    .Y(_0044_));
 sg13g2_nand2b_1 _1386_ (.Y(_0595_),
    .B(\vga_image_generator.counter[20] ),
    .A_N(\vga_image_generator.counter[21] ));
 sg13g2_inv_1 _1387_ (.Y(_0596_),
    .A(_0595_));
 sg13g2_a21oi_1 _1388_ (.A1(_0589_),
    .A2(_0596_),
    .Y(_0597_),
    .B1(net110));
 sg13g2_nor2_1 _1389_ (.A(net272),
    .B(_0597_),
    .Y(_0045_));
 sg13g2_nor2_1 _1390_ (.A(\vga_image_generator.counter[20] ),
    .B(\vga_image_generator.counter[21] ),
    .Y(_0598_));
 sg13g2_a21oi_1 _1391_ (.A1(_0589_),
    .A2(_0598_),
    .Y(_0599_),
    .B1(net117));
 sg13g2_nor2_1 _1392_ (.A(net274),
    .B(net118),
    .Y(_0046_));
 sg13g2_nor2b_2 _1393_ (.A(net246),
    .B_N(\vga_image_generator.counter[23] ),
    .Y(_0600_));
 sg13g2_and2_1 _1394_ (.A(_0118_),
    .B(_0590_),
    .X(_0601_));
 sg13g2_a21oi_1 _1395_ (.A1(_0600_),
    .A2(_0601_),
    .Y(_0602_),
    .B1(net160));
 sg13g2_nor2_1 _1396_ (.A(net272),
    .B(net161),
    .Y(_0047_));
 sg13g2_nor2_1 _1397_ (.A(\vga_image_generator.counter[24] ),
    .B(_0592_),
    .Y(_0603_));
 sg13g2_a21oi_1 _1398_ (.A1(_0600_),
    .A2(_0603_),
    .Y(_0604_),
    .B1(net158));
 sg13g2_nor2_1 _1399_ (.A(net274),
    .B(net159),
    .Y(_0048_));
 sg13g2_nor2_1 _1400_ (.A(\vga_image_generator.counter[24] ),
    .B(_0595_),
    .Y(_0605_));
 sg13g2_a21oi_1 _1401_ (.A1(_0600_),
    .A2(_0605_),
    .Y(_0606_),
    .B1(net150));
 sg13g2_nor2_1 _1402_ (.A(net272),
    .B(net151),
    .Y(_0049_));
 sg13g2_nor3_2 _1403_ (.A(\vga_image_generator.counter[20] ),
    .B(\vga_image_generator.counter[21] ),
    .C(\vga_image_generator.counter[24] ),
    .Y(_0607_));
 sg13g2_a21oi_1 _1404_ (.A1(_0600_),
    .A2(_0607_),
    .Y(_0608_),
    .B1(net121));
 sg13g2_nor2_1 _1405_ (.A(net272),
    .B(net122),
    .Y(_0050_));
 sg13g2_nor2b_2 _1406_ (.A(\vga_image_generator.counter[23] ),
    .B_N(net247),
    .Y(_0609_));
 sg13g2_a21oi_1 _1407_ (.A1(_0601_),
    .A2(_0609_),
    .Y(_0610_),
    .B1(net156));
 sg13g2_nor2_1 _1408_ (.A(net273),
    .B(net157),
    .Y(_0051_));
 sg13g2_a21oi_1 _1409_ (.A1(_0603_),
    .A2(_0609_),
    .Y(_0611_),
    .B1(net103));
 sg13g2_nor2_1 _1410_ (.A(net272),
    .B(net104),
    .Y(_0052_));
 sg13g2_a21oi_1 _1411_ (.A1(_0605_),
    .A2(_0609_),
    .Y(_0612_),
    .B1(net115));
 sg13g2_nor2_1 _1412_ (.A(net273),
    .B(net116),
    .Y(_0053_));
 sg13g2_a21oi_1 _1413_ (.A1(_0607_),
    .A2(_0609_),
    .Y(_0613_),
    .B1(net105));
 sg13g2_nor2_1 _1414_ (.A(net274),
    .B(net106),
    .Y(_0054_));
 sg13g2_nor2_1 _1415_ (.A(net246),
    .B(net245),
    .Y(_0614_));
 sg13g2_a21oi_1 _1416_ (.A1(_0601_),
    .A2(_0614_),
    .Y(_0615_),
    .B1(net155));
 sg13g2_nor2_1 _1417_ (.A(net273),
    .B(_0615_),
    .Y(_0055_));
 sg13g2_nor4_1 _1418_ (.A(net246),
    .B(net245),
    .C(\vga_image_generator.counter[24] ),
    .D(_0592_),
    .Y(_0616_));
 sg13g2_o21ai_1 _1419_ (.B1(net280),
    .Y(_0617_),
    .A1(net177),
    .A2(_0616_));
 sg13g2_inv_1 _1420_ (.Y(_0056_),
    .A(net178));
 sg13g2_nor4_1 _1421_ (.A(net246),
    .B(net245),
    .C(\vga_image_generator.counter[24] ),
    .D(_0595_),
    .Y(_0618_));
 sg13g2_o21ai_1 _1422_ (.B1(net280),
    .Y(_0619_),
    .A1(net188),
    .A2(_0618_));
 sg13g2_inv_1 _1423_ (.Y(_0057_),
    .A(net189));
 sg13g2_a21oi_1 _1424_ (.A1(_0607_),
    .A2(_0614_),
    .Y(_0620_),
    .B1(net111));
 sg13g2_nor2_1 _1425_ (.A(net273),
    .B(net112),
    .Y(_0058_));
 sg13g2_and2_1 _1426_ (.A(net1),
    .B(net99),
    .X(_0059_));
 sg13g2_o21ai_1 _1427_ (.B1(net281),
    .Y(_0621_),
    .A1(net162),
    .A2(\vga_image_generator.counter[0] ));
 sg13g2_a21oi_1 _1428_ (.A1(net162),
    .A2(\vga_image_generator.counter[0] ),
    .Y(_0060_),
    .B1(_0621_));
 sg13g2_a21oi_1 _1429_ (.A1(\vga_image_generator.counter[1] ),
    .A2(\vga_image_generator.counter[0] ),
    .Y(_0622_),
    .B1(net144));
 sg13g2_nand3_1 _1430_ (.B(\vga_image_generator.counter[0] ),
    .C(net144),
    .A(\vga_image_generator.counter[1] ),
    .Y(_0623_));
 sg13g2_nand2_1 _1431_ (.Y(_0624_),
    .A(net281),
    .B(_0623_));
 sg13g2_nor2_1 _1432_ (.A(net145),
    .B(_0624_),
    .Y(_0061_));
 sg13g2_nor2b_1 _1433_ (.A(net147),
    .B_N(_0623_),
    .Y(_0625_));
 sg13g2_and4_2 _1434_ (.A(net162),
    .B(\vga_image_generator.counter[0] ),
    .C(net144),
    .D(net147),
    .X(_0626_));
 sg13g2_nor3_1 _1435_ (.A(_0119_),
    .B(net148),
    .C(_0626_),
    .Y(_0062_));
 sg13g2_and2_1 _1436_ (.A(net179),
    .B(_0626_),
    .X(_0627_));
 sg13g2_o21ai_1 _1437_ (.B1(net279),
    .Y(_0628_),
    .A1(net179),
    .A2(_0626_));
 sg13g2_nor2_1 _1438_ (.A(_0627_),
    .B(net180),
    .Y(_0063_));
 sg13g2_xnor2_1 _1439_ (.Y(_0629_),
    .A(net172),
    .B(_0627_));
 sg13g2_nor2_1 _1440_ (.A(net272),
    .B(net173),
    .Y(_0064_));
 sg13g2_a21oi_1 _1441_ (.A1(\vga_image_generator.counter[5] ),
    .A2(_0627_),
    .Y(_0630_),
    .B1(net107));
 sg13g2_nand4_1 _1442_ (.B(net172),
    .C(net107),
    .A(net179),
    .Y(_0631_),
    .D(_0626_));
 sg13g2_nand2_1 _1443_ (.Y(_0632_),
    .A(net279),
    .B(_0631_));
 sg13g2_nor2_1 _1444_ (.A(net108),
    .B(_0632_),
    .Y(_0065_));
 sg13g2_and2_1 _1445_ (.A(_0116_),
    .B(_0631_),
    .X(_0633_));
 sg13g2_nor2_1 _1446_ (.A(_0116_),
    .B(_0631_),
    .Y(_0634_));
 sg13g2_nor3_1 _1447_ (.A(net271),
    .B(_0633_),
    .C(_0634_),
    .Y(_0066_));
 sg13g2_and2_1 _1448_ (.A(net184),
    .B(_0634_),
    .X(_0635_));
 sg13g2_o21ai_1 _1449_ (.B1(net278),
    .Y(_0636_),
    .A1(net184),
    .A2(_0634_));
 sg13g2_nor2_1 _1450_ (.A(_0635_),
    .B(net185),
    .Y(_0067_));
 sg13g2_o21ai_1 _1451_ (.B1(net278),
    .Y(_0637_),
    .A1(net132),
    .A2(_0635_));
 sg13g2_a21oi_1 _1452_ (.A1(net132),
    .A2(_0635_),
    .Y(_0068_),
    .B1(_0637_));
 sg13g2_a21oi_1 _1453_ (.A1(net132),
    .A2(_0635_),
    .Y(_0638_),
    .B1(net136));
 sg13g2_nand3_1 _1454_ (.B(net132),
    .C(net136),
    .A(\vga_image_generator.counter[8] ),
    .Y(_0639_));
 sg13g2_nor3_1 _1455_ (.A(_0116_),
    .B(_0631_),
    .C(_0639_),
    .Y(_0640_));
 sg13g2_nor3_1 _1456_ (.A(net271),
    .B(net137),
    .C(_0640_),
    .Y(_0069_));
 sg13g2_nor2_1 _1457_ (.A(net164),
    .B(_0640_),
    .Y(_0641_));
 sg13g2_nor4_2 _1458_ (.A(_0116_),
    .B(_0117_),
    .C(_0631_),
    .Y(_0642_),
    .D(_0639_));
 sg13g2_nor3_1 _1459_ (.A(net271),
    .B(net165),
    .C(_0642_),
    .Y(_0070_));
 sg13g2_o21ai_1 _1460_ (.B1(net278),
    .Y(_0643_),
    .A1(net139),
    .A2(_0642_));
 sg13g2_a21oi_1 _1461_ (.A1(net139),
    .A2(_0642_),
    .Y(_0071_),
    .B1(_0643_));
 sg13g2_a21oi_1 _1462_ (.A1(\vga_image_generator.counter[12] ),
    .A2(_0642_),
    .Y(_0644_),
    .B1(net126));
 sg13g2_and3_1 _1463_ (.X(_0645_),
    .A(net139),
    .B(net126),
    .C(_0642_));
 sg13g2_nor3_1 _1464_ (.A(net271),
    .B(net127),
    .C(_0645_),
    .Y(_0072_));
 sg13g2_xnor2_1 _1465_ (.Y(_0646_),
    .A(net174),
    .B(_0645_));
 sg13g2_nor2_1 _1466_ (.A(net271),
    .B(_0646_),
    .Y(_0073_));
 sg13g2_a21oi_1 _1467_ (.A1(\vga_image_generator.counter[14] ),
    .A2(_0645_),
    .Y(_0647_),
    .B1(net141));
 sg13g2_and3_1 _1468_ (.X(_0648_),
    .A(\vga_image_generator.counter[14] ),
    .B(net141),
    .C(_0645_));
 sg13g2_nor3_1 _1469_ (.A(net271),
    .B(net142),
    .C(_0648_),
    .Y(_0074_));
 sg13g2_o21ai_1 _1470_ (.B1(net278),
    .Y(_0649_),
    .A1(net134),
    .A2(_0648_));
 sg13g2_a21oi_1 _1471_ (.A1(net134),
    .A2(_0648_),
    .Y(_0075_),
    .B1(_0649_));
 sg13g2_a21oi_1 _1472_ (.A1(\vga_image_generator.counter[16] ),
    .A2(_0648_),
    .Y(_0650_),
    .B1(net123));
 sg13g2_and2_1 _1473_ (.A(\vga_image_generator.counter[16] ),
    .B(\vga_image_generator.counter[17] ),
    .X(_0651_));
 sg13g2_and4_2 _1474_ (.A(\vga_image_generator.counter[14] ),
    .B(net141),
    .C(_0645_),
    .D(_0651_),
    .X(_0652_));
 sg13g2_nor3_1 _1475_ (.A(net271),
    .B(net124),
    .C(_0652_),
    .Y(_0076_));
 sg13g2_o21ai_1 _1476_ (.B1(net278),
    .Y(_0653_),
    .A1(net152),
    .A2(_0652_));
 sg13g2_a21oi_1 _1477_ (.A1(net152),
    .A2(_0652_),
    .Y(_0077_),
    .B1(_0653_));
 sg13g2_a21oi_1 _1478_ (.A1(\vga_image_generator.counter[18] ),
    .A2(_0652_),
    .Y(_0654_),
    .B1(net129));
 sg13g2_and3_2 _1479_ (.X(_0655_),
    .A(net152),
    .B(net129),
    .C(_0652_));
 sg13g2_nor3_1 _1480_ (.A(net271),
    .B(net130),
    .C(_0655_),
    .Y(_0078_));
 sg13g2_o21ai_1 _1481_ (.B1(net278),
    .Y(_0656_),
    .A1(net192),
    .A2(_0655_));
 sg13g2_a21oi_1 _1482_ (.A1(net192),
    .A2(_0655_),
    .Y(_0079_),
    .B1(_0656_));
 sg13g2_a21o_1 _1483_ (.A2(_0655_),
    .A1(net192),
    .B1(net206),
    .X(_0657_));
 sg13g2_nand2_1 _1484_ (.Y(_0658_),
    .A(_0590_),
    .B(_0655_));
 sg13g2_and3_1 _1485_ (.X(_0080_),
    .A(net278),
    .B(_0657_),
    .C(_0658_));
 sg13g2_nand2b_1 _1486_ (.Y(_0659_),
    .B(_0658_),
    .A_N(net246));
 sg13g2_nand3_1 _1487_ (.B(_0590_),
    .C(_0655_),
    .A(net246),
    .Y(_0660_));
 sg13g2_and3_1 _1488_ (.X(_0081_),
    .A(net279),
    .B(_0659_),
    .C(_0660_));
 sg13g2_nand2b_1 _1489_ (.Y(_0661_),
    .B(_0660_),
    .A_N(net245));
 sg13g2_nand4_1 _1490_ (.B(net245),
    .C(_0590_),
    .A(net246),
    .Y(_0662_),
    .D(_0655_));
 sg13g2_and3_1 _1491_ (.X(_0082_),
    .A(net279),
    .B(_0661_),
    .C(_0662_));
 sg13g2_o21ai_1 _1492_ (.B1(net279),
    .Y(_0663_),
    .A1(_0118_),
    .A2(_0662_));
 sg13g2_a21oi_1 _1493_ (.A1(_0118_),
    .A2(_0662_),
    .Y(_0083_),
    .B1(_0663_));
 sg13g2_nor4_1 _1494_ (.A(net247),
    .B(net245),
    .C(net167),
    .D(_0592_),
    .Y(_0664_));
 sg13g2_o21ai_1 _1495_ (.B1(net278),
    .Y(_0665_),
    .A1(net170),
    .A2(_0664_));
 sg13g2_inv_1 _1496_ (.Y(_0084_),
    .A(net171));
 sg13g2_and2_1 _1497_ (.A(net98),
    .B(_0563_),
    .X(_0085_));
 sg13g2_nor3_1 _1498_ (.A(net274),
    .B(_0154_),
    .C(_0214_),
    .Y(_0086_));
 sg13g2_nor3_1 _1499_ (.A(net274),
    .B(_0155_),
    .C(_0173_),
    .Y(_0087_));
 sg13g2_o21ai_1 _1500_ (.B1(net281),
    .Y(_0666_),
    .A1(net240),
    .A2(_0173_));
 sg13g2_nor2_1 _1501_ (.A(net214),
    .B(_0666_),
    .Y(_0088_));
 sg13g2_o21ai_1 _1502_ (.B1(net281),
    .Y(_0667_),
    .A1(net236),
    .A2(_0175_));
 sg13g2_nor2_1 _1503_ (.A(_0176_),
    .B(_0667_),
    .Y(_0089_));
 sg13g2_xnor2_1 _1504_ (.Y(_0668_),
    .A(net233),
    .B(_0176_));
 sg13g2_nor2_1 _1505_ (.A(_0564_),
    .B(_0668_),
    .Y(_0090_));
 sg13g2_a21oi_1 _1506_ (.A1(net219),
    .A2(_0175_),
    .Y(_0669_),
    .B1(net231));
 sg13g2_and2_1 _1507_ (.A(_0175_),
    .B(_0261_),
    .X(_0670_));
 sg13g2_nor3_1 _1508_ (.A(_0564_),
    .B(_0669_),
    .C(_0670_),
    .Y(_0091_));
 sg13g2_nor2_1 _1509_ (.A(net228),
    .B(_0670_),
    .Y(_0671_));
 sg13g2_and2_1 _1510_ (.A(net228),
    .B(_0670_),
    .X(_0672_));
 sg13g2_nor3_1 _1511_ (.A(_0564_),
    .B(_0671_),
    .C(_0672_),
    .Y(_0092_));
 sg13g2_o21ai_1 _1512_ (.B1(_0563_),
    .Y(_0673_),
    .A1(net226),
    .A2(_0672_));
 sg13g2_a21oi_1 _1513_ (.A1(net226),
    .A2(_0672_),
    .Y(_0093_),
    .B1(_0673_));
 sg13g2_and2_1 _1514_ (.A(_0112_),
    .B(_0672_),
    .X(_0674_));
 sg13g2_o21ai_1 _1515_ (.B1(_0563_),
    .Y(_0675_),
    .A1(net224),
    .A2(_0674_));
 sg13g2_a21oi_1 _1516_ (.A1(net224),
    .A2(_0674_),
    .Y(_0094_),
    .B1(_0675_));
 sg13g2_nor4_1 _1517_ (.A(net247),
    .B(net245),
    .C(net167),
    .D(_0595_),
    .Y(_0676_));
 sg13g2_o21ai_1 _1518_ (.B1(net281),
    .Y(_0677_),
    .A1(\vga_image_generator.character_hold[16] ),
    .A2(net168));
 sg13g2_inv_1 _1519_ (.Y(_0095_),
    .A(net169));
 sg13g2_dfrbp_1 _1520_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net10),
    .D(_0028_),
    .Q_N(_0027_),
    .Q(\bnc_image_generator.counter[0] ));
 sg13g2_dfrbp_1 _1521_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net18),
    .D(_0029_),
    .Q_N(_0026_),
    .Q(\bnc_image_generator.counter[1] ));
 sg13g2_dfrbp_1 _1522_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net17),
    .D(_0030_),
    .Q_N(_0025_),
    .Q(\bnc_image_generator.counter[2] ));
 sg13g2_dfrbp_1 _1523_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net16),
    .D(net176),
    .Q_N(_0024_),
    .Q(\BNC1_out[0] ));
 sg13g2_dfrbp_1 _1524_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net21),
    .D(_0032_),
    .Q_N(_0735_),
    .Q(\bnc_image_generator.counter[4] ));
 sg13g2_dfrbp_1 _1525_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net15),
    .D(net194),
    .Q_N(_0734_),
    .Q(hsync));
 sg13g2_dfrbp_1 _1526_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net14),
    .D(net102),
    .Q_N(_0023_),
    .Q(\hvsync_gen.vpos[0] ));
 sg13g2_dfrbp_1 _1527_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net12),
    .D(_0034_),
    .Q_N(_0733_),
    .Q(\hvsync_gen.vpos[1] ));
 sg13g2_dfrbp_1 _1528_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net9),
    .D(_0035_),
    .Q_N(_0732_),
    .Q(\hvsync_gen.vpos[2] ));
 sg13g2_dfrbp_1 _1529_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net7),
    .D(_0036_),
    .Q_N(_0731_),
    .Q(\hvsync_gen.vpos[3] ));
 sg13g2_dfrbp_1 _1530_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net5),
    .D(_0037_),
    .Q_N(_0730_),
    .Q(\hvsync_gen.vpos[4] ));
 sg13g2_dfrbp_1 _1531_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net73),
    .D(_0038_),
    .Q_N(_0729_),
    .Q(\hvsync_gen.vpos[5] ));
 sg13g2_dfrbp_1 _1532_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net71),
    .D(_0039_),
    .Q_N(_0728_),
    .Q(\hvsync_gen.vpos[6] ));
 sg13g2_dfrbp_1 _1533_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net69),
    .D(_0040_),
    .Q_N(_0727_),
    .Q(\hvsync_gen.vpos[7] ));
 sg13g2_dfrbp_1 _1534_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net67),
    .D(_0041_),
    .Q_N(_0022_),
    .Q(\hvsync_gen.vpos[8] ));
 sg13g2_dfrbp_1 _1535_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net75),
    .D(net187),
    .Q_N(_0736_),
    .Q(\hvsync_gen.vpos[9] ));
 sg13g2_dfrbp_1 _1536_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net65),
    .D(net191),
    .Q_N(_0726_),
    .Q(\hvsync_gen.vsync ));
 sg13g2_dfrbp_1 _1537_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net63),
    .D(_0043_),
    .Q_N(_0725_),
    .Q(\vga_image_generator.character_hold[15] ));
 sg13g2_dfrbp_1 _1538_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net61),
    .D(_0044_),
    .Q_N(_0724_),
    .Q(\vga_image_generator.character_hold[14] ));
 sg13g2_dfrbp_1 _1539_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net59),
    .D(_0045_),
    .Q_N(_0723_),
    .Q(\vga_image_generator.character_hold[13] ));
 sg13g2_dfrbp_1 _1540_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net57),
    .D(_0046_),
    .Q_N(_0722_),
    .Q(\vga_image_generator.character_hold[12] ));
 sg13g2_dfrbp_1 _1541_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net55),
    .D(_0047_),
    .Q_N(_0721_),
    .Q(\vga_image_generator.character_hold[11] ));
 sg13g2_dfrbp_1 _1542_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net53),
    .D(_0048_),
    .Q_N(_0720_),
    .Q(\vga_image_generator.character_hold[10] ));
 sg13g2_dfrbp_1 _1543_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net51),
    .D(_0049_),
    .Q_N(_0719_),
    .Q(\vga_image_generator.character_hold[9] ));
 sg13g2_dfrbp_1 _1544_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net49),
    .D(_0050_),
    .Q_N(_0718_),
    .Q(\vga_image_generator.character_hold[8] ));
 sg13g2_dfrbp_1 _1545_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net47),
    .D(_0051_),
    .Q_N(_0717_),
    .Q(\vga_image_generator.character_hold[7] ));
 sg13g2_dfrbp_1 _1546_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net45),
    .D(_0052_),
    .Q_N(_0716_),
    .Q(\vga_image_generator.character_hold[6] ));
 sg13g2_dfrbp_1 _1547_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net43),
    .D(_0053_),
    .Q_N(_0715_),
    .Q(\vga_image_generator.character_hold[5] ));
 sg13g2_dfrbp_1 _1548_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net41),
    .D(_0054_),
    .Q_N(_0714_),
    .Q(\vga_image_generator.character_hold[4] ));
 sg13g2_dfrbp_1 _1549_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net39),
    .D(_0055_),
    .Q_N(_0713_),
    .Q(\vga_image_generator.character_hold[3] ));
 sg13g2_dfrbp_1 _1550_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net37),
    .D(_0056_),
    .Q_N(_0712_),
    .Q(\vga_image_generator.character_hold[2] ));
 sg13g2_dfrbp_1 _1551_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net35),
    .D(_0057_),
    .Q_N(_0711_),
    .Q(\vga_image_generator.character_hold[1] ));
 sg13g2_dfrbp_1 _1552_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net33),
    .D(_0058_),
    .Q_N(_0710_),
    .Q(\vga_image_generator.character_hold[0] ));
 sg13g2_dfrbp_1 _1553_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net31),
    .D(_0059_),
    .Q_N(_0021_),
    .Q(\vga_image_generator.counter[0] ));
 sg13g2_dfrbp_1 _1554_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net30),
    .D(net163),
    .Q_N(_0709_),
    .Q(\vga_image_generator.counter[1] ));
 sg13g2_dfrbp_1 _1555_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net29),
    .D(net146),
    .Q_N(_0708_),
    .Q(\vga_image_generator.counter[2] ));
 sg13g2_dfrbp_1 _1556_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net28),
    .D(net149),
    .Q_N(_0707_),
    .Q(\vga_image_generator.counter[3] ));
 sg13g2_dfrbp_1 _1557_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net27),
    .D(_0063_),
    .Q_N(_0706_),
    .Q(\vga_image_generator.counter[4] ));
 sg13g2_dfrbp_1 _1558_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net26),
    .D(_0064_),
    .Q_N(_0705_),
    .Q(\vga_image_generator.counter[5] ));
 sg13g2_dfrbp_1 _1559_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net25),
    .D(net109),
    .Q_N(_0704_),
    .Q(\vga_image_generator.counter[6] ));
 sg13g2_dfrbp_1 _1560_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net24),
    .D(_0066_),
    .Q_N(_0703_),
    .Q(\vga_image_generator.counter[7] ));
 sg13g2_dfrbp_1 _1561_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net23),
    .D(_0067_),
    .Q_N(_0702_),
    .Q(\vga_image_generator.counter[8] ));
 sg13g2_dfrbp_1 _1562_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net22),
    .D(net133),
    .Q_N(_0701_),
    .Q(\vga_image_generator.counter[9] ));
 sg13g2_dfrbp_1 _1563_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net20),
    .D(net138),
    .Q_N(_0700_),
    .Q(\vga_image_generator.counter[10] ));
 sg13g2_dfrbp_1 _1564_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net19),
    .D(net166),
    .Q_N(_0699_),
    .Q(\vga_image_generator.counter[11] ));
 sg13g2_dfrbp_1 _1565_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net13),
    .D(net140),
    .Q_N(_0698_),
    .Q(\vga_image_generator.counter[12] ));
 sg13g2_dfrbp_1 _1566_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net11),
    .D(net128),
    .Q_N(_0697_),
    .Q(\vga_image_generator.counter[13] ));
 sg13g2_dfrbp_1 _1567_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net8),
    .D(_0073_),
    .Q_N(_0696_),
    .Q(\vga_image_generator.counter[14] ));
 sg13g2_dfrbp_1 _1568_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net6),
    .D(net143),
    .Q_N(_0695_),
    .Q(\vga_image_generator.counter[15] ));
 sg13g2_dfrbp_1 _1569_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net74),
    .D(net135),
    .Q_N(_0694_),
    .Q(\vga_image_generator.counter[16] ));
 sg13g2_dfrbp_1 _1570_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net72),
    .D(net125),
    .Q_N(_0693_),
    .Q(\vga_image_generator.counter[17] ));
 sg13g2_dfrbp_1 _1571_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net70),
    .D(net153),
    .Q_N(_0692_),
    .Q(\vga_image_generator.counter[18] ));
 sg13g2_dfrbp_1 _1572_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net68),
    .D(net131),
    .Q_N(_0691_),
    .Q(\vga_image_generator.counter[19] ));
 sg13g2_dfrbp_1 _1573_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net66),
    .D(_0079_),
    .Q_N(_0690_),
    .Q(\vga_image_generator.counter[20] ));
 sg13g2_dfrbp_1 _1574_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net64),
    .D(_0080_),
    .Q_N(_0689_),
    .Q(\vga_image_generator.counter[21] ));
 sg13g2_dfrbp_1 _1575_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net62),
    .D(_0081_),
    .Q_N(_0688_),
    .Q(\vga_image_generator.counter[22] ));
 sg13g2_dfrbp_1 _1576_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net60),
    .D(_0082_),
    .Q_N(_0687_),
    .Q(\vga_image_generator.counter[23] ));
 sg13g2_dfrbp_1 _1577_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net58),
    .D(net197),
    .Q_N(_0020_),
    .Q(\vga_image_generator.counter[24] ));
 sg13g2_dfrbp_1 _1578_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net56),
    .D(_0084_),
    .Q_N(_0686_),
    .Q(\vga_image_generator.character_hold[17] ));
 sg13g2_dfrbp_1 _1579_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net52),
    .D(_0085_),
    .Q_N(_0019_),
    .Q(\hvsync_gen.hpos[0] ));
 sg13g2_dfrbp_1 _1580_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net50),
    .D(net205),
    .Q_N(_0685_),
    .Q(\hvsync_gen.hpos[1] ));
 sg13g2_dfrbp_1 _1581_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net48),
    .D(_0087_),
    .Q_N(_0684_),
    .Q(\hvsync_gen.hpos[2] ));
 sg13g2_dfrbp_1 _1582_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net46),
    .D(_0088_),
    .Q_N(_0683_),
    .Q(\hvsync_gen.hpos[3] ));
 sg13g2_dfrbp_1 _1583_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net44),
    .D(_0089_),
    .Q_N(_0682_),
    .Q(\hvsync_gen.hpos[4] ));
 sg13g2_dfrbp_1 _1584_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net42),
    .D(_0090_),
    .Q_N(_0681_),
    .Q(\hvsync_gen.hpos[5] ));
 sg13g2_dfrbp_1 _1585_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net40),
    .D(_0091_),
    .Q_N(_0680_),
    .Q(\hvsync_gen.hpos[6] ));
 sg13g2_dfrbp_1 _1586_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net38),
    .D(_0092_),
    .Q_N(_0679_),
    .Q(\hvsync_gen.hpos[7] ));
 sg13g2_dfrbp_1 _1587_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net36),
    .D(_0093_),
    .Q_N(_0018_),
    .Q(\hvsync_gen.hpos[8] ));
 sg13g2_dfrbp_1 _1588_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net34),
    .D(_0094_),
    .Q_N(_0017_),
    .Q(\hvsync_gen.hpos[9] ));
 sg13g2_dfrbp_1 _1589_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net76),
    .D(_0095_),
    .Q_N(_0737_),
    .Q(\vga_image_generator.character_hold[16] ));
 sg13g2_dfrbp_1 _1590_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net77),
    .D(_0008_),
    .Q_N(_0738_),
    .Q(\BNC2Y_out[0] ));
 sg13g2_dfrbp_1 _1591_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net78),
    .D(_0009_),
    .Q_N(_0739_),
    .Q(\BNC2Y_out[4] ));
 sg13g2_dfrbp_1 _1592_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net79),
    .D(_0010_),
    .Q_N(_0740_),
    .Q(\BNC2Y_out[1] ));
 sg13g2_dfrbp_1 _1593_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net80),
    .D(_0011_),
    .Q_N(_0741_),
    .Q(\BNC2Y_out[5] ));
 sg13g2_dfrbp_1 _1594_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net81),
    .D(_0012_),
    .Q_N(_0742_),
    .Q(\BNC1_out[5] ));
 sg13g2_dfrbp_1 _1595_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net82),
    .D(_0013_),
    .Q_N(_0743_),
    .Q(\BNC1_out[1] ));
 sg13g2_dfrbp_1 _1596_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net83),
    .D(net120),
    .Q_N(_0744_),
    .Q(\BNC1_out[4] ));
 sg13g2_dfrbp_1 _1597_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net84),
    .D(_0000_),
    .Q_N(_0745_),
    .Q(\BNC2X_out[0] ));
 sg13g2_dfrbp_1 _1598_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net85),
    .D(_0001_),
    .Q_N(_0746_),
    .Q(\BNC2X_out[4] ));
 sg13g2_dfrbp_1 _1599_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net86),
    .D(net183),
    .Q_N(_0747_),
    .Q(\BNC2X_out[1] ));
 sg13g2_dfrbp_1 _1600_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net87),
    .D(_0003_),
    .Q_N(_0748_),
    .Q(\BNC2X_out[5] ));
 sg13g2_dfrbp_1 _1601_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net88),
    .D(_0004_),
    .Q_N(_0749_),
    .Q(\BNC1_out[7] ));
 sg13g2_dfrbp_1 _1602_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net89),
    .D(_0005_),
    .Q_N(_0750_),
    .Q(\BNC1_out[3] ));
 sg13g2_dfrbp_1 _1603_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net54),
    .D(_0006_),
    .Q_N(_0751_),
    .Q(\BNC1_out[6] ));
 sg13g2_dfrbp_1 _1604_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net32),
    .D(_0007_),
    .Q_N(_0678_),
    .Q(\BNC1_out[2] ));
 sg13g2_tiehi _1568__6 (.L_HI(net6));
 sg13g2_tiehi _1529__7 (.L_HI(net7));
 sg13g2_tiehi _1567__8 (.L_HI(net8));
 sg13g2_tiehi _1528__9 (.L_HI(net9));
 sg13g2_tiehi _1520__10 (.L_HI(net10));
 sg13g2_tiehi _1566__11 (.L_HI(net11));
 sg13g2_tiehi _1527__12 (.L_HI(net12));
 sg13g2_tiehi _1565__13 (.L_HI(net13));
 sg13g2_tiehi _1526__14 (.L_HI(net14));
 sg13g2_tiehi _1525__15 (.L_HI(net15));
 sg13g2_tiehi _1523__16 (.L_HI(net16));
 sg13g2_tiehi _1522__17 (.L_HI(net17));
 sg13g2_tiehi _1521__18 (.L_HI(net18));
 sg13g2_tiehi _1564__19 (.L_HI(net19));
 sg13g2_tiehi _1563__20 (.L_HI(net20));
 sg13g2_tiehi _1524__21 (.L_HI(net21));
 sg13g2_tiehi _1562__22 (.L_HI(net22));
 sg13g2_tiehi _1561__23 (.L_HI(net23));
 sg13g2_tiehi _1560__24 (.L_HI(net24));
 sg13g2_tiehi _1559__25 (.L_HI(net25));
 sg13g2_tiehi _1558__26 (.L_HI(net26));
 sg13g2_tiehi _1557__27 (.L_HI(net27));
 sg13g2_tiehi _1556__28 (.L_HI(net28));
 sg13g2_tiehi _1555__29 (.L_HI(net29));
 sg13g2_tiehi _1554__30 (.L_HI(net30));
 sg13g2_tiehi _1553__31 (.L_HI(net31));
 sg13g2_tiehi _1604__32 (.L_HI(net32));
 sg13g2_tiehi _1552__33 (.L_HI(net33));
 sg13g2_tiehi _1588__34 (.L_HI(net34));
 sg13g2_tiehi _1551__35 (.L_HI(net35));
 sg13g2_tiehi _1587__36 (.L_HI(net36));
 sg13g2_tiehi _1550__37 (.L_HI(net37));
 sg13g2_tiehi _1586__38 (.L_HI(net38));
 sg13g2_tiehi _1549__39 (.L_HI(net39));
 sg13g2_tiehi _1585__40 (.L_HI(net40));
 sg13g2_tiehi _1548__41 (.L_HI(net41));
 sg13g2_tiehi _1584__42 (.L_HI(net42));
 sg13g2_tiehi _1547__43 (.L_HI(net43));
 sg13g2_tiehi _1583__44 (.L_HI(net44));
 sg13g2_tiehi _1546__45 (.L_HI(net45));
 sg13g2_tiehi _1582__46 (.L_HI(net46));
 sg13g2_tiehi _1545__47 (.L_HI(net47));
 sg13g2_tiehi _1581__48 (.L_HI(net48));
 sg13g2_tiehi _1544__49 (.L_HI(net49));
 sg13g2_tiehi _1580__50 (.L_HI(net50));
 sg13g2_tiehi _1543__51 (.L_HI(net51));
 sg13g2_tiehi _1579__52 (.L_HI(net52));
 sg13g2_tiehi _1542__53 (.L_HI(net53));
 sg13g2_tiehi _1603__54 (.L_HI(net54));
 sg13g2_tiehi _1541__55 (.L_HI(net55));
 sg13g2_tiehi _1578__56 (.L_HI(net56));
 sg13g2_tiehi _1540__57 (.L_HI(net57));
 sg13g2_tiehi _1577__58 (.L_HI(net58));
 sg13g2_tiehi _1539__59 (.L_HI(net59));
 sg13g2_tiehi _1576__60 (.L_HI(net60));
 sg13g2_tiehi _1538__61 (.L_HI(net61));
 sg13g2_tiehi _1575__62 (.L_HI(net62));
 sg13g2_tiehi _1537__63 (.L_HI(net63));
 sg13g2_tiehi _1574__64 (.L_HI(net64));
 sg13g2_tiehi _1536__65 (.L_HI(net65));
 sg13g2_tiehi _1573__66 (.L_HI(net66));
 sg13g2_tiehi _1534__67 (.L_HI(net67));
 sg13g2_tiehi _1572__68 (.L_HI(net68));
 sg13g2_tiehi _1533__69 (.L_HI(net69));
 sg13g2_tiehi _1571__70 (.L_HI(net70));
 sg13g2_tiehi _1532__71 (.L_HI(net71));
 sg13g2_tiehi _1570__72 (.L_HI(net72));
 sg13g2_tiehi _1531__73 (.L_HI(net73));
 sg13g2_tiehi _1569__74 (.L_HI(net74));
 sg13g2_tiehi _1535__75 (.L_HI(net75));
 sg13g2_tiehi _1589__76 (.L_HI(net76));
 sg13g2_tiehi _1590__77 (.L_HI(net77));
 sg13g2_tiehi _1591__78 (.L_HI(net78));
 sg13g2_tiehi _1592__79 (.L_HI(net79));
 sg13g2_tiehi _1593__80 (.L_HI(net80));
 sg13g2_tiehi _1594__81 (.L_HI(net81));
 sg13g2_tiehi _1595__82 (.L_HI(net82));
 sg13g2_tiehi _1596__83 (.L_HI(net83));
 sg13g2_tiehi _1597__84 (.L_HI(net84));
 sg13g2_tiehi _1598__85 (.L_HI(net85));
 sg13g2_tiehi _1599__86 (.L_HI(net86));
 sg13g2_tiehi _1600__87 (.L_HI(net87));
 sg13g2_tiehi _1601__88 (.L_HI(net88));
 sg13g2_tiehi _1602__89 (.L_HI(net89));
 sg13g2_tiehi tt_um_NicklausThompson_SkyKing_90 (.L_HI(net90));
 sg13g2_tiehi tt_um_NicklausThompson_SkyKing_91 (.L_HI(net91));
 sg13g2_tiehi tt_um_NicklausThompson_SkyKing_92 (.L_HI(net92));
 sg13g2_tiehi tt_um_NicklausThompson_SkyKing_93 (.L_HI(net93));
 sg13g2_tiehi tt_um_NicklausThompson_SkyKing_94 (.L_HI(net94));
 sg13g2_tiehi tt_um_NicklausThompson_SkyKing_95 (.L_HI(net95));
 sg13g2_tiehi tt_um_NicklausThompson_SkyKing_96 (.L_HI(net96));
 sg13g2_tiehi tt_um_NicklausThompson_SkyKing_97 (.L_HI(net97));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_2 fanout216 (.A(_0276_),
    .X(net216));
 sg13g2_buf_2 fanout217 (.A(_0205_),
    .X(net217));
 sg13g2_buf_2 fanout218 (.A(_0152_),
    .X(net218));
 sg13g2_buf_1 fanout219 (.A(_0152_),
    .X(net219));
 sg13g2_buf_2 fanout220 (.A(net221),
    .X(net220));
 sg13g2_buf_2 fanout221 (.A(_0115_),
    .X(net221));
 sg13g2_buf_2 fanout222 (.A(net193),
    .X(net222));
 sg13g2_buf_2 fanout223 (.A(_0017_),
    .X(net223));
 sg13g2_buf_2 fanout224 (.A(net211),
    .X(net224));
 sg13g2_buf_2 fanout225 (.A(\hvsync_gen.hpos[9] ),
    .X(net225));
 sg13g2_buf_4 fanout226 (.X(net226),
    .A(net215));
 sg13g2_buf_2 fanout227 (.A(\hvsync_gen.hpos[8] ),
    .X(net227));
 sg13g2_buf_2 fanout228 (.A(net229),
    .X(net228));
 sg13g2_buf_4 fanout229 (.X(net229),
    .A(\hvsync_gen.hpos[7] ));
 sg13g2_buf_2 fanout230 (.A(net232),
    .X(net230));
 sg13g2_buf_4 fanout231 (.X(net231),
    .A(net232));
 sg13g2_buf_2 fanout232 (.A(\hvsync_gen.hpos[6] ),
    .X(net232));
 sg13g2_buf_2 fanout233 (.A(net284),
    .X(net233));
 sg13g2_buf_4 fanout234 (.X(net234),
    .A(\hvsync_gen.hpos[5] ));
 sg13g2_buf_2 fanout235 (.A(net236),
    .X(net235));
 sg13g2_buf_2 fanout236 (.A(net237),
    .X(net236));
 sg13g2_buf_2 fanout237 (.A(\hvsync_gen.hpos[4] ),
    .X(net237));
 sg13g2_buf_2 fanout238 (.A(net241),
    .X(net238));
 sg13g2_buf_1 fanout239 (.A(net241),
    .X(net239));
 sg13g2_buf_2 fanout240 (.A(net241),
    .X(net240));
 sg13g2_buf_2 fanout241 (.A(\hvsync_gen.hpos[3] ),
    .X(net241));
 sg13g2_buf_2 fanout242 (.A(net243),
    .X(net242));
 sg13g2_buf_2 fanout243 (.A(net210),
    .X(net243));
 sg13g2_buf_2 fanout244 (.A(\hvsync_gen.hpos[1] ),
    .X(net244));
 sg13g2_buf_2 fanout245 (.A(\vga_image_generator.counter[23] ),
    .X(net245));
 sg13g2_buf_2 fanout246 (.A(net247),
    .X(net246));
 sg13g2_buf_2 fanout247 (.A(\vga_image_generator.counter[22] ),
    .X(net247));
 sg13g2_buf_4 fanout248 (.X(net248),
    .A(net198));
 sg13g2_buf_4 fanout249 (.X(net249),
    .A(net212));
 sg13g2_buf_2 fanout250 (.A(net283),
    .X(net250));
 sg13g2_buf_2 fanout251 (.A(net207),
    .X(net251));
 sg13g2_buf_2 fanout252 (.A(\hvsync_gen.vpos[4] ),
    .X(net252));
 sg13g2_buf_4 fanout253 (.X(net253),
    .A(\hvsync_gen.vpos[3] ));
 sg13g2_buf_2 fanout254 (.A(net208),
    .X(net254));
 sg13g2_buf_2 fanout255 (.A(net209),
    .X(net255));
 sg13g2_buf_1 fanout256 (.A(\hvsync_gen.vpos[2] ),
    .X(net256));
 sg13g2_buf_2 fanout257 (.A(net258),
    .X(net257));
 sg13g2_buf_2 fanout258 (.A(net181),
    .X(net258));
 sg13g2_buf_2 fanout259 (.A(net260),
    .X(net259));
 sg13g2_buf_2 fanout260 (.A(\BNC1_out[0] ),
    .X(net260));
 sg13g2_buf_2 fanout261 (.A(net202),
    .X(net261));
 sg13g2_buf_2 fanout262 (.A(net263),
    .X(net262));
 sg13g2_buf_2 fanout263 (.A(net202),
    .X(net263));
 sg13g2_buf_2 fanout264 (.A(net267),
    .X(net264));
 sg13g2_buf_2 fanout265 (.A(net267),
    .X(net265));
 sg13g2_buf_1 fanout266 (.A(net267),
    .X(net266));
 sg13g2_buf_1 fanout267 (.A(net195),
    .X(net267));
 sg13g2_buf_2 fanout268 (.A(\bnc_image_generator.counter[1] ),
    .X(net268));
 sg13g2_buf_2 fanout269 (.A(\bnc_image_generator.counter[1] ),
    .X(net269));
 sg13g2_buf_2 fanout270 (.A(\bnc_image_generator.counter[0] ),
    .X(net270));
 sg13g2_buf_2 fanout271 (.A(net273),
    .X(net271));
 sg13g2_buf_2 fanout272 (.A(net273),
    .X(net272));
 sg13g2_buf_4 fanout273 (.X(net273),
    .A(net274));
 sg13g2_buf_4 fanout274 (.X(net274),
    .A(_0119_));
 sg13g2_buf_2 fanout275 (.A(net3),
    .X(net275));
 sg13g2_buf_2 fanout276 (.A(net3),
    .X(net276));
 sg13g2_buf_2 fanout277 (.A(net2),
    .X(net277));
 sg13g2_buf_4 fanout278 (.X(net278),
    .A(net280));
 sg13g2_buf_1 fanout279 (.A(net280),
    .X(net279));
 sg13g2_buf_4 fanout280 (.X(net280),
    .A(net281));
 sg13g2_buf_4 fanout281 (.X(net281),
    .A(net1));
 sg13g2_buf_2 input1 (.A(rst_n),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[0]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[1]),
    .X(net3));
 sg13g2_buf_4 input4 (.X(net4),
    .A(ui_in[3]));
 sg13g2_tiehi _1530__5 (.L_HI(net5));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_4_1_0_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_4_3_0_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_4_5_0_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_4_6_0_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_4_7_0_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_4_9_0_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_4_10_0_clk));
 sg13g2_inv_1 clkload7 (.A(clknet_4_11_0_clk));
 sg13g2_inv_1 clkload8 (.A(clknet_4_13_0_clk));
 sg13g2_inv_1 clkload9 (.A(clknet_4_14_0_clk));
 sg13g2_inv_1 clkload10 (.A(clknet_4_15_0_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(_0019_),
    .X(net98));
 sg13g2_dlygate4sd3_1 hold2 (.A(_0021_),
    .X(net99));
 sg13g2_dlygate4sd3_1 hold3 (.A(_0027_),
    .X(net100));
 sg13g2_dlygate4sd3_1 hold4 (.A(_0023_),
    .X(net101));
 sg13g2_dlygate4sd3_1 hold5 (.A(_0033_),
    .X(net102));
 sg13g2_dlygate4sd3_1 hold6 (.A(\vga_image_generator.character_hold[6] ),
    .X(net103));
 sg13g2_dlygate4sd3_1 hold7 (.A(_0611_),
    .X(net104));
 sg13g2_dlygate4sd3_1 hold8 (.A(\vga_image_generator.character_hold[4] ),
    .X(net105));
 sg13g2_dlygate4sd3_1 hold9 (.A(_0613_),
    .X(net106));
 sg13g2_dlygate4sd3_1 hold10 (.A(\vga_image_generator.counter[6] ),
    .X(net107));
 sg13g2_dlygate4sd3_1 hold11 (.A(_0630_),
    .X(net108));
 sg13g2_dlygate4sd3_1 hold12 (.A(_0065_),
    .X(net109));
 sg13g2_dlygate4sd3_1 hold13 (.A(\vga_image_generator.character_hold[13] ),
    .X(net110));
 sg13g2_dlygate4sd3_1 hold14 (.A(\vga_image_generator.character_hold[0] ),
    .X(net111));
 sg13g2_dlygate4sd3_1 hold15 (.A(_0620_),
    .X(net112));
 sg13g2_dlygate4sd3_1 hold16 (.A(\vga_image_generator.character_hold[14] ),
    .X(net113));
 sg13g2_dlygate4sd3_1 hold17 (.A(_0594_),
    .X(net114));
 sg13g2_dlygate4sd3_1 hold18 (.A(\vga_image_generator.character_hold[5] ),
    .X(net115));
 sg13g2_dlygate4sd3_1 hold19 (.A(_0612_),
    .X(net116));
 sg13g2_dlygate4sd3_1 hold20 (.A(\vga_image_generator.character_hold[12] ),
    .X(net117));
 sg13g2_dlygate4sd3_1 hold21 (.A(_0599_),
    .X(net118));
 sg13g2_dlygate4sd3_1 hold22 (.A(_0024_),
    .X(net119));
 sg13g2_dlygate4sd3_1 hold23 (.A(_0014_),
    .X(net120));
 sg13g2_dlygate4sd3_1 hold24 (.A(\vga_image_generator.character_hold[8] ),
    .X(net121));
 sg13g2_dlygate4sd3_1 hold25 (.A(_0608_),
    .X(net122));
 sg13g2_dlygate4sd3_1 hold26 (.A(\vga_image_generator.counter[17] ),
    .X(net123));
 sg13g2_dlygate4sd3_1 hold27 (.A(_0650_),
    .X(net124));
 sg13g2_dlygate4sd3_1 hold28 (.A(_0076_),
    .X(net125));
 sg13g2_dlygate4sd3_1 hold29 (.A(\vga_image_generator.counter[13] ),
    .X(net126));
 sg13g2_dlygate4sd3_1 hold30 (.A(_0644_),
    .X(net127));
 sg13g2_dlygate4sd3_1 hold31 (.A(_0072_),
    .X(net128));
 sg13g2_dlygate4sd3_1 hold32 (.A(\vga_image_generator.counter[19] ),
    .X(net129));
 sg13g2_dlygate4sd3_1 hold33 (.A(_0654_),
    .X(net130));
 sg13g2_dlygate4sd3_1 hold34 (.A(_0078_),
    .X(net131));
 sg13g2_dlygate4sd3_1 hold35 (.A(\vga_image_generator.counter[9] ),
    .X(net132));
 sg13g2_dlygate4sd3_1 hold36 (.A(_0068_),
    .X(net133));
 sg13g2_dlygate4sd3_1 hold37 (.A(\vga_image_generator.counter[16] ),
    .X(net134));
 sg13g2_dlygate4sd3_1 hold38 (.A(_0075_),
    .X(net135));
 sg13g2_dlygate4sd3_1 hold39 (.A(\vga_image_generator.counter[10] ),
    .X(net136));
 sg13g2_dlygate4sd3_1 hold40 (.A(_0638_),
    .X(net137));
 sg13g2_dlygate4sd3_1 hold41 (.A(_0069_),
    .X(net138));
 sg13g2_dlygate4sd3_1 hold42 (.A(\vga_image_generator.counter[12] ),
    .X(net139));
 sg13g2_dlygate4sd3_1 hold43 (.A(_0071_),
    .X(net140));
 sg13g2_dlygate4sd3_1 hold44 (.A(\vga_image_generator.counter[15] ),
    .X(net141));
 sg13g2_dlygate4sd3_1 hold45 (.A(_0647_),
    .X(net142));
 sg13g2_dlygate4sd3_1 hold46 (.A(_0074_),
    .X(net143));
 sg13g2_dlygate4sd3_1 hold47 (.A(\vga_image_generator.counter[2] ),
    .X(net144));
 sg13g2_dlygate4sd3_1 hold48 (.A(_0622_),
    .X(net145));
 sg13g2_dlygate4sd3_1 hold49 (.A(_0061_),
    .X(net146));
 sg13g2_dlygate4sd3_1 hold50 (.A(\vga_image_generator.counter[3] ),
    .X(net147));
 sg13g2_dlygate4sd3_1 hold51 (.A(_0625_),
    .X(net148));
 sg13g2_dlygate4sd3_1 hold52 (.A(_0062_),
    .X(net149));
 sg13g2_dlygate4sd3_1 hold53 (.A(\vga_image_generator.character_hold[9] ),
    .X(net150));
 sg13g2_dlygate4sd3_1 hold54 (.A(_0606_),
    .X(net151));
 sg13g2_dlygate4sd3_1 hold55 (.A(\vga_image_generator.counter[18] ),
    .X(net152));
 sg13g2_dlygate4sd3_1 hold56 (.A(_0077_),
    .X(net153));
 sg13g2_dlygate4sd3_1 hold57 (.A(\vga_image_generator.character_hold[15] ),
    .X(net154));
 sg13g2_dlygate4sd3_1 hold58 (.A(\vga_image_generator.character_hold[3] ),
    .X(net155));
 sg13g2_dlygate4sd3_1 hold59 (.A(\vga_image_generator.character_hold[7] ),
    .X(net156));
 sg13g2_dlygate4sd3_1 hold60 (.A(_0610_),
    .X(net157));
 sg13g2_dlygate4sd3_1 hold61 (.A(\vga_image_generator.character_hold[10] ),
    .X(net158));
 sg13g2_dlygate4sd3_1 hold62 (.A(_0604_),
    .X(net159));
 sg13g2_dlygate4sd3_1 hold63 (.A(\vga_image_generator.character_hold[11] ),
    .X(net160));
 sg13g2_dlygate4sd3_1 hold64 (.A(_0602_),
    .X(net161));
 sg13g2_dlygate4sd3_1 hold65 (.A(\vga_image_generator.counter[1] ),
    .X(net162));
 sg13g2_dlygate4sd3_1 hold66 (.A(_0060_),
    .X(net163));
 sg13g2_dlygate4sd3_1 hold67 (.A(\vga_image_generator.counter[11] ),
    .X(net164));
 sg13g2_dlygate4sd3_1 hold68 (.A(_0641_),
    .X(net165));
 sg13g2_dlygate4sd3_1 hold69 (.A(_0070_),
    .X(net166));
 sg13g2_dlygate4sd3_1 hold70 (.A(_0020_),
    .X(net167));
 sg13g2_dlygate4sd3_1 hold71 (.A(_0676_),
    .X(net168));
 sg13g2_dlygate4sd3_1 hold72 (.A(_0677_),
    .X(net169));
 sg13g2_dlygate4sd3_1 hold73 (.A(\vga_image_generator.character_hold[17] ),
    .X(net170));
 sg13g2_dlygate4sd3_1 hold74 (.A(_0665_),
    .X(net171));
 sg13g2_dlygate4sd3_1 hold75 (.A(\vga_image_generator.counter[5] ),
    .X(net172));
 sg13g2_dlygate4sd3_1 hold76 (.A(_0629_),
    .X(net173));
 sg13g2_dlygate4sd3_1 hold77 (.A(\vga_image_generator.counter[14] ),
    .X(net174));
 sg13g2_dlygate4sd3_1 hold78 (.A(_0025_),
    .X(net175));
 sg13g2_dlygate4sd3_1 hold79 (.A(_0031_),
    .X(net176));
 sg13g2_dlygate4sd3_1 hold80 (.A(\vga_image_generator.character_hold[2] ),
    .X(net177));
 sg13g2_dlygate4sd3_1 hold81 (.A(_0617_),
    .X(net178));
 sg13g2_dlygate4sd3_1 hold82 (.A(\vga_image_generator.counter[4] ),
    .X(net179));
 sg13g2_dlygate4sd3_1 hold83 (.A(_0628_),
    .X(net180));
 sg13g2_dlygate4sd3_1 hold84 (.A(\bnc_image_generator.counter[4] ),
    .X(net181));
 sg13g2_dlygate4sd3_1 hold85 (.A(_0534_),
    .X(net182));
 sg13g2_dlygate4sd3_1 hold86 (.A(_0002_),
    .X(net183));
 sg13g2_dlygate4sd3_1 hold87 (.A(\vga_image_generator.counter[8] ),
    .X(net184));
 sg13g2_dlygate4sd3_1 hold88 (.A(_0636_),
    .X(net185));
 sg13g2_dlygate4sd3_1 hold89 (.A(\hvsync_gen.vpos[9] ),
    .X(net186));
 sg13g2_dlygate4sd3_1 hold90 (.A(_0042_),
    .X(net187));
 sg13g2_dlygate4sd3_1 hold91 (.A(\vga_image_generator.character_hold[1] ),
    .X(net188));
 sg13g2_dlygate4sd3_1 hold92 (.A(_0619_),
    .X(net189));
 sg13g2_dlygate4sd3_1 hold93 (.A(\hvsync_gen.vpos[1] ),
    .X(net190));
 sg13g2_dlygate4sd3_1 hold94 (.A(_0016_),
    .X(net191));
 sg13g2_dlygate4sd3_1 hold95 (.A(\vga_image_generator.counter[20] ),
    .X(net192));
 sg13g2_dlygate4sd3_1 hold96 (.A(_0017_),
    .X(net193));
 sg13g2_dlygate4sd3_1 hold97 (.A(_0015_),
    .X(net194));
 sg13g2_dlygate4sd3_1 hold98 (.A(\bnc_image_generator.counter[2] ),
    .X(net195));
 sg13g2_dlygate4sd3_1 hold99 (.A(\vga_image_generator.counter[24] ),
    .X(net196));
 sg13g2_dlygate4sd3_1 hold100 (.A(_0083_),
    .X(net197));
 sg13g2_dlygate4sd3_1 hold101 (.A(\hvsync_gen.vpos[7] ),
    .X(net198));
 sg13g2_dlygate4sd3_1 hold102 (.A(_0582_),
    .X(net199));
 sg13g2_dlygate4sd3_1 hold103 (.A(\vga_image_generator.counter[7] ),
    .X(net200));
 sg13g2_dlygate4sd3_1 hold104 (.A(\bnc_image_generator.counter[0] ),
    .X(net201));
 sg13g2_dlygate4sd3_1 hold105 (.A(\BNC1_out[0] ),
    .X(net202));
 sg13g2_dlygate4sd3_1 hold106 (.A(\hvsync_gen.vpos[1] ),
    .X(net203));
 sg13g2_dlygate4sd3_1 hold107 (.A(\hvsync_gen.hpos[0] ),
    .X(net204));
 sg13g2_dlygate4sd3_1 hold108 (.A(_0086_),
    .X(net205));
 sg13g2_dlygate4sd3_1 hold109 (.A(\vga_image_generator.counter[21] ),
    .X(net206));
 sg13g2_dlygate4sd3_1 hold110 (.A(\hvsync_gen.vpos[4] ),
    .X(net207));
 sg13g2_dlygate4sd3_1 hold111 (.A(\hvsync_gen.vpos[3] ),
    .X(net208));
 sg13g2_dlygate4sd3_1 hold112 (.A(\hvsync_gen.vpos[2] ),
    .X(net209));
 sg13g2_dlygate4sd3_1 hold113 (.A(\hvsync_gen.hpos[2] ),
    .X(net210));
 sg13g2_dlygate4sd3_1 hold114 (.A(\hvsync_gen.hpos[9] ),
    .X(net211));
 sg13g2_dlygate4sd3_1 hold115 (.A(\hvsync_gen.vpos[6] ),
    .X(net212));
 sg13g2_dlygate4sd3_1 hold116 (.A(\hvsync_gen.hpos[1] ),
    .X(net213));
 sg13g2_dlygate4sd3_1 hold117 (.A(_0175_),
    .X(net214));
 sg13g2_dlygate4sd3_1 hold118 (.A(\hvsync_gen.hpos[8] ),
    .X(net215));
 sg13g2_dlygate4sd3_1 hold119 (.A(_0026_),
    .X(net282));
 sg13g2_dlygate4sd3_1 hold120 (.A(\hvsync_gen.vpos[5] ),
    .X(net283));
 sg13g2_dlygate4sd3_1 hold121 (.A(\hvsync_gen.hpos[5] ),
    .X(net284));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_fill_1 FILLER_6_84 ();
 sg13g2_fill_2 FILLER_6_89 ();
 sg13g2_decap_8 FILLER_6_95 ();
 sg13g2_decap_8 FILLER_6_102 ();
 sg13g2_decap_8 FILLER_6_109 ();
 sg13g2_decap_8 FILLER_6_116 ();
 sg13g2_decap_8 FILLER_6_123 ();
 sg13g2_decap_8 FILLER_6_130 ();
 sg13g2_decap_8 FILLER_6_137 ();
 sg13g2_decap_8 FILLER_6_144 ();
 sg13g2_decap_8 FILLER_6_151 ();
 sg13g2_decap_8 FILLER_6_158 ();
 sg13g2_decap_8 FILLER_6_165 ();
 sg13g2_decap_8 FILLER_6_172 ();
 sg13g2_decap_8 FILLER_6_179 ();
 sg13g2_decap_8 FILLER_6_186 ();
 sg13g2_decap_8 FILLER_6_193 ();
 sg13g2_decap_8 FILLER_6_200 ();
 sg13g2_decap_8 FILLER_6_207 ();
 sg13g2_decap_8 FILLER_6_214 ();
 sg13g2_decap_8 FILLER_6_221 ();
 sg13g2_decap_8 FILLER_6_228 ();
 sg13g2_decap_8 FILLER_6_235 ();
 sg13g2_decap_8 FILLER_6_242 ();
 sg13g2_decap_8 FILLER_6_249 ();
 sg13g2_decap_8 FILLER_6_256 ();
 sg13g2_decap_8 FILLER_6_263 ();
 sg13g2_decap_8 FILLER_6_270 ();
 sg13g2_decap_8 FILLER_6_277 ();
 sg13g2_decap_8 FILLER_6_284 ();
 sg13g2_decap_8 FILLER_6_291 ();
 sg13g2_decap_8 FILLER_6_298 ();
 sg13g2_decap_8 FILLER_6_305 ();
 sg13g2_decap_8 FILLER_6_312 ();
 sg13g2_decap_8 FILLER_6_319 ();
 sg13g2_decap_8 FILLER_6_326 ();
 sg13g2_decap_8 FILLER_6_333 ();
 sg13g2_decap_8 FILLER_6_340 ();
 sg13g2_decap_8 FILLER_6_347 ();
 sg13g2_decap_8 FILLER_6_354 ();
 sg13g2_decap_8 FILLER_6_361 ();
 sg13g2_decap_8 FILLER_6_368 ();
 sg13g2_decap_8 FILLER_6_375 ();
 sg13g2_decap_8 FILLER_6_382 ();
 sg13g2_decap_8 FILLER_6_389 ();
 sg13g2_decap_8 FILLER_6_396 ();
 sg13g2_decap_4 FILLER_6_403 ();
 sg13g2_fill_2 FILLER_6_407 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_fill_2 FILLER_7_28 ();
 sg13g2_fill_1 FILLER_7_30 ();
 sg13g2_fill_2 FILLER_7_35 ();
 sg13g2_fill_1 FILLER_7_37 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_fill_1 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_68 ();
 sg13g2_fill_2 FILLER_7_92 ();
 sg13g2_fill_1 FILLER_7_94 ();
 sg13g2_fill_2 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_111 ();
 sg13g2_decap_8 FILLER_7_118 ();
 sg13g2_decap_8 FILLER_7_125 ();
 sg13g2_decap_8 FILLER_7_132 ();
 sg13g2_decap_8 FILLER_7_139 ();
 sg13g2_decap_8 FILLER_7_146 ();
 sg13g2_decap_8 FILLER_7_153 ();
 sg13g2_decap_8 FILLER_7_160 ();
 sg13g2_decap_8 FILLER_7_167 ();
 sg13g2_decap_8 FILLER_7_174 ();
 sg13g2_decap_8 FILLER_7_181 ();
 sg13g2_decap_8 FILLER_7_188 ();
 sg13g2_decap_8 FILLER_7_195 ();
 sg13g2_decap_8 FILLER_7_202 ();
 sg13g2_decap_8 FILLER_7_209 ();
 sg13g2_decap_8 FILLER_7_216 ();
 sg13g2_decap_8 FILLER_7_223 ();
 sg13g2_decap_8 FILLER_7_230 ();
 sg13g2_decap_8 FILLER_7_237 ();
 sg13g2_decap_8 FILLER_7_244 ();
 sg13g2_decap_8 FILLER_7_251 ();
 sg13g2_decap_8 FILLER_7_258 ();
 sg13g2_decap_8 FILLER_7_265 ();
 sg13g2_decap_8 FILLER_7_272 ();
 sg13g2_decap_8 FILLER_7_279 ();
 sg13g2_decap_8 FILLER_7_286 ();
 sg13g2_decap_8 FILLER_7_293 ();
 sg13g2_decap_8 FILLER_7_300 ();
 sg13g2_decap_8 FILLER_7_307 ();
 sg13g2_decap_8 FILLER_7_314 ();
 sg13g2_decap_8 FILLER_7_321 ();
 sg13g2_decap_8 FILLER_7_328 ();
 sg13g2_decap_8 FILLER_7_335 ();
 sg13g2_decap_8 FILLER_7_342 ();
 sg13g2_decap_8 FILLER_7_349 ();
 sg13g2_decap_8 FILLER_7_356 ();
 sg13g2_decap_8 FILLER_7_363 ();
 sg13g2_decap_8 FILLER_7_370 ();
 sg13g2_decap_8 FILLER_7_377 ();
 sg13g2_decap_8 FILLER_7_384 ();
 sg13g2_decap_8 FILLER_7_391 ();
 sg13g2_decap_8 FILLER_7_398 ();
 sg13g2_decap_4 FILLER_7_405 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_fill_2 FILLER_8_21 ();
 sg13g2_fill_2 FILLER_8_54 ();
 sg13g2_fill_1 FILLER_8_56 ();
 sg13g2_fill_1 FILLER_8_71 ();
 sg13g2_decap_8 FILLER_8_125 ();
 sg13g2_decap_8 FILLER_8_132 ();
 sg13g2_decap_8 FILLER_8_139 ();
 sg13g2_decap_8 FILLER_8_146 ();
 sg13g2_decap_8 FILLER_8_153 ();
 sg13g2_decap_8 FILLER_8_160 ();
 sg13g2_decap_8 FILLER_8_167 ();
 sg13g2_decap_8 FILLER_8_174 ();
 sg13g2_decap_8 FILLER_8_181 ();
 sg13g2_decap_8 FILLER_8_188 ();
 sg13g2_decap_8 FILLER_8_195 ();
 sg13g2_decap_8 FILLER_8_202 ();
 sg13g2_decap_8 FILLER_8_209 ();
 sg13g2_decap_8 FILLER_8_216 ();
 sg13g2_decap_8 FILLER_8_223 ();
 sg13g2_decap_8 FILLER_8_230 ();
 sg13g2_decap_8 FILLER_8_237 ();
 sg13g2_decap_8 FILLER_8_244 ();
 sg13g2_decap_8 FILLER_8_251 ();
 sg13g2_decap_8 FILLER_8_258 ();
 sg13g2_decap_8 FILLER_8_265 ();
 sg13g2_decap_8 FILLER_8_272 ();
 sg13g2_decap_8 FILLER_8_279 ();
 sg13g2_decap_8 FILLER_8_286 ();
 sg13g2_decap_8 FILLER_8_293 ();
 sg13g2_decap_8 FILLER_8_300 ();
 sg13g2_decap_8 FILLER_8_307 ();
 sg13g2_decap_8 FILLER_8_314 ();
 sg13g2_decap_8 FILLER_8_321 ();
 sg13g2_decap_8 FILLER_8_328 ();
 sg13g2_decap_8 FILLER_8_335 ();
 sg13g2_decap_8 FILLER_8_342 ();
 sg13g2_decap_8 FILLER_8_349 ();
 sg13g2_decap_8 FILLER_8_356 ();
 sg13g2_decap_8 FILLER_8_363 ();
 sg13g2_decap_8 FILLER_8_370 ();
 sg13g2_decap_8 FILLER_8_377 ();
 sg13g2_decap_8 FILLER_8_384 ();
 sg13g2_decap_8 FILLER_8_391 ();
 sg13g2_decap_8 FILLER_8_398 ();
 sg13g2_decap_4 FILLER_8_405 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_fill_2 FILLER_9_50 ();
 sg13g2_fill_1 FILLER_9_52 ();
 sg13g2_decap_8 FILLER_9_136 ();
 sg13g2_decap_8 FILLER_9_143 ();
 sg13g2_decap_8 FILLER_9_150 ();
 sg13g2_decap_8 FILLER_9_157 ();
 sg13g2_decap_8 FILLER_9_164 ();
 sg13g2_decap_8 FILLER_9_171 ();
 sg13g2_decap_8 FILLER_9_178 ();
 sg13g2_decap_8 FILLER_9_185 ();
 sg13g2_decap_8 FILLER_9_192 ();
 sg13g2_decap_8 FILLER_9_199 ();
 sg13g2_decap_8 FILLER_9_206 ();
 sg13g2_decap_8 FILLER_9_213 ();
 sg13g2_decap_8 FILLER_9_220 ();
 sg13g2_decap_8 FILLER_9_227 ();
 sg13g2_decap_8 FILLER_9_234 ();
 sg13g2_decap_8 FILLER_9_241 ();
 sg13g2_decap_8 FILLER_9_248 ();
 sg13g2_decap_8 FILLER_9_255 ();
 sg13g2_decap_8 FILLER_9_262 ();
 sg13g2_decap_8 FILLER_9_269 ();
 sg13g2_decap_8 FILLER_9_276 ();
 sg13g2_decap_8 FILLER_9_283 ();
 sg13g2_decap_8 FILLER_9_290 ();
 sg13g2_decap_8 FILLER_9_297 ();
 sg13g2_decap_8 FILLER_9_304 ();
 sg13g2_decap_8 FILLER_9_311 ();
 sg13g2_decap_8 FILLER_9_318 ();
 sg13g2_decap_8 FILLER_9_325 ();
 sg13g2_decap_8 FILLER_9_332 ();
 sg13g2_decap_8 FILLER_9_339 ();
 sg13g2_decap_8 FILLER_9_346 ();
 sg13g2_decap_8 FILLER_9_353 ();
 sg13g2_decap_8 FILLER_9_360 ();
 sg13g2_decap_8 FILLER_9_367 ();
 sg13g2_decap_8 FILLER_9_374 ();
 sg13g2_decap_8 FILLER_9_381 ();
 sg13g2_decap_8 FILLER_9_388 ();
 sg13g2_decap_8 FILLER_9_395 ();
 sg13g2_decap_8 FILLER_9_402 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_fill_1 FILLER_10_61 ();
 sg13g2_fill_2 FILLER_10_106 ();
 sg13g2_fill_1 FILLER_10_108 ();
 sg13g2_fill_2 FILLER_10_118 ();
 sg13g2_decap_8 FILLER_10_146 ();
 sg13g2_decap_8 FILLER_10_153 ();
 sg13g2_decap_8 FILLER_10_160 ();
 sg13g2_decap_8 FILLER_10_167 ();
 sg13g2_decap_8 FILLER_10_174 ();
 sg13g2_decap_8 FILLER_10_181 ();
 sg13g2_decap_8 FILLER_10_188 ();
 sg13g2_decap_8 FILLER_10_195 ();
 sg13g2_decap_8 FILLER_10_202 ();
 sg13g2_decap_8 FILLER_10_209 ();
 sg13g2_decap_8 FILLER_10_216 ();
 sg13g2_decap_8 FILLER_10_223 ();
 sg13g2_decap_8 FILLER_10_230 ();
 sg13g2_decap_8 FILLER_10_237 ();
 sg13g2_decap_8 FILLER_10_244 ();
 sg13g2_decap_8 FILLER_10_251 ();
 sg13g2_decap_8 FILLER_10_258 ();
 sg13g2_decap_8 FILLER_10_265 ();
 sg13g2_decap_8 FILLER_10_272 ();
 sg13g2_decap_8 FILLER_10_279 ();
 sg13g2_decap_8 FILLER_10_286 ();
 sg13g2_decap_8 FILLER_10_293 ();
 sg13g2_decap_8 FILLER_10_300 ();
 sg13g2_decap_8 FILLER_10_307 ();
 sg13g2_decap_8 FILLER_10_314 ();
 sg13g2_decap_8 FILLER_10_321 ();
 sg13g2_decap_8 FILLER_10_328 ();
 sg13g2_decap_8 FILLER_10_335 ();
 sg13g2_decap_8 FILLER_10_342 ();
 sg13g2_decap_8 FILLER_10_349 ();
 sg13g2_decap_8 FILLER_10_356 ();
 sg13g2_decap_8 FILLER_10_363 ();
 sg13g2_decap_8 FILLER_10_370 ();
 sg13g2_decap_8 FILLER_10_377 ();
 sg13g2_decap_8 FILLER_10_384 ();
 sg13g2_decap_8 FILLER_10_391 ();
 sg13g2_decap_8 FILLER_10_398 ();
 sg13g2_decap_4 FILLER_10_405 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_4 FILLER_11_14 ();
 sg13g2_fill_2 FILLER_11_118 ();
 sg13g2_fill_1 FILLER_11_120 ();
 sg13g2_decap_8 FILLER_11_151 ();
 sg13g2_decap_8 FILLER_11_158 ();
 sg13g2_decap_8 FILLER_11_165 ();
 sg13g2_decap_8 FILLER_11_172 ();
 sg13g2_decap_8 FILLER_11_179 ();
 sg13g2_decap_8 FILLER_11_186 ();
 sg13g2_fill_2 FILLER_11_193 ();
 sg13g2_decap_8 FILLER_11_200 ();
 sg13g2_decap_4 FILLER_11_212 ();
 sg13g2_decap_8 FILLER_11_220 ();
 sg13g2_decap_8 FILLER_11_227 ();
 sg13g2_decap_8 FILLER_11_234 ();
 sg13g2_decap_8 FILLER_11_241 ();
 sg13g2_decap_8 FILLER_11_248 ();
 sg13g2_decap_8 FILLER_11_255 ();
 sg13g2_decap_8 FILLER_11_262 ();
 sg13g2_decap_8 FILLER_11_269 ();
 sg13g2_decap_8 FILLER_11_276 ();
 sg13g2_decap_8 FILLER_11_283 ();
 sg13g2_decap_8 FILLER_11_290 ();
 sg13g2_decap_8 FILLER_11_297 ();
 sg13g2_decap_8 FILLER_11_304 ();
 sg13g2_decap_8 FILLER_11_311 ();
 sg13g2_decap_8 FILLER_11_318 ();
 sg13g2_decap_8 FILLER_11_325 ();
 sg13g2_decap_8 FILLER_11_332 ();
 sg13g2_decap_8 FILLER_11_339 ();
 sg13g2_decap_8 FILLER_11_346 ();
 sg13g2_decap_8 FILLER_11_353 ();
 sg13g2_decap_8 FILLER_11_360 ();
 sg13g2_decap_8 FILLER_11_367 ();
 sg13g2_decap_8 FILLER_11_374 ();
 sg13g2_decap_8 FILLER_11_381 ();
 sg13g2_decap_8 FILLER_11_388 ();
 sg13g2_decap_8 FILLER_11_395 ();
 sg13g2_decap_8 FILLER_11_402 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_fill_2 FILLER_12_7 ();
 sg13g2_fill_1 FILLER_12_9 ();
 sg13g2_fill_1 FILLER_12_36 ();
 sg13g2_fill_2 FILLER_12_62 ();
 sg13g2_decap_8 FILLER_12_162 ();
 sg13g2_decap_8 FILLER_12_169 ();
 sg13g2_decap_8 FILLER_12_176 ();
 sg13g2_decap_8 FILLER_12_183 ();
 sg13g2_fill_2 FILLER_12_190 ();
 sg13g2_fill_2 FILLER_12_201 ();
 sg13g2_decap_4 FILLER_12_230 ();
 sg13g2_decap_8 FILLER_12_243 ();
 sg13g2_decap_8 FILLER_12_250 ();
 sg13g2_decap_8 FILLER_12_257 ();
 sg13g2_decap_8 FILLER_12_264 ();
 sg13g2_decap_8 FILLER_12_271 ();
 sg13g2_decap_8 FILLER_12_278 ();
 sg13g2_decap_8 FILLER_12_285 ();
 sg13g2_decap_8 FILLER_12_292 ();
 sg13g2_decap_8 FILLER_12_299 ();
 sg13g2_decap_8 FILLER_12_306 ();
 sg13g2_decap_8 FILLER_12_313 ();
 sg13g2_decap_8 FILLER_12_320 ();
 sg13g2_decap_8 FILLER_12_327 ();
 sg13g2_decap_8 FILLER_12_334 ();
 sg13g2_decap_8 FILLER_12_341 ();
 sg13g2_decap_8 FILLER_12_348 ();
 sg13g2_decap_8 FILLER_12_355 ();
 sg13g2_decap_8 FILLER_12_362 ();
 sg13g2_decap_8 FILLER_12_369 ();
 sg13g2_decap_8 FILLER_12_376 ();
 sg13g2_decap_8 FILLER_12_383 ();
 sg13g2_decap_8 FILLER_12_390 ();
 sg13g2_decap_8 FILLER_12_397 ();
 sg13g2_decap_4 FILLER_12_404 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_4 FILLER_13_7 ();
 sg13g2_fill_1 FILLER_13_11 ();
 sg13g2_fill_1 FILLER_13_57 ();
 sg13g2_fill_2 FILLER_13_63 ();
 sg13g2_fill_1 FILLER_13_65 ();
 sg13g2_fill_2 FILLER_13_92 ();
 sg13g2_fill_2 FILLER_13_129 ();
 sg13g2_fill_1 FILLER_13_131 ();
 sg13g2_decap_8 FILLER_13_167 ();
 sg13g2_decap_8 FILLER_13_174 ();
 sg13g2_decap_4 FILLER_13_181 ();
 sg13g2_fill_1 FILLER_13_185 ();
 sg13g2_decap_8 FILLER_13_247 ();
 sg13g2_decap_8 FILLER_13_254 ();
 sg13g2_decap_8 FILLER_13_261 ();
 sg13g2_decap_8 FILLER_13_268 ();
 sg13g2_decap_8 FILLER_13_275 ();
 sg13g2_decap_8 FILLER_13_282 ();
 sg13g2_decap_8 FILLER_13_289 ();
 sg13g2_decap_8 FILLER_13_296 ();
 sg13g2_decap_8 FILLER_13_303 ();
 sg13g2_decap_8 FILLER_13_310 ();
 sg13g2_decap_8 FILLER_13_317 ();
 sg13g2_decap_8 FILLER_13_324 ();
 sg13g2_decap_8 FILLER_13_331 ();
 sg13g2_decap_8 FILLER_13_338 ();
 sg13g2_decap_8 FILLER_13_345 ();
 sg13g2_decap_8 FILLER_13_352 ();
 sg13g2_decap_8 FILLER_13_359 ();
 sg13g2_decap_8 FILLER_13_366 ();
 sg13g2_decap_8 FILLER_13_373 ();
 sg13g2_decap_8 FILLER_13_380 ();
 sg13g2_decap_8 FILLER_13_387 ();
 sg13g2_decap_8 FILLER_13_394 ();
 sg13g2_decap_8 FILLER_13_401 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_4 FILLER_14_14 ();
 sg13g2_fill_2 FILLER_14_44 ();
 sg13g2_fill_2 FILLER_14_60 ();
 sg13g2_fill_1 FILLER_14_144 ();
 sg13g2_fill_2 FILLER_14_149 ();
 sg13g2_fill_2 FILLER_14_184 ();
 sg13g2_fill_1 FILLER_14_186 ();
 sg13g2_fill_2 FILLER_14_199 ();
 sg13g2_fill_1 FILLER_14_201 ();
 sg13g2_fill_2 FILLER_14_228 ();
 sg13g2_decap_8 FILLER_14_265 ();
 sg13g2_decap_8 FILLER_14_272 ();
 sg13g2_decap_8 FILLER_14_279 ();
 sg13g2_decap_8 FILLER_14_286 ();
 sg13g2_decap_8 FILLER_14_293 ();
 sg13g2_decap_8 FILLER_14_300 ();
 sg13g2_decap_8 FILLER_14_307 ();
 sg13g2_decap_8 FILLER_14_314 ();
 sg13g2_decap_8 FILLER_14_321 ();
 sg13g2_decap_8 FILLER_14_328 ();
 sg13g2_decap_8 FILLER_14_335 ();
 sg13g2_decap_8 FILLER_14_342 ();
 sg13g2_decap_8 FILLER_14_349 ();
 sg13g2_decap_8 FILLER_14_356 ();
 sg13g2_decap_8 FILLER_14_363 ();
 sg13g2_decap_8 FILLER_14_370 ();
 sg13g2_decap_8 FILLER_14_377 ();
 sg13g2_decap_8 FILLER_14_384 ();
 sg13g2_decap_8 FILLER_14_391 ();
 sg13g2_decap_8 FILLER_14_398 ();
 sg13g2_decap_4 FILLER_14_405 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_4 FILLER_15_21 ();
 sg13g2_fill_2 FILLER_15_25 ();
 sg13g2_fill_2 FILLER_15_109 ();
 sg13g2_fill_1 FILLER_15_111 ();
 sg13g2_fill_2 FILLER_15_166 ();
 sg13g2_fill_1 FILLER_15_179 ();
 sg13g2_fill_1 FILLER_15_194 ();
 sg13g2_fill_2 FILLER_15_207 ();
 sg13g2_fill_1 FILLER_15_209 ();
 sg13g2_decap_4 FILLER_15_236 ();
 sg13g2_fill_2 FILLER_15_249 ();
 sg13g2_fill_1 FILLER_15_251 ();
 sg13g2_decap_8 FILLER_15_261 ();
 sg13g2_decap_8 FILLER_15_268 ();
 sg13g2_decap_8 FILLER_15_275 ();
 sg13g2_decap_8 FILLER_15_282 ();
 sg13g2_decap_8 FILLER_15_289 ();
 sg13g2_decap_8 FILLER_15_296 ();
 sg13g2_decap_8 FILLER_15_303 ();
 sg13g2_decap_8 FILLER_15_310 ();
 sg13g2_decap_8 FILLER_15_317 ();
 sg13g2_decap_8 FILLER_15_324 ();
 sg13g2_decap_8 FILLER_15_331 ();
 sg13g2_decap_8 FILLER_15_338 ();
 sg13g2_decap_8 FILLER_15_345 ();
 sg13g2_decap_8 FILLER_15_352 ();
 sg13g2_decap_8 FILLER_15_359 ();
 sg13g2_decap_8 FILLER_15_366 ();
 sg13g2_decap_8 FILLER_15_373 ();
 sg13g2_decap_8 FILLER_15_380 ();
 sg13g2_decap_8 FILLER_15_387 ();
 sg13g2_decap_8 FILLER_15_394 ();
 sg13g2_decap_8 FILLER_15_401 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_4 FILLER_16_28 ();
 sg13g2_fill_2 FILLER_16_32 ();
 sg13g2_fill_2 FILLER_16_98 ();
 sg13g2_fill_2 FILLER_16_104 ();
 sg13g2_fill_1 FILLER_16_106 ();
 sg13g2_fill_1 FILLER_16_114 ();
 sg13g2_fill_2 FILLER_16_149 ();
 sg13g2_fill_1 FILLER_16_172 ();
 sg13g2_decap_8 FILLER_16_199 ();
 sg13g2_fill_1 FILLER_16_206 ();
 sg13g2_fill_2 FILLER_16_211 ();
 sg13g2_fill_1 FILLER_16_213 ();
 sg13g2_fill_2 FILLER_16_223 ();
 sg13g2_decap_4 FILLER_16_244 ();
 sg13g2_fill_1 FILLER_16_248 ();
 sg13g2_decap_8 FILLER_16_253 ();
 sg13g2_decap_8 FILLER_16_260 ();
 sg13g2_decap_8 FILLER_16_267 ();
 sg13g2_decap_8 FILLER_16_274 ();
 sg13g2_decap_8 FILLER_16_281 ();
 sg13g2_decap_8 FILLER_16_288 ();
 sg13g2_decap_8 FILLER_16_295 ();
 sg13g2_decap_8 FILLER_16_302 ();
 sg13g2_decap_8 FILLER_16_309 ();
 sg13g2_decap_8 FILLER_16_316 ();
 sg13g2_decap_8 FILLER_16_323 ();
 sg13g2_decap_8 FILLER_16_330 ();
 sg13g2_decap_8 FILLER_16_337 ();
 sg13g2_decap_8 FILLER_16_344 ();
 sg13g2_decap_8 FILLER_16_351 ();
 sg13g2_decap_8 FILLER_16_358 ();
 sg13g2_decap_8 FILLER_16_365 ();
 sg13g2_decap_8 FILLER_16_372 ();
 sg13g2_decap_8 FILLER_16_379 ();
 sg13g2_decap_8 FILLER_16_386 ();
 sg13g2_decap_8 FILLER_16_393 ();
 sg13g2_decap_8 FILLER_16_400 ();
 sg13g2_fill_2 FILLER_16_407 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_fill_1 FILLER_17_126 ();
 sg13g2_fill_1 FILLER_17_170 ();
 sg13g2_fill_1 FILLER_17_180 ();
 sg13g2_fill_2 FILLER_17_194 ();
 sg13g2_decap_4 FILLER_17_222 ();
 sg13g2_fill_1 FILLER_17_226 ();
 sg13g2_fill_1 FILLER_17_249 ();
 sg13g2_decap_8 FILLER_17_263 ();
 sg13g2_decap_8 FILLER_17_270 ();
 sg13g2_decap_8 FILLER_17_277 ();
 sg13g2_decap_8 FILLER_17_284 ();
 sg13g2_decap_8 FILLER_17_291 ();
 sg13g2_decap_8 FILLER_17_298 ();
 sg13g2_fill_2 FILLER_17_305 ();
 sg13g2_decap_8 FILLER_17_311 ();
 sg13g2_decap_8 FILLER_17_318 ();
 sg13g2_decap_8 FILLER_17_325 ();
 sg13g2_decap_8 FILLER_17_332 ();
 sg13g2_decap_8 FILLER_17_339 ();
 sg13g2_decap_8 FILLER_17_346 ();
 sg13g2_decap_8 FILLER_17_353 ();
 sg13g2_decap_8 FILLER_17_360 ();
 sg13g2_decap_8 FILLER_17_367 ();
 sg13g2_decap_8 FILLER_17_374 ();
 sg13g2_decap_8 FILLER_17_381 ();
 sg13g2_decap_8 FILLER_17_388 ();
 sg13g2_decap_8 FILLER_17_395 ();
 sg13g2_decap_8 FILLER_17_402 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_4 FILLER_18_77 ();
 sg13g2_fill_2 FILLER_18_81 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_fill_2 FILLER_18_98 ();
 sg13g2_fill_2 FILLER_18_113 ();
 sg13g2_fill_1 FILLER_18_115 ();
 sg13g2_fill_2 FILLER_18_271 ();
 sg13g2_decap_8 FILLER_18_277 ();
 sg13g2_fill_2 FILLER_18_284 ();
 sg13g2_fill_2 FILLER_18_296 ();
 sg13g2_fill_1 FILLER_18_298 ();
 sg13g2_fill_1 FILLER_18_325 ();
 sg13g2_decap_8 FILLER_18_352 ();
 sg13g2_decap_8 FILLER_18_359 ();
 sg13g2_decap_8 FILLER_18_366 ();
 sg13g2_decap_8 FILLER_18_373 ();
 sg13g2_decap_8 FILLER_18_380 ();
 sg13g2_decap_8 FILLER_18_387 ();
 sg13g2_decap_8 FILLER_18_394 ();
 sg13g2_decap_8 FILLER_18_401 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_4 FILLER_19_91 ();
 sg13g2_fill_1 FILLER_19_151 ();
 sg13g2_fill_1 FILLER_19_163 ();
 sg13g2_fill_2 FILLER_19_169 ();
 sg13g2_fill_1 FILLER_19_176 ();
 sg13g2_fill_2 FILLER_19_211 ();
 sg13g2_fill_1 FILLER_19_213 ();
 sg13g2_fill_2 FILLER_19_231 ();
 sg13g2_fill_1 FILLER_19_233 ();
 sg13g2_decap_4 FILLER_19_256 ();
 sg13g2_fill_2 FILLER_19_260 ();
 sg13g2_fill_2 FILLER_19_288 ();
 sg13g2_fill_1 FILLER_19_298 ();
 sg13g2_fill_2 FILLER_19_308 ();
 sg13g2_fill_1 FILLER_19_310 ();
 sg13g2_fill_2 FILLER_19_316 ();
 sg13g2_fill_1 FILLER_19_318 ();
 sg13g2_decap_8 FILLER_19_327 ();
 sg13g2_fill_2 FILLER_19_334 ();
 sg13g2_fill_1 FILLER_19_336 ();
 sg13g2_fill_2 FILLER_19_341 ();
 sg13g2_fill_1 FILLER_19_343 ();
 sg13g2_fill_2 FILLER_19_349 ();
 sg13g2_decap_8 FILLER_19_381 ();
 sg13g2_fill_2 FILLER_19_388 ();
 sg13g2_decap_8 FILLER_19_399 ();
 sg13g2_fill_2 FILLER_19_406 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_fill_2 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_fill_2 FILLER_20_135 ();
 sg13g2_fill_2 FILLER_20_142 ();
 sg13g2_fill_1 FILLER_20_149 ();
 sg13g2_fill_1 FILLER_20_161 ();
 sg13g2_fill_2 FILLER_20_230 ();
 sg13g2_fill_1 FILLER_20_232 ();
 sg13g2_fill_2 FILLER_20_247 ();
 sg13g2_fill_1 FILLER_20_249 ();
 sg13g2_fill_1 FILLER_20_260 ();
 sg13g2_fill_1 FILLER_20_274 ();
 sg13g2_fill_2 FILLER_20_335 ();
 sg13g2_decap_4 FILLER_20_345 ();
 sg13g2_fill_1 FILLER_20_349 ();
 sg13g2_fill_2 FILLER_20_354 ();
 sg13g2_fill_1 FILLER_20_356 ();
 sg13g2_fill_1 FILLER_20_375 ();
 sg13g2_fill_2 FILLER_20_407 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_4 FILLER_21_98 ();
 sg13g2_fill_2 FILLER_21_133 ();
 sg13g2_fill_2 FILLER_21_166 ();
 sg13g2_fill_1 FILLER_21_168 ();
 sg13g2_decap_8 FILLER_21_195 ();
 sg13g2_fill_1 FILLER_21_217 ();
 sg13g2_fill_2 FILLER_21_229 ();
 sg13g2_fill_1 FILLER_21_231 ();
 sg13g2_fill_1 FILLER_21_248 ();
 sg13g2_fill_2 FILLER_21_255 ();
 sg13g2_fill_1 FILLER_21_257 ();
 sg13g2_fill_2 FILLER_21_280 ();
 sg13g2_decap_8 FILLER_21_286 ();
 sg13g2_fill_2 FILLER_21_330 ();
 sg13g2_fill_1 FILLER_21_332 ();
 sg13g2_fill_2 FILLER_21_343 ();
 sg13g2_fill_1 FILLER_21_345 ();
 sg13g2_fill_1 FILLER_21_389 ();
 sg13g2_decap_4 FILLER_21_403 ();
 sg13g2_fill_2 FILLER_21_407 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_fill_1 FILLER_22_105 ();
 sg13g2_fill_1 FILLER_22_123 ();
 sg13g2_fill_1 FILLER_22_213 ();
 sg13g2_fill_2 FILLER_22_230 ();
 sg13g2_decap_4 FILLER_22_236 ();
 sg13g2_fill_2 FILLER_22_240 ();
 sg13g2_fill_1 FILLER_22_252 ();
 sg13g2_decap_4 FILLER_22_257 ();
 sg13g2_fill_2 FILLER_22_276 ();
 sg13g2_decap_8 FILLER_22_282 ();
 sg13g2_fill_2 FILLER_22_289 ();
 sg13g2_fill_1 FILLER_22_291 ();
 sg13g2_fill_2 FILLER_22_326 ();
 sg13g2_fill_2 FILLER_22_333 ();
 sg13g2_fill_2 FILLER_22_361 ();
 sg13g2_fill_1 FILLER_22_363 ();
 sg13g2_decap_8 FILLER_22_369 ();
 sg13g2_decap_8 FILLER_22_376 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_fill_2 FILLER_23_98 ();
 sg13g2_fill_1 FILLER_23_100 ();
 sg13g2_fill_2 FILLER_23_139 ();
 sg13g2_fill_1 FILLER_23_185 ();
 sg13g2_decap_4 FILLER_23_218 ();
 sg13g2_fill_1 FILLER_23_222 ();
 sg13g2_fill_1 FILLER_23_228 ();
 sg13g2_fill_1 FILLER_23_240 ();
 sg13g2_fill_1 FILLER_23_257 ();
 sg13g2_fill_2 FILLER_23_270 ();
 sg13g2_decap_4 FILLER_23_282 ();
 sg13g2_fill_1 FILLER_23_286 ();
 sg13g2_decap_4 FILLER_23_306 ();
 sg13g2_decap_8 FILLER_23_315 ();
 sg13g2_fill_2 FILLER_23_322 ();
 sg13g2_fill_1 FILLER_23_324 ();
 sg13g2_fill_2 FILLER_23_330 ();
 sg13g2_decap_4 FILLER_23_341 ();
 sg13g2_decap_8 FILLER_23_352 ();
 sg13g2_decap_4 FILLER_23_359 ();
 sg13g2_decap_4 FILLER_23_370 ();
 sg13g2_fill_2 FILLER_23_374 ();
 sg13g2_fill_1 FILLER_23_385 ();
 sg13g2_fill_2 FILLER_23_391 ();
 sg13g2_fill_1 FILLER_23_393 ();
 sg13g2_decap_4 FILLER_23_403 ();
 sg13g2_fill_2 FILLER_23_407 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_decap_4 FILLER_24_98 ();
 sg13g2_fill_1 FILLER_24_127 ();
 sg13g2_fill_1 FILLER_24_159 ();
 sg13g2_fill_1 FILLER_24_178 ();
 sg13g2_fill_2 FILLER_24_194 ();
 sg13g2_fill_1 FILLER_24_211 ();
 sg13g2_decap_8 FILLER_24_218 ();
 sg13g2_decap_8 FILLER_24_225 ();
 sg13g2_decap_8 FILLER_24_232 ();
 sg13g2_decap_4 FILLER_24_258 ();
 sg13g2_fill_2 FILLER_24_262 ();
 sg13g2_decap_8 FILLER_24_275 ();
 sg13g2_decap_4 FILLER_24_282 ();
 sg13g2_decap_8 FILLER_24_292 ();
 sg13g2_fill_2 FILLER_24_299 ();
 sg13g2_fill_1 FILLER_24_301 ();
 sg13g2_decap_8 FILLER_24_310 ();
 sg13g2_fill_2 FILLER_24_317 ();
 sg13g2_decap_4 FILLER_24_324 ();
 sg13g2_fill_2 FILLER_24_348 ();
 sg13g2_fill_1 FILLER_24_350 ();
 sg13g2_decap_4 FILLER_24_375 ();
 sg13g2_fill_2 FILLER_24_379 ();
 sg13g2_fill_1 FILLER_24_387 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_8 FILLER_25_91 ();
 sg13g2_decap_4 FILLER_25_98 ();
 sg13g2_fill_2 FILLER_25_128 ();
 sg13g2_fill_2 FILLER_25_139 ();
 sg13g2_fill_1 FILLER_25_193 ();
 sg13g2_fill_2 FILLER_25_198 ();
 sg13g2_fill_1 FILLER_25_200 ();
 sg13g2_fill_2 FILLER_25_207 ();
 sg13g2_decap_4 FILLER_25_216 ();
 sg13g2_fill_2 FILLER_25_234 ();
 sg13g2_fill_2 FILLER_25_255 ();
 sg13g2_fill_1 FILLER_25_257 ();
 sg13g2_decap_4 FILLER_25_280 ();
 sg13g2_fill_1 FILLER_25_305 ();
 sg13g2_fill_1 FILLER_25_322 ();
 sg13g2_decap_4 FILLER_25_329 ();
 sg13g2_fill_2 FILLER_25_338 ();
 sg13g2_fill_1 FILLER_25_340 ();
 sg13g2_fill_2 FILLER_25_370 ();
 sg13g2_fill_1 FILLER_25_372 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_decap_4 FILLER_26_91 ();
 sg13g2_fill_1 FILLER_26_95 ();
 sg13g2_decap_4 FILLER_26_99 ();
 sg13g2_fill_2 FILLER_26_168 ();
 sg13g2_fill_2 FILLER_26_179 ();
 sg13g2_fill_1 FILLER_26_181 ();
 sg13g2_fill_1 FILLER_26_198 ();
 sg13g2_fill_1 FILLER_26_208 ();
 sg13g2_decap_4 FILLER_26_226 ();
 sg13g2_fill_1 FILLER_26_247 ();
 sg13g2_fill_1 FILLER_26_254 ();
 sg13g2_fill_2 FILLER_26_268 ();
 sg13g2_fill_1 FILLER_26_279 ();
 sg13g2_fill_2 FILLER_26_285 ();
 sg13g2_fill_1 FILLER_26_287 ();
 sg13g2_decap_8 FILLER_26_292 ();
 sg13g2_fill_2 FILLER_26_314 ();
 sg13g2_fill_1 FILLER_26_316 ();
 sg13g2_fill_1 FILLER_26_323 ();
 sg13g2_decap_8 FILLER_26_344 ();
 sg13g2_decap_4 FILLER_26_351 ();
 sg13g2_fill_2 FILLER_26_355 ();
 sg13g2_fill_2 FILLER_26_360 ();
 sg13g2_fill_1 FILLER_26_362 ();
 sg13g2_decap_4 FILLER_26_370 ();
 sg13g2_fill_1 FILLER_26_374 ();
 sg13g2_fill_2 FILLER_26_381 ();
 sg13g2_fill_1 FILLER_26_408 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_fill_2 FILLER_27_56 ();
 sg13g2_fill_1 FILLER_27_58 ();
 sg13g2_decap_4 FILLER_27_85 ();
 sg13g2_fill_1 FILLER_27_191 ();
 sg13g2_fill_1 FILLER_27_202 ();
 sg13g2_fill_2 FILLER_27_223 ();
 sg13g2_decap_8 FILLER_27_228 ();
 sg13g2_decap_8 FILLER_27_245 ();
 sg13g2_decap_8 FILLER_27_252 ();
 sg13g2_decap_8 FILLER_27_271 ();
 sg13g2_fill_2 FILLER_27_278 ();
 sg13g2_fill_1 FILLER_27_280 ();
 sg13g2_decap_4 FILLER_27_285 ();
 sg13g2_fill_1 FILLER_27_299 ();
 sg13g2_fill_2 FILLER_27_310 ();
 sg13g2_fill_1 FILLER_27_312 ();
 sg13g2_decap_4 FILLER_27_345 ();
 sg13g2_fill_2 FILLER_27_355 ();
 sg13g2_decap_4 FILLER_27_378 ();
 sg13g2_fill_2 FILLER_27_407 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_fill_1 FILLER_28_42 ();
 sg13g2_fill_2 FILLER_28_48 ();
 sg13g2_decap_8 FILLER_28_53 ();
 sg13g2_fill_2 FILLER_28_60 ();
 sg13g2_fill_1 FILLER_28_66 ();
 sg13g2_fill_1 FILLER_28_115 ();
 sg13g2_fill_2 FILLER_28_191 ();
 sg13g2_fill_1 FILLER_28_226 ();
 sg13g2_fill_1 FILLER_28_251 ();
 sg13g2_fill_2 FILLER_28_265 ();
 sg13g2_fill_1 FILLER_28_267 ();
 sg13g2_fill_2 FILLER_28_284 ();
 sg13g2_fill_1 FILLER_28_286 ();
 sg13g2_fill_1 FILLER_28_291 ();
 sg13g2_decap_4 FILLER_28_297 ();
 sg13g2_fill_1 FILLER_28_311 ();
 sg13g2_fill_1 FILLER_28_321 ();
 sg13g2_fill_2 FILLER_28_330 ();
 sg13g2_fill_2 FILLER_28_353 ();
 sg13g2_fill_2 FILLER_28_398 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_fill_2 FILLER_29_28 ();
 sg13g2_fill_1 FILLER_29_30 ();
 sg13g2_fill_2 FILLER_29_35 ();
 sg13g2_fill_1 FILLER_29_46 ();
 sg13g2_fill_2 FILLER_29_117 ();
 sg13g2_fill_1 FILLER_29_119 ();
 sg13g2_fill_2 FILLER_29_138 ();
 sg13g2_fill_1 FILLER_29_140 ();
 sg13g2_fill_2 FILLER_29_146 ();
 sg13g2_fill_2 FILLER_29_170 ();
 sg13g2_fill_1 FILLER_29_172 ();
 sg13g2_decap_8 FILLER_29_199 ();
 sg13g2_fill_1 FILLER_29_206 ();
 sg13g2_decap_4 FILLER_29_224 ();
 sg13g2_fill_1 FILLER_29_228 ();
 sg13g2_fill_1 FILLER_29_238 ();
 sg13g2_fill_2 FILLER_29_259 ();
 sg13g2_decap_8 FILLER_29_266 ();
 sg13g2_decap_8 FILLER_29_273 ();
 sg13g2_fill_2 FILLER_29_297 ();
 sg13g2_fill_1 FILLER_29_305 ();
 sg13g2_fill_1 FILLER_29_316 ();
 sg13g2_fill_2 FILLER_29_327 ();
 sg13g2_fill_2 FILLER_29_339 ();
 sg13g2_fill_1 FILLER_29_341 ();
 sg13g2_fill_2 FILLER_29_354 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_4 FILLER_30_14 ();
 sg13g2_fill_2 FILLER_30_18 ();
 sg13g2_decap_4 FILLER_30_55 ();
 sg13g2_fill_2 FILLER_30_67 ();
 sg13g2_fill_1 FILLER_30_73 ();
 sg13g2_fill_1 FILLER_30_134 ();
 sg13g2_fill_1 FILLER_30_159 ();
 sg13g2_fill_2 FILLER_30_164 ();
 sg13g2_decap_8 FILLER_30_174 ();
 sg13g2_fill_2 FILLER_30_181 ();
 sg13g2_fill_1 FILLER_30_183 ();
 sg13g2_decap_8 FILLER_30_188 ();
 sg13g2_fill_1 FILLER_30_195 ();
 sg13g2_decap_8 FILLER_30_200 ();
 sg13g2_fill_1 FILLER_30_207 ();
 sg13g2_decap_8 FILLER_30_213 ();
 sg13g2_decap_8 FILLER_30_220 ();
 sg13g2_fill_2 FILLER_30_227 ();
 sg13g2_decap_4 FILLER_30_233 ();
 sg13g2_fill_1 FILLER_30_237 ();
 sg13g2_fill_2 FILLER_30_253 ();
 sg13g2_fill_1 FILLER_30_255 ();
 sg13g2_fill_1 FILLER_30_278 ();
 sg13g2_fill_2 FILLER_30_282 ();
 sg13g2_fill_1 FILLER_30_284 ();
 sg13g2_fill_1 FILLER_30_295 ();
 sg13g2_decap_8 FILLER_30_301 ();
 sg13g2_decap_8 FILLER_30_308 ();
 sg13g2_decap_8 FILLER_30_320 ();
 sg13g2_fill_1 FILLER_30_327 ();
 sg13g2_decap_8 FILLER_30_336 ();
 sg13g2_fill_1 FILLER_30_343 ();
 sg13g2_decap_8 FILLER_30_351 ();
 sg13g2_decap_4 FILLER_30_358 ();
 sg13g2_decap_8 FILLER_30_372 ();
 sg13g2_fill_2 FILLER_30_391 ();
 sg13g2_fill_1 FILLER_30_393 ();
 sg13g2_decap_4 FILLER_30_404 ();
 sg13g2_fill_1 FILLER_30_408 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_fill_2 FILLER_31_51 ();
 sg13g2_fill_1 FILLER_31_53 ();
 sg13g2_decap_8 FILLER_31_60 ();
 sg13g2_decap_4 FILLER_31_67 ();
 sg13g2_fill_2 FILLER_31_71 ();
 sg13g2_fill_2 FILLER_31_88 ();
 sg13g2_fill_1 FILLER_31_102 ();
 sg13g2_fill_2 FILLER_31_148 ();
 sg13g2_fill_1 FILLER_31_150 ();
 sg13g2_fill_2 FILLER_31_157 ();
 sg13g2_fill_1 FILLER_31_211 ();
 sg13g2_decap_4 FILLER_31_215 ();
 sg13g2_fill_2 FILLER_31_254 ();
 sg13g2_decap_4 FILLER_31_298 ();
 sg13g2_decap_4 FILLER_31_331 ();
 sg13g2_fill_1 FILLER_31_335 ();
 sg13g2_fill_2 FILLER_31_354 ();
 sg13g2_fill_1 FILLER_31_376 ();
 sg13g2_fill_2 FILLER_31_380 ();
 sg13g2_fill_1 FILLER_31_382 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_4 FILLER_32_35 ();
 sg13g2_fill_2 FILLER_32_54 ();
 sg13g2_fill_1 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_89 ();
 sg13g2_fill_2 FILLER_32_96 ();
 sg13g2_fill_2 FILLER_32_147 ();
 sg13g2_fill_1 FILLER_32_149 ();
 sg13g2_decap_8 FILLER_32_164 ();
 sg13g2_decap_4 FILLER_32_171 ();
 sg13g2_decap_8 FILLER_32_183 ();
 sg13g2_fill_2 FILLER_32_190 ();
 sg13g2_fill_1 FILLER_32_192 ();
 sg13g2_fill_1 FILLER_32_220 ();
 sg13g2_decap_4 FILLER_32_225 ();
 sg13g2_fill_2 FILLER_32_229 ();
 sg13g2_fill_1 FILLER_32_254 ();
 sg13g2_decap_8 FILLER_32_277 ();
 sg13g2_fill_2 FILLER_32_284 ();
 sg13g2_fill_1 FILLER_32_286 ();
 sg13g2_decap_8 FILLER_32_299 ();
 sg13g2_decap_4 FILLER_32_306 ();
 sg13g2_fill_1 FILLER_32_310 ();
 sg13g2_fill_1 FILLER_32_315 ();
 sg13g2_fill_1 FILLER_32_321 ();
 sg13g2_fill_2 FILLER_32_334 ();
 sg13g2_fill_2 FILLER_32_342 ();
 sg13g2_fill_1 FILLER_32_344 ();
 sg13g2_fill_2 FILLER_32_360 ();
 sg13g2_fill_1 FILLER_32_390 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_fill_1 FILLER_33_28 ();
 sg13g2_fill_1 FILLER_33_44 ();
 sg13g2_fill_2 FILLER_33_61 ();
 sg13g2_fill_1 FILLER_33_63 ();
 sg13g2_fill_1 FILLER_33_73 ();
 sg13g2_fill_1 FILLER_33_99 ();
 sg13g2_fill_2 FILLER_33_105 ();
 sg13g2_fill_2 FILLER_33_112 ();
 sg13g2_fill_1 FILLER_33_114 ();
 sg13g2_fill_1 FILLER_33_119 ();
 sg13g2_fill_1 FILLER_33_150 ();
 sg13g2_decap_8 FILLER_33_156 ();
 sg13g2_fill_2 FILLER_33_163 ();
 sg13g2_fill_2 FILLER_33_191 ();
 sg13g2_decap_8 FILLER_33_232 ();
 sg13g2_fill_2 FILLER_33_239 ();
 sg13g2_fill_1 FILLER_33_241 ();
 sg13g2_fill_1 FILLER_33_259 ();
 sg13g2_fill_1 FILLER_33_263 ();
 sg13g2_decap_8 FILLER_33_278 ();
 sg13g2_fill_2 FILLER_33_285 ();
 sg13g2_fill_2 FILLER_33_293 ();
 sg13g2_fill_2 FILLER_33_300 ();
 sg13g2_fill_2 FILLER_33_307 ();
 sg13g2_fill_2 FILLER_33_352 ();
 sg13g2_fill_2 FILLER_33_373 ();
 sg13g2_fill_1 FILLER_33_382 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_fill_2 FILLER_34_35 ();
 sg13g2_fill_2 FILLER_34_59 ();
 sg13g2_fill_2 FILLER_34_70 ();
 sg13g2_fill_1 FILLER_34_72 ();
 sg13g2_fill_1 FILLER_34_83 ();
 sg13g2_fill_1 FILLER_34_103 ();
 sg13g2_fill_2 FILLER_34_110 ();
 sg13g2_fill_1 FILLER_34_154 ();
 sg13g2_decap_4 FILLER_34_158 ();
 sg13g2_fill_2 FILLER_34_162 ();
 sg13g2_decap_4 FILLER_34_190 ();
 sg13g2_fill_1 FILLER_34_194 ();
 sg13g2_decap_4 FILLER_34_200 ();
 sg13g2_decap_8 FILLER_34_222 ();
 sg13g2_decap_8 FILLER_34_229 ();
 sg13g2_decap_4 FILLER_34_236 ();
 sg13g2_fill_2 FILLER_34_240 ();
 sg13g2_decap_8 FILLER_34_274 ();
 sg13g2_fill_1 FILLER_34_281 ();
 sg13g2_fill_1 FILLER_34_307 ();
 sg13g2_fill_2 FILLER_34_349 ();
 sg13g2_fill_1 FILLER_34_351 ();
 sg13g2_fill_2 FILLER_34_369 ();
 sg13g2_fill_2 FILLER_34_376 ();
 sg13g2_fill_1 FILLER_34_378 ();
 sg13g2_fill_1 FILLER_34_393 ();
 sg13g2_decap_8 FILLER_34_402 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_fill_2 FILLER_35_35 ();
 sg13g2_fill_2 FILLER_35_62 ();
 sg13g2_fill_1 FILLER_35_64 ();
 sg13g2_fill_1 FILLER_35_86 ();
 sg13g2_fill_1 FILLER_35_91 ();
 sg13g2_fill_2 FILLER_35_108 ();
 sg13g2_fill_2 FILLER_35_116 ();
 sg13g2_fill_1 FILLER_35_118 ();
 sg13g2_decap_4 FILLER_35_127 ();
 sg13g2_fill_1 FILLER_35_131 ();
 sg13g2_fill_2 FILLER_35_146 ();
 sg13g2_fill_1 FILLER_35_148 ();
 sg13g2_decap_8 FILLER_35_183 ();
 sg13g2_fill_2 FILLER_35_190 ();
 sg13g2_fill_2 FILLER_35_202 ();
 sg13g2_fill_2 FILLER_35_229 ();
 sg13g2_fill_2 FILLER_35_236 ();
 sg13g2_fill_2 FILLER_35_264 ();
 sg13g2_fill_2 FILLER_35_282 ();
 sg13g2_fill_2 FILLER_35_293 ();
 sg13g2_fill_1 FILLER_35_295 ();
 sg13g2_fill_1 FILLER_35_312 ();
 sg13g2_fill_1 FILLER_35_317 ();
 sg13g2_decap_4 FILLER_35_327 ();
 sg13g2_fill_2 FILLER_35_368 ();
 sg13g2_fill_1 FILLER_35_370 ();
 sg13g2_fill_2 FILLER_35_375 ();
 sg13g2_fill_1 FILLER_35_377 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_4 FILLER_36_35 ();
 sg13g2_fill_2 FILLER_36_39 ();
 sg13g2_fill_2 FILLER_36_50 ();
 sg13g2_fill_1 FILLER_36_52 ();
 sg13g2_decap_8 FILLER_36_67 ();
 sg13g2_decap_4 FILLER_36_74 ();
 sg13g2_fill_1 FILLER_36_95 ();
 sg13g2_fill_1 FILLER_36_100 ();
 sg13g2_fill_1 FILLER_36_105 ();
 sg13g2_decap_8 FILLER_36_110 ();
 sg13g2_fill_2 FILLER_36_117 ();
 sg13g2_fill_2 FILLER_36_145 ();
 sg13g2_fill_1 FILLER_36_147 ();
 sg13g2_decap_8 FILLER_36_152 ();
 sg13g2_fill_1 FILLER_36_159 ();
 sg13g2_decap_4 FILLER_36_164 ();
 sg13g2_fill_2 FILLER_36_198 ();
 sg13g2_fill_2 FILLER_36_218 ();
 sg13g2_fill_1 FILLER_36_220 ();
 sg13g2_decap_8 FILLER_36_226 ();
 sg13g2_fill_1 FILLER_36_233 ();
 sg13g2_decap_4 FILLER_36_239 ();
 sg13g2_fill_1 FILLER_36_273 ();
 sg13g2_decap_8 FILLER_36_330 ();
 sg13g2_fill_2 FILLER_36_337 ();
 sg13g2_fill_1 FILLER_36_359 ();
 sg13g2_decap_4 FILLER_36_405 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_4 FILLER_37_42 ();
 sg13g2_fill_1 FILLER_37_46 ();
 sg13g2_fill_2 FILLER_37_73 ();
 sg13g2_decap_4 FILLER_37_111 ();
 sg13g2_decap_8 FILLER_37_123 ();
 sg13g2_fill_2 FILLER_37_134 ();
 sg13g2_fill_1 FILLER_37_136 ();
 sg13g2_decap_8 FILLER_37_167 ();
 sg13g2_decap_8 FILLER_37_174 ();
 sg13g2_decap_8 FILLER_37_181 ();
 sg13g2_fill_2 FILLER_37_188 ();
 sg13g2_fill_2 FILLER_37_199 ();
 sg13g2_fill_2 FILLER_37_308 ();
 sg13g2_fill_1 FILLER_37_310 ();
 sg13g2_fill_2 FILLER_37_332 ();
 sg13g2_decap_8 FILLER_37_401 ();
 sg13g2_fill_1 FILLER_37_408 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_135 ();
 sg13g2_decap_8 FILLER_38_142 ();
 sg13g2_fill_1 FILLER_38_178 ();
 sg13g2_fill_1 FILLER_38_205 ();
 sg13g2_decap_4 FILLER_38_211 ();
 sg13g2_fill_1 FILLER_38_215 ();
 sg13g2_decap_8 FILLER_38_221 ();
 sg13g2_fill_2 FILLER_38_228 ();
 sg13g2_fill_1 FILLER_38_230 ();
 sg13g2_decap_8 FILLER_38_235 ();
 sg13g2_decap_8 FILLER_38_242 ();
 sg13g2_fill_1 FILLER_38_249 ();
 sg13g2_decap_8 FILLER_38_254 ();
 sg13g2_decap_8 FILLER_38_261 ();
 sg13g2_fill_2 FILLER_38_268 ();
 sg13g2_fill_1 FILLER_38_322 ();
 sg13g2_fill_1 FILLER_38_349 ();
 sg13g2_decap_8 FILLER_38_401 ();
 sg13g2_fill_1 FILLER_38_408 ();
 assign uio_oe[0] = net90;
 assign uio_oe[1] = net91;
 assign uio_oe[2] = net92;
 assign uio_oe[3] = net93;
 assign uio_oe[4] = net94;
 assign uio_oe[5] = net95;
 assign uio_oe[6] = net96;
 assign uio_oe[7] = net97;
endmodule

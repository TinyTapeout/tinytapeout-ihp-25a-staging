module tt_um_uart_mvm_sys (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire \MVM_UART_SYSTEM.AXIS_MVM.MATVEC.cen ;
 wire \MVM_UART_SYSTEM.AXIS_MVM.MATVEC.k_pad[0][0] ;
 wire \MVM_UART_SYSTEM.AXIS_MVM.MATVEC.k_pad[0][1] ;
 wire \MVM_UART_SYSTEM.AXIS_MVM.MATVEC.k_pad[1][0] ;
 wire \MVM_UART_SYSTEM.AXIS_MVM.MATVEC.k_pad[1][1] ;
 wire \MVM_UART_SYSTEM.AXIS_MVM.MATVEC.k_pad[2][0] ;
 wire \MVM_UART_SYSTEM.AXIS_MVM.MATVEC.k_pad[2][1] ;
 wire \MVM_UART_SYSTEM.AXIS_MVM.MATVEC.k_pad[3][0] ;
 wire \MVM_UART_SYSTEM.AXIS_MVM.MATVEC.k_pad[3][1] ;
 wire \MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[0][0] ;
 wire \MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[0][1] ;
 wire \MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[0][2] ;
 wire \MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[0][3] ;
 wire \MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[0][4] ;
 wire \MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[0][5] ;
 wire \MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[1][0] ;
 wire \MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[1][1] ;
 wire \MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[1][2] ;
 wire \MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[1][3] ;
 wire \MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[1][4] ;
 wire \MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[1][5] ;
 wire \MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[2][0] ;
 wire \MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[2][1] ;
 wire \MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[2][2] ;
 wire \MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[2][3] ;
 wire \MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[2][4] ;
 wire \MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[2][5] ;
 wire \MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[2][6] ;
 wire \MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[4][0] ;
 wire \MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[4][1] ;
 wire \MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[4][2] ;
 wire \MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[4][3] ;
 wire \MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[4][4] ;
 wire \MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[4][5] ;
 wire \MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[5][0] ;
 wire \MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[5][1] ;
 wire \MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[5][2] ;
 wire \MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[5][3] ;
 wire \MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[5][4] ;
 wire \MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[5][5] ;
 wire \MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[6][0] ;
 wire \MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[6][1] ;
 wire \MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[6][2] ;
 wire \MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[6][3] ;
 wire \MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[6][4] ;
 wire \MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[6][5] ;
 wire \MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[6][6] ;
 wire \MVM_UART_SYSTEM.AXIS_MVM.MATVEC.x_pad[0][0] ;
 wire \MVM_UART_SYSTEM.AXIS_MVM.MATVEC.x_pad[0][1] ;
 wire \MVM_UART_SYSTEM.AXIS_MVM.MATVEC.x_pad[0][2] ;
 wire \MVM_UART_SYSTEM.AXIS_MVM.MATVEC.x_pad[0][3] ;
 wire \MVM_UART_SYSTEM.AXIS_MVM.MATVEC.x_pad[1][0] ;
 wire \MVM_UART_SYSTEM.AXIS_MVM.MATVEC.x_pad[1][1] ;
 wire \MVM_UART_SYSTEM.AXIS_MVM.MATVEC.x_pad[1][2] ;
 wire \MVM_UART_SYSTEM.AXIS_MVM.MATVEC.x_pad[1][3] ;
 wire \MVM_UART_SYSTEM.AXIS_MVM.SKID.buffer[0] ;
 wire \MVM_UART_SYSTEM.AXIS_MVM.SKID.buffer[10] ;
 wire \MVM_UART_SYSTEM.AXIS_MVM.SKID.buffer[11] ;
 wire \MVM_UART_SYSTEM.AXIS_MVM.SKID.buffer[12] ;
 wire \MVM_UART_SYSTEM.AXIS_MVM.SKID.buffer[13] ;
 wire \MVM_UART_SYSTEM.AXIS_MVM.SKID.buffer[1] ;
 wire \MVM_UART_SYSTEM.AXIS_MVM.SKID.buffer[2] ;
 wire \MVM_UART_SYSTEM.AXIS_MVM.SKID.buffer[3] ;
 wire \MVM_UART_SYSTEM.AXIS_MVM.SKID.buffer[4] ;
 wire \MVM_UART_SYSTEM.AXIS_MVM.SKID.buffer[5] ;
 wire \MVM_UART_SYSTEM.AXIS_MVM.SKID.buffer[6] ;
 wire \MVM_UART_SYSTEM.AXIS_MVM.SKID.buffer[7] ;
 wire \MVM_UART_SYSTEM.AXIS_MVM.SKID.buffer[8] ;
 wire \MVM_UART_SYSTEM.AXIS_MVM.SKID.buffer[9] ;
 wire \MVM_UART_SYSTEM.AXIS_MVM.SKID.m_data[0] ;
 wire \MVM_UART_SYSTEM.AXIS_MVM.SKID.m_data[10] ;
 wire \MVM_UART_SYSTEM.AXIS_MVM.SKID.m_data[11] ;
 wire \MVM_UART_SYSTEM.AXIS_MVM.SKID.m_data[12] ;
 wire \MVM_UART_SYSTEM.AXIS_MVM.SKID.m_data[13] ;
 wire \MVM_UART_SYSTEM.AXIS_MVM.SKID.m_data[1] ;
 wire \MVM_UART_SYSTEM.AXIS_MVM.SKID.m_data[2] ;
 wire \MVM_UART_SYSTEM.AXIS_MVM.SKID.m_data[3] ;
 wire \MVM_UART_SYSTEM.AXIS_MVM.SKID.m_data[4] ;
 wire \MVM_UART_SYSTEM.AXIS_MVM.SKID.m_data[5] ;
 wire \MVM_UART_SYSTEM.AXIS_MVM.SKID.m_data[6] ;
 wire \MVM_UART_SYSTEM.AXIS_MVM.SKID.m_data[7] ;
 wire \MVM_UART_SYSTEM.AXIS_MVM.SKID.m_data[8] ;
 wire \MVM_UART_SYSTEM.AXIS_MVM.SKID.m_data[9] ;
 wire \MVM_UART_SYSTEM.AXIS_MVM.SKID.m_valid ;
 wire \MVM_UART_SYSTEM.AXIS_MVM.SKID.s_valid ;
 wire \MVM_UART_SYSTEM.AXIS_MVM.SKID.state[0] ;
 wire \MVM_UART_SYSTEM.AXIS_MVM.SKID.state[1] ;
 wire \MVM_UART_SYSTEM.AXIS_MVM.SKID.state_next[0] ;
 wire \MVM_UART_SYSTEM.AXIS_MVM.SKID.state_next[1] ;
 wire \MVM_UART_SYSTEM.AXIS_MVM.s_axis_kx_tvalid ;
 wire \MVM_UART_SYSTEM.AXIS_MVM.shift ;
 wire \MVM_UART_SYSTEM.UART_RX.c_bits[0] ;
 wire \MVM_UART_SYSTEM.UART_RX.c_bits[1] ;
 wire \MVM_UART_SYSTEM.UART_RX.c_bits[2] ;
 wire \MVM_UART_SYSTEM.UART_RX.c_clocks[0] ;
 wire \MVM_UART_SYSTEM.UART_RX.c_clocks[10] ;
 wire \MVM_UART_SYSTEM.UART_RX.c_clocks[11] ;
 wire \MVM_UART_SYSTEM.UART_RX.c_clocks[1] ;
 wire \MVM_UART_SYSTEM.UART_RX.c_clocks[2] ;
 wire \MVM_UART_SYSTEM.UART_RX.c_clocks[3] ;
 wire \MVM_UART_SYSTEM.UART_RX.c_clocks[4] ;
 wire \MVM_UART_SYSTEM.UART_RX.c_clocks[5] ;
 wire \MVM_UART_SYSTEM.UART_RX.c_clocks[6] ;
 wire \MVM_UART_SYSTEM.UART_RX.c_clocks[7] ;
 wire \MVM_UART_SYSTEM.UART_RX.c_clocks[8] ;
 wire \MVM_UART_SYSTEM.UART_RX.c_clocks[9] ;
 wire \MVM_UART_SYSTEM.UART_RX.c_words ;
 wire \MVM_UART_SYSTEM.UART_RX.state[0] ;
 wire \MVM_UART_SYSTEM.UART_RX.state[1] ;
 wire \MVM_UART_SYSTEM.UART_RX.state[2] ;
 wire \MVM_UART_SYSTEM.UART_RX.state[3] ;
 wire \MVM_UART_SYSTEM.UART_TX.c_clocks[0] ;
 wire \MVM_UART_SYSTEM.UART_TX.c_clocks[10] ;
 wire \MVM_UART_SYSTEM.UART_TX.c_clocks[11] ;
 wire \MVM_UART_SYSTEM.UART_TX.c_clocks[1] ;
 wire \MVM_UART_SYSTEM.UART_TX.c_clocks[2] ;
 wire \MVM_UART_SYSTEM.UART_TX.c_clocks[3] ;
 wire \MVM_UART_SYSTEM.UART_TX.c_clocks[4] ;
 wire \MVM_UART_SYSTEM.UART_TX.c_clocks[5] ;
 wire \MVM_UART_SYSTEM.UART_TX.c_clocks[6] ;
 wire \MVM_UART_SYSTEM.UART_TX.c_clocks[7] ;
 wire \MVM_UART_SYSTEM.UART_TX.c_clocks[8] ;
 wire \MVM_UART_SYSTEM.UART_TX.c_clocks[9] ;
 wire \MVM_UART_SYSTEM.UART_TX.c_pulses[0] ;
 wire \MVM_UART_SYSTEM.UART_TX.c_pulses[1] ;
 wire \MVM_UART_SYSTEM.UART_TX.c_pulses[2] ;
 wire \MVM_UART_SYSTEM.UART_TX.c_pulses[3] ;
 wire \MVM_UART_SYSTEM.UART_TX.c_pulses[4] ;
 wire \MVM_UART_SYSTEM.UART_TX.m_packets[0] ;
 wire \MVM_UART_SYSTEM.UART_TX.m_packets[10] ;
 wire \MVM_UART_SYSTEM.UART_TX.m_packets[11] ;
 wire \MVM_UART_SYSTEM.UART_TX.m_packets[12] ;
 wire \MVM_UART_SYSTEM.UART_TX.m_packets[13] ;
 wire \MVM_UART_SYSTEM.UART_TX.m_packets[14] ;
 wire \MVM_UART_SYSTEM.UART_TX.m_packets[15] ;
 wire \MVM_UART_SYSTEM.UART_TX.m_packets[16] ;
 wire \MVM_UART_SYSTEM.UART_TX.m_packets[17] ;
 wire \MVM_UART_SYSTEM.UART_TX.m_packets[18] ;
 wire \MVM_UART_SYSTEM.UART_TX.m_packets[19] ;
 wire \MVM_UART_SYSTEM.UART_TX.m_packets[1] ;
 wire \MVM_UART_SYSTEM.UART_TX.m_packets[20] ;
 wire \MVM_UART_SYSTEM.UART_TX.m_packets[21] ;
 wire \MVM_UART_SYSTEM.UART_TX.m_packets[22] ;
 wire \MVM_UART_SYSTEM.UART_TX.m_packets[23] ;
 wire \MVM_UART_SYSTEM.UART_TX.m_packets[24] ;
 wire \MVM_UART_SYSTEM.UART_TX.m_packets[25] ;
 wire \MVM_UART_SYSTEM.UART_TX.m_packets[2] ;
 wire \MVM_UART_SYSTEM.UART_TX.m_packets[3] ;
 wire \MVM_UART_SYSTEM.UART_TX.m_packets[4] ;
 wire \MVM_UART_SYSTEM.UART_TX.m_packets[5] ;
 wire \MVM_UART_SYSTEM.UART_TX.m_packets[6] ;
 wire \MVM_UART_SYSTEM.UART_TX.m_packets[7] ;
 wire \MVM_UART_SYSTEM.UART_TX.m_packets[8] ;
 wire \MVM_UART_SYSTEM.UART_TX.m_packets[9] ;
 wire \MVM_UART_SYSTEM.UART_TX.state ;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire clknet_0_clk;
 wire _0712_;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net1;
 wire net2;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_5_0__leaf_clk;
 wire clknet_5_1__leaf_clk;
 wire clknet_5_2__leaf_clk;
 wire clknet_5_3__leaf_clk;
 wire clknet_5_4__leaf_clk;
 wire clknet_5_5__leaf_clk;
 wire clknet_5_6__leaf_clk;
 wire clknet_5_7__leaf_clk;
 wire clknet_5_8__leaf_clk;
 wire clknet_5_9__leaf_clk;
 wire clknet_5_10__leaf_clk;
 wire clknet_5_11__leaf_clk;
 wire clknet_5_12__leaf_clk;
 wire clknet_5_13__leaf_clk;
 wire clknet_5_14__leaf_clk;
 wire clknet_5_15__leaf_clk;
 wire clknet_5_16__leaf_clk;
 wire clknet_5_17__leaf_clk;
 wire clknet_5_18__leaf_clk;
 wire clknet_5_19__leaf_clk;
 wire clknet_5_20__leaf_clk;
 wire clknet_5_21__leaf_clk;
 wire clknet_5_22__leaf_clk;
 wire clknet_5_23__leaf_clk;
 wire clknet_5_24__leaf_clk;
 wire clknet_5_25__leaf_clk;
 wire clknet_5_26__leaf_clk;
 wire clknet_5_27__leaf_clk;
 wire clknet_5_28__leaf_clk;
 wire clknet_5_29__leaf_clk;
 wire clknet_5_30__leaf_clk;
 wire clknet_5_31__leaf_clk;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;

 sg13g2_inv_1 _0713_ (.Y(_0181_),
    .A(_0032_));
 sg13g2_inv_1 _0714_ (.Y(_0182_),
    .A(_0031_));
 sg13g2_inv_1 _0715_ (.Y(_0183_),
    .A(_0024_));
 sg13g2_inv_1 _0716_ (.Y(_0184_),
    .A(_0019_));
 sg13g2_inv_1 _0717_ (.Y(_0185_),
    .A(_0018_));
 sg13g2_inv_1 _0718_ (.Y(_0186_),
    .A(_0011_));
 sg13g2_inv_2 _0719_ (.Y(_0187_),
    .A(net199));
 sg13g2_inv_1 _0720_ (.Y(_0188_),
    .A(\MVM_UART_SYSTEM.UART_RX.state[3] ));
 sg13g2_inv_1 _0721_ (.Y(_0189_),
    .A(net373));
 sg13g2_inv_1 _0722_ (.Y(_0190_),
    .A(net377));
 sg13g2_inv_1 _0723_ (.Y(_0191_),
    .A(net303));
 sg13g2_inv_1 _0724_ (.Y(_0192_),
    .A(\MVM_UART_SYSTEM.UART_TX.c_clocks[5] ));
 sg13g2_inv_1 _0725_ (.Y(_0193_),
    .A(\MVM_UART_SYSTEM.UART_TX.c_clocks[9] ));
 sg13g2_inv_1 _0726_ (.Y(_0194_),
    .A(\MVM_UART_SYSTEM.UART_TX.c_clocks[11] ));
 sg13g2_inv_1 _0727_ (.Y(_0195_),
    .A(net92));
 sg13g2_inv_1 _0728_ (.Y(_0196_),
    .A(net384));
 sg13g2_inv_1 _0729_ (.Y(_0197_),
    .A(net261));
 sg13g2_inv_1 _0730_ (.Y(_0198_),
    .A(_0009_));
 sg13g2_inv_1 _0731_ (.Y(_0199_),
    .A(\MVM_UART_SYSTEM.AXIS_MVM.SKID.m_data[6] ));
 sg13g2_inv_1 _0732_ (.Y(_0200_),
    .A(\MVM_UART_SYSTEM.AXIS_MVM.SKID.m_data[13] ));
 sg13g2_inv_1 _0733_ (.Y(_0201_),
    .A(net241));
 sg13g2_inv_1 _0734_ (.Y(_0202_),
    .A(net271));
 sg13g2_inv_1 _0735_ (.Y(_0203_),
    .A(net345));
 sg13g2_inv_1 _0736_ (.Y(_0204_),
    .A(net318));
 sg13g2_inv_1 _0737_ (.Y(_0205_),
    .A(net330));
 sg13g2_inv_1 _0738_ (.Y(_0206_),
    .A(net344));
 sg13g2_inv_1 _0739_ (.Y(_0207_),
    .A(net356));
 sg13g2_inv_1 _0740_ (.Y(_0208_),
    .A(net311));
 sg13g2_inv_1 _0741_ (.Y(_0209_),
    .A(net335));
 sg13g2_inv_1 _0742_ (.Y(_0210_),
    .A(net334));
 sg13g2_inv_1 _0743_ (.Y(_0211_),
    .A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.x_pad[0][3] ));
 sg13g2_inv_1 _0744_ (.Y(_0212_),
    .A(net395));
 sg13g2_nand4_1 _0745_ (.B(net331),
    .C(_0191_),
    .A(_0190_),
    .Y(_0213_),
    .D(\MVM_UART_SYSTEM.UART_RX.c_clocks[11] ));
 sg13g2_or2_1 _0746_ (.X(_0214_),
    .B(\MVM_UART_SYSTEM.UART_RX.c_clocks[6] ),
    .A(net224));
 sg13g2_nand2_1 _0747_ (.Y(_0215_),
    .A(net282),
    .B(net347));
 sg13g2_nand2_1 _0748_ (.Y(_0216_),
    .A(\MVM_UART_SYSTEM.UART_RX.c_clocks[3] ),
    .B(net327));
 sg13g2_or2_1 _0749_ (.X(_0217_),
    .B(_0215_),
    .A(_0214_));
 sg13g2_or3_1 _0750_ (.A(\MVM_UART_SYSTEM.UART_RX.c_clocks[2] ),
    .B(\MVM_UART_SYSTEM.UART_RX.c_clocks[4] ),
    .C(_0216_),
    .X(_0218_));
 sg13g2_nor3_2 _0751_ (.A(_0213_),
    .B(_0217_),
    .C(_0218_),
    .Y(_0219_));
 sg13g2_inv_1 _0752_ (.Y(_0220_),
    .A(_0219_));
 sg13g2_nor3_1 _0753_ (.A(_0213_),
    .B(_0217_),
    .C(_0218_),
    .Y(_0221_));
 sg13g2_nand2_1 _0754_ (.Y(_0222_),
    .A(\MVM_UART_SYSTEM.UART_RX.state[3] ),
    .B(_0221_));
 sg13g2_a22oi_1 _0755_ (.Y(_0037_),
    .B1(_0219_),
    .B2(\MVM_UART_SYSTEM.UART_RX.state[3] ),
    .A2(net1),
    .A1(net81));
 sg13g2_nand2b_1 _0756_ (.Y(_0223_),
    .B(net291),
    .A_N(\MVM_UART_SYSTEM.AXIS_MVM.SKID.state[1] ));
 sg13g2_nand2_1 _0757_ (.Y(_0224_),
    .A(net342),
    .B(net199));
 sg13g2_nor2_1 _0758_ (.A(_0223_),
    .B(_0224_),
    .Y(_0225_));
 sg13g2_nand2_1 _0759_ (.Y(_0226_),
    .A(net400),
    .B(_0187_));
 sg13g2_nand3_1 _0760_ (.B(_0224_),
    .C(_0226_),
    .A(_0223_),
    .Y(_0227_));
 sg13g2_nor2b_1 _0761_ (.A(net183),
    .B_N(_0227_),
    .Y(\MVM_UART_SYSTEM.AXIS_MVM.SKID.state_next[0] ));
 sg13g2_nor2b_1 _0762_ (.A(\MVM_UART_SYSTEM.AXIS_MVM.SKID.state[0] ),
    .B_N(\MVM_UART_SYSTEM.AXIS_MVM.SKID.state[1] ),
    .Y(_0228_));
 sg13g2_a21oi_1 _0763_ (.A1(net199),
    .A2(net185),
    .Y(_0003_),
    .B1(net182));
 sg13g2_nand3b_1 _0764_ (.B(net342),
    .C(\MVM_UART_SYSTEM.AXIS_MVM.SKID.state[1] ),
    .Y(_0229_),
    .A_N(net291));
 sg13g2_nand2_1 _0765_ (.Y(\MVM_UART_SYSTEM.AXIS_MVM.SKID.state_next[1] ),
    .A(_0003_),
    .B(net343));
 sg13g2_nand2_1 _0766_ (.Y(_0230_),
    .A(\MVM_UART_SYSTEM.UART_TX.c_pulses[3] ),
    .B(\MVM_UART_SYSTEM.UART_TX.c_pulses[4] ));
 sg13g2_nor4_2 _0767_ (.A(\MVM_UART_SYSTEM.UART_TX.c_pulses[1] ),
    .B(_0196_),
    .C(\MVM_UART_SYSTEM.UART_TX.c_pulses[2] ),
    .Y(_0231_),
    .D(_0230_));
 sg13g2_nor4_1 _0768_ (.A(\MVM_UART_SYSTEM.UART_TX.c_clocks[4] ),
    .B(_0192_),
    .C(net100),
    .D(\MVM_UART_SYSTEM.UART_TX.c_clocks[6] ),
    .Y(_0232_));
 sg13g2_nand3b_1 _0769_ (.B(_0232_),
    .C(\MVM_UART_SYSTEM.UART_TX.c_clocks[3] ),
    .Y(_0233_),
    .A_N(\MVM_UART_SYSTEM.UART_TX.c_clocks[2] ));
 sg13g2_nor4_1 _0770_ (.A(\MVM_UART_SYSTEM.UART_TX.c_clocks[8] ),
    .B(_0193_),
    .C(\MVM_UART_SYSTEM.UART_TX.c_clocks[10] ),
    .D(_0194_),
    .Y(_0234_));
 sg13g2_nand3_1 _0771_ (.B(net399),
    .C(net367),
    .A(net200),
    .Y(_0235_));
 sg13g2_nand4_1 _0772_ (.B(\MVM_UART_SYSTEM.UART_TX.c_clocks[1] ),
    .C(\MVM_UART_SYSTEM.UART_TX.c_clocks[0] ),
    .A(net200),
    .Y(_0236_),
    .D(_0234_));
 sg13g2_nor2_2 _0773_ (.A(_0233_),
    .B(_0236_),
    .Y(_0237_));
 sg13g2_and2_1 _0774_ (.A(_0231_),
    .B(_0237_),
    .X(_0238_));
 sg13g2_nand3_1 _0775_ (.B(\MVM_UART_SYSTEM.UART_TX.c_clocks[0] ),
    .C(\MVM_UART_SYSTEM.UART_TX.c_clocks[3] ),
    .A(\MVM_UART_SYSTEM.UART_TX.c_clocks[1] ),
    .Y(_0239_));
 sg13g2_nor2_1 _0776_ (.A(\MVM_UART_SYSTEM.UART_TX.c_clocks[2] ),
    .B(_0239_),
    .Y(_0240_));
 sg13g2_and4_1 _0777_ (.A(net200),
    .B(_0232_),
    .C(_0234_),
    .D(_0240_),
    .X(_0241_));
 sg13g2_nand2_1 _0778_ (.Y(_0242_),
    .A(_0231_),
    .B(net178));
 sg13g2_a21oi_1 _0779_ (.A1(_0187_),
    .A2(_0195_),
    .Y(_0712_),
    .B1(_0238_));
 sg13g2_nand3_1 _0780_ (.B(\MVM_UART_SYSTEM.UART_RX.c_bits[0] ),
    .C(\MVM_UART_SYSTEM.UART_RX.c_bits[2] ),
    .A(\MVM_UART_SYSTEM.UART_RX.c_bits[1] ),
    .Y(_0243_));
 sg13g2_and2_1 _0781_ (.A(\MVM_UART_SYSTEM.UART_RX.state[1] ),
    .B(_0219_),
    .X(_0244_));
 sg13g2_nand3b_1 _0782_ (.B(net373),
    .C(net385),
    .Y(_0245_),
    .A_N(net374));
 sg13g2_nand2b_1 _0783_ (.Y(_0246_),
    .B(net347),
    .A_N(net282));
 sg13g2_nor4_1 _0784_ (.A(net327),
    .B(_0214_),
    .C(_0245_),
    .D(_0246_),
    .Y(_0247_));
 sg13g2_nor4_1 _0785_ (.A(_0190_),
    .B(\MVM_UART_SYSTEM.UART_RX.c_clocks[9] ),
    .C(_0191_),
    .D(\MVM_UART_SYSTEM.UART_RX.c_clocks[11] ),
    .Y(_0248_));
 sg13g2_and2_2 _0786_ (.A(_0247_),
    .B(_0248_),
    .X(_0249_));
 sg13g2_nand2_2 _0787_ (.Y(_0250_),
    .A(\MVM_UART_SYSTEM.UART_RX.state[1] ),
    .B(_0221_));
 sg13g2_inv_1 _0788_ (.Y(_0251_),
    .A(_0250_));
 sg13g2_a22oi_1 _0789_ (.Y(_0252_),
    .B1(_0249_),
    .B2(\MVM_UART_SYSTEM.UART_RX.state[2] ),
    .A2(net175),
    .A1(_0243_));
 sg13g2_o21ai_1 _0790_ (.B1(_0252_),
    .Y(_0000_),
    .A1(net79),
    .A2(_0219_));
 sg13g2_nand2b_1 _0791_ (.Y(_0253_),
    .B(net81),
    .A_N(net1));
 sg13g2_o21ai_1 _0792_ (.B1(_0253_),
    .Y(_0001_),
    .A1(net83),
    .A2(_0249_));
 sg13g2_nand3_1 _0793_ (.B(net360),
    .C(net175),
    .A(net361),
    .Y(_0254_));
 sg13g2_nand4_1 _0794_ (.B(net360),
    .C(net150),
    .A(net361),
    .Y(_0255_),
    .D(net175));
 sg13g2_o21ai_1 _0795_ (.B1(_0255_),
    .Y(_0002_),
    .A1(_0188_),
    .A2(_0219_));
 sg13g2_or2_1 _0796_ (.X(_0004_),
    .B(\MVM_UART_SYSTEM.AXIS_MVM.SKID.state_next[1] ),
    .A(_0227_));
 sg13g2_nor2_1 _0797_ (.A(net63),
    .B(_0255_),
    .Y(_0005_));
 sg13g2_xor2_1 _0798_ (.B(net175),
    .A(net360),
    .X(_0038_));
 sg13g2_a21o_1 _0799_ (.A2(net175),
    .A1(net360),
    .B1(net361),
    .X(_0256_));
 sg13g2_and2_1 _0800_ (.A(_0254_),
    .B(_0256_),
    .X(_0039_));
 sg13g2_xnor2_1 _0801_ (.Y(_0040_),
    .A(net150),
    .B(_0254_));
 sg13g2_xor2_1 _0802_ (.B(net367),
    .A(net200),
    .X(_0041_));
 sg13g2_a21o_1 _0803_ (.A2(net367),
    .A1(net199),
    .B1(net399),
    .X(_0257_));
 sg13g2_and2_1 _0804_ (.A(_0235_),
    .B(_0257_),
    .X(_0042_));
 sg13g2_and4_1 _0805_ (.A(net200),
    .B(net402),
    .C(\MVM_UART_SYSTEM.UART_TX.c_clocks[0] ),
    .D(net338),
    .X(_0258_));
 sg13g2_nor2b_1 _0806_ (.A(net338),
    .B_N(_0235_),
    .Y(_0259_));
 sg13g2_nor3_1 _0807_ (.A(_0241_),
    .B(net403),
    .C(net339),
    .Y(_0043_));
 sg13g2_and2_1 _0808_ (.A(net365),
    .B(_0258_),
    .X(_0260_));
 sg13g2_nor2_1 _0809_ (.A(net365),
    .B(_0258_),
    .Y(_0261_));
 sg13g2_nor3_1 _0810_ (.A(_0241_),
    .B(_0260_),
    .C(net366),
    .Y(_0044_));
 sg13g2_xor2_1 _0811_ (.B(_0260_),
    .A(net280),
    .X(_0045_));
 sg13g2_a21oi_1 _0812_ (.A1(\MVM_UART_SYSTEM.UART_TX.c_clocks[4] ),
    .A2(_0260_),
    .Y(_0262_),
    .B1(net244));
 sg13g2_and4_1 _0813_ (.A(\MVM_UART_SYSTEM.UART_TX.c_clocks[3] ),
    .B(\MVM_UART_SYSTEM.UART_TX.c_clocks[4] ),
    .C(net244),
    .D(_0258_),
    .X(_0263_));
 sg13g2_nor3_1 _0814_ (.A(net178),
    .B(net245),
    .C(_0263_),
    .Y(_0046_));
 sg13g2_xor2_1 _0815_ (.B(_0263_),
    .A(net266),
    .X(_0047_));
 sg13g2_and3_1 _0816_ (.X(_0264_),
    .A(net100),
    .B(net266),
    .C(_0263_));
 sg13g2_a21oi_1 _0817_ (.A1(\MVM_UART_SYSTEM.UART_TX.c_clocks[6] ),
    .A2(_0263_),
    .Y(_0265_),
    .B1(net100));
 sg13g2_nor2_1 _0818_ (.A(_0264_),
    .B(net101),
    .Y(_0048_));
 sg13g2_xor2_1 _0819_ (.B(_0264_),
    .A(net290),
    .X(_0049_));
 sg13g2_a21oi_1 _0820_ (.A1(\MVM_UART_SYSTEM.UART_TX.c_clocks[8] ),
    .A2(_0264_),
    .Y(_0266_),
    .B1(net158));
 sg13g2_and3_1 _0821_ (.X(_0267_),
    .A(\MVM_UART_SYSTEM.UART_TX.c_clocks[8] ),
    .B(net158),
    .C(_0264_));
 sg13g2_nor3_1 _0822_ (.A(net178),
    .B(net159),
    .C(_0267_),
    .Y(_0050_));
 sg13g2_and2_1 _0823_ (.A(net114),
    .B(_0267_),
    .X(_0268_));
 sg13g2_xor2_1 _0824_ (.B(_0267_),
    .A(net114),
    .X(_0051_));
 sg13g2_nor2_1 _0825_ (.A(net317),
    .B(_0268_),
    .Y(_0269_));
 sg13g2_a21oi_1 _0826_ (.A1(net317),
    .A2(_0268_),
    .Y(_0270_),
    .B1(net178));
 sg13g2_nor2b_1 _0827_ (.A(_0269_),
    .B_N(_0270_),
    .Y(_0052_));
 sg13g2_mux2_1 _0828_ (.A0(net229),
    .A1(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[2][0] ),
    .S(net183),
    .X(_0053_));
 sg13g2_mux2_1 _0829_ (.A0(net163),
    .A1(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[2][1] ),
    .S(net181),
    .X(_0054_));
 sg13g2_nor2_1 _0830_ (.A(\MVM_UART_SYSTEM.AXIS_MVM.SKID.buffer[2] ),
    .B(net181),
    .Y(_0271_));
 sg13g2_a21oi_1 _0831_ (.A1(_0201_),
    .A2(net181),
    .Y(_0055_),
    .B1(_0271_));
 sg13g2_mux2_1 _0832_ (.A0(net142),
    .A1(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[2][3] ),
    .S(net181),
    .X(_0056_));
 sg13g2_mux2_1 _0833_ (.A0(net268),
    .A1(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[2][4] ),
    .S(net181),
    .X(_0057_));
 sg13g2_mux2_1 _0834_ (.A0(net265),
    .A1(net110),
    .S(net181),
    .X(_0058_));
 sg13g2_mux2_1 _0835_ (.A0(net243),
    .A1(net235),
    .S(net181),
    .X(_0059_));
 sg13g2_mux2_1 _0836_ (.A0(net165),
    .A1(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[6][0] ),
    .S(net182),
    .X(_0060_));
 sg13g2_mux2_1 _0837_ (.A0(net132),
    .A1(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[6][1] ),
    .S(net181),
    .X(_0061_));
 sg13g2_nor2_1 _0838_ (.A(net118),
    .B(net182),
    .Y(_0272_));
 sg13g2_a21oi_1 _0839_ (.A1(_0202_),
    .A2(net182),
    .Y(_0062_),
    .B1(_0272_));
 sg13g2_mux2_1 _0840_ (.A0(net128),
    .A1(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[6][3] ),
    .S(net182),
    .X(_0063_));
 sg13g2_mux2_1 _0841_ (.A0(net233),
    .A1(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[6][4] ),
    .S(net182),
    .X(_0064_));
 sg13g2_mux2_1 _0842_ (.A0(net260),
    .A1(net237),
    .S(net182),
    .X(_0065_));
 sg13g2_mux2_1 _0843_ (.A0(net130),
    .A1(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[6][6] ),
    .S(net182),
    .X(_0066_));
 sg13g2_nor2_1 _0844_ (.A(\MVM_UART_SYSTEM.UART_RX.state[3] ),
    .B(\MVM_UART_SYSTEM.UART_RX.state[1] ),
    .Y(_0273_));
 sg13g2_or2_1 _0845_ (.X(_0274_),
    .B(\MVM_UART_SYSTEM.UART_RX.state[1] ),
    .A(\MVM_UART_SYSTEM.UART_RX.state[3] ));
 sg13g2_nand2_1 _0846_ (.Y(_0275_),
    .A(net83),
    .B(_0273_));
 sg13g2_nand2_1 _0847_ (.Y(_0276_),
    .A(\MVM_UART_SYSTEM.UART_RX.c_clocks[0] ),
    .B(net180));
 sg13g2_xor2_1 _0848_ (.B(net180),
    .A(net347),
    .X(_0067_));
 sg13g2_nand2_1 _0849_ (.Y(_0277_),
    .A(net282),
    .B(_0276_));
 sg13g2_and2_1 _0850_ (.A(_0249_),
    .B(_0273_),
    .X(_0278_));
 sg13g2_nand2b_1 _0851_ (.Y(_0279_),
    .B(net180),
    .A_N(_0246_));
 sg13g2_o21ai_1 _0852_ (.B1(net283),
    .Y(_0068_),
    .A1(_0278_),
    .A2(_0279_));
 sg13g2_nand2b_1 _0853_ (.Y(_0280_),
    .B(net179),
    .A_N(_0215_));
 sg13g2_nand3_1 _0854_ (.B(\MVM_UART_SYSTEM.UART_RX.c_clocks[0] ),
    .C(net373),
    .A(net282),
    .Y(_0281_));
 sg13g2_inv_1 _0855_ (.Y(_0282_),
    .A(_0281_));
 sg13g2_a21oi_1 _0856_ (.A1(net83),
    .A2(_0273_),
    .Y(_0283_),
    .B1(_0281_));
 sg13g2_nand2_2 _0857_ (.Y(_0284_),
    .A(_0222_),
    .B(_0250_));
 sg13g2_or3_1 _0858_ (.A(_0278_),
    .B(_0282_),
    .C(_0284_),
    .X(_0285_));
 sg13g2_a22oi_1 _0859_ (.Y(_0069_),
    .B1(_0285_),
    .B2(net180),
    .A2(_0280_),
    .A1(_0189_));
 sg13g2_nor2_1 _0860_ (.A(net374),
    .B(_0283_),
    .Y(_0286_));
 sg13g2_and2_1 _0861_ (.A(net374),
    .B(_0283_),
    .X(_0287_));
 sg13g2_nor3_1 _0862_ (.A(_0284_),
    .B(net375),
    .C(_0287_),
    .Y(_0070_));
 sg13g2_nor2_1 _0863_ (.A(net385),
    .B(net179),
    .Y(_0288_));
 sg13g2_a21oi_1 _0864_ (.A1(net374),
    .A2(_0282_),
    .Y(_0289_),
    .B1(net385));
 sg13g2_a221oi_1 _0865_ (.B2(net385),
    .C1(_0289_),
    .B1(_0287_),
    .A1(_0249_),
    .Y(_0290_),
    .A2(net179));
 sg13g2_a21oi_1 _0866_ (.A1(_0247_),
    .A2(_0274_),
    .Y(_0291_),
    .B1(_0290_));
 sg13g2_nor2_1 _0867_ (.A(_0288_),
    .B(_0291_),
    .Y(_0071_));
 sg13g2_a21oi_1 _0868_ (.A1(\MVM_UART_SYSTEM.UART_RX.c_clocks[4] ),
    .A2(_0287_),
    .Y(_0292_),
    .B1(net327));
 sg13g2_and3_1 _0869_ (.X(_0293_),
    .A(net401),
    .B(net327),
    .C(_0287_));
 sg13g2_nor3_1 _0870_ (.A(_0284_),
    .B(net328),
    .C(_0293_),
    .Y(_0072_));
 sg13g2_xor2_1 _0871_ (.B(_0293_),
    .A(net353),
    .X(_0073_));
 sg13g2_a21oi_1 _0872_ (.A1(\MVM_UART_SYSTEM.UART_RX.c_clocks[6] ),
    .A2(_0293_),
    .Y(_0294_),
    .B1(net224));
 sg13g2_nand3_1 _0873_ (.B(net353),
    .C(_0293_),
    .A(net224),
    .Y(_0295_));
 sg13g2_nor2b_1 _0874_ (.A(net225),
    .B_N(_0295_),
    .Y(_0074_));
 sg13g2_nand4_1 _0875_ (.B(net224),
    .C(\MVM_UART_SYSTEM.UART_RX.c_clocks[6] ),
    .A(\MVM_UART_SYSTEM.UART_RX.c_clocks[4] ),
    .Y(_0296_),
    .D(\MVM_UART_SYSTEM.UART_RX.c_clocks[8] ));
 sg13g2_nor3_2 _0876_ (.A(_0216_),
    .B(_0281_),
    .C(_0296_),
    .Y(_0297_));
 sg13g2_or2_1 _0877_ (.X(_0298_),
    .B(_0297_),
    .A(_0278_));
 sg13g2_a22oi_1 _0878_ (.Y(_0075_),
    .B1(_0298_),
    .B2(net179),
    .A2(_0295_),
    .A1(_0190_));
 sg13g2_a21oi_1 _0879_ (.A1(net179),
    .A2(_0297_),
    .Y(_0299_),
    .B1(net331));
 sg13g2_and3_1 _0880_ (.X(_0300_),
    .A(net331),
    .B(net179),
    .C(_0297_));
 sg13g2_nand2_1 _0881_ (.Y(_0301_),
    .A(\MVM_UART_SYSTEM.UART_RX.c_clocks[9] ),
    .B(_0297_));
 sg13g2_nor3_1 _0882_ (.A(_0284_),
    .B(net332),
    .C(_0300_),
    .Y(_0076_));
 sg13g2_nor2_1 _0883_ (.A(net303),
    .B(net179),
    .Y(_0302_));
 sg13g2_a22oi_1 _0884_ (.Y(_0303_),
    .B1(_0301_),
    .B2(_0191_),
    .A2(net179),
    .A1(_0249_));
 sg13g2_nand2_1 _0885_ (.Y(_0304_),
    .A(net303),
    .B(_0300_));
 sg13g2_a22oi_1 _0886_ (.Y(_0305_),
    .B1(_0303_),
    .B2(_0304_),
    .A2(_0274_),
    .A1(_0248_));
 sg13g2_nor2_1 _0887_ (.A(_0302_),
    .B(_0305_),
    .Y(_0077_));
 sg13g2_xor2_1 _0888_ (.B(_0304_),
    .A(net370),
    .X(_0306_));
 sg13g2_nor2_1 _0889_ (.A(_0284_),
    .B(_0306_),
    .Y(_0078_));
 sg13g2_mux2_1 _0890_ (.A0(net397),
    .A1(net394),
    .S(net173),
    .X(_0079_));
 sg13g2_mux2_1 _0891_ (.A0(net394),
    .A1(net389),
    .S(net173),
    .X(_0080_));
 sg13g2_nor2_1 _0892_ (.A(net389),
    .B(net173),
    .Y(_0307_));
 sg13g2_a21oi_1 _0893_ (.A1(_0211_),
    .A2(net173),
    .Y(_0081_),
    .B1(_0307_));
 sg13g2_nand2_1 _0894_ (.Y(_0308_),
    .A(net380),
    .B(_0251_));
 sg13g2_o21ai_1 _0895_ (.B1(net381),
    .Y(_0082_),
    .A1(_0211_),
    .A2(_0251_));
 sg13g2_mux2_1 _0896_ (.A0(net380),
    .A1(net387),
    .S(net174),
    .X(_0083_));
 sg13g2_mux2_1 _0897_ (.A0(net387),
    .A1(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.x_pad[1][2] ),
    .S(net174),
    .X(_0084_));
 sg13g2_nor2_1 _0898_ (.A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.x_pad[1][2] ),
    .B(net174),
    .Y(_0309_));
 sg13g2_a21oi_1 _0899_ (.A1(_0212_),
    .A2(net174),
    .Y(_0085_),
    .B1(_0309_));
 sg13g2_nand2_1 _0900_ (.Y(_0310_),
    .A(net348),
    .B(_0251_));
 sg13g2_o21ai_1 _0901_ (.B1(net349),
    .Y(_0086_),
    .A1(_0212_),
    .A2(_0251_));
 sg13g2_mux2_1 _0902_ (.A0(net348),
    .A1(net378),
    .S(net173),
    .X(_0087_));
 sg13g2_mux2_1 _0903_ (.A0(net378),
    .A1(net391),
    .S(net173),
    .X(_0088_));
 sg13g2_mux2_1 _0904_ (.A0(net391),
    .A1(net320),
    .S(net174),
    .X(_0089_));
 sg13g2_mux2_1 _0905_ (.A0(net320),
    .A1(net379),
    .S(net174),
    .X(_0090_));
 sg13g2_mux2_1 _0906_ (.A0(net379),
    .A1(net383),
    .S(net173),
    .X(_0091_));
 sg13g2_mux2_1 _0907_ (.A0(net383),
    .A1(net392),
    .S(net173),
    .X(_0092_));
 sg13g2_mux2_1 _0908_ (.A0(net392),
    .A1(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.k_pad[0][1] ),
    .S(net174),
    .X(_0093_));
 sg13g2_mux2_1 _0909_ (.A0(net398),
    .A1(net1),
    .S(net175),
    .X(_0094_));
 sg13g2_xnor2_1 _0910_ (.Y(_0095_),
    .A(_0196_),
    .B(net178));
 sg13g2_a21oi_1 _0911_ (.A1(\MVM_UART_SYSTEM.UART_TX.c_pulses[0] ),
    .A2(net178),
    .Y(_0311_),
    .B1(net287));
 sg13g2_and3_1 _0912_ (.X(_0312_),
    .A(net287),
    .B(\MVM_UART_SYSTEM.UART_TX.c_pulses[0] ),
    .C(net178));
 sg13g2_nor3_1 _0913_ (.A(_0238_),
    .B(net288),
    .C(_0312_),
    .Y(_0096_));
 sg13g2_xor2_1 _0914_ (.B(_0312_),
    .A(net315),
    .X(_0097_));
 sg13g2_a21oi_1 _0915_ (.A1(\MVM_UART_SYSTEM.UART_TX.c_pulses[2] ),
    .A2(_0312_),
    .Y(_0313_),
    .B1(net105));
 sg13g2_nand3_1 _0916_ (.B(net105),
    .C(_0312_),
    .A(\MVM_UART_SYSTEM.UART_TX.c_pulses[2] ),
    .Y(_0314_));
 sg13g2_nand2_1 _0917_ (.Y(_0315_),
    .A(_0242_),
    .B(_0314_));
 sg13g2_nor2_1 _0918_ (.A(net106),
    .B(_0315_),
    .Y(_0098_));
 sg13g2_a21oi_1 _0919_ (.A1(_0242_),
    .A2(_0314_),
    .Y(_0316_),
    .B1(_0197_));
 sg13g2_a21oi_1 _0920_ (.A1(_0197_),
    .A2(_0314_),
    .Y(_0099_),
    .B1(_0316_));
 sg13g2_a21oi_1 _0921_ (.A1(_0187_),
    .A2(net92),
    .Y(_0317_),
    .B1(net178));
 sg13g2_or2_1 _0922_ (.X(_0318_),
    .B(_0231_),
    .A(net103));
 sg13g2_a22oi_1 _0923_ (.Y(_0100_),
    .B1(_0318_),
    .B2(_0237_),
    .A2(net171),
    .A1(_0186_));
 sg13g2_nand2b_1 _0924_ (.Y(_0319_),
    .B(net200),
    .A_N(_0231_));
 sg13g2_or2_1 _0925_ (.X(_0320_),
    .B(net108),
    .A(net198));
 sg13g2_o21ai_1 _0926_ (.B1(_0320_),
    .Y(_0321_),
    .A1(\MVM_UART_SYSTEM.UART_TX.m_packets[2] ),
    .A2(net176));
 sg13g2_mux2_1 _0927_ (.A0(_0321_),
    .A1(net239),
    .S(net170),
    .X(_0101_));
 sg13g2_or2_1 _0928_ (.X(_0322_),
    .B(net122),
    .A(net198));
 sg13g2_o21ai_1 _0929_ (.B1(_0322_),
    .Y(_0323_),
    .A1(\MVM_UART_SYSTEM.UART_TX.m_packets[3] ),
    .A2(net176));
 sg13g2_mux2_1 _0930_ (.A0(_0323_),
    .A1(net247),
    .S(net168),
    .X(_0102_));
 sg13g2_or2_1 _0931_ (.X(_0324_),
    .B(net136),
    .A(net198));
 sg13g2_o21ai_1 _0932_ (.B1(_0324_),
    .Y(_0325_),
    .A1(\MVM_UART_SYSTEM.UART_TX.m_packets[4] ),
    .A2(net176));
 sg13g2_mux2_1 _0933_ (.A0(_0325_),
    .A1(net154),
    .S(net168),
    .X(_0103_));
 sg13g2_or2_1 _0934_ (.X(_0326_),
    .B(\MVM_UART_SYSTEM.AXIS_MVM.SKID.m_data[3] ),
    .A(net201));
 sg13g2_o21ai_1 _0935_ (.B1(_0326_),
    .Y(_0327_),
    .A1(\MVM_UART_SYSTEM.UART_TX.m_packets[5] ),
    .A2(net176));
 sg13g2_mux2_1 _0936_ (.A0(_0327_),
    .A1(net263),
    .S(net168),
    .X(_0104_));
 sg13g2_or2_1 _0937_ (.X(_0328_),
    .B(\MVM_UART_SYSTEM.AXIS_MVM.SKID.m_data[4] ),
    .A(net198));
 sg13g2_o21ai_1 _0938_ (.B1(_0328_),
    .Y(_0329_),
    .A1(\MVM_UART_SYSTEM.UART_TX.m_packets[6] ),
    .A2(net176));
 sg13g2_mux2_1 _0939_ (.A0(_0329_),
    .A1(net252),
    .S(net169),
    .X(_0105_));
 sg13g2_or2_1 _0940_ (.X(_0330_),
    .B(net126),
    .A(net198));
 sg13g2_o21ai_1 _0941_ (.B1(_0330_),
    .Y(_0331_),
    .A1(\MVM_UART_SYSTEM.UART_TX.m_packets[7] ),
    .A2(net176));
 sg13g2_mux2_1 _0942_ (.A0(_0331_),
    .A1(net227),
    .S(net169),
    .X(_0106_));
 sg13g2_or2_1 _0943_ (.X(_0332_),
    .B(net176),
    .A(net86));
 sg13g2_a21oi_2 _0944_ (.B1(net168),
    .Y(_0333_),
    .A2(_0199_),
    .A1(_0187_));
 sg13g2_a22oi_1 _0945_ (.Y(_0107_),
    .B1(_0332_),
    .B2(_0333_),
    .A2(net169),
    .A1(_0185_));
 sg13g2_or2_1 _0946_ (.X(_0334_),
    .B(net176),
    .A(net94));
 sg13g2_a22oi_1 _0947_ (.Y(_0108_),
    .B1(_0333_),
    .B2(_0334_),
    .A2(net169),
    .A1(_0184_));
 sg13g2_nand2_1 _0948_ (.Y(_0335_),
    .A(_0020_),
    .B(net169));
 sg13g2_or3_2 _0949_ (.A(_0009_),
    .B(_0231_),
    .C(net170),
    .X(_0336_));
 sg13g2_o21ai_1 _0950_ (.B1(_0335_),
    .Y(_0109_),
    .A1(net77),
    .A2(_0336_));
 sg13g2_nand2_1 _0951_ (.Y(_0337_),
    .A(_0021_),
    .B(net168));
 sg13g2_o21ai_1 _0952_ (.B1(_0337_),
    .Y(_0110_),
    .A1(net71),
    .A2(_0336_));
 sg13g2_nand2_1 _0953_ (.Y(_0338_),
    .A(_0022_),
    .B(net171));
 sg13g2_o21ai_1 _0954_ (.B1(_0338_),
    .Y(_0111_),
    .A1(net67),
    .A2(_0336_));
 sg13g2_nand2_1 _0955_ (.Y(_0339_),
    .A(_0023_),
    .B(net171));
 sg13g2_o21ai_1 _0956_ (.B1(_0339_),
    .Y(_0112_),
    .A1(net75),
    .A2(_0336_));
 sg13g2_or2_1 _0957_ (.X(_0340_),
    .B(_0231_),
    .A(net98));
 sg13g2_a22oi_1 _0958_ (.Y(_0113_),
    .B1(_0340_),
    .B2(_0237_),
    .A2(net172),
    .A1(_0183_));
 sg13g2_or2_1 _0959_ (.X(_0341_),
    .B(net146),
    .A(net198));
 sg13g2_o21ai_1 _0960_ (.B1(_0341_),
    .Y(_0342_),
    .A1(\MVM_UART_SYSTEM.UART_TX.m_packets[15] ),
    .A2(net177));
 sg13g2_mux2_1 _0961_ (.A0(_0342_),
    .A1(net156),
    .S(net170),
    .X(_0114_));
 sg13g2_or2_1 _0962_ (.X(_0343_),
    .B(net112),
    .A(net198));
 sg13g2_o21ai_1 _0963_ (.B1(_0343_),
    .Y(_0344_),
    .A1(\MVM_UART_SYSTEM.UART_TX.m_packets[16] ),
    .A2(net177));
 sg13g2_mux2_1 _0964_ (.A0(_0344_),
    .A1(net152),
    .S(net168),
    .X(_0115_));
 sg13g2_or2_1 _0965_ (.X(_0345_),
    .B(net134),
    .A(net198));
 sg13g2_o21ai_1 _0966_ (.B1(_0345_),
    .Y(_0346_),
    .A1(\MVM_UART_SYSTEM.UART_TX.m_packets[17] ),
    .A2(net177));
 sg13g2_mux2_1 _0967_ (.A0(_0346_),
    .A1(net140),
    .S(net168),
    .X(_0116_));
 sg13g2_or2_1 _0968_ (.X(_0347_),
    .B(net120),
    .A(net199));
 sg13g2_o21ai_1 _0969_ (.B1(_0347_),
    .Y(_0348_),
    .A1(\MVM_UART_SYSTEM.UART_TX.m_packets[18] ),
    .A2(net177));
 sg13g2_mux2_1 _0970_ (.A0(_0348_),
    .A1(net256),
    .S(net168),
    .X(_0117_));
 sg13g2_or2_1 _0971_ (.X(_0349_),
    .B(net124),
    .A(net199));
 sg13g2_o21ai_1 _0972_ (.B1(_0349_),
    .Y(_0350_),
    .A1(\MVM_UART_SYSTEM.UART_TX.m_packets[19] ),
    .A2(net177));
 sg13g2_mux2_1 _0973_ (.A0(_0350_),
    .A1(net254),
    .S(net170),
    .X(_0118_));
 sg13g2_or2_1 _0974_ (.X(_0351_),
    .B(net116),
    .A(net199));
 sg13g2_o21ai_1 _0975_ (.B1(_0351_),
    .Y(_0352_),
    .A1(\MVM_UART_SYSTEM.UART_TX.m_packets[20] ),
    .A2(net177));
 sg13g2_mux2_1 _0976_ (.A0(_0352_),
    .A1(net148),
    .S(net170),
    .X(_0119_));
 sg13g2_or2_1 _0977_ (.X(_0353_),
    .B(net177),
    .A(net90));
 sg13g2_a21oi_1 _0978_ (.A1(_0187_),
    .A2(_0200_),
    .Y(_0354_),
    .B1(net170));
 sg13g2_a22oi_1 _0979_ (.Y(_0120_),
    .B1(_0353_),
    .B2(_0354_),
    .A2(net170),
    .A1(_0182_));
 sg13g2_or2_1 _0980_ (.X(_0355_),
    .B(net177),
    .A(net96));
 sg13g2_a22oi_1 _0981_ (.Y(_0121_),
    .B1(_0354_),
    .B2(_0355_),
    .A2(net170),
    .A1(_0181_));
 sg13g2_nand2_1 _0982_ (.Y(_0356_),
    .A(_0033_),
    .B(net171));
 sg13g2_o21ai_1 _0983_ (.B1(_0356_),
    .Y(_0122_),
    .A1(net69),
    .A2(_0336_));
 sg13g2_nand2_1 _0984_ (.Y(_0357_),
    .A(_0034_),
    .B(net171));
 sg13g2_o21ai_1 _0985_ (.B1(_0357_),
    .Y(_0123_),
    .A1(net73),
    .A2(_0336_));
 sg13g2_nand2_1 _0986_ (.Y(_0358_),
    .A(_0035_),
    .B(net171));
 sg13g2_o21ai_1 _0987_ (.B1(_0358_),
    .Y(_0124_),
    .A1(net65),
    .A2(_0336_));
 sg13g2_nand2_1 _0988_ (.Y(_0359_),
    .A(net84),
    .B(net171));
 sg13g2_nand2_1 _0989_ (.Y(_0125_),
    .A(_0336_),
    .B(_0359_));
 sg13g2_nor3_1 _0990_ (.A(net79),
    .B(_0220_),
    .C(_0243_),
    .Y(_0360_));
 sg13g2_mux2_1 _0991_ (.A0(net88),
    .A1(net63),
    .S(_0360_),
    .X(_0126_));
 sg13g2_mux2_1 _0992_ (.A0(\MVM_UART_SYSTEM.AXIS_MVM.shift ),
    .A1(net231),
    .S(net196),
    .X(_0127_));
 sg13g2_nand3_1 _0993_ (.B(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.x_pad[1][0] ),
    .C(net188),
    .A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.k_pad[2][0] ),
    .Y(_0361_));
 sg13g2_o21ai_1 _0994_ (.B1(_0361_),
    .Y(_0128_),
    .A1(_0207_),
    .A2(net195));
 sg13g2_nor2_1 _0995_ (.A(net305),
    .B(net192),
    .Y(_0362_));
 sg13g2_nand2_1 _0996_ (.Y(_0363_),
    .A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.k_pad[2][0] ),
    .B(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.x_pad[1][1] ));
 sg13g2_nand2_1 _0997_ (.Y(_0364_),
    .A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.x_pad[1][0] ),
    .B(net320));
 sg13g2_xnor2_1 _0998_ (.Y(_0365_),
    .A(_0363_),
    .B(net321));
 sg13g2_a21oi_1 _0999_ (.A1(net187),
    .A2(net322),
    .Y(_0129_),
    .B1(_0362_));
 sg13g2_nand2b_1 _1000_ (.Y(_0366_),
    .B(net309),
    .A_N(net187));
 sg13g2_nand2_1 _1001_ (.Y(_0367_),
    .A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.x_pad[1][0] ),
    .B(_0363_));
 sg13g2_nor2b_1 _1002_ (.A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.x_pad[1][1] ),
    .B_N(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.k_pad[2][1] ),
    .Y(_0368_));
 sg13g2_nand2_1 _1003_ (.Y(_0369_),
    .A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.k_pad[2][0] ),
    .B(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.x_pad[1][2] ));
 sg13g2_nand3_1 _1004_ (.B(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.x_pad[1][2] ),
    .C(_0368_),
    .A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.k_pad[2][0] ),
    .Y(_0370_));
 sg13g2_xnor2_1 _1005_ (.Y(_0371_),
    .A(_0368_),
    .B(_0369_));
 sg13g2_a21oi_1 _1006_ (.A1(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.k_pad[2][1] ),
    .A2(_0367_),
    .Y(_0372_),
    .B1(_0371_));
 sg13g2_nand3_1 _1007_ (.B(_0367_),
    .C(_0371_),
    .A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.k_pad[2][1] ),
    .Y(_0373_));
 sg13g2_nand2_1 _1008_ (.Y(_0374_),
    .A(net187),
    .B(_0373_));
 sg13g2_o21ai_1 _1009_ (.B1(_0366_),
    .Y(_0130_),
    .A1(_0372_),
    .A2(_0374_));
 sg13g2_nor2_1 _1010_ (.A(net351),
    .B(net187),
    .Y(_0375_));
 sg13g2_nor2b_1 _1011_ (.A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.x_pad[1][2] ),
    .B_N(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.k_pad[2][1] ),
    .Y(_0376_));
 sg13g2_and2_1 _1012_ (.A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.k_pad[2][0] ),
    .B(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.x_pad[1][3] ),
    .X(_0377_));
 sg13g2_xnor2_1 _1013_ (.Y(_0378_),
    .A(_0376_),
    .B(_0377_));
 sg13g2_or2_1 _1014_ (.X(_0379_),
    .B(_0378_),
    .A(_0370_));
 sg13g2_xnor2_1 _1015_ (.Y(_0380_),
    .A(_0370_),
    .B(_0378_));
 sg13g2_or2_1 _1016_ (.X(_0381_),
    .B(_0380_),
    .A(_0373_));
 sg13g2_xnor2_1 _1017_ (.Y(_0382_),
    .A(_0373_),
    .B(_0380_));
 sg13g2_a21oi_1 _1018_ (.A1(net187),
    .A2(_0382_),
    .Y(_0131_),
    .B1(_0375_));
 sg13g2_a21oi_1 _1019_ (.A1(_0212_),
    .A2(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.k_pad[2][1] ),
    .Y(_0383_),
    .B1(_0377_));
 sg13g2_a21o_1 _1020_ (.A2(_0377_),
    .A1(_0376_),
    .B1(_0383_),
    .X(_0384_));
 sg13g2_nand3_1 _1021_ (.B(_0381_),
    .C(_0384_),
    .A(_0379_),
    .Y(_0385_));
 sg13g2_a21o_1 _1022_ (.A2(_0381_),
    .A1(_0379_),
    .B1(_0384_),
    .X(_0386_));
 sg13g2_nand3_1 _1023_ (.B(_0385_),
    .C(_0386_),
    .A(net187),
    .Y(_0387_));
 sg13g2_o21ai_1 _1024_ (.B1(_0387_),
    .Y(_0132_),
    .A1(_0209_),
    .A2(net192));
 sg13g2_nand2b_1 _1025_ (.Y(_0388_),
    .B(net297),
    .A_N(net192));
 sg13g2_o21ai_1 _1026_ (.B1(_0388_),
    .Y(_0133_),
    .A1(_0383_),
    .A2(_0387_));
 sg13g2_nand2_1 _1027_ (.Y(_0389_),
    .A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[1][0] ),
    .B(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[0][0] ));
 sg13g2_xnor2_1 _1028_ (.Y(_0390_),
    .A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[1][0] ),
    .B(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[0][0] ));
 sg13g2_nor2_1 _1029_ (.A(net258),
    .B(net194),
    .Y(_0391_));
 sg13g2_a21oi_1 _1030_ (.A1(net194),
    .A2(_0390_),
    .Y(_0134_),
    .B1(_0391_));
 sg13g2_nor2_1 _1031_ (.A(net276),
    .B(net194),
    .Y(_0392_));
 sg13g2_nand2_1 _1032_ (.Y(_0393_),
    .A(net305),
    .B(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[0][1] ));
 sg13g2_xnor2_1 _1033_ (.Y(_0394_),
    .A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[1][1] ),
    .B(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[0][1] ));
 sg13g2_or2_1 _1034_ (.X(_0395_),
    .B(_0394_),
    .A(_0389_));
 sg13g2_xnor2_1 _1035_ (.Y(_0396_),
    .A(_0389_),
    .B(_0394_));
 sg13g2_a21oi_1 _1036_ (.A1(net192),
    .A2(_0396_),
    .Y(_0135_),
    .B1(_0392_));
 sg13g2_nand2_1 _1037_ (.Y(_0397_),
    .A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[1][2] ),
    .B(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[0][2] ));
 sg13g2_xnor2_1 _1038_ (.Y(_0398_),
    .A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[1][2] ),
    .B(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[0][2] ));
 sg13g2_nand3_1 _1039_ (.B(_0395_),
    .C(_0398_),
    .A(net306),
    .Y(_0399_));
 sg13g2_a21o_1 _1040_ (.A2(_0395_),
    .A1(_0393_),
    .B1(_0398_),
    .X(_0400_));
 sg13g2_nand3_1 _1041_ (.B(_0399_),
    .C(_0400_),
    .A(net192),
    .Y(_0401_));
 sg13g2_o21ai_1 _1042_ (.B1(_0401_),
    .Y(_0136_),
    .A1(_0201_),
    .A2(net192));
 sg13g2_nor2_1 _1043_ (.A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[1][3] ),
    .B(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[0][3] ),
    .Y(_0402_));
 sg13g2_xor2_1 _1044_ (.B(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[0][3] ),
    .A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[1][3] ),
    .X(_0403_));
 sg13g2_nand2_1 _1045_ (.Y(_0404_),
    .A(_0397_),
    .B(_0400_));
 sg13g2_xnor2_1 _1046_ (.Y(_0405_),
    .A(_0403_),
    .B(_0404_));
 sg13g2_nor2_1 _1047_ (.A(net299),
    .B(net193),
    .Y(_0406_));
 sg13g2_a21oi_1 _1048_ (.A1(net193),
    .A2(_0405_),
    .Y(_0137_),
    .B1(_0406_));
 sg13g2_a22oi_1 _1049_ (.Y(_0407_),
    .B1(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[1][3] ),
    .B2(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[0][3] ),
    .A2(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[0][2] ),
    .A1(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[1][2] ));
 sg13g2_a21oi_1 _1050_ (.A1(_0400_),
    .A2(_0407_),
    .Y(_0408_),
    .B1(_0402_));
 sg13g2_nor2_1 _1051_ (.A(_0209_),
    .B(_0210_),
    .Y(_0409_));
 sg13g2_xor2_1 _1052_ (.B(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[0][4] ),
    .A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[1][4] ),
    .X(_0410_));
 sg13g2_xnor2_1 _1053_ (.Y(_0411_),
    .A(_0408_),
    .B(_0410_));
 sg13g2_nor2_1 _1054_ (.A(net295),
    .B(net193),
    .Y(_0412_));
 sg13g2_a21oi_1 _1055_ (.A1(net193),
    .A2(_0411_),
    .Y(_0138_),
    .B1(_0412_));
 sg13g2_nor2_1 _1056_ (.A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[1][5] ),
    .B(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[0][5] ),
    .Y(_0413_));
 sg13g2_xnor2_1 _1057_ (.Y(_0414_),
    .A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[1][5] ),
    .B(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[0][5] ));
 sg13g2_a21oi_1 _1058_ (.A1(_0408_),
    .A2(_0410_),
    .Y(_0415_),
    .B1(_0409_));
 sg13g2_and2_1 _1059_ (.A(_0414_),
    .B(_0415_),
    .X(_0416_));
 sg13g2_o21ai_1 _1060_ (.B1(net193),
    .Y(_0417_),
    .A1(_0414_),
    .A2(_0415_));
 sg13g2_nand2b_1 _1061_ (.Y(_0418_),
    .B(net110),
    .A_N(net193));
 sg13g2_o21ai_1 _1062_ (.B1(_0418_),
    .Y(_0139_),
    .A1(_0416_),
    .A2(_0417_));
 sg13g2_nand2b_1 _1063_ (.Y(_0419_),
    .B(net235),
    .A_N(net193));
 sg13g2_o21ai_1 _1064_ (.B1(_0419_),
    .Y(_0140_),
    .A1(_0413_),
    .A2(_0417_));
 sg13g2_nand3_1 _1065_ (.B(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.k_pad[1][0] ),
    .C(net186),
    .A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.x_pad[0][0] ),
    .Y(_0420_));
 sg13g2_o21ai_1 _1066_ (.B1(_0420_),
    .Y(_0141_),
    .A1(_0204_),
    .A2(net195));
 sg13g2_nor2_1 _1067_ (.A(net336),
    .B(net189),
    .Y(_0421_));
 sg13g2_nand2_1 _1068_ (.Y(_0422_),
    .A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.k_pad[1][0] ),
    .B(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.x_pad[0][1] ));
 sg13g2_nand2_1 _1069_ (.Y(_0423_),
    .A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.x_pad[0][0] ),
    .B(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.k_pad[1][1] ));
 sg13g2_xnor2_1 _1070_ (.Y(_0424_),
    .A(_0422_),
    .B(_0423_));
 sg13g2_a21oi_1 _1071_ (.A1(net188),
    .A2(_0424_),
    .Y(_0142_),
    .B1(_0421_));
 sg13g2_nand2b_1 _1072_ (.Y(_0425_),
    .B(net354),
    .A_N(net190));
 sg13g2_nand2_1 _1073_ (.Y(_0426_),
    .A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.x_pad[0][0] ),
    .B(_0422_));
 sg13g2_nand2_1 _1074_ (.Y(_0427_),
    .A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.k_pad[1][0] ),
    .B(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.x_pad[0][2] ));
 sg13g2_nor2b_1 _1075_ (.A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.x_pad[0][1] ),
    .B_N(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.k_pad[1][1] ),
    .Y(_0428_));
 sg13g2_nand2b_1 _1076_ (.Y(_0429_),
    .B(_0428_),
    .A_N(_0427_));
 sg13g2_xnor2_1 _1077_ (.Y(_0430_),
    .A(_0427_),
    .B(_0428_));
 sg13g2_nand3_1 _1078_ (.B(_0426_),
    .C(_0430_),
    .A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.k_pad[1][1] ),
    .Y(_0431_));
 sg13g2_a21oi_1 _1079_ (.A1(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.k_pad[1][1] ),
    .A2(_0426_),
    .Y(_0432_),
    .B1(_0430_));
 sg13g2_nand2_1 _1080_ (.Y(_0433_),
    .A(net190),
    .B(_0431_));
 sg13g2_o21ai_1 _1081_ (.B1(_0425_),
    .Y(_0143_),
    .A1(_0432_),
    .A2(_0433_));
 sg13g2_nor2_1 _1082_ (.A(net372),
    .B(net190),
    .Y(_0434_));
 sg13g2_and2_1 _1083_ (.A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.k_pad[1][0] ),
    .B(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.x_pad[0][3] ),
    .X(_0435_));
 sg13g2_nor2b_1 _1084_ (.A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.x_pad[0][2] ),
    .B_N(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.k_pad[1][1] ),
    .Y(_0436_));
 sg13g2_xnor2_1 _1085_ (.Y(_0437_),
    .A(_0435_),
    .B(_0436_));
 sg13g2_or2_1 _1086_ (.X(_0438_),
    .B(_0437_),
    .A(_0429_));
 sg13g2_xnor2_1 _1087_ (.Y(_0439_),
    .A(_0429_),
    .B(_0437_));
 sg13g2_xnor2_1 _1088_ (.Y(_0440_),
    .A(_0431_),
    .B(_0439_));
 sg13g2_a21oi_1 _1089_ (.A1(net190),
    .A2(_0440_),
    .Y(_0144_),
    .B1(_0434_));
 sg13g2_a21oi_1 _1090_ (.A1(_0211_),
    .A2(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.k_pad[1][1] ),
    .Y(_0441_),
    .B1(_0435_));
 sg13g2_a21oi_1 _1091_ (.A1(_0435_),
    .A2(_0436_),
    .Y(_0442_),
    .B1(_0441_));
 sg13g2_o21ai_1 _1092_ (.B1(_0438_),
    .Y(_0443_),
    .A1(_0431_),
    .A2(_0439_));
 sg13g2_nor2_1 _1093_ (.A(_0442_),
    .B(_0443_),
    .Y(_0444_));
 sg13g2_nand2_1 _1094_ (.Y(_0445_),
    .A(_0442_),
    .B(_0443_));
 sg13g2_nand3b_1 _1095_ (.B(_0445_),
    .C(net190),
    .Y(_0446_),
    .A_N(_0444_));
 sg13g2_o21ai_1 _1096_ (.B1(_0446_),
    .Y(_0145_),
    .A1(_0206_),
    .A2(net190));
 sg13g2_nand2b_1 _1097_ (.Y(_0447_),
    .B(net293),
    .A_N(net190));
 sg13g2_o21ai_1 _1098_ (.B1(_0447_),
    .Y(_0146_),
    .A1(_0441_),
    .A2(_0446_));
 sg13g2_nand3_1 _1099_ (.B(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.k_pad[0][0] ),
    .C(net187),
    .A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.x_pad[1][0] ),
    .Y(_0448_));
 sg13g2_o21ai_1 _1100_ (.B1(_0448_),
    .Y(_0147_),
    .A1(_0203_),
    .A2(net192));
 sg13g2_nor2_1 _1101_ (.A(net325),
    .B(net196),
    .Y(_0449_));
 sg13g2_nand2_1 _1102_ (.Y(_0450_),
    .A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.k_pad[0][0] ),
    .B(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.x_pad[1][1] ));
 sg13g2_nand2_1 _1103_ (.Y(_0451_),
    .A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.x_pad[1][0] ),
    .B(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.k_pad[0][1] ));
 sg13g2_xnor2_1 _1104_ (.Y(_0452_),
    .A(_0450_),
    .B(_0451_));
 sg13g2_a21oi_1 _1105_ (.A1(net189),
    .A2(_0452_),
    .Y(_0148_),
    .B1(_0449_));
 sg13g2_nand2b_1 _1106_ (.Y(_0453_),
    .B(net323),
    .A_N(net189));
 sg13g2_nand2_1 _1107_ (.Y(_0454_),
    .A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.x_pad[1][0] ),
    .B(_0450_));
 sg13g2_nor2b_1 _1108_ (.A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.x_pad[1][1] ),
    .B_N(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.k_pad[0][1] ),
    .Y(_0455_));
 sg13g2_nand2_1 _1109_ (.Y(_0456_),
    .A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.k_pad[0][0] ),
    .B(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.x_pad[1][2] ));
 sg13g2_nand3_1 _1110_ (.B(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.x_pad[1][2] ),
    .C(_0455_),
    .A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.k_pad[0][0] ),
    .Y(_0457_));
 sg13g2_xnor2_1 _1111_ (.Y(_0458_),
    .A(_0455_),
    .B(_0456_));
 sg13g2_nand3_1 _1112_ (.B(_0454_),
    .C(_0458_),
    .A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.k_pad[0][1] ),
    .Y(_0459_));
 sg13g2_a21oi_1 _1113_ (.A1(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.k_pad[0][1] ),
    .A2(_0454_),
    .Y(_0460_),
    .B1(_0458_));
 sg13g2_nand2_1 _1114_ (.Y(_0461_),
    .A(net189),
    .B(_0459_));
 sg13g2_o21ai_1 _1115_ (.B1(_0453_),
    .Y(_0149_),
    .A1(_0460_),
    .A2(_0461_));
 sg13g2_nor2_1 _1116_ (.A(net358),
    .B(net191),
    .Y(_0462_));
 sg13g2_nor2b_1 _1117_ (.A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.x_pad[1][2] ),
    .B_N(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.k_pad[0][1] ),
    .Y(_0463_));
 sg13g2_and2_1 _1118_ (.A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.k_pad[0][0] ),
    .B(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.x_pad[1][3] ),
    .X(_0464_));
 sg13g2_xnor2_1 _1119_ (.Y(_0465_),
    .A(_0463_),
    .B(_0464_));
 sg13g2_or2_1 _1120_ (.X(_0466_),
    .B(_0465_),
    .A(_0457_));
 sg13g2_xnor2_1 _1121_ (.Y(_0467_),
    .A(_0457_),
    .B(_0465_));
 sg13g2_or2_1 _1122_ (.X(_0468_),
    .B(_0467_),
    .A(_0459_));
 sg13g2_xnor2_1 _1123_ (.Y(_0469_),
    .A(_0459_),
    .B(_0467_));
 sg13g2_a21oi_1 _1124_ (.A1(net189),
    .A2(_0469_),
    .Y(_0150_),
    .B1(net359));
 sg13g2_a21oi_1 _1125_ (.A1(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.k_pad[0][1] ),
    .A2(_0212_),
    .Y(_0470_),
    .B1(_0464_));
 sg13g2_a21o_1 _1126_ (.A2(_0464_),
    .A1(_0463_),
    .B1(_0470_),
    .X(_0471_));
 sg13g2_nand3_1 _1127_ (.B(_0468_),
    .C(_0471_),
    .A(_0466_),
    .Y(_0472_));
 sg13g2_a21o_1 _1128_ (.A2(_0468_),
    .A1(_0466_),
    .B1(_0471_),
    .X(_0473_));
 sg13g2_nand3_1 _1129_ (.B(_0472_),
    .C(_0473_),
    .A(net189),
    .Y(_0474_));
 sg13g2_o21ai_1 _1130_ (.B1(_0474_),
    .Y(_0151_),
    .A1(_0205_),
    .A2(net189));
 sg13g2_nand2b_1 _1131_ (.Y(_0475_),
    .B(net307),
    .A_N(net189));
 sg13g2_o21ai_1 _1132_ (.B1(_0475_),
    .Y(_0152_),
    .A1(_0470_),
    .A2(_0474_));
 sg13g2_nand2_1 _1133_ (.Y(_0476_),
    .A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[5][0] ),
    .B(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[4][0] ));
 sg13g2_xnor2_1 _1134_ (.Y(_0477_),
    .A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[5][0] ),
    .B(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[4][0] ));
 sg13g2_nor2_1 _1135_ (.A(net273),
    .B(net197),
    .Y(_0478_));
 sg13g2_a21oi_1 _1136_ (.A1(net197),
    .A2(_0477_),
    .Y(_0153_),
    .B1(net274));
 sg13g2_nor2_1 _1137_ (.A(net301),
    .B(net194),
    .Y(_0479_));
 sg13g2_nand2_1 _1138_ (.Y(_0480_),
    .A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[5][1] ),
    .B(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[4][1] ));
 sg13g2_xnor2_1 _1139_ (.Y(_0481_),
    .A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[5][1] ),
    .B(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[4][1] ));
 sg13g2_or2_1 _1140_ (.X(_0482_),
    .B(_0481_),
    .A(_0476_));
 sg13g2_xnor2_1 _1141_ (.Y(_0483_),
    .A(_0476_),
    .B(_0481_));
 sg13g2_a21oi_1 _1142_ (.A1(net193),
    .A2(_0483_),
    .Y(_0154_),
    .B1(_0479_));
 sg13g2_nand2_1 _1143_ (.Y(_0484_),
    .A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[5][2] ),
    .B(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[4][2] ));
 sg13g2_xnor2_1 _1144_ (.Y(_0485_),
    .A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[5][2] ),
    .B(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[4][2] ));
 sg13g2_nand3_1 _1145_ (.B(_0482_),
    .C(_0485_),
    .A(_0480_),
    .Y(_0486_));
 sg13g2_a21o_1 _1146_ (.A2(_0482_),
    .A1(_0480_),
    .B1(_0485_),
    .X(_0487_));
 sg13g2_nand3_1 _1147_ (.B(_0486_),
    .C(_0487_),
    .A(net196),
    .Y(_0488_));
 sg13g2_o21ai_1 _1148_ (.B1(_0488_),
    .Y(_0155_),
    .A1(_0202_),
    .A2(net196));
 sg13g2_nor2_1 _1149_ (.A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[5][3] ),
    .B(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[4][3] ),
    .Y(_0489_));
 sg13g2_xor2_1 _1150_ (.B(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[4][3] ),
    .A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[5][3] ),
    .X(_0490_));
 sg13g2_nand2_1 _1151_ (.Y(_0491_),
    .A(_0484_),
    .B(_0487_));
 sg13g2_xnor2_1 _1152_ (.Y(_0492_),
    .A(_0490_),
    .B(_0491_));
 sg13g2_nor2_1 _1153_ (.A(net161),
    .B(net196),
    .Y(_0493_));
 sg13g2_a21oi_1 _1154_ (.A1(net196),
    .A2(_0492_),
    .Y(_0156_),
    .B1(_0493_));
 sg13g2_nor2_1 _1155_ (.A(net249),
    .B(net197),
    .Y(_0494_));
 sg13g2_a22oi_1 _1156_ (.Y(_0495_),
    .B1(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[5][3] ),
    .B2(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[4][3] ),
    .A2(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[4][2] ),
    .A1(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[5][2] ));
 sg13g2_a21oi_1 _1157_ (.A1(_0487_),
    .A2(_0495_),
    .Y(_0496_),
    .B1(_0489_));
 sg13g2_nor2_1 _1158_ (.A(_0205_),
    .B(_0206_),
    .Y(_0497_));
 sg13g2_xor2_1 _1159_ (.B(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[4][4] ),
    .A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[5][4] ),
    .X(_0498_));
 sg13g2_xnor2_1 _1160_ (.Y(_0499_),
    .A(_0496_),
    .B(_0498_));
 sg13g2_a21oi_1 _1161_ (.A1(net197),
    .A2(_0499_),
    .Y(_0157_),
    .B1(net250));
 sg13g2_nor2_1 _1162_ (.A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[5][5] ),
    .B(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[4][5] ),
    .Y(_0500_));
 sg13g2_xnor2_1 _1163_ (.Y(_0501_),
    .A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[5][5] ),
    .B(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[4][5] ));
 sg13g2_a21oi_1 _1164_ (.A1(_0496_),
    .A2(_0498_),
    .Y(_0502_),
    .B1(_0497_));
 sg13g2_and2_1 _1165_ (.A(_0501_),
    .B(_0502_),
    .X(_0503_));
 sg13g2_o21ai_1 _1166_ (.B1(net190),
    .Y(_0504_),
    .A1(_0501_),
    .A2(_0502_));
 sg13g2_nand2b_1 _1167_ (.Y(_0505_),
    .B(net237),
    .A_N(net196));
 sg13g2_o21ai_1 _1168_ (.B1(_0505_),
    .Y(_0158_),
    .A1(_0503_),
    .A2(_0504_));
 sg13g2_nand2b_1 _1169_ (.Y(_0506_),
    .B(net138),
    .A_N(net196));
 sg13g2_o21ai_1 _1170_ (.B1(_0506_),
    .Y(_0159_),
    .A1(_0500_),
    .A2(_0504_));
 sg13g2_mux2_1 _1171_ (.A0(net291),
    .A1(\MVM_UART_SYSTEM.AXIS_MVM.shift ),
    .S(net197),
    .X(_0160_));
 sg13g2_nand3_1 _1172_ (.B(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.x_pad[0][0] ),
    .C(net188),
    .A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.k_pad[3][0] ),
    .Y(_0507_));
 sg13g2_o21ai_1 _1173_ (.B1(_0507_),
    .Y(_0161_),
    .A1(_0208_),
    .A2(net195));
 sg13g2_nor2_1 _1174_ (.A(net340),
    .B(net186),
    .Y(_0508_));
 sg13g2_nand2_1 _1175_ (.Y(_0509_),
    .A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.k_pad[3][0] ),
    .B(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.x_pad[0][1] ));
 sg13g2_nand2_1 _1176_ (.Y(_0510_),
    .A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.x_pad[0][0] ),
    .B(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.k_pad[3][1] ));
 sg13g2_xnor2_1 _1177_ (.Y(_0511_),
    .A(_0509_),
    .B(_0510_));
 sg13g2_a21oi_1 _1178_ (.A1(net186),
    .A2(_0511_),
    .Y(_0162_),
    .B1(_0508_));
 sg13g2_nand2b_1 _1179_ (.Y(_0512_),
    .B(net363),
    .A_N(net186));
 sg13g2_nand2_1 _1180_ (.Y(_0513_),
    .A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.x_pad[0][0] ),
    .B(_0509_));
 sg13g2_nand2_1 _1181_ (.Y(_0514_),
    .A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.k_pad[3][0] ),
    .B(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.x_pad[0][2] ));
 sg13g2_nor2b_1 _1182_ (.A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.x_pad[0][1] ),
    .B_N(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.k_pad[3][1] ),
    .Y(_0515_));
 sg13g2_nand2b_1 _1183_ (.Y(_0516_),
    .B(_0515_),
    .A_N(_0514_));
 sg13g2_xnor2_1 _1184_ (.Y(_0517_),
    .A(_0514_),
    .B(_0515_));
 sg13g2_a21oi_1 _1185_ (.A1(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.k_pad[3][1] ),
    .A2(_0513_),
    .Y(_0518_),
    .B1(_0517_));
 sg13g2_nand3_1 _1186_ (.B(_0513_),
    .C(_0517_),
    .A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.k_pad[3][1] ),
    .Y(_0519_));
 sg13g2_nand2_1 _1187_ (.Y(_0520_),
    .A(net186),
    .B(_0519_));
 sg13g2_o21ai_1 _1188_ (.B1(_0512_),
    .Y(_0163_),
    .A1(_0518_),
    .A2(_0520_));
 sg13g2_nor2_1 _1189_ (.A(net369),
    .B(net186),
    .Y(_0521_));
 sg13g2_and2_1 _1190_ (.A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.k_pad[3][0] ),
    .B(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.x_pad[0][3] ),
    .X(_0522_));
 sg13g2_nor2b_1 _1191_ (.A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.x_pad[0][2] ),
    .B_N(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.k_pad[3][1] ),
    .Y(_0523_));
 sg13g2_xnor2_1 _1192_ (.Y(_0524_),
    .A(_0522_),
    .B(_0523_));
 sg13g2_or2_1 _1193_ (.X(_0525_),
    .B(_0524_),
    .A(_0516_));
 sg13g2_xnor2_1 _1194_ (.Y(_0526_),
    .A(_0516_),
    .B(_0524_));
 sg13g2_xnor2_1 _1195_ (.Y(_0527_),
    .A(_0519_),
    .B(_0526_));
 sg13g2_a21oi_1 _1196_ (.A1(net186),
    .A2(_0527_),
    .Y(_0164_),
    .B1(_0521_));
 sg13g2_a21oi_1 _1197_ (.A1(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.k_pad[3][1] ),
    .A2(_0211_),
    .Y(_0528_),
    .B1(_0522_));
 sg13g2_a21oi_1 _1198_ (.A1(_0522_),
    .A2(_0523_),
    .Y(_0529_),
    .B1(_0528_));
 sg13g2_o21ai_1 _1199_ (.B1(_0525_),
    .Y(_0530_),
    .A1(_0519_),
    .A2(_0526_));
 sg13g2_nor2_1 _1200_ (.A(_0529_),
    .B(_0530_),
    .Y(_0531_));
 sg13g2_nand2_1 _1201_ (.Y(_0532_),
    .A(_0529_),
    .B(_0530_));
 sg13g2_nand3b_1 _1202_ (.B(_0532_),
    .C(net186),
    .Y(_0533_),
    .A_N(_0531_));
 sg13g2_o21ai_1 _1203_ (.B1(_0533_),
    .Y(_0165_),
    .A1(_0210_),
    .A2(net192));
 sg13g2_nand2b_1 _1204_ (.Y(_0534_),
    .B(net313),
    .A_N(net187));
 sg13g2_o21ai_1 _1205_ (.B1(_0534_),
    .Y(_0166_),
    .A1(_0528_),
    .A2(_0533_));
 sg13g2_a21o_1 _1206_ (.A2(_0198_),
    .A1(\MVM_UART_SYSTEM.AXIS_MVM.SKID.state[1] ),
    .B1(\MVM_UART_SYSTEM.AXIS_MVM.SKID.state[0] ),
    .X(_0535_));
 sg13g2_o21ai_1 _1207_ (.B1(_0535_),
    .Y(_0536_),
    .A1(net199),
    .A2(_0223_));
 sg13g2_and2_1 _1208_ (.A(_0004_),
    .B(_0536_),
    .X(_0537_));
 sg13g2_mux2_1 _1209_ (.A0(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[2][0] ),
    .A1(\MVM_UART_SYSTEM.AXIS_MVM.SKID.buffer[0] ),
    .S(net184),
    .X(_0538_));
 sg13g2_mux2_1 _1210_ (.A0(net108),
    .A1(_0538_),
    .S(net166),
    .X(_0167_));
 sg13g2_mux2_1 _1211_ (.A0(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[2][1] ),
    .A1(\MVM_UART_SYSTEM.AXIS_MVM.SKID.buffer[1] ),
    .S(net184),
    .X(_0539_));
 sg13g2_mux2_1 _1212_ (.A0(net122),
    .A1(_0539_),
    .S(net166),
    .X(_0168_));
 sg13g2_mux2_1 _1213_ (.A0(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[2][2] ),
    .A1(\MVM_UART_SYSTEM.AXIS_MVM.SKID.buffer[2] ),
    .S(net184),
    .X(_0540_));
 sg13g2_mux2_1 _1214_ (.A0(net136),
    .A1(_0540_),
    .S(net166),
    .X(_0169_));
 sg13g2_mux2_1 _1215_ (.A0(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[2][3] ),
    .A1(net142),
    .S(net184),
    .X(_0541_));
 sg13g2_mux2_1 _1216_ (.A0(net278),
    .A1(_0541_),
    .S(net166),
    .X(_0170_));
 sg13g2_mux2_1 _1217_ (.A0(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[2][4] ),
    .A1(net268),
    .S(net184),
    .X(_0542_));
 sg13g2_mux2_1 _1218_ (.A0(net285),
    .A1(_0542_),
    .S(net166),
    .X(_0171_));
 sg13g2_mux2_1 _1219_ (.A0(net110),
    .A1(\MVM_UART_SYSTEM.AXIS_MVM.SKID.buffer[5] ),
    .S(net184),
    .X(_0543_));
 sg13g2_mux2_1 _1220_ (.A0(net126),
    .A1(_0543_),
    .S(net166),
    .X(_0172_));
 sg13g2_mux2_1 _1221_ (.A0(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[2][6] ),
    .A1(\MVM_UART_SYSTEM.AXIS_MVM.SKID.buffer[6] ),
    .S(net184),
    .X(_0544_));
 sg13g2_mux2_1 _1222_ (.A0(net144),
    .A1(_0544_),
    .S(net166),
    .X(_0173_));
 sg13g2_mux2_1 _1223_ (.A0(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[6][0] ),
    .A1(\MVM_UART_SYSTEM.AXIS_MVM.SKID.buffer[7] ),
    .S(net185),
    .X(_0545_));
 sg13g2_mux2_1 _1224_ (.A0(net146),
    .A1(_0545_),
    .S(net167),
    .X(_0174_));
 sg13g2_mux2_1 _1225_ (.A0(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[6][1] ),
    .A1(\MVM_UART_SYSTEM.AXIS_MVM.SKID.buffer[8] ),
    .S(net184),
    .X(_0546_));
 sg13g2_mux2_1 _1226_ (.A0(net112),
    .A1(_0546_),
    .S(net166),
    .X(_0175_));
 sg13g2_mux2_1 _1227_ (.A0(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[6][2] ),
    .A1(net118),
    .S(net185),
    .X(_0547_));
 sg13g2_mux2_1 _1228_ (.A0(net134),
    .A1(_0547_),
    .S(net167),
    .X(_0176_));
 sg13g2_mux2_1 _1229_ (.A0(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[6][3] ),
    .A1(\MVM_UART_SYSTEM.AXIS_MVM.SKID.buffer[10] ),
    .S(net185),
    .X(_0548_));
 sg13g2_mux2_1 _1230_ (.A0(net120),
    .A1(_0548_),
    .S(net167),
    .X(_0177_));
 sg13g2_mux2_1 _1231_ (.A0(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[6][4] ),
    .A1(\MVM_UART_SYSTEM.AXIS_MVM.SKID.buffer[11] ),
    .S(net185),
    .X(_0549_));
 sg13g2_mux2_1 _1232_ (.A0(net124),
    .A1(_0549_),
    .S(net167),
    .X(_0178_));
 sg13g2_mux2_1 _1233_ (.A0(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[6][5] ),
    .A1(\MVM_UART_SYSTEM.AXIS_MVM.SKID.buffer[12] ),
    .S(net185),
    .X(_0550_));
 sg13g2_mux2_1 _1234_ (.A0(net116),
    .A1(_0550_),
    .S(net167),
    .X(_0179_));
 sg13g2_mux2_1 _1235_ (.A0(net138),
    .A1(net130),
    .S(net185),
    .X(_0551_));
 sg13g2_mux2_1 _1236_ (.A0(net270),
    .A1(_0551_),
    .S(net167),
    .X(_0180_));
 sg13g2_dfrbp_1 _1237_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net207),
    .D(_0038_),
    .Q_N(_0667_),
    .Q(\MVM_UART_SYSTEM.UART_RX.c_bits[0] ));
 sg13g2_dfrbp_1 _1238_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net207),
    .D(_0039_),
    .Q_N(_0666_),
    .Q(\MVM_UART_SYSTEM.UART_RX.c_bits[1] ));
 sg13g2_dfrbp_1 _1239_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net207),
    .D(net151),
    .Q_N(_0665_),
    .Q(\MVM_UART_SYSTEM.UART_RX.c_bits[2] ));
 sg13g2_dfrbp_1 _1240_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net220),
    .D(net368),
    .Q_N(_0664_),
    .Q(\MVM_UART_SYSTEM.UART_TX.c_clocks[0] ));
 sg13g2_dfrbp_1 _1241_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net220),
    .D(_0042_),
    .Q_N(_0663_),
    .Q(\MVM_UART_SYSTEM.UART_TX.c_clocks[1] ));
 sg13g2_dfrbp_1 _1242_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net220),
    .D(_0043_),
    .Q_N(_0662_),
    .Q(\MVM_UART_SYSTEM.UART_TX.c_clocks[2] ));
 sg13g2_dfrbp_1 _1243_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net220),
    .D(_0044_),
    .Q_N(_0661_),
    .Q(\MVM_UART_SYSTEM.UART_TX.c_clocks[3] ));
 sg13g2_dfrbp_1 _1244_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net219),
    .D(net281),
    .Q_N(_0660_),
    .Q(\MVM_UART_SYSTEM.UART_TX.c_clocks[4] ));
 sg13g2_dfrbp_1 _1245_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net219),
    .D(net246),
    .Q_N(_0659_),
    .Q(\MVM_UART_SYSTEM.UART_TX.c_clocks[5] ));
 sg13g2_dfrbp_1 _1246_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net219),
    .D(net267),
    .Q_N(_0658_),
    .Q(\MVM_UART_SYSTEM.UART_TX.c_clocks[6] ));
 sg13g2_dfrbp_1 _1247_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net220),
    .D(net102),
    .Q_N(_0657_),
    .Q(\MVM_UART_SYSTEM.UART_TX.c_clocks[7] ));
 sg13g2_dfrbp_1 _1248_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net219),
    .D(_0049_),
    .Q_N(_0656_),
    .Q(\MVM_UART_SYSTEM.UART_TX.c_clocks[8] ));
 sg13g2_dfrbp_1 _1249_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net219),
    .D(net160),
    .Q_N(_0655_),
    .Q(\MVM_UART_SYSTEM.UART_TX.c_clocks[9] ));
 sg13g2_dfrbp_1 _1250_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net219),
    .D(net115),
    .Q_N(_0654_),
    .Q(\MVM_UART_SYSTEM.UART_TX.c_clocks[10] ));
 sg13g2_dfrbp_1 _1251_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net215),
    .D(_0052_),
    .Q_N(_0668_),
    .Q(\MVM_UART_SYSTEM.UART_TX.c_clocks[11] ));
 sg13g2_dfrbp_1 _1252_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net208),
    .D(net64),
    .Q_N(_0653_),
    .Q(\MVM_UART_SYSTEM.AXIS_MVM.s_axis_kx_tvalid ));
 sg13g2_dfrbp_1 _1253_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net210),
    .D(net230),
    .Q_N(_0652_),
    .Q(\MVM_UART_SYSTEM.AXIS_MVM.SKID.buffer[0] ));
 sg13g2_dfrbp_1 _1254_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net209),
    .D(net164),
    .Q_N(_0651_),
    .Q(\MVM_UART_SYSTEM.AXIS_MVM.SKID.buffer[1] ));
 sg13g2_dfrbp_1 _1255_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net209),
    .D(net242),
    .Q_N(_0650_),
    .Q(\MVM_UART_SYSTEM.AXIS_MVM.SKID.buffer[2] ));
 sg13g2_dfrbp_1 _1256_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net209),
    .D(net143),
    .Q_N(_0649_),
    .Q(\MVM_UART_SYSTEM.AXIS_MVM.SKID.buffer[3] ));
 sg13g2_dfrbp_1 _1257_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net211),
    .D(net269),
    .Q_N(_0648_),
    .Q(\MVM_UART_SYSTEM.AXIS_MVM.SKID.buffer[4] ));
 sg13g2_dfrbp_1 _1258_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net209),
    .D(_0058_),
    .Q_N(_0647_),
    .Q(\MVM_UART_SYSTEM.AXIS_MVM.SKID.buffer[5] ));
 sg13g2_dfrbp_1 _1259_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net209),
    .D(_0059_),
    .Q_N(_0646_),
    .Q(\MVM_UART_SYSTEM.AXIS_MVM.SKID.buffer[6] ));
 sg13g2_dfrbp_1 _1260_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net210),
    .D(net223),
    .Q_N(_0645_),
    .Q(\MVM_UART_SYSTEM.AXIS_MVM.SKID.buffer[7] ));
 sg13g2_dfrbp_1 _1261_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net210),
    .D(net133),
    .Q_N(_0644_),
    .Q(\MVM_UART_SYSTEM.AXIS_MVM.SKID.buffer[8] ));
 sg13g2_dfrbp_1 _1262_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net210),
    .D(net119),
    .Q_N(_0643_),
    .Q(\MVM_UART_SYSTEM.AXIS_MVM.SKID.buffer[9] ));
 sg13g2_dfrbp_1 _1263_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net214),
    .D(net129),
    .Q_N(_0642_),
    .Q(\MVM_UART_SYSTEM.AXIS_MVM.SKID.buffer[10] ));
 sg13g2_dfrbp_1 _1264_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net214),
    .D(net234),
    .Q_N(_0641_),
    .Q(\MVM_UART_SYSTEM.AXIS_MVM.SKID.buffer[11] ));
 sg13g2_dfrbp_1 _1265_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net215),
    .D(_0065_),
    .Q_N(_0640_),
    .Q(\MVM_UART_SYSTEM.AXIS_MVM.SKID.buffer[12] ));
 sg13g2_dfrbp_1 _1266_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net214),
    .D(net131),
    .Q_N(_0639_),
    .Q(\MVM_UART_SYSTEM.AXIS_MVM.SKID.buffer[13] ));
 sg13g2_dfrbp_1 _1267_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net208),
    .D(_0067_),
    .Q_N(_0638_),
    .Q(\MVM_UART_SYSTEM.UART_RX.c_clocks[0] ));
 sg13g2_dfrbp_1 _1268_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net206),
    .D(net284),
    .Q_N(_0637_),
    .Q(\MVM_UART_SYSTEM.UART_RX.c_clocks[1] ));
 sg13g2_dfrbp_1 _1269_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net206),
    .D(_0069_),
    .Q_N(_0636_),
    .Q(\MVM_UART_SYSTEM.UART_RX.c_clocks[2] ));
 sg13g2_dfrbp_1 _1270_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net206),
    .D(net376),
    .Q_N(_0635_),
    .Q(\MVM_UART_SYSTEM.UART_RX.c_clocks[3] ));
 sg13g2_dfrbp_1 _1271_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net205),
    .D(net386),
    .Q_N(_0634_),
    .Q(\MVM_UART_SYSTEM.UART_RX.c_clocks[4] ));
 sg13g2_dfrbp_1 _1272_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net205),
    .D(net329),
    .Q_N(_0633_),
    .Q(\MVM_UART_SYSTEM.UART_RX.c_clocks[5] ));
 sg13g2_dfrbp_1 _1273_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net205),
    .D(_0073_),
    .Q_N(_0632_),
    .Q(\MVM_UART_SYSTEM.UART_RX.c_clocks[6] ));
 sg13g2_dfrbp_1 _1274_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net205),
    .D(net226),
    .Q_N(_0631_),
    .Q(\MVM_UART_SYSTEM.UART_RX.c_clocks[7] ));
 sg13g2_dfrbp_1 _1275_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net205),
    .D(_0075_),
    .Q_N(_0630_),
    .Q(\MVM_UART_SYSTEM.UART_RX.c_clocks[8] ));
 sg13g2_dfrbp_1 _1276_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net205),
    .D(net333),
    .Q_N(_0629_),
    .Q(\MVM_UART_SYSTEM.UART_RX.c_clocks[9] ));
 sg13g2_dfrbp_1 _1277_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net205),
    .D(net304),
    .Q_N(_0628_),
    .Q(\MVM_UART_SYSTEM.UART_RX.c_clocks[10] ));
 sg13g2_dfrbp_1 _1278_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net205),
    .D(net371),
    .Q_N(_0627_),
    .Q(\MVM_UART_SYSTEM.UART_RX.c_clocks[11] ));
 sg13g2_dfrbp_1 _1279_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net202),
    .D(_0079_),
    .Q_N(_0626_),
    .Q(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.x_pad[0][0] ));
 sg13g2_dfrbp_1 _1280_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net202),
    .D(_0080_),
    .Q_N(_0625_),
    .Q(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.x_pad[0][1] ));
 sg13g2_dfrbp_1 _1281_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net203),
    .D(net390),
    .Q_N(_0624_),
    .Q(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.x_pad[0][2] ));
 sg13g2_dfrbp_1 _1282_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net203),
    .D(net382),
    .Q_N(_0623_),
    .Q(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.x_pad[0][3] ));
 sg13g2_dfrbp_1 _1283_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net204),
    .D(_0083_),
    .Q_N(_0622_),
    .Q(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.x_pad[1][0] ));
 sg13g2_dfrbp_1 _1284_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net204),
    .D(net388),
    .Q_N(_0621_),
    .Q(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.x_pad[1][1] ));
 sg13g2_dfrbp_1 _1285_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net203),
    .D(net396),
    .Q_N(_0620_),
    .Q(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.x_pad[1][2] ));
 sg13g2_dfrbp_1 _1286_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net202),
    .D(net350),
    .Q_N(_0619_),
    .Q(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.x_pad[1][3] ));
 sg13g2_dfrbp_1 _1287_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net202),
    .D(_0087_),
    .Q_N(_0618_),
    .Q(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.k_pad[3][0] ));
 sg13g2_dfrbp_1 _1288_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net202),
    .D(_0088_),
    .Q_N(_0617_),
    .Q(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.k_pad[3][1] ));
 sg13g2_dfrbp_1 _1289_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net202),
    .D(_0089_),
    .Q_N(_0616_),
    .Q(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.k_pad[2][0] ));
 sg13g2_dfrbp_1 _1290_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net202),
    .D(_0090_),
    .Q_N(_0615_),
    .Q(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.k_pad[2][1] ));
 sg13g2_dfrbp_1 _1291_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net203),
    .D(_0091_),
    .Q_N(_0614_),
    .Q(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.k_pad[1][0] ));
 sg13g2_dfrbp_1 _1292_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net202),
    .D(_0092_),
    .Q_N(_0613_),
    .Q(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.k_pad[1][1] ));
 sg13g2_dfrbp_1 _1293_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net203),
    .D(net393),
    .Q_N(_0612_),
    .Q(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.k_pad[0][0] ));
 sg13g2_dfrbp_1 _1294_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net222),
    .D(_0094_),
    .Q_N(_0611_),
    .Q(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.k_pad[0][1] ));
 sg13g2_dfrbp_1 _1295_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net208),
    .D(net82),
    .Q_N(\MVM_UART_SYSTEM.UART_RX.state[0] ),
    .Q(_0010_));
 sg13g2_dfrbp_1 _1296_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net207),
    .D(net80),
    .Q_N(_0008_),
    .Q(\MVM_UART_SYSTEM.UART_RX.state[1] ));
 sg13g2_dfrbp_1 _1297_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net206),
    .D(_0001_),
    .Q_N(_0007_),
    .Q(\MVM_UART_SYSTEM.UART_RX.state[2] ));
 sg13g2_dfrbp_1 _1298_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net206),
    .D(net362),
    .Q_N(_0669_),
    .Q(\MVM_UART_SYSTEM.UART_RX.state[3] ));
 sg13g2_dfrbp_1 _1299_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net219),
    .D(net93),
    .Q_N(_0009_),
    .Q(\MVM_UART_SYSTEM.UART_TX.state ));
 sg13g2_dfrbp_1 _1300_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net215),
    .D(_0095_),
    .Q_N(_0610_),
    .Q(\MVM_UART_SYSTEM.UART_TX.c_pulses[0] ));
 sg13g2_dfrbp_1 _1301_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net215),
    .D(net289),
    .Q_N(_0609_),
    .Q(\MVM_UART_SYSTEM.UART_TX.c_pulses[1] ));
 sg13g2_dfrbp_1 _1302_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net215),
    .D(net316),
    .Q_N(_0608_),
    .Q(\MVM_UART_SYSTEM.UART_TX.c_pulses[2] ));
 sg13g2_dfrbp_1 _1303_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net208),
    .D(net107),
    .Q_N(_0607_),
    .Q(\MVM_UART_SYSTEM.UART_TX.c_pulses[3] ));
 sg13g2_dfrbp_1 _1304_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net208),
    .D(net262),
    .Q_N(_0606_),
    .Q(\MVM_UART_SYSTEM.UART_TX.c_pulses[4] ));
 sg13g2_dfrbp_1 _1305_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net215),
    .D(net104),
    .Q_N(\MVM_UART_SYSTEM.UART_TX.m_packets[0] ),
    .Q(_0011_));
 sg13g2_dfrbp_1 _1306_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net219),
    .D(net240),
    .Q_N(\MVM_UART_SYSTEM.UART_TX.m_packets[1] ),
    .Q(_0012_));
 sg13g2_dfrbp_1 _1307_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net213),
    .D(net248),
    .Q_N(\MVM_UART_SYSTEM.UART_TX.m_packets[2] ),
    .Q(_0013_));
 sg13g2_dfrbp_1 _1308_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net211),
    .D(net155),
    .Q_N(\MVM_UART_SYSTEM.UART_TX.m_packets[3] ),
    .Q(_0014_));
 sg13g2_dfrbp_1 _1309_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net211),
    .D(net264),
    .Q_N(\MVM_UART_SYSTEM.UART_TX.m_packets[4] ),
    .Q(_0015_));
 sg13g2_dfrbp_1 _1310_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net211),
    .D(net253),
    .Q_N(\MVM_UART_SYSTEM.UART_TX.m_packets[5] ),
    .Q(_0016_));
 sg13g2_dfrbp_1 _1311_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net212),
    .D(net228),
    .Q_N(\MVM_UART_SYSTEM.UART_TX.m_packets[6] ),
    .Q(_0017_));
 sg13g2_dfrbp_1 _1312_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net212),
    .D(net87),
    .Q_N(\MVM_UART_SYSTEM.UART_TX.m_packets[7] ),
    .Q(_0018_));
 sg13g2_dfrbp_1 _1313_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net212),
    .D(net95),
    .Q_N(\MVM_UART_SYSTEM.UART_TX.m_packets[8] ),
    .Q(_0019_));
 sg13g2_dfrbp_1 _1314_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net212),
    .D(net78),
    .Q_N(\MVM_UART_SYSTEM.UART_TX.m_packets[9] ),
    .Q(_0020_));
 sg13g2_dfrbp_1 _1315_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net218),
    .D(net72),
    .Q_N(\MVM_UART_SYSTEM.UART_TX.m_packets[10] ),
    .Q(_0021_));
 sg13g2_dfrbp_1 _1316_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net218),
    .D(net68),
    .Q_N(\MVM_UART_SYSTEM.UART_TX.m_packets[11] ),
    .Q(_0022_));
 sg13g2_dfrbp_1 _1317_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net218),
    .D(net76),
    .Q_N(\MVM_UART_SYSTEM.UART_TX.m_packets[12] ),
    .Q(_0023_));
 sg13g2_dfrbp_1 _1318_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net218),
    .D(net99),
    .Q_N(\MVM_UART_SYSTEM.UART_TX.m_packets[13] ),
    .Q(_0024_));
 sg13g2_dfrbp_1 _1319_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net217),
    .D(net157),
    .Q_N(\MVM_UART_SYSTEM.UART_TX.m_packets[14] ),
    .Q(_0025_));
 sg13g2_dfrbp_1 _1320_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net212),
    .D(net153),
    .Q_N(\MVM_UART_SYSTEM.UART_TX.m_packets[15] ),
    .Q(_0026_));
 sg13g2_dfrbp_1 _1321_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net212),
    .D(net141),
    .Q_N(\MVM_UART_SYSTEM.UART_TX.m_packets[16] ),
    .Q(_0027_));
 sg13g2_dfrbp_1 _1322_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net217),
    .D(net257),
    .Q_N(\MVM_UART_SYSTEM.UART_TX.m_packets[17] ),
    .Q(_0028_));
 sg13g2_dfrbp_1 _1323_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net214),
    .D(net255),
    .Q_N(\MVM_UART_SYSTEM.UART_TX.m_packets[18] ),
    .Q(_0029_));
 sg13g2_dfrbp_1 _1324_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net214),
    .D(net149),
    .Q_N(\MVM_UART_SYSTEM.UART_TX.m_packets[19] ),
    .Q(_0030_));
 sg13g2_dfrbp_1 _1325_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net217),
    .D(net91),
    .Q_N(\MVM_UART_SYSTEM.UART_TX.m_packets[20] ),
    .Q(_0031_));
 sg13g2_dfrbp_1 _1326_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net217),
    .D(net97),
    .Q_N(\MVM_UART_SYSTEM.UART_TX.m_packets[21] ),
    .Q(_0032_));
 sg13g2_dfrbp_1 _1327_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net217),
    .D(net70),
    .Q_N(\MVM_UART_SYSTEM.UART_TX.m_packets[22] ),
    .Q(_0033_));
 sg13g2_dfrbp_1 _1328_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net217),
    .D(net74),
    .Q_N(\MVM_UART_SYSTEM.UART_TX.m_packets[23] ),
    .Q(_0034_));
 sg13g2_dfrbp_1 _1329_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net217),
    .D(net66),
    .Q_N(\MVM_UART_SYSTEM.UART_TX.m_packets[24] ),
    .Q(_0035_));
 sg13g2_dfrbp_1 _1330_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net217),
    .D(net85),
    .Q_N(\MVM_UART_SYSTEM.UART_TX.m_packets[25] ),
    .Q(_0036_));
 sg13g2_dfrbp_1 _1331_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net207),
    .D(net89),
    .Q_N(_0006_),
    .Q(\MVM_UART_SYSTEM.UART_RX.c_words ));
 sg13g2_dfrbp_1 _1332_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net208),
    .D(net232),
    .Q_N(_0605_),
    .Q(\MVM_UART_SYSTEM.AXIS_MVM.shift ));
 sg13g2_dfrbp_1 _1333_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net52),
    .D(net357),
    .Q_N(_0604_),
    .Q(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[1][0] ));
 sg13g2_dfrbp_1 _1334_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net51),
    .D(_0129_),
    .Q_N(_0603_),
    .Q(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[1][1] ));
 sg13g2_dfrbp_1 _1335_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net50),
    .D(net310),
    .Q_N(_0602_),
    .Q(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[1][2] ));
 sg13g2_dfrbp_1 _1336_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net49),
    .D(net352),
    .Q_N(_0601_),
    .Q(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[1][3] ));
 sg13g2_dfrbp_1 _1337_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net48),
    .D(_0132_),
    .Q_N(_0600_),
    .Q(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[1][4] ));
 sg13g2_dfrbp_1 _1338_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net47),
    .D(net298),
    .Q_N(_0599_),
    .Q(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[1][5] ));
 sg13g2_dfrbp_1 _1339_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net46),
    .D(net259),
    .Q_N(_0598_),
    .Q(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[2][0] ));
 sg13g2_dfrbp_1 _1340_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net45),
    .D(net277),
    .Q_N(_0597_),
    .Q(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[2][1] ));
 sg13g2_dfrbp_1 _1341_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net44),
    .D(_0136_),
    .Q_N(_0596_),
    .Q(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[2][2] ));
 sg13g2_dfrbp_1 _1342_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net43),
    .D(net300),
    .Q_N(_0595_),
    .Q(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[2][3] ));
 sg13g2_dfrbp_1 _1343_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net42),
    .D(net296),
    .Q_N(_0594_),
    .Q(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[2][4] ));
 sg13g2_dfrbp_1 _1344_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net41),
    .D(net111),
    .Q_N(_0593_),
    .Q(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[2][5] ));
 sg13g2_dfrbp_1 _1345_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net40),
    .D(net236),
    .Q_N(_0592_),
    .Q(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[2][6] ));
 sg13g2_dfrbp_1 _1346_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net39),
    .D(net319),
    .Q_N(_0591_),
    .Q(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[4][0] ));
 sg13g2_dfrbp_1 _1347_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net38),
    .D(net337),
    .Q_N(_0590_),
    .Q(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[4][1] ));
 sg13g2_dfrbp_1 _1348_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net37),
    .D(net355),
    .Q_N(_0589_),
    .Q(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[4][2] ));
 sg13g2_dfrbp_1 _1349_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net36),
    .D(_0144_),
    .Q_N(_0588_),
    .Q(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[4][3] ));
 sg13g2_dfrbp_1 _1350_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net35),
    .D(_0145_),
    .Q_N(_0587_),
    .Q(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[4][4] ));
 sg13g2_dfrbp_1 _1351_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net34),
    .D(net294),
    .Q_N(_0586_),
    .Q(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[4][5] ));
 sg13g2_dfrbp_1 _1352_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net33),
    .D(net346),
    .Q_N(_0585_),
    .Q(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[5][0] ));
 sg13g2_dfrbp_1 _1353_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net32),
    .D(net326),
    .Q_N(_0584_),
    .Q(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[5][1] ));
 sg13g2_dfrbp_1 _1354_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net31),
    .D(net324),
    .Q_N(_0583_),
    .Q(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[5][2] ));
 sg13g2_dfrbp_1 _1355_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net30),
    .D(_0150_),
    .Q_N(_0582_),
    .Q(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[5][3] ));
 sg13g2_dfrbp_1 _1356_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net29),
    .D(_0151_),
    .Q_N(_0581_),
    .Q(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[5][4] ));
 sg13g2_dfrbp_1 _1357_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net28),
    .D(net308),
    .Q_N(_0580_),
    .Q(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[5][5] ));
 sg13g2_dfrbp_1 _1358_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net27),
    .D(net275),
    .Q_N(_0579_),
    .Q(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[6][0] ));
 sg13g2_dfrbp_1 _1359_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net26),
    .D(net302),
    .Q_N(_0578_),
    .Q(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[6][1] ));
 sg13g2_dfrbp_1 _1360_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net25),
    .D(net272),
    .Q_N(_0577_),
    .Q(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[6][2] ));
 sg13g2_dfrbp_1 _1361_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net61),
    .D(net162),
    .Q_N(_0576_),
    .Q(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[6][3] ));
 sg13g2_dfrbp_1 _1362_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net60),
    .D(net251),
    .Q_N(_0575_),
    .Q(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[6][4] ));
 sg13g2_dfrbp_1 _1363_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net59),
    .D(net238),
    .Q_N(_0574_),
    .Q(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[6][5] ));
 sg13g2_dfrbp_1 _1364_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net58),
    .D(net139),
    .Q_N(_0573_),
    .Q(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[6][6] ));
 sg13g2_dfrbp_1 _1365_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net208),
    .D(net292),
    .Q_N(_0572_),
    .Q(\MVM_UART_SYSTEM.AXIS_MVM.SKID.s_valid ));
 sg13g2_dfrbp_1 _1366_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net57),
    .D(net312),
    .Q_N(_0571_),
    .Q(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[0][0] ));
 sg13g2_dfrbp_1 _1367_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net56),
    .D(net341),
    .Q_N(_0570_),
    .Q(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[0][1] ));
 sg13g2_dfrbp_1 _1368_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net55),
    .D(net364),
    .Q_N(_0569_),
    .Q(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[0][2] ));
 sg13g2_dfrbp_1 _1369_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net54),
    .D(_0164_),
    .Q_N(_0568_),
    .Q(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[0][3] ));
 sg13g2_dfrbp_1 _1370_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net53),
    .D(_0165_),
    .Q_N(_0567_),
    .Q(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[0][4] ));
 sg13g2_dfrbp_1 _1371_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net62),
    .D(net314),
    .Q_N(_0670_),
    .Q(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[0][5] ));
 sg13g2_dfrbp_1 _1372_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net215),
    .D(_0003_),
    .Q_N(_0566_),
    .Q(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.cen ));
 sg13g2_dfrbp_1 _1373_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net210),
    .D(net109),
    .Q_N(_0565_),
    .Q(\MVM_UART_SYSTEM.AXIS_MVM.SKID.m_data[0] ));
 sg13g2_dfrbp_1 _1374_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net209),
    .D(net123),
    .Q_N(_0564_),
    .Q(\MVM_UART_SYSTEM.AXIS_MVM.SKID.m_data[1] ));
 sg13g2_dfrbp_1 _1375_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net209),
    .D(net137),
    .Q_N(_0563_),
    .Q(\MVM_UART_SYSTEM.AXIS_MVM.SKID.m_data[2] ));
 sg13g2_dfrbp_1 _1376_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net211),
    .D(net279),
    .Q_N(_0562_),
    .Q(\MVM_UART_SYSTEM.AXIS_MVM.SKID.m_data[3] ));
 sg13g2_dfrbp_1 _1377_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net211),
    .D(net286),
    .Q_N(_0561_),
    .Q(\MVM_UART_SYSTEM.AXIS_MVM.SKID.m_data[4] ));
 sg13g2_dfrbp_1 _1378_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net211),
    .D(net127),
    .Q_N(_0560_),
    .Q(\MVM_UART_SYSTEM.AXIS_MVM.SKID.m_data[5] ));
 sg13g2_dfrbp_1 _1379_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net211),
    .D(net145),
    .Q_N(_0559_),
    .Q(\MVM_UART_SYSTEM.AXIS_MVM.SKID.m_data[6] ));
 sg13g2_dfrbp_1 _1380_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net213),
    .D(net147),
    .Q_N(_0558_),
    .Q(\MVM_UART_SYSTEM.AXIS_MVM.SKID.m_data[7] ));
 sg13g2_dfrbp_1 _1381_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net212),
    .D(net113),
    .Q_N(_0557_),
    .Q(\MVM_UART_SYSTEM.AXIS_MVM.SKID.m_data[8] ));
 sg13g2_dfrbp_1 _1382_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net209),
    .D(net135),
    .Q_N(_0556_),
    .Q(\MVM_UART_SYSTEM.AXIS_MVM.SKID.m_data[9] ));
 sg13g2_dfrbp_1 _1383_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net214),
    .D(net121),
    .Q_N(_0555_),
    .Q(\MVM_UART_SYSTEM.AXIS_MVM.SKID.m_data[10] ));
 sg13g2_dfrbp_1 _1384_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net216),
    .D(net125),
    .Q_N(_0554_),
    .Q(\MVM_UART_SYSTEM.AXIS_MVM.SKID.m_data[11] ));
 sg13g2_dfrbp_1 _1385_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net214),
    .D(net117),
    .Q_N(_0553_),
    .Q(\MVM_UART_SYSTEM.AXIS_MVM.SKID.m_data[12] ));
 sg13g2_dfrbp_1 _1386_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net214),
    .D(_0180_),
    .Q_N(_0671_),
    .Q(\MVM_UART_SYSTEM.AXIS_MVM.SKID.m_data[13] ));
 sg13g2_dfrbp_1 _1387_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net215),
    .D(_0004_),
    .Q_N(_0672_),
    .Q(\MVM_UART_SYSTEM.AXIS_MVM.SKID.m_valid ));
 sg13g2_dfrbp_1 _1388_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net216),
    .D(\MVM_UART_SYSTEM.AXIS_MVM.SKID.state_next[0] ),
    .Q_N(_0673_),
    .Q(\MVM_UART_SYSTEM.AXIS_MVM.SKID.state[0] ));
 sg13g2_dfrbp_1 _1389_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net216),
    .D(\MVM_UART_SYSTEM.AXIS_MVM.SKID.state_next[1] ),
    .Q_N(_0552_),
    .Q(\MVM_UART_SYSTEM.AXIS_MVM.SKID.state[1] ));
 sg13g2_tiehi _1359__26 (.L_HI(net26));
 sg13g2_tiehi _1358__27 (.L_HI(net27));
 sg13g2_tiehi _1357__28 (.L_HI(net28));
 sg13g2_tiehi _1356__29 (.L_HI(net29));
 sg13g2_tiehi _1355__30 (.L_HI(net30));
 sg13g2_tiehi _1354__31 (.L_HI(net31));
 sg13g2_tiehi _1353__32 (.L_HI(net32));
 sg13g2_tiehi _1352__33 (.L_HI(net33));
 sg13g2_tiehi _1351__34 (.L_HI(net34));
 sg13g2_tiehi _1350__35 (.L_HI(net35));
 sg13g2_tiehi _1349__36 (.L_HI(net36));
 sg13g2_tiehi _1348__37 (.L_HI(net37));
 sg13g2_tiehi _1347__38 (.L_HI(net38));
 sg13g2_tiehi _1346__39 (.L_HI(net39));
 sg13g2_tiehi _1345__40 (.L_HI(net40));
 sg13g2_tiehi _1344__41 (.L_HI(net41));
 sg13g2_tiehi _1343__42 (.L_HI(net42));
 sg13g2_tiehi _1342__43 (.L_HI(net43));
 sg13g2_tiehi _1341__44 (.L_HI(net44));
 sg13g2_tiehi _1340__45 (.L_HI(net45));
 sg13g2_tiehi _1339__46 (.L_HI(net46));
 sg13g2_tiehi _1338__47 (.L_HI(net47));
 sg13g2_tiehi _1337__48 (.L_HI(net48));
 sg13g2_tiehi _1336__49 (.L_HI(net49));
 sg13g2_tiehi _1335__50 (.L_HI(net50));
 sg13g2_tiehi _1334__51 (.L_HI(net51));
 sg13g2_tiehi _1333__52 (.L_HI(net52));
 sg13g2_tiehi _1370__53 (.L_HI(net53));
 sg13g2_tiehi _1369__54 (.L_HI(net54));
 sg13g2_tiehi _1368__55 (.L_HI(net55));
 sg13g2_tiehi _1367__56 (.L_HI(net56));
 sg13g2_tiehi _1366__57 (.L_HI(net57));
 sg13g2_tiehi _1364__58 (.L_HI(net58));
 sg13g2_tiehi _1363__59 (.L_HI(net59));
 sg13g2_tiehi _1362__60 (.L_HI(net60));
 sg13g2_tiehi _1361__61 (.L_HI(net61));
 sg13g2_tiehi _1371__62 (.L_HI(net62));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_uart_mvm_sys_3 (.L_LO(net3));
 sg13g2_tielo tt_um_uart_mvm_sys_4 (.L_LO(net4));
 sg13g2_tielo tt_um_uart_mvm_sys_5 (.L_LO(net5));
 sg13g2_tielo tt_um_uart_mvm_sys_6 (.L_LO(net6));
 sg13g2_tielo tt_um_uart_mvm_sys_7 (.L_LO(net7));
 sg13g2_tielo tt_um_uart_mvm_sys_8 (.L_LO(net8));
 sg13g2_tielo tt_um_uart_mvm_sys_9 (.L_LO(net9));
 sg13g2_tielo tt_um_uart_mvm_sys_10 (.L_LO(net10));
 sg13g2_tielo tt_um_uart_mvm_sys_11 (.L_LO(net11));
 sg13g2_tielo tt_um_uart_mvm_sys_12 (.L_LO(net12));
 sg13g2_tielo tt_um_uart_mvm_sys_13 (.L_LO(net13));
 sg13g2_tielo tt_um_uart_mvm_sys_14 (.L_LO(net14));
 sg13g2_tielo tt_um_uart_mvm_sys_15 (.L_LO(net15));
 sg13g2_tielo tt_um_uart_mvm_sys_16 (.L_LO(net16));
 sg13g2_tielo tt_um_uart_mvm_sys_17 (.L_LO(net17));
 sg13g2_tielo tt_um_uart_mvm_sys_18 (.L_LO(net18));
 sg13g2_tielo tt_um_uart_mvm_sys_19 (.L_LO(net19));
 sg13g2_tielo tt_um_uart_mvm_sys_20 (.L_LO(net20));
 sg13g2_tielo tt_um_uart_mvm_sys_21 (.L_LO(net21));
 sg13g2_tielo tt_um_uart_mvm_sys_22 (.L_LO(net22));
 sg13g2_tielo tt_um_uart_mvm_sys_23 (.L_LO(net23));
 sg13g2_tielo tt_um_uart_mvm_sys_24 (.L_LO(net24));
 sg13g2_tiehi _1360__25 (.L_HI(net25));
 sg13g2_buf_1 _1451_ (.A(\MVM_UART_SYSTEM.UART_TX.m_packets[0] ),
    .X(uo_out[0]));
 sg13g2_buf_4 fanout166 (.X(net166),
    .A(_0537_));
 sg13g2_buf_2 fanout167 (.A(_0537_),
    .X(net167));
 sg13g2_buf_4 fanout168 (.X(net168),
    .A(net172));
 sg13g2_buf_2 fanout169 (.A(net172),
    .X(net169));
 sg13g2_buf_2 fanout170 (.A(net171),
    .X(net170));
 sg13g2_buf_2 fanout171 (.A(net172),
    .X(net171));
 sg13g2_buf_2 fanout172 (.A(_0317_),
    .X(net172));
 sg13g2_buf_4 fanout173 (.X(net173),
    .A(net175));
 sg13g2_buf_2 fanout174 (.A(net175),
    .X(net174));
 sg13g2_buf_4 fanout175 (.X(net175),
    .A(_0244_));
 sg13g2_buf_2 fanout176 (.A(_0319_),
    .X(net176));
 sg13g2_buf_2 fanout177 (.A(_0319_),
    .X(net177));
 sg13g2_buf_2 fanout178 (.A(_0241_),
    .X(net178));
 sg13g2_buf_2 fanout179 (.A(_0275_),
    .X(net179));
 sg13g2_buf_1 fanout180 (.A(_0275_),
    .X(net180));
 sg13g2_buf_4 fanout181 (.X(net181),
    .A(net183));
 sg13g2_buf_4 fanout182 (.X(net182),
    .A(net183));
 sg13g2_buf_2 fanout183 (.A(_0225_),
    .X(net183));
 sg13g2_buf_4 fanout184 (.X(net184),
    .A(_0228_));
 sg13g2_buf_2 fanout185 (.A(_0228_),
    .X(net185));
 sg13g2_buf_2 fanout186 (.A(net188),
    .X(net186));
 sg13g2_buf_2 fanout187 (.A(net188),
    .X(net187));
 sg13g2_buf_2 fanout188 (.A(net191),
    .X(net188));
 sg13g2_buf_2 fanout189 (.A(net191),
    .X(net189));
 sg13g2_buf_2 fanout190 (.A(net191),
    .X(net190));
 sg13g2_buf_1 fanout191 (.A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.cen ),
    .X(net191));
 sg13g2_buf_2 fanout192 (.A(net195),
    .X(net192));
 sg13g2_buf_2 fanout193 (.A(net195),
    .X(net193));
 sg13g2_buf_1 fanout194 (.A(net195),
    .X(net194));
 sg13g2_buf_2 fanout195 (.A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.cen ),
    .X(net195));
 sg13g2_buf_2 fanout196 (.A(net197),
    .X(net196));
 sg13g2_buf_2 fanout197 (.A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.cen ),
    .X(net197));
 sg13g2_buf_2 fanout198 (.A(net201),
    .X(net198));
 sg13g2_buf_2 fanout199 (.A(net201),
    .X(net199));
 sg13g2_buf_2 fanout200 (.A(net201),
    .X(net200));
 sg13g2_buf_2 fanout201 (.A(\MVM_UART_SYSTEM.UART_TX.state ),
    .X(net201));
 sg13g2_buf_4 fanout202 (.X(net202),
    .A(net204));
 sg13g2_buf_2 fanout203 (.A(net204),
    .X(net203));
 sg13g2_buf_2 fanout204 (.A(net222),
    .X(net204));
 sg13g2_buf_4 fanout205 (.X(net205),
    .A(net207));
 sg13g2_buf_2 fanout206 (.A(net207),
    .X(net206));
 sg13g2_buf_4 fanout207 (.X(net207),
    .A(net208));
 sg13g2_buf_4 fanout208 (.X(net208),
    .A(net222));
 sg13g2_buf_4 fanout209 (.X(net209),
    .A(net213));
 sg13g2_buf_2 fanout210 (.A(net213),
    .X(net210));
 sg13g2_buf_4 fanout211 (.X(net211),
    .A(net212));
 sg13g2_buf_4 fanout212 (.X(net212),
    .A(net213));
 sg13g2_buf_2 fanout213 (.A(net222),
    .X(net213));
 sg13g2_buf_4 fanout214 (.X(net214),
    .A(net216));
 sg13g2_buf_4 fanout215 (.X(net215),
    .A(net216));
 sg13g2_buf_2 fanout216 (.A(net222),
    .X(net216));
 sg13g2_buf_4 fanout217 (.X(net217),
    .A(net221));
 sg13g2_buf_2 fanout218 (.A(net221),
    .X(net218));
 sg13g2_buf_4 fanout219 (.X(net219),
    .A(net221));
 sg13g2_buf_2 fanout220 (.A(net221),
    .X(net220));
 sg13g2_buf_1 fanout221 (.A(net222),
    .X(net221));
 sg13g2_buf_4 fanout222 (.X(net222),
    .A(rst_n));
 sg13g2_buf_2 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_tielo tt_um_uart_mvm_sys_2 (.L_LO(net2));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_buf_2 clkbuf_5_0__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_0__leaf_clk));
 sg13g2_buf_2 clkbuf_5_1__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_1__leaf_clk));
 sg13g2_buf_2 clkbuf_5_2__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_2__leaf_clk));
 sg13g2_buf_2 clkbuf_5_3__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_3__leaf_clk));
 sg13g2_buf_2 clkbuf_5_4__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_4__leaf_clk));
 sg13g2_buf_2 clkbuf_5_5__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_5__leaf_clk));
 sg13g2_buf_2 clkbuf_5_6__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_6__leaf_clk));
 sg13g2_buf_2 clkbuf_5_7__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_7__leaf_clk));
 sg13g2_buf_2 clkbuf_5_8__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_8__leaf_clk));
 sg13g2_buf_2 clkbuf_5_9__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_9__leaf_clk));
 sg13g2_buf_2 clkbuf_5_10__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_10__leaf_clk));
 sg13g2_buf_2 clkbuf_5_11__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_11__leaf_clk));
 sg13g2_buf_2 clkbuf_5_12__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_12__leaf_clk));
 sg13g2_buf_2 clkbuf_5_13__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_13__leaf_clk));
 sg13g2_buf_2 clkbuf_5_14__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_14__leaf_clk));
 sg13g2_buf_2 clkbuf_5_15__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_15__leaf_clk));
 sg13g2_buf_2 clkbuf_5_16__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_16__leaf_clk));
 sg13g2_buf_2 clkbuf_5_17__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_17__leaf_clk));
 sg13g2_buf_2 clkbuf_5_18__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_18__leaf_clk));
 sg13g2_buf_2 clkbuf_5_19__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_19__leaf_clk));
 sg13g2_buf_2 clkbuf_5_20__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_20__leaf_clk));
 sg13g2_buf_2 clkbuf_5_21__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_21__leaf_clk));
 sg13g2_buf_2 clkbuf_5_22__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_22__leaf_clk));
 sg13g2_buf_2 clkbuf_5_23__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_23__leaf_clk));
 sg13g2_buf_2 clkbuf_5_24__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_24__leaf_clk));
 sg13g2_buf_2 clkbuf_5_25__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_25__leaf_clk));
 sg13g2_buf_2 clkbuf_5_26__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_26__leaf_clk));
 sg13g2_buf_2 clkbuf_5_27__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_27__leaf_clk));
 sg13g2_buf_2 clkbuf_5_28__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_28__leaf_clk));
 sg13g2_buf_2 clkbuf_5_29__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_29__leaf_clk));
 sg13g2_buf_2 clkbuf_5_30__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_30__leaf_clk));
 sg13g2_buf_2 clkbuf_5_31__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_31__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_5_7__leaf_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_5_11__leaf_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_5_15__leaf_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_5_19__leaf_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_5_23__leaf_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_5_27__leaf_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_5_31__leaf_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(_0006_),
    .X(net63));
 sg13g2_dlygate4sd3_1 hold2 (.A(_0005_),
    .X(net64));
 sg13g2_dlygate4sd3_1 hold3 (.A(\MVM_UART_SYSTEM.UART_TX.m_packets[25] ),
    .X(net65));
 sg13g2_dlygate4sd3_1 hold4 (.A(_0124_),
    .X(net66));
 sg13g2_dlygate4sd3_1 hold5 (.A(\MVM_UART_SYSTEM.UART_TX.m_packets[12] ),
    .X(net67));
 sg13g2_dlygate4sd3_1 hold6 (.A(_0111_),
    .X(net68));
 sg13g2_dlygate4sd3_1 hold7 (.A(\MVM_UART_SYSTEM.UART_TX.m_packets[23] ),
    .X(net69));
 sg13g2_dlygate4sd3_1 hold8 (.A(_0122_),
    .X(net70));
 sg13g2_dlygate4sd3_1 hold9 (.A(\MVM_UART_SYSTEM.UART_TX.m_packets[11] ),
    .X(net71));
 sg13g2_dlygate4sd3_1 hold10 (.A(_0110_),
    .X(net72));
 sg13g2_dlygate4sd3_1 hold11 (.A(\MVM_UART_SYSTEM.UART_TX.m_packets[24] ),
    .X(net73));
 sg13g2_dlygate4sd3_1 hold12 (.A(_0123_),
    .X(net74));
 sg13g2_dlygate4sd3_1 hold13 (.A(\MVM_UART_SYSTEM.UART_TX.m_packets[13] ),
    .X(net75));
 sg13g2_dlygate4sd3_1 hold14 (.A(_0112_),
    .X(net76));
 sg13g2_dlygate4sd3_1 hold15 (.A(\MVM_UART_SYSTEM.UART_TX.m_packets[10] ),
    .X(net77));
 sg13g2_dlygate4sd3_1 hold16 (.A(_0109_),
    .X(net78));
 sg13g2_dlygate4sd3_1 hold17 (.A(_0008_),
    .X(net79));
 sg13g2_dlygate4sd3_1 hold18 (.A(_0000_),
    .X(net80));
 sg13g2_dlygate4sd3_1 hold19 (.A(\MVM_UART_SYSTEM.UART_RX.state[0] ),
    .X(net81));
 sg13g2_dlygate4sd3_1 hold20 (.A(_0037_),
    .X(net82));
 sg13g2_dlygate4sd3_1 hold21 (.A(_0007_),
    .X(net83));
 sg13g2_dlygate4sd3_1 hold22 (.A(_0036_),
    .X(net84));
 sg13g2_dlygate4sd3_1 hold23 (.A(_0125_),
    .X(net85));
 sg13g2_dlygate4sd3_1 hold24 (.A(\MVM_UART_SYSTEM.UART_TX.m_packets[8] ),
    .X(net86));
 sg13g2_dlygate4sd3_1 hold25 (.A(_0107_),
    .X(net87));
 sg13g2_dlygate4sd3_1 hold26 (.A(\MVM_UART_SYSTEM.UART_RX.c_words ),
    .X(net88));
 sg13g2_dlygate4sd3_1 hold27 (.A(_0126_),
    .X(net89));
 sg13g2_dlygate4sd3_1 hold28 (.A(\MVM_UART_SYSTEM.UART_TX.m_packets[21] ),
    .X(net90));
 sg13g2_dlygate4sd3_1 hold29 (.A(_0120_),
    .X(net91));
 sg13g2_dlygate4sd3_1 hold30 (.A(\MVM_UART_SYSTEM.AXIS_MVM.SKID.m_valid ),
    .X(net92));
 sg13g2_dlygate4sd3_1 hold31 (.A(_0712_),
    .X(net93));
 sg13g2_dlygate4sd3_1 hold32 (.A(\MVM_UART_SYSTEM.UART_TX.m_packets[9] ),
    .X(net94));
 sg13g2_dlygate4sd3_1 hold33 (.A(_0108_),
    .X(net95));
 sg13g2_dlygate4sd3_1 hold34 (.A(\MVM_UART_SYSTEM.UART_TX.m_packets[22] ),
    .X(net96));
 sg13g2_dlygate4sd3_1 hold35 (.A(_0121_),
    .X(net97));
 sg13g2_dlygate4sd3_1 hold36 (.A(\MVM_UART_SYSTEM.UART_TX.m_packets[14] ),
    .X(net98));
 sg13g2_dlygate4sd3_1 hold37 (.A(_0113_),
    .X(net99));
 sg13g2_dlygate4sd3_1 hold38 (.A(\MVM_UART_SYSTEM.UART_TX.c_clocks[7] ),
    .X(net100));
 sg13g2_dlygate4sd3_1 hold39 (.A(_0265_),
    .X(net101));
 sg13g2_dlygate4sd3_1 hold40 (.A(_0048_),
    .X(net102));
 sg13g2_dlygate4sd3_1 hold41 (.A(\MVM_UART_SYSTEM.UART_TX.m_packets[1] ),
    .X(net103));
 sg13g2_dlygate4sd3_1 hold42 (.A(_0100_),
    .X(net104));
 sg13g2_dlygate4sd3_1 hold43 (.A(\MVM_UART_SYSTEM.UART_TX.c_pulses[3] ),
    .X(net105));
 sg13g2_dlygate4sd3_1 hold44 (.A(_0313_),
    .X(net106));
 sg13g2_dlygate4sd3_1 hold45 (.A(_0098_),
    .X(net107));
 sg13g2_dlygate4sd3_1 hold46 (.A(\MVM_UART_SYSTEM.AXIS_MVM.SKID.m_data[0] ),
    .X(net108));
 sg13g2_dlygate4sd3_1 hold47 (.A(_0167_),
    .X(net109));
 sg13g2_dlygate4sd3_1 hold48 (.A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[2][5] ),
    .X(net110));
 sg13g2_dlygate4sd3_1 hold49 (.A(_0139_),
    .X(net111));
 sg13g2_dlygate4sd3_1 hold50 (.A(\MVM_UART_SYSTEM.AXIS_MVM.SKID.m_data[8] ),
    .X(net112));
 sg13g2_dlygate4sd3_1 hold51 (.A(_0175_),
    .X(net113));
 sg13g2_dlygate4sd3_1 hold52 (.A(\MVM_UART_SYSTEM.UART_TX.c_clocks[10] ),
    .X(net114));
 sg13g2_dlygate4sd3_1 hold53 (.A(_0051_),
    .X(net115));
 sg13g2_dlygate4sd3_1 hold54 (.A(\MVM_UART_SYSTEM.AXIS_MVM.SKID.m_data[12] ),
    .X(net116));
 sg13g2_dlygate4sd3_1 hold55 (.A(_0179_),
    .X(net117));
 sg13g2_dlygate4sd3_1 hold56 (.A(\MVM_UART_SYSTEM.AXIS_MVM.SKID.buffer[9] ),
    .X(net118));
 sg13g2_dlygate4sd3_1 hold57 (.A(_0062_),
    .X(net119));
 sg13g2_dlygate4sd3_1 hold58 (.A(\MVM_UART_SYSTEM.AXIS_MVM.SKID.m_data[10] ),
    .X(net120));
 sg13g2_dlygate4sd3_1 hold59 (.A(_0177_),
    .X(net121));
 sg13g2_dlygate4sd3_1 hold60 (.A(\MVM_UART_SYSTEM.AXIS_MVM.SKID.m_data[1] ),
    .X(net122));
 sg13g2_dlygate4sd3_1 hold61 (.A(_0168_),
    .X(net123));
 sg13g2_dlygate4sd3_1 hold62 (.A(\MVM_UART_SYSTEM.AXIS_MVM.SKID.m_data[11] ),
    .X(net124));
 sg13g2_dlygate4sd3_1 hold63 (.A(_0178_),
    .X(net125));
 sg13g2_dlygate4sd3_1 hold64 (.A(\MVM_UART_SYSTEM.AXIS_MVM.SKID.m_data[5] ),
    .X(net126));
 sg13g2_dlygate4sd3_1 hold65 (.A(_0172_),
    .X(net127));
 sg13g2_dlygate4sd3_1 hold66 (.A(\MVM_UART_SYSTEM.AXIS_MVM.SKID.buffer[10] ),
    .X(net128));
 sg13g2_dlygate4sd3_1 hold67 (.A(_0063_),
    .X(net129));
 sg13g2_dlygate4sd3_1 hold68 (.A(\MVM_UART_SYSTEM.AXIS_MVM.SKID.buffer[13] ),
    .X(net130));
 sg13g2_dlygate4sd3_1 hold69 (.A(_0066_),
    .X(net131));
 sg13g2_dlygate4sd3_1 hold70 (.A(\MVM_UART_SYSTEM.AXIS_MVM.SKID.buffer[8] ),
    .X(net132));
 sg13g2_dlygate4sd3_1 hold71 (.A(_0061_),
    .X(net133));
 sg13g2_dlygate4sd3_1 hold72 (.A(\MVM_UART_SYSTEM.AXIS_MVM.SKID.m_data[9] ),
    .X(net134));
 sg13g2_dlygate4sd3_1 hold73 (.A(_0176_),
    .X(net135));
 sg13g2_dlygate4sd3_1 hold74 (.A(\MVM_UART_SYSTEM.AXIS_MVM.SKID.m_data[2] ),
    .X(net136));
 sg13g2_dlygate4sd3_1 hold75 (.A(_0169_),
    .X(net137));
 sg13g2_dlygate4sd3_1 hold76 (.A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[6][6] ),
    .X(net138));
 sg13g2_dlygate4sd3_1 hold77 (.A(_0159_),
    .X(net139));
 sg13g2_dlygate4sd3_1 hold78 (.A(_0027_),
    .X(net140));
 sg13g2_dlygate4sd3_1 hold79 (.A(_0116_),
    .X(net141));
 sg13g2_dlygate4sd3_1 hold80 (.A(\MVM_UART_SYSTEM.AXIS_MVM.SKID.buffer[3] ),
    .X(net142));
 sg13g2_dlygate4sd3_1 hold81 (.A(_0056_),
    .X(net143));
 sg13g2_dlygate4sd3_1 hold82 (.A(\MVM_UART_SYSTEM.AXIS_MVM.SKID.m_data[6] ),
    .X(net144));
 sg13g2_dlygate4sd3_1 hold83 (.A(_0173_),
    .X(net145));
 sg13g2_dlygate4sd3_1 hold84 (.A(\MVM_UART_SYSTEM.AXIS_MVM.SKID.m_data[7] ),
    .X(net146));
 sg13g2_dlygate4sd3_1 hold85 (.A(_0174_),
    .X(net147));
 sg13g2_dlygate4sd3_1 hold86 (.A(_0030_),
    .X(net148));
 sg13g2_dlygate4sd3_1 hold87 (.A(_0119_),
    .X(net149));
 sg13g2_dlygate4sd3_1 hold88 (.A(\MVM_UART_SYSTEM.UART_RX.c_bits[2] ),
    .X(net150));
 sg13g2_dlygate4sd3_1 hold89 (.A(_0040_),
    .X(net151));
 sg13g2_dlygate4sd3_1 hold90 (.A(_0026_),
    .X(net152));
 sg13g2_dlygate4sd3_1 hold91 (.A(_0115_),
    .X(net153));
 sg13g2_dlygate4sd3_1 hold92 (.A(_0014_),
    .X(net154));
 sg13g2_dlygate4sd3_1 hold93 (.A(_0103_),
    .X(net155));
 sg13g2_dlygate4sd3_1 hold94 (.A(_0025_),
    .X(net156));
 sg13g2_dlygate4sd3_1 hold95 (.A(_0114_),
    .X(net157));
 sg13g2_dlygate4sd3_1 hold96 (.A(\MVM_UART_SYSTEM.UART_TX.c_clocks[9] ),
    .X(net158));
 sg13g2_dlygate4sd3_1 hold97 (.A(_0266_),
    .X(net159));
 sg13g2_dlygate4sd3_1 hold98 (.A(_0050_),
    .X(net160));
 sg13g2_dlygate4sd3_1 hold99 (.A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[6][3] ),
    .X(net161));
 sg13g2_dlygate4sd3_1 hold100 (.A(_0156_),
    .X(net162));
 sg13g2_dlygate4sd3_1 hold101 (.A(\MVM_UART_SYSTEM.AXIS_MVM.SKID.buffer[1] ),
    .X(net163));
 sg13g2_dlygate4sd3_1 hold102 (.A(_0054_),
    .X(net164));
 sg13g2_dlygate4sd3_1 hold103 (.A(\MVM_UART_SYSTEM.AXIS_MVM.SKID.buffer[7] ),
    .X(net165));
 sg13g2_dlygate4sd3_1 hold104 (.A(_0060_),
    .X(net223));
 sg13g2_dlygate4sd3_1 hold105 (.A(\MVM_UART_SYSTEM.UART_RX.c_clocks[7] ),
    .X(net224));
 sg13g2_dlygate4sd3_1 hold106 (.A(_0294_),
    .X(net225));
 sg13g2_dlygate4sd3_1 hold107 (.A(_0074_),
    .X(net226));
 sg13g2_dlygate4sd3_1 hold108 (.A(_0017_),
    .X(net227));
 sg13g2_dlygate4sd3_1 hold109 (.A(_0106_),
    .X(net228));
 sg13g2_dlygate4sd3_1 hold110 (.A(\MVM_UART_SYSTEM.AXIS_MVM.SKID.buffer[0] ),
    .X(net229));
 sg13g2_dlygate4sd3_1 hold111 (.A(_0053_),
    .X(net230));
 sg13g2_dlygate4sd3_1 hold112 (.A(\MVM_UART_SYSTEM.AXIS_MVM.s_axis_kx_tvalid ),
    .X(net231));
 sg13g2_dlygate4sd3_1 hold113 (.A(_0127_),
    .X(net232));
 sg13g2_dlygate4sd3_1 hold114 (.A(\MVM_UART_SYSTEM.AXIS_MVM.SKID.buffer[11] ),
    .X(net233));
 sg13g2_dlygate4sd3_1 hold115 (.A(_0064_),
    .X(net234));
 sg13g2_dlygate4sd3_1 hold116 (.A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[2][6] ),
    .X(net235));
 sg13g2_dlygate4sd3_1 hold117 (.A(_0140_),
    .X(net236));
 sg13g2_dlygate4sd3_1 hold118 (.A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[6][5] ),
    .X(net237));
 sg13g2_dlygate4sd3_1 hold119 (.A(_0158_),
    .X(net238));
 sg13g2_dlygate4sd3_1 hold120 (.A(_0012_),
    .X(net239));
 sg13g2_dlygate4sd3_1 hold121 (.A(_0101_),
    .X(net240));
 sg13g2_dlygate4sd3_1 hold122 (.A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[2][2] ),
    .X(net241));
 sg13g2_dlygate4sd3_1 hold123 (.A(_0055_),
    .X(net242));
 sg13g2_dlygate4sd3_1 hold124 (.A(\MVM_UART_SYSTEM.AXIS_MVM.SKID.buffer[6] ),
    .X(net243));
 sg13g2_dlygate4sd3_1 hold125 (.A(\MVM_UART_SYSTEM.UART_TX.c_clocks[5] ),
    .X(net244));
 sg13g2_dlygate4sd3_1 hold126 (.A(_0262_),
    .X(net245));
 sg13g2_dlygate4sd3_1 hold127 (.A(_0046_),
    .X(net246));
 sg13g2_dlygate4sd3_1 hold128 (.A(_0013_),
    .X(net247));
 sg13g2_dlygate4sd3_1 hold129 (.A(_0102_),
    .X(net248));
 sg13g2_dlygate4sd3_1 hold130 (.A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[6][4] ),
    .X(net249));
 sg13g2_dlygate4sd3_1 hold131 (.A(_0494_),
    .X(net250));
 sg13g2_dlygate4sd3_1 hold132 (.A(_0157_),
    .X(net251));
 sg13g2_dlygate4sd3_1 hold133 (.A(_0016_),
    .X(net252));
 sg13g2_dlygate4sd3_1 hold134 (.A(_0105_),
    .X(net253));
 sg13g2_dlygate4sd3_1 hold135 (.A(_0029_),
    .X(net254));
 sg13g2_dlygate4sd3_1 hold136 (.A(_0118_),
    .X(net255));
 sg13g2_dlygate4sd3_1 hold137 (.A(_0028_),
    .X(net256));
 sg13g2_dlygate4sd3_1 hold138 (.A(_0117_),
    .X(net257));
 sg13g2_dlygate4sd3_1 hold139 (.A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[2][0] ),
    .X(net258));
 sg13g2_dlygate4sd3_1 hold140 (.A(_0134_),
    .X(net259));
 sg13g2_dlygate4sd3_1 hold141 (.A(\MVM_UART_SYSTEM.AXIS_MVM.SKID.buffer[12] ),
    .X(net260));
 sg13g2_dlygate4sd3_1 hold142 (.A(\MVM_UART_SYSTEM.UART_TX.c_pulses[4] ),
    .X(net261));
 sg13g2_dlygate4sd3_1 hold143 (.A(_0099_),
    .X(net262));
 sg13g2_dlygate4sd3_1 hold144 (.A(_0015_),
    .X(net263));
 sg13g2_dlygate4sd3_1 hold145 (.A(_0104_),
    .X(net264));
 sg13g2_dlygate4sd3_1 hold146 (.A(\MVM_UART_SYSTEM.AXIS_MVM.SKID.buffer[5] ),
    .X(net265));
 sg13g2_dlygate4sd3_1 hold147 (.A(\MVM_UART_SYSTEM.UART_TX.c_clocks[6] ),
    .X(net266));
 sg13g2_dlygate4sd3_1 hold148 (.A(_0047_),
    .X(net267));
 sg13g2_dlygate4sd3_1 hold149 (.A(\MVM_UART_SYSTEM.AXIS_MVM.SKID.buffer[4] ),
    .X(net268));
 sg13g2_dlygate4sd3_1 hold150 (.A(_0057_),
    .X(net269));
 sg13g2_dlygate4sd3_1 hold151 (.A(\MVM_UART_SYSTEM.AXIS_MVM.SKID.m_data[13] ),
    .X(net270));
 sg13g2_dlygate4sd3_1 hold152 (.A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[6][2] ),
    .X(net271));
 sg13g2_dlygate4sd3_1 hold153 (.A(_0155_),
    .X(net272));
 sg13g2_dlygate4sd3_1 hold154 (.A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[6][0] ),
    .X(net273));
 sg13g2_dlygate4sd3_1 hold155 (.A(_0478_),
    .X(net274));
 sg13g2_dlygate4sd3_1 hold156 (.A(_0153_),
    .X(net275));
 sg13g2_dlygate4sd3_1 hold157 (.A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[2][1] ),
    .X(net276));
 sg13g2_dlygate4sd3_1 hold158 (.A(_0135_),
    .X(net277));
 sg13g2_dlygate4sd3_1 hold159 (.A(\MVM_UART_SYSTEM.AXIS_MVM.SKID.m_data[3] ),
    .X(net278));
 sg13g2_dlygate4sd3_1 hold160 (.A(_0170_),
    .X(net279));
 sg13g2_dlygate4sd3_1 hold161 (.A(\MVM_UART_SYSTEM.UART_TX.c_clocks[4] ),
    .X(net280));
 sg13g2_dlygate4sd3_1 hold162 (.A(_0045_),
    .X(net281));
 sg13g2_dlygate4sd3_1 hold163 (.A(\MVM_UART_SYSTEM.UART_RX.c_clocks[1] ),
    .X(net282));
 sg13g2_dlygate4sd3_1 hold164 (.A(_0277_),
    .X(net283));
 sg13g2_dlygate4sd3_1 hold165 (.A(_0068_),
    .X(net284));
 sg13g2_dlygate4sd3_1 hold166 (.A(\MVM_UART_SYSTEM.AXIS_MVM.SKID.m_data[4] ),
    .X(net285));
 sg13g2_dlygate4sd3_1 hold167 (.A(_0171_),
    .X(net286));
 sg13g2_dlygate4sd3_1 hold168 (.A(\MVM_UART_SYSTEM.UART_TX.c_pulses[1] ),
    .X(net287));
 sg13g2_dlygate4sd3_1 hold169 (.A(_0311_),
    .X(net288));
 sg13g2_dlygate4sd3_1 hold170 (.A(_0096_),
    .X(net289));
 sg13g2_dlygate4sd3_1 hold171 (.A(\MVM_UART_SYSTEM.UART_TX.c_clocks[8] ),
    .X(net290));
 sg13g2_dlygate4sd3_1 hold172 (.A(\MVM_UART_SYSTEM.AXIS_MVM.SKID.s_valid ),
    .X(net291));
 sg13g2_dlygate4sd3_1 hold173 (.A(_0160_),
    .X(net292));
 sg13g2_dlygate4sd3_1 hold174 (.A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[4][5] ),
    .X(net293));
 sg13g2_dlygate4sd3_1 hold175 (.A(_0146_),
    .X(net294));
 sg13g2_dlygate4sd3_1 hold176 (.A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[2][4] ),
    .X(net295));
 sg13g2_dlygate4sd3_1 hold177 (.A(_0138_),
    .X(net296));
 sg13g2_dlygate4sd3_1 hold178 (.A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[1][5] ),
    .X(net297));
 sg13g2_dlygate4sd3_1 hold179 (.A(_0133_),
    .X(net298));
 sg13g2_dlygate4sd3_1 hold180 (.A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[2][3] ),
    .X(net299));
 sg13g2_dlygate4sd3_1 hold181 (.A(_0137_),
    .X(net300));
 sg13g2_dlygate4sd3_1 hold182 (.A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[6][1] ),
    .X(net301));
 sg13g2_dlygate4sd3_1 hold183 (.A(_0154_),
    .X(net302));
 sg13g2_dlygate4sd3_1 hold184 (.A(\MVM_UART_SYSTEM.UART_RX.c_clocks[10] ),
    .X(net303));
 sg13g2_dlygate4sd3_1 hold185 (.A(_0077_),
    .X(net304));
 sg13g2_dlygate4sd3_1 hold186 (.A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[1][1] ),
    .X(net305));
 sg13g2_dlygate4sd3_1 hold187 (.A(_0393_),
    .X(net306));
 sg13g2_dlygate4sd3_1 hold188 (.A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[5][5] ),
    .X(net307));
 sg13g2_dlygate4sd3_1 hold189 (.A(_0152_),
    .X(net308));
 sg13g2_dlygate4sd3_1 hold190 (.A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[1][2] ),
    .X(net309));
 sg13g2_dlygate4sd3_1 hold191 (.A(_0130_),
    .X(net310));
 sg13g2_dlygate4sd3_1 hold192 (.A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[0][0] ),
    .X(net311));
 sg13g2_dlygate4sd3_1 hold193 (.A(_0161_),
    .X(net312));
 sg13g2_dlygate4sd3_1 hold194 (.A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[0][5] ),
    .X(net313));
 sg13g2_dlygate4sd3_1 hold195 (.A(_0166_),
    .X(net314));
 sg13g2_dlygate4sd3_1 hold196 (.A(\MVM_UART_SYSTEM.UART_TX.c_pulses[2] ),
    .X(net315));
 sg13g2_dlygate4sd3_1 hold197 (.A(_0097_),
    .X(net316));
 sg13g2_dlygate4sd3_1 hold198 (.A(\MVM_UART_SYSTEM.UART_TX.c_clocks[11] ),
    .X(net317));
 sg13g2_dlygate4sd3_1 hold199 (.A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[4][0] ),
    .X(net318));
 sg13g2_dlygate4sd3_1 hold200 (.A(_0141_),
    .X(net319));
 sg13g2_dlygate4sd3_1 hold201 (.A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.k_pad[2][1] ),
    .X(net320));
 sg13g2_dlygate4sd3_1 hold202 (.A(_0364_),
    .X(net321));
 sg13g2_dlygate4sd3_1 hold203 (.A(_0365_),
    .X(net322));
 sg13g2_dlygate4sd3_1 hold204 (.A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[5][2] ),
    .X(net323));
 sg13g2_dlygate4sd3_1 hold205 (.A(_0149_),
    .X(net324));
 sg13g2_dlygate4sd3_1 hold206 (.A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[5][1] ),
    .X(net325));
 sg13g2_dlygate4sd3_1 hold207 (.A(_0148_),
    .X(net326));
 sg13g2_dlygate4sd3_1 hold208 (.A(\MVM_UART_SYSTEM.UART_RX.c_clocks[5] ),
    .X(net327));
 sg13g2_dlygate4sd3_1 hold209 (.A(_0292_),
    .X(net328));
 sg13g2_dlygate4sd3_1 hold210 (.A(_0072_),
    .X(net329));
 sg13g2_dlygate4sd3_1 hold211 (.A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[5][4] ),
    .X(net330));
 sg13g2_dlygate4sd3_1 hold212 (.A(\MVM_UART_SYSTEM.UART_RX.c_clocks[9] ),
    .X(net331));
 sg13g2_dlygate4sd3_1 hold213 (.A(_0299_),
    .X(net332));
 sg13g2_dlygate4sd3_1 hold214 (.A(_0076_),
    .X(net333));
 sg13g2_dlygate4sd3_1 hold215 (.A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[0][4] ),
    .X(net334));
 sg13g2_dlygate4sd3_1 hold216 (.A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[1][4] ),
    .X(net335));
 sg13g2_dlygate4sd3_1 hold217 (.A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[4][1] ),
    .X(net336));
 sg13g2_dlygate4sd3_1 hold218 (.A(_0142_),
    .X(net337));
 sg13g2_dlygate4sd3_1 hold219 (.A(\MVM_UART_SYSTEM.UART_TX.c_clocks[2] ),
    .X(net338));
 sg13g2_dlygate4sd3_1 hold220 (.A(_0259_),
    .X(net339));
 sg13g2_dlygate4sd3_1 hold221 (.A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[0][1] ),
    .X(net340));
 sg13g2_dlygate4sd3_1 hold222 (.A(_0162_),
    .X(net341));
 sg13g2_dlygate4sd3_1 hold223 (.A(\MVM_UART_SYSTEM.AXIS_MVM.SKID.state[0] ),
    .X(net342));
 sg13g2_dlygate4sd3_1 hold224 (.A(_0229_),
    .X(net343));
 sg13g2_dlygate4sd3_1 hold225 (.A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[4][4] ),
    .X(net344));
 sg13g2_dlygate4sd3_1 hold226 (.A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[5][0] ),
    .X(net345));
 sg13g2_dlygate4sd3_1 hold227 (.A(_0147_),
    .X(net346));
 sg13g2_dlygate4sd3_1 hold228 (.A(\MVM_UART_SYSTEM.UART_RX.c_clocks[0] ),
    .X(net347));
 sg13g2_dlygate4sd3_1 hold229 (.A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.k_pad[3][0] ),
    .X(net348));
 sg13g2_dlygate4sd3_1 hold230 (.A(_0310_),
    .X(net349));
 sg13g2_dlygate4sd3_1 hold231 (.A(_0086_),
    .X(net350));
 sg13g2_dlygate4sd3_1 hold232 (.A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[1][3] ),
    .X(net351));
 sg13g2_dlygate4sd3_1 hold233 (.A(_0131_),
    .X(net352));
 sg13g2_dlygate4sd3_1 hold234 (.A(\MVM_UART_SYSTEM.UART_RX.c_clocks[6] ),
    .X(net353));
 sg13g2_dlygate4sd3_1 hold235 (.A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[4][2] ),
    .X(net354));
 sg13g2_dlygate4sd3_1 hold236 (.A(_0143_),
    .X(net355));
 sg13g2_dlygate4sd3_1 hold237 (.A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[1][0] ),
    .X(net356));
 sg13g2_dlygate4sd3_1 hold238 (.A(_0128_),
    .X(net357));
 sg13g2_dlygate4sd3_1 hold239 (.A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[5][3] ),
    .X(net358));
 sg13g2_dlygate4sd3_1 hold240 (.A(_0462_),
    .X(net359));
 sg13g2_dlygate4sd3_1 hold241 (.A(\MVM_UART_SYSTEM.UART_RX.c_bits[0] ),
    .X(net360));
 sg13g2_dlygate4sd3_1 hold242 (.A(\MVM_UART_SYSTEM.UART_RX.c_bits[1] ),
    .X(net361));
 sg13g2_dlygate4sd3_1 hold243 (.A(_0002_),
    .X(net362));
 sg13g2_dlygate4sd3_1 hold244 (.A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[0][2] ),
    .X(net363));
 sg13g2_dlygate4sd3_1 hold245 (.A(_0163_),
    .X(net364));
 sg13g2_dlygate4sd3_1 hold246 (.A(\MVM_UART_SYSTEM.UART_TX.c_clocks[3] ),
    .X(net365));
 sg13g2_dlygate4sd3_1 hold247 (.A(_0261_),
    .X(net366));
 sg13g2_dlygate4sd3_1 hold248 (.A(\MVM_UART_SYSTEM.UART_TX.c_clocks[0] ),
    .X(net367));
 sg13g2_dlygate4sd3_1 hold249 (.A(_0041_),
    .X(net368));
 sg13g2_dlygate4sd3_1 hold250 (.A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[0][3] ),
    .X(net369));
 sg13g2_dlygate4sd3_1 hold251 (.A(\MVM_UART_SYSTEM.UART_RX.c_clocks[11] ),
    .X(net370));
 sg13g2_dlygate4sd3_1 hold252 (.A(_0078_),
    .X(net371));
 sg13g2_dlygate4sd3_1 hold253 (.A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.tree[4][3] ),
    .X(net372));
 sg13g2_dlygate4sd3_1 hold254 (.A(\MVM_UART_SYSTEM.UART_RX.c_clocks[2] ),
    .X(net373));
 sg13g2_dlygate4sd3_1 hold255 (.A(\MVM_UART_SYSTEM.UART_RX.c_clocks[3] ),
    .X(net374));
 sg13g2_dlygate4sd3_1 hold256 (.A(_0286_),
    .X(net375));
 sg13g2_dlygate4sd3_1 hold257 (.A(_0070_),
    .X(net376));
 sg13g2_dlygate4sd3_1 hold258 (.A(\MVM_UART_SYSTEM.UART_RX.c_clocks[8] ),
    .X(net377));
 sg13g2_dlygate4sd3_1 hold259 (.A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.k_pad[3][1] ),
    .X(net378));
 sg13g2_dlygate4sd3_1 hold260 (.A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.k_pad[1][0] ),
    .X(net379));
 sg13g2_dlygate4sd3_1 hold261 (.A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.x_pad[1][0] ),
    .X(net380));
 sg13g2_dlygate4sd3_1 hold262 (.A(_0308_),
    .X(net381));
 sg13g2_dlygate4sd3_1 hold263 (.A(_0082_),
    .X(net382));
 sg13g2_dlygate4sd3_1 hold264 (.A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.k_pad[1][1] ),
    .X(net383));
 sg13g2_dlygate4sd3_1 hold265 (.A(\MVM_UART_SYSTEM.UART_TX.c_pulses[0] ),
    .X(net384));
 sg13g2_dlygate4sd3_1 hold266 (.A(\MVM_UART_SYSTEM.UART_RX.c_clocks[4] ),
    .X(net385));
 sg13g2_dlygate4sd3_1 hold267 (.A(_0071_),
    .X(net386));
 sg13g2_dlygate4sd3_1 hold268 (.A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.x_pad[1][1] ),
    .X(net387));
 sg13g2_dlygate4sd3_1 hold269 (.A(_0084_),
    .X(net388));
 sg13g2_dlygate4sd3_1 hold270 (.A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.x_pad[0][2] ),
    .X(net389));
 sg13g2_dlygate4sd3_1 hold271 (.A(_0081_),
    .X(net390));
 sg13g2_dlygate4sd3_1 hold272 (.A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.k_pad[2][0] ),
    .X(net391));
 sg13g2_dlygate4sd3_1 hold273 (.A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.k_pad[0][0] ),
    .X(net392));
 sg13g2_dlygate4sd3_1 hold274 (.A(_0093_),
    .X(net393));
 sg13g2_dlygate4sd3_1 hold275 (.A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.x_pad[0][1] ),
    .X(net394));
 sg13g2_dlygate4sd3_1 hold276 (.A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.x_pad[1][3] ),
    .X(net395));
 sg13g2_dlygate4sd3_1 hold277 (.A(_0085_),
    .X(net396));
 sg13g2_dlygate4sd3_1 hold278 (.A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.x_pad[0][0] ),
    .X(net397));
 sg13g2_dlygate4sd3_1 hold279 (.A(\MVM_UART_SYSTEM.AXIS_MVM.MATVEC.k_pad[0][1] ),
    .X(net398));
 sg13g2_dlygate4sd3_1 hold280 (.A(\MVM_UART_SYSTEM.UART_TX.c_clocks[1] ),
    .X(net399));
 sg13g2_dlygate4sd3_1 hold281 (.A(\MVM_UART_SYSTEM.AXIS_MVM.SKID.state[1] ),
    .X(net400));
 sg13g2_dlygate4sd3_1 hold282 (.A(\MVM_UART_SYSTEM.UART_RX.c_clocks[4] ),
    .X(net401));
 sg13g2_dlygate4sd3_1 hold283 (.A(\MVM_UART_SYSTEM.UART_TX.c_clocks[1] ),
    .X(net402));
 sg13g2_dlygate4sd3_1 hold284 (.A(_0258_),
    .X(net403));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_fill_2 FILLER_8_245 ();
 sg13g2_fill_1 FILLER_8_247 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_4 FILLER_9_70 ();
 sg13g2_fill_2 FILLER_9_74 ();
 sg13g2_decap_8 FILLER_9_80 ();
 sg13g2_decap_8 FILLER_9_87 ();
 sg13g2_decap_8 FILLER_9_94 ();
 sg13g2_decap_8 FILLER_9_101 ();
 sg13g2_decap_8 FILLER_9_108 ();
 sg13g2_decap_8 FILLER_9_115 ();
 sg13g2_decap_8 FILLER_9_122 ();
 sg13g2_decap_8 FILLER_9_129 ();
 sg13g2_fill_1 FILLER_9_136 ();
 sg13g2_decap_4 FILLER_9_145 ();
 sg13g2_decap_8 FILLER_9_153 ();
 sg13g2_decap_8 FILLER_9_164 ();
 sg13g2_decap_8 FILLER_9_171 ();
 sg13g2_decap_8 FILLER_9_178 ();
 sg13g2_decap_8 FILLER_9_185 ();
 sg13g2_decap_8 FILLER_9_192 ();
 sg13g2_decap_8 FILLER_9_202 ();
 sg13g2_decap_8 FILLER_9_209 ();
 sg13g2_decap_8 FILLER_9_225 ();
 sg13g2_fill_2 FILLER_9_232 ();
 sg13g2_fill_2 FILLER_9_251 ();
 sg13g2_fill_1 FILLER_9_253 ();
 sg13g2_decap_8 FILLER_9_263 ();
 sg13g2_decap_8 FILLER_9_270 ();
 sg13g2_decap_8 FILLER_9_277 ();
 sg13g2_decap_8 FILLER_9_284 ();
 sg13g2_decap_8 FILLER_9_291 ();
 sg13g2_decap_8 FILLER_9_298 ();
 sg13g2_decap_8 FILLER_9_305 ();
 sg13g2_decap_8 FILLER_9_312 ();
 sg13g2_decap_8 FILLER_9_319 ();
 sg13g2_decap_8 FILLER_9_326 ();
 sg13g2_decap_8 FILLER_9_333 ();
 sg13g2_decap_8 FILLER_9_340 ();
 sg13g2_decap_8 FILLER_9_347 ();
 sg13g2_decap_8 FILLER_9_354 ();
 sg13g2_decap_8 FILLER_9_361 ();
 sg13g2_decap_8 FILLER_9_368 ();
 sg13g2_decap_8 FILLER_9_375 ();
 sg13g2_decap_8 FILLER_9_382 ();
 sg13g2_decap_8 FILLER_9_389 ();
 sg13g2_decap_8 FILLER_9_396 ();
 sg13g2_decap_4 FILLER_9_403 ();
 sg13g2_fill_2 FILLER_9_407 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_fill_2 FILLER_10_63 ();
 sg13g2_fill_1 FILLER_10_83 ();
 sg13g2_fill_2 FILLER_10_93 ();
 sg13g2_decap_8 FILLER_10_104 ();
 sg13g2_decap_8 FILLER_10_111 ();
 sg13g2_decap_4 FILLER_10_118 ();
 sg13g2_fill_2 FILLER_10_122 ();
 sg13g2_fill_1 FILLER_10_150 ();
 sg13g2_fill_2 FILLER_10_165 ();
 sg13g2_fill_2 FILLER_10_171 ();
 sg13g2_fill_1 FILLER_10_199 ();
 sg13g2_fill_2 FILLER_10_209 ();
 sg13g2_decap_8 FILLER_10_268 ();
 sg13g2_fill_2 FILLER_10_275 ();
 sg13g2_fill_1 FILLER_10_277 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_4 FILLER_11_49 ();
 sg13g2_fill_2 FILLER_11_53 ();
 sg13g2_fill_1 FILLER_11_60 ();
 sg13g2_fill_1 FILLER_11_113 ();
 sg13g2_fill_2 FILLER_11_137 ();
 sg13g2_fill_1 FILLER_11_139 ();
 sg13g2_fill_1 FILLER_11_167 ();
 sg13g2_decap_4 FILLER_11_178 ();
 sg13g2_fill_2 FILLER_11_182 ();
 sg13g2_fill_1 FILLER_11_192 ();
 sg13g2_decap_4 FILLER_11_213 ();
 sg13g2_fill_1 FILLER_11_257 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_fill_2 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_fill_1 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_341 ();
 sg13g2_decap_8 FILLER_11_348 ();
 sg13g2_fill_2 FILLER_11_355 ();
 sg13g2_decap_8 FILLER_11_361 ();
 sg13g2_fill_1 FILLER_11_368 ();
 sg13g2_decap_8 FILLER_11_373 ();
 sg13g2_decap_8 FILLER_11_380 ();
 sg13g2_decap_8 FILLER_11_387 ();
 sg13g2_decap_8 FILLER_11_394 ();
 sg13g2_decap_8 FILLER_11_401 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_fill_2 FILLER_12_49 ();
 sg13g2_fill_2 FILLER_12_67 ();
 sg13g2_fill_1 FILLER_12_69 ();
 sg13g2_fill_1 FILLER_12_126 ();
 sg13g2_fill_1 FILLER_12_136 ();
 sg13g2_fill_2 FILLER_12_146 ();
 sg13g2_fill_2 FILLER_12_170 ();
 sg13g2_fill_1 FILLER_12_172 ();
 sg13g2_fill_1 FILLER_12_199 ();
 sg13g2_fill_2 FILLER_12_224 ();
 sg13g2_fill_1 FILLER_12_226 ();
 sg13g2_fill_1 FILLER_12_232 ();
 sg13g2_fill_2 FILLER_12_264 ();
 sg13g2_fill_1 FILLER_12_266 ();
 sg13g2_decap_4 FILLER_12_316 ();
 sg13g2_fill_1 FILLER_12_320 ();
 sg13g2_decap_4 FILLER_12_326 ();
 sg13g2_fill_1 FILLER_12_330 ();
 sg13g2_fill_2 FILLER_12_368 ();
 sg13g2_fill_1 FILLER_12_370 ();
 sg13g2_fill_1 FILLER_12_376 ();
 sg13g2_decap_8 FILLER_12_390 ();
 sg13g2_decap_8 FILLER_12_401 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_fill_2 FILLER_13_35 ();
 sg13g2_decap_4 FILLER_13_50 ();
 sg13g2_fill_2 FILLER_13_62 ();
 sg13g2_fill_1 FILLER_13_64 ();
 sg13g2_fill_2 FILLER_13_80 ();
 sg13g2_fill_1 FILLER_13_91 ();
 sg13g2_fill_1 FILLER_13_136 ();
 sg13g2_fill_2 FILLER_13_163 ();
 sg13g2_fill_1 FILLER_13_165 ();
 sg13g2_fill_2 FILLER_13_190 ();
 sg13g2_fill_1 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_4 FILLER_14_28 ();
 sg13g2_fill_2 FILLER_14_41 ();
 sg13g2_fill_2 FILLER_14_67 ();
 sg13g2_fill_2 FILLER_14_108 ();
 sg13g2_fill_1 FILLER_14_110 ();
 sg13g2_fill_2 FILLER_14_146 ();
 sg13g2_decap_4 FILLER_14_177 ();
 sg13g2_fill_1 FILLER_14_207 ();
 sg13g2_fill_2 FILLER_14_276 ();
 sg13g2_fill_1 FILLER_14_278 ();
 sg13g2_fill_1 FILLER_14_304 ();
 sg13g2_fill_2 FILLER_14_330 ();
 sg13g2_fill_2 FILLER_14_388 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_4 FILLER_15_21 ();
 sg13g2_fill_1 FILLER_15_25 ();
 sg13g2_fill_1 FILLER_15_61 ();
 sg13g2_fill_1 FILLER_15_67 ();
 sg13g2_fill_1 FILLER_15_80 ();
 sg13g2_fill_1 FILLER_15_98 ();
 sg13g2_fill_1 FILLER_15_124 ();
 sg13g2_fill_1 FILLER_15_135 ();
 sg13g2_fill_2 FILLER_15_208 ();
 sg13g2_fill_1 FILLER_15_210 ();
 sg13g2_fill_2 FILLER_15_220 ();
 sg13g2_fill_2 FILLER_15_248 ();
 sg13g2_fill_2 FILLER_15_386 ();
 sg13g2_fill_1 FILLER_15_388 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_fill_1 FILLER_16_21 ();
 sg13g2_fill_1 FILLER_16_42 ();
 sg13g2_fill_1 FILLER_16_113 ();
 sg13g2_fill_2 FILLER_16_127 ();
 sg13g2_fill_1 FILLER_16_129 ();
 sg13g2_fill_1 FILLER_16_161 ();
 sg13g2_fill_1 FILLER_16_193 ();
 sg13g2_fill_1 FILLER_16_225 ();
 sg13g2_fill_2 FILLER_16_273 ();
 sg13g2_fill_2 FILLER_16_330 ();
 sg13g2_fill_1 FILLER_16_332 ();
 sg13g2_fill_2 FILLER_16_361 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_4 FILLER_17_21 ();
 sg13g2_fill_2 FILLER_17_25 ();
 sg13g2_fill_1 FILLER_17_56 ();
 sg13g2_fill_1 FILLER_17_65 ();
 sg13g2_fill_2 FILLER_17_80 ();
 sg13g2_fill_1 FILLER_17_108 ();
 sg13g2_fill_1 FILLER_17_123 ();
 sg13g2_fill_2 FILLER_17_133 ();
 sg13g2_fill_1 FILLER_17_135 ();
 sg13g2_fill_2 FILLER_17_218 ();
 sg13g2_fill_1 FILLER_17_220 ();
 sg13g2_fill_2 FILLER_17_280 ();
 sg13g2_fill_2 FILLER_17_308 ();
 sg13g2_fill_2 FILLER_17_402 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_fill_2 FILLER_18_21 ();
 sg13g2_fill_1 FILLER_18_83 ();
 sg13g2_fill_1 FILLER_18_99 ();
 sg13g2_fill_1 FILLER_18_140 ();
 sg13g2_fill_2 FILLER_18_203 ();
 sg13g2_fill_2 FILLER_18_210 ();
 sg13g2_fill_1 FILLER_18_280 ();
 sg13g2_fill_2 FILLER_18_360 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_4 FILLER_19_14 ();
 sg13g2_fill_1 FILLER_19_18 ();
 sg13g2_fill_2 FILLER_19_51 ();
 sg13g2_fill_1 FILLER_19_62 ();
 sg13g2_fill_1 FILLER_19_139 ();
 sg13g2_fill_1 FILLER_19_145 ();
 sg13g2_fill_2 FILLER_19_207 ();
 sg13g2_fill_1 FILLER_19_209 ();
 sg13g2_fill_2 FILLER_19_245 ();
 sg13g2_fill_1 FILLER_19_247 ();
 sg13g2_fill_2 FILLER_19_258 ();
 sg13g2_fill_1 FILLER_19_260 ();
 sg13g2_fill_1 FILLER_19_312 ();
 sg13g2_fill_2 FILLER_19_328 ();
 sg13g2_fill_1 FILLER_19_330 ();
 sg13g2_fill_1 FILLER_19_349 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_4 FILLER_20_14 ();
 sg13g2_fill_2 FILLER_20_105 ();
 sg13g2_fill_2 FILLER_20_152 ();
 sg13g2_fill_1 FILLER_20_158 ();
 sg13g2_fill_1 FILLER_20_163 ();
 sg13g2_fill_2 FILLER_20_187 ();
 sg13g2_fill_1 FILLER_20_189 ();
 sg13g2_fill_2 FILLER_20_370 ();
 sg13g2_fill_2 FILLER_20_407 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_4 FILLER_21_14 ();
 sg13g2_fill_2 FILLER_21_18 ();
 sg13g2_fill_1 FILLER_21_61 ();
 sg13g2_fill_2 FILLER_21_116 ();
 sg13g2_fill_1 FILLER_21_118 ();
 sg13g2_fill_2 FILLER_21_124 ();
 sg13g2_fill_1 FILLER_21_126 ();
 sg13g2_fill_2 FILLER_21_132 ();
 sg13g2_fill_1 FILLER_21_134 ();
 sg13g2_fill_1 FILLER_21_147 ();
 sg13g2_fill_1 FILLER_21_174 ();
 sg13g2_fill_1 FILLER_21_182 ();
 sg13g2_fill_2 FILLER_21_205 ();
 sg13g2_fill_2 FILLER_21_212 ();
 sg13g2_decap_8 FILLER_21_218 ();
 sg13g2_fill_1 FILLER_21_287 ();
 sg13g2_fill_1 FILLER_21_311 ();
 sg13g2_fill_2 FILLER_21_329 ();
 sg13g2_fill_1 FILLER_21_354 ();
 sg13g2_fill_1 FILLER_21_365 ();
 sg13g2_fill_1 FILLER_21_376 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_fill_2 FILLER_22_57 ();
 sg13g2_fill_1 FILLER_22_84 ();
 sg13g2_fill_1 FILLER_22_94 ();
 sg13g2_fill_2 FILLER_22_114 ();
 sg13g2_fill_1 FILLER_22_133 ();
 sg13g2_fill_2 FILLER_22_190 ();
 sg13g2_fill_2 FILLER_22_201 ();
 sg13g2_fill_2 FILLER_22_281 ();
 sg13g2_fill_1 FILLER_22_384 ();
 sg13g2_fill_1 FILLER_22_399 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_fill_2 FILLER_23_21 ();
 sg13g2_fill_1 FILLER_23_23 ();
 sg13g2_decap_4 FILLER_23_36 ();
 sg13g2_fill_2 FILLER_23_49 ();
 sg13g2_fill_1 FILLER_23_51 ();
 sg13g2_fill_1 FILLER_23_108 ();
 sg13g2_fill_1 FILLER_23_117 ();
 sg13g2_fill_2 FILLER_23_123 ();
 sg13g2_fill_1 FILLER_23_125 ();
 sg13g2_fill_1 FILLER_23_136 ();
 sg13g2_fill_1 FILLER_23_157 ();
 sg13g2_fill_1 FILLER_23_163 ();
 sg13g2_fill_2 FILLER_23_177 ();
 sg13g2_fill_1 FILLER_23_224 ();
 sg13g2_fill_2 FILLER_23_268 ();
 sg13g2_fill_1 FILLER_23_270 ();
 sg13g2_fill_1 FILLER_23_307 ();
 sg13g2_fill_2 FILLER_23_333 ();
 sg13g2_fill_1 FILLER_23_335 ();
 sg13g2_fill_1 FILLER_23_373 ();
 sg13g2_fill_2 FILLER_23_393 ();
 sg13g2_fill_1 FILLER_23_395 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_fill_2 FILLER_24_44 ();
 sg13g2_fill_1 FILLER_24_51 ();
 sg13g2_fill_2 FILLER_24_60 ();
 sg13g2_fill_1 FILLER_24_81 ();
 sg13g2_fill_1 FILLER_24_99 ();
 sg13g2_fill_2 FILLER_24_192 ();
 sg13g2_fill_2 FILLER_24_311 ();
 sg13g2_fill_1 FILLER_24_313 ();
 sg13g2_fill_2 FILLER_24_371 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_fill_2 FILLER_25_35 ();
 sg13g2_fill_1 FILLER_25_37 ();
 sg13g2_fill_2 FILLER_25_54 ();
 sg13g2_fill_1 FILLER_25_56 ();
 sg13g2_fill_1 FILLER_25_66 ();
 sg13g2_fill_1 FILLER_25_111 ();
 sg13g2_fill_2 FILLER_25_151 ();
 sg13g2_fill_1 FILLER_25_162 ();
 sg13g2_fill_2 FILLER_25_213 ();
 sg13g2_fill_2 FILLER_25_327 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_4 FILLER_26_21 ();
 sg13g2_fill_1 FILLER_26_25 ();
 sg13g2_fill_2 FILLER_26_43 ();
 sg13g2_fill_1 FILLER_26_50 ();
 sg13g2_fill_2 FILLER_26_80 ();
 sg13g2_fill_1 FILLER_26_82 ();
 sg13g2_fill_1 FILLER_26_121 ();
 sg13g2_fill_2 FILLER_26_190 ();
 sg13g2_fill_1 FILLER_26_192 ();
 sg13g2_fill_2 FILLER_26_255 ();
 sg13g2_fill_1 FILLER_26_267 ();
 sg13g2_fill_1 FILLER_26_299 ();
 sg13g2_fill_1 FILLER_26_408 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_fill_2 FILLER_27_21 ();
 sg13g2_fill_1 FILLER_27_23 ();
 sg13g2_fill_2 FILLER_27_99 ();
 sg13g2_fill_1 FILLER_27_115 ();
 sg13g2_fill_1 FILLER_27_142 ();
 sg13g2_fill_2 FILLER_27_157 ();
 sg13g2_fill_1 FILLER_27_159 ();
 sg13g2_fill_2 FILLER_27_407 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_fill_2 FILLER_28_42 ();
 sg13g2_fill_2 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_60 ();
 sg13g2_fill_1 FILLER_28_67 ();
 sg13g2_fill_1 FILLER_28_158 ();
 sg13g2_fill_1 FILLER_28_258 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_4 FILLER_29_28 ();
 sg13g2_fill_2 FILLER_29_152 ();
 sg13g2_fill_2 FILLER_29_197 ();
 sg13g2_fill_1 FILLER_29_199 ();
 sg13g2_fill_2 FILLER_29_267 ();
 sg13g2_fill_1 FILLER_29_278 ();
 sg13g2_fill_1 FILLER_29_375 ();
 sg13g2_fill_2 FILLER_29_407 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_4 FILLER_30_28 ();
 sg13g2_fill_1 FILLER_30_32 ();
 sg13g2_fill_2 FILLER_30_76 ();
 sg13g2_fill_1 FILLER_30_78 ();
 sg13g2_fill_1 FILLER_30_112 ();
 sg13g2_fill_1 FILLER_30_123 ();
 sg13g2_fill_2 FILLER_30_170 ();
 sg13g2_fill_1 FILLER_30_172 ();
 sg13g2_fill_2 FILLER_30_202 ();
 sg13g2_fill_1 FILLER_30_317 ();
 sg13g2_fill_2 FILLER_30_357 ();
 sg13g2_fill_1 FILLER_30_408 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_4 FILLER_31_21 ();
 sg13g2_fill_2 FILLER_31_25 ();
 sg13g2_fill_2 FILLER_31_65 ();
 sg13g2_fill_1 FILLER_31_67 ();
 sg13g2_fill_1 FILLER_31_94 ();
 sg13g2_fill_2 FILLER_31_212 ();
 sg13g2_fill_1 FILLER_31_214 ();
 sg13g2_fill_1 FILLER_31_275 ();
 sg13g2_fill_2 FILLER_31_297 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_4 FILLER_32_28 ();
 sg13g2_fill_1 FILLER_32_50 ();
 sg13g2_fill_2 FILLER_32_75 ();
 sg13g2_fill_1 FILLER_32_104 ();
 sg13g2_fill_1 FILLER_32_201 ();
 sg13g2_fill_1 FILLER_32_212 ();
 sg13g2_fill_2 FILLER_32_255 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_fill_2 FILLER_33_92 ();
 sg13g2_fill_1 FILLER_33_94 ();
 sg13g2_fill_2 FILLER_33_137 ();
 sg13g2_fill_2 FILLER_33_148 ();
 sg13g2_fill_2 FILLER_33_282 ();
 sg13g2_fill_1 FILLER_33_315 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_fill_2 FILLER_34_21 ();
 sg13g2_fill_2 FILLER_34_61 ();
 sg13g2_fill_1 FILLER_34_63 ();
 sg13g2_fill_2 FILLER_34_110 ();
 sg13g2_fill_1 FILLER_34_112 ();
 sg13g2_fill_1 FILLER_34_118 ();
 sg13g2_fill_1 FILLER_34_164 ();
 sg13g2_fill_2 FILLER_34_248 ();
 sg13g2_fill_1 FILLER_34_286 ();
 sg13g2_fill_1 FILLER_34_330 ();
 sg13g2_fill_2 FILLER_34_407 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_4 FILLER_35_21 ();
 sg13g2_fill_1 FILLER_35_25 ();
 sg13g2_fill_1 FILLER_35_62 ();
 sg13g2_fill_2 FILLER_35_106 ();
 sg13g2_fill_2 FILLER_35_144 ();
 sg13g2_fill_2 FILLER_35_191 ();
 sg13g2_fill_1 FILLER_35_193 ();
 sg13g2_fill_1 FILLER_35_252 ();
 sg13g2_fill_2 FILLER_35_291 ();
 sg13g2_fill_2 FILLER_35_336 ();
 sg13g2_fill_1 FILLER_35_355 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_fill_2 FILLER_36_21 ();
 sg13g2_fill_1 FILLER_36_23 ();
 sg13g2_fill_2 FILLER_36_85 ();
 sg13g2_fill_1 FILLER_36_123 ();
 sg13g2_fill_1 FILLER_36_163 ();
 sg13g2_fill_1 FILLER_36_226 ();
 sg13g2_fill_2 FILLER_36_246 ();
 sg13g2_fill_1 FILLER_36_296 ();
 sg13g2_fill_2 FILLER_36_335 ();
 sg13g2_fill_1 FILLER_36_408 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_fill_2 FILLER_37_14 ();
 sg13g2_fill_2 FILLER_37_147 ();
 sg13g2_fill_1 FILLER_37_163 ();
 sg13g2_fill_2 FILLER_37_178 ();
 sg13g2_fill_1 FILLER_37_304 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_fill_2 FILLER_38_7 ();
 sg13g2_fill_1 FILLER_38_9 ();
 sg13g2_fill_1 FILLER_38_90 ();
 sg13g2_fill_1 FILLER_38_286 ();
 sg13g2_fill_1 FILLER_38_329 ();
 assign uio_oe[0] = net2;
 assign uio_oe[1] = net3;
 assign uio_oe[2] = net4;
 assign uio_oe[3] = net5;
 assign uio_oe[4] = net6;
 assign uio_oe[5] = net7;
 assign uio_oe[6] = net8;
 assign uio_oe[7] = net9;
 assign uio_out[0] = net10;
 assign uio_out[1] = net11;
 assign uio_out[2] = net12;
 assign uio_out[3] = net13;
 assign uio_out[4] = net14;
 assign uio_out[5] = net15;
 assign uio_out[6] = net16;
 assign uio_out[7] = net17;
 assign uo_out[1] = net18;
 assign uo_out[2] = net19;
 assign uo_out[3] = net20;
 assign uo_out[4] = net21;
 assign uo_out[5] = net22;
 assign uo_out[6] = net23;
 assign uo_out[7] = net24;
endmodule

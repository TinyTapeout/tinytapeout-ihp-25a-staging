module tt_um_stochastic_integrator_tt9_CL123abc (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire clknet_leaf_0_clk;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire \clk_counter[0] ;
 wire \clk_counter[10] ;
 wire \clk_counter[11] ;
 wire \clk_counter[12] ;
 wire \clk_counter[13] ;
 wire \clk_counter[14] ;
 wire \clk_counter[15] ;
 wire \clk_counter[16] ;
 wire \clk_counter[17] ;
 wire \clk_counter[1] ;
 wire \clk_counter[2] ;
 wire \clk_counter[3] ;
 wire \clk_counter[4] ;
 wire \clk_counter[5] ;
 wire \clk_counter[6] ;
 wire \clk_counter[7] ;
 wire \clk_counter[8] ;
 wire \clk_counter[9] ;
 wire \input_a_sng_comparator.bits_a[0] ;
 wire \input_a_sng_comparator.bits_a[1] ;
 wire \input_a_sng_comparator.bits_a[2] ;
 wire \input_a_sng_comparator.bits_a[3] ;
 wire \input_a_sng_comparator.bits_a[4] ;
 wire \input_a_sng_comparator.bits_a[5] ;
 wire \input_a_sng_comparator.bits_a[6] ;
 wire \input_a_sng_comparator.bits_a[7] ;
 wire \input_a_sng_comparator.bits_a[8] ;
 wire \input_a_sng_comparator.bits_b[0] ;
 wire \input_a_sng_comparator.bits_b[1] ;
 wire \input_a_sng_comparator.bits_b[2] ;
 wire \input_a_sng_comparator.bits_b[3] ;
 wire \input_a_sng_comparator.bits_b[4] ;
 wire \input_a_sng_comparator.bits_b[5] ;
 wire \input_a_sng_comparator.bits_b[6] ;
 wire \input_a_sng_comparator.bits_b[7] ;
 wire \input_a_sng_comparator.bits_b[8] ;
 wire \input_b_sng_comparator.bits_a[0] ;
 wire \input_b_sng_comparator.bits_a[1] ;
 wire \input_b_sng_comparator.bits_a[2] ;
 wire \input_b_sng_comparator.bits_a[3] ;
 wire \input_b_sng_comparator.bits_a[4] ;
 wire \input_b_sng_comparator.bits_a[5] ;
 wire \input_b_sng_comparator.bits_a[6] ;
 wire \input_b_sng_comparator.bits_a[7] ;
 wire \input_b_sng_comparator.bits_a[8] ;
 wire \input_b_sng_comparator.bits_b[0] ;
 wire \input_b_sng_comparator.bits_b[1] ;
 wire \input_b_sng_comparator.bits_b[2] ;
 wire \input_halfprob1_sng_comparator.bits_b[0] ;
 wire \input_halfprob1_sng_comparator.bits_b[1] ;
 wire \input_halfprob1_sng_comparator.bits_b[6] ;
 wire \input_halfprob1_sng_comparator.bits_b[7] ;
 wire \input_halfprob1_sng_comparator.bits_b[8] ;
 wire \input_halfprob2_sng_comparator.bits_b[1] ;
 wire \input_halfprob2_sng_comparator.bits_b[2] ;
 wire \input_halfprob2_sng_comparator.bits_b[3] ;
 wire \input_halfprob2_sng_comparator.bits_b[4] ;
 wire \input_halfprob2_sng_comparator.bits_b[5] ;
 wire \input_halfprob2_sng_comparator.bits_b[6] ;
 wire \input_halfprob2_sng_comparator.bits_b[7] ;
 wire \input_halfprob2_sng_comparator.bits_b[8] ;
 wire \integrator_a_counter.value_output[0] ;
 wire \integrator_a_counter.value_output[1] ;
 wire \integrator_a_counter.value_output[2] ;
 wire \integrator_a_counter.value_output[3] ;
 wire \integrator_a_counter.value_output[4] ;
 wire \integrator_a_counter.value_output[5] ;
 wire \integrator_a_counter.value_output[6] ;
 wire \integrator_a_counter.value_output[7] ;
 wire \integrator_a_counter.value_output[8] ;
 wire \integrator_a_output.bitseq[0] ;
 wire \integrator_a_output.bitseq[1] ;
 wire \integrator_a_output.bitseq[2] ;
 wire \integrator_a_output.bitseq[3] ;
 wire \integrator_a_output.bitseq[4] ;
 wire \integrator_a_output.bitseq[5] ;
 wire \integrator_a_output.bitseq[6] ;
 wire \integrator_a_output.bitseq[7] ;
 wire \integrator_a_output.counter[0] ;
 wire \integrator_a_output.counter[1] ;
 wire \integrator_a_output.counter[2] ;
 wire \integrator_a_output.counter[3] ;
 wire \integrator_a_output.input_bits[0] ;
 wire \integrator_a_output.input_bits[1] ;
 wire \integrator_a_output.input_bits[2] ;
 wire \integrator_a_output.input_bits[3] ;
 wire \integrator_a_output.input_bits[4] ;
 wire \integrator_a_output.input_bits[5] ;
 wire \integrator_a_output.input_bits[6] ;
 wire \integrator_a_output.input_bits[7] ;
 wire \integrator_a_output.input_bits[8] ;
 wire \integrator_a_output.output_bit ;
 wire \integrator_a_sng_comparator.bits_b[1] ;
 wire \integrator_b_counter.value_output[0] ;
 wire \integrator_b_counter.value_output[1] ;
 wire \integrator_b_counter.value_output[2] ;
 wire \integrator_b_counter.value_output[3] ;
 wire \integrator_b_counter.value_output[4] ;
 wire \integrator_b_counter.value_output[5] ;
 wire \integrator_b_counter.value_output[6] ;
 wire \integrator_b_counter.value_output[7] ;
 wire \integrator_b_counter.value_output[8] ;
 wire \integrator_b_output.bitseq[0] ;
 wire \integrator_b_output.bitseq[1] ;
 wire \integrator_b_output.bitseq[2] ;
 wire \integrator_b_output.bitseq[3] ;
 wire \integrator_b_output.bitseq[4] ;
 wire \integrator_b_output.bitseq[5] ;
 wire \integrator_b_output.bitseq[6] ;
 wire \integrator_b_output.bitseq[7] ;
 wire \integrator_b_output.counter[0] ;
 wire \integrator_b_output.counter[1] ;
 wire \integrator_b_output.counter[2] ;
 wire \integrator_b_output.counter[3] ;
 wire \integrator_b_output.input_bits[0] ;
 wire \integrator_b_output.input_bits[1] ;
 wire \integrator_b_output.input_bits[2] ;
 wire \integrator_b_output.input_bits[3] ;
 wire \integrator_b_output.input_bits[4] ;
 wire \integrator_b_output.input_bits[5] ;
 wire \integrator_b_output.input_bits[6] ;
 wire \integrator_b_output.input_bits[7] ;
 wire \integrator_b_output.input_bits[8] ;
 wire \integrator_b_output.output_bit ;
 wire \integrator_b_sng_comparator.bits_b[6] ;
 wire \integrator_b_sng_comparator.bits_b[7] ;
 wire \integrator_b_sng_comparator.bits_b[8] ;
 wire \integrator_c_counter.value_output[0] ;
 wire \integrator_c_counter.value_output[1] ;
 wire \integrator_c_counter.value_output[2] ;
 wire \integrator_c_counter.value_output[3] ;
 wire \integrator_c_counter.value_output[4] ;
 wire \integrator_c_counter.value_output[5] ;
 wire \integrator_c_counter.value_output[6] ;
 wire \integrator_c_counter.value_output[7] ;
 wire \integrator_c_counter.value_output[8] ;
 wire \integrator_c_output.bitseq[0] ;
 wire \integrator_c_output.bitseq[1] ;
 wire \integrator_c_output.bitseq[2] ;
 wire \integrator_c_output.bitseq[3] ;
 wire \integrator_c_output.bitseq[4] ;
 wire \integrator_c_output.bitseq[5] ;
 wire \integrator_c_output.bitseq[6] ;
 wire \integrator_c_output.bitseq[7] ;
 wire \integrator_c_output.counter[0] ;
 wire \integrator_c_output.counter[1] ;
 wire \integrator_c_output.counter[2] ;
 wire \integrator_c_output.counter[3] ;
 wire \integrator_c_output.input_bits[0] ;
 wire \integrator_c_output.input_bits[1] ;
 wire \integrator_c_output.input_bits[2] ;
 wire \integrator_c_output.input_bits[3] ;
 wire \integrator_c_output.input_bits[4] ;
 wire \integrator_c_output.input_bits[5] ;
 wire \integrator_c_output.input_bits[6] ;
 wire \integrator_c_output.input_bits[7] ;
 wire \integrator_c_output.input_bits[8] ;
 wire \integrator_c_output.output_bit ;
 wire integrator_c_sn_bit;
 wire \integrator_c_sng_comparator.bits_b[0] ;
 wire \integrator_c_sng_comparator.bits_b[3] ;
 wire \serial_input.adjustment[0] ;
 wire \serial_input.adjustment[1] ;
 wire \serial_input.adjustment[2] ;
 wire \serial_input.adjustment[3] ;
 wire \serial_input.adjustment[4] ;
 wire \serial_input.loop ;
 wire \serial_input.output_bitcounter_1[0] ;
 wire \serial_input.output_bitcounter_1[1] ;
 wire \serial_input.output_bitcounter_1[2] ;
 wire \serial_input.output_bitcounter_1[3] ;
 wire \serial_input.output_bitcounter_1[4] ;
 wire \serial_input.output_bitcounter_1[5] ;
 wire \serial_input.output_bitcounter_1[6] ;
 wire \serial_input.output_bitcounter_1[7] ;
 wire \serial_input.output_bitcounter_1[8] ;
 wire \serial_input.output_bitcounter_2[0] ;
 wire \serial_input.output_bitcounter_2[1] ;
 wire \serial_input.output_bitcounter_2[2] ;
 wire \serial_input.output_bitcounter_2[3] ;
 wire \serial_input.output_bitcounter_2[4] ;
 wire \serial_input.output_bitcounter_2[5] ;
 wire \serial_input.output_bitcounter_2[6] ;
 wire \serial_input.output_bitcounter_2[7] ;
 wire \serial_input.output_bitcounter_2[8] ;
 wire \serial_input.output_case[0] ;
 wire \serial_input.output_case[1] ;
 wire \serial_input.output_case[2] ;
 wire \serial_input.output_case[3] ;
 wire \system_integrator_a_counter.init_flag ;
 wire \system_integrator_a_counter.value_output[0] ;
 wire \system_integrator_a_counter.value_output[1] ;
 wire \system_integrator_a_counter.value_output[2] ;
 wire \system_integrator_a_counter.value_output[3] ;
 wire \system_integrator_a_counter.value_output[4] ;
 wire \system_integrator_a_counter.value_output[5] ;
 wire \system_integrator_a_counter.value_output[6] ;
 wire \system_integrator_a_counter.value_output[7] ;
 wire \system_integrator_a_counter.value_output[8] ;
 wire \system_integrator_a_output.bitseq[0] ;
 wire \system_integrator_a_output.bitseq[1] ;
 wire \system_integrator_a_output.bitseq[2] ;
 wire \system_integrator_a_output.bitseq[3] ;
 wire \system_integrator_a_output.bitseq[4] ;
 wire \system_integrator_a_output.bitseq[5] ;
 wire \system_integrator_a_output.bitseq[6] ;
 wire \system_integrator_a_output.bitseq[7] ;
 wire \system_integrator_a_output.counter[0] ;
 wire \system_integrator_a_output.counter[1] ;
 wire \system_integrator_a_output.counter[2] ;
 wire \system_integrator_a_output.counter[3] ;
 wire \system_integrator_a_output.input_bits[0] ;
 wire \system_integrator_a_output.input_bits[1] ;
 wire \system_integrator_a_output.input_bits[2] ;
 wire \system_integrator_a_output.input_bits[3] ;
 wire \system_integrator_a_output.input_bits[4] ;
 wire \system_integrator_a_output.input_bits[5] ;
 wire \system_integrator_a_output.input_bits[6] ;
 wire \system_integrator_a_output.input_bits[7] ;
 wire \system_integrator_a_output.input_bits[8] ;
 wire \system_integrator_a_output.output_bit ;
 wire \system_integrator_b_counter.value_output[0] ;
 wire \system_integrator_b_counter.value_output[1] ;
 wire \system_integrator_b_counter.value_output[2] ;
 wire \system_integrator_b_counter.value_output[3] ;
 wire \system_integrator_b_counter.value_output[4] ;
 wire \system_integrator_b_counter.value_output[5] ;
 wire \system_integrator_b_counter.value_output[6] ;
 wire \system_integrator_b_counter.value_output[7] ;
 wire \system_integrator_b_counter.value_output[8] ;
 wire \system_integrator_b_output.bitseq[0] ;
 wire \system_integrator_b_output.bitseq[1] ;
 wire \system_integrator_b_output.bitseq[2] ;
 wire \system_integrator_b_output.bitseq[3] ;
 wire \system_integrator_b_output.bitseq[4] ;
 wire \system_integrator_b_output.bitseq[5] ;
 wire \system_integrator_b_output.bitseq[6] ;
 wire \system_integrator_b_output.bitseq[7] ;
 wire \system_integrator_b_output.counter[0] ;
 wire \system_integrator_b_output.counter[1] ;
 wire \system_integrator_b_output.counter[2] ;
 wire \system_integrator_b_output.counter[3] ;
 wire \system_integrator_b_output.input_bits[0] ;
 wire \system_integrator_b_output.input_bits[1] ;
 wire \system_integrator_b_output.input_bits[2] ;
 wire \system_integrator_b_output.input_bits[3] ;
 wire \system_integrator_b_output.input_bits[4] ;
 wire \system_integrator_b_output.input_bits[5] ;
 wire \system_integrator_b_output.input_bits[6] ;
 wire \system_integrator_b_output.input_bits[7] ;
 wire \system_integrator_b_output.input_bits[8] ;
 wire \system_integrator_b_output.output_bit ;
 wire \test_integrator_a_counter.value_output[0] ;
 wire \test_integrator_a_counter.value_output[1] ;
 wire \test_integrator_a_counter.value_output[2] ;
 wire \test_integrator_a_counter.value_output[3] ;
 wire \test_integrator_a_counter.value_output[4] ;
 wire \test_integrator_a_counter.value_output[5] ;
 wire \test_integrator_a_counter.value_output[6] ;
 wire \test_integrator_a_counter.value_output[7] ;
 wire \test_integrator_a_counter.value_output[8] ;
 wire \test_integrator_a_output.bitseq[0] ;
 wire \test_integrator_a_output.bitseq[1] ;
 wire \test_integrator_a_output.bitseq[2] ;
 wire \test_integrator_a_output.bitseq[3] ;
 wire \test_integrator_a_output.bitseq[4] ;
 wire \test_integrator_a_output.bitseq[5] ;
 wire \test_integrator_a_output.bitseq[6] ;
 wire \test_integrator_a_output.bitseq[7] ;
 wire \test_integrator_a_output.counter[0] ;
 wire \test_integrator_a_output.counter[1] ;
 wire \test_integrator_a_output.counter[2] ;
 wire \test_integrator_a_output.counter[3] ;
 wire \test_integrator_a_output.input_bits[0] ;
 wire \test_integrator_a_output.input_bits[1] ;
 wire \test_integrator_a_output.input_bits[2] ;
 wire \test_integrator_a_output.input_bits[3] ;
 wire \test_integrator_a_output.input_bits[4] ;
 wire \test_integrator_a_output.input_bits[5] ;
 wire \test_integrator_a_output.input_bits[6] ;
 wire \test_integrator_a_output.input_bits[7] ;
 wire \test_integrator_a_output.input_bits[8] ;
 wire \test_integrator_a_output.output_bit ;
 wire \test_integrator_b_counter.value_output[0] ;
 wire \test_integrator_b_counter.value_output[1] ;
 wire \test_integrator_b_counter.value_output[2] ;
 wire \test_integrator_b_counter.value_output[3] ;
 wire \test_integrator_b_counter.value_output[4] ;
 wire \test_integrator_b_counter.value_output[5] ;
 wire \test_integrator_b_counter.value_output[6] ;
 wire \test_integrator_b_counter.value_output[7] ;
 wire \test_integrator_b_counter.value_output[8] ;
 wire \test_integrator_b_output.bitseq[0] ;
 wire \test_integrator_b_output.bitseq[1] ;
 wire \test_integrator_b_output.bitseq[2] ;
 wire \test_integrator_b_output.bitseq[3] ;
 wire \test_integrator_b_output.bitseq[4] ;
 wire \test_integrator_b_output.bitseq[5] ;
 wire \test_integrator_b_output.bitseq[6] ;
 wire \test_integrator_b_output.bitseq[7] ;
 wire \test_integrator_b_output.counter[0] ;
 wire \test_integrator_b_output.counter[1] ;
 wire \test_integrator_b_output.counter[2] ;
 wire \test_integrator_b_output.counter[3] ;
 wire \test_integrator_b_output.input_bits[0] ;
 wire \test_integrator_b_output.input_bits[1] ;
 wire \test_integrator_b_output.input_bits[2] ;
 wire \test_integrator_b_output.input_bits[3] ;
 wire \test_integrator_b_output.input_bits[4] ;
 wire \test_integrator_b_output.input_bits[5] ;
 wire \test_integrator_b_output.input_bits[6] ;
 wire \test_integrator_b_output.input_bits[7] ;
 wire \test_integrator_b_output.input_bits[8] ;
 wire \test_integrator_b_output.output_bit ;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net1;
 wire net2;
 wire net3;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;

 sg13g2_inv_1 _1936_ (.Y(_1613_),
    .A(net325));
 sg13g2_inv_1 _1937_ (.Y(_1614_),
    .A(\input_b_sng_comparator.bits_a[0] ));
 sg13g2_inv_1 _1938_ (.Y(_1615_),
    .A(\input_a_sng_comparator.bits_a[0] ));
 sg13g2_inv_2 _1939_ (.Y(_1616_),
    .A(\test_integrator_a_counter.value_output[8] ));
 sg13g2_inv_2 _1940_ (.Y(_1617_),
    .A(net467));
 sg13g2_inv_1 _1941_ (.Y(_1618_),
    .A(net497));
 sg13g2_inv_1 _1942_ (.Y(_1619_),
    .A(net501));
 sg13g2_inv_2 _1943_ (.Y(_1620_),
    .A(net488));
 sg13g2_inv_2 _1944_ (.Y(_1621_),
    .A(net496));
 sg13g2_inv_2 _1945_ (.Y(_1622_),
    .A(net491));
 sg13g2_inv_1 _1946_ (.Y(_1623_),
    .A(\test_integrator_a_counter.value_output[1] ));
 sg13g2_inv_2 _1947_ (.Y(_1624_),
    .A(net470));
 sg13g2_inv_1 _1948_ (.Y(_1625_),
    .A(net500));
 sg13g2_inv_2 _1949_ (.Y(_1626_),
    .A(net486));
 sg13g2_inv_1 _1950_ (.Y(_1627_),
    .A(net502));
 sg13g2_inv_2 _1951_ (.Y(_1628_),
    .A(net472));
 sg13g2_inv_1 _1952_ (.Y(_1629_),
    .A(net503));
 sg13g2_inv_1 _1953_ (.Y(_1630_),
    .A(net478));
 sg13g2_inv_1 _1954_ (.Y(_1631_),
    .A(\system_integrator_a_counter.value_output[4] ));
 sg13g2_inv_2 _1955_ (.Y(_1632_),
    .A(net312));
 sg13g2_inv_2 _1956_ (.Y(_1633_),
    .A(\integrator_c_counter.value_output[7] ));
 sg13g2_inv_2 _1957_ (.Y(_1634_),
    .A(net473));
 sg13g2_inv_1 _1958_ (.Y(_1635_),
    .A(\integrator_c_counter.value_output[5] ));
 sg13g2_inv_1 _1959_ (.Y(_1636_),
    .A(\integrator_c_counter.value_output[4] ));
 sg13g2_inv_1 _1960_ (.Y(_1637_),
    .A(\integrator_c_counter.value_output[3] ));
 sg13g2_inv_2 _1961_ (.Y(_1638_),
    .A(net456));
 sg13g2_inv_1 _1962_ (.Y(_1639_),
    .A(\integrator_c_counter.value_output[1] ));
 sg13g2_inv_2 _1963_ (.Y(_1640_),
    .A(net391));
 sg13g2_inv_2 _1964_ (.Y(_1641_),
    .A(\integrator_b_counter.value_output[7] ));
 sg13g2_inv_1 _1965_ (.Y(_1642_),
    .A(\integrator_b_counter.value_output[4] ));
 sg13g2_inv_1 _1966_ (.Y(_1643_),
    .A(\integrator_b_counter.value_output[0] ));
 sg13g2_inv_1 _1967_ (.Y(_1644_),
    .A(\integrator_a_counter.value_output[7] ));
 sg13g2_inv_1 _1968_ (.Y(_1645_),
    .A(\integrator_a_counter.value_output[4] ));
 sg13g2_inv_2 _1969_ (.Y(_1646_),
    .A(\integrator_a_counter.value_output[0] ));
 sg13g2_inv_1 _1970_ (.Y(_1647_),
    .A(\test_integrator_b_counter.value_output[7] ));
 sg13g2_inv_1 _1971_ (.Y(_1648_),
    .A(\test_integrator_b_counter.value_output[4] ));
 sg13g2_inv_1 _1972_ (.Y(_1649_),
    .A(\test_integrator_b_counter.value_output[3] ));
 sg13g2_inv_1 _1973_ (.Y(_1650_),
    .A(net495));
 sg13g2_inv_1 _1974_ (.Y(_1651_),
    .A(net213));
 sg13g2_inv_1 _1975_ (.Y(_0124_),
    .A(net25));
 sg13g2_inv_1 _1976_ (.Y(_0122_),
    .A(net26));
 sg13g2_inv_1 _1977_ (.Y(_0120_),
    .A(net33));
 sg13g2_inv_1 _1978_ (.Y(_1652_),
    .A(\input_a_sng_comparator.bits_b[7] ));
 sg13g2_inv_1 _1979_ (.Y(_1653_),
    .A(net601));
 sg13g2_inv_1 _1980_ (.Y(_0111_),
    .A(net412));
 sg13g2_inv_1 _1981_ (.Y(_1654_),
    .A(net585));
 sg13g2_inv_1 _1982_ (.Y(_1655_),
    .A(\input_a_sng_comparator.bits_b[6] ));
 sg13g2_inv_1 _1983_ (.Y(_1656_),
    .A(net600));
 sg13g2_inv_1 _1984_ (.Y(_0633_),
    .A(net603));
 sg13g2_inv_1 _1985_ (.Y(_0634_),
    .A(\integrator_b_sng_comparator.bits_b[6] ));
 sg13g2_inv_1 _1986_ (.Y(_0635_),
    .A(net594));
 sg13g2_inv_1 _1987_ (.Y(_0636_),
    .A(_0050_));
 sg13g2_inv_1 _1988_ (.Y(_0637_),
    .A(\input_halfprob2_sng_comparator.bits_b[3] ));
 sg13g2_inv_1 _1989_ (.Y(_0638_),
    .A(\input_halfprob2_sng_comparator.bits_b[2] ));
 sg13g2_inv_1 _1990_ (.Y(_0639_),
    .A(\input_halfprob1_sng_comparator.bits_b[0] ));
 sg13g2_inv_1 _1991_ (.Y(_0640_),
    .A(\integrator_a_sng_comparator.bits_b[1] ));
 sg13g2_inv_2 _1992_ (.Y(_0641_),
    .A(\input_halfprob2_sng_comparator.bits_b[8] ));
 sg13g2_inv_1 _1993_ (.Y(_0642_),
    .A(net421));
 sg13g2_inv_1 _1994_ (.Y(_0643_),
    .A(net468));
 sg13g2_inv_1 _1995_ (.Y(_0644_),
    .A(net253));
 sg13g2_inv_1 _1996_ (.Y(_0645_),
    .A(\clk_counter[10] ));
 sg13g2_inv_1 _1997_ (.Y(_0646_),
    .A(net306));
 sg13g2_inv_1 _1998_ (.Y(_0647_),
    .A(\serial_input.adjustment[3] ));
 sg13g2_inv_1 _1999_ (.Y(_0000_),
    .A(net363));
 sg13g2_inv_1 _2000_ (.Y(_0648_),
    .A(net364));
 sg13g2_inv_1 _2001_ (.Y(_0004_),
    .A(net383));
 sg13g2_inv_1 _2002_ (.Y(_0649_),
    .A(net337));
 sg13g2_inv_1 _2003_ (.Y(_0008_),
    .A(net382));
 sg13g2_inv_1 _2004_ (.Y(_0650_),
    .A(net303));
 sg13g2_inv_1 _2005_ (.Y(_0013_),
    .A(net352));
 sg13g2_inv_1 _2006_ (.Y(_0651_),
    .A(net308));
 sg13g2_inv_1 _2007_ (.Y(_0017_),
    .A(net347));
 sg13g2_inv_1 _2008_ (.Y(_0652_),
    .A(net320));
 sg13g2_inv_1 _2009_ (.Y(_0653_),
    .A(\input_halfprob1_sng_comparator.bits_b[8] ));
 sg13g2_inv_1 _2010_ (.Y(_0021_),
    .A(net355));
 sg13g2_inv_1 _2011_ (.Y(_0654_),
    .A(net356));
 sg13g2_inv_1 _2012_ (.Y(_0025_),
    .A(net394));
 sg13g2_inv_1 _2013_ (.Y(_0655_),
    .A(net392));
 sg13g2_inv_1 _2014_ (.Y(_0656_),
    .A(_0034_));
 sg13g2_inv_1 _2015_ (.Y(_0657_),
    .A(_0036_));
 sg13g2_inv_1 _2016_ (.Y(_0658_),
    .A(net431));
 sg13g2_inv_1 _2017_ (.Y(_0659_),
    .A(_0047_));
 sg13g2_inv_1 _2018_ (.Y(_0660_),
    .A(_0048_));
 sg13g2_inv_1 _2019_ (.Y(_0087_),
    .A(net655));
 sg13g2_nor2_1 _2020_ (.A(\serial_input.adjustment[4] ),
    .B(_0643_),
    .Y(_0661_));
 sg13g2_nor2b_1 _2021_ (.A(\clk_counter[0] ),
    .B_N(\serial_input.adjustment[0] ),
    .Y(_0662_));
 sg13g2_nor2b_1 _2022_ (.A(\serial_input.adjustment[0] ),
    .B_N(\clk_counter[0] ),
    .Y(_0663_));
 sg13g2_xnor2_1 _2023_ (.Y(_0664_),
    .A(net213),
    .B(\clk_counter[2] ));
 sg13g2_nor2_1 _2024_ (.A(\clk_counter[3] ),
    .B(_0647_),
    .Y(_0665_));
 sg13g2_nor4_1 _2025_ (.A(net585),
    .B(_0661_),
    .C(_0662_),
    .D(_0665_),
    .Y(_0666_));
 sg13g2_xnor2_1 _2026_ (.Y(_0667_),
    .A(\serial_input.adjustment[1] ),
    .B(\clk_counter[1] ));
 sg13g2_a221oi_1 _2027_ (.B2(\clk_counter[3] ),
    .C1(_0663_),
    .B1(_0647_),
    .A1(\serial_input.adjustment[4] ),
    .Y(_0668_),
    .A2(_0643_));
 sg13g2_nand4_1 _2028_ (.B(_0666_),
    .C(_0667_),
    .A(_0664_),
    .Y(_0669_),
    .D(_0668_));
 sg13g2_nor2_1 _2029_ (.A(\serial_input.output_bitcounter_2[8] ),
    .B(net535),
    .Y(_0670_));
 sg13g2_a21oi_1 _2030_ (.A1(_1613_),
    .A2(net535),
    .Y(_0632_),
    .B1(_0670_));
 sg13g2_mux2_1 _2031_ (.A0(net327),
    .A1(net331),
    .S(net535),
    .X(_0631_));
 sg13g2_mux2_1 _2032_ (.A0(net348),
    .A1(\input_b_sng_comparator.bits_a[6] ),
    .S(net534),
    .X(_0630_));
 sg13g2_mux2_1 _2033_ (.A0(net358),
    .A1(\input_b_sng_comparator.bits_a[5] ),
    .S(net534),
    .X(_0629_));
 sg13g2_mux2_1 _2034_ (.A0(net313),
    .A1(\input_b_sng_comparator.bits_a[4] ),
    .S(net534),
    .X(_0628_));
 sg13g2_mux2_1 _2035_ (.A0(net360),
    .A1(net386),
    .S(net535),
    .X(_0627_));
 sg13g2_mux2_1 _2036_ (.A0(net258),
    .A1(\input_b_sng_comparator.bits_a[2] ),
    .S(net535),
    .X(_0626_));
 sg13g2_mux2_1 _2037_ (.A0(net284),
    .A1(\input_b_sng_comparator.bits_a[1] ),
    .S(net535),
    .X(_0625_));
 sg13g2_nor2_1 _2038_ (.A(net268),
    .B(net535),
    .Y(_0671_));
 sg13g2_a21oi_1 _2039_ (.A1(_1614_),
    .A2(_0669_),
    .Y(_0624_),
    .B1(_0671_));
 sg13g2_nand2_1 _2040_ (.Y(_0672_),
    .A(\integrator_b_output.counter[0] ),
    .B(net337));
 sg13g2_nor3_2 _2041_ (.A(\integrator_b_output.counter[1] ),
    .B(\integrator_b_output.counter[2] ),
    .C(_0672_),
    .Y(_0673_));
 sg13g2_nor4_2 _2042_ (.A(\integrator_b_output.counter[0] ),
    .B(\integrator_b_output.counter[1] ),
    .C(\integrator_b_output.counter[2] ),
    .Y(_0674_),
    .D(\integrator_b_output.counter[3] ));
 sg13g2_a22oi_1 _2043_ (.Y(_0675_),
    .B1(net580),
    .B2(net43),
    .A2(net549),
    .A1(\integrator_b_output.bitseq[7] ));
 sg13g2_inv_1 _2044_ (.Y(_0623_),
    .A(net44));
 sg13g2_nand2_1 _2045_ (.Y(_0676_),
    .A(net116),
    .B(net549));
 sg13g2_nand2b_1 _2046_ (.Y(_0677_),
    .B(net580),
    .A_N(\integrator_b_output.input_bits[7] ));
 sg13g2_o21ai_1 _2047_ (.B1(_0677_),
    .Y(_0678_),
    .A1(\integrator_b_output.bitseq[7] ),
    .A2(net580));
 sg13g2_o21ai_1 _2048_ (.B1(_0676_),
    .Y(_0622_),
    .A1(net549),
    .A2(_0678_));
 sg13g2_nand2_1 _2049_ (.Y(_0679_),
    .A(net80),
    .B(net549));
 sg13g2_nand2b_1 _2050_ (.Y(_0680_),
    .B(net580),
    .A_N(\integrator_b_output.input_bits[6] ));
 sg13g2_o21ai_1 _2051_ (.B1(_0680_),
    .Y(_0681_),
    .A1(\integrator_b_output.bitseq[6] ),
    .A2(net580));
 sg13g2_o21ai_1 _2052_ (.B1(_0679_),
    .Y(_0621_),
    .A1(net549),
    .A2(_0681_));
 sg13g2_nand2_1 _2053_ (.Y(_0682_),
    .A(net108),
    .B(net549));
 sg13g2_nand2b_1 _2054_ (.Y(_0683_),
    .B(net580),
    .A_N(\integrator_b_output.input_bits[5] ));
 sg13g2_o21ai_1 _2055_ (.B1(_0683_),
    .Y(_0684_),
    .A1(net80),
    .A2(net580));
 sg13g2_o21ai_1 _2056_ (.B1(_0682_),
    .Y(_0620_),
    .A1(net549),
    .A2(_0684_));
 sg13g2_nand2_1 _2057_ (.Y(_0685_),
    .A(net114),
    .B(net548));
 sg13g2_nand2b_1 _2058_ (.Y(_0686_),
    .B(net580),
    .A_N(\integrator_b_output.input_bits[4] ));
 sg13g2_o21ai_1 _2059_ (.B1(_0686_),
    .Y(_0687_),
    .A1(net108),
    .A2(net579));
 sg13g2_o21ai_1 _2060_ (.B1(_0685_),
    .Y(_0619_),
    .A1(net548),
    .A2(_0687_));
 sg13g2_nand2_1 _2061_ (.Y(_0688_),
    .A(net85),
    .B(_0673_));
 sg13g2_nand2b_1 _2062_ (.Y(_0689_),
    .B(net579),
    .A_N(\integrator_b_output.input_bits[3] ));
 sg13g2_o21ai_1 _2063_ (.B1(_0689_),
    .Y(_0690_),
    .A1(\integrator_b_output.bitseq[3] ),
    .A2(net579));
 sg13g2_o21ai_1 _2064_ (.B1(net86),
    .Y(_0618_),
    .A1(net548),
    .A2(_0690_));
 sg13g2_nand2_1 _2065_ (.Y(_0691_),
    .A(net128),
    .B(net548));
 sg13g2_nand2b_1 _2066_ (.Y(_0692_),
    .B(net579),
    .A_N(\integrator_b_output.input_bits[2] ));
 sg13g2_o21ai_1 _2067_ (.B1(_0692_),
    .Y(_0693_),
    .A1(net85),
    .A2(_0674_));
 sg13g2_o21ai_1 _2068_ (.B1(_0691_),
    .Y(_0617_),
    .A1(net548),
    .A2(_0693_));
 sg13g2_nand2_1 _2069_ (.Y(_0694_),
    .A(net176),
    .B(net548));
 sg13g2_nand2b_1 _2070_ (.Y(_0695_),
    .B(net579),
    .A_N(net146));
 sg13g2_o21ai_1 _2071_ (.B1(_0695_),
    .Y(_0696_),
    .A1(net128),
    .A2(net579));
 sg13g2_o21ai_1 _2072_ (.B1(_0694_),
    .Y(_0616_),
    .A1(net548),
    .A2(_0696_));
 sg13g2_mux2_1 _2073_ (.A0(net404),
    .A1(\input_a_sng_comparator.bits_a[8] ),
    .S(net533),
    .X(_0615_));
 sg13g2_mux2_1 _2074_ (.A0(net310),
    .A1(net409),
    .S(net533),
    .X(_0614_));
 sg13g2_mux2_1 _2075_ (.A0(net290),
    .A1(net324),
    .S(net533),
    .X(_0613_));
 sg13g2_mux2_1 _2076_ (.A0(net333),
    .A1(net351),
    .S(net533),
    .X(_0612_));
 sg13g2_mux2_1 _2077_ (.A0(net211),
    .A1(net242),
    .S(net534),
    .X(_0611_));
 sg13g2_mux2_1 _2078_ (.A0(net332),
    .A1(net370),
    .S(net534),
    .X(_0610_));
 sg13g2_mux2_1 _2079_ (.A0(net300),
    .A1(net350),
    .S(net533),
    .X(_0609_));
 sg13g2_mux2_1 _2080_ (.A0(net120),
    .A1(\input_a_sng_comparator.bits_a[1] ),
    .S(net533),
    .X(_0608_));
 sg13g2_nor2_1 _2081_ (.A(net59),
    .B(net533),
    .Y(_0697_));
 sg13g2_a21oi_1 _2082_ (.A1(_1615_),
    .A2(net533),
    .Y(_0607_),
    .B1(_0697_));
 sg13g2_nor4_2 _2083_ (.A(\clk_counter[1] ),
    .B(\clk_counter[0] ),
    .C(\clk_counter[3] ),
    .Y(_0698_),
    .D(\clk_counter[2] ));
 sg13g2_nor2_1 _2084_ (.A(net366),
    .B(net570),
    .Y(_0699_));
 sg13g2_a21oi_1 _2085_ (.A1(_1616_),
    .A2(net570),
    .Y(_0606_),
    .B1(_0699_));
 sg13g2_nor2_1 _2086_ (.A(net264),
    .B(net570),
    .Y(_0700_));
 sg13g2_a21oi_1 _2087_ (.A1(_1617_),
    .A2(net570),
    .Y(_0605_),
    .B1(_0700_));
 sg13g2_nor2_1 _2088_ (.A(net295),
    .B(net570),
    .Y(_0701_));
 sg13g2_a21oi_1 _2089_ (.A1(_1618_),
    .A2(net570),
    .Y(_0604_),
    .B1(_0701_));
 sg13g2_nor2_1 _2090_ (.A(net361),
    .B(net571),
    .Y(_0702_));
 sg13g2_a21oi_1 _2091_ (.A1(_1619_),
    .A2(net570),
    .Y(_0603_),
    .B1(_0702_));
 sg13g2_nor2_1 _2092_ (.A(net329),
    .B(net570),
    .Y(_0703_));
 sg13g2_a21oi_1 _2093_ (.A1(_1620_),
    .A2(net571),
    .Y(_0602_),
    .B1(_0703_));
 sg13g2_nor2_1 _2094_ (.A(net339),
    .B(net572),
    .Y(_0704_));
 sg13g2_a21oi_1 _2095_ (.A1(_1621_),
    .A2(net572),
    .Y(_0601_),
    .B1(_0704_));
 sg13g2_nor2_1 _2096_ (.A(net282),
    .B(net572),
    .Y(_0705_));
 sg13g2_a21oi_1 _2097_ (.A1(_1622_),
    .A2(net572),
    .Y(_0600_),
    .B1(_0705_));
 sg13g2_nor2_1 _2098_ (.A(net221),
    .B(net572),
    .Y(_0706_));
 sg13g2_a21oi_1 _2099_ (.A1(_1623_),
    .A2(net572),
    .Y(_0599_),
    .B1(_0706_));
 sg13g2_mux2_1 _2100_ (.A0(net49),
    .A1(net234),
    .S(net572),
    .X(_0598_));
 sg13g2_mux2_1 _2101_ (.A0(net39),
    .A1(net292),
    .S(net562),
    .X(_0597_));
 sg13g2_nor2_1 _2102_ (.A(net280),
    .B(net562),
    .Y(_0707_));
 sg13g2_a21oi_1 _2103_ (.A1(_1624_),
    .A2(net562),
    .Y(_0596_),
    .B1(_0707_));
 sg13g2_nor2_1 _2104_ (.A(net260),
    .B(net562),
    .Y(_0708_));
 sg13g2_a21oi_1 _2105_ (.A1(_1625_),
    .A2(net562),
    .Y(_0595_),
    .B1(_0708_));
 sg13g2_nor2_1 _2106_ (.A(net272),
    .B(net562),
    .Y(_0709_));
 sg13g2_a21oi_1 _2107_ (.A1(_1626_),
    .A2(net562),
    .Y(_0594_),
    .B1(_0709_));
 sg13g2_nor2_1 _2108_ (.A(net334),
    .B(net562),
    .Y(_0710_));
 sg13g2_a21oi_1 _2109_ (.A1(_1627_),
    .A2(net563),
    .Y(_0593_),
    .B1(_0710_));
 sg13g2_nor2_1 _2110_ (.A(net353),
    .B(net563),
    .Y(_0711_));
 sg13g2_a21oi_1 _2111_ (.A1(_1628_),
    .A2(net563),
    .Y(_0592_),
    .B1(_0711_));
 sg13g2_nor2_1 _2112_ (.A(net343),
    .B(net563),
    .Y(_0712_));
 sg13g2_a21oi_1 _2113_ (.A1(_1629_),
    .A2(net563),
    .Y(_0591_),
    .B1(_0712_));
 sg13g2_nor2_1 _2114_ (.A(net293),
    .B(net563),
    .Y(_0713_));
 sg13g2_a21oi_1 _2115_ (.A1(_1630_),
    .A2(net563),
    .Y(_0590_),
    .B1(_0713_));
 sg13g2_mux2_1 _2116_ (.A0(net286),
    .A1(\system_integrator_b_counter.value_output[0] ),
    .S(net563),
    .X(_0589_));
 sg13g2_mux2_1 _2117_ (.A0(net52),
    .A1(net257),
    .S(net575),
    .X(_0588_));
 sg13g2_mux2_1 _2118_ (.A0(net215),
    .A1(\system_integrator_a_counter.value_output[7] ),
    .S(net575),
    .X(_0587_));
 sg13g2_mux2_1 _2119_ (.A0(net288),
    .A1(\system_integrator_a_counter.value_output[6] ),
    .S(net575),
    .X(_0586_));
 sg13g2_mux2_1 _2120_ (.A0(net207),
    .A1(\system_integrator_a_counter.value_output[5] ),
    .S(net575),
    .X(_0585_));
 sg13g2_nor2_1 _2121_ (.A(net276),
    .B(net575),
    .Y(_0714_));
 sg13g2_a21oi_1 _2122_ (.A1(_1631_),
    .A2(net575),
    .Y(_0584_),
    .B1(_0714_));
 sg13g2_mux2_1 _2123_ (.A0(net246),
    .A1(\system_integrator_a_counter.value_output[3] ),
    .S(net571),
    .X(_0583_));
 sg13g2_mux2_1 _2124_ (.A0(net200),
    .A1(net588),
    .S(net571),
    .X(_0582_));
 sg13g2_mux2_1 _2125_ (.A0(net232),
    .A1(\system_integrator_a_counter.value_output[1] ),
    .S(net571),
    .X(_0581_));
 sg13g2_mux2_1 _2126_ (.A0(net239),
    .A1(net252),
    .S(net571),
    .X(_0580_));
 sg13g2_nor2_1 _2127_ (.A(net165),
    .B(net573),
    .Y(_0715_));
 sg13g2_a21oi_1 _2128_ (.A1(_1632_),
    .A2(net573),
    .Y(_0579_),
    .B1(_0715_));
 sg13g2_nor2_1 _2129_ (.A(net255),
    .B(net573),
    .Y(_0716_));
 sg13g2_a21oi_1 _2130_ (.A1(_1633_),
    .A2(net574),
    .Y(_0578_),
    .B1(_0716_));
 sg13g2_nor2_1 _2131_ (.A(net322),
    .B(net573),
    .Y(_0717_));
 sg13g2_a21oi_1 _2132_ (.A1(_1634_),
    .A2(net572),
    .Y(_0577_),
    .B1(_0717_));
 sg13g2_nor2_1 _2133_ (.A(net315),
    .B(net577),
    .Y(_0718_));
 sg13g2_a21oi_1 _2134_ (.A1(_1635_),
    .A2(net574),
    .Y(_0576_),
    .B1(_0718_));
 sg13g2_nor2_1 _2135_ (.A(net345),
    .B(net577),
    .Y(_0719_));
 sg13g2_a21oi_1 _2136_ (.A1(_1636_),
    .A2(net576),
    .Y(_0575_),
    .B1(_0719_));
 sg13g2_nor2_1 _2137_ (.A(net278),
    .B(net576),
    .Y(_0720_));
 sg13g2_a21oi_1 _2138_ (.A1(_1637_),
    .A2(net576),
    .Y(_0574_),
    .B1(_0720_));
 sg13g2_nor2_1 _2139_ (.A(net167),
    .B(net576),
    .Y(_0721_));
 sg13g2_a21oi_1 _2140_ (.A1(_1638_),
    .A2(net577),
    .Y(_0573_),
    .B1(_0721_));
 sg13g2_nor2_1 _2141_ (.A(net266),
    .B(net576),
    .Y(_0722_));
 sg13g2_a21oi_1 _2142_ (.A1(_1639_),
    .A2(net576),
    .Y(_0572_),
    .B1(_0722_));
 sg13g2_nor2_1 _2143_ (.A(net172),
    .B(net576),
    .Y(_0723_));
 sg13g2_a21oi_1 _2144_ (.A1(_1640_),
    .A2(net576),
    .Y(_0571_),
    .B1(_0723_));
 sg13g2_mux2_1 _2145_ (.A0(net43),
    .A1(net231),
    .S(net568),
    .X(_0570_));
 sg13g2_nor2_1 _2146_ (.A(net118),
    .B(net568),
    .Y(_0724_));
 sg13g2_a21oi_1 _2147_ (.A1(_1641_),
    .A2(net568),
    .Y(_0569_),
    .B1(_0724_));
 sg13g2_mux2_1 _2148_ (.A0(net132),
    .A1(net589),
    .S(net568),
    .X(_0568_));
 sg13g2_mux2_1 _2149_ (.A0(net182),
    .A1(\integrator_b_counter.value_output[5] ),
    .S(net569),
    .X(_0567_));
 sg13g2_nor2_1 _2150_ (.A(net179),
    .B(net578),
    .Y(_0725_));
 sg13g2_a21oi_1 _2151_ (.A1(_1642_),
    .A2(net569),
    .Y(_0566_),
    .B1(net180));
 sg13g2_mux2_1 _2152_ (.A0(net192),
    .A1(\integrator_b_counter.value_output[3] ),
    .S(net569),
    .X(_0565_));
 sg13g2_mux2_1 _2153_ (.A0(net198),
    .A1(\integrator_b_counter.value_output[2] ),
    .S(net569),
    .X(_0564_));
 sg13g2_mux2_1 _2154_ (.A0(net146),
    .A1(\integrator_b_counter.value_output[1] ),
    .S(net569),
    .X(_0563_));
 sg13g2_nor2_1 _2155_ (.A(net219),
    .B(net569),
    .Y(_0726_));
 sg13g2_a21oi_1 _2156_ (.A1(_1643_),
    .A2(net569),
    .Y(_0562_),
    .B1(_0726_));
 sg13g2_mux2_1 _2157_ (.A0(net54),
    .A1(net243),
    .S(net565),
    .X(_0561_));
 sg13g2_nor2_1 _2158_ (.A(net262),
    .B(net565),
    .Y(_0727_));
 sg13g2_a21oi_1 _2159_ (.A1(_1644_),
    .A2(net565),
    .Y(_0560_),
    .B1(_0727_));
 sg13g2_mux2_1 _2160_ (.A0(net194),
    .A1(net590),
    .S(net564),
    .X(_0559_));
 sg13g2_mux2_1 _2161_ (.A0(net248),
    .A1(\integrator_a_counter.value_output[5] ),
    .S(net564),
    .X(_0558_));
 sg13g2_nor2_1 _2162_ (.A(net156),
    .B(net564),
    .Y(_0728_));
 sg13g2_a21oi_1 _2163_ (.A1(_1645_),
    .A2(net564),
    .Y(_0557_),
    .B1(_0728_));
 sg13g2_mux2_1 _2164_ (.A0(net274),
    .A1(\integrator_a_counter.value_output[3] ),
    .S(net564),
    .X(_0556_));
 sg13g2_mux2_1 _2165_ (.A0(net196),
    .A1(\integrator_a_counter.value_output[2] ),
    .S(net565),
    .X(_0555_));
 sg13g2_mux2_1 _2166_ (.A0(net202),
    .A1(\integrator_a_counter.value_output[1] ),
    .S(net565),
    .X(_0554_));
 sg13g2_nor2_1 _2167_ (.A(net341),
    .B(net565),
    .Y(_0729_));
 sg13g2_a21oi_1 _2168_ (.A1(_1646_),
    .A2(net565),
    .Y(_0553_),
    .B1(_0729_));
 sg13g2_nand2_1 _2169_ (.Y(_0730_),
    .A(net355),
    .B(net356));
 sg13g2_nor3_2 _2170_ (.A(\test_integrator_a_output.counter[1] ),
    .B(\test_integrator_a_output.counter[2] ),
    .C(_0730_),
    .Y(_0731_));
 sg13g2_nor4_2 _2171_ (.A(\test_integrator_a_output.counter[0] ),
    .B(\test_integrator_a_output.counter[1] ),
    .C(\test_integrator_a_output.counter[2] ),
    .Y(_0732_),
    .D(\test_integrator_a_output.counter[3] ));
 sg13g2_a22oi_1 _2172_ (.Y(_0733_),
    .B1(net560),
    .B2(\test_integrator_a_output.input_bits[8] ),
    .A2(net546),
    .A1(net229));
 sg13g2_inv_1 _2173_ (.Y(_0552_),
    .A(net230));
 sg13g2_nand2_1 _2174_ (.Y(_0734_),
    .A(net237),
    .B(net546));
 sg13g2_nand2b_1 _2175_ (.Y(_0735_),
    .B(net560),
    .A_N(\test_integrator_a_output.input_bits[7] ));
 sg13g2_o21ai_1 _2176_ (.B1(_0735_),
    .Y(_0736_),
    .A1(net229),
    .A2(net560));
 sg13g2_o21ai_1 _2177_ (.B1(_0734_),
    .Y(_0551_),
    .A1(net546),
    .A2(_0736_));
 sg13g2_nand2_1 _2178_ (.Y(_0737_),
    .A(net130),
    .B(net546));
 sg13g2_nand2b_1 _2179_ (.Y(_0738_),
    .B(net560),
    .A_N(\test_integrator_a_output.input_bits[6] ));
 sg13g2_o21ai_1 _2180_ (.B1(_0738_),
    .Y(_0739_),
    .A1(\test_integrator_a_output.bitseq[6] ),
    .A2(net560));
 sg13g2_o21ai_1 _2181_ (.B1(_0737_),
    .Y(_0550_),
    .A1(net546),
    .A2(_0739_));
 sg13g2_nand2_1 _2182_ (.Y(_0740_),
    .A(net150),
    .B(net546));
 sg13g2_nand2b_1 _2183_ (.Y(_0741_),
    .B(net560),
    .A_N(\test_integrator_a_output.input_bits[5] ));
 sg13g2_o21ai_1 _2184_ (.B1(_0741_),
    .Y(_0742_),
    .A1(net130),
    .A2(net561));
 sg13g2_o21ai_1 _2185_ (.B1(_0740_),
    .Y(_0549_),
    .A1(net546),
    .A2(_0742_));
 sg13g2_nand2_1 _2186_ (.Y(_0743_),
    .A(net67),
    .B(net547));
 sg13g2_nand2b_1 _2187_ (.Y(_0744_),
    .B(net561),
    .A_N(\test_integrator_a_output.input_bits[4] ));
 sg13g2_o21ai_1 _2188_ (.B1(_0744_),
    .Y(_0745_),
    .A1(\test_integrator_a_output.bitseq[4] ),
    .A2(net560));
 sg13g2_o21ai_1 _2189_ (.B1(_0743_),
    .Y(_0548_),
    .A1(net547),
    .A2(_0745_));
 sg13g2_nand2_1 _2190_ (.Y(_0746_),
    .A(net88),
    .B(_0731_));
 sg13g2_nand2b_1 _2191_ (.Y(_0747_),
    .B(_0732_),
    .A_N(\test_integrator_a_output.input_bits[3] ));
 sg13g2_o21ai_1 _2192_ (.B1(_0747_),
    .Y(_0748_),
    .A1(net67),
    .A2(net560));
 sg13g2_o21ai_1 _2193_ (.B1(net89),
    .Y(_0547_),
    .A1(net547),
    .A2(_0748_));
 sg13g2_nand2_1 _2194_ (.Y(_0749_),
    .A(net154),
    .B(net547));
 sg13g2_nand2b_1 _2195_ (.Y(_0750_),
    .B(_0732_),
    .A_N(\test_integrator_a_output.input_bits[2] ));
 sg13g2_o21ai_1 _2196_ (.B1(_0750_),
    .Y(_0751_),
    .A1(net88),
    .A2(net561));
 sg13g2_o21ai_1 _2197_ (.B1(_0749_),
    .Y(_0546_),
    .A1(net547),
    .A2(_0751_));
 sg13g2_nand2_1 _2198_ (.Y(_0752_),
    .A(net244),
    .B(net547));
 sg13g2_nand2b_1 _2199_ (.Y(_0753_),
    .B(net561),
    .A_N(net221));
 sg13g2_o21ai_1 _2200_ (.B1(_0753_),
    .Y(_0754_),
    .A1(net154),
    .A2(net561));
 sg13g2_o21ai_1 _2201_ (.B1(_0752_),
    .Y(_0545_),
    .A1(_0731_),
    .A2(_0754_));
 sg13g2_nor2b_1 _2202_ (.A(net597),
    .B_N(\input_a_sng_comparator.bits_a[6] ),
    .Y(_0755_));
 sg13g2_a21oi_1 _2203_ (.A1(\input_a_sng_comparator.bits_a[7] ),
    .A2(_1652_),
    .Y(_0756_),
    .B1(_0755_));
 sg13g2_a21o_1 _2204_ (.A2(_1652_),
    .A1(\input_a_sng_comparator.bits_a[7] ),
    .B1(_0755_),
    .X(_0757_));
 sg13g2_nor2b_1 _2205_ (.A(\input_a_sng_comparator.bits_a[5] ),
    .B_N(net598),
    .Y(_0758_));
 sg13g2_nor2b_1 _2206_ (.A(\input_a_sng_comparator.bits_a[7] ),
    .B_N(\input_a_sng_comparator.bits_b[7] ),
    .Y(_0759_));
 sg13g2_nor2b_1 _2207_ (.A(\input_a_sng_comparator.bits_a[6] ),
    .B_N(net597),
    .Y(_0760_));
 sg13g2_or3_1 _2208_ (.A(_0758_),
    .B(_0759_),
    .C(_0760_),
    .X(_0761_));
 sg13g2_nor2_1 _2209_ (.A(_0757_),
    .B(_0761_),
    .Y(_0762_));
 sg13g2_nor2b_1 _2210_ (.A(net598),
    .B_N(\input_a_sng_comparator.bits_a[5] ),
    .Y(_0763_));
 sg13g2_a21o_1 _2211_ (.A2(_1656_),
    .A1(\input_a_sng_comparator.bits_a[4] ),
    .B1(_0763_),
    .X(_0764_));
 sg13g2_nor2_1 _2212_ (.A(\input_a_sng_comparator.bits_a[4] ),
    .B(_1656_),
    .Y(_0765_));
 sg13g2_nor4_1 _2213_ (.A(_0757_),
    .B(_0761_),
    .C(_0764_),
    .D(_0765_),
    .Y(_0766_));
 sg13g2_nor2b_1 _2214_ (.A(net602),
    .B_N(\input_a_sng_comparator.bits_a[2] ),
    .Y(_0767_));
 sg13g2_nor2b_1 _2215_ (.A(\input_a_sng_comparator.bits_b[3] ),
    .B_N(\input_a_sng_comparator.bits_a[3] ),
    .Y(_0768_));
 sg13g2_nor2b_1 _2216_ (.A(\input_a_sng_comparator.bits_a[3] ),
    .B_N(\input_a_sng_comparator.bits_b[3] ),
    .Y(_0769_));
 sg13g2_nand2b_1 _2217_ (.Y(_0770_),
    .B(net601),
    .A_N(\input_a_sng_comparator.bits_a[3] ));
 sg13g2_nor2b_1 _2218_ (.A(\input_a_sng_comparator.bits_a[2] ),
    .B_N(net602),
    .Y(_0771_));
 sg13g2_or4_1 _2219_ (.A(_0767_),
    .B(_0768_),
    .C(_0769_),
    .D(_0771_),
    .X(_0772_));
 sg13g2_nor2b_1 _2220_ (.A(\input_a_sng_comparator.bits_b[1] ),
    .B_N(\input_a_sng_comparator.bits_a[1] ),
    .Y(_0773_));
 sg13g2_nand2b_1 _2221_ (.Y(_0774_),
    .B(net603),
    .A_N(\input_a_sng_comparator.bits_a[1] ));
 sg13g2_nand2b_1 _2222_ (.Y(_0775_),
    .B(\input_a_sng_comparator.bits_b[0] ),
    .A_N(\input_a_sng_comparator.bits_a[0] ));
 sg13g2_nand2_1 _2223_ (.Y(_0776_),
    .A(_0774_),
    .B(_0775_));
 sg13g2_a21oi_1 _2224_ (.A1(_0774_),
    .A2(_0775_),
    .Y(_0777_),
    .B1(_0773_));
 sg13g2_o21ai_1 _2225_ (.B1(_0770_),
    .Y(_0778_),
    .A1(_0767_),
    .A2(_0768_));
 sg13g2_o21ai_1 _2226_ (.B1(_0778_),
    .Y(_0779_),
    .A1(_0772_),
    .A2(_0777_));
 sg13g2_nand2b_1 _2227_ (.Y(_0780_),
    .B(\input_a_sng_comparator.bits_a[8] ),
    .A_N(\input_a_sng_comparator.bits_b[8] ));
 sg13g2_o21ai_1 _2228_ (.B1(_0780_),
    .Y(_0781_),
    .A1(_0756_),
    .A2(_0759_));
 sg13g2_a221oi_1 _2229_ (.B2(_0779_),
    .C1(_0781_),
    .B1(_0766_),
    .A1(_0762_),
    .Y(_0782_),
    .A2(_0764_));
 sg13g2_o21ai_1 _2230_ (.B1(_0780_),
    .Y(_0783_),
    .A1(_1615_),
    .A2(\input_a_sng_comparator.bits_b[0] ));
 sg13g2_nor4_1 _2231_ (.A(_0772_),
    .B(_0773_),
    .C(_0776_),
    .D(_0783_),
    .Y(_0784_));
 sg13g2_nor2_1 _2232_ (.A(\input_a_sng_comparator.bits_a[8] ),
    .B(_0120_),
    .Y(_0785_));
 sg13g2_a21o_1 _2233_ (.A2(_0784_),
    .A1(_0766_),
    .B1(_0785_),
    .X(_0786_));
 sg13g2_or2_2 _2234_ (.X(_0787_),
    .B(_0786_),
    .A(_0782_));
 sg13g2_nand2b_1 _2235_ (.Y(_0788_),
    .B(\test_integrator_b_counter.value_output[6] ),
    .A_N(\integrator_b_sng_comparator.bits_b[6] ));
 sg13g2_o21ai_1 _2236_ (.B1(_0788_),
    .Y(_0789_),
    .A1(_1647_),
    .A2(net596));
 sg13g2_nand2b_1 _2237_ (.Y(_0790_),
    .B(\integrator_b_sng_comparator.bits_b[6] ),
    .A_N(\test_integrator_b_counter.value_output[6] ));
 sg13g2_nand2b_1 _2238_ (.Y(_0791_),
    .B(net596),
    .A_N(\test_integrator_b_counter.value_output[7] ));
 sg13g2_nand2b_1 _2239_ (.Y(_0792_),
    .B(net597),
    .A_N(\test_integrator_b_counter.value_output[5] ));
 sg13g2_nand3_1 _2240_ (.B(_0791_),
    .C(_0792_),
    .A(_0790_),
    .Y(_0793_));
 sg13g2_nor2_1 _2241_ (.A(_0789_),
    .B(_0793_),
    .Y(_0794_));
 sg13g2_nand2b_1 _2242_ (.Y(_0795_),
    .B(\test_integrator_b_counter.value_output[5] ),
    .A_N(net597));
 sg13g2_o21ai_1 _2243_ (.B1(_0795_),
    .Y(_0796_),
    .A1(_1648_),
    .A2(net598));
 sg13g2_nor2b_1 _2244_ (.A(\test_integrator_b_counter.value_output[4] ),
    .B_N(net598),
    .Y(_0797_));
 sg13g2_nand2b_1 _2245_ (.Y(_0798_),
    .B(net599),
    .A_N(\test_integrator_b_counter.value_output[3] ));
 sg13g2_nand2b_1 _2246_ (.Y(_0799_),
    .B(_0798_),
    .A_N(_0797_));
 sg13g2_or4_1 _2247_ (.A(_0789_),
    .B(_0793_),
    .C(_0796_),
    .D(_0797_),
    .X(_0800_));
 sg13g2_nor4_1 _2248_ (.A(_0789_),
    .B(_0793_),
    .C(_0796_),
    .D(_0799_),
    .Y(_0801_));
 sg13g2_a22oi_1 _2249_ (.Y(_0802_),
    .B1(_1656_),
    .B2(\test_integrator_b_counter.value_output[3] ),
    .A2(_1653_),
    .A1(\test_integrator_b_counter.value_output[2] ));
 sg13g2_nor2b_1 _2250_ (.A(net602),
    .B_N(net592),
    .Y(_0803_));
 sg13g2_nand2b_1 _2251_ (.Y(_0804_),
    .B(net601),
    .A_N(net591));
 sg13g2_inv_1 _2252_ (.Y(_0805_),
    .A(_0804_));
 sg13g2_xnor2_1 _2253_ (.Y(_0806_),
    .A(net592),
    .B(net602));
 sg13g2_nand2b_1 _2254_ (.Y(_0807_),
    .B(net603),
    .A_N(\test_integrator_b_counter.value_output[0] ));
 sg13g2_nor2b_1 _2255_ (.A(\integrator_b_sng_comparator.bits_b[8] ),
    .B_N(\test_integrator_b_counter.value_output[8] ),
    .Y(_0808_));
 sg13g2_a21o_1 _2256_ (.A2(_0791_),
    .A1(_0789_),
    .B1(_0808_),
    .X(_0809_));
 sg13g2_and2_1 _2257_ (.A(_0806_),
    .B(_0807_),
    .X(_0810_));
 sg13g2_a21oi_1 _2258_ (.A1(_0806_),
    .A2(_0807_),
    .Y(_0811_),
    .B1(_0803_));
 sg13g2_o21ai_1 _2259_ (.B1(_0802_),
    .Y(_0812_),
    .A1(_0805_),
    .A2(_0811_));
 sg13g2_and2_1 _2260_ (.A(_0798_),
    .B(_0804_),
    .X(_0813_));
 sg13g2_a221oi_1 _2261_ (.B2(_0812_),
    .C1(_0809_),
    .B1(_0801_),
    .A1(_0794_),
    .Y(_0814_),
    .A2(_0796_));
 sg13g2_a21oi_1 _2262_ (.A1(\test_integrator_b_counter.value_output[0] ),
    .A2(_0633_),
    .Y(_0815_),
    .B1(_0808_));
 sg13g2_nand4_1 _2263_ (.B(_0810_),
    .C(_0813_),
    .A(_0802_),
    .Y(_0816_),
    .D(_0815_));
 sg13g2_nand2b_1 _2264_ (.Y(_0817_),
    .B(\integrator_b_sng_comparator.bits_b[8] ),
    .A_N(\test_integrator_b_counter.value_output[8] ));
 sg13g2_o21ai_1 _2265_ (.B1(_0817_),
    .Y(_0818_),
    .A1(_0800_),
    .A2(_0816_));
 sg13g2_nor2_2 _2266_ (.A(_0814_),
    .B(_0818_),
    .Y(_0819_));
 sg13g2_nor4_1 _2267_ (.A(_0782_),
    .B(_0786_),
    .C(_0814_),
    .D(_0818_),
    .Y(_0820_));
 sg13g2_nor4_1 _2268_ (.A(\test_integrator_a_counter.value_output[7] ),
    .B(\test_integrator_a_counter.value_output[6] ),
    .C(\test_integrator_a_counter.value_output[5] ),
    .D(\test_integrator_a_counter.value_output[4] ),
    .Y(_0821_));
 sg13g2_nor4_1 _2269_ (.A(\test_integrator_a_counter.value_output[2] ),
    .B(\test_integrator_a_counter.value_output[1] ),
    .C(\test_integrator_a_counter.value_output[0] ),
    .D(net594),
    .Y(_0822_));
 sg13g2_nand4_1 _2270_ (.B(_1621_),
    .C(_0821_),
    .A(_1616_),
    .Y(_0823_),
    .D(_0822_));
 sg13g2_nand4_1 _2271_ (.B(\test_integrator_a_counter.value_output[0] ),
    .C(net582),
    .A(\test_integrator_a_counter.value_output[1] ),
    .Y(_0824_),
    .D(_0636_));
 sg13g2_nand4_1 _2272_ (.B(\test_integrator_a_counter.value_output[6] ),
    .C(\test_integrator_a_counter.value_output[5] ),
    .A(\test_integrator_a_counter.value_output[7] ),
    .Y(_0825_),
    .D(\test_integrator_a_counter.value_output[2] ));
 sg13g2_nor4_1 _2273_ (.A(_1620_),
    .B(_1621_),
    .C(_0824_),
    .D(_0825_),
    .Y(_0826_));
 sg13g2_nor2_1 _2274_ (.A(_0819_),
    .B(_0826_),
    .Y(_0827_));
 sg13g2_a22oi_1 _2275_ (.Y(_0828_),
    .B1(_0827_),
    .B2(_0787_),
    .A2(_0823_),
    .A1(net532));
 sg13g2_xnor2_1 _2276_ (.Y(_0829_),
    .A(\test_integrator_a_counter.value_output[4] ),
    .B(net530));
 sg13g2_nor2_2 _2277_ (.A(\test_integrator_a_counter.value_output[3] ),
    .B(net530),
    .Y(_0830_));
 sg13g2_and2_1 _2278_ (.A(\test_integrator_a_counter.value_output[3] ),
    .B(net530),
    .X(_0831_));
 sg13g2_and2_1 _2279_ (.A(\test_integrator_a_counter.value_output[2] ),
    .B(net531),
    .X(_0832_));
 sg13g2_xnor2_1 _2280_ (.Y(_0833_),
    .A(\test_integrator_a_counter.value_output[2] ),
    .B(net530));
 sg13g2_nor2_1 _2281_ (.A(_0656_),
    .B(net531),
    .Y(_0834_));
 sg13g2_a21oi_1 _2282_ (.A1(_0656_),
    .A2(net531),
    .Y(_0835_),
    .B1(\test_integrator_a_counter.value_output[0] ));
 sg13g2_nor3_2 _2283_ (.A(_0833_),
    .B(_0834_),
    .C(_0835_),
    .Y(_0836_));
 sg13g2_nor2_1 _2284_ (.A(_0832_),
    .B(_0836_),
    .Y(_0837_));
 sg13g2_nor3_2 _2285_ (.A(_0831_),
    .B(_0832_),
    .C(_0836_),
    .Y(_0838_));
 sg13g2_nor3_1 _2286_ (.A(_0829_),
    .B(_0830_),
    .C(_0838_),
    .Y(_0839_));
 sg13g2_xnor2_1 _2287_ (.Y(_0840_),
    .A(\test_integrator_a_counter.value_output[5] ),
    .B(net530));
 sg13g2_nor4_2 _2288_ (.A(_0829_),
    .B(_0830_),
    .C(_0838_),
    .Y(_0841_),
    .D(_0840_));
 sg13g2_nor2_1 _2289_ (.A(\test_integrator_a_counter.value_output[6] ),
    .B(net532),
    .Y(_0842_));
 sg13g2_nand2_1 _2290_ (.Y(_0843_),
    .A(\test_integrator_a_counter.value_output[6] ),
    .B(net532));
 sg13g2_nor2b_1 _2291_ (.A(_0842_),
    .B_N(_0843_),
    .Y(_0844_));
 sg13g2_xnor2_1 _2292_ (.Y(_0845_),
    .A(_1617_),
    .B(net532));
 sg13g2_nand3_1 _2293_ (.B(_0844_),
    .C(_0845_),
    .A(_0841_),
    .Y(_0846_));
 sg13g2_nand2_1 _2294_ (.Y(_0847_),
    .A(net532),
    .B(_0821_));
 sg13g2_mux2_1 _2295_ (.A0(net532),
    .A1(_0847_),
    .S(_0846_),
    .X(_0848_));
 sg13g2_nand2b_1 _2296_ (.Y(_0849_),
    .B(net374),
    .A_N(_0848_));
 sg13g2_nand2b_1 _2297_ (.Y(_0850_),
    .B(_0848_),
    .A_N(net374));
 sg13g2_nor2_2 _2298_ (.A(net594),
    .B(net519),
    .Y(_0851_));
 sg13g2_and2_1 _2299_ (.A(_0849_),
    .B(_0851_),
    .X(_0852_));
 sg13g2_a22oi_1 _2300_ (.Y(_0544_),
    .B1(_0850_),
    .B2(_0852_),
    .A2(net519),
    .A1(_1616_));
 sg13g2_o21ai_1 _2301_ (.B1(net530),
    .Y(_0853_),
    .A1(\test_integrator_a_counter.value_output[5] ),
    .A2(\test_integrator_a_counter.value_output[4] ));
 sg13g2_nor2b_1 _2302_ (.A(_0841_),
    .B_N(_0853_),
    .Y(_0854_));
 sg13g2_o21ai_1 _2303_ (.B1(_0843_),
    .Y(_0855_),
    .A1(_0842_),
    .A2(_0854_));
 sg13g2_xnor2_1 _2304_ (.Y(_0856_),
    .A(_0845_),
    .B(_0855_));
 sg13g2_a22oi_1 _2305_ (.Y(_0543_),
    .B1(_0851_),
    .B2(_0856_),
    .A2(net519),
    .A1(_1617_));
 sg13g2_xor2_1 _2306_ (.B(_0854_),
    .A(_0844_),
    .X(_0857_));
 sg13g2_a22oi_1 _2307_ (.Y(_0542_),
    .B1(_0851_),
    .B2(_0857_),
    .A2(net519),
    .A1(_1618_));
 sg13g2_a21oi_1 _2308_ (.A1(\test_integrator_a_counter.value_output[4] ),
    .A2(net530),
    .Y(_0858_),
    .B1(_0839_));
 sg13g2_xnor2_1 _2309_ (.Y(_0859_),
    .A(_0840_),
    .B(_0858_));
 sg13g2_a22oi_1 _2310_ (.Y(_0541_),
    .B1(_0851_),
    .B2(_0859_),
    .A2(_0828_),
    .A1(_1619_));
 sg13g2_o21ai_1 _2311_ (.B1(_0829_),
    .Y(_0860_),
    .A1(_0830_),
    .A2(_0838_));
 sg13g2_nand2b_1 _2312_ (.Y(_0861_),
    .B(_0860_),
    .A_N(_0839_));
 sg13g2_a22oi_1 _2313_ (.Y(_0540_),
    .B1(_0851_),
    .B2(_0861_),
    .A2(net519),
    .A1(_1620_));
 sg13g2_or2_1 _2314_ (.X(_0862_),
    .B(_0831_),
    .A(_0830_));
 sg13g2_xnor2_1 _2315_ (.Y(_0863_),
    .A(_0837_),
    .B(_0862_));
 sg13g2_a22oi_1 _2316_ (.Y(_0539_),
    .B1(_0851_),
    .B2(_0863_),
    .A2(net519),
    .A1(_1621_));
 sg13g2_o21ai_1 _2317_ (.B1(_0833_),
    .Y(_0864_),
    .A1(_0834_),
    .A2(_0835_));
 sg13g2_nand2b_1 _2318_ (.Y(_0865_),
    .B(_0864_),
    .A_N(_0836_));
 sg13g2_a22oi_1 _2319_ (.Y(_0538_),
    .B1(_0851_),
    .B2(_0865_),
    .A2(net519),
    .A1(_1622_));
 sg13g2_xnor2_1 _2320_ (.Y(_0866_),
    .A(_0034_),
    .B(net531));
 sg13g2_xor2_1 _2321_ (.B(_0866_),
    .A(net417),
    .X(_0867_));
 sg13g2_a22oi_1 _2322_ (.Y(_0537_),
    .B1(_0851_),
    .B2(net418),
    .A2(net519),
    .A1(_1623_));
 sg13g2_nand2_1 _2323_ (.Y(_0868_),
    .A(net582),
    .B(net417));
 sg13g2_o21ai_1 _2324_ (.B1(_0868_),
    .Y(_0869_),
    .A1(net582),
    .A2(net530));
 sg13g2_mux2_1 _2325_ (.A0(_0869_),
    .A1(net234),
    .S(_0828_),
    .X(_0536_));
 sg13g2_nand2b_1 _2326_ (.Y(_0870_),
    .B(\system_integrator_a_counter.value_output[6] ),
    .A_N(\input_halfprob2_sng_comparator.bits_b[3] ));
 sg13g2_nand2b_1 _2327_ (.Y(_0871_),
    .B(\system_integrator_a_counter.value_output[7] ),
    .A_N(\input_halfprob2_sng_comparator.bits_b[4] ));
 sg13g2_nand2_1 _2328_ (.Y(_0872_),
    .A(_0870_),
    .B(_0871_));
 sg13g2_nand2b_1 _2329_ (.Y(_0873_),
    .B(\input_halfprob2_sng_comparator.bits_b[4] ),
    .A_N(\system_integrator_a_counter.value_output[7] ));
 sg13g2_nand2b_1 _2330_ (.Y(_0874_),
    .B(\input_halfprob2_sng_comparator.bits_b[3] ),
    .A_N(\system_integrator_a_counter.value_output[6] ));
 sg13g2_and4_1 _2331_ (.A(_0870_),
    .B(_0871_),
    .C(_0873_),
    .D(_0874_),
    .X(_0875_));
 sg13g2_nand2b_1 _2332_ (.Y(_0876_),
    .B(\system_integrator_a_counter.value_output[5] ),
    .A_N(\input_halfprob2_sng_comparator.bits_b[2] ));
 sg13g2_nand2b_1 _2333_ (.Y(_0877_),
    .B(\system_integrator_a_counter.value_output[4] ),
    .A_N(\input_halfprob2_sng_comparator.bits_b[1] ));
 sg13g2_nor2b_1 _2334_ (.A(\system_integrator_a_counter.value_output[5] ),
    .B_N(\input_halfprob2_sng_comparator.bits_b[2] ),
    .Y(_0878_));
 sg13g2_a21oi_1 _2335_ (.A1(_1631_),
    .A2(\input_halfprob2_sng_comparator.bits_b[1] ),
    .Y(_0879_),
    .B1(_0878_));
 sg13g2_nand4_1 _2336_ (.B(_0876_),
    .C(_0877_),
    .A(_0875_),
    .Y(_0880_),
    .D(_0879_));
 sg13g2_nand2b_1 _2337_ (.Y(_0881_),
    .B(\system_integrator_a_counter.value_output[2] ),
    .A_N(\input_halfprob1_sng_comparator.bits_b[0] ));
 sg13g2_nand2b_1 _2338_ (.Y(_0882_),
    .B(\system_integrator_a_counter.value_output[3] ),
    .A_N(\input_halfprob1_sng_comparator.bits_b[1] ));
 sg13g2_nand2_1 _2339_ (.Y(_0883_),
    .A(_0881_),
    .B(_0882_));
 sg13g2_nand2b_1 _2340_ (.Y(_0884_),
    .B(\input_halfprob1_sng_comparator.bits_b[1] ),
    .A_N(\system_integrator_a_counter.value_output[3] ));
 sg13g2_nand2b_1 _2341_ (.Y(_0885_),
    .B(\input_halfprob1_sng_comparator.bits_b[0] ),
    .A_N(net588));
 sg13g2_and4_1 _2342_ (.A(_0881_),
    .B(_0882_),
    .C(_0884_),
    .D(_0885_),
    .X(_0886_));
 sg13g2_nand2b_1 _2343_ (.Y(_0887_),
    .B(\system_integrator_a_counter.value_output[1] ),
    .A_N(\integrator_a_sng_comparator.bits_b[1] ));
 sg13g2_nor2b_1 _2344_ (.A(\system_integrator_a_counter.value_output[0] ),
    .B_N(net595),
    .Y(_0888_));
 sg13g2_xor2_1 _2345_ (.B(\integrator_a_sng_comparator.bits_b[1] ),
    .A(\system_integrator_a_counter.value_output[1] ),
    .X(_0889_));
 sg13g2_o21ai_1 _2346_ (.B1(_0887_),
    .Y(_0890_),
    .A1(_0888_),
    .A2(_0889_));
 sg13g2_a22oi_1 _2347_ (.Y(_0891_),
    .B1(_0886_),
    .B2(_0890_),
    .A2(_0884_),
    .A1(_0883_));
 sg13g2_a21oi_1 _2348_ (.A1(_0876_),
    .A2(_0877_),
    .Y(_0892_),
    .B1(_0878_));
 sg13g2_nor2b_1 _2349_ (.A(\input_halfprob2_sng_comparator.bits_b[5] ),
    .B_N(\system_integrator_a_counter.value_output[8] ),
    .Y(_0893_));
 sg13g2_a221oi_1 _2350_ (.B2(_0892_),
    .C1(_0893_),
    .B1(_0875_),
    .A1(_0872_),
    .Y(_0894_),
    .A2(_0873_));
 sg13g2_o21ai_1 _2351_ (.B1(_0894_),
    .Y(_0895_),
    .A1(_0880_),
    .A2(_0891_));
 sg13g2_nand2_1 _2352_ (.Y(_0896_),
    .A(\system_integrator_a_counter.value_output[0] ),
    .B(_0641_));
 sg13g2_nand3b_1 _2353_ (.B(_0896_),
    .C(_0886_),
    .Y(_0897_),
    .A_N(_0893_));
 sg13g2_or4_1 _2354_ (.A(_0880_),
    .B(_0888_),
    .C(_0889_),
    .D(_0897_),
    .X(_0898_));
 sg13g2_nand2b_1 _2355_ (.Y(_0899_),
    .B(\input_halfprob2_sng_comparator.bits_b[5] ),
    .A_N(\system_integrator_a_counter.value_output[8] ));
 sg13g2_nand3_1 _2356_ (.B(_0898_),
    .C(_0899_),
    .A(_0895_),
    .Y(_0900_));
 sg13g2_and4_1 _2357_ (.A(net595),
    .B(_0895_),
    .C(_0898_),
    .D(_0899_),
    .X(_0901_));
 sg13g2_nand4_1 _2358_ (.B(_0895_),
    .C(_0898_),
    .A(net595),
    .Y(_0902_),
    .D(_0899_));
 sg13g2_nand2_1 _2359_ (.Y(_0903_),
    .A(_0641_),
    .B(_0900_));
 sg13g2_nor3_1 _2360_ (.A(\system_integrator_b_counter.value_output[7] ),
    .B(\system_integrator_b_counter.value_output[5] ),
    .C(\system_integrator_b_counter.value_output[4] ),
    .Y(_0904_));
 sg13g2_nor2_1 _2361_ (.A(\system_integrator_b_counter.value_output[8] ),
    .B(\system_integrator_b_counter.value_output[6] ),
    .Y(_0905_));
 sg13g2_nor4_1 _2362_ (.A(\system_integrator_b_counter.value_output[3] ),
    .B(\system_integrator_b_counter.value_output[2] ),
    .C(\system_integrator_b_counter.value_output[1] ),
    .D(net587),
    .Y(_0906_));
 sg13g2_nand4_1 _2363_ (.B(_0904_),
    .C(_0905_),
    .A(net529),
    .Y(_0907_),
    .D(_0906_));
 sg13g2_nand2_1 _2364_ (.Y(_0908_),
    .A(\system_integrator_b_counter.value_output[1] ),
    .B(net587));
 sg13g2_nand4_1 _2365_ (.B(\system_integrator_b_counter.value_output[6] ),
    .C(\system_integrator_b_counter.value_output[5] ),
    .A(\system_integrator_b_counter.value_output[7] ),
    .Y(_0909_),
    .D(\system_integrator_b_counter.value_output[2] ));
 sg13g2_nor4_1 _2366_ (.A(net595),
    .B(_0029_),
    .C(_0908_),
    .D(_0909_),
    .Y(_0910_));
 sg13g2_nand3_1 _2367_ (.B(\system_integrator_b_counter.value_output[3] ),
    .C(_0910_),
    .A(\system_integrator_b_counter.value_output[4] ),
    .Y(_0911_));
 sg13g2_a21oi_1 _2368_ (.A1(_0907_),
    .A2(_0911_),
    .Y(_0912_),
    .B1(net593));
 sg13g2_a21o_1 _2369_ (.A2(_0903_),
    .A1(_0902_),
    .B1(_0912_),
    .X(_0913_));
 sg13g2_xnor2_1 _2370_ (.Y(_0914_),
    .A(_1628_),
    .B(net528));
 sg13g2_inv_1 _2371_ (.Y(_0915_),
    .A(_0914_));
 sg13g2_nor2_1 _2372_ (.A(_0032_),
    .B(_0902_),
    .Y(_0916_));
 sg13g2_xnor2_1 _2373_ (.Y(_0917_),
    .A(_0032_),
    .B(net528));
 sg13g2_a21oi_2 _2374_ (.B1(_0916_),
    .Y(_0918_),
    .A2(_0917_),
    .A1(net587));
 sg13g2_nand2_1 _2375_ (.Y(_0919_),
    .A(\system_integrator_b_counter.value_output[2] ),
    .B(net528));
 sg13g2_xnor2_1 _2376_ (.Y(_0920_),
    .A(\system_integrator_b_counter.value_output[2] ),
    .B(net528));
 sg13g2_nor3_1 _2377_ (.A(_0915_),
    .B(_0918_),
    .C(_0920_),
    .Y(_0921_));
 sg13g2_a21oi_1 _2378_ (.A1(_1628_),
    .A2(_1629_),
    .Y(_0922_),
    .B1(_0902_));
 sg13g2_nor2_1 _2379_ (.A(_0921_),
    .B(_0922_),
    .Y(_0923_));
 sg13g2_xnor2_1 _2380_ (.Y(_0924_),
    .A(\system_integrator_b_counter.value_output[4] ),
    .B(net528));
 sg13g2_xnor2_1 _2381_ (.Y(_0925_),
    .A(\system_integrator_b_counter.value_output[5] ),
    .B(net528));
 sg13g2_nor2_1 _2382_ (.A(_0924_),
    .B(_0925_),
    .Y(_0926_));
 sg13g2_o21ai_1 _2383_ (.B1(_0926_),
    .Y(_0927_),
    .A1(_0921_),
    .A2(_0922_));
 sg13g2_xnor2_1 _2384_ (.Y(_0928_),
    .A(\system_integrator_b_counter.value_output[6] ),
    .B(net529));
 sg13g2_xnor2_1 _2385_ (.Y(_0929_),
    .A(\system_integrator_b_counter.value_output[7] ),
    .B(net529));
 sg13g2_or2_1 _2386_ (.X(_0930_),
    .B(_0929_),
    .A(_0928_));
 sg13g2_a21o_1 _2387_ (.A2(_0904_),
    .A1(_1625_),
    .B1(_0902_),
    .X(_0931_));
 sg13g2_o21ai_1 _2388_ (.B1(_0931_),
    .Y(_0932_),
    .A1(_0927_),
    .A2(_0930_));
 sg13g2_o21ai_1 _2389_ (.B1(net581),
    .Y(_0933_),
    .A1(net445),
    .A2(_0932_));
 sg13g2_a21oi_1 _2390_ (.A1(net445),
    .A2(_0932_),
    .Y(_0934_),
    .B1(_0933_));
 sg13g2_xnor2_1 _2391_ (.Y(_0935_),
    .A(_0902_),
    .B(_0934_));
 sg13g2_nand2_1 _2392_ (.Y(_0936_),
    .A(net292),
    .B(net514));
 sg13g2_o21ai_1 _2393_ (.B1(_0936_),
    .Y(_0535_),
    .A1(net514),
    .A2(_0935_));
 sg13g2_a21oi_2 _2394_ (.B1(net513),
    .Y(_0937_),
    .A2(net528),
    .A1(net593));
 sg13g2_o21ai_1 _2395_ (.B1(net529),
    .Y(_0938_),
    .A1(\system_integrator_b_counter.value_output[5] ),
    .A2(\system_integrator_b_counter.value_output[4] ));
 sg13g2_a21oi_1 _2396_ (.A1(_0927_),
    .A2(_0938_),
    .Y(_0939_),
    .B1(_0928_));
 sg13g2_a21oi_1 _2397_ (.A1(\system_integrator_b_counter.value_output[6] ),
    .A2(net529),
    .Y(_0940_),
    .B1(_0939_));
 sg13g2_o21ai_1 _2398_ (.B1(net581),
    .Y(_0941_),
    .A1(_0929_),
    .A2(_0940_));
 sg13g2_a21o_1 _2399_ (.A2(_0940_),
    .A1(_0929_),
    .B1(_0941_),
    .X(_0942_));
 sg13g2_a22oi_1 _2400_ (.Y(_0534_),
    .B1(_0937_),
    .B2(_0942_),
    .A2(net513),
    .A1(_1624_));
 sg13g2_nand3_1 _2401_ (.B(_0928_),
    .C(_0938_),
    .A(_0927_),
    .Y(_0943_));
 sg13g2_nor2_1 _2402_ (.A(net593),
    .B(_0939_),
    .Y(_0944_));
 sg13g2_nand2_1 _2403_ (.Y(_0945_),
    .A(_0943_),
    .B(_0944_));
 sg13g2_a22oi_1 _2404_ (.Y(_0533_),
    .B1(_0937_),
    .B2(_0945_),
    .A2(net513),
    .A1(_1625_));
 sg13g2_nor2_1 _2405_ (.A(_0923_),
    .B(_0924_),
    .Y(_0946_));
 sg13g2_a21oi_1 _2406_ (.A1(\system_integrator_b_counter.value_output[4] ),
    .A2(net528),
    .Y(_0947_),
    .B1(_0946_));
 sg13g2_xor2_1 _2407_ (.B(_0947_),
    .A(_0925_),
    .X(_0948_));
 sg13g2_nand2_1 _2408_ (.Y(_0949_),
    .A(net581),
    .B(_0948_));
 sg13g2_a22oi_1 _2409_ (.Y(_0532_),
    .B1(_0937_),
    .B2(_0949_),
    .A2(net513),
    .A1(_1626_));
 sg13g2_and2_1 _2410_ (.A(_0923_),
    .B(_0924_),
    .X(_0950_));
 sg13g2_or3_1 _2411_ (.A(net593),
    .B(_0946_),
    .C(_0950_),
    .X(_0951_));
 sg13g2_a22oi_1 _2412_ (.Y(_0531_),
    .B1(_0937_),
    .B2(_0951_),
    .A2(net513),
    .A1(_1627_));
 sg13g2_o21ai_1 _2413_ (.B1(_0919_),
    .Y(_0952_),
    .A1(_0918_),
    .A2(_0920_));
 sg13g2_xnor2_1 _2414_ (.Y(_0953_),
    .A(_0915_),
    .B(_0952_));
 sg13g2_nand2_1 _2415_ (.Y(_0954_),
    .A(net581),
    .B(_0953_));
 sg13g2_a22oi_1 _2416_ (.Y(_0530_),
    .B1(_0937_),
    .B2(_0954_),
    .A2(net513),
    .A1(_1628_));
 sg13g2_o21ai_1 _2417_ (.B1(net581),
    .Y(_0955_),
    .A1(_0918_),
    .A2(_0920_));
 sg13g2_a21o_1 _2418_ (.A2(_0920_),
    .A1(_0918_),
    .B1(_0955_),
    .X(_0956_));
 sg13g2_a22oi_1 _2419_ (.Y(_0529_),
    .B1(_0937_),
    .B2(_0956_),
    .A2(net513),
    .A1(_1629_));
 sg13g2_a21oi_1 _2420_ (.A1(net587),
    .A2(_0917_),
    .Y(_0957_),
    .B1(net593));
 sg13g2_o21ai_1 _2421_ (.B1(_0957_),
    .Y(_0958_),
    .A1(net587),
    .A2(_0917_));
 sg13g2_a22oi_1 _2422_ (.Y(_0528_),
    .B1(_0937_),
    .B2(_0958_),
    .A2(net513),
    .A1(_1630_));
 sg13g2_a21oi_1 _2423_ (.A1(net587),
    .A2(net581),
    .Y(_0959_),
    .B1(net514));
 sg13g2_a21o_1 _2424_ (.A2(net514),
    .A1(net587),
    .B1(_0959_),
    .X(_0527_));
 sg13g2_nand2b_1 _2425_ (.Y(_0960_),
    .B(\system_integrator_b_counter.value_output[6] ),
    .A_N(\integrator_b_sng_comparator.bits_b[6] ));
 sg13g2_o21ai_1 _2426_ (.B1(_0960_),
    .Y(_0961_),
    .A1(_1624_),
    .A2(net596));
 sg13g2_nand2b_1 _2427_ (.Y(_0962_),
    .B(\integrator_b_sng_comparator.bits_b[6] ),
    .A_N(\system_integrator_b_counter.value_output[6] ));
 sg13g2_nand2b_1 _2428_ (.Y(_0963_),
    .B(net596),
    .A_N(\system_integrator_b_counter.value_output[7] ));
 sg13g2_nand2b_1 _2429_ (.Y(_0964_),
    .B(net597),
    .A_N(\system_integrator_b_counter.value_output[5] ));
 sg13g2_nand3_1 _2430_ (.B(_0963_),
    .C(_0964_),
    .A(_0962_),
    .Y(_0965_));
 sg13g2_nor2_1 _2431_ (.A(_0961_),
    .B(_0965_),
    .Y(_0966_));
 sg13g2_nand2b_1 _2432_ (.Y(_0967_),
    .B(\system_integrator_b_counter.value_output[4] ),
    .A_N(net598));
 sg13g2_o21ai_1 _2433_ (.B1(_0967_),
    .Y(_0968_),
    .A1(_1626_),
    .A2(net597));
 sg13g2_nor2b_1 _2434_ (.A(\system_integrator_b_counter.value_output[4] ),
    .B_N(net598),
    .Y(_0969_));
 sg13g2_nor4_1 _2435_ (.A(_0961_),
    .B(_0965_),
    .C(_0968_),
    .D(_0969_),
    .Y(_0970_));
 sg13g2_nor2b_1 _2436_ (.A(net601),
    .B_N(\system_integrator_b_counter.value_output[2] ),
    .Y(_0971_));
 sg13g2_nor2b_1 _2437_ (.A(net599),
    .B_N(\system_integrator_b_counter.value_output[3] ),
    .Y(_0972_));
 sg13g2_nor2b_1 _2438_ (.A(\system_integrator_b_counter.value_output[3] ),
    .B_N(net599),
    .Y(_0973_));
 sg13g2_nand2b_1 _2439_ (.Y(_0974_),
    .B(net599),
    .A_N(\system_integrator_b_counter.value_output[3] ));
 sg13g2_nor2b_1 _2440_ (.A(\system_integrator_b_counter.value_output[2] ),
    .B_N(net601),
    .Y(_0975_));
 sg13g2_or4_1 _2441_ (.A(_0971_),
    .B(_0972_),
    .C(_0973_),
    .D(_0975_),
    .X(_0976_));
 sg13g2_nor2b_1 _2442_ (.A(net602),
    .B_N(\system_integrator_b_counter.value_output[1] ),
    .Y(_0977_));
 sg13g2_nand2b_1 _2443_ (.Y(_0978_),
    .B(net603),
    .A_N(\system_integrator_b_counter.value_output[0] ));
 sg13g2_xnor2_1 _2444_ (.Y(_0979_),
    .A(\system_integrator_b_counter.value_output[1] ),
    .B(net602));
 sg13g2_nand2_1 _2445_ (.Y(_0980_),
    .A(_0978_),
    .B(_0979_));
 sg13g2_a21oi_1 _2446_ (.A1(_0978_),
    .A2(_0979_),
    .Y(_0981_),
    .B1(_0977_));
 sg13g2_o21ai_1 _2447_ (.B1(_0974_),
    .Y(_0982_),
    .A1(_0971_),
    .A2(_0972_));
 sg13g2_o21ai_1 _2448_ (.B1(_0982_),
    .Y(_0983_),
    .A1(_0976_),
    .A2(_0981_));
 sg13g2_nor2b_1 _2449_ (.A(\integrator_b_sng_comparator.bits_b[8] ),
    .B_N(\system_integrator_b_counter.value_output[8] ),
    .Y(_0984_));
 sg13g2_a21o_1 _2450_ (.A2(_0963_),
    .A1(_0961_),
    .B1(_0984_),
    .X(_0985_));
 sg13g2_a221oi_1 _2451_ (.B2(_0983_),
    .C1(_0985_),
    .B1(_0970_),
    .A1(_0966_),
    .Y(_0986_),
    .A2(_0968_));
 sg13g2_nor2b_1 _2452_ (.A(net603),
    .B_N(net587),
    .Y(_0987_));
 sg13g2_nor4_1 _2453_ (.A(_0976_),
    .B(_0980_),
    .C(_0984_),
    .D(_0987_),
    .Y(_0988_));
 sg13g2_nor2b_1 _2454_ (.A(\system_integrator_b_counter.value_output[8] ),
    .B_N(\integrator_b_sng_comparator.bits_b[8] ),
    .Y(_0989_));
 sg13g2_a21o_1 _2455_ (.A2(_0988_),
    .A1(_0970_),
    .B1(_0989_),
    .X(_0990_));
 sg13g2_or2_1 _2456_ (.X(_0991_),
    .B(_0990_),
    .A(_0986_));
 sg13g2_and2_2 _2457_ (.A(_0653_),
    .B(_0991_),
    .X(_0992_));
 sg13g2_o21ai_1 _2458_ (.B1(_0653_),
    .Y(_0993_),
    .A1(_0986_),
    .A2(_0990_));
 sg13g2_nor2_1 _2459_ (.A(\system_integrator_a_counter.value_output[8] ),
    .B(\system_integrator_a_counter.value_output[3] ),
    .Y(_0994_));
 sg13g2_nor4_1 _2460_ (.A(net588),
    .B(\system_integrator_a_counter.value_output[1] ),
    .C(\system_integrator_a_counter.value_output[0] ),
    .D(net594),
    .Y(_0995_));
 sg13g2_nand3_1 _2461_ (.B(\system_integrator_a_counter.value_output[1] ),
    .C(\system_integrator_a_counter.value_output[0] ),
    .A(net588),
    .Y(_0996_));
 sg13g2_nand4_1 _2462_ (.B(\system_integrator_a_counter.value_output[7] ),
    .C(\system_integrator_a_counter.value_output[6] ),
    .A(\system_integrator_a_counter.value_output[8] ),
    .Y(_0997_),
    .D(\system_integrator_a_counter.value_output[3] ));
 sg13g2_nand2_1 _2463_ (.Y(_0998_),
    .A(\system_integrator_a_counter.value_output[5] ),
    .B(\system_integrator_a_counter.value_output[4] ));
 sg13g2_nor4_1 _2464_ (.A(net594),
    .B(_0996_),
    .C(_0997_),
    .D(_0998_),
    .Y(_0999_));
 sg13g2_nor2_1 _2465_ (.A(_0991_),
    .B(_0999_),
    .Y(_1000_));
 sg13g2_nor4_1 _2466_ (.A(\system_integrator_a_counter.value_output[7] ),
    .B(\system_integrator_a_counter.value_output[6] ),
    .C(\system_integrator_a_counter.value_output[5] ),
    .D(\system_integrator_a_counter.value_output[4] ),
    .Y(_1001_));
 sg13g2_nor2_1 _2467_ (.A(net527),
    .B(_1001_),
    .Y(_1002_));
 sg13g2_nand3_1 _2468_ (.B(_0995_),
    .C(_1001_),
    .A(_0994_),
    .Y(_1003_));
 sg13g2_a22oi_1 _2469_ (.Y(_1004_),
    .B1(_1003_),
    .B2(_0992_),
    .A2(_1000_),
    .A1(net31));
 sg13g2_nand2_1 _2470_ (.Y(_1005_),
    .A(net257),
    .B(net518));
 sg13g2_xnor2_1 _2471_ (.Y(_1006_),
    .A(\system_integrator_a_counter.value_output[4] ),
    .B(net527));
 sg13g2_and2_1 _2472_ (.A(\system_integrator_a_counter.value_output[3] ),
    .B(_0992_),
    .X(_1007_));
 sg13g2_nand2b_1 _2473_ (.Y(_1008_),
    .B(_0993_),
    .A_N(\system_integrator_a_counter.value_output[3] ));
 sg13g2_nand2_1 _2474_ (.Y(_1009_),
    .A(net588),
    .B(_0992_));
 sg13g2_nor2_1 _2475_ (.A(_0031_),
    .B(net527),
    .Y(_1010_));
 sg13g2_xor2_1 _2476_ (.B(net527),
    .A(_0031_),
    .X(_1011_));
 sg13g2_a21oi_2 _2477_ (.B1(_1010_),
    .Y(_1012_),
    .A2(_1011_),
    .A1(\system_integrator_a_counter.value_output[0] ));
 sg13g2_nor2_1 _2478_ (.A(net588),
    .B(_0992_),
    .Y(_1013_));
 sg13g2_xnor2_1 _2479_ (.Y(_1014_),
    .A(net588),
    .B(_0993_));
 sg13g2_nor2b_1 _2480_ (.A(_1012_),
    .B_N(_1014_),
    .Y(_1015_));
 sg13g2_o21ai_1 _2481_ (.B1(_1009_),
    .Y(_1016_),
    .A1(_1012_),
    .A2(_1013_));
 sg13g2_a21o_1 _2482_ (.A2(_1016_),
    .A1(_1008_),
    .B1(_1007_),
    .X(_1017_));
 sg13g2_and2_1 _2483_ (.A(_1006_),
    .B(_1017_),
    .X(_1018_));
 sg13g2_xnor2_1 _2484_ (.Y(_1019_),
    .A(\system_integrator_a_counter.value_output[5] ),
    .B(net527));
 sg13g2_nand3_1 _2485_ (.B(_1017_),
    .C(_1019_),
    .A(_1006_),
    .Y(_1020_));
 sg13g2_xnor2_1 _2486_ (.Y(_1021_),
    .A(\system_integrator_a_counter.value_output[7] ),
    .B(net527));
 sg13g2_xnor2_1 _2487_ (.Y(_1022_),
    .A(\system_integrator_a_counter.value_output[6] ),
    .B(net527));
 sg13g2_inv_1 _2488_ (.Y(_1023_),
    .A(_1022_));
 sg13g2_nor2_1 _2489_ (.A(_1020_),
    .B(_1023_),
    .Y(_1024_));
 sg13g2_a21oi_1 _2490_ (.A1(_1021_),
    .A2(_1024_),
    .Y(_1025_),
    .B1(_1002_));
 sg13g2_xor2_1 _2491_ (.B(net527),
    .A(\system_integrator_a_counter.value_output[8] ),
    .X(_1026_));
 sg13g2_or2_2 _2492_ (.X(_1027_),
    .B(net518),
    .A(net594));
 sg13g2_xnor2_1 _2493_ (.Y(_1028_),
    .A(_1025_),
    .B(_1026_));
 sg13g2_o21ai_1 _2494_ (.B1(_1005_),
    .Y(_0526_),
    .A1(_1027_),
    .A2(_1028_));
 sg13g2_nand2_1 _2495_ (.Y(_1029_),
    .A(net453),
    .B(net518));
 sg13g2_o21ai_1 _2496_ (.B1(_0992_),
    .Y(_1030_),
    .A1(\system_integrator_a_counter.value_output[5] ),
    .A2(\system_integrator_a_counter.value_output[4] ));
 sg13g2_a21oi_1 _2497_ (.A1(_1020_),
    .A2(_1030_),
    .Y(_1031_),
    .B1(_1023_));
 sg13g2_a21o_1 _2498_ (.A2(_0992_),
    .A1(\system_integrator_a_counter.value_output[6] ),
    .B1(_1031_),
    .X(_1032_));
 sg13g2_nor2_1 _2499_ (.A(_1021_),
    .B(_1032_),
    .Y(_1033_));
 sg13g2_a21o_1 _2500_ (.A2(_1032_),
    .A1(_1021_),
    .B1(_1027_),
    .X(_1034_));
 sg13g2_o21ai_1 _2501_ (.B1(_1029_),
    .Y(_0525_),
    .A1(_1033_),
    .A2(_1034_));
 sg13g2_nand2_1 _2502_ (.Y(_1035_),
    .A(net459),
    .B(net518));
 sg13g2_nand3_1 _2503_ (.B(_1023_),
    .C(_1030_),
    .A(_1020_),
    .Y(_1036_));
 sg13g2_nand2b_1 _2504_ (.Y(_1037_),
    .B(_1036_),
    .A_N(_1031_));
 sg13g2_o21ai_1 _2505_ (.B1(_1035_),
    .Y(_0524_),
    .A1(_1027_),
    .A2(_1037_));
 sg13g2_nand2_1 _2506_ (.Y(_1038_),
    .A(net460),
    .B(net518));
 sg13g2_a21oi_1 _2507_ (.A1(\system_integrator_a_counter.value_output[4] ),
    .A2(_0992_),
    .Y(_1039_),
    .B1(_1018_));
 sg13g2_xor2_1 _2508_ (.B(_1039_),
    .A(_1019_),
    .X(_1040_));
 sg13g2_o21ai_1 _2509_ (.B1(_1038_),
    .Y(_0523_),
    .A1(_1027_),
    .A2(_1040_));
 sg13g2_nor2_1 _2510_ (.A(_1006_),
    .B(_1017_),
    .Y(_1041_));
 sg13g2_nor3_1 _2511_ (.A(_1018_),
    .B(_1027_),
    .C(_1041_),
    .Y(_1042_));
 sg13g2_a21o_1 _2512_ (.A2(net518),
    .A1(net471),
    .B1(_1042_),
    .X(_0522_));
 sg13g2_nand2_1 _2513_ (.Y(_1043_),
    .A(net463),
    .B(_1004_));
 sg13g2_nor2b_1 _2514_ (.A(_1007_),
    .B_N(_1008_),
    .Y(_1044_));
 sg13g2_nor2_1 _2515_ (.A(_1016_),
    .B(_1044_),
    .Y(_1045_));
 sg13g2_a21o_1 _2516_ (.A2(_1044_),
    .A1(_1016_),
    .B1(_1027_),
    .X(_1046_));
 sg13g2_o21ai_1 _2517_ (.B1(_1043_),
    .Y(_0521_),
    .A1(_1045_),
    .A2(_1046_));
 sg13g2_nand2b_1 _2518_ (.Y(_1047_),
    .B(_1012_),
    .A_N(_1014_));
 sg13g2_nor2_1 _2519_ (.A(_1015_),
    .B(_1027_),
    .Y(_1048_));
 sg13g2_a22oi_1 _2520_ (.Y(_1049_),
    .B1(_1047_),
    .B2(_1048_),
    .A2(_1004_),
    .A1(net588));
 sg13g2_inv_1 _2521_ (.Y(_0520_),
    .A(net490));
 sg13g2_nand2_1 _2522_ (.Y(_1050_),
    .A(net461),
    .B(_1004_));
 sg13g2_xnor2_1 _2523_ (.Y(_1051_),
    .A(net252),
    .B(_1011_));
 sg13g2_o21ai_1 _2524_ (.B1(_1050_),
    .Y(_0519_),
    .A1(_1027_),
    .A2(_1051_));
 sg13g2_nor2_1 _2525_ (.A(net582),
    .B(_0992_),
    .Y(_1052_));
 sg13g2_a21oi_1 _2526_ (.A1(net582),
    .A2(net102),
    .Y(_1053_),
    .B1(_1052_));
 sg13g2_nand2_1 _2527_ (.Y(_1054_),
    .A(\system_integrator_a_counter.value_output[0] ),
    .B(net518));
 sg13g2_o21ai_1 _2528_ (.B1(_1054_),
    .Y(_0518_),
    .A1(net518),
    .A2(_1053_));
 sg13g2_nand2b_1 _2529_ (.Y(_1055_),
    .B(\input_b_sng_comparator.bits_a[6] ),
    .A_N(net601));
 sg13g2_nand2b_1 _2530_ (.Y(_1056_),
    .B(\input_b_sng_comparator.bits_a[7] ),
    .A_N(net600));
 sg13g2_nand2_1 _2531_ (.Y(_1057_),
    .A(_1055_),
    .B(_1056_));
 sg13g2_nand2b_1 _2532_ (.Y(_1058_),
    .B(net600),
    .A_N(\input_b_sng_comparator.bits_a[7] ));
 sg13g2_nand2b_1 _2533_ (.Y(_1059_),
    .B(\input_a_sng_comparator.bits_b[3] ),
    .A_N(\input_b_sng_comparator.bits_a[6] ));
 sg13g2_nand4_1 _2534_ (.B(_1056_),
    .C(_1058_),
    .A(_1055_),
    .Y(_1060_),
    .D(_1059_));
 sg13g2_nor2b_1 _2535_ (.A(net603),
    .B_N(\input_b_sng_comparator.bits_a[4] ),
    .Y(_1061_));
 sg13g2_nor2b_1 _2536_ (.A(\input_a_sng_comparator.bits_b[2] ),
    .B_N(\input_b_sng_comparator.bits_a[5] ),
    .Y(_1062_));
 sg13g2_nand2b_1 _2537_ (.Y(_1063_),
    .B(\input_a_sng_comparator.bits_b[2] ),
    .A_N(\input_b_sng_comparator.bits_a[5] ));
 sg13g2_o21ai_1 _2538_ (.B1(_1063_),
    .Y(_1064_),
    .A1(\input_b_sng_comparator.bits_a[4] ),
    .A2(_0633_));
 sg13g2_nor4_1 _2539_ (.A(_1060_),
    .B(_1061_),
    .C(_1062_),
    .D(_1064_),
    .Y(_1065_));
 sg13g2_nor2b_1 _2540_ (.A(\input_b_sng_comparator.bits_b[2] ),
    .B_N(\input_b_sng_comparator.bits_a[2] ),
    .Y(_1066_));
 sg13g2_nor2b_1 _2541_ (.A(\input_a_sng_comparator.bits_b[0] ),
    .B_N(\input_b_sng_comparator.bits_a[3] ),
    .Y(_1067_));
 sg13g2_nor2b_1 _2542_ (.A(\input_b_sng_comparator.bits_a[3] ),
    .B_N(\input_a_sng_comparator.bits_b[0] ),
    .Y(_1068_));
 sg13g2_nand2b_1 _2543_ (.Y(_1069_),
    .B(\input_a_sng_comparator.bits_b[0] ),
    .A_N(\input_b_sng_comparator.bits_a[3] ));
 sg13g2_nor2b_1 _2544_ (.A(\input_b_sng_comparator.bits_a[2] ),
    .B_N(\input_b_sng_comparator.bits_b[2] ),
    .Y(_1070_));
 sg13g2_or4_1 _2545_ (.A(_1066_),
    .B(_1067_),
    .C(_1068_),
    .D(_1070_),
    .X(_1071_));
 sg13g2_nor2b_1 _2546_ (.A(\input_b_sng_comparator.bits_b[1] ),
    .B_N(\input_b_sng_comparator.bits_a[1] ),
    .Y(_1072_));
 sg13g2_nand2b_1 _2547_ (.Y(_1073_),
    .B(\input_b_sng_comparator.bits_b[0] ),
    .A_N(\input_b_sng_comparator.bits_a[0] ));
 sg13g2_nand2b_1 _2548_ (.Y(_1074_),
    .B(\input_b_sng_comparator.bits_b[1] ),
    .A_N(\input_b_sng_comparator.bits_a[1] ));
 sg13g2_nand2_1 _2549_ (.Y(_1075_),
    .A(_1073_),
    .B(_1074_));
 sg13g2_a21oi_1 _2550_ (.A1(_1073_),
    .A2(_1074_),
    .Y(_1076_),
    .B1(_1072_));
 sg13g2_o21ai_1 _2551_ (.B1(_1069_),
    .Y(_1077_),
    .A1(_1066_),
    .A2(_1067_));
 sg13g2_o21ai_1 _2552_ (.B1(_1077_),
    .Y(_1078_),
    .A1(_1071_),
    .A2(_1076_));
 sg13g2_a21oi_1 _2553_ (.A1(_1061_),
    .A2(_1063_),
    .Y(_1079_),
    .B1(_1062_));
 sg13g2_nand2b_1 _2554_ (.Y(_1080_),
    .B(\input_b_sng_comparator.bits_a[8] ),
    .A_N(\input_a_sng_comparator.bits_b[5] ));
 sg13g2_o21ai_1 _2555_ (.B1(_1080_),
    .Y(_1081_),
    .A1(_1060_),
    .A2(_1079_));
 sg13g2_a221oi_1 _2556_ (.B2(_1078_),
    .C1(_1081_),
    .B1(_1065_),
    .A1(_1057_),
    .Y(_1082_),
    .A2(_1058_));
 sg13g2_o21ai_1 _2557_ (.B1(_1080_),
    .Y(_1083_),
    .A1(_1614_),
    .A2(\input_b_sng_comparator.bits_b[0] ));
 sg13g2_nor4_1 _2558_ (.A(_1071_),
    .B(_1072_),
    .C(_1075_),
    .D(_1083_),
    .Y(_1084_));
 sg13g2_a221oi_1 _2559_ (.B2(_1084_),
    .C1(_1082_),
    .B1(_1065_),
    .A1(_1613_),
    .Y(_1085_),
    .A2(\input_a_sng_comparator.bits_b[5] ));
 sg13g2_nand2b_1 _2560_ (.Y(_1086_),
    .B(net589),
    .A_N(\integrator_b_sng_comparator.bits_b[6] ));
 sg13g2_o21ai_1 _2561_ (.B1(_1086_),
    .Y(_1087_),
    .A1(_1641_),
    .A2(net596));
 sg13g2_nor2_1 _2562_ (.A(net589),
    .B(_0634_),
    .Y(_1088_));
 sg13g2_nand2b_1 _2563_ (.Y(_1089_),
    .B(net596),
    .A_N(\integrator_b_counter.value_output[7] ));
 sg13g2_o21ai_1 _2564_ (.B1(_1089_),
    .Y(_1090_),
    .A1(\integrator_b_counter.value_output[5] ),
    .A2(_1655_));
 sg13g2_nor3_1 _2565_ (.A(_1087_),
    .B(_1088_),
    .C(_1090_),
    .Y(_1091_));
 sg13g2_nand2b_1 _2566_ (.Y(_1092_),
    .B(\integrator_b_counter.value_output[5] ),
    .A_N(net597));
 sg13g2_nand2b_1 _2567_ (.Y(_1093_),
    .B(\integrator_b_counter.value_output[4] ),
    .A_N(net598));
 sg13g2_nand2_1 _2568_ (.Y(_1094_),
    .A(_1092_),
    .B(_1093_));
 sg13g2_nand2b_1 _2569_ (.Y(_1095_),
    .B(net598),
    .A_N(\integrator_b_counter.value_output[4] ));
 sg13g2_nand3_1 _2570_ (.B(_1093_),
    .C(_1095_),
    .A(_1092_),
    .Y(_1096_));
 sg13g2_nor4_1 _2571_ (.A(_1087_),
    .B(_1088_),
    .C(_1090_),
    .D(_1096_),
    .Y(_1097_));
 sg13g2_nor2b_1 _2572_ (.A(net601),
    .B_N(\integrator_b_counter.value_output[2] ),
    .Y(_1098_));
 sg13g2_nor2b_1 _2573_ (.A(net599),
    .B_N(\integrator_b_counter.value_output[3] ),
    .Y(_1099_));
 sg13g2_nor2b_1 _2574_ (.A(\integrator_b_counter.value_output[3] ),
    .B_N(net599),
    .Y(_1100_));
 sg13g2_nand2b_1 _2575_ (.Y(_1101_),
    .B(net599),
    .A_N(\integrator_b_counter.value_output[3] ));
 sg13g2_nor2b_1 _2576_ (.A(\integrator_b_counter.value_output[2] ),
    .B_N(net601),
    .Y(_1102_));
 sg13g2_or4_1 _2577_ (.A(_1098_),
    .B(_1099_),
    .C(_1100_),
    .D(_1102_),
    .X(_1103_));
 sg13g2_nor2b_1 _2578_ (.A(net602),
    .B_N(\integrator_b_counter.value_output[1] ),
    .Y(_1104_));
 sg13g2_nand2b_1 _2579_ (.Y(_1105_),
    .B(net603),
    .A_N(\integrator_b_counter.value_output[0] ));
 sg13g2_xnor2_1 _2580_ (.Y(_1106_),
    .A(\integrator_b_counter.value_output[1] ),
    .B(net602));
 sg13g2_a21oi_1 _2581_ (.A1(_1105_),
    .A2(_1106_),
    .Y(_1107_),
    .B1(_1104_));
 sg13g2_o21ai_1 _2582_ (.B1(_1101_),
    .Y(_1108_),
    .A1(_1098_),
    .A2(_1099_));
 sg13g2_o21ai_1 _2583_ (.B1(_1108_),
    .Y(_1109_),
    .A1(_1103_),
    .A2(_1107_));
 sg13g2_nor2b_1 _2584_ (.A(\integrator_b_sng_comparator.bits_b[8] ),
    .B_N(\integrator_b_counter.value_output[8] ),
    .Y(_1110_));
 sg13g2_a21o_1 _2585_ (.A2(_1089_),
    .A1(_1087_),
    .B1(_1110_),
    .X(_1111_));
 sg13g2_a221oi_1 _2586_ (.B2(_1109_),
    .C1(_1111_),
    .B1(_1097_),
    .A1(_1091_),
    .Y(_1112_),
    .A2(_1094_));
 sg13g2_nor2_1 _2587_ (.A(_1643_),
    .B(net603),
    .Y(_1113_));
 sg13g2_nor3_1 _2588_ (.A(_1103_),
    .B(_1110_),
    .C(_1113_),
    .Y(_1114_));
 sg13g2_nand4_1 _2589_ (.B(_1105_),
    .C(_1106_),
    .A(_1097_),
    .Y(_1115_),
    .D(_1114_));
 sg13g2_nand2b_1 _2590_ (.Y(_1116_),
    .B(\integrator_b_sng_comparator.bits_b[8] ),
    .A_N(\integrator_b_counter.value_output[8] ));
 sg13g2_nand3b_1 _2591_ (.B(_1115_),
    .C(_1116_),
    .Y(_1117_),
    .A_N(_1112_));
 sg13g2_and2_1 _2592_ (.A(net526),
    .B(_1117_),
    .X(_1118_));
 sg13g2_nand2_1 _2593_ (.Y(_1119_),
    .A(net526),
    .B(_1117_));
 sg13g2_nor3_1 _2594_ (.A(\integrator_c_counter.value_output[2] ),
    .B(\integrator_c_counter.value_output[1] ),
    .C(\integrator_c_counter.value_output[0] ),
    .Y(_1120_));
 sg13g2_nor4_1 _2595_ (.A(\integrator_c_counter.value_output[6] ),
    .B(\integrator_c_counter.value_output[5] ),
    .C(\integrator_c_counter.value_output[4] ),
    .D(\integrator_c_counter.value_output[3] ),
    .Y(_1121_));
 sg13g2_nand4_1 _2596_ (.B(_1633_),
    .C(_1120_),
    .A(_1632_),
    .Y(_1122_),
    .D(_1121_));
 sg13g2_nand3b_1 _2597_ (.B(\integrator_c_counter.value_output[0] ),
    .C(\integrator_c_counter.value_output[1] ),
    .Y(_1123_),
    .A_N(_0053_));
 sg13g2_nand4_1 _2598_ (.B(\integrator_c_counter.value_output[4] ),
    .C(\integrator_c_counter.value_output[3] ),
    .A(\integrator_c_counter.value_output[5] ),
    .Y(_1124_),
    .D(\integrator_c_counter.value_output[2] ));
 sg13g2_nor4_1 _2599_ (.A(_1633_),
    .B(_1634_),
    .C(_1123_),
    .D(_1124_),
    .Y(_1125_));
 sg13g2_nor3_1 _2600_ (.A(net526),
    .B(_1117_),
    .C(_1125_),
    .Y(_1126_));
 sg13g2_a21o_1 _2601_ (.A2(_1122_),
    .A1(net524),
    .B1(_1126_),
    .X(_1127_));
 sg13g2_nor2_1 _2602_ (.A(net312),
    .B(net517),
    .Y(_1128_));
 sg13g2_a21o_1 _2603_ (.A2(_0049_),
    .A1(_1636_),
    .B1(_1119_),
    .X(_1129_));
 sg13g2_o21ai_1 _2604_ (.B1(net524),
    .Y(_1130_),
    .A1(\integrator_c_counter.value_output[7] ),
    .A2(\integrator_c_counter.value_output[6] ));
 sg13g2_xnor2_1 _2605_ (.Y(_1131_),
    .A(\integrator_c_counter.value_output[4] ),
    .B(net525));
 sg13g2_nor2_1 _2606_ (.A(_0660_),
    .B(net525),
    .Y(_1132_));
 sg13g2_nor2_1 _2607_ (.A(_1638_),
    .B(_1119_),
    .Y(_1133_));
 sg13g2_xnor2_1 _2608_ (.Y(_1134_),
    .A(_1638_),
    .B(net525));
 sg13g2_nand3_1 _2609_ (.B(net526),
    .C(_1117_),
    .A(_0659_),
    .Y(_1135_));
 sg13g2_a21oi_1 _2610_ (.A1(net526),
    .A2(_1117_),
    .Y(_1136_),
    .B1(_0659_));
 sg13g2_a21oi_2 _2611_ (.B1(_1136_),
    .Y(_1137_),
    .A2(_1135_),
    .A1(_1640_));
 sg13g2_nand2_1 _2612_ (.Y(_1138_),
    .A(_1134_),
    .B(_1137_));
 sg13g2_nand2b_1 _2613_ (.Y(_1139_),
    .B(_1138_),
    .A_N(_1133_));
 sg13g2_a221oi_1 _2614_ (.B2(_1137_),
    .C1(_1133_),
    .B1(_1134_),
    .A1(_0660_),
    .Y(_1140_),
    .A2(net525));
 sg13g2_nor3_1 _2615_ (.A(_1131_),
    .B(_1132_),
    .C(_1140_),
    .Y(_1141_));
 sg13g2_xnor2_1 _2616_ (.Y(_1142_),
    .A(_0049_),
    .B(net524));
 sg13g2_nand2_1 _2617_ (.Y(_1143_),
    .A(_1141_),
    .B(_1142_));
 sg13g2_xnor2_1 _2618_ (.Y(_1144_),
    .A(\integrator_c_counter.value_output[7] ),
    .B(net524));
 sg13g2_xnor2_1 _2619_ (.Y(_1145_),
    .A(\integrator_c_counter.value_output[6] ),
    .B(net524));
 sg13g2_or3_1 _2620_ (.A(_1143_),
    .B(_1144_),
    .C(_1145_),
    .X(_1146_));
 sg13g2_nand3_1 _2621_ (.B(_1130_),
    .C(_1146_),
    .A(_1129_),
    .Y(_1147_));
 sg13g2_xnor2_1 _2622_ (.Y(_1148_),
    .A(net402),
    .B(net524));
 sg13g2_xnor2_1 _2623_ (.Y(_1149_),
    .A(_1147_),
    .B(_1148_));
 sg13g2_a21oi_1 _2624_ (.A1(net517),
    .A2(_1149_),
    .Y(_0517_),
    .B1(_1128_));
 sg13g2_a21oi_1 _2625_ (.A1(_1129_),
    .A2(_1143_),
    .Y(_1150_),
    .B1(_1145_));
 sg13g2_inv_1 _2626_ (.Y(_1151_),
    .A(_1150_));
 sg13g2_a21oi_1 _2627_ (.A1(net506),
    .A2(net524),
    .Y(_1152_),
    .B1(_1150_));
 sg13g2_xnor2_1 _2628_ (.Y(_1153_),
    .A(_1144_),
    .B(_1152_));
 sg13g2_nor2_1 _2629_ (.A(net433),
    .B(net515),
    .Y(_1154_));
 sg13g2_a21oi_1 _2630_ (.A1(net515),
    .A2(_1153_),
    .Y(_0516_),
    .B1(_1154_));
 sg13g2_nand3_1 _2631_ (.B(_1143_),
    .C(_1145_),
    .A(_1129_),
    .Y(_1155_));
 sg13g2_nand3_1 _2632_ (.B(_1151_),
    .C(_1155_),
    .A(net515),
    .Y(_1156_));
 sg13g2_o21ai_1 _2633_ (.B1(_1156_),
    .Y(_0515_),
    .A1(_1634_),
    .A2(net515));
 sg13g2_nor2_1 _2634_ (.A(net410),
    .B(net516),
    .Y(_1157_));
 sg13g2_a21oi_1 _2635_ (.A1(\integrator_c_counter.value_output[4] ),
    .A2(net525),
    .Y(_1158_),
    .B1(_1141_));
 sg13g2_xor2_1 _2636_ (.B(_1158_),
    .A(_1142_),
    .X(_1159_));
 sg13g2_a21oi_1 _2637_ (.A1(net515),
    .A2(_1159_),
    .Y(_0514_),
    .B1(_1157_));
 sg13g2_nor2_1 _2638_ (.A(net442),
    .B(net516),
    .Y(_1160_));
 sg13g2_o21ai_1 _2639_ (.B1(_1131_),
    .Y(_1161_),
    .A1(_1132_),
    .A2(_1140_));
 sg13g2_nand2b_1 _2640_ (.Y(_1162_),
    .B(_1161_),
    .A_N(_1141_));
 sg13g2_a21oi_1 _2641_ (.A1(net515),
    .A2(_1162_),
    .Y(_0513_),
    .B1(_1160_));
 sg13g2_xnor2_1 _2642_ (.Y(_1163_),
    .A(_0048_),
    .B(net524));
 sg13g2_xnor2_1 _2643_ (.Y(_1164_),
    .A(_1139_),
    .B(_1163_));
 sg13g2_nor2_1 _2644_ (.A(net407),
    .B(net515),
    .Y(_1165_));
 sg13g2_a21oi_1 _2645_ (.A1(net515),
    .A2(_1164_),
    .Y(_0512_),
    .B1(_1165_));
 sg13g2_and2_1 _2646_ (.A(net516),
    .B(_1138_),
    .X(_1166_));
 sg13g2_o21ai_1 _2647_ (.B1(_1166_),
    .Y(_1167_),
    .A1(_1134_),
    .A2(_1137_));
 sg13g2_o21ai_1 _2648_ (.B1(_1167_),
    .Y(_0511_),
    .A1(_1638_),
    .A2(net516));
 sg13g2_nor2_1 _2649_ (.A(net415),
    .B(net517),
    .Y(_1168_));
 sg13g2_xnor2_1 _2650_ (.Y(_1169_),
    .A(_0659_),
    .B(net525));
 sg13g2_xnor2_1 _2651_ (.Y(_1170_),
    .A(net47),
    .B(_1169_));
 sg13g2_a21oi_1 _2652_ (.A1(net517),
    .A2(_1170_),
    .Y(_0510_),
    .B1(_1168_));
 sg13g2_nand2_1 _2653_ (.Y(_1171_),
    .A(net47),
    .B(net517));
 sg13g2_o21ai_1 _2654_ (.B1(_1171_),
    .Y(_0509_),
    .A1(_1640_),
    .A2(net517));
 sg13g2_nand2b_1 _2655_ (.Y(_1172_),
    .B(\integrator_a_counter.value_output[6] ),
    .A_N(\input_halfprob2_sng_comparator.bits_b[3] ));
 sg13g2_o21ai_1 _2656_ (.B1(_1172_),
    .Y(_1173_),
    .A1(_1644_),
    .A2(\input_halfprob2_sng_comparator.bits_b[4] ));
 sg13g2_nor2_1 _2657_ (.A(\integrator_a_counter.value_output[5] ),
    .B(_0638_),
    .Y(_1174_));
 sg13g2_nand2b_1 _2658_ (.Y(_1175_),
    .B(\input_halfprob2_sng_comparator.bits_b[4] ),
    .A_N(\integrator_a_counter.value_output[7] ));
 sg13g2_o21ai_1 _2659_ (.B1(_1175_),
    .Y(_1176_),
    .A1(net590),
    .A2(_0637_));
 sg13g2_nor3_1 _2660_ (.A(_1173_),
    .B(_1174_),
    .C(_1176_),
    .Y(_1177_));
 sg13g2_nand2b_1 _2661_ (.Y(_1178_),
    .B(\integrator_a_counter.value_output[5] ),
    .A_N(\input_halfprob2_sng_comparator.bits_b[2] ));
 sg13g2_nand2b_1 _2662_ (.Y(_1179_),
    .B(\integrator_a_counter.value_output[4] ),
    .A_N(\input_halfprob2_sng_comparator.bits_b[1] ));
 sg13g2_nand2_1 _2663_ (.Y(_1180_),
    .A(_1178_),
    .B(_1179_));
 sg13g2_nand2b_1 _2664_ (.Y(_1181_),
    .B(\input_halfprob2_sng_comparator.bits_b[1] ),
    .A_N(\integrator_a_counter.value_output[4] ));
 sg13g2_nand3_1 _2665_ (.B(_1179_),
    .C(_1181_),
    .A(_1178_),
    .Y(_1182_));
 sg13g2_nor4_1 _2666_ (.A(_1173_),
    .B(_1174_),
    .C(_1176_),
    .D(_1182_),
    .Y(_1183_));
 sg13g2_nor2b_1 _2667_ (.A(\input_halfprob1_sng_comparator.bits_b[0] ),
    .B_N(\integrator_a_counter.value_output[2] ),
    .Y(_1184_));
 sg13g2_nor2b_1 _2668_ (.A(\input_halfprob1_sng_comparator.bits_b[1] ),
    .B_N(\integrator_a_counter.value_output[3] ),
    .Y(_1185_));
 sg13g2_nor2b_1 _2669_ (.A(\integrator_a_counter.value_output[3] ),
    .B_N(\input_halfprob1_sng_comparator.bits_b[1] ),
    .Y(_1186_));
 sg13g2_nand2b_1 _2670_ (.Y(_1187_),
    .B(\input_halfprob1_sng_comparator.bits_b[1] ),
    .A_N(\integrator_a_counter.value_output[3] ));
 sg13g2_nor2b_1 _2671_ (.A(\integrator_a_counter.value_output[2] ),
    .B_N(\input_halfprob1_sng_comparator.bits_b[0] ),
    .Y(_1188_));
 sg13g2_or4_1 _2672_ (.A(_1184_),
    .B(_1185_),
    .C(_1186_),
    .D(_1188_),
    .X(_1189_));
 sg13g2_nor2b_1 _2673_ (.A(\integrator_a_sng_comparator.bits_b[1] ),
    .B_N(\integrator_a_counter.value_output[1] ),
    .Y(_1190_));
 sg13g2_nand2b_1 _2674_ (.Y(_1191_),
    .B(net595),
    .A_N(\integrator_a_counter.value_output[0] ));
 sg13g2_xnor2_1 _2675_ (.Y(_1192_),
    .A(\integrator_a_counter.value_output[1] ),
    .B(\integrator_a_sng_comparator.bits_b[1] ));
 sg13g2_a21oi_1 _2676_ (.A1(_1191_),
    .A2(_1192_),
    .Y(_1193_),
    .B1(_1190_));
 sg13g2_o21ai_1 _2677_ (.B1(_1187_),
    .Y(_1194_),
    .A1(_1184_),
    .A2(_1185_));
 sg13g2_o21ai_1 _2678_ (.B1(_1194_),
    .Y(_1195_),
    .A1(_1189_),
    .A2(_1193_));
 sg13g2_nor2b_1 _2679_ (.A(\input_halfprob2_sng_comparator.bits_b[5] ),
    .B_N(\integrator_a_counter.value_output[8] ),
    .Y(_1196_));
 sg13g2_a21o_1 _2680_ (.A2(_1175_),
    .A1(_1173_),
    .B1(_1196_),
    .X(_1197_));
 sg13g2_a221oi_1 _2681_ (.B2(_1195_),
    .C1(_1197_),
    .B1(_1183_),
    .A1(_1177_),
    .Y(_1198_),
    .A2(_1180_));
 sg13g2_nor2_1 _2682_ (.A(_1646_),
    .B(net595),
    .Y(_1199_));
 sg13g2_nor3_1 _2683_ (.A(_1189_),
    .B(_1196_),
    .C(_1199_),
    .Y(_1200_));
 sg13g2_nand4_1 _2684_ (.B(_1191_),
    .C(_1192_),
    .A(_1183_),
    .Y(_1201_),
    .D(_1200_));
 sg13g2_nand2b_1 _2685_ (.Y(_1202_),
    .B(\input_halfprob2_sng_comparator.bits_b[5] ),
    .A_N(\integrator_a_counter.value_output[8] ));
 sg13g2_nand3b_1 _2686_ (.B(_1201_),
    .C(_1202_),
    .Y(_1203_),
    .A_N(_1198_));
 sg13g2_nand2_1 _2687_ (.Y(_1204_),
    .A(_1085_),
    .B(_1203_));
 sg13g2_inv_1 _2688_ (.Y(_1205_),
    .A(net522));
 sg13g2_nor4_1 _2689_ (.A(\integrator_b_counter.value_output[6] ),
    .B(\integrator_b_counter.value_output[5] ),
    .C(\integrator_b_counter.value_output[4] ),
    .D(\integrator_b_counter.value_output[3] ),
    .Y(_1206_));
 sg13g2_nand3b_1 _2690_ (.B(_1641_),
    .C(_1206_),
    .Y(_1207_),
    .A_N(\integrator_b_counter.value_output[8] ));
 sg13g2_nor4_1 _2691_ (.A(\integrator_b_counter.value_output[2] ),
    .B(\integrator_b_counter.value_output[1] ),
    .C(\integrator_b_counter.value_output[0] ),
    .D(_1207_),
    .Y(_1208_));
 sg13g2_nor2b_1 _2692_ (.A(_0051_),
    .B_N(\integrator_b_counter.value_output[1] ),
    .Y(_1209_));
 sg13g2_nand4_1 _2693_ (.B(net589),
    .C(\integrator_b_counter.value_output[5] ),
    .A(\integrator_b_counter.value_output[7] ),
    .Y(_1210_),
    .D(\integrator_b_counter.value_output[2] ));
 sg13g2_nand4_1 _2694_ (.B(\integrator_b_counter.value_output[3] ),
    .C(\integrator_b_counter.value_output[0] ),
    .A(\integrator_b_counter.value_output[4] ),
    .Y(_1211_),
    .D(_1209_));
 sg13g2_nor2_1 _2695_ (.A(net526),
    .B(_1203_),
    .Y(_1212_));
 sg13g2_o21ai_1 _2696_ (.B1(_1212_),
    .Y(_1213_),
    .A1(_1210_),
    .A2(_1211_));
 sg13g2_o21ai_1 _2697_ (.B1(_1213_),
    .Y(_1214_),
    .A1(net523),
    .A2(_1208_));
 sg13g2_nor2_1 _2698_ (.A(net231),
    .B(net511),
    .Y(_1215_));
 sg13g2_nor2_1 _2699_ (.A(_1642_),
    .B(net523),
    .Y(_1216_));
 sg13g2_xnor2_1 _2700_ (.Y(_1217_),
    .A(_1642_),
    .B(net523));
 sg13g2_inv_1 _2701_ (.Y(_1218_),
    .A(_1217_));
 sg13g2_or2_1 _2702_ (.X(_1219_),
    .B(net522),
    .A(_0045_));
 sg13g2_nand2_1 _2703_ (.Y(_1220_),
    .A(_0045_),
    .B(net522));
 sg13g2_nand2_1 _2704_ (.Y(_1221_),
    .A(\integrator_b_counter.value_output[2] ),
    .B(_1205_));
 sg13g2_xor2_1 _2705_ (.B(net523),
    .A(\integrator_b_counter.value_output[2] ),
    .X(_1222_));
 sg13g2_nand2_1 _2706_ (.Y(_1223_),
    .A(_0044_),
    .B(net523));
 sg13g2_o21ai_1 _2707_ (.B1(_1643_),
    .Y(_1224_),
    .A1(_0044_),
    .A2(net523));
 sg13g2_nand2_1 _2708_ (.Y(_1225_),
    .A(_1223_),
    .B(_1224_));
 sg13g2_nand3b_1 _2709_ (.B(_1223_),
    .C(_1224_),
    .Y(_1226_),
    .A_N(_1222_));
 sg13g2_nand2_1 _2710_ (.Y(_1227_),
    .A(_1221_),
    .B(_1226_));
 sg13g2_nand3_1 _2711_ (.B(_1221_),
    .C(_1226_),
    .A(_1219_),
    .Y(_1228_));
 sg13g2_and2_1 _2712_ (.A(_1220_),
    .B(_1228_),
    .X(_1229_));
 sg13g2_xor2_1 _2713_ (.B(net522),
    .A(_0046_),
    .X(_1230_));
 sg13g2_nand4_1 _2714_ (.B(_1220_),
    .C(_1228_),
    .A(_1218_),
    .Y(_1231_),
    .D(_1230_));
 sg13g2_xor2_1 _2715_ (.B(net522),
    .A(net589),
    .X(_1232_));
 sg13g2_xnor2_1 _2716_ (.Y(_1233_),
    .A(_1641_),
    .B(net522));
 sg13g2_or3_1 _2717_ (.A(_1231_),
    .B(_1232_),
    .C(_1233_),
    .X(_1234_));
 sg13g2_a21o_1 _2718_ (.A2(_0046_),
    .A1(_1642_),
    .B1(net522),
    .X(_1235_));
 sg13g2_o21ai_1 _2719_ (.B1(_1205_),
    .Y(_1236_),
    .A1(\integrator_b_counter.value_output[7] ),
    .A2(net589));
 sg13g2_nand3_1 _2720_ (.B(_1235_),
    .C(_1236_),
    .A(_1234_),
    .Y(_1237_));
 sg13g2_xor2_1 _2721_ (.B(net522),
    .A(net434),
    .X(_1238_));
 sg13g2_xnor2_1 _2722_ (.Y(_1239_),
    .A(_1237_),
    .B(_1238_));
 sg13g2_a21oi_1 _2723_ (.A1(net511),
    .A2(_1239_),
    .Y(_0508_),
    .B1(_1215_));
 sg13g2_a21oi_1 _2724_ (.A1(_1231_),
    .A2(_1235_),
    .Y(_1240_),
    .B1(_1232_));
 sg13g2_a21oi_1 _2725_ (.A1(net589),
    .A2(_1205_),
    .Y(_1241_),
    .B1(_1240_));
 sg13g2_nor2_1 _2726_ (.A(net435),
    .B(net511),
    .Y(_1242_));
 sg13g2_xnor2_1 _2727_ (.Y(_1243_),
    .A(_1233_),
    .B(_1241_));
 sg13g2_a21oi_1 _2728_ (.A1(net511),
    .A2(_1243_),
    .Y(_0507_),
    .B1(_1242_));
 sg13g2_nand3_1 _2729_ (.B(_1232_),
    .C(_1235_),
    .A(_1231_),
    .Y(_1244_));
 sg13g2_nor2b_1 _2730_ (.A(_1240_),
    .B_N(_1244_),
    .Y(_1245_));
 sg13g2_mux2_1 _2731_ (.A0(net589),
    .A1(_1245_),
    .S(net511),
    .X(_0506_));
 sg13g2_a21oi_1 _2732_ (.A1(_1218_),
    .A2(_1229_),
    .Y(_1246_),
    .B1(_1216_));
 sg13g2_xor2_1 _2733_ (.B(_1246_),
    .A(_1230_),
    .X(_1247_));
 sg13g2_nor2_1 _2734_ (.A(net448),
    .B(net511),
    .Y(_1248_));
 sg13g2_a21oi_1 _2735_ (.A1(net512),
    .A2(_1247_),
    .Y(_0505_),
    .B1(_1248_));
 sg13g2_nor2_1 _2736_ (.A(net436),
    .B(net511),
    .Y(_1249_));
 sg13g2_xnor2_1 _2737_ (.Y(_1250_),
    .A(_1218_),
    .B(_1229_));
 sg13g2_a21oi_1 _2738_ (.A1(net511),
    .A2(_1250_),
    .Y(_0504_),
    .B1(_1249_));
 sg13g2_nand2_1 _2739_ (.Y(_1251_),
    .A(_1219_),
    .B(_1220_));
 sg13g2_xnor2_1 _2740_ (.Y(_1252_),
    .A(_1227_),
    .B(_1251_));
 sg13g2_mux2_1 _2741_ (.A0(net437),
    .A1(_1252_),
    .S(net512),
    .X(_0503_));
 sg13g2_xor2_1 _2742_ (.B(_1225_),
    .A(_1222_),
    .X(_1253_));
 sg13g2_mux2_1 _2743_ (.A0(net466),
    .A1(_1253_),
    .S(net512),
    .X(_0502_));
 sg13g2_nor2_1 _2744_ (.A(net387),
    .B(net512),
    .Y(_1254_));
 sg13g2_xnor2_1 _2745_ (.Y(_1255_),
    .A(_0044_),
    .B(net523));
 sg13g2_xnor2_1 _2746_ (.Y(_1256_),
    .A(net57),
    .B(_1255_));
 sg13g2_a21oi_1 _2747_ (.A1(net512),
    .A2(_1256_),
    .Y(_0501_),
    .B1(_1254_));
 sg13g2_nand2_1 _2748_ (.Y(_1257_),
    .A(net57),
    .B(net512));
 sg13g2_o21ai_1 _2749_ (.B1(_1257_),
    .Y(_0500_),
    .A1(_1643_),
    .A2(net512));
 sg13g2_nand2_1 _2750_ (.Y(_1258_),
    .A(_0787_),
    .B(net526));
 sg13g2_inv_1 _2751_ (.Y(_1259_),
    .A(net520));
 sg13g2_or2_1 _2752_ (.X(_1260_),
    .B(\integrator_a_counter.value_output[0] ),
    .A(\integrator_a_counter.value_output[2] ));
 sg13g2_nor4_1 _2753_ (.A(\integrator_a_counter.value_output[8] ),
    .B(\integrator_a_counter.value_output[7] ),
    .C(net590),
    .D(\integrator_a_counter.value_output[3] ),
    .Y(_1261_));
 sg13g2_nor4_1 _2754_ (.A(\integrator_a_counter.value_output[5] ),
    .B(\integrator_a_counter.value_output[4] ),
    .C(\integrator_a_counter.value_output[1] ),
    .D(_1260_),
    .Y(_1262_));
 sg13g2_a21oi_1 _2755_ (.A1(_1261_),
    .A2(_1262_),
    .Y(_1263_),
    .B1(net521));
 sg13g2_nand2b_1 _2756_ (.Y(_1264_),
    .B(\integrator_a_counter.value_output[1] ),
    .A_N(_0054_));
 sg13g2_nand2_1 _2757_ (.Y(_1265_),
    .A(\integrator_a_counter.value_output[7] ),
    .B(net590));
 sg13g2_nand4_1 _2758_ (.B(\integrator_a_counter.value_output[4] ),
    .C(\integrator_a_counter.value_output[3] ),
    .A(\integrator_a_counter.value_output[5] ),
    .Y(_1266_),
    .D(\integrator_a_counter.value_output[2] ));
 sg13g2_nor4_1 _2759_ (.A(_1646_),
    .B(_1264_),
    .C(_1265_),
    .D(_1266_),
    .Y(_1267_));
 sg13g2_nor3_1 _2760_ (.A(_0787_),
    .B(net526),
    .C(_1267_),
    .Y(_1268_));
 sg13g2_or2_1 _2761_ (.X(_1269_),
    .B(_1268_),
    .A(_1263_));
 sg13g2_nor2_1 _2762_ (.A(net243),
    .B(net509),
    .Y(_1270_));
 sg13g2_xor2_1 _2763_ (.B(net520),
    .A(_0043_),
    .X(_1271_));
 sg13g2_nor2_1 _2764_ (.A(_1645_),
    .B(net520),
    .Y(_1272_));
 sg13g2_xnor2_1 _2765_ (.Y(_1273_),
    .A(_1645_),
    .B(net520));
 sg13g2_inv_1 _2766_ (.Y(_1274_),
    .A(_1273_));
 sg13g2_nand2_1 _2767_ (.Y(_1275_),
    .A(_0042_),
    .B(net520));
 sg13g2_or2_1 _2768_ (.X(_1276_),
    .B(net520),
    .A(_0042_));
 sg13g2_nand2_1 _2769_ (.Y(_1277_),
    .A(\integrator_a_counter.value_output[2] ),
    .B(_1259_));
 sg13g2_xor2_1 _2770_ (.B(net521),
    .A(\integrator_a_counter.value_output[2] ),
    .X(_1278_));
 sg13g2_nand2_1 _2771_ (.Y(_1279_),
    .A(_0041_),
    .B(net521));
 sg13g2_o21ai_1 _2772_ (.B1(_1646_),
    .Y(_1280_),
    .A1(_0041_),
    .A2(net521));
 sg13g2_nand2_1 _2773_ (.Y(_1281_),
    .A(_1279_),
    .B(_1280_));
 sg13g2_nand3b_1 _2774_ (.B(_1279_),
    .C(_1280_),
    .Y(_1282_),
    .A_N(_1278_));
 sg13g2_nand2_1 _2775_ (.Y(_1283_),
    .A(_1277_),
    .B(_1282_));
 sg13g2_nand3_1 _2776_ (.B(_1277_),
    .C(_1282_),
    .A(_1276_),
    .Y(_1284_));
 sg13g2_and2_1 _2777_ (.A(_1275_),
    .B(_1284_),
    .X(_1285_));
 sg13g2_nand4_1 _2778_ (.B(_1274_),
    .C(_1275_),
    .A(_1271_),
    .Y(_1286_),
    .D(_1284_));
 sg13g2_xor2_1 _2779_ (.B(net520),
    .A(net590),
    .X(_1287_));
 sg13g2_xnor2_1 _2780_ (.Y(_1288_),
    .A(_1644_),
    .B(net521));
 sg13g2_or3_1 _2781_ (.A(_1286_),
    .B(_1287_),
    .C(_1288_),
    .X(_1289_));
 sg13g2_a21o_1 _2782_ (.A2(_0043_),
    .A1(_1645_),
    .B1(net520),
    .X(_1290_));
 sg13g2_o21ai_1 _2783_ (.B1(_1259_),
    .Y(_1291_),
    .A1(\integrator_a_counter.value_output[7] ),
    .A2(net590));
 sg13g2_nand3_1 _2784_ (.B(_1290_),
    .C(_1291_),
    .A(_1289_),
    .Y(_1292_));
 sg13g2_xor2_1 _2785_ (.B(net521),
    .A(net420),
    .X(_1293_));
 sg13g2_xnor2_1 _2786_ (.Y(_1294_),
    .A(_1292_),
    .B(_1293_));
 sg13g2_a21oi_1 _2787_ (.A1(_1269_),
    .A2(_1294_),
    .Y(_0499_),
    .B1(_1270_));
 sg13g2_a21oi_1 _2788_ (.A1(_1286_),
    .A2(_1290_),
    .Y(_1295_),
    .B1(_1287_));
 sg13g2_a21oi_1 _2789_ (.A1(net590),
    .A2(_1259_),
    .Y(_1296_),
    .B1(_1295_));
 sg13g2_xnor2_1 _2790_ (.Y(_1297_),
    .A(_1288_),
    .B(_1296_));
 sg13g2_nor2_1 _2791_ (.A(net443),
    .B(net509),
    .Y(_1298_));
 sg13g2_a21oi_1 _2792_ (.A1(net509),
    .A2(_1297_),
    .Y(_0498_),
    .B1(_1298_));
 sg13g2_nor2_1 _2793_ (.A(net590),
    .B(net510),
    .Y(_1299_));
 sg13g2_nand3_1 _2794_ (.B(_1287_),
    .C(_1290_),
    .A(_1286_),
    .Y(_1300_));
 sg13g2_nand2b_1 _2795_ (.Y(_1301_),
    .B(_1300_),
    .A_N(_1295_));
 sg13g2_a21oi_1 _2796_ (.A1(net510),
    .A2(_1301_),
    .Y(_0497_),
    .B1(_1299_));
 sg13g2_a21oi_1 _2797_ (.A1(_1274_),
    .A2(_1285_),
    .Y(_1302_),
    .B1(_1272_));
 sg13g2_xor2_1 _2798_ (.B(_1302_),
    .A(_1271_),
    .X(_1303_));
 sg13g2_nor2_1 _2799_ (.A(net464),
    .B(net510),
    .Y(_1304_));
 sg13g2_a21oi_1 _2800_ (.A1(net510),
    .A2(_1303_),
    .Y(_0496_),
    .B1(_1304_));
 sg13g2_nor2_1 _2801_ (.A(net446),
    .B(net510),
    .Y(_1305_));
 sg13g2_xnor2_1 _2802_ (.Y(_1306_),
    .A(_1274_),
    .B(_1285_));
 sg13g2_a21oi_1 _2803_ (.A1(net510),
    .A2(_1306_),
    .Y(_0495_),
    .B1(_1305_));
 sg13g2_nand2_1 _2804_ (.Y(_1307_),
    .A(_1275_),
    .B(_1276_));
 sg13g2_xnor2_1 _2805_ (.Y(_1308_),
    .A(_1283_),
    .B(_1307_));
 sg13g2_mux2_1 _2806_ (.A0(net474),
    .A1(_1308_),
    .S(net510),
    .X(_0494_));
 sg13g2_xor2_1 _2807_ (.B(_1281_),
    .A(_1278_),
    .X(_1309_));
 sg13g2_mux2_1 _2808_ (.A0(net480),
    .A1(_1309_),
    .S(net509),
    .X(_0493_));
 sg13g2_nor2_1 _2809_ (.A(net397),
    .B(net509),
    .Y(_1310_));
 sg13g2_xnor2_1 _2810_ (.Y(_1311_),
    .A(_0041_),
    .B(net521));
 sg13g2_xnor2_1 _2811_ (.Y(_1312_),
    .A(net45),
    .B(_1311_));
 sg13g2_a21oi_1 _2812_ (.A1(net509),
    .A2(_1312_),
    .Y(_0492_),
    .B1(_1310_));
 sg13g2_nand2_1 _2813_ (.Y(_1313_),
    .A(net45),
    .B(net509));
 sg13g2_o21ai_1 _2814_ (.B1(_1313_),
    .Y(_0491_),
    .A1(_1646_),
    .A2(net509));
 sg13g2_mux2_1 _2815_ (.A0(net73),
    .A1(net189),
    .S(net566),
    .X(_0490_));
 sg13g2_nor2_1 _2816_ (.A(net318),
    .B(net566),
    .Y(_1314_));
 sg13g2_a21oi_1 _2817_ (.A1(_1647_),
    .A2(net566),
    .Y(_0489_),
    .B1(_1314_));
 sg13g2_mux2_1 _2818_ (.A0(net235),
    .A1(\test_integrator_b_counter.value_output[6] ),
    .S(net566),
    .X(_0488_));
 sg13g2_mux2_1 _2819_ (.A0(net223),
    .A1(\test_integrator_b_counter.value_output[5] ),
    .S(net566),
    .X(_0487_));
 sg13g2_nor2_1 _2820_ (.A(net204),
    .B(net567),
    .Y(_1315_));
 sg13g2_a21oi_1 _2821_ (.A1(_1648_),
    .A2(net567),
    .Y(_0486_),
    .B1(_1315_));
 sg13g2_nor2_1 _2822_ (.A(net217),
    .B(net567),
    .Y(_1316_));
 sg13g2_a21oi_1 _2823_ (.A1(_1649_),
    .A2(net567),
    .Y(_0485_),
    .B1(_1316_));
 sg13g2_mux2_1 _2824_ (.A0(net250),
    .A1(net591),
    .S(net567),
    .X(_0484_));
 sg13g2_mux2_1 _2825_ (.A0(net177),
    .A1(net592),
    .S(net566),
    .X(_0483_));
 sg13g2_nor2_1 _2826_ (.A(net174),
    .B(net566),
    .Y(_1317_));
 sg13g2_a21oi_1 _2827_ (.A1(_1650_),
    .A2(net566),
    .Y(_0482_),
    .B1(_1317_));
 sg13g2_nand2_1 _2828_ (.Y(_1318_),
    .A(\system_integrator_b_output.counter[0] ),
    .B(net320));
 sg13g2_nor3_2 _2829_ (.A(\system_integrator_b_output.counter[1] ),
    .B(\system_integrator_b_output.counter[2] ),
    .C(_1318_),
    .Y(_1319_));
 sg13g2_nor4_2 _2830_ (.A(\system_integrator_b_output.counter[0] ),
    .B(\system_integrator_b_output.counter[1] ),
    .C(\system_integrator_b_output.counter[2] ),
    .Y(_1320_),
    .D(\system_integrator_b_output.counter[3] ));
 sg13g2_a22oi_1 _2831_ (.Y(_1321_),
    .B1(net558),
    .B2(net39),
    .A2(net544),
    .A1(\system_integrator_b_output.bitseq[7] ));
 sg13g2_inv_1 _2832_ (.Y(_0481_),
    .A(net40));
 sg13g2_nand2_1 _2833_ (.Y(_1322_),
    .A(net69),
    .B(net544));
 sg13g2_nand2b_1 _2834_ (.Y(_1323_),
    .B(net559),
    .A_N(\system_integrator_b_output.input_bits[7] ));
 sg13g2_o21ai_1 _2835_ (.B1(_1323_),
    .Y(_1324_),
    .A1(\system_integrator_b_output.bitseq[7] ),
    .A2(net558));
 sg13g2_o21ai_1 _2836_ (.B1(_1322_),
    .Y(_0480_),
    .A1(net544),
    .A2(_1324_));
 sg13g2_nand2_1 _2837_ (.Y(_1325_),
    .A(net126),
    .B(net545));
 sg13g2_nand2b_1 _2838_ (.Y(_1326_),
    .B(net559),
    .A_N(\system_integrator_b_output.input_bits[6] ));
 sg13g2_o21ai_1 _2839_ (.B1(_1326_),
    .Y(_1327_),
    .A1(net69),
    .A2(net558));
 sg13g2_o21ai_1 _2840_ (.B1(_1325_),
    .Y(_0479_),
    .A1(net544),
    .A2(_1327_));
 sg13g2_nand2_1 _2841_ (.Y(_1328_),
    .A(net209),
    .B(net545));
 sg13g2_nand2b_1 _2842_ (.Y(_1329_),
    .B(net558),
    .A_N(\system_integrator_b_output.input_bits[5] ));
 sg13g2_o21ai_1 _2843_ (.B1(_1329_),
    .Y(_1330_),
    .A1(net126),
    .A2(net558));
 sg13g2_o21ai_1 _2844_ (.B1(_1328_),
    .Y(_0478_),
    .A1(net544),
    .A2(_1330_));
 sg13g2_nand2_1 _2845_ (.Y(_1331_),
    .A(net112),
    .B(net544));
 sg13g2_nand2b_1 _2846_ (.Y(_1332_),
    .B(net558),
    .A_N(\system_integrator_b_output.input_bits[4] ));
 sg13g2_o21ai_1 _2847_ (.B1(_1332_),
    .Y(_1333_),
    .A1(\system_integrator_b_output.bitseq[4] ),
    .A2(net558));
 sg13g2_o21ai_1 _2848_ (.B1(_1331_),
    .Y(_0477_),
    .A1(net544),
    .A2(_1333_));
 sg13g2_nand2_1 _2849_ (.Y(_1334_),
    .A(net160),
    .B(_1319_));
 sg13g2_nand2b_1 _2850_ (.Y(_1335_),
    .B(net559),
    .A_N(\system_integrator_b_output.input_bits[3] ));
 sg13g2_o21ai_1 _2851_ (.B1(_1335_),
    .Y(_1336_),
    .A1(net112),
    .A2(net558));
 sg13g2_o21ai_1 _2852_ (.B1(net161),
    .Y(_0476_),
    .A1(net545),
    .A2(_1336_));
 sg13g2_nand2_1 _2853_ (.Y(_1337_),
    .A(net143),
    .B(_1319_));
 sg13g2_nand2b_1 _2854_ (.Y(_1338_),
    .B(_1320_),
    .A_N(\system_integrator_b_output.input_bits[2] ));
 sg13g2_o21ai_1 _2855_ (.B1(_1338_),
    .Y(_1339_),
    .A1(\system_integrator_b_output.bitseq[2] ),
    .A2(net559));
 sg13g2_o21ai_1 _2856_ (.B1(net144),
    .Y(_0475_),
    .A1(net545),
    .A2(_1339_));
 sg13g2_nand2_1 _2857_ (.Y(_1340_),
    .A(net104),
    .B(net545));
 sg13g2_nand2b_1 _2858_ (.Y(_1341_),
    .B(net559),
    .A_N(\system_integrator_b_output.input_bits[1] ));
 sg13g2_o21ai_1 _2859_ (.B1(_1341_),
    .Y(_1342_),
    .A1(\system_integrator_b_output.bitseq[1] ),
    .A2(_1320_));
 sg13g2_o21ai_1 _2860_ (.B1(_1340_),
    .Y(_0474_),
    .A1(net545),
    .A2(_1342_));
 sg13g2_nand2_1 _2861_ (.Y(_1343_),
    .A(_1616_),
    .B(\input_halfprob2_sng_comparator.bits_b[5] ));
 sg13g2_nor2_1 _2862_ (.A(\test_integrator_a_counter.value_output[1] ),
    .B(_0640_),
    .Y(_1344_));
 sg13g2_nand2_1 _2863_ (.Y(_1345_),
    .A(\test_integrator_a_counter.value_output[0] ),
    .B(_0641_));
 sg13g2_a22oi_1 _2864_ (.Y(_1346_),
    .B1(_0640_),
    .B2(\test_integrator_a_counter.value_output[1] ),
    .A2(_0639_),
    .A1(\test_integrator_a_counter.value_output[2] ));
 sg13g2_o21ai_1 _2865_ (.B1(_1346_),
    .Y(_1347_),
    .A1(_1344_),
    .A2(_1345_));
 sg13g2_a22oi_1 _2866_ (.Y(_1348_),
    .B1(\input_halfprob1_sng_comparator.bits_b[0] ),
    .B2(_1622_),
    .A2(\input_halfprob1_sng_comparator.bits_b[1] ),
    .A1(_1621_));
 sg13g2_nand2b_1 _2867_ (.Y(_1349_),
    .B(\test_integrator_a_counter.value_output[3] ),
    .A_N(\input_halfprob1_sng_comparator.bits_b[1] ));
 sg13g2_o21ai_1 _2868_ (.B1(_1349_),
    .Y(_1350_),
    .A1(_1620_),
    .A2(\input_halfprob2_sng_comparator.bits_b[1] ));
 sg13g2_a21oi_1 _2869_ (.A1(_1347_),
    .A2(_1348_),
    .Y(_1351_),
    .B1(_1350_));
 sg13g2_a221oi_1 _2870_ (.B2(_1620_),
    .C1(_1351_),
    .B1(\input_halfprob2_sng_comparator.bits_b[1] ),
    .A1(_1619_),
    .Y(_1352_),
    .A2(\input_halfprob2_sng_comparator.bits_b[2] ));
 sg13g2_a221oi_1 _2871_ (.B2(\test_integrator_a_counter.value_output[5] ),
    .C1(_1352_),
    .B1(_0638_),
    .A1(\test_integrator_a_counter.value_output[6] ),
    .Y(_1353_),
    .A2(_0637_));
 sg13g2_a221oi_1 _2872_ (.B2(_1618_),
    .C1(_1353_),
    .B1(\input_halfprob2_sng_comparator.bits_b[3] ),
    .A1(_1617_),
    .Y(_1354_),
    .A2(\input_halfprob2_sng_comparator.bits_b[4] ));
 sg13g2_nand2b_1 _2873_ (.Y(_1355_),
    .B(\test_integrator_a_counter.value_output[7] ),
    .A_N(\input_halfprob2_sng_comparator.bits_b[4] ));
 sg13g2_o21ai_1 _2874_ (.B1(_1355_),
    .Y(_1356_),
    .A1(_1616_),
    .A2(\input_halfprob2_sng_comparator.bits_b[5] ));
 sg13g2_o21ai_1 _2875_ (.B1(_1343_),
    .Y(_1357_),
    .A1(_1354_),
    .A2(_1356_));
 sg13g2_nand3_1 _2876_ (.B(\test_integrator_b_counter.value_output[1] ),
    .C(\test_integrator_b_counter.value_output[0] ),
    .A(net591),
    .Y(_1358_));
 sg13g2_nor2_1 _2877_ (.A(_1649_),
    .B(_1358_),
    .Y(_1359_));
 sg13g2_and3_1 _2878_ (.X(_1360_),
    .A(\test_integrator_b_counter.value_output[5] ),
    .B(\test_integrator_b_counter.value_output[4] ),
    .C(_1359_));
 sg13g2_nor2b_1 _2879_ (.A(net593),
    .B_N(\test_integrator_b_counter.value_output[8] ),
    .Y(_1361_));
 sg13g2_nand4_1 _2880_ (.B(\test_integrator_b_counter.value_output[6] ),
    .C(_1360_),
    .A(\test_integrator_b_counter.value_output[7] ),
    .Y(_1362_),
    .D(_1361_));
 sg13g2_nor2b_1 _2881_ (.A(_0819_),
    .B_N(_1362_),
    .Y(_1363_));
 sg13g2_nand2b_1 _2882_ (.Y(_1364_),
    .B(_1363_),
    .A_N(_1357_));
 sg13g2_nand2_1 _2883_ (.Y(_1365_),
    .A(net495),
    .B(net581));
 sg13g2_and2_2 _2884_ (.A(_0819_),
    .B(_1357_),
    .X(_1366_));
 sg13g2_nand2_2 _2885_ (.Y(_1367_),
    .A(_0819_),
    .B(_1357_));
 sg13g2_nand2_1 _2886_ (.Y(_1368_),
    .A(_1365_),
    .B(_1366_));
 sg13g2_o21ai_1 _2887_ (.B1(_1368_),
    .Y(_1369_),
    .A1(_1364_),
    .A2(_1365_));
 sg13g2_a21oi_1 _2888_ (.A1(_1650_),
    .A2(_1364_),
    .Y(_0473_),
    .B1(_1369_));
 sg13g2_nand2_1 _2889_ (.Y(_1370_),
    .A(\system_integrator_a_output.counter[0] ),
    .B(net308));
 sg13g2_nor3_2 _2890_ (.A(\system_integrator_a_output.counter[1] ),
    .B(\system_integrator_a_output.counter[2] ),
    .C(_1370_),
    .Y(_1371_));
 sg13g2_nor4_2 _2891_ (.A(\system_integrator_a_output.counter[0] ),
    .B(\system_integrator_a_output.counter[1] ),
    .C(\system_integrator_a_output.counter[2] ),
    .Y(_1372_),
    .D(\system_integrator_a_output.counter[3] ));
 sg13g2_a22oi_1 _2892_ (.Y(_1373_),
    .B1(net556),
    .B2(net52),
    .A2(net543),
    .A1(\system_integrator_a_output.bitseq[7] ));
 sg13g2_inv_1 _2893_ (.Y(_0472_),
    .A(net53));
 sg13g2_nand2_1 _2894_ (.Y(_1374_),
    .A(net106),
    .B(net543));
 sg13g2_nand2b_1 _2895_ (.Y(_1375_),
    .B(net556),
    .A_N(\system_integrator_a_output.input_bits[7] ));
 sg13g2_o21ai_1 _2896_ (.B1(_1375_),
    .Y(_1376_),
    .A1(\system_integrator_a_output.bitseq[7] ),
    .A2(net556));
 sg13g2_o21ai_1 _2897_ (.B1(_1374_),
    .Y(_0471_),
    .A1(net543),
    .A2(_1376_));
 sg13g2_nand2_1 _2898_ (.Y(_1377_),
    .A(net75),
    .B(net543));
 sg13g2_nand2b_1 _2899_ (.Y(_1378_),
    .B(net556),
    .A_N(\system_integrator_a_output.input_bits[6] ));
 sg13g2_o21ai_1 _2900_ (.B1(_1378_),
    .Y(_1379_),
    .A1(\system_integrator_a_output.bitseq[6] ),
    .A2(net556));
 sg13g2_o21ai_1 _2901_ (.B1(_1377_),
    .Y(_0470_),
    .A1(net543),
    .A2(_1379_));
 sg13g2_nand2_1 _2902_ (.Y(_1380_),
    .A(net93),
    .B(net543));
 sg13g2_nand2b_1 _2903_ (.Y(_1381_),
    .B(net557),
    .A_N(\system_integrator_a_output.input_bits[5] ));
 sg13g2_o21ai_1 _2904_ (.B1(_1381_),
    .Y(_1382_),
    .A1(net75),
    .A2(net556));
 sg13g2_o21ai_1 _2905_ (.B1(_1380_),
    .Y(_0469_),
    .A1(net543),
    .A2(_1382_));
 sg13g2_nand2_1 _2906_ (.Y(_1383_),
    .A(net169),
    .B(net542));
 sg13g2_nand2b_1 _2907_ (.Y(_1384_),
    .B(net556),
    .A_N(\system_integrator_a_output.input_bits[4] ));
 sg13g2_o21ai_1 _2908_ (.B1(_1384_),
    .Y(_1385_),
    .A1(net93),
    .A2(net556));
 sg13g2_o21ai_1 _2909_ (.B1(_1383_),
    .Y(_0468_),
    .A1(net542),
    .A2(_1385_));
 sg13g2_nand2_1 _2910_ (.Y(_1386_),
    .A(net148),
    .B(net542));
 sg13g2_nand2b_1 _2911_ (.Y(_1387_),
    .B(_1372_),
    .A_N(\system_integrator_a_output.input_bits[3] ));
 sg13g2_o21ai_1 _2912_ (.B1(_1387_),
    .Y(_1388_),
    .A1(\system_integrator_a_output.bitseq[3] ),
    .A2(net557));
 sg13g2_o21ai_1 _2913_ (.B1(_1386_),
    .Y(_0467_),
    .A1(net542),
    .A2(_1388_));
 sg13g2_nand2_1 _2914_ (.Y(_1389_),
    .A(net71),
    .B(net542));
 sg13g2_nand2b_1 _2915_ (.Y(_1390_),
    .B(_1372_),
    .A_N(\system_integrator_a_output.input_bits[2] ));
 sg13g2_o21ai_1 _2916_ (.B1(_1390_),
    .Y(_1391_),
    .A1(\system_integrator_a_output.bitseq[2] ),
    .A2(net557));
 sg13g2_o21ai_1 _2917_ (.B1(_1389_),
    .Y(_0466_),
    .A1(net542),
    .A2(_1391_));
 sg13g2_nand2_1 _2918_ (.Y(_1392_),
    .A(net77),
    .B(_1371_));
 sg13g2_nand2b_1 _2919_ (.Y(_1393_),
    .B(net557),
    .A_N(\system_integrator_a_output.input_bits[1] ));
 sg13g2_o21ai_1 _2920_ (.B1(_1393_),
    .Y(_1394_),
    .A1(net71),
    .A2(net557));
 sg13g2_o21ai_1 _2921_ (.B1(net78),
    .Y(_0465_),
    .A1(net542),
    .A2(_1394_));
 sg13g2_nand2_1 _2922_ (.Y(_1395_),
    .A(\test_integrator_b_output.counter[0] ),
    .B(net392));
 sg13g2_nor3_2 _2923_ (.A(\test_integrator_b_output.counter[1] ),
    .B(\test_integrator_b_output.counter[2] ),
    .C(_1395_),
    .Y(_1396_));
 sg13g2_nor4_2 _2924_ (.A(\test_integrator_b_output.counter[0] ),
    .B(\test_integrator_b_output.counter[1] ),
    .C(\test_integrator_b_output.counter[2] ),
    .Y(_1397_),
    .D(\test_integrator_b_output.counter[3] ));
 sg13g2_a22oi_1 _2925_ (.Y(_1398_),
    .B1(net555),
    .B2(net73),
    .A2(net541),
    .A1(\test_integrator_b_output.bitseq[7] ));
 sg13g2_inv_1 _2926_ (.Y(_0464_),
    .A(net74));
 sg13g2_nand2_1 _2927_ (.Y(_1399_),
    .A(net61),
    .B(net541));
 sg13g2_nand2b_1 _2928_ (.Y(_1400_),
    .B(net555),
    .A_N(\test_integrator_b_output.input_bits[7] ));
 sg13g2_o21ai_1 _2929_ (.B1(_1400_),
    .Y(_1401_),
    .A1(\test_integrator_b_output.bitseq[7] ),
    .A2(net555));
 sg13g2_o21ai_1 _2930_ (.B1(_1399_),
    .Y(_0463_),
    .A1(net541),
    .A2(_1401_));
 sg13g2_nand2_1 _2931_ (.Y(_1402_),
    .A(net122),
    .B(net540));
 sg13g2_nand2b_1 _2932_ (.Y(_1403_),
    .B(net555),
    .A_N(\test_integrator_b_output.input_bits[6] ));
 sg13g2_o21ai_1 _2933_ (.B1(_1403_),
    .Y(_1404_),
    .A1(net61),
    .A2(net555));
 sg13g2_o21ai_1 _2934_ (.B1(_1402_),
    .Y(_0462_),
    .A1(net541),
    .A2(_1404_));
 sg13g2_nand2_1 _2935_ (.Y(_1405_),
    .A(net184),
    .B(net540));
 sg13g2_nand2b_1 _2936_ (.Y(_1406_),
    .B(net554),
    .A_N(\test_integrator_b_output.input_bits[5] ));
 sg13g2_o21ai_1 _2937_ (.B1(_1406_),
    .Y(_1407_),
    .A1(net122),
    .A2(net554));
 sg13g2_o21ai_1 _2938_ (.B1(_1405_),
    .Y(_0461_),
    .A1(net540),
    .A2(_1407_));
 sg13g2_nand2_1 _2939_ (.Y(_1408_),
    .A(net82),
    .B(net540));
 sg13g2_nand2b_1 _2940_ (.Y(_1409_),
    .B(net554),
    .A_N(\test_integrator_b_output.input_bits[4] ));
 sg13g2_o21ai_1 _2941_ (.B1(_1409_),
    .Y(_1410_),
    .A1(\test_integrator_b_output.bitseq[4] ),
    .A2(_1397_));
 sg13g2_o21ai_1 _2942_ (.B1(_1408_),
    .Y(_0460_),
    .A1(_1396_),
    .A2(_1410_));
 sg13g2_nand2_1 _2943_ (.Y(_1411_),
    .A(net158),
    .B(net540));
 sg13g2_nand2b_1 _2944_ (.Y(_1412_),
    .B(net554),
    .A_N(\test_integrator_b_output.input_bits[3] ));
 sg13g2_o21ai_1 _2945_ (.B1(_1412_),
    .Y(_1413_),
    .A1(net82),
    .A2(_1397_));
 sg13g2_o21ai_1 _2946_ (.B1(_1411_),
    .Y(_0459_),
    .A1(_1396_),
    .A2(_1413_));
 sg13g2_nand2_1 _2947_ (.Y(_1414_),
    .A(net139),
    .B(net540));
 sg13g2_nand2b_1 _2948_ (.Y(_1415_),
    .B(net554),
    .A_N(\test_integrator_b_output.input_bits[2] ));
 sg13g2_o21ai_1 _2949_ (.B1(_1415_),
    .Y(_1416_),
    .A1(\test_integrator_b_output.bitseq[2] ),
    .A2(net554));
 sg13g2_o21ai_1 _2950_ (.B1(_1414_),
    .Y(_0458_),
    .A1(net540),
    .A2(_1416_));
 sg13g2_nand2_1 _2951_ (.Y(_1417_),
    .A(net124),
    .B(net541));
 sg13g2_nand2b_1 _2952_ (.Y(_1418_),
    .B(net554),
    .A_N(\test_integrator_b_output.input_bits[1] ));
 sg13g2_o21ai_1 _2953_ (.B1(_1418_),
    .Y(_1419_),
    .A1(\test_integrator_b_output.bitseq[1] ),
    .A2(net554));
 sg13g2_o21ai_1 _2954_ (.B1(_1417_),
    .Y(_0457_),
    .A1(net541),
    .A2(_1419_));
 sg13g2_and2_1 _2955_ (.A(_1364_),
    .B(_1367_),
    .X(_1420_));
 sg13g2_inv_1 _2956_ (.Y(_1421_),
    .A(_1420_));
 sg13g2_nand2_1 _2957_ (.Y(_1422_),
    .A(net189),
    .B(net508));
 sg13g2_nor3_1 _2958_ (.A(\test_integrator_b_counter.value_output[3] ),
    .B(net591),
    .C(net592),
    .Y(_1423_));
 sg13g2_and2_1 _2959_ (.A(_1648_),
    .B(_1423_),
    .X(_1424_));
 sg13g2_nand2b_1 _2960_ (.Y(_1425_),
    .B(_1424_),
    .A_N(\test_integrator_b_counter.value_output[5] ));
 sg13g2_or3_1 _2961_ (.A(\test_integrator_b_counter.value_output[6] ),
    .B(_1367_),
    .C(_1425_),
    .X(_1426_));
 sg13g2_nand4_1 _2962_ (.B(\test_integrator_b_counter.value_output[6] ),
    .C(_1360_),
    .A(\test_integrator_b_counter.value_output[7] ),
    .Y(_1427_),
    .D(_1367_));
 sg13g2_o21ai_1 _2963_ (.B1(_1427_),
    .Y(_1428_),
    .A1(\test_integrator_b_counter.value_output[7] ),
    .A2(_1426_));
 sg13g2_and2_1 _2964_ (.A(_0658_),
    .B(_1428_),
    .X(_1429_));
 sg13g2_nor2_2 _2965_ (.A(net593),
    .B(net508),
    .Y(_1430_));
 sg13g2_nand2_2 _2966_ (.Y(_1431_),
    .A(net581),
    .B(_1421_));
 sg13g2_o21ai_1 _2967_ (.B1(_1430_),
    .Y(_1432_),
    .A1(_0658_),
    .A2(_1428_));
 sg13g2_o21ai_1 _2968_ (.B1(_1422_),
    .Y(_0456_),
    .A1(_1429_),
    .A2(net432));
 sg13g2_nand2b_1 _2969_ (.Y(_1433_),
    .B(_1360_),
    .A_N(net372));
 sg13g2_o21ai_1 _2970_ (.B1(_1426_),
    .Y(_1434_),
    .A1(_1366_),
    .A2(_1433_));
 sg13g2_xor2_1 _2971_ (.B(_1434_),
    .A(net384),
    .X(_1435_));
 sg13g2_nand2_1 _2972_ (.Y(_1436_),
    .A(\test_integrator_b_counter.value_output[7] ),
    .B(net508));
 sg13g2_o21ai_1 _2973_ (.B1(_1436_),
    .Y(_0455_),
    .A1(_1431_),
    .A2(_1435_));
 sg13g2_nand2_1 _2974_ (.Y(_1437_),
    .A(\test_integrator_b_counter.value_output[6] ),
    .B(net508));
 sg13g2_nor2_1 _2975_ (.A(_1367_),
    .B(_1425_),
    .Y(_1438_));
 sg13g2_a21oi_1 _2976_ (.A1(_1360_),
    .A2(_1367_),
    .Y(_1439_),
    .B1(_1438_));
 sg13g2_xnor2_1 _2977_ (.Y(_1440_),
    .A(net372),
    .B(_1439_));
 sg13g2_o21ai_1 _2978_ (.B1(_1437_),
    .Y(_0454_),
    .A1(_1431_),
    .A2(_1440_));
 sg13g2_nand2_1 _2979_ (.Y(_1441_),
    .A(\test_integrator_b_counter.value_output[5] ),
    .B(net508));
 sg13g2_and2_1 _2980_ (.A(_1359_),
    .B(_1367_),
    .X(_1442_));
 sg13g2_a22oi_1 _2981_ (.Y(_1443_),
    .B1(_1442_),
    .B2(_0657_),
    .A2(_1424_),
    .A1(_1366_));
 sg13g2_xnor2_1 _2982_ (.Y(_1444_),
    .A(net297),
    .B(_1443_));
 sg13g2_o21ai_1 _2983_ (.B1(_1441_),
    .Y(_0453_),
    .A1(_1431_),
    .A2(net298));
 sg13g2_nand2_1 _2984_ (.Y(_1445_),
    .A(net399),
    .B(net508));
 sg13g2_a21oi_1 _2985_ (.A1(_1366_),
    .A2(_1423_),
    .Y(_1446_),
    .B1(_1442_));
 sg13g2_and2_1 _2986_ (.A(_0036_),
    .B(_1446_),
    .X(_1447_));
 sg13g2_o21ai_1 _2987_ (.B1(_1430_),
    .Y(_1448_),
    .A1(_0036_),
    .A2(_1446_));
 sg13g2_o21ai_1 _2988_ (.B1(_1445_),
    .Y(_0452_),
    .A1(_1447_),
    .A2(_1448_));
 sg13g2_nand2_1 _2989_ (.Y(_1449_),
    .A(\test_integrator_b_counter.value_output[3] ),
    .B(net508));
 sg13g2_nand2_1 _2990_ (.Y(_1450_),
    .A(_1358_),
    .B(_1367_));
 sg13g2_o21ai_1 _2991_ (.B1(_1366_),
    .Y(_1451_),
    .A1(net591),
    .A2(net592));
 sg13g2_nand2_1 _2992_ (.Y(_1452_),
    .A(_1450_),
    .B(_1451_));
 sg13g2_and2_1 _2993_ (.A(net395),
    .B(_1452_),
    .X(_1453_));
 sg13g2_o21ai_1 _2994_ (.B1(_1430_),
    .Y(_1454_),
    .A1(net395),
    .A2(_1452_));
 sg13g2_o21ai_1 _2995_ (.B1(_1449_),
    .Y(_0451_),
    .A1(_1453_),
    .A2(_1454_));
 sg13g2_xnor2_1 _2996_ (.Y(_1455_),
    .A(net591),
    .B(net592));
 sg13g2_a21oi_1 _2997_ (.A1(net592),
    .A2(\test_integrator_b_counter.value_output[0] ),
    .Y(_1456_),
    .B1(net591));
 sg13g2_nor2_1 _2998_ (.A(_1450_),
    .B(_1456_),
    .Y(_1457_));
 sg13g2_a21oi_1 _2999_ (.A1(_1366_),
    .A2(_1455_),
    .Y(_1458_),
    .B1(_1457_));
 sg13g2_nand2_1 _3000_ (.Y(_1459_),
    .A(net591),
    .B(net508));
 sg13g2_o21ai_1 _3001_ (.B1(_1459_),
    .Y(_0450_),
    .A1(_1431_),
    .A2(_1458_));
 sg13g2_o21ai_1 _3002_ (.B1(_1367_),
    .Y(_1460_),
    .A1(_1650_),
    .A2(_1364_));
 sg13g2_xnor2_1 _3003_ (.Y(_1461_),
    .A(net592),
    .B(_1460_));
 sg13g2_a21oi_1 _3004_ (.A1(net593),
    .A2(_1421_),
    .Y(_0449_),
    .B1(_1461_));
 sg13g2_nand2_1 _3005_ (.Y(_1462_),
    .A(\integrator_c_output.counter[0] ),
    .B(net303));
 sg13g2_nor3_1 _3006_ (.A(\integrator_c_output.counter[1] ),
    .B(\integrator_c_output.counter[2] ),
    .C(_1462_),
    .Y(_1463_));
 sg13g2_nor4_2 _3007_ (.A(\integrator_c_output.counter[0] ),
    .B(\integrator_c_output.counter[1] ),
    .C(\integrator_c_output.counter[2] ),
    .Y(_1464_),
    .D(\integrator_c_output.counter[3] ));
 sg13g2_a22oi_1 _3008_ (.Y(_1465_),
    .B1(net553),
    .B2(net165),
    .A2(net539),
    .A1(\integrator_c_output.bitseq[7] ));
 sg13g2_inv_1 _3009_ (.Y(_0448_),
    .A(net166));
 sg13g2_nand2_1 _3010_ (.Y(_1466_),
    .A(net137),
    .B(net539));
 sg13g2_nand2b_1 _3011_ (.Y(_1467_),
    .B(net553),
    .A_N(\integrator_c_output.input_bits[7] ));
 sg13g2_o21ai_1 _3012_ (.B1(_1467_),
    .Y(_1468_),
    .A1(\integrator_c_output.bitseq[7] ),
    .A2(net553));
 sg13g2_o21ai_1 _3013_ (.B1(_1466_),
    .Y(_0447_),
    .A1(net539),
    .A2(_1468_));
 sg13g2_nand2_1 _3014_ (.Y(_1469_),
    .A(net63),
    .B(net539));
 sg13g2_nand2b_1 _3015_ (.Y(_1470_),
    .B(net553),
    .A_N(\integrator_c_output.input_bits[6] ));
 sg13g2_o21ai_1 _3016_ (.B1(_1470_),
    .Y(_1471_),
    .A1(\integrator_c_output.bitseq[6] ),
    .A2(net553));
 sg13g2_o21ai_1 _3017_ (.B1(_1469_),
    .Y(_0446_),
    .A1(net539),
    .A2(_1471_));
 sg13g2_nand2_1 _3018_ (.Y(_1472_),
    .A(net190),
    .B(net538));
 sg13g2_nand2b_1 _3019_ (.Y(_1473_),
    .B(net553),
    .A_N(\integrator_c_output.input_bits[5] ));
 sg13g2_o21ai_1 _3020_ (.B1(_1473_),
    .Y(_1474_),
    .A1(net63),
    .A2(net553));
 sg13g2_o21ai_1 _3021_ (.B1(_1472_),
    .Y(_0445_),
    .A1(net539),
    .A2(_1474_));
 sg13g2_nand2_1 _3022_ (.Y(_1475_),
    .A(net152),
    .B(net538));
 sg13g2_nand2b_1 _3023_ (.Y(_1476_),
    .B(net552),
    .A_N(\integrator_c_output.input_bits[4] ));
 sg13g2_o21ai_1 _3024_ (.B1(_1476_),
    .Y(_1477_),
    .A1(\integrator_c_output.bitseq[4] ),
    .A2(_1464_));
 sg13g2_o21ai_1 _3025_ (.B1(_1475_),
    .Y(_0444_),
    .A1(net538),
    .A2(_1477_));
 sg13g2_nand2_1 _3026_ (.Y(_1478_),
    .A(net163),
    .B(net538));
 sg13g2_nand2b_1 _3027_ (.Y(_1479_),
    .B(net552),
    .A_N(\integrator_c_output.input_bits[3] ));
 sg13g2_o21ai_1 _3028_ (.B1(_1479_),
    .Y(_1480_),
    .A1(net152),
    .A2(net552));
 sg13g2_o21ai_1 _3029_ (.B1(_1478_),
    .Y(_0443_),
    .A1(_1463_),
    .A2(_1480_));
 sg13g2_nand2_1 _3030_ (.Y(_1481_),
    .A(net100),
    .B(net538));
 sg13g2_nand2b_1 _3031_ (.Y(_1482_),
    .B(net552),
    .A_N(\integrator_c_output.input_bits[2] ));
 sg13g2_o21ai_1 _3032_ (.B1(_1482_),
    .Y(_1483_),
    .A1(\integrator_c_output.bitseq[2] ),
    .A2(net552));
 sg13g2_o21ai_1 _3033_ (.B1(_1481_),
    .Y(_0442_),
    .A1(net538),
    .A2(_1483_));
 sg13g2_nand2_1 _3034_ (.Y(_1484_),
    .A(net65),
    .B(net538));
 sg13g2_nand2b_1 _3035_ (.Y(_1485_),
    .B(net552),
    .A_N(\integrator_c_output.input_bits[1] ));
 sg13g2_o21ai_1 _3036_ (.B1(_1485_),
    .Y(_1486_),
    .A1(\integrator_c_output.bitseq[1] ),
    .A2(net552));
 sg13g2_o21ai_1 _3037_ (.B1(_1484_),
    .Y(_0441_),
    .A1(net538),
    .A2(_1486_));
 sg13g2_nor2_2 _3038_ (.A(net389),
    .B(net430),
    .Y(_1487_));
 sg13g2_nor2b_1 _3039_ (.A(_1487_),
    .B_N(\serial_input.output_case[3] ),
    .Y(_1488_));
 sg13g2_nor4_1 _3040_ (.A(\clk_counter[13] ),
    .B(\clk_counter[12] ),
    .C(\clk_counter[15] ),
    .D(\clk_counter[14] ),
    .Y(_1489_));
 sg13g2_nor4_2 _3041_ (.A(\clk_counter[9] ),
    .B(\clk_counter[8] ),
    .C(\clk_counter[11] ),
    .Y(_1490_),
    .D(\clk_counter[10] ));
 sg13g2_nor4_1 _3042_ (.A(\clk_counter[5] ),
    .B(\clk_counter[4] ),
    .C(\clk_counter[7] ),
    .D(\clk_counter[6] ),
    .Y(_1491_));
 sg13g2_nand4_1 _3043_ (.B(_1489_),
    .C(_1490_),
    .A(net578),
    .Y(_1492_),
    .D(_1491_));
 sg13g2_inv_1 _3044_ (.Y(_1493_),
    .A(_1492_));
 sg13g2_nor3_1 _3045_ (.A(\clk_counter[16] ),
    .B(\clk_counter[17] ),
    .C(_1488_),
    .Y(_1494_));
 sg13g2_nand3_1 _3046_ (.B(_1493_),
    .C(_1494_),
    .A(_0052_),
    .Y(_1495_));
 sg13g2_and2_1 _3047_ (.A(net389),
    .B(net505),
    .X(_1496_));
 sg13g2_o21ai_1 _3048_ (.B1(\serial_input.output_case[0] ),
    .Y(_1497_),
    .A1(_1487_),
    .A2(_1496_));
 sg13g2_and2_1 _3049_ (.A(\serial_input.output_case[3] ),
    .B(\serial_input.output_case[2] ),
    .X(_1498_));
 sg13g2_nor2_1 _3050_ (.A(\serial_input.output_case[3] ),
    .B(\serial_input.output_case[2] ),
    .Y(_1499_));
 sg13g2_nor3_1 _3051_ (.A(\serial_input.output_case[1] ),
    .B(_1498_),
    .C(_1499_),
    .Y(_1500_));
 sg13g2_nand2b_1 _3052_ (.Y(_1501_),
    .B(_1500_),
    .A_N(\serial_input.output_case[0] ));
 sg13g2_o21ai_1 _3053_ (.B1(_1501_),
    .Y(_1502_),
    .A1(\serial_input.output_case[3] ),
    .A2(_1497_));
 sg13g2_nor2b_1 _3054_ (.A(_1495_),
    .B_N(_1502_),
    .Y(_1503_));
 sg13g2_a21o_1 _3055_ (.A2(_1495_),
    .A1(net376),
    .B1(_1503_),
    .X(_0440_));
 sg13g2_a21o_1 _3056_ (.A2(_1495_),
    .A1(net141),
    .B1(_1503_),
    .X(_0439_));
 sg13g2_nor2b_1 _3057_ (.A(\serial_input.output_case[0] ),
    .B_N(\serial_input.output_case[1] ),
    .Y(_1504_));
 sg13g2_a221oi_1 _3058_ (.B2(_1499_),
    .C1(_1495_),
    .B1(_1504_),
    .A1(\serial_input.output_case[0] ),
    .Y(_1505_),
    .A2(_1500_));
 sg13g2_a21oi_1 _3059_ (.A1(_1651_),
    .A2(_1495_),
    .Y(_0438_),
    .B1(_1505_));
 sg13g2_nor2_1 _3060_ (.A(\serial_input.output_case[0] ),
    .B(_1496_),
    .Y(_1506_));
 sg13g2_nor4_1 _3061_ (.A(\serial_input.output_case[3] ),
    .B(_1487_),
    .C(_1495_),
    .D(_1506_),
    .Y(_1507_));
 sg13g2_a21o_1 _3062_ (.A2(_1495_),
    .A1(net380),
    .B1(_1507_),
    .X(_0437_));
 sg13g2_mux2_1 _3063_ (.A0(\serial_input.output_case[0] ),
    .A1(net227),
    .S(_1495_),
    .X(_0436_));
 sg13g2_nand2_1 _3064_ (.Y(_1508_),
    .A(net363),
    .B(net364));
 sg13g2_nor3_2 _3065_ (.A(\integrator_a_output.counter[1] ),
    .B(\integrator_a_output.counter[2] ),
    .C(_1508_),
    .Y(_1509_));
 sg13g2_nor4_2 _3066_ (.A(\integrator_a_output.counter[0] ),
    .B(\integrator_a_output.counter[1] ),
    .C(\integrator_a_output.counter[2] ),
    .Y(_1510_),
    .D(\integrator_a_output.counter[3] ));
 sg13g2_a22oi_1 _3067_ (.Y(_1511_),
    .B1(_1510_),
    .B2(net54),
    .A2(net537),
    .A1(\integrator_a_output.bitseq[7] ));
 sg13g2_inv_1 _3068_ (.Y(_0435_),
    .A(net55));
 sg13g2_nand2_1 _3069_ (.Y(_1512_),
    .A(net186),
    .B(_1509_));
 sg13g2_nand2b_1 _3070_ (.Y(_1513_),
    .B(net550),
    .A_N(\integrator_a_output.input_bits[7] ));
 sg13g2_o21ai_1 _3071_ (.B1(_1513_),
    .Y(_1514_),
    .A1(\integrator_a_output.bitseq[7] ),
    .A2(net550));
 sg13g2_o21ai_1 _3072_ (.B1(net187),
    .Y(_0434_),
    .A1(_1509_),
    .A2(_1514_));
 sg13g2_nand2_1 _3073_ (.Y(_1515_),
    .A(net91),
    .B(net537));
 sg13g2_nand2b_1 _3074_ (.Y(_1516_),
    .B(net551),
    .A_N(\integrator_a_output.input_bits[6] ));
 sg13g2_o21ai_1 _3075_ (.B1(_1516_),
    .Y(_1517_),
    .A1(\integrator_a_output.bitseq[6] ),
    .A2(net551));
 sg13g2_o21ai_1 _3076_ (.B1(_1515_),
    .Y(_0433_),
    .A1(net536),
    .A2(_1517_));
 sg13g2_nand2_1 _3077_ (.Y(_1518_),
    .A(net135),
    .B(net536));
 sg13g2_nand2b_1 _3078_ (.Y(_1519_),
    .B(net551),
    .A_N(\integrator_a_output.input_bits[5] ));
 sg13g2_o21ai_1 _3079_ (.B1(_1519_),
    .Y(_1520_),
    .A1(net91),
    .A2(net551));
 sg13g2_o21ai_1 _3080_ (.B1(_1518_),
    .Y(_0432_),
    .A1(net536),
    .A2(_1520_));
 sg13g2_nand2_1 _3081_ (.Y(_1521_),
    .A(net171),
    .B(net536));
 sg13g2_nand2b_1 _3082_ (.Y(_1522_),
    .B(net551),
    .A_N(net156));
 sg13g2_o21ai_1 _3083_ (.B1(_1522_),
    .Y(_1523_),
    .A1(net135),
    .A2(net551));
 sg13g2_o21ai_1 _3084_ (.B1(_1521_),
    .Y(_0431_),
    .A1(net536),
    .A2(_1523_));
 sg13g2_nand2_1 _3085_ (.Y(_1524_),
    .A(net225),
    .B(net536));
 sg13g2_nand2b_1 _3086_ (.Y(_1525_),
    .B(net551),
    .A_N(\integrator_a_output.input_bits[3] ));
 sg13g2_o21ai_1 _3087_ (.B1(_1525_),
    .Y(_1526_),
    .A1(net171),
    .A2(net551));
 sg13g2_o21ai_1 _3088_ (.B1(_1524_),
    .Y(_0430_),
    .A1(net536),
    .A2(_1526_));
 sg13g2_nand2_1 _3089_ (.Y(_1527_),
    .A(net110),
    .B(net537));
 sg13g2_nand2b_1 _3090_ (.Y(_1528_),
    .B(net550),
    .A_N(\integrator_a_output.input_bits[2] ));
 sg13g2_o21ai_1 _3091_ (.B1(_1528_),
    .Y(_1529_),
    .A1(\integrator_a_output.bitseq[2] ),
    .A2(net550));
 sg13g2_o21ai_1 _3092_ (.B1(_1527_),
    .Y(_0429_),
    .A1(net537),
    .A2(_1529_));
 sg13g2_nand2_1 _3093_ (.Y(_1530_),
    .A(net98),
    .B(net537));
 sg13g2_nand2b_1 _3094_ (.Y(_1531_),
    .B(net550),
    .A_N(\integrator_a_output.input_bits[1] ));
 sg13g2_o21ai_1 _3095_ (.B1(_1531_),
    .Y(_1532_),
    .A1(\integrator_a_output.bitseq[1] ),
    .A2(net550));
 sg13g2_o21ai_1 _3096_ (.B1(_1530_),
    .Y(_0428_),
    .A1(net537),
    .A2(_1532_));
 sg13g2_xnor2_1 _3097_ (.Y(_0109_),
    .A(net441),
    .B(net84));
 sg13g2_nor3_2 _3098_ (.A(net499),
    .B(_0646_),
    .C(_1492_),
    .Y(_1533_));
 sg13g2_and3_2 _3099_ (.X(_1534_),
    .A(\serial_input.output_case[0] ),
    .B(net585),
    .C(_1533_));
 sg13g2_nand2_1 _3100_ (.Y(_1535_),
    .A(_1487_),
    .B(_1534_));
 sg13g2_a22oi_1 _3101_ (.Y(_1536_),
    .B1(_1535_),
    .B2(net428),
    .A2(_1534_),
    .A1(_1496_));
 sg13g2_nand3_1 _3102_ (.B(_1498_),
    .C(_1534_),
    .A(\serial_input.output_case[1] ),
    .Y(_1537_));
 sg13g2_nor2b_1 _3103_ (.A(_1536_),
    .B_N(_1537_),
    .Y(_0427_));
 sg13g2_a21oi_1 _3104_ (.A1(\serial_input.output_case[1] ),
    .A2(_1534_),
    .Y(_1538_),
    .B1(net389));
 sg13g2_a21oi_1 _3105_ (.A1(_1496_),
    .A2(_1534_),
    .Y(_0426_),
    .B1(net390));
 sg13g2_xnor2_1 _3106_ (.Y(_1539_),
    .A(net430),
    .B(_1534_));
 sg13g2_a21oi_1 _3107_ (.A1(net428),
    .A2(_1487_),
    .Y(_0425_),
    .B1(_1539_));
 sg13g2_a21oi_1 _3108_ (.A1(net585),
    .A2(_1533_),
    .Y(_1540_),
    .B1(net413));
 sg13g2_nor2_1 _3109_ (.A(_1534_),
    .B(net414),
    .Y(_0424_));
 sg13g2_mux2_1 _3110_ (.A0(net1),
    .A1(net404),
    .S(net585),
    .X(_0423_));
 sg13g2_mux2_1 _3111_ (.A0(\serial_input.output_bitcounter_1[8] ),
    .A1(net310),
    .S(net583),
    .X(_0422_));
 sg13g2_mux2_1 _3112_ (.A0(net310),
    .A1(net290),
    .S(net583),
    .X(_0421_));
 sg13g2_mux2_1 _3113_ (.A0(net290),
    .A1(\serial_input.output_bitcounter_1[5] ),
    .S(net583),
    .X(_0420_));
 sg13g2_mux2_1 _3114_ (.A0(net333),
    .A1(net211),
    .S(net583),
    .X(_0419_));
 sg13g2_mux2_1 _3115_ (.A0(net211),
    .A1(\serial_input.output_bitcounter_1[3] ),
    .S(net583),
    .X(_0418_));
 sg13g2_mux2_1 _3116_ (.A0(net332),
    .A1(net300),
    .S(net583),
    .X(_0417_));
 sg13g2_mux2_1 _3117_ (.A0(net300),
    .A1(net120),
    .S(net583),
    .X(_0416_));
 sg13g2_mux2_1 _3118_ (.A0(net120),
    .A1(net59),
    .S(net583),
    .X(_0415_));
 sg13g2_mux2_1 _3119_ (.A0(net2),
    .A1(net336),
    .S(net585),
    .X(_0414_));
 sg13g2_mux2_1 _3120_ (.A0(net336),
    .A1(net327),
    .S(net584),
    .X(_0413_));
 sg13g2_mux2_1 _3121_ (.A0(net327),
    .A1(\serial_input.output_bitcounter_2[6] ),
    .S(net584),
    .X(_0412_));
 sg13g2_mux2_1 _3122_ (.A0(net348),
    .A1(net358),
    .S(net584),
    .X(_0411_));
 sg13g2_mux2_1 _3123_ (.A0(net358),
    .A1(net313),
    .S(net584),
    .X(_0410_));
 sg13g2_mux2_1 _3124_ (.A0(net313),
    .A1(net360),
    .S(net585),
    .X(_0409_));
 sg13g2_mux2_1 _3125_ (.A0(net360),
    .A1(net258),
    .S(net585),
    .X(_0408_));
 sg13g2_mux2_1 _3126_ (.A0(net258),
    .A1(net284),
    .S(net586),
    .X(_0407_));
 sg13g2_mux2_1 _3127_ (.A0(net284),
    .A1(net268),
    .S(net586),
    .X(_0406_));
 sg13g2_o21ai_1 _3128_ (.B1(net535),
    .Y(_0012_),
    .A1(_1654_),
    .A2(_1533_));
 sg13g2_xnor2_1 _3129_ (.Y(_1541_),
    .A(net363),
    .B(net447));
 sg13g2_nor2_1 _3130_ (.A(net536),
    .B(_1541_),
    .Y(_0001_));
 sg13g2_nand3_1 _3131_ (.B(net447),
    .C(net484),
    .A(net363),
    .Y(_1542_));
 sg13g2_a21o_1 _3132_ (.A2(net447),
    .A1(net363),
    .B1(net484),
    .X(_1543_));
 sg13g2_and2_1 _3133_ (.A(_1542_),
    .B(_1543_),
    .X(_0002_));
 sg13g2_nor2_1 _3134_ (.A(_1508_),
    .B(_0002_),
    .Y(_1544_));
 sg13g2_a21oi_1 _3135_ (.A1(_0648_),
    .A2(_1542_),
    .Y(_0003_),
    .B1(_1544_));
 sg13g2_xnor2_1 _3136_ (.Y(_1545_),
    .A(net383),
    .B(net425));
 sg13g2_nor2_1 _3137_ (.A(net549),
    .B(_1545_),
    .Y(_0005_));
 sg13g2_nand3_1 _3138_ (.B(net425),
    .C(net493),
    .A(net383),
    .Y(_1546_));
 sg13g2_a21o_1 _3139_ (.A2(net425),
    .A1(net383),
    .B1(net493),
    .X(_1547_));
 sg13g2_and2_1 _3140_ (.A(_1546_),
    .B(_1547_),
    .X(_0006_));
 sg13g2_nor2_1 _3141_ (.A(_0672_),
    .B(_0006_),
    .Y(_1548_));
 sg13g2_a21oi_1 _3142_ (.A1(_0649_),
    .A2(_1546_),
    .Y(_0007_),
    .B1(_1548_));
 sg13g2_xnor2_1 _3143_ (.Y(_1549_),
    .A(net382),
    .B(net444));
 sg13g2_nor2_1 _3144_ (.A(net539),
    .B(_1549_),
    .Y(_0009_));
 sg13g2_nand3_1 _3145_ (.B(net444),
    .C(net481),
    .A(net382),
    .Y(_1550_));
 sg13g2_a21o_1 _3146_ (.A2(net444),
    .A1(net382),
    .B1(net481),
    .X(_1551_));
 sg13g2_and2_1 _3147_ (.A(_1550_),
    .B(_1551_),
    .X(_0010_));
 sg13g2_nor2_1 _3148_ (.A(_1462_),
    .B(_0010_),
    .Y(_1552_));
 sg13g2_a21oi_1 _3149_ (.A1(_0650_),
    .A2(_1550_),
    .Y(_0011_),
    .B1(_1552_));
 sg13g2_xnor2_1 _3150_ (.Y(_1553_),
    .A(net352),
    .B(net452));
 sg13g2_nor2_1 _3151_ (.A(net542),
    .B(_1553_),
    .Y(_0014_));
 sg13g2_nand3_1 _3152_ (.B(net452),
    .C(net487),
    .A(net352),
    .Y(_1554_));
 sg13g2_a21o_1 _3153_ (.A2(net452),
    .A1(net352),
    .B1(net487),
    .X(_1555_));
 sg13g2_and2_1 _3154_ (.A(_1554_),
    .B(_1555_),
    .X(_0015_));
 sg13g2_nor2_1 _3155_ (.A(_1370_),
    .B(_0015_),
    .Y(_1556_));
 sg13g2_a21oi_1 _3156_ (.A1(_0651_),
    .A2(_1554_),
    .Y(_0016_),
    .B1(_1556_));
 sg13g2_xnor2_1 _3157_ (.Y(_1557_),
    .A(net347),
    .B(net450));
 sg13g2_nor2_1 _3158_ (.A(net544),
    .B(_1557_),
    .Y(_0018_));
 sg13g2_nand3_1 _3159_ (.B(net450),
    .C(net485),
    .A(net347),
    .Y(_1558_));
 sg13g2_a21o_1 _3160_ (.A2(net450),
    .A1(net347),
    .B1(net485),
    .X(_1559_));
 sg13g2_and2_1 _3161_ (.A(_1558_),
    .B(_1559_),
    .X(_0019_));
 sg13g2_nor2_1 _3162_ (.A(_1318_),
    .B(_0019_),
    .Y(_1560_));
 sg13g2_a21oi_1 _3163_ (.A1(_0652_),
    .A2(_1558_),
    .Y(_0020_),
    .B1(_1560_));
 sg13g2_xnor2_1 _3164_ (.Y(_1561_),
    .A(net355),
    .B(net455));
 sg13g2_nor2_1 _3165_ (.A(net546),
    .B(_1561_),
    .Y(_0022_));
 sg13g2_nand3_1 _3166_ (.B(net455),
    .C(net492),
    .A(net355),
    .Y(_1562_));
 sg13g2_a21o_1 _3167_ (.A2(net455),
    .A1(net355),
    .B1(net492),
    .X(_1563_));
 sg13g2_and2_1 _3168_ (.A(_1562_),
    .B(_1563_),
    .X(_0023_));
 sg13g2_nor2_1 _3169_ (.A(_0730_),
    .B(_0023_),
    .Y(_1564_));
 sg13g2_a21oi_1 _3170_ (.A1(_0654_),
    .A2(_1562_),
    .Y(_0024_),
    .B1(_1564_));
 sg13g2_xnor2_1 _3171_ (.Y(_1565_),
    .A(net394),
    .B(net454));
 sg13g2_nor2_1 _3172_ (.A(net540),
    .B(_1565_),
    .Y(_0026_));
 sg13g2_nand3_1 _3173_ (.B(net454),
    .C(net494),
    .A(net394),
    .Y(_1566_));
 sg13g2_a21o_1 _3174_ (.A2(net454),
    .A1(net394),
    .B1(net494),
    .X(_1567_));
 sg13g2_and2_1 _3175_ (.A(_1566_),
    .B(_1567_),
    .X(_0027_));
 sg13g2_nor2_1 _3176_ (.A(_1395_),
    .B(_0027_),
    .Y(_1568_));
 sg13g2_a21oi_1 _3177_ (.A1(_0655_),
    .A2(_1566_),
    .Y(_0028_),
    .B1(_1568_));
 sg13g2_nand2_1 _3178_ (.Y(_1569_),
    .A(net341),
    .B(net550));
 sg13g2_nand2b_1 _3179_ (.Y(_1570_),
    .B(net98),
    .A_N(net550));
 sg13g2_o21ai_1 _3180_ (.B1(_1569_),
    .Y(_1929_),
    .A1(net537),
    .A2(_1570_));
 sg13g2_nand2_1 _3181_ (.Y(_1571_),
    .A(net219),
    .B(net579));
 sg13g2_nand2b_1 _3182_ (.Y(_1572_),
    .B(net176),
    .A_N(net579));
 sg13g2_o21ai_1 _3183_ (.B1(_1571_),
    .Y(_1930_),
    .A1(net548),
    .A2(_1572_));
 sg13g2_nand2_1 _3184_ (.Y(_1573_),
    .A(net172),
    .B(net552));
 sg13g2_nand2b_1 _3185_ (.Y(_1574_),
    .B(net65),
    .A_N(_1464_));
 sg13g2_o21ai_1 _3186_ (.B1(_1573_),
    .Y(_1931_),
    .A1(net539),
    .A2(_1574_));
 sg13g2_nand2_1 _3187_ (.Y(_1575_),
    .A(net239),
    .B(net557));
 sg13g2_nand2b_1 _3188_ (.Y(_1576_),
    .B(net77),
    .A_N(net557));
 sg13g2_o21ai_1 _3189_ (.B1(_1575_),
    .Y(_1932_),
    .A1(_1371_),
    .A2(_1576_));
 sg13g2_nand2_1 _3190_ (.Y(_1577_),
    .A(net286),
    .B(net559));
 sg13g2_nand2b_1 _3191_ (.Y(_1578_),
    .B(net104),
    .A_N(net559));
 sg13g2_o21ai_1 _3192_ (.B1(_1577_),
    .Y(_1933_),
    .A1(net545),
    .A2(_1578_));
 sg13g2_nand2_1 _3193_ (.Y(_1579_),
    .A(net49),
    .B(net561));
 sg13g2_nand2b_1 _3194_ (.Y(_1580_),
    .B(\test_integrator_a_output.bitseq[0] ),
    .A_N(net561));
 sg13g2_o21ai_1 _3195_ (.B1(net50),
    .Y(_1934_),
    .A1(net547),
    .A2(_1580_));
 sg13g2_nand2_1 _3196_ (.Y(_1581_),
    .A(net174),
    .B(net555));
 sg13g2_nand2b_1 _3197_ (.Y(_1582_),
    .B(net124),
    .A_N(net555));
 sg13g2_o21ai_1 _3198_ (.B1(_1581_),
    .Y(_1935_),
    .A1(net541),
    .A2(_1582_));
 sg13g2_nand2_1 _3199_ (.Y(_1583_),
    .A(\integrator_c_counter.value_output[6] ),
    .B(_0641_));
 sg13g2_nand2_1 _3200_ (.Y(_1584_),
    .A(\integrator_c_counter.value_output[1] ),
    .B(_0634_));
 sg13g2_o21ai_1 _3201_ (.B1(_1584_),
    .Y(_1585_),
    .A1(_1640_),
    .A2(\integrator_c_sng_comparator.bits_b[0] ));
 sg13g2_a22oi_1 _3202_ (.Y(_1586_),
    .B1(\integrator_b_sng_comparator.bits_b[6] ),
    .B2(_1639_),
    .A2(net596),
    .A1(_1638_));
 sg13g2_nand2b_1 _3203_ (.Y(_1587_),
    .B(\integrator_c_counter.value_output[2] ),
    .A_N(net596));
 sg13g2_o21ai_1 _3204_ (.B1(_1587_),
    .Y(_1588_),
    .A1(_1637_),
    .A2(\integrator_c_sng_comparator.bits_b[3] ));
 sg13g2_a21oi_1 _3205_ (.A1(_1585_),
    .A2(_1586_),
    .Y(_1589_),
    .B1(_1588_));
 sg13g2_a221oi_1 _3206_ (.B2(_1637_),
    .C1(_1589_),
    .B1(\integrator_c_sng_comparator.bits_b[3] ),
    .A1(_1636_),
    .Y(_1590_),
    .A2(\input_halfprob2_sng_comparator.bits_b[6] ));
 sg13g2_nand2b_1 _3207_ (.Y(_1591_),
    .B(\integrator_c_counter.value_output[5] ),
    .A_N(\input_halfprob2_sng_comparator.bits_b[7] ));
 sg13g2_o21ai_1 _3208_ (.B1(_1591_),
    .Y(_1592_),
    .A1(_1636_),
    .A2(\input_halfprob2_sng_comparator.bits_b[6] ));
 sg13g2_a22oi_1 _3209_ (.Y(_1593_),
    .B1(\input_halfprob2_sng_comparator.bits_b[7] ),
    .B2(_1635_),
    .A2(net595),
    .A1(_1634_));
 sg13g2_o21ai_1 _3210_ (.B1(_1593_),
    .Y(_1594_),
    .A1(_1590_),
    .A2(_1592_));
 sg13g2_a22oi_1 _3211_ (.Y(_1595_),
    .B1(_1583_),
    .B2(_1594_),
    .A2(\integrator_a_sng_comparator.bits_b[1] ),
    .A1(_1633_));
 sg13g2_a221oi_1 _3212_ (.B2(\integrator_c_counter.value_output[7] ),
    .C1(_1595_),
    .B1(_0640_),
    .A1(\integrator_c_counter.value_output[8] ),
    .Y(_1596_),
    .A2(_0639_));
 sg13g2_a21oi_1 _3213_ (.A1(_1632_),
    .A2(\input_halfprob1_sng_comparator.bits_b[0] ),
    .Y(integrator_c_sn_bit),
    .B1(_1596_));
 sg13g2_xor2_1 _3214_ (.B(\clk_counter[0] ),
    .A(net423),
    .X(_0063_));
 sg13g2_nand3_1 _3215_ (.B(\clk_counter[0] ),
    .C(net475),
    .A(\clk_counter[1] ),
    .Y(_1597_));
 sg13g2_a21o_1 _3216_ (.A2(\clk_counter[0] ),
    .A1(net423),
    .B1(net475),
    .X(_1598_));
 sg13g2_and2_1 _3217_ (.A(_1597_),
    .B(net476),
    .X(_0064_));
 sg13g2_nor2_2 _3218_ (.A(_0642_),
    .B(_1597_),
    .Y(_1599_));
 sg13g2_xnor2_1 _3219_ (.Y(_0065_),
    .A(net421),
    .B(_1597_));
 sg13g2_xnor2_1 _3220_ (.Y(_0066_),
    .A(_0643_),
    .B(_1599_));
 sg13g2_nand3_1 _3221_ (.B(net468),
    .C(_1599_),
    .A(net469),
    .Y(_1600_));
 sg13g2_a21o_1 _3222_ (.A2(_1599_),
    .A1(net468),
    .B1(net469),
    .X(_1601_));
 sg13g2_and2_1 _3223_ (.A(_1600_),
    .B(_1601_),
    .X(_0067_));
 sg13g2_nand4_1 _3224_ (.B(\clk_counter[4] ),
    .C(net301),
    .A(\clk_counter[5] ),
    .Y(_1602_),
    .D(_1599_));
 sg13g2_xnor2_1 _3225_ (.Y(_0068_),
    .A(net301),
    .B(_1600_));
 sg13g2_nor2_2 _3226_ (.A(_0644_),
    .B(_1602_),
    .Y(_1603_));
 sg13g2_xnor2_1 _3227_ (.Y(_0069_),
    .A(net253),
    .B(_1602_));
 sg13g2_xor2_1 _3228_ (.B(_1603_),
    .A(net378),
    .X(_0070_));
 sg13g2_nand3_1 _3229_ (.B(net378),
    .C(_1603_),
    .A(net458),
    .Y(_1604_));
 sg13g2_a21o_1 _3230_ (.A2(_1603_),
    .A1(net378),
    .B1(net458),
    .X(_1605_));
 sg13g2_and2_1 _3231_ (.A(_1604_),
    .B(_1605_),
    .X(_0071_));
 sg13g2_nor2_1 _3232_ (.A(_0645_),
    .B(_1604_),
    .Y(_1606_));
 sg13g2_xnor2_1 _3233_ (.Y(_0055_),
    .A(net368),
    .B(_1604_));
 sg13g2_and2_1 _3234_ (.A(net270),
    .B(_1606_),
    .X(_1607_));
 sg13g2_xor2_1 _3235_ (.B(_1606_),
    .A(net270),
    .X(_0056_));
 sg13g2_xor2_1 _3236_ (.B(_1607_),
    .A(net371),
    .X(_0057_));
 sg13g2_and3_2 _3237_ (.X(_1608_),
    .A(net95),
    .B(net371),
    .C(_1607_));
 sg13g2_a21oi_1 _3238_ (.A1(\clk_counter[12] ),
    .A2(_1607_),
    .Y(_1609_),
    .B1(net95));
 sg13g2_nor2_1 _3239_ (.A(_1608_),
    .B(net96),
    .Y(_0058_));
 sg13g2_xor2_1 _3240_ (.B(_1608_),
    .A(net406),
    .X(_0059_));
 sg13g2_nand3_1 _3241_ (.B(net406),
    .C(_1608_),
    .A(net426),
    .Y(_1610_));
 sg13g2_a21o_1 _3242_ (.A2(_1608_),
    .A1(net406),
    .B1(net426),
    .X(_1611_));
 sg13g2_and2_1 _3243_ (.A(_1610_),
    .B(_1611_),
    .X(_0060_));
 sg13g2_nand4_1 _3244_ (.B(\clk_counter[14] ),
    .C(\clk_counter[16] ),
    .A(\clk_counter[15] ),
    .Y(_1612_),
    .D(_1608_));
 sg13g2_xnor2_1 _3245_ (.Y(_0061_),
    .A(\clk_counter[16] ),
    .B(_1610_));
 sg13g2_xnor2_1 _3246_ (.Y(_0062_),
    .A(net306),
    .B(_1612_));
 sg13g2_inv_1 _3247_ (.Y(_0088_),
    .A(net651));
 sg13g2_inv_1 _3248_ (.Y(_0089_),
    .A(net654));
 sg13g2_inv_1 _3249_ (.Y(_0090_),
    .A(net654));
 sg13g2_inv_1 _3250_ (.Y(_0091_),
    .A(net648));
 sg13g2_inv_1 _3251_ (.Y(_0092_),
    .A(net648));
 sg13g2_inv_1 _3252_ (.Y(_0093_),
    .A(net648));
 sg13g2_inv_1 _3253_ (.Y(_0094_),
    .A(net648));
 sg13g2_inv_1 _3254_ (.Y(_0095_),
    .A(net655));
 sg13g2_inv_1 _3255_ (.Y(_0096_),
    .A(net646));
 sg13g2_inv_1 _3256_ (.Y(_0097_),
    .A(net646));
 sg13g2_inv_1 _3257_ (.Y(_0098_),
    .A(net646));
 sg13g2_inv_1 _3258_ (.Y(_0099_),
    .A(net646));
 sg13g2_inv_1 _3259_ (.Y(_0100_),
    .A(net649));
 sg13g2_inv_1 _3260_ (.Y(_0101_),
    .A(net646));
 sg13g2_inv_1 _3261_ (.Y(_0102_),
    .A(net646));
 sg13g2_inv_1 _3262_ (.Y(_0103_),
    .A(net646));
 sg13g2_inv_1 _3263_ (.Y(_0104_),
    .A(net655));
 sg13g2_inv_1 _3264_ (.Y(_0105_),
    .A(net654));
 sg13g2_inv_1 _3265_ (.Y(_0106_),
    .A(net654));
 sg13g2_inv_1 _3266_ (.Y(_0107_),
    .A(net654));
 sg13g2_inv_1 _3267_ (.Y(_0108_),
    .A(net654));
 sg13g2_inv_1 _3268_ (.Y(_0110_),
    .A(net632));
 sg13g2_inv_1 _3269_ (.Y(_0112_),
    .A(net645));
 sg13g2_inv_1 _3270_ (.Y(_0113_),
    .A(net642));
 sg13g2_inv_1 _3271_ (.Y(_0114_),
    .A(net642));
 sg13g2_inv_1 _3272_ (.Y(_0115_),
    .A(net642));
 sg13g2_inv_1 _3273_ (.Y(_0116_),
    .A(net622));
 sg13g2_inv_1 _3274_ (.Y(_0117_),
    .A(net626));
 sg13g2_inv_1 _3275_ (.Y(_0118_),
    .A(net622));
 sg13g2_inv_1 _3276_ (.Y(_0119_),
    .A(net626));
 sg13g2_inv_1 _3277_ (.Y(_0121_),
    .A(net622));
 sg13g2_inv_1 _3278_ (.Y(_0123_),
    .A(net642));
 sg13g2_inv_1 _3279_ (.Y(_0125_),
    .A(net632));
 sg13g2_inv_1 _3280_ (.Y(_0126_),
    .A(net642));
 sg13g2_inv_1 _3281_ (.Y(_0127_),
    .A(net642));
 sg13g2_inv_1 _3282_ (.Y(_0128_),
    .A(net642));
 sg13g2_inv_1 _3283_ (.Y(_0129_),
    .A(net645));
 sg13g2_inv_1 _3284_ (.Y(_0130_),
    .A(net644));
 sg13g2_inv_1 _3285_ (.Y(_0131_),
    .A(net644));
 sg13g2_inv_1 _3286_ (.Y(_0132_),
    .A(net644));
 sg13g2_inv_1 _3287_ (.Y(_0133_),
    .A(net643));
 sg13g2_inv_1 _3288_ (.Y(_0134_),
    .A(net643));
 sg13g2_inv_1 _3289_ (.Y(_0135_),
    .A(net631));
 sg13g2_inv_1 _3290_ (.Y(_0136_),
    .A(net632));
 sg13g2_inv_1 _3291_ (.Y(_0137_),
    .A(net613));
 sg13g2_inv_1 _3292_ (.Y(_0138_),
    .A(net632));
 sg13g2_inv_1 _3293_ (.Y(_0139_),
    .A(net632));
 sg13g2_inv_1 _3294_ (.Y(_0140_),
    .A(net632));
 sg13g2_inv_1 _3295_ (.Y(_0141_),
    .A(net632));
 sg13g2_inv_1 _3296_ (.Y(_0142_),
    .A(net630));
 sg13g2_inv_1 _3297_ (.Y(_0143_),
    .A(net611));
 sg13g2_inv_1 _3298_ (.Y(_0144_),
    .A(net613));
 sg13g2_inv_1 _3299_ (.Y(_0145_),
    .A(net610));
 sg13g2_inv_1 _3300_ (.Y(_0146_),
    .A(net610));
 sg13g2_inv_1 _3301_ (.Y(_0147_),
    .A(net610));
 sg13g2_inv_1 _3302_ (.Y(_0148_),
    .A(net604));
 sg13g2_inv_1 _3303_ (.Y(_0149_),
    .A(net604));
 sg13g2_inv_1 _3304_ (.Y(_0150_),
    .A(net604));
 sg13g2_inv_1 _3305_ (.Y(_0151_),
    .A(net610));
 sg13g2_inv_1 _3306_ (.Y(_0152_),
    .A(net610));
 sg13g2_inv_1 _3307_ (.Y(_0153_),
    .A(net655));
 sg13g2_inv_1 _3308_ (.Y(_0154_),
    .A(net655));
 sg13g2_inv_1 _3309_ (.Y(_0155_),
    .A(net656));
 sg13g2_inv_1 _3310_ (.Y(_0156_),
    .A(net655));
 sg13g2_inv_1 _3311_ (.Y(_0157_),
    .A(net656));
 sg13g2_inv_1 _3312_ (.Y(_0159_),
    .A(net604));
 sg13g2_inv_1 _3313_ (.Y(_0160_),
    .A(net651));
 sg13g2_inv_1 _3314_ (.Y(_0161_),
    .A(net652));
 sg13g2_inv_1 _3315_ (.Y(_0162_),
    .A(net652));
 sg13g2_inv_1 _3316_ (.Y(_0163_),
    .A(net651));
 sg13g2_inv_1 _3317_ (.Y(_0164_),
    .A(net651));
 sg13g2_inv_1 _3318_ (.Y(_0165_),
    .A(net651));
 sg13g2_inv_1 _3319_ (.Y(_0166_),
    .A(net651));
 sg13g2_inv_1 _3320_ (.Y(_0167_),
    .A(net638));
 sg13g2_inv_1 _3321_ (.Y(_0168_),
    .A(net617));
 sg13g2_inv_1 _3322_ (.Y(_0169_),
    .A(net617));
 sg13g2_inv_1 _3323_ (.Y(_0170_),
    .A(net622));
 sg13g2_inv_1 _3324_ (.Y(_0171_),
    .A(net622));
 sg13g2_inv_1 _3325_ (.Y(_0172_),
    .A(net617));
 sg13g2_inv_1 _3326_ (.Y(_0173_),
    .A(net617));
 sg13g2_inv_1 _3327_ (.Y(_0174_),
    .A(net617));
 sg13g2_inv_1 _3328_ (.Y(_0175_),
    .A(net617));
 sg13g2_inv_1 _3329_ (.Y(_0176_),
    .A(net616));
 sg13g2_inv_1 _3330_ (.Y(_0177_),
    .A(net616));
 sg13g2_inv_1 _3331_ (.Y(_0178_),
    .A(net616));
 sg13g2_inv_1 _3332_ (.Y(_0179_),
    .A(net616));
 sg13g2_inv_1 _3333_ (.Y(_0180_),
    .A(net616));
 sg13g2_inv_1 _3334_ (.Y(_0181_),
    .A(net616));
 sg13g2_inv_1 _3335_ (.Y(_0182_),
    .A(net615));
 sg13g2_inv_1 _3336_ (.Y(_0183_),
    .A(net615));
 sg13g2_inv_1 _3337_ (.Y(_0184_),
    .A(net633));
 sg13g2_inv_1 _3338_ (.Y(_0185_),
    .A(net634));
 sg13g2_inv_1 _3339_ (.Y(_0186_),
    .A(net633));
 sg13g2_inv_1 _3340_ (.Y(_0187_),
    .A(net633));
 sg13g2_inv_1 _3341_ (.Y(_0188_),
    .A(net629));
 sg13g2_inv_1 _3342_ (.Y(_0189_),
    .A(net629));
 sg13g2_inv_1 _3343_ (.Y(_0190_),
    .A(net629));
 sg13g2_inv_1 _3344_ (.Y(_0191_),
    .A(net628));
 sg13g2_inv_1 _3345_ (.Y(_0192_),
    .A(net622));
 sg13g2_inv_1 _3346_ (.Y(_0193_),
    .A(net606));
 sg13g2_inv_1 _3347_ (.Y(_0194_),
    .A(net606));
 sg13g2_inv_1 _3348_ (.Y(_0195_),
    .A(net606));
 sg13g2_inv_1 _3349_ (.Y(_0196_),
    .A(net606));
 sg13g2_inv_1 _3350_ (.Y(_0197_),
    .A(net607));
 sg13g2_inv_1 _3351_ (.Y(_0198_),
    .A(net607));
 sg13g2_inv_1 _3352_ (.Y(_0199_),
    .A(net607));
 sg13g2_inv_1 _3353_ (.Y(_0200_),
    .A(net607));
 sg13g2_inv_1 _3354_ (.Y(_0201_),
    .A(net615));
 sg13g2_inv_1 _3355_ (.Y(_0202_),
    .A(net615));
 sg13g2_inv_1 _3356_ (.Y(_0203_),
    .A(net617));
 sg13g2_inv_1 _3357_ (.Y(_0204_),
    .A(net618));
 sg13g2_inv_1 _3358_ (.Y(_0205_),
    .A(net618));
 sg13g2_inv_1 _3359_ (.Y(_0206_),
    .A(net615));
 sg13g2_inv_1 _3360_ (.Y(_0207_),
    .A(net615));
 sg13g2_inv_1 _3361_ (.Y(_0208_),
    .A(net615));
 sg13g2_inv_1 _3362_ (.Y(_0209_),
    .A(net615));
 sg13g2_inv_1 _3363_ (.Y(_0210_),
    .A(net639));
 sg13g2_inv_1 _3364_ (.Y(_0211_),
    .A(net604));
 sg13g2_inv_1 _3365_ (.Y(_0212_),
    .A(net604));
 sg13g2_inv_1 _3366_ (.Y(_0213_),
    .A(net604));
 sg13g2_inv_1 _3367_ (.Y(_0214_),
    .A(net604));
 sg13g2_inv_1 _3368_ (.Y(_0215_),
    .A(net611));
 sg13g2_inv_1 _3369_ (.Y(_0216_),
    .A(net611));
 sg13g2_inv_1 _3370_ (.Y(_0217_),
    .A(net612));
 sg13g2_inv_1 _3371_ (.Y(_0218_),
    .A(net608));
 sg13g2_inv_1 _3372_ (.Y(_0219_),
    .A(net612));
 sg13g2_inv_1 _3373_ (.Y(_0220_),
    .A(net605));
 sg13g2_inv_1 _3374_ (.Y(_0221_),
    .A(net610));
 sg13g2_inv_1 _3375_ (.Y(_0222_),
    .A(net610));
 sg13g2_inv_1 _3376_ (.Y(_0223_),
    .A(net611));
 sg13g2_inv_1 _3377_ (.Y(_0224_),
    .A(net651));
 sg13g2_inv_1 _3378_ (.Y(_0225_),
    .A(net620));
 sg13g2_inv_1 _3379_ (.Y(_0226_),
    .A(net619));
 sg13g2_inv_1 _3380_ (.Y(_0227_),
    .A(net619));
 sg13g2_inv_1 _3381_ (.Y(_0228_),
    .A(net619));
 sg13g2_inv_1 _3382_ (.Y(_0229_),
    .A(net623));
 sg13g2_inv_1 _3383_ (.Y(_0230_),
    .A(net623));
 sg13g2_inv_1 _3384_ (.Y(_0231_),
    .A(net623));
 sg13g2_inv_1 _3385_ (.Y(_0232_),
    .A(net623));
 sg13g2_inv_1 _3386_ (.Y(_0233_),
    .A(net619));
 sg13g2_inv_1 _3387_ (.Y(_0234_),
    .A(net619));
 sg13g2_inv_1 _3388_ (.Y(_0235_),
    .A(net619));
 sg13g2_inv_1 _3389_ (.Y(_0236_),
    .A(net617));
 sg13g2_inv_1 _3390_ (.Y(_0237_),
    .A(net622));
 sg13g2_inv_1 _3391_ (.Y(_0238_),
    .A(net651));
 sg13g2_inv_1 _3392_ (.Y(_0239_),
    .A(net652));
 sg13g2_inv_1 _3393_ (.Y(_0240_),
    .A(net652));
 sg13g2_inv_1 _3394_ (.Y(_0241_),
    .A(net652));
 sg13g2_inv_1 _3395_ (.Y(_0242_),
    .A(net652));
 sg13g2_inv_1 _3396_ (.Y(_0243_),
    .A(net643));
 sg13g2_inv_1 _3397_ (.Y(_0244_),
    .A(net643));
 sg13g2_inv_1 _3398_ (.Y(_0245_),
    .A(net643));
 sg13g2_inv_1 _3399_ (.Y(_0246_),
    .A(net643));
 sg13g2_inv_1 _3400_ (.Y(_0247_),
    .A(net640));
 sg13g2_inv_1 _3401_ (.Y(_0248_),
    .A(net631));
 sg13g2_inv_1 _3402_ (.Y(_0249_),
    .A(net631));
 sg13g2_inv_1 _3403_ (.Y(_0250_),
    .A(net631));
 sg13g2_inv_1 _3404_ (.Y(_0251_),
    .A(net631));
 sg13g2_inv_1 _3405_ (.Y(_0252_),
    .A(net639));
 sg13g2_inv_1 _3406_ (.Y(_0253_),
    .A(net634));
 sg13g2_inv_1 _3407_ (.Y(_0254_),
    .A(net634));
 sg13g2_inv_1 _3408_ (.Y(_0255_),
    .A(net633));
 sg13g2_inv_1 _3409_ (.Y(_0256_),
    .A(net633));
 sg13g2_inv_1 _3410_ (.Y(_0257_),
    .A(net629));
 sg13g2_inv_1 _3411_ (.Y(_0258_),
    .A(net630));
 sg13g2_inv_1 _3412_ (.Y(_0259_),
    .A(net630));
 sg13g2_inv_1 _3413_ (.Y(_0260_),
    .A(net629));
 sg13g2_inv_1 _3414_ (.Y(_0261_),
    .A(net628));
 sg13g2_inv_1 _3415_ (.Y(_0262_),
    .A(net628));
 sg13g2_inv_1 _3416_ (.Y(_0263_),
    .A(net628));
 sg13g2_inv_1 _3417_ (.Y(_0264_),
    .A(net628));
 sg13g2_inv_1 _3418_ (.Y(_0265_),
    .A(net630));
 sg13g2_inv_1 _3419_ (.Y(_0266_),
    .A(net639));
 sg13g2_inv_1 _3420_ (.Y(_0267_),
    .A(net606));
 sg13g2_inv_1 _3421_ (.Y(_0268_),
    .A(net606));
 sg13g2_inv_1 _3422_ (.Y(_0269_),
    .A(net606));
 sg13g2_inv_1 _3423_ (.Y(_0270_),
    .A(net606));
 sg13g2_inv_1 _3424_ (.Y(_0271_),
    .A(net613));
 sg13g2_inv_1 _3425_ (.Y(_0272_),
    .A(net612));
 sg13g2_inv_1 _3426_ (.Y(_0273_),
    .A(net612));
 sg13g2_inv_1 _3427_ (.Y(_0274_),
    .A(net613));
 sg13g2_inv_1 _3428_ (.Y(_0275_),
    .A(net612));
 sg13g2_inv_1 _3429_ (.Y(_0276_),
    .A(net612));
 sg13g2_inv_1 _3430_ (.Y(_0277_),
    .A(net612));
 sg13g2_inv_1 _3431_ (.Y(_0278_),
    .A(net612));
 sg13g2_inv_1 _3432_ (.Y(_0279_),
    .A(net613));
 sg13g2_inv_1 _3433_ (.Y(_0280_),
    .A(net639));
 sg13g2_inv_1 _3434_ (.Y(_0281_),
    .A(net635));
 sg13g2_inv_1 _3435_ (.Y(_0282_),
    .A(net635));
 sg13g2_inv_1 _3436_ (.Y(_0283_),
    .A(net635));
 sg13g2_inv_1 _3437_ (.Y(_0284_),
    .A(net635));
 sg13g2_inv_1 _3438_ (.Y(_0285_),
    .A(net637));
 sg13g2_inv_1 _3439_ (.Y(_0286_),
    .A(net637));
 sg13g2_inv_1 _3440_ (.Y(_0287_),
    .A(net637));
 sg13g2_inv_1 _3441_ (.Y(_0288_),
    .A(net637));
 sg13g2_inv_1 _3442_ (.Y(_0289_),
    .A(net637));
 sg13g2_inv_1 _3443_ (.Y(_0290_),
    .A(net637));
 sg13g2_inv_1 _3444_ (.Y(_0291_),
    .A(net631));
 sg13g2_inv_1 _3445_ (.Y(_0292_),
    .A(net631));
 sg13g2_inv_1 _3446_ (.Y(_0293_),
    .A(net631));
 sg13g2_inv_1 _3447_ (.Y(_0294_),
    .A(net638));
 sg13g2_inv_1 _3448_ (.Y(_0295_),
    .A(net621));
 sg13g2_inv_1 _3449_ (.Y(_0296_),
    .A(net621));
 sg13g2_inv_1 _3450_ (.Y(_0297_),
    .A(net621));
 sg13g2_inv_1 _3451_ (.Y(_0298_),
    .A(net621));
 sg13g2_inv_1 _3452_ (.Y(_0299_),
    .A(net638));
 sg13g2_inv_1 _3453_ (.Y(_0300_),
    .A(net638));
 sg13g2_inv_1 _3454_ (.Y(_0301_),
    .A(net638));
 sg13g2_inv_1 _3455_ (.Y(_0302_),
    .A(net635));
 sg13g2_inv_1 _3456_ (.Y(_0303_),
    .A(net635));
 sg13g2_inv_1 _3457_ (.Y(_0304_),
    .A(net635));
 sg13g2_inv_1 _3458_ (.Y(_0305_),
    .A(net636));
 sg13g2_inv_1 _3459_ (.Y(_0306_),
    .A(net635));
 sg13g2_inv_1 _3460_ (.Y(_0307_),
    .A(net610));
 sg13g2_inv_1 _3461_ (.Y(_0308_),
    .A(net611));
 sg13g2_inv_1 _3462_ (.Y(_0309_),
    .A(net611));
 sg13g2_inv_1 _3463_ (.Y(_0310_),
    .A(net605));
 sg13g2_inv_1 _3464_ (.Y(_0311_),
    .A(net605));
 sg13g2_inv_1 _3465_ (.Y(_0312_),
    .A(net605));
 sg13g2_inv_1 _3466_ (.Y(_0313_),
    .A(net605));
 sg13g2_inv_1 _3467_ (.Y(_0314_),
    .A(net614));
 sg13g2_inv_1 _3468_ (.Y(_0315_),
    .A(net611));
 sg13g2_inv_1 _3469_ (.Y(_0316_),
    .A(net624));
 sg13g2_inv_1 _3470_ (.Y(_0317_),
    .A(net625));
 sg13g2_inv_1 _3471_ (.Y(_0318_),
    .A(net625));
 sg13g2_inv_1 _3472_ (.Y(_0319_),
    .A(net623));
 sg13g2_inv_1 _3473_ (.Y(_0320_),
    .A(net625));
 sg13g2_inv_1 _3474_ (.Y(_0321_),
    .A(net623));
 sg13g2_inv_1 _3475_ (.Y(_0322_),
    .A(net620));
 sg13g2_inv_1 _3476_ (.Y(_0323_),
    .A(net619));
 sg13g2_inv_1 _3477_ (.Y(_0324_),
    .A(net619));
 sg13g2_inv_1 _3478_ (.Y(_0325_),
    .A(net650));
 sg13g2_inv_1 _3479_ (.Y(_0326_),
    .A(net644));
 sg13g2_inv_1 _3480_ (.Y(_0327_),
    .A(net650));
 sg13g2_inv_1 _3481_ (.Y(_0328_),
    .A(net650));
 sg13g2_inv_1 _3482_ (.Y(_0329_),
    .A(net650));
 sg13g2_inv_1 _3483_ (.Y(_0330_),
    .A(net650));
 sg13g2_inv_1 _3484_ (.Y(_0331_),
    .A(net637));
 sg13g2_inv_1 _3485_ (.Y(_0332_),
    .A(net640));
 sg13g2_inv_1 _3486_ (.Y(_0333_),
    .A(net637));
 sg13g2_inv_1 _3487_ (.Y(_0334_),
    .A(net633));
 sg13g2_inv_1 _3488_ (.Y(_0335_),
    .A(net633));
 sg13g2_inv_1 _3489_ (.Y(_0336_),
    .A(net633));
 sg13g2_inv_1 _3490_ (.Y(_0337_),
    .A(net629));
 sg13g2_inv_1 _3491_ (.Y(_0338_),
    .A(net629));
 sg13g2_inv_1 _3492_ (.Y(_0339_),
    .A(net629));
 sg13g2_inv_1 _3493_ (.Y(_0340_),
    .A(net628));
 sg13g2_inv_1 _3494_ (.Y(_0341_),
    .A(net628));
 sg13g2_inv_1 _3495_ (.Y(_0342_),
    .A(net628));
 sg13g2_inv_1 _3496_ (.Y(_0343_),
    .A(net609));
 sg13g2_inv_1 _3497_ (.Y(_0344_),
    .A(net608));
 sg13g2_inv_1 _3498_ (.Y(_0345_),
    .A(net608));
 sg13g2_inv_1 _3499_ (.Y(_0346_),
    .A(net608));
 sg13g2_inv_1 _3500_ (.Y(_0347_),
    .A(net608));
 sg13g2_inv_1 _3501_ (.Y(_0348_),
    .A(net607));
 sg13g2_inv_1 _3502_ (.Y(_0349_),
    .A(net608));
 sg13g2_inv_1 _3503_ (.Y(_0350_),
    .A(net607));
 sg13g2_inv_1 _3504_ (.Y(_0351_),
    .A(net607));
 sg13g2_inv_1 _3505_ (.Y(_0352_),
    .A(net639));
 sg13g2_inv_1 _3506_ (.Y(_0353_),
    .A(net638));
 sg13g2_inv_1 _3507_ (.Y(_0354_),
    .A(net638));
 sg13g2_inv_1 _3508_ (.Y(_0355_),
    .A(net638));
 sg13g2_inv_1 _3509_ (.Y(_0356_),
    .A(net636));
 sg13g2_inv_1 _3510_ (.Y(_0357_),
    .A(net634));
 sg13g2_inv_1 _3511_ (.Y(_0358_),
    .A(net634));
 sg13g2_inv_1 _3512_ (.Y(_0359_),
    .A(net634));
 sg13g2_inv_1 _3513_ (.Y(_0360_),
    .A(net634));
 sg13g2_inv_1 _3514_ (.Y(_0361_),
    .A(net655));
 sg13g2_inv_1 _3515_ (.Y(_0362_),
    .A(net656));
 sg13g2_inv_1 _3516_ (.Y(_0363_),
    .A(net655));
 sg13g2_inv_1 _3517_ (.Y(_0364_),
    .A(net656));
 sg13g2_inv_1 _3518_ (.Y(_0365_),
    .A(net656));
 sg13g2_inv_1 _3519_ (.Y(_0366_),
    .A(net656));
 sg13g2_inv_1 _3520_ (.Y(_0367_),
    .A(net657));
 sg13g2_inv_1 _3521_ (.Y(_0368_),
    .A(net654));
 sg13g2_inv_1 _3522_ (.Y(_0369_),
    .A(net647));
 sg13g2_inv_1 _3523_ (.Y(_0370_),
    .A(net647));
 sg13g2_inv_1 _3524_ (.Y(_0371_),
    .A(net647));
 sg13g2_inv_1 _3525_ (.Y(_0372_),
    .A(net647));
 sg13g2_inv_1 _3526_ (.Y(_0373_),
    .A(net649));
 sg13g2_inv_1 _3527_ (.Y(_0374_),
    .A(net647));
 sg13g2_inv_1 _3528_ (.Y(_0375_),
    .A(net647));
 sg13g2_inv_1 _3529_ (.Y(_0376_),
    .A(net647));
 sg13g2_inv_1 _3530_ (.Y(_0377_),
    .A(net647));
 sg13g2_inv_1 _3531_ (.Y(_0378_),
    .A(net657));
 sg13g2_inv_1 _3532_ (.Y(_0379_),
    .A(net645));
 sg13g2_inv_1 _3533_ (.Y(_0380_),
    .A(net646));
 sg13g2_inv_1 _3534_ (.Y(_0381_),
    .A(net649));
 sg13g2_inv_1 _3535_ (.Y(_0382_),
    .A(net649));
 sg13g2_inv_1 _3536_ (.Y(_0383_),
    .A(net624));
 sg13g2_inv_1 _3537_ (.Y(_0384_),
    .A(net624));
 sg13g2_inv_1 _3538_ (.Y(_0385_),
    .A(net624));
 sg13g2_inv_1 _3539_ (.Y(_0386_),
    .A(net622));
 sg13g2_inv_1 _3540_ (.Y(_0387_),
    .A(net642));
 sg13g2_inv_1 _3541_ (.Y(_0388_),
    .A(net654));
 sg13g2_inv_1 _3542_ (.Y(_0389_),
    .A(net624));
 sg13g2_inv_1 _3543_ (.Y(_0390_),
    .A(net624));
 sg13g2_inv_1 _3544_ (.Y(_0391_),
    .A(net624));
 sg13g2_inv_1 _3545_ (.Y(_0392_),
    .A(net624));
 sg13g2_inv_1 _3546_ (.Y(_0393_),
    .A(net623));
 sg13g2_inv_1 _3547_ (.Y(_0394_),
    .A(net623));
 sg13g2_inv_1 _3548_ (.Y(_0395_),
    .A(net620));
 sg13g2_inv_1 _3549_ (.Y(_0396_),
    .A(net620));
 sg13g2_inv_1 _3550_ (.Y(_0397_),
    .A(net650));
 sg13g2_inv_1 _3551_ (.Y(_0398_),
    .A(net650));
 sg13g2_inv_1 _3552_ (.Y(_0399_),
    .A(net650));
 sg13g2_inv_1 _3553_ (.Y(_0400_),
    .A(net653));
 sg13g2_inv_1 _3554_ (.Y(_0401_),
    .A(net643));
 sg13g2_inv_1 _3555_ (.Y(_0402_),
    .A(net648));
 sg13g2_inv_1 _3556_ (.Y(_0403_),
    .A(net648));
 sg13g2_inv_1 _3557_ (.Y(_0404_),
    .A(net648));
 sg13g2_inv_1 _3558_ (.Y(_0405_),
    .A(net643));
 sg13g2_dfrbp_1 _3559_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(_0087_),
    .D(_0406_),
    .Q_N(_1928_),
    .Q(\serial_input.output_bitcounter_2[0] ));
 sg13g2_dfrbp_1 _3560_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(_0088_),
    .D(_0407_),
    .Q_N(_1927_),
    .Q(\serial_input.output_bitcounter_2[1] ));
 sg13g2_dfrbp_1 _3561_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(_0089_),
    .D(_0408_),
    .Q_N(_1926_),
    .Q(\serial_input.output_bitcounter_2[2] ));
 sg13g2_dfrbp_1 _3562_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(_0090_),
    .D(_0409_),
    .Q_N(_1925_),
    .Q(\serial_input.output_bitcounter_2[3] ));
 sg13g2_dfrbp_1 _3563_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(_0091_),
    .D(_0410_),
    .Q_N(_1924_),
    .Q(\serial_input.output_bitcounter_2[4] ));
 sg13g2_dfrbp_1 _3564_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(_0092_),
    .D(_0411_),
    .Q_N(_1923_),
    .Q(\serial_input.output_bitcounter_2[5] ));
 sg13g2_dfrbp_1 _3565_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(_0093_),
    .D(net328),
    .Q_N(_1922_),
    .Q(\serial_input.output_bitcounter_2[6] ));
 sg13g2_dfrbp_1 _3566_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(_0094_),
    .D(_0413_),
    .Q_N(_1921_),
    .Q(\serial_input.output_bitcounter_2[7] ));
 sg13g2_dfrbp_1 _3567_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(_0095_),
    .D(_0414_),
    .Q_N(_1920_),
    .Q(\serial_input.output_bitcounter_2[8] ));
 sg13g2_dfrbp_1 _3568_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(_0096_),
    .D(_0415_),
    .Q_N(_1919_),
    .Q(\serial_input.output_bitcounter_1[0] ));
 sg13g2_dfrbp_1 _3569_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(_0097_),
    .D(_0416_),
    .Q_N(_1918_),
    .Q(\serial_input.output_bitcounter_1[1] ));
 sg13g2_dfrbp_1 _3570_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(_0098_),
    .D(_0417_),
    .Q_N(_1917_),
    .Q(\serial_input.output_bitcounter_1[2] ));
 sg13g2_dfrbp_1 _3571_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(_0099_),
    .D(net212),
    .Q_N(_1916_),
    .Q(\serial_input.output_bitcounter_1[3] ));
 sg13g2_dfrbp_1 _3572_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(_0100_),
    .D(_0419_),
    .Q_N(_1915_),
    .Q(\serial_input.output_bitcounter_1[4] ));
 sg13g2_dfrbp_1 _3573_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(_0101_),
    .D(net291),
    .Q_N(_1914_),
    .Q(\serial_input.output_bitcounter_1[5] ));
 sg13g2_dfrbp_1 _3574_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(_0102_),
    .D(_0421_),
    .Q_N(_1913_),
    .Q(\serial_input.output_bitcounter_1[6] ));
 sg13g2_dfrbp_1 _3575_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(_0103_),
    .D(net311),
    .Q_N(_1912_),
    .Q(\serial_input.output_bitcounter_1[7] ));
 sg13g2_dfrbp_1 _3576_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(_0104_),
    .D(_0423_),
    .Q_N(_1911_),
    .Q(\serial_input.output_bitcounter_1[8] ));
 sg13g2_dfrbp_1 _3577_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(_0105_),
    .D(_0424_),
    .Q_N(_1910_),
    .Q(\serial_input.output_case[0] ));
 sg13g2_dfrbp_1 _3578_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(_0106_),
    .D(_0425_),
    .Q_N(_1909_),
    .Q(\serial_input.output_case[1] ));
 sg13g2_dfrbp_1 _3579_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(_0107_),
    .D(_0426_),
    .Q_N(_1908_),
    .Q(\serial_input.output_case[2] ));
 sg13g2_dfrbp_1 _3580_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(_0108_),
    .D(net429),
    .Q_N(_1907_),
    .Q(\serial_input.output_case[3] ));
 sg13g2_dfrbp_1 _3581_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(_0110_),
    .D(_0109_),
    .Q_N(\input_a_sng_comparator.bits_b[0] ),
    .Q(_0075_));
 sg13g2_dfrbp_1 _3582_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(_0112_),
    .D(_0111_),
    .Q_N(\input_a_sng_comparator.bits_b[1] ),
    .Q(_0076_));
 sg13g2_dfrbp_1 _3583_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(_0113_),
    .D(net28),
    .Q_N(_1906_),
    .Q(\input_a_sng_comparator.bits_b[2] ));
 sg13g2_dfrbp_1 _3584_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(_0114_),
    .D(net37),
    .Q_N(_1905_),
    .Q(\input_a_sng_comparator.bits_b[3] ));
 sg13g2_dfrbp_1 _3585_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(_0115_),
    .D(net22),
    .Q_N(\input_a_sng_comparator.bits_b[4] ),
    .Q(_0077_));
 sg13g2_dfrbp_1 _3586_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(_0116_),
    .D(net599),
    .Q_N(_1904_),
    .Q(\input_a_sng_comparator.bits_b[5] ));
 sg13g2_dfrbp_1 _3587_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(_0117_),
    .D(net20),
    .Q_N(\input_a_sng_comparator.bits_b[6] ),
    .Q(_0078_));
 sg13g2_dfrbp_1 _3588_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(_0118_),
    .D(net597),
    .Q_N(_1903_),
    .Q(\input_a_sng_comparator.bits_b[7] ));
 sg13g2_dfrbp_1 _3589_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(_0119_),
    .D(net21),
    .Q_N(\input_a_sng_comparator.bits_b[8] ),
    .Q(_0079_));
 sg13g2_dfrbp_1 _3590_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(_0121_),
    .D(_0120_),
    .Q_N(\input_halfprob1_sng_comparator.bits_b[6] ),
    .Q(_0080_));
 sg13g2_dfrbp_1 _3591_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(_0123_),
    .D(_0122_),
    .Q_N(\input_halfprob1_sng_comparator.bits_b[7] ),
    .Q(_0081_));
 sg13g2_dfrbp_1 _3592_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(_0125_),
    .D(_0124_),
    .Q_N(\input_halfprob1_sng_comparator.bits_b[8] ),
    .Q(_0082_));
 sg13g2_dfrbp_1 _3593_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(_0126_),
    .D(net31),
    .Q_N(_1902_),
    .Q(\integrator_c_sng_comparator.bits_b[0] ));
 sg13g2_dfrbp_1 _3594_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(_0127_),
    .D(net32),
    .Q_N(_1901_),
    .Q(\integrator_b_sng_comparator.bits_b[6] ));
 sg13g2_dfrbp_1 _3595_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(_0128_),
    .D(net241),
    .Q_N(_1900_),
    .Q(\integrator_b_sng_comparator.bits_b[7] ));
 sg13g2_dfrbp_1 _3596_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(_0129_),
    .D(net29),
    .Q_N(_1899_),
    .Q(\integrator_b_sng_comparator.bits_b[8] ));
 sg13g2_dfrbp_1 _3597_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(_0130_),
    .D(net401),
    .Q_N(_1898_),
    .Q(\input_b_sng_comparator.bits_b[0] ));
 sg13g2_dfrbp_1 _3598_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(_0131_),
    .D(net24),
    .Q_N(\input_b_sng_comparator.bits_b[1] ),
    .Q(_0083_));
 sg13g2_dfrbp_1 _3599_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(_0132_),
    .D(net27),
    .Q_N(_1897_),
    .Q(\input_b_sng_comparator.bits_b[2] ));
 sg13g2_dfrbp_1 _3600_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(_0133_),
    .D(net35),
    .Q_N(_1896_),
    .Q(\integrator_c_sng_comparator.bits_b[3] ));
 sg13g2_dfrbp_1 _3601_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(_0134_),
    .D(net34),
    .Q_N(_1895_),
    .Q(\input_halfprob2_sng_comparator.bits_b[6] ));
 sg13g2_dfrbp_1 _3602_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(_0135_),
    .D(net30),
    .Q_N(_1894_),
    .Q(\input_halfprob2_sng_comparator.bits_b[7] ));
 sg13g2_dfrbp_1 _3603_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(_0136_),
    .D(net36),
    .Q_N(_1893_),
    .Q(\input_halfprob2_sng_comparator.bits_b[8] ));
 sg13g2_dfrbp_1 _3604_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(_0137_),
    .D(net595),
    .Q_N(_1892_),
    .Q(\integrator_a_sng_comparator.bits_b[1] ));
 sg13g2_dfrbp_1 _3605_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(_0138_),
    .D(net317),
    .Q_N(_1891_),
    .Q(\input_halfprob1_sng_comparator.bits_b[0] ));
 sg13g2_dfrbp_1 _3606_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(_0139_),
    .D(net134),
    .Q_N(_1890_),
    .Q(\input_halfprob1_sng_comparator.bits_b[1] ));
 sg13g2_dfrbp_1 _3607_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(_0140_),
    .D(net56),
    .Q_N(_1889_),
    .Q(\input_halfprob2_sng_comparator.bits_b[1] ));
 sg13g2_dfrbp_1 _3608_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(_0141_),
    .D(net42),
    .Q_N(_1888_),
    .Q(\input_halfprob2_sng_comparator.bits_b[2] ));
 sg13g2_dfrbp_1 _3609_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(_0142_),
    .D(net84),
    .Q_N(_1887_),
    .Q(\input_halfprob2_sng_comparator.bits_b[3] ));
 sg13g2_dfrbp_1 _3610_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(_0143_),
    .D(net38),
    .Q_N(_1886_),
    .Q(\input_halfprob2_sng_comparator.bits_b[4] ));
 sg13g2_dfrbp_1 _3611_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(_0144_),
    .D(net41),
    .Q_N(_1885_),
    .Q(\input_halfprob2_sng_comparator.bits_b[5] ));
 sg13g2_dfrbp_1 _3612_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(_0145_),
    .D(net99),
    .Q_N(_1884_),
    .Q(\integrator_a_output.bitseq[0] ));
 sg13g2_dfrbp_1 _3613_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(_0146_),
    .D(net111),
    .Q_N(_1883_),
    .Q(\integrator_a_output.bitseq[1] ));
 sg13g2_dfrbp_1 _3614_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(_0147_),
    .D(net226),
    .Q_N(_1882_),
    .Q(\integrator_a_output.bitseq[2] ));
 sg13g2_dfrbp_1 _3615_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(_0148_),
    .D(_0431_),
    .Q_N(_1881_),
    .Q(\integrator_a_output.bitseq[3] ));
 sg13g2_dfrbp_1 _3616_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(_0149_),
    .D(net136),
    .Q_N(_1880_),
    .Q(\integrator_a_output.bitseq[4] ));
 sg13g2_dfrbp_1 _3617_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(_0150_),
    .D(net92),
    .Q_N(_1879_),
    .Q(\integrator_a_output.bitseq[5] ));
 sg13g2_dfrbp_1 _3618_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(_0151_),
    .D(net188),
    .Q_N(_1878_),
    .Q(\integrator_a_output.bitseq[6] ));
 sg13g2_dfrbp_1 _3619_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(_0152_),
    .D(_0435_),
    .Q_N(_1877_),
    .Q(\integrator_a_output.bitseq[7] ));
 sg13g2_dfrbp_1 _3620_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(_0153_),
    .D(net228),
    .Q_N(\serial_input.adjustment[0] ),
    .Q(_0084_));
 sg13g2_dfrbp_1 _3621_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(_0154_),
    .D(net381),
    .Q_N(_1876_),
    .Q(\serial_input.adjustment[1] ));
 sg13g2_dfrbp_1 _3622_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(_0155_),
    .D(net214),
    .Q_N(_1875_),
    .Q(\serial_input.adjustment[2] ));
 sg13g2_dfrbp_1 _3623_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(_0156_),
    .D(net142),
    .Q_N(\serial_input.adjustment[3] ),
    .Q(_0085_));
 sg13g2_dfrbp_1 _3624_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(_0157_),
    .D(net377),
    .Q_N(_1874_),
    .Q(\serial_input.adjustment[4] ));
 sg13g2_dfrbp_1 _3625_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(_0159_),
    .D(net19),
    .Q_N(\system_integrator_a_counter.init_flag ),
    .Q(_0086_));
 sg13g2_dfrbp_1 _3626_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(_0160_),
    .D(net66),
    .Q_N(_1873_),
    .Q(\integrator_c_output.bitseq[0] ));
 sg13g2_dfrbp_1 _3627_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(_0161_),
    .D(net101),
    .Q_N(_1872_),
    .Q(\integrator_c_output.bitseq[1] ));
 sg13g2_dfrbp_1 _3628_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(_0162_),
    .D(net164),
    .Q_N(_1871_),
    .Q(\integrator_c_output.bitseq[2] ));
 sg13g2_dfrbp_1 _3629_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(_0163_),
    .D(net153),
    .Q_N(_1870_),
    .Q(\integrator_c_output.bitseq[3] ));
 sg13g2_dfrbp_1 _3630_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(_0164_),
    .D(net191),
    .Q_N(_1869_),
    .Q(\integrator_c_output.bitseq[4] ));
 sg13g2_dfrbp_1 _3631_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(_0165_),
    .D(net64),
    .Q_N(_1868_),
    .Q(\integrator_c_output.bitseq[5] ));
 sg13g2_dfrbp_1 _3632_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(_0166_),
    .D(net138),
    .Q_N(_1867_),
    .Q(\integrator_c_output.bitseq[6] ));
 sg13g2_dfrbp_1 _3633_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(_0167_),
    .D(_0448_),
    .Q_N(_1866_),
    .Q(\integrator_c_output.bitseq[7] ));
 sg13g2_dfrbp_1 _3634_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(_0168_),
    .D(net440),
    .Q_N(_1865_),
    .Q(\test_integrator_b_counter.value_output[1] ));
 sg13g2_dfrbp_1 _3635_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(_0169_),
    .D(net483),
    .Q_N(_1864_),
    .Q(\test_integrator_b_counter.value_output[2] ));
 sg13g2_dfrbp_1 _3636_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(_0170_),
    .D(net396),
    .Q_N(_0035_),
    .Q(\test_integrator_b_counter.value_output[3] ));
 sg13g2_dfrbp_1 _3637_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(_0171_),
    .D(net400),
    .Q_N(_0036_),
    .Q(\test_integrator_b_counter.value_output[4] ));
 sg13g2_dfrbp_1 _3638_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(_0172_),
    .D(net299),
    .Q_N(_0037_),
    .Q(\test_integrator_b_counter.value_output[5] ));
 sg13g2_dfrbp_1 _3639_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(_0173_),
    .D(net373),
    .Q_N(_0038_),
    .Q(\test_integrator_b_counter.value_output[6] ));
 sg13g2_dfrbp_1 _3640_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(_0174_),
    .D(net385),
    .Q_N(_0039_),
    .Q(\test_integrator_b_counter.value_output[7] ));
 sg13g2_dfrbp_1 _3641_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(_0175_),
    .D(_0456_),
    .Q_N(_0040_),
    .Q(\test_integrator_b_counter.value_output[8] ));
 sg13g2_dfrbp_1 _3642_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(_0176_),
    .D(net125),
    .Q_N(_1863_),
    .Q(\test_integrator_b_output.bitseq[0] ));
 sg13g2_dfrbp_1 _3643_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(_0177_),
    .D(net140),
    .Q_N(_1862_),
    .Q(\test_integrator_b_output.bitseq[1] ));
 sg13g2_dfrbp_1 _3644_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(_0178_),
    .D(net159),
    .Q_N(_1861_),
    .Q(\test_integrator_b_output.bitseq[2] ));
 sg13g2_dfrbp_1 _3645_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(_0179_),
    .D(net83),
    .Q_N(_1860_),
    .Q(\test_integrator_b_output.bitseq[3] ));
 sg13g2_dfrbp_1 _3646_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(_0180_),
    .D(net185),
    .Q_N(_1859_),
    .Q(\test_integrator_b_output.bitseq[4] ));
 sg13g2_dfrbp_1 _3647_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(_0181_),
    .D(net123),
    .Q_N(_1858_),
    .Q(\test_integrator_b_output.bitseq[5] ));
 sg13g2_dfrbp_1 _3648_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(_0182_),
    .D(net62),
    .Q_N(_1857_),
    .Q(\test_integrator_b_output.bitseq[6] ));
 sg13g2_dfrbp_1 _3649_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(_0183_),
    .D(_0464_),
    .Q_N(_1856_),
    .Q(\test_integrator_b_output.bitseq[7] ));
 sg13g2_dfrbp_1 _3650_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(_0184_),
    .D(net79),
    .Q_N(_1855_),
    .Q(\system_integrator_a_output.bitseq[0] ));
 sg13g2_dfrbp_1 _3651_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(_0185_),
    .D(net72),
    .Q_N(_1854_),
    .Q(\system_integrator_a_output.bitseq[1] ));
 sg13g2_dfrbp_1 _3652_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(_0186_),
    .D(net149),
    .Q_N(_1853_),
    .Q(\system_integrator_a_output.bitseq[2] ));
 sg13g2_dfrbp_1 _3653_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(_0187_),
    .D(net170),
    .Q_N(_1852_),
    .Q(\system_integrator_a_output.bitseq[3] ));
 sg13g2_dfrbp_1 _3654_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(_0188_),
    .D(net94),
    .Q_N(_1851_),
    .Q(\system_integrator_a_output.bitseq[4] ));
 sg13g2_dfrbp_1 _3655_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(_0189_),
    .D(net76),
    .Q_N(_1850_),
    .Q(\system_integrator_a_output.bitseq[5] ));
 sg13g2_dfrbp_1 _3656_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(_0190_),
    .D(net107),
    .Q_N(_1849_),
    .Q(\system_integrator_a_output.bitseq[6] ));
 sg13g2_dfrbp_1 _3657_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(_0191_),
    .D(_0472_),
    .Q_N(_1848_),
    .Q(\system_integrator_a_output.bitseq[7] ));
 sg13g2_dfrbp_1 _3658_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(_0192_),
    .D(_0473_),
    .Q_N(_1847_),
    .Q(\test_integrator_b_counter.value_output[0] ));
 sg13g2_dfrbp_1 _3659_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(_0193_),
    .D(net105),
    .Q_N(_1846_),
    .Q(\system_integrator_b_output.bitseq[0] ));
 sg13g2_dfrbp_1 _3660_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(_0194_),
    .D(net145),
    .Q_N(_1845_),
    .Q(\system_integrator_b_output.bitseq[1] ));
 sg13g2_dfrbp_1 _3661_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(_0195_),
    .D(net162),
    .Q_N(_1844_),
    .Q(\system_integrator_b_output.bitseq[2] ));
 sg13g2_dfrbp_1 _3662_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(_0196_),
    .D(net113),
    .Q_N(_1843_),
    .Q(\system_integrator_b_output.bitseq[3] ));
 sg13g2_dfrbp_1 _3663_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(_0197_),
    .D(net210),
    .Q_N(_1842_),
    .Q(\system_integrator_b_output.bitseq[4] ));
 sg13g2_dfrbp_1 _3664_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(_0198_),
    .D(net127),
    .Q_N(_1841_),
    .Q(\system_integrator_b_output.bitseq[5] ));
 sg13g2_dfrbp_1 _3665_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(_0199_),
    .D(net70),
    .Q_N(_1840_),
    .Q(\system_integrator_b_output.bitseq[6] ));
 sg13g2_dfrbp_1 _3666_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(_0200_),
    .D(_0481_),
    .Q_N(_1839_),
    .Q(\system_integrator_b_output.bitseq[7] ));
 sg13g2_dfrbp_1 _3667_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(_0201_),
    .D(net175),
    .Q_N(_1838_),
    .Q(\test_integrator_b_output.input_bits[0] ));
 sg13g2_dfrbp_1 _3668_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(_0202_),
    .D(net178),
    .Q_N(_1837_),
    .Q(\test_integrator_b_output.input_bits[1] ));
 sg13g2_dfrbp_1 _3669_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(_0203_),
    .D(net251),
    .Q_N(_1836_),
    .Q(\test_integrator_b_output.input_bits[2] ));
 sg13g2_dfrbp_1 _3670_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(_0204_),
    .D(net218),
    .Q_N(_1835_),
    .Q(\test_integrator_b_output.input_bits[3] ));
 sg13g2_dfrbp_1 _3671_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(_0205_),
    .D(net205),
    .Q_N(_1834_),
    .Q(\test_integrator_b_output.input_bits[4] ));
 sg13g2_dfrbp_1 _3672_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(_0206_),
    .D(net224),
    .Q_N(_1833_),
    .Q(\test_integrator_b_output.input_bits[5] ));
 sg13g2_dfrbp_1 _3673_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(_0207_),
    .D(net236),
    .Q_N(_1832_),
    .Q(\test_integrator_b_output.input_bits[6] ));
 sg13g2_dfrbp_1 _3674_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(_0208_),
    .D(net319),
    .Q_N(_1831_),
    .Q(\test_integrator_b_output.input_bits[7] ));
 sg13g2_dfrbp_1 _3675_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(_0209_),
    .D(_0490_),
    .Q_N(_1830_),
    .Q(\test_integrator_b_output.input_bits[8] ));
 sg13g2_dfrbp_1 _3676_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(_0210_),
    .D(_1929_),
    .Q_N(_1829_),
    .Q(\integrator_a_output.output_bit ));
 sg13g2_dfrbp_1 _3677_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(_0211_),
    .D(_0000_),
    .Q_N(_1828_),
    .Q(\integrator_a_output.counter[0] ));
 sg13g2_dfrbp_1 _3678_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(_0212_),
    .D(_0001_),
    .Q_N(_1827_),
    .Q(\integrator_a_output.counter[1] ));
 sg13g2_dfrbp_1 _3679_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(_0213_),
    .D(_0002_),
    .Q_N(_1826_),
    .Q(\integrator_a_output.counter[2] ));
 sg13g2_dfrbp_1 _3680_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(_0214_),
    .D(net365),
    .Q_N(_1825_),
    .Q(\integrator_a_output.counter[3] ));
 sg13g2_dfrbp_1 _3681_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(_0215_),
    .D(net46),
    .Q_N(_0074_),
    .Q(\integrator_a_counter.value_output[0] ));
 sg13g2_dfrbp_1 _3682_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(_0216_),
    .D(net398),
    .Q_N(_0041_),
    .Q(\integrator_a_counter.value_output[1] ));
 sg13g2_dfrbp_1 _3683_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(_0217_),
    .D(_0493_),
    .Q_N(_1824_),
    .Q(\integrator_a_counter.value_output[2] ));
 sg13g2_dfrbp_1 _3684_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(_0218_),
    .D(_0494_),
    .Q_N(_0042_),
    .Q(\integrator_a_counter.value_output[3] ));
 sg13g2_dfrbp_1 _3685_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(_0219_),
    .D(_0495_),
    .Q_N(_1823_),
    .Q(\integrator_a_counter.value_output[4] ));
 sg13g2_dfrbp_1 _3686_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(_0220_),
    .D(net465),
    .Q_N(_0043_),
    .Q(\integrator_a_counter.value_output[5] ));
 sg13g2_dfrbp_1 _3687_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(_0221_),
    .D(_0497_),
    .Q_N(_1822_),
    .Q(\integrator_a_counter.value_output[6] ));
 sg13g2_dfrbp_1 _3688_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(_0222_),
    .D(_0498_),
    .Q_N(_1821_),
    .Q(\integrator_a_counter.value_output[7] ));
 sg13g2_dfrbp_1 _3689_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(_0223_),
    .D(_0499_),
    .Q_N(_0054_),
    .Q(\integrator_a_counter.value_output[8] ));
 sg13g2_dfrbp_1 _3690_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(_0224_),
    .D(_1930_),
    .Q_N(_1820_),
    .Q(\integrator_b_output.output_bit ));
 sg13g2_dfrbp_1 _3691_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(_0225_),
    .D(_0004_),
    .Q_N(_1819_),
    .Q(\integrator_b_output.counter[0] ));
 sg13g2_dfrbp_1 _3692_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(_0226_),
    .D(_0005_),
    .Q_N(_1818_),
    .Q(\integrator_b_output.counter[1] ));
 sg13g2_dfrbp_1 _3693_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(_0227_),
    .D(_0006_),
    .Q_N(_1817_),
    .Q(\integrator_b_output.counter[2] ));
 sg13g2_dfrbp_1 _3694_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(_0228_),
    .D(net338),
    .Q_N(_1816_),
    .Q(\integrator_b_output.counter[3] ));
 sg13g2_dfrbp_1 _3695_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(_0229_),
    .D(net58),
    .Q_N(_0073_),
    .Q(\integrator_b_counter.value_output[0] ));
 sg13g2_dfrbp_1 _3696_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(_0230_),
    .D(net388),
    .Q_N(_0044_),
    .Q(\integrator_b_counter.value_output[1] ));
 sg13g2_dfrbp_1 _3697_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(_0231_),
    .D(_0502_),
    .Q_N(_1815_),
    .Q(\integrator_b_counter.value_output[2] ));
 sg13g2_dfrbp_1 _3698_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(_0232_),
    .D(net438),
    .Q_N(_0045_),
    .Q(\integrator_b_counter.value_output[3] ));
 sg13g2_dfrbp_1 _3699_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(_0233_),
    .D(_0504_),
    .Q_N(_1814_),
    .Q(\integrator_b_counter.value_output[4] ));
 sg13g2_dfrbp_1 _3700_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(_0234_),
    .D(net449),
    .Q_N(_0046_),
    .Q(\integrator_b_counter.value_output[5] ));
 sg13g2_dfrbp_1 _3701_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(_0235_),
    .D(_0506_),
    .Q_N(_1813_),
    .Q(\integrator_b_counter.value_output[6] ));
 sg13g2_dfrbp_1 _3702_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(_0236_),
    .D(_0507_),
    .Q_N(_1812_),
    .Q(\integrator_b_counter.value_output[7] ));
 sg13g2_dfrbp_1 _3703_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(_0237_),
    .D(_0508_),
    .Q_N(_0051_),
    .Q(\integrator_b_counter.value_output[8] ));
 sg13g2_dfrbp_1 _3704_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(_0238_),
    .D(net173),
    .Q_N(_1811_),
    .Q(\integrator_c_output.output_bit ));
 sg13g2_dfrbp_1 _3705_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(_0239_),
    .D(_0008_),
    .Q_N(_1810_),
    .Q(\integrator_c_output.counter[0] ));
 sg13g2_dfrbp_1 _3706_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(_0240_),
    .D(_0009_),
    .Q_N(_1809_),
    .Q(\integrator_c_output.counter[1] ));
 sg13g2_dfrbp_1 _3707_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(_0241_),
    .D(_0010_),
    .Q_N(_1808_),
    .Q(\integrator_c_output.counter[2] ));
 sg13g2_dfrbp_1 _3708_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(_0242_),
    .D(net304),
    .Q_N(_1807_),
    .Q(\integrator_c_output.counter[3] ));
 sg13g2_dfrbp_1 _3709_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(_0243_),
    .D(net48),
    .Q_N(_0072_),
    .Q(\integrator_c_counter.value_output[0] ));
 sg13g2_dfrbp_1 _3710_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(_0244_),
    .D(net416),
    .Q_N(_0047_),
    .Q(\integrator_c_counter.value_output[1] ));
 sg13g2_dfrbp_1 _3711_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(_0245_),
    .D(net457),
    .Q_N(_1806_),
    .Q(\integrator_c_counter.value_output[2] ));
 sg13g2_dfrbp_1 _3712_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(_0246_),
    .D(net408),
    .Q_N(_0048_),
    .Q(\integrator_c_counter.value_output[3] ));
 sg13g2_dfrbp_1 _3713_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(_0247_),
    .D(_0513_),
    .Q_N(_1805_),
    .Q(\integrator_c_counter.value_output[4] ));
 sg13g2_dfrbp_1 _3714_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(_0248_),
    .D(net411),
    .Q_N(_0049_),
    .Q(\integrator_c_counter.value_output[5] ));
 sg13g2_dfrbp_1 _3715_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(_0249_),
    .D(_0515_),
    .Q_N(_1804_),
    .Q(\integrator_c_counter.value_output[6] ));
 sg13g2_dfrbp_1 _3716_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(_0250_),
    .D(_0516_),
    .Q_N(_1803_),
    .Q(\integrator_c_counter.value_output[7] ));
 sg13g2_dfrbp_1 _3717_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(_0251_),
    .D(_0517_),
    .Q_N(_0053_),
    .Q(\integrator_c_counter.value_output[8] ));
 sg13g2_dfrbp_1 _3718_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(_0252_),
    .D(net240),
    .Q_N(_1802_),
    .Q(\system_integrator_a_output.output_bit ));
 sg13g2_dfrbp_1 _3719_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(_0253_),
    .D(_0013_),
    .Q_N(_1801_),
    .Q(\system_integrator_a_output.counter[0] ));
 sg13g2_dfrbp_1 _3720_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(_0254_),
    .D(_0014_),
    .Q_N(_1800_),
    .Q(\system_integrator_a_output.counter[1] ));
 sg13g2_dfrbp_1 _3721_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(_0255_),
    .D(_0015_),
    .Q_N(_1799_),
    .Q(\system_integrator_a_output.counter[2] ));
 sg13g2_dfrbp_1 _3722_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(_0256_),
    .D(net309),
    .Q_N(_1798_),
    .Q(\system_integrator_a_output.counter[3] ));
 sg13g2_dfrbp_1 _3723_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(_0257_),
    .D(net103),
    .Q_N(_0030_),
    .Q(\system_integrator_a_counter.value_output[0] ));
 sg13g2_dfrbp_1 _3724_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(_0258_),
    .D(net462),
    .Q_N(_0031_),
    .Q(\system_integrator_a_counter.value_output[1] ));
 sg13g2_dfrbp_1 _3725_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(_0259_),
    .D(_0520_),
    .Q_N(_1797_),
    .Q(\system_integrator_a_counter.value_output[2] ));
 sg13g2_dfrbp_1 _3726_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(_0260_),
    .D(_0521_),
    .Q_N(_1796_),
    .Q(\system_integrator_a_counter.value_output[3] ));
 sg13g2_dfrbp_1 _3727_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(_0261_),
    .D(_0522_),
    .Q_N(_1795_),
    .Q(\system_integrator_a_counter.value_output[4] ));
 sg13g2_dfrbp_1 _3728_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(_0262_),
    .D(_0523_),
    .Q_N(_1794_),
    .Q(\system_integrator_a_counter.value_output[5] ));
 sg13g2_dfrbp_1 _3729_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(_0263_),
    .D(_0524_),
    .Q_N(_1793_),
    .Q(\system_integrator_a_counter.value_output[6] ));
 sg13g2_dfrbp_1 _3730_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(_0264_),
    .D(_0525_),
    .Q_N(_1792_),
    .Q(\system_integrator_a_counter.value_output[7] ));
 sg13g2_dfrbp_1 _3731_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(_0265_),
    .D(_0526_),
    .Q_N(_1791_),
    .Q(\system_integrator_a_counter.value_output[8] ));
 sg13g2_dfrbp_1 _3732_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(_0266_),
    .D(_1933_),
    .Q_N(_1790_),
    .Q(\system_integrator_b_output.output_bit ));
 sg13g2_dfrbp_1 _3733_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(_0267_),
    .D(_0017_),
    .Q_N(_1789_),
    .Q(\system_integrator_b_output.counter[0] ));
 sg13g2_dfrbp_1 _3734_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(_0268_),
    .D(_0018_),
    .Q_N(_1788_),
    .Q(\system_integrator_b_output.counter[1] ));
 sg13g2_dfrbp_1 _3735_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(_0269_),
    .D(_0019_),
    .Q_N(_1787_),
    .Q(\system_integrator_b_output.counter[2] ));
 sg13g2_dfrbp_1 _3736_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(_0270_),
    .D(net321),
    .Q_N(_1786_),
    .Q(\system_integrator_b_output.counter[3] ));
 sg13g2_dfrbp_1 _3737_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(_0271_),
    .D(_0527_),
    .Q_N(_1785_),
    .Q(\system_integrator_b_counter.value_output[0] ));
 sg13g2_dfrbp_1 _3738_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(_0272_),
    .D(net479),
    .Q_N(_0032_),
    .Q(\system_integrator_b_counter.value_output[1] ));
 sg13g2_dfrbp_1 _3739_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(_0273_),
    .D(_0529_),
    .Q_N(_1784_),
    .Q(\system_integrator_b_counter.value_output[2] ));
 sg13g2_dfrbp_1 _3740_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(_0274_),
    .D(_0530_),
    .Q_N(_1783_),
    .Q(\system_integrator_b_counter.value_output[3] ));
 sg13g2_dfrbp_1 _3741_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(_0275_),
    .D(_0531_),
    .Q_N(_1782_),
    .Q(\system_integrator_b_counter.value_output[4] ));
 sg13g2_dfrbp_1 _3742_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(_0276_),
    .D(_0532_),
    .Q_N(_1781_),
    .Q(\system_integrator_b_counter.value_output[5] ));
 sg13g2_dfrbp_1 _3743_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(_0277_),
    .D(_0533_),
    .Q_N(_1780_),
    .Q(\system_integrator_b_counter.value_output[6] ));
 sg13g2_dfrbp_1 _3744_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(_0278_),
    .D(_0534_),
    .Q_N(_1779_),
    .Q(\system_integrator_b_counter.value_output[7] ));
 sg13g2_dfrbp_1 _3745_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(_0279_),
    .D(_0535_),
    .Q_N(_0029_),
    .Q(\system_integrator_b_counter.value_output[8] ));
 sg13g2_dfrbp_1 _3746_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(_0280_),
    .D(net51),
    .Q_N(_1778_),
    .Q(\test_integrator_a_output.output_bit ));
 sg13g2_dfrbp_1 _3747_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(_0281_),
    .D(_0021_),
    .Q_N(_1777_),
    .Q(\test_integrator_a_output.counter[0] ));
 sg13g2_dfrbp_1 _3748_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(_0282_),
    .D(_0022_),
    .Q_N(_1776_),
    .Q(\test_integrator_a_output.counter[1] ));
 sg13g2_dfrbp_1 _3749_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(_0283_),
    .D(_0023_),
    .Q_N(_1775_),
    .Q(\test_integrator_a_output.counter[2] ));
 sg13g2_dfrbp_1 _3750_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(_0284_),
    .D(net357),
    .Q_N(_1774_),
    .Q(\test_integrator_a_output.counter[3] ));
 sg13g2_dfrbp_1 _3751_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(_0285_),
    .D(_0536_),
    .Q_N(_0033_),
    .Q(\test_integrator_a_counter.value_output[0] ));
 sg13g2_dfrbp_1 _3752_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(_0286_),
    .D(net419),
    .Q_N(_0034_),
    .Q(\test_integrator_a_counter.value_output[1] ));
 sg13g2_dfrbp_1 _3753_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(_0287_),
    .D(_0538_),
    .Q_N(_1773_),
    .Q(\test_integrator_a_counter.value_output[2] ));
 sg13g2_dfrbp_1 _3754_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(_0288_),
    .D(_0539_),
    .Q_N(_1772_),
    .Q(\test_integrator_a_counter.value_output[3] ));
 sg13g2_dfrbp_1 _3755_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(_0289_),
    .D(_0540_),
    .Q_N(_1771_),
    .Q(\test_integrator_a_counter.value_output[4] ));
 sg13g2_dfrbp_1 _3756_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(_0290_),
    .D(_0541_),
    .Q_N(_1770_),
    .Q(\test_integrator_a_counter.value_output[5] ));
 sg13g2_dfrbp_1 _3757_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(_0291_),
    .D(_0542_),
    .Q_N(_1769_),
    .Q(\test_integrator_a_counter.value_output[6] ));
 sg13g2_dfrbp_1 _3758_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(_0292_),
    .D(_0543_),
    .Q_N(_1768_),
    .Q(\test_integrator_a_counter.value_output[7] ));
 sg13g2_dfrbp_1 _3759_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(_0293_),
    .D(net375),
    .Q_N(_0050_),
    .Q(\test_integrator_a_counter.value_output[8] ));
 sg13g2_dfrbp_1 _3760_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(_0294_),
    .D(_1935_),
    .Q_N(_1767_),
    .Q(\test_integrator_b_output.output_bit ));
 sg13g2_dfrbp_1 _3761_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(_0295_),
    .D(_0025_),
    .Q_N(_1766_),
    .Q(\test_integrator_b_output.counter[0] ));
 sg13g2_dfrbp_1 _3762_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(_0296_),
    .D(_0026_),
    .Q_N(_1765_),
    .Q(\test_integrator_b_output.counter[1] ));
 sg13g2_dfrbp_1 _3763_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(_0297_),
    .D(_0027_),
    .Q_N(_1764_),
    .Q(\test_integrator_b_output.counter[2] ));
 sg13g2_dfrbp_1 _3764_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(_0298_),
    .D(net393),
    .Q_N(_1763_),
    .Q(\test_integrator_b_output.counter[3] ));
 sg13g2_dfrbp_1 _3765_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(_0299_),
    .D(net245),
    .Q_N(_1762_),
    .Q(\test_integrator_a_output.bitseq[0] ));
 sg13g2_dfrbp_1 _3766_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(_0300_),
    .D(net155),
    .Q_N(_1761_),
    .Q(\test_integrator_a_output.bitseq[1] ));
 sg13g2_dfrbp_1 _3767_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(_0301_),
    .D(net90),
    .Q_N(_1760_),
    .Q(\test_integrator_a_output.bitseq[2] ));
 sg13g2_dfrbp_1 _3768_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(_0302_),
    .D(net68),
    .Q_N(_1759_),
    .Q(\test_integrator_a_output.bitseq[3] ));
 sg13g2_dfrbp_1 _3769_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(_0303_),
    .D(net151),
    .Q_N(_1758_),
    .Q(\test_integrator_a_output.bitseq[4] ));
 sg13g2_dfrbp_1 _3770_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(_0304_),
    .D(net131),
    .Q_N(_1757_),
    .Q(\test_integrator_a_output.bitseq[5] ));
 sg13g2_dfrbp_1 _3771_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(_0305_),
    .D(net238),
    .Q_N(_1756_),
    .Q(\test_integrator_a_output.bitseq[6] ));
 sg13g2_dfrbp_1 _3772_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(_0306_),
    .D(_0552_),
    .Q_N(_1755_),
    .Q(\test_integrator_a_output.bitseq[7] ));
 sg13g2_dfrbp_1 _3773_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(_0307_),
    .D(net342),
    .Q_N(_1754_),
    .Q(\integrator_a_output.input_bits[0] ));
 sg13g2_dfrbp_1 _3774_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(_0308_),
    .D(net203),
    .Q_N(_1753_),
    .Q(\integrator_a_output.input_bits[1] ));
 sg13g2_dfrbp_1 _3775_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(_0309_),
    .D(net197),
    .Q_N(_1752_),
    .Q(\integrator_a_output.input_bits[2] ));
 sg13g2_dfrbp_1 _3776_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(_0310_),
    .D(net275),
    .Q_N(_1751_),
    .Q(\integrator_a_output.input_bits[3] ));
 sg13g2_dfrbp_1 _3777_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(_0311_),
    .D(net157),
    .Q_N(_1750_),
    .Q(\integrator_a_output.input_bits[4] ));
 sg13g2_dfrbp_1 _3778_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(_0312_),
    .D(net249),
    .Q_N(_1749_),
    .Q(\integrator_a_output.input_bits[5] ));
 sg13g2_dfrbp_1 _3779_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(_0313_),
    .D(net195),
    .Q_N(_1748_),
    .Q(\integrator_a_output.input_bits[6] ));
 sg13g2_dfrbp_1 _3780_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(_0314_),
    .D(net263),
    .Q_N(_1747_),
    .Q(\integrator_a_output.input_bits[7] ));
 sg13g2_dfrbp_1 _3781_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(_0315_),
    .D(_0561_),
    .Q_N(_1746_),
    .Q(\integrator_a_output.input_bits[8] ));
 sg13g2_dfrbp_1 _3782_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(_0316_),
    .D(net220),
    .Q_N(_1745_),
    .Q(\integrator_b_output.input_bits[0] ));
 sg13g2_dfrbp_1 _3783_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(_0317_),
    .D(net147),
    .Q_N(_1744_),
    .Q(\integrator_b_output.input_bits[1] ));
 sg13g2_dfrbp_1 _3784_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(_0318_),
    .D(net199),
    .Q_N(_1743_),
    .Q(\integrator_b_output.input_bits[2] ));
 sg13g2_dfrbp_1 _3785_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(_0319_),
    .D(net193),
    .Q_N(_1742_),
    .Q(\integrator_b_output.input_bits[3] ));
 sg13g2_dfrbp_1 _3786_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(_0320_),
    .D(net181),
    .Q_N(_1741_),
    .Q(\integrator_b_output.input_bits[4] ));
 sg13g2_dfrbp_1 _3787_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(_0321_),
    .D(net183),
    .Q_N(_1740_),
    .Q(\integrator_b_output.input_bits[5] ));
 sg13g2_dfrbp_1 _3788_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(_0322_),
    .D(net133),
    .Q_N(_1739_),
    .Q(\integrator_b_output.input_bits[6] ));
 sg13g2_dfrbp_1 _3789_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(_0323_),
    .D(net119),
    .Q_N(_1738_),
    .Q(\integrator_b_output.input_bits[7] ));
 sg13g2_dfrbp_1 _3790_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(_0324_),
    .D(_0570_),
    .Q_N(_1737_),
    .Q(\integrator_b_output.input_bits[8] ));
 sg13g2_dfrbp_1 _3791_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(_0325_),
    .D(_0571_),
    .Q_N(_1736_),
    .Q(\integrator_c_output.input_bits[0] ));
 sg13g2_dfrbp_1 _3792_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(_0326_),
    .D(net267),
    .Q_N(_1735_),
    .Q(\integrator_c_output.input_bits[1] ));
 sg13g2_dfrbp_1 _3793_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(_0327_),
    .D(net168),
    .Q_N(_1734_),
    .Q(\integrator_c_output.input_bits[2] ));
 sg13g2_dfrbp_1 _3794_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(_0328_),
    .D(net279),
    .Q_N(_1733_),
    .Q(\integrator_c_output.input_bits[3] ));
 sg13g2_dfrbp_1 _3795_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(_0329_),
    .D(net346),
    .Q_N(_1732_),
    .Q(\integrator_c_output.input_bits[4] ));
 sg13g2_dfrbp_1 _3796_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(_0330_),
    .D(net316),
    .Q_N(_1731_),
    .Q(\integrator_c_output.input_bits[5] ));
 sg13g2_dfrbp_1 _3797_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(_0331_),
    .D(net323),
    .Q_N(_1730_),
    .Q(\integrator_c_output.input_bits[6] ));
 sg13g2_dfrbp_1 _3798_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(_0332_),
    .D(net256),
    .Q_N(_1729_),
    .Q(\integrator_c_output.input_bits[7] ));
 sg13g2_dfrbp_1 _3799_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(_0333_),
    .D(_0579_),
    .Q_N(_1728_),
    .Q(\integrator_c_output.input_bits[8] ));
 sg13g2_dfrbp_1 _3800_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(_0334_),
    .D(_0580_),
    .Q_N(_1727_),
    .Q(\system_integrator_a_output.input_bits[0] ));
 sg13g2_dfrbp_1 _3801_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(_0335_),
    .D(net233),
    .Q_N(_1726_),
    .Q(\system_integrator_a_output.input_bits[1] ));
 sg13g2_dfrbp_1 _3802_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(_0336_),
    .D(net201),
    .Q_N(_1725_),
    .Q(\system_integrator_a_output.input_bits[2] ));
 sg13g2_dfrbp_1 _3803_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(_0337_),
    .D(net247),
    .Q_N(_1724_),
    .Q(\system_integrator_a_output.input_bits[3] ));
 sg13g2_dfrbp_1 _3804_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(_0338_),
    .D(net277),
    .Q_N(_1723_),
    .Q(\system_integrator_a_output.input_bits[4] ));
 sg13g2_dfrbp_1 _3805_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(_0339_),
    .D(net208),
    .Q_N(_1722_),
    .Q(\system_integrator_a_output.input_bits[5] ));
 sg13g2_dfrbp_1 _3806_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(_0340_),
    .D(net289),
    .Q_N(_1721_),
    .Q(\system_integrator_a_output.input_bits[6] ));
 sg13g2_dfrbp_1 _3807_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(_0341_),
    .D(net216),
    .Q_N(_1720_),
    .Q(\system_integrator_a_output.input_bits[7] ));
 sg13g2_dfrbp_1 _3808_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(_0342_),
    .D(_0588_),
    .Q_N(_1719_),
    .Q(\system_integrator_a_output.input_bits[8] ));
 sg13g2_dfrbp_1 _3809_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(_0343_),
    .D(net287),
    .Q_N(_1718_),
    .Q(\system_integrator_b_output.input_bits[0] ));
 sg13g2_dfrbp_1 _3810_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(_0344_),
    .D(net294),
    .Q_N(_1717_),
    .Q(\system_integrator_b_output.input_bits[1] ));
 sg13g2_dfrbp_1 _3811_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(_0345_),
    .D(net344),
    .Q_N(_1716_),
    .Q(\system_integrator_b_output.input_bits[2] ));
 sg13g2_dfrbp_1 _3812_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(_0346_),
    .D(net354),
    .Q_N(_1715_),
    .Q(\system_integrator_b_output.input_bits[3] ));
 sg13g2_dfrbp_1 _3813_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(_0347_),
    .D(net335),
    .Q_N(_1714_),
    .Q(\system_integrator_b_output.input_bits[4] ));
 sg13g2_dfrbp_1 _3814_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(_0348_),
    .D(net273),
    .Q_N(_1713_),
    .Q(\system_integrator_b_output.input_bits[5] ));
 sg13g2_dfrbp_1 _3815_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(_0349_),
    .D(net261),
    .Q_N(_1712_),
    .Q(\system_integrator_b_output.input_bits[6] ));
 sg13g2_dfrbp_1 _3816_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(_0350_),
    .D(net281),
    .Q_N(_1711_),
    .Q(\system_integrator_b_output.input_bits[7] ));
 sg13g2_dfrbp_1 _3817_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(_0351_),
    .D(_0597_),
    .Q_N(_1710_),
    .Q(\system_integrator_b_output.input_bits[8] ));
 sg13g2_dfrbp_1 _3818_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(_0352_),
    .D(_0598_),
    .Q_N(_1709_),
    .Q(\test_integrator_a_output.input_bits[0] ));
 sg13g2_dfrbp_1 _3819_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(_0353_),
    .D(net222),
    .Q_N(_1708_),
    .Q(\test_integrator_a_output.input_bits[1] ));
 sg13g2_dfrbp_1 _3820_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(_0354_),
    .D(net283),
    .Q_N(_1707_),
    .Q(\test_integrator_a_output.input_bits[2] ));
 sg13g2_dfrbp_1 _3821_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(_0355_),
    .D(net340),
    .Q_N(_1706_),
    .Q(\test_integrator_a_output.input_bits[3] ));
 sg13g2_dfrbp_1 _3822_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(_0356_),
    .D(net330),
    .Q_N(_1705_),
    .Q(\test_integrator_a_output.input_bits[4] ));
 sg13g2_dfrbp_1 _3823_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(_0357_),
    .D(net362),
    .Q_N(_1704_),
    .Q(\test_integrator_a_output.input_bits[5] ));
 sg13g2_dfrbp_1 _3824_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(_0358_),
    .D(net296),
    .Q_N(_1703_),
    .Q(\test_integrator_a_output.input_bits[6] ));
 sg13g2_dfrbp_1 _3825_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(_0359_),
    .D(net265),
    .Q_N(_1702_),
    .Q(\test_integrator_a_output.input_bits[7] ));
 sg13g2_dfrbp_1 _3826_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(_0360_),
    .D(net367),
    .Q_N(_1701_),
    .Q(\test_integrator_a_output.input_bits[8] ));
 sg13g2_dfrbp_1 _3827_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(_0361_),
    .D(net23),
    .Q_N(_1657_),
    .Q(\clk_counter[0] ));
 sg13g2_dfrbp_1 _3828_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(_0362_),
    .D(net424),
    .Q_N(_1700_),
    .Q(\clk_counter[1] ));
 sg13g2_dfrbp_1 _3829_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(_0363_),
    .D(net477),
    .Q_N(_1699_),
    .Q(\clk_counter[2] ));
 sg13g2_dfrbp_1 _3830_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(_0364_),
    .D(net422),
    .Q_N(_1698_),
    .Q(\clk_counter[3] ));
 sg13g2_dfrbp_1 _3831_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(_0365_),
    .D(_0066_),
    .Q_N(_1697_),
    .Q(\clk_counter[4] ));
 sg13g2_dfrbp_1 _3832_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(_0366_),
    .D(_0067_),
    .Q_N(_1696_),
    .Q(\clk_counter[5] ));
 sg13g2_dfrbp_1 _3833_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(_0367_),
    .D(net302),
    .Q_N(_1695_),
    .Q(\clk_counter[6] ));
 sg13g2_dfrbp_1 _3834_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(_0368_),
    .D(net254),
    .Q_N(_1694_),
    .Q(\clk_counter[7] ));
 sg13g2_dfrbp_1 _3835_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(_0369_),
    .D(net379),
    .Q_N(_1693_),
    .Q(\clk_counter[8] ));
 sg13g2_dfrbp_1 _3836_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(_0370_),
    .D(_0071_),
    .Q_N(_1692_),
    .Q(\clk_counter[9] ));
 sg13g2_dfrbp_1 _3837_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(_0371_),
    .D(net369),
    .Q_N(_1691_),
    .Q(\clk_counter[10] ));
 sg13g2_dfrbp_1 _3838_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(_0372_),
    .D(net271),
    .Q_N(_1690_),
    .Q(\clk_counter[11] ));
 sg13g2_dfrbp_1 _3839_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(_0373_),
    .D(_0057_),
    .Q_N(_1689_),
    .Q(\clk_counter[12] ));
 sg13g2_dfrbp_1 _3840_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(_0374_),
    .D(net97),
    .Q_N(_1688_),
    .Q(\clk_counter[13] ));
 sg13g2_dfrbp_1 _3841_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(_0375_),
    .D(_0059_),
    .Q_N(_1687_),
    .Q(\clk_counter[14] ));
 sg13g2_dfrbp_1 _3842_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(_0376_),
    .D(_0060_),
    .Q_N(_1686_),
    .Q(\clk_counter[15] ));
 sg13g2_dfrbp_1 _3843_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(_0377_),
    .D(net427),
    .Q_N(_1685_),
    .Q(\clk_counter[16] ));
 sg13g2_dfrbp_1 _3844_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(_0378_),
    .D(net307),
    .Q_N(_1684_),
    .Q(\clk_counter[17] ));
 sg13g2_dfrbp_1 _3845_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(_0379_),
    .D(net60),
    .Q_N(_1683_),
    .Q(\input_a_sng_comparator.bits_a[0] ));
 sg13g2_dfrbp_1 _3846_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(_0380_),
    .D(net121),
    .Q_N(_1682_),
    .Q(\input_a_sng_comparator.bits_a[1] ));
 sg13g2_dfrbp_1 _3847_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(_0381_),
    .D(_0609_),
    .Q_N(_1681_),
    .Q(\input_a_sng_comparator.bits_a[2] ));
 sg13g2_dfrbp_1 _3848_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(_0382_),
    .D(_0610_),
    .Q_N(_1680_),
    .Q(\input_a_sng_comparator.bits_a[3] ));
 sg13g2_dfrbp_1 _3849_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(_0383_),
    .D(_0611_),
    .Q_N(_1679_),
    .Q(\input_a_sng_comparator.bits_a[4] ));
 sg13g2_dfrbp_1 _3850_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(_0384_),
    .D(_0612_),
    .Q_N(_1678_),
    .Q(\input_a_sng_comparator.bits_a[5] ));
 sg13g2_dfrbp_1 _3851_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(_0385_),
    .D(_0613_),
    .Q_N(_1677_),
    .Q(\input_a_sng_comparator.bits_a[6] ));
 sg13g2_dfrbp_1 _3852_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(_0386_),
    .D(_0614_),
    .Q_N(_1676_),
    .Q(\input_a_sng_comparator.bits_a[7] ));
 sg13g2_dfrbp_1 _3853_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(_0387_),
    .D(net405),
    .Q_N(_1675_),
    .Q(\input_a_sng_comparator.bits_a[8] ));
 sg13g2_dfrbp_1 _3854_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(_0388_),
    .D(_0012_),
    .Q_N(_0052_),
    .Q(\serial_input.loop ));
 sg13g2_dfrbp_1 _3855_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(_0389_),
    .D(_0616_),
    .Q_N(_1674_),
    .Q(\integrator_b_output.bitseq[0] ));
 sg13g2_dfrbp_1 _3856_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(_0390_),
    .D(net129),
    .Q_N(_1673_),
    .Q(\integrator_b_output.bitseq[1] ));
 sg13g2_dfrbp_1 _3857_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(_0391_),
    .D(net87),
    .Q_N(_1672_),
    .Q(\integrator_b_output.bitseq[2] ));
 sg13g2_dfrbp_1 _3858_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(_0392_),
    .D(net115),
    .Q_N(_1671_),
    .Q(\integrator_b_output.bitseq[3] ));
 sg13g2_dfrbp_1 _3859_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(_0393_),
    .D(net109),
    .Q_N(_1670_),
    .Q(\integrator_b_output.bitseq[4] ));
 sg13g2_dfrbp_1 _3860_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(_0394_),
    .D(net81),
    .Q_N(_1669_),
    .Q(\integrator_b_output.bitseq[5] ));
 sg13g2_dfrbp_1 _3861_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(_0395_),
    .D(net117),
    .Q_N(_1668_),
    .Q(\integrator_b_output.bitseq[6] ));
 sg13g2_dfrbp_1 _3862_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(_0396_),
    .D(_0623_),
    .Q_N(_1667_),
    .Q(\integrator_b_output.bitseq[7] ));
 sg13g2_dfrbp_1 _3863_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(_0397_),
    .D(net269),
    .Q_N(_1666_),
    .Q(\input_b_sng_comparator.bits_a[0] ));
 sg13g2_dfrbp_1 _3864_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(_0398_),
    .D(net285),
    .Q_N(_1665_),
    .Q(\input_b_sng_comparator.bits_a[1] ));
 sg13g2_dfrbp_1 _3865_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(_0399_),
    .D(net259),
    .Q_N(_1664_),
    .Q(\input_b_sng_comparator.bits_a[2] ));
 sg13g2_dfrbp_1 _3866_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(_0400_),
    .D(_0627_),
    .Q_N(_1663_),
    .Q(\input_b_sng_comparator.bits_a[3] ));
 sg13g2_dfrbp_1 _3867_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(_0401_),
    .D(net314),
    .Q_N(_1662_),
    .Q(\input_b_sng_comparator.bits_a[4] ));
 sg13g2_dfrbp_1 _3868_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(_0402_),
    .D(net359),
    .Q_N(_1661_),
    .Q(\input_b_sng_comparator.bits_a[5] ));
 sg13g2_dfrbp_1 _3869_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(_0403_),
    .D(net349),
    .Q_N(_1660_),
    .Q(\input_b_sng_comparator.bits_a[6] ));
 sg13g2_dfrbp_1 _3870_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(_0404_),
    .D(_0631_),
    .Q_N(_1659_),
    .Q(\input_b_sng_comparator.bits_a[7] ));
 sg13g2_dfrbp_1 _3871_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(_0405_),
    .D(net326),
    .Q_N(_1658_),
    .Q(\input_b_sng_comparator.bits_a[8] ));
 sg13g2_buf_2 clkbuf_leaf_0_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_tielo tt_um_stochastic_integrator_tt9_CL123abc_4 (.L_LO(net4));
 sg13g2_tielo tt_um_stochastic_integrator_tt9_CL123abc_5 (.L_LO(net5));
 sg13g2_tielo tt_um_stochastic_integrator_tt9_CL123abc_6 (.L_LO(net6));
 sg13g2_tielo tt_um_stochastic_integrator_tt9_CL123abc_7 (.L_LO(net7));
 sg13g2_tielo tt_um_stochastic_integrator_tt9_CL123abc_8 (.L_LO(net8));
 sg13g2_tielo tt_um_stochastic_integrator_tt9_CL123abc_9 (.L_LO(net9));
 sg13g2_tielo tt_um_stochastic_integrator_tt9_CL123abc_10 (.L_LO(net10));
 sg13g2_tielo tt_um_stochastic_integrator_tt9_CL123abc_11 (.L_LO(net11));
 sg13g2_tielo tt_um_stochastic_integrator_tt9_CL123abc_12 (.L_LO(net12));
 sg13g2_tielo tt_um_stochastic_integrator_tt9_CL123abc_13 (.L_LO(net13));
 sg13g2_tielo tt_um_stochastic_integrator_tt9_CL123abc_14 (.L_LO(net14));
 sg13g2_tielo tt_um_stochastic_integrator_tt9_CL123abc_15 (.L_LO(net15));
 sg13g2_tielo tt_um_stochastic_integrator_tt9_CL123abc_16 (.L_LO(net16));
 sg13g2_tielo tt_um_stochastic_integrator_tt9_CL123abc_17 (.L_LO(net17));
 sg13g2_tielo tt_um_stochastic_integrator_tt9_CL123abc_18 (.L_LO(net18));
 sg13g2_tiehi _3625__19 (.L_HI(net19));
 sg13g2_buf_2 _3889_ (.A(\integrator_a_output.output_bit ),
    .X(uo_out[0]));
 sg13g2_buf_2 _3890_ (.A(\integrator_b_output.output_bit ),
    .X(uo_out[1]));
 sg13g2_buf_1 _3891_ (.A(\integrator_c_output.output_bit ),
    .X(uo_out[2]));
 sg13g2_buf_1 _3892_ (.A(\system_integrator_a_output.output_bit ),
    .X(uo_out[3]));
 sg13g2_buf_1 _3893_ (.A(\system_integrator_b_output.output_bit ),
    .X(uo_out[4]));
 sg13g2_buf_1 _3894_ (.A(\test_integrator_a_output.output_bit ),
    .X(uo_out[5]));
 sg13g2_buf_1 _3895_ (.A(\test_integrator_b_output.output_bit ),
    .X(uo_out[6]));
 sg13g2_buf_2 _3896_ (.A(integrator_c_sn_bit),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout508 (.A(_1420_),
    .X(net508));
 sg13g2_buf_2 fanout509 (.A(net510),
    .X(net509));
 sg13g2_buf_2 fanout510 (.A(_1269_),
    .X(net510));
 sg13g2_buf_2 fanout511 (.A(net512),
    .X(net511));
 sg13g2_buf_2 fanout512 (.A(_1214_),
    .X(net512));
 sg13g2_buf_2 fanout513 (.A(_0913_),
    .X(net513));
 sg13g2_buf_1 fanout514 (.A(_0913_),
    .X(net514));
 sg13g2_buf_2 fanout515 (.A(net517),
    .X(net515));
 sg13g2_buf_1 fanout516 (.A(net517),
    .X(net516));
 sg13g2_buf_2 fanout517 (.A(_1127_),
    .X(net517));
 sg13g2_buf_2 fanout518 (.A(_1004_),
    .X(net518));
 sg13g2_buf_2 fanout519 (.A(_0828_),
    .X(net519));
 sg13g2_buf_2 fanout520 (.A(_1258_),
    .X(net520));
 sg13g2_buf_2 fanout521 (.A(_1258_),
    .X(net521));
 sg13g2_buf_2 fanout522 (.A(net523),
    .X(net522));
 sg13g2_buf_2 fanout523 (.A(_1204_),
    .X(net523));
 sg13g2_buf_4 fanout524 (.X(net524),
    .A(_1118_));
 sg13g2_buf_2 fanout525 (.A(_1118_),
    .X(net525));
 sg13g2_buf_4 fanout526 (.X(net526),
    .A(_1085_));
 sg13g2_buf_4 fanout527 (.X(net527),
    .A(_0993_));
 sg13g2_buf_4 fanout528 (.X(net528),
    .A(_0901_));
 sg13g2_buf_2 fanout529 (.A(_0901_),
    .X(net529));
 sg13g2_buf_2 fanout530 (.A(net532),
    .X(net530));
 sg13g2_buf_1 fanout531 (.A(net532),
    .X(net531));
 sg13g2_buf_2 fanout532 (.A(_0820_),
    .X(net532));
 sg13g2_buf_4 fanout533 (.X(net533),
    .A(net534));
 sg13g2_buf_4 fanout534 (.X(net534),
    .A(_0669_));
 sg13g2_buf_2 fanout535 (.A(_0669_),
    .X(net535));
 sg13g2_buf_2 fanout536 (.A(net537),
    .X(net536));
 sg13g2_buf_2 fanout537 (.A(_1509_),
    .X(net537));
 sg13g2_buf_2 fanout538 (.A(_1463_),
    .X(net538));
 sg13g2_buf_2 fanout539 (.A(_1463_),
    .X(net539));
 sg13g2_buf_2 fanout540 (.A(net541),
    .X(net540));
 sg13g2_buf_2 fanout541 (.A(_1396_),
    .X(net541));
 sg13g2_buf_2 fanout542 (.A(net543),
    .X(net542));
 sg13g2_buf_2 fanout543 (.A(_1371_),
    .X(net543));
 sg13g2_buf_2 fanout544 (.A(net545),
    .X(net544));
 sg13g2_buf_2 fanout545 (.A(_1319_),
    .X(net545));
 sg13g2_buf_2 fanout546 (.A(net547),
    .X(net546));
 sg13g2_buf_2 fanout547 (.A(_0731_),
    .X(net547));
 sg13g2_buf_2 fanout548 (.A(_0673_),
    .X(net548));
 sg13g2_buf_2 fanout549 (.A(_0673_),
    .X(net549));
 sg13g2_buf_2 fanout550 (.A(_1510_),
    .X(net550));
 sg13g2_buf_2 fanout551 (.A(_1510_),
    .X(net551));
 sg13g2_buf_2 fanout552 (.A(net553),
    .X(net552));
 sg13g2_buf_2 fanout553 (.A(_1464_),
    .X(net553));
 sg13g2_buf_2 fanout554 (.A(net555),
    .X(net554));
 sg13g2_buf_2 fanout555 (.A(_1397_),
    .X(net555));
 sg13g2_buf_2 fanout556 (.A(net557),
    .X(net556));
 sg13g2_buf_2 fanout557 (.A(_1372_),
    .X(net557));
 sg13g2_buf_2 fanout558 (.A(net559),
    .X(net558));
 sg13g2_buf_2 fanout559 (.A(_1320_),
    .X(net559));
 sg13g2_buf_2 fanout560 (.A(net561),
    .X(net560));
 sg13g2_buf_2 fanout561 (.A(_0732_),
    .X(net561));
 sg13g2_buf_2 fanout562 (.A(net564),
    .X(net562));
 sg13g2_buf_2 fanout563 (.A(net564),
    .X(net563));
 sg13g2_buf_2 fanout564 (.A(net565),
    .X(net564));
 sg13g2_buf_2 fanout565 (.A(net578),
    .X(net565));
 sg13g2_buf_2 fanout566 (.A(net567),
    .X(net566));
 sg13g2_buf_2 fanout567 (.A(net568),
    .X(net567));
 sg13g2_buf_2 fanout568 (.A(net569),
    .X(net568));
 sg13g2_buf_4 fanout569 (.X(net569),
    .A(net578));
 sg13g2_buf_2 fanout570 (.A(net571),
    .X(net570));
 sg13g2_buf_2 fanout571 (.A(net575),
    .X(net571));
 sg13g2_buf_2 fanout572 (.A(net574),
    .X(net572));
 sg13g2_buf_1 fanout573 (.A(net574),
    .X(net573));
 sg13g2_buf_1 fanout574 (.A(net575),
    .X(net574));
 sg13g2_buf_4 fanout575 (.X(net575),
    .A(net578));
 sg13g2_buf_2 fanout576 (.A(net577),
    .X(net576));
 sg13g2_buf_1 fanout577 (.A(net578),
    .X(net577));
 sg13g2_buf_8 fanout578 (.A(_0698_),
    .X(net578));
 sg13g2_buf_2 fanout579 (.A(_0674_),
    .X(net579));
 sg13g2_buf_2 fanout580 (.A(_0674_),
    .X(net580));
 sg13g2_buf_4 fanout581 (.X(net581),
    .A(_0635_));
 sg13g2_buf_2 fanout582 (.A(_0635_),
    .X(net582));
 sg13g2_buf_4 fanout583 (.X(net583),
    .A(net586));
 sg13g2_buf_2 fanout584 (.A(net586),
    .X(net584));
 sg13g2_buf_2 fanout585 (.A(net586),
    .X(net585));
 sg13g2_buf_2 fanout586 (.A(net305),
    .X(net586));
 sg13g2_buf_2 fanout587 (.A(\system_integrator_b_counter.value_output[0] ),
    .X(net587));
 sg13g2_buf_2 fanout588 (.A(net489),
    .X(net588));
 sg13g2_buf_2 fanout589 (.A(net504),
    .X(net589));
 sg13g2_buf_4 fanout590 (.X(net590),
    .A(net498));
 sg13g2_buf_2 fanout591 (.A(net482),
    .X(net591));
 sg13g2_buf_4 fanout592 (.X(net592),
    .A(\test_integrator_b_counter.value_output[1] ));
 sg13g2_buf_4 fanout593 (.X(net593),
    .A(net439));
 sg13g2_buf_4 fanout594 (.X(net594),
    .A(net439));
 sg13g2_buf_4 fanout595 (.X(net595),
    .A(net403));
 sg13g2_buf_4 fanout596 (.X(net596),
    .A(\integrator_b_sng_comparator.bits_b[7] ));
 sg13g2_buf_2 fanout597 (.A(net206),
    .X(net597));
 sg13g2_buf_2 fanout598 (.A(\input_a_sng_comparator.bits_b[5] ),
    .X(net598));
 sg13g2_buf_2 fanout599 (.A(net600),
    .X(net599));
 sg13g2_buf_2 fanout600 (.A(net451),
    .X(net600));
 sg13g2_buf_4 fanout601 (.X(net601),
    .A(\input_a_sng_comparator.bits_b[3] ));
 sg13g2_buf_4 fanout602 (.X(net602),
    .A(\input_a_sng_comparator.bits_b[2] ));
 sg13g2_buf_4 fanout603 (.X(net603),
    .A(\input_a_sng_comparator.bits_b[1] ));
 sg13g2_buf_2 fanout604 (.A(net609),
    .X(net604));
 sg13g2_buf_1 fanout605 (.A(net609),
    .X(net605));
 sg13g2_buf_2 fanout606 (.A(net608),
    .X(net606));
 sg13g2_buf_2 fanout607 (.A(net608),
    .X(net607));
 sg13g2_buf_2 fanout608 (.A(net609),
    .X(net608));
 sg13g2_buf_1 fanout609 (.A(net627),
    .X(net609));
 sg13g2_buf_2 fanout610 (.A(net611),
    .X(net610));
 sg13g2_buf_2 fanout611 (.A(net614),
    .X(net611));
 sg13g2_buf_2 fanout612 (.A(net614),
    .X(net612));
 sg13g2_buf_2 fanout613 (.A(net614),
    .X(net613));
 sg13g2_buf_1 fanout614 (.A(net627),
    .X(net614));
 sg13g2_buf_2 fanout615 (.A(net618),
    .X(net615));
 sg13g2_buf_2 fanout616 (.A(net618),
    .X(net616));
 sg13g2_buf_2 fanout617 (.A(net618),
    .X(net617));
 sg13g2_buf_2 fanout618 (.A(net627),
    .X(net618));
 sg13g2_buf_2 fanout619 (.A(net621),
    .X(net619));
 sg13g2_buf_1 fanout620 (.A(net621),
    .X(net620));
 sg13g2_buf_2 fanout621 (.A(net627),
    .X(net621));
 sg13g2_buf_4 fanout622 (.X(net622),
    .A(net626));
 sg13g2_buf_2 fanout623 (.A(net625),
    .X(net623));
 sg13g2_buf_2 fanout624 (.A(net625),
    .X(net624));
 sg13g2_buf_2 fanout625 (.A(net626),
    .X(net625));
 sg13g2_buf_2 fanout626 (.A(net627),
    .X(net626));
 sg13g2_buf_4 fanout627 (.X(net627),
    .A(rst_n));
 sg13g2_buf_2 fanout628 (.A(net630),
    .X(net628));
 sg13g2_buf_2 fanout629 (.A(net630),
    .X(net629));
 sg13g2_buf_2 fanout630 (.A(net641),
    .X(net630));
 sg13g2_buf_2 fanout631 (.A(net632),
    .X(net631));
 sg13g2_buf_2 fanout632 (.A(net641),
    .X(net632));
 sg13g2_buf_2 fanout633 (.A(net634),
    .X(net633));
 sg13g2_buf_2 fanout634 (.A(net636),
    .X(net634));
 sg13g2_buf_2 fanout635 (.A(net636),
    .X(net635));
 sg13g2_buf_1 fanout636 (.A(net641),
    .X(net636));
 sg13g2_buf_2 fanout637 (.A(net640),
    .X(net637));
 sg13g2_buf_2 fanout638 (.A(net640),
    .X(net638));
 sg13g2_buf_2 fanout639 (.A(net640),
    .X(net639));
 sg13g2_buf_2 fanout640 (.A(net641),
    .X(net640));
 sg13g2_buf_2 fanout641 (.A(rst_n),
    .X(net641));
 sg13g2_buf_2 fanout642 (.A(net645),
    .X(net642));
 sg13g2_buf_2 fanout643 (.A(net645),
    .X(net643));
 sg13g2_buf_1 fanout644 (.A(net645),
    .X(net644));
 sg13g2_buf_2 fanout645 (.A(net658),
    .X(net645));
 sg13g2_buf_2 fanout646 (.A(net649),
    .X(net646));
 sg13g2_buf_2 fanout647 (.A(net648),
    .X(net647));
 sg13g2_buf_2 fanout648 (.A(net649),
    .X(net648));
 sg13g2_buf_2 fanout649 (.A(net658),
    .X(net649));
 sg13g2_buf_2 fanout650 (.A(net653),
    .X(net650));
 sg13g2_buf_4 fanout651 (.X(net651),
    .A(net653));
 sg13g2_buf_2 fanout652 (.A(net653),
    .X(net652));
 sg13g2_buf_1 fanout653 (.A(net658),
    .X(net653));
 sg13g2_buf_2 fanout654 (.A(net657),
    .X(net654));
 sg13g2_buf_2 fanout655 (.A(net657),
    .X(net655));
 sg13g2_buf_2 fanout656 (.A(net657),
    .X(net656));
 sg13g2_buf_2 fanout657 (.A(net658),
    .X(net657));
 sg13g2_buf_2 fanout658 (.A(rst_n),
    .X(net658));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_tielo tt_um_stochastic_integrator_tt9_CL123abc_3 (.L_LO(net3));
 sg13g2_buf_2 clkbuf_leaf_1_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_2 clkbuf_leaf_2_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_2 clkbuf_leaf_3_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_2 clkbuf_leaf_4_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_2 clkbuf_leaf_5_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_2 clkbuf_leaf_6_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_2 clkbuf_leaf_7_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_2 clkbuf_leaf_8_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_2 clkbuf_leaf_9_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_2 clkbuf_leaf_10_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_2 clkbuf_leaf_11_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_2 clkbuf_leaf_12_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_2 clkbuf_leaf_13_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_2 clkbuf_leaf_14_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_2 clkbuf_leaf_15_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_2 clkbuf_leaf_16_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_2 clkbuf_leaf_17_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_2 clkbuf_leaf_18_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_2 clkbuf_leaf_19_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_2 clkbuf_leaf_20_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_2 clkbuf_leaf_21_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_2 clkbuf_leaf_22_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_2 clkbuf_leaf_23_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_2 clkbuf_leaf_24_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_2 clkbuf_leaf_25_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_2 clkbuf_leaf_26_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_2 clkbuf_leaf_27_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_2 clkbuf_leaf_28_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_2 clkbuf_leaf_29_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_2 clkbuf_leaf_30_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_2 clkbuf_leaf_31_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_31_clk));
 sg13g2_buf_2 clkbuf_leaf_32_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_32_clk));
 sg13g2_buf_2 clkbuf_leaf_33_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_33_clk));
 sg13g2_buf_2 clkbuf_leaf_34_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_34_clk));
 sg13g2_buf_2 clkbuf_leaf_35_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_35_clk));
 sg13g2_buf_2 clkbuf_leaf_36_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_36_clk));
 sg13g2_buf_2 clkbuf_leaf_37_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_37_clk));
 sg13g2_buf_2 clkbuf_leaf_38_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_38_clk));
 sg13g2_buf_2 clkbuf_leaf_39_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_39_clk));
 sg13g2_buf_2 clkbuf_leaf_40_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_40_clk));
 sg13g2_buf_2 clkbuf_leaf_41_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_41_clk));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_2 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sg13g2_buf_2 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sg13g2_buf_2 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sg13g2_buf_2 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sg13g2_buf_2 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sg13g2_buf_2 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sg13g2_buf_2 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sg13g2_buf_2 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sg13g2_buf_2 clkload0 (.A(clknet_3_1__leaf_clk));
 sg13g2_buf_2 clkload1 (.A(clknet_3_2__leaf_clk));
 sg13g2_buf_2 clkload2 (.A(clknet_3_3__leaf_clk));
 sg13g2_buf_2 clkload3 (.A(clknet_3_5__leaf_clk));
 sg13g2_buf_2 clkload4 (.A(clknet_3_6__leaf_clk));
 sg13g2_buf_2 clkload5 (.A(clknet_3_7__leaf_clk));
 sg13g2_inv_4 clkload6 (.A(clknet_leaf_41_clk));
 sg13g2_inv_1 clkload7 (.A(clknet_leaf_1_clk));
 sg13g2_inv_4 clkload8 (.A(clknet_leaf_4_clk));
 sg13g2_inv_2 clkload9 (.A(clknet_leaf_36_clk));
 sg13g2_inv_1 clkload10 (.A(clknet_leaf_32_clk));
 sg13g2_inv_4 clkload11 (.A(clknet_leaf_27_clk));
 sg13g2_inv_2 clkload12 (.A(clknet_leaf_28_clk));
 sg13g2_inv_4 clkload13 (.A(clknet_leaf_5_clk));
 sg13g2_inv_1 clkload14 (.A(clknet_leaf_11_clk));
 sg13g2_inv_1 clkload15 (.A(clknet_leaf_14_clk));
 sg13g2_inv_1 clkload16 (.A(clknet_leaf_9_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(_1904_),
    .X(net20));
 sg13g2_dlygate4sd3_1 hold2 (.A(_1903_),
    .X(net21));
 sg13g2_dlygate4sd3_1 hold3 (.A(_1905_),
    .X(net22));
 sg13g2_dlygate4sd3_1 hold4 (.A(_1657_),
    .X(net23));
 sg13g2_dlygate4sd3_1 hold5 (.A(_1898_),
    .X(net24));
 sg13g2_dlygate4sd3_1 hold6 (.A(\input_halfprob1_sng_comparator.bits_b[7] ),
    .X(net25));
 sg13g2_dlygate4sd3_1 hold7 (.A(\input_halfprob1_sng_comparator.bits_b[6] ),
    .X(net26));
 sg13g2_dlygate4sd3_1 hold8 (.A(\input_b_sng_comparator.bits_b[1] ),
    .X(net27));
 sg13g2_dlygate4sd3_1 hold9 (.A(\input_a_sng_comparator.bits_b[1] ),
    .X(net28));
 sg13g2_dlygate4sd3_1 hold10 (.A(\integrator_b_sng_comparator.bits_b[7] ),
    .X(net29));
 sg13g2_dlygate4sd3_1 hold11 (.A(\input_halfprob2_sng_comparator.bits_b[6] ),
    .X(net30));
 sg13g2_dlygate4sd3_1 hold12 (.A(\input_halfprob1_sng_comparator.bits_b[8] ),
    .X(net31));
 sg13g2_dlygate4sd3_1 hold13 (.A(\integrator_c_sng_comparator.bits_b[0] ),
    .X(net32));
 sg13g2_dlygate4sd3_1 hold14 (.A(\input_a_sng_comparator.bits_b[8] ),
    .X(net33));
 sg13g2_dlygate4sd3_1 hold15 (.A(\integrator_c_sng_comparator.bits_b[3] ),
    .X(net34));
 sg13g2_dlygate4sd3_1 hold16 (.A(\input_b_sng_comparator.bits_b[2] ),
    .X(net35));
 sg13g2_dlygate4sd3_1 hold17 (.A(\input_halfprob2_sng_comparator.bits_b[7] ),
    .X(net36));
 sg13g2_dlygate4sd3_1 hold18 (.A(\input_a_sng_comparator.bits_b[2] ),
    .X(net37));
 sg13g2_dlygate4sd3_1 hold19 (.A(\input_halfprob2_sng_comparator.bits_b[3] ),
    .X(net38));
 sg13g2_dlygate4sd3_1 hold20 (.A(\system_integrator_b_output.input_bits[8] ),
    .X(net39));
 sg13g2_dlygate4sd3_1 hold21 (.A(_1321_),
    .X(net40));
 sg13g2_dlygate4sd3_1 hold22 (.A(\input_halfprob2_sng_comparator.bits_b[4] ),
    .X(net41));
 sg13g2_dlygate4sd3_1 hold23 (.A(\input_halfprob2_sng_comparator.bits_b[1] ),
    .X(net42));
 sg13g2_dlygate4sd3_1 hold24 (.A(\integrator_b_output.input_bits[8] ),
    .X(net43));
 sg13g2_dlygate4sd3_1 hold25 (.A(_0675_),
    .X(net44));
 sg13g2_dlygate4sd3_1 hold26 (.A(_0074_),
    .X(net45));
 sg13g2_dlygate4sd3_1 hold27 (.A(_0491_),
    .X(net46));
 sg13g2_dlygate4sd3_1 hold28 (.A(_0072_),
    .X(net47));
 sg13g2_dlygate4sd3_1 hold29 (.A(_0509_),
    .X(net48));
 sg13g2_dlygate4sd3_1 hold30 (.A(\test_integrator_a_output.input_bits[0] ),
    .X(net49));
 sg13g2_dlygate4sd3_1 hold31 (.A(_1579_),
    .X(net50));
 sg13g2_dlygate4sd3_1 hold32 (.A(_1934_),
    .X(net51));
 sg13g2_dlygate4sd3_1 hold33 (.A(\system_integrator_a_output.input_bits[8] ),
    .X(net52));
 sg13g2_dlygate4sd3_1 hold34 (.A(_1373_),
    .X(net53));
 sg13g2_dlygate4sd3_1 hold35 (.A(\integrator_a_output.input_bits[8] ),
    .X(net54));
 sg13g2_dlygate4sd3_1 hold36 (.A(_1511_),
    .X(net55));
 sg13g2_dlygate4sd3_1 hold37 (.A(\input_halfprob1_sng_comparator.bits_b[1] ),
    .X(net56));
 sg13g2_dlygate4sd3_1 hold38 (.A(_0073_),
    .X(net57));
 sg13g2_dlygate4sd3_1 hold39 (.A(_0500_),
    .X(net58));
 sg13g2_dlygate4sd3_1 hold40 (.A(\serial_input.output_bitcounter_1[0] ),
    .X(net59));
 sg13g2_dlygate4sd3_1 hold41 (.A(_0607_),
    .X(net60));
 sg13g2_dlygate4sd3_1 hold42 (.A(\test_integrator_b_output.bitseq[6] ),
    .X(net61));
 sg13g2_dlygate4sd3_1 hold43 (.A(_0463_),
    .X(net62));
 sg13g2_dlygate4sd3_1 hold44 (.A(\integrator_c_output.bitseq[5] ),
    .X(net63));
 sg13g2_dlygate4sd3_1 hold45 (.A(_0446_),
    .X(net64));
 sg13g2_dlygate4sd3_1 hold46 (.A(\integrator_c_output.bitseq[0] ),
    .X(net65));
 sg13g2_dlygate4sd3_1 hold47 (.A(_0441_),
    .X(net66));
 sg13g2_dlygate4sd3_1 hold48 (.A(\test_integrator_a_output.bitseq[3] ),
    .X(net67));
 sg13g2_dlygate4sd3_1 hold49 (.A(_0548_),
    .X(net68));
 sg13g2_dlygate4sd3_1 hold50 (.A(\system_integrator_b_output.bitseq[6] ),
    .X(net69));
 sg13g2_dlygate4sd3_1 hold51 (.A(_0480_),
    .X(net70));
 sg13g2_dlygate4sd3_1 hold52 (.A(\system_integrator_a_output.bitseq[1] ),
    .X(net71));
 sg13g2_dlygate4sd3_1 hold53 (.A(_0466_),
    .X(net72));
 sg13g2_dlygate4sd3_1 hold54 (.A(\test_integrator_b_output.input_bits[8] ),
    .X(net73));
 sg13g2_dlygate4sd3_1 hold55 (.A(_1398_),
    .X(net74));
 sg13g2_dlygate4sd3_1 hold56 (.A(\system_integrator_a_output.bitseq[5] ),
    .X(net75));
 sg13g2_dlygate4sd3_1 hold57 (.A(_0470_),
    .X(net76));
 sg13g2_dlygate4sd3_1 hold58 (.A(\system_integrator_a_output.bitseq[0] ),
    .X(net77));
 sg13g2_dlygate4sd3_1 hold59 (.A(_1392_),
    .X(net78));
 sg13g2_dlygate4sd3_1 hold60 (.A(_0465_),
    .X(net79));
 sg13g2_dlygate4sd3_1 hold61 (.A(\integrator_b_output.bitseq[5] ),
    .X(net80));
 sg13g2_dlygate4sd3_1 hold62 (.A(_0621_),
    .X(net81));
 sg13g2_dlygate4sd3_1 hold63 (.A(\test_integrator_b_output.bitseq[3] ),
    .X(net82));
 sg13g2_dlygate4sd3_1 hold64 (.A(_0460_),
    .X(net83));
 sg13g2_dlygate4sd3_1 hold65 (.A(\input_halfprob2_sng_comparator.bits_b[2] ),
    .X(net84));
 sg13g2_dlygate4sd3_1 hold66 (.A(\integrator_b_output.bitseq[2] ),
    .X(net85));
 sg13g2_dlygate4sd3_1 hold67 (.A(_0688_),
    .X(net86));
 sg13g2_dlygate4sd3_1 hold68 (.A(_0618_),
    .X(net87));
 sg13g2_dlygate4sd3_1 hold69 (.A(\test_integrator_a_output.bitseq[2] ),
    .X(net88));
 sg13g2_dlygate4sd3_1 hold70 (.A(_0746_),
    .X(net89));
 sg13g2_dlygate4sd3_1 hold71 (.A(_0547_),
    .X(net90));
 sg13g2_dlygate4sd3_1 hold72 (.A(\integrator_a_output.bitseq[5] ),
    .X(net91));
 sg13g2_dlygate4sd3_1 hold73 (.A(_0433_),
    .X(net92));
 sg13g2_dlygate4sd3_1 hold74 (.A(\system_integrator_a_output.bitseq[4] ),
    .X(net93));
 sg13g2_dlygate4sd3_1 hold75 (.A(_0469_),
    .X(net94));
 sg13g2_dlygate4sd3_1 hold76 (.A(\clk_counter[13] ),
    .X(net95));
 sg13g2_dlygate4sd3_1 hold77 (.A(_1609_),
    .X(net96));
 sg13g2_dlygate4sd3_1 hold78 (.A(_0058_),
    .X(net97));
 sg13g2_dlygate4sd3_1 hold79 (.A(\integrator_a_output.bitseq[0] ),
    .X(net98));
 sg13g2_dlygate4sd3_1 hold80 (.A(_0428_),
    .X(net99));
 sg13g2_dlygate4sd3_1 hold81 (.A(\integrator_c_output.bitseq[1] ),
    .X(net100));
 sg13g2_dlygate4sd3_1 hold82 (.A(_0442_),
    .X(net101));
 sg13g2_dlygate4sd3_1 hold83 (.A(_0030_),
    .X(net102));
 sg13g2_dlygate4sd3_1 hold84 (.A(_0518_),
    .X(net103));
 sg13g2_dlygate4sd3_1 hold85 (.A(\system_integrator_b_output.bitseq[0] ),
    .X(net104));
 sg13g2_dlygate4sd3_1 hold86 (.A(_0474_),
    .X(net105));
 sg13g2_dlygate4sd3_1 hold87 (.A(\system_integrator_a_output.bitseq[6] ),
    .X(net106));
 sg13g2_dlygate4sd3_1 hold88 (.A(_0471_),
    .X(net107));
 sg13g2_dlygate4sd3_1 hold89 (.A(\integrator_b_output.bitseq[4] ),
    .X(net108));
 sg13g2_dlygate4sd3_1 hold90 (.A(_0620_),
    .X(net109));
 sg13g2_dlygate4sd3_1 hold91 (.A(\integrator_a_output.bitseq[1] ),
    .X(net110));
 sg13g2_dlygate4sd3_1 hold92 (.A(_0429_),
    .X(net111));
 sg13g2_dlygate4sd3_1 hold93 (.A(\system_integrator_b_output.bitseq[3] ),
    .X(net112));
 sg13g2_dlygate4sd3_1 hold94 (.A(_0477_),
    .X(net113));
 sg13g2_dlygate4sd3_1 hold95 (.A(\integrator_b_output.bitseq[3] ),
    .X(net114));
 sg13g2_dlygate4sd3_1 hold96 (.A(_0619_),
    .X(net115));
 sg13g2_dlygate4sd3_1 hold97 (.A(\integrator_b_output.bitseq[6] ),
    .X(net116));
 sg13g2_dlygate4sd3_1 hold98 (.A(_0622_),
    .X(net117));
 sg13g2_dlygate4sd3_1 hold99 (.A(\integrator_b_output.input_bits[7] ),
    .X(net118));
 sg13g2_dlygate4sd3_1 hold100 (.A(_0569_),
    .X(net119));
 sg13g2_dlygate4sd3_1 hold101 (.A(\serial_input.output_bitcounter_1[1] ),
    .X(net120));
 sg13g2_dlygate4sd3_1 hold102 (.A(_0608_),
    .X(net121));
 sg13g2_dlygate4sd3_1 hold103 (.A(\test_integrator_b_output.bitseq[5] ),
    .X(net122));
 sg13g2_dlygate4sd3_1 hold104 (.A(_0462_),
    .X(net123));
 sg13g2_dlygate4sd3_1 hold105 (.A(\test_integrator_b_output.bitseq[0] ),
    .X(net124));
 sg13g2_dlygate4sd3_1 hold106 (.A(_0457_),
    .X(net125));
 sg13g2_dlygate4sd3_1 hold107 (.A(\system_integrator_b_output.bitseq[5] ),
    .X(net126));
 sg13g2_dlygate4sd3_1 hold108 (.A(_0479_),
    .X(net127));
 sg13g2_dlygate4sd3_1 hold109 (.A(\integrator_b_output.bitseq[1] ),
    .X(net128));
 sg13g2_dlygate4sd3_1 hold110 (.A(_0617_),
    .X(net129));
 sg13g2_dlygate4sd3_1 hold111 (.A(\test_integrator_a_output.bitseq[5] ),
    .X(net130));
 sg13g2_dlygate4sd3_1 hold112 (.A(_0550_),
    .X(net131));
 sg13g2_dlygate4sd3_1 hold113 (.A(\integrator_b_output.input_bits[6] ),
    .X(net132));
 sg13g2_dlygate4sd3_1 hold114 (.A(_0568_),
    .X(net133));
 sg13g2_dlygate4sd3_1 hold115 (.A(\input_halfprob1_sng_comparator.bits_b[0] ),
    .X(net134));
 sg13g2_dlygate4sd3_1 hold116 (.A(\integrator_a_output.bitseq[4] ),
    .X(net135));
 sg13g2_dlygate4sd3_1 hold117 (.A(_0432_),
    .X(net136));
 sg13g2_dlygate4sd3_1 hold118 (.A(\integrator_c_output.bitseq[6] ),
    .X(net137));
 sg13g2_dlygate4sd3_1 hold119 (.A(_0447_),
    .X(net138));
 sg13g2_dlygate4sd3_1 hold120 (.A(\test_integrator_b_output.bitseq[1] ),
    .X(net139));
 sg13g2_dlygate4sd3_1 hold121 (.A(_0458_),
    .X(net140));
 sg13g2_dlygate4sd3_1 hold122 (.A(_0085_),
    .X(net141));
 sg13g2_dlygate4sd3_1 hold123 (.A(_0439_),
    .X(net142));
 sg13g2_dlygate4sd3_1 hold124 (.A(\system_integrator_b_output.bitseq[1] ),
    .X(net143));
 sg13g2_dlygate4sd3_1 hold125 (.A(_1337_),
    .X(net144));
 sg13g2_dlygate4sd3_1 hold126 (.A(_0475_),
    .X(net145));
 sg13g2_dlygate4sd3_1 hold127 (.A(\integrator_b_output.input_bits[1] ),
    .X(net146));
 sg13g2_dlygate4sd3_1 hold128 (.A(_0563_),
    .X(net147));
 sg13g2_dlygate4sd3_1 hold129 (.A(\system_integrator_a_output.bitseq[2] ),
    .X(net148));
 sg13g2_dlygate4sd3_1 hold130 (.A(_0467_),
    .X(net149));
 sg13g2_dlygate4sd3_1 hold131 (.A(\test_integrator_a_output.bitseq[4] ),
    .X(net150));
 sg13g2_dlygate4sd3_1 hold132 (.A(_0549_),
    .X(net151));
 sg13g2_dlygate4sd3_1 hold133 (.A(\integrator_c_output.bitseq[3] ),
    .X(net152));
 sg13g2_dlygate4sd3_1 hold134 (.A(_0444_),
    .X(net153));
 sg13g2_dlygate4sd3_1 hold135 (.A(\test_integrator_a_output.bitseq[1] ),
    .X(net154));
 sg13g2_dlygate4sd3_1 hold136 (.A(_0546_),
    .X(net155));
 sg13g2_dlygate4sd3_1 hold137 (.A(\integrator_a_output.input_bits[4] ),
    .X(net156));
 sg13g2_dlygate4sd3_1 hold138 (.A(_0557_),
    .X(net157));
 sg13g2_dlygate4sd3_1 hold139 (.A(\test_integrator_b_output.bitseq[2] ),
    .X(net158));
 sg13g2_dlygate4sd3_1 hold140 (.A(_0459_),
    .X(net159));
 sg13g2_dlygate4sd3_1 hold141 (.A(\system_integrator_b_output.bitseq[2] ),
    .X(net160));
 sg13g2_dlygate4sd3_1 hold142 (.A(_1334_),
    .X(net161));
 sg13g2_dlygate4sd3_1 hold143 (.A(_0476_),
    .X(net162));
 sg13g2_dlygate4sd3_1 hold144 (.A(\integrator_c_output.bitseq[2] ),
    .X(net163));
 sg13g2_dlygate4sd3_1 hold145 (.A(_0443_),
    .X(net164));
 sg13g2_dlygate4sd3_1 hold146 (.A(\integrator_c_output.input_bits[8] ),
    .X(net165));
 sg13g2_dlygate4sd3_1 hold147 (.A(_1465_),
    .X(net166));
 sg13g2_dlygate4sd3_1 hold148 (.A(\integrator_c_output.input_bits[2] ),
    .X(net167));
 sg13g2_dlygate4sd3_1 hold149 (.A(_0573_),
    .X(net168));
 sg13g2_dlygate4sd3_1 hold150 (.A(\system_integrator_a_output.bitseq[3] ),
    .X(net169));
 sg13g2_dlygate4sd3_1 hold151 (.A(_0468_),
    .X(net170));
 sg13g2_dlygate4sd3_1 hold152 (.A(\integrator_a_output.bitseq[3] ),
    .X(net171));
 sg13g2_dlygate4sd3_1 hold153 (.A(\integrator_c_output.input_bits[0] ),
    .X(net172));
 sg13g2_dlygate4sd3_1 hold154 (.A(_1931_),
    .X(net173));
 sg13g2_dlygate4sd3_1 hold155 (.A(\test_integrator_b_output.input_bits[0] ),
    .X(net174));
 sg13g2_dlygate4sd3_1 hold156 (.A(_0482_),
    .X(net175));
 sg13g2_dlygate4sd3_1 hold157 (.A(\integrator_b_output.bitseq[0] ),
    .X(net176));
 sg13g2_dlygate4sd3_1 hold158 (.A(\test_integrator_b_output.input_bits[1] ),
    .X(net177));
 sg13g2_dlygate4sd3_1 hold159 (.A(_0483_),
    .X(net178));
 sg13g2_dlygate4sd3_1 hold160 (.A(\integrator_b_output.input_bits[4] ),
    .X(net179));
 sg13g2_dlygate4sd3_1 hold161 (.A(_0725_),
    .X(net180));
 sg13g2_dlygate4sd3_1 hold162 (.A(_0566_),
    .X(net181));
 sg13g2_dlygate4sd3_1 hold163 (.A(\integrator_b_output.input_bits[5] ),
    .X(net182));
 sg13g2_dlygate4sd3_1 hold164 (.A(_0567_),
    .X(net183));
 sg13g2_dlygate4sd3_1 hold165 (.A(\test_integrator_b_output.bitseq[4] ),
    .X(net184));
 sg13g2_dlygate4sd3_1 hold166 (.A(_0461_),
    .X(net185));
 sg13g2_dlygate4sd3_1 hold167 (.A(\integrator_a_output.bitseq[6] ),
    .X(net186));
 sg13g2_dlygate4sd3_1 hold168 (.A(_1512_),
    .X(net187));
 sg13g2_dlygate4sd3_1 hold169 (.A(_0434_),
    .X(net188));
 sg13g2_dlygate4sd3_1 hold170 (.A(\test_integrator_b_counter.value_output[8] ),
    .X(net189));
 sg13g2_dlygate4sd3_1 hold171 (.A(\integrator_c_output.bitseq[4] ),
    .X(net190));
 sg13g2_dlygate4sd3_1 hold172 (.A(_0445_),
    .X(net191));
 sg13g2_dlygate4sd3_1 hold173 (.A(\integrator_b_output.input_bits[3] ),
    .X(net192));
 sg13g2_dlygate4sd3_1 hold174 (.A(_0565_),
    .X(net193));
 sg13g2_dlygate4sd3_1 hold175 (.A(\integrator_a_output.input_bits[6] ),
    .X(net194));
 sg13g2_dlygate4sd3_1 hold176 (.A(_0559_),
    .X(net195));
 sg13g2_dlygate4sd3_1 hold177 (.A(\integrator_a_output.input_bits[2] ),
    .X(net196));
 sg13g2_dlygate4sd3_1 hold178 (.A(_0555_),
    .X(net197));
 sg13g2_dlygate4sd3_1 hold179 (.A(\integrator_b_output.input_bits[2] ),
    .X(net198));
 sg13g2_dlygate4sd3_1 hold180 (.A(_0564_),
    .X(net199));
 sg13g2_dlygate4sd3_1 hold181 (.A(\system_integrator_a_output.input_bits[2] ),
    .X(net200));
 sg13g2_dlygate4sd3_1 hold182 (.A(_0582_),
    .X(net201));
 sg13g2_dlygate4sd3_1 hold183 (.A(\integrator_a_output.input_bits[1] ),
    .X(net202));
 sg13g2_dlygate4sd3_1 hold184 (.A(_0554_),
    .X(net203));
 sg13g2_dlygate4sd3_1 hold185 (.A(\test_integrator_b_output.input_bits[4] ),
    .X(net204));
 sg13g2_dlygate4sd3_1 hold186 (.A(_0486_),
    .X(net205));
 sg13g2_dlygate4sd3_1 hold187 (.A(\input_a_sng_comparator.bits_b[6] ),
    .X(net206));
 sg13g2_dlygate4sd3_1 hold188 (.A(\system_integrator_a_output.input_bits[5] ),
    .X(net207));
 sg13g2_dlygate4sd3_1 hold189 (.A(_0585_),
    .X(net208));
 sg13g2_dlygate4sd3_1 hold190 (.A(\system_integrator_b_output.bitseq[4] ),
    .X(net209));
 sg13g2_dlygate4sd3_1 hold191 (.A(_0478_),
    .X(net210));
 sg13g2_dlygate4sd3_1 hold192 (.A(\serial_input.output_bitcounter_1[4] ),
    .X(net211));
 sg13g2_dlygate4sd3_1 hold193 (.A(_0418_),
    .X(net212));
 sg13g2_dlygate4sd3_1 hold194 (.A(\serial_input.adjustment[2] ),
    .X(net213));
 sg13g2_dlygate4sd3_1 hold195 (.A(_0438_),
    .X(net214));
 sg13g2_dlygate4sd3_1 hold196 (.A(\system_integrator_a_output.input_bits[7] ),
    .X(net215));
 sg13g2_dlygate4sd3_1 hold197 (.A(_0587_),
    .X(net216));
 sg13g2_dlygate4sd3_1 hold198 (.A(\test_integrator_b_output.input_bits[3] ),
    .X(net217));
 sg13g2_dlygate4sd3_1 hold199 (.A(_0485_),
    .X(net218));
 sg13g2_dlygate4sd3_1 hold200 (.A(\integrator_b_output.input_bits[0] ),
    .X(net219));
 sg13g2_dlygate4sd3_1 hold201 (.A(_0562_),
    .X(net220));
 sg13g2_dlygate4sd3_1 hold202 (.A(\test_integrator_a_output.input_bits[1] ),
    .X(net221));
 sg13g2_dlygate4sd3_1 hold203 (.A(_0599_),
    .X(net222));
 sg13g2_dlygate4sd3_1 hold204 (.A(\test_integrator_b_output.input_bits[5] ),
    .X(net223));
 sg13g2_dlygate4sd3_1 hold205 (.A(_0487_),
    .X(net224));
 sg13g2_dlygate4sd3_1 hold206 (.A(\integrator_a_output.bitseq[2] ),
    .X(net225));
 sg13g2_dlygate4sd3_1 hold207 (.A(_0430_),
    .X(net226));
 sg13g2_dlygate4sd3_1 hold208 (.A(_0084_),
    .X(net227));
 sg13g2_dlygate4sd3_1 hold209 (.A(_0436_),
    .X(net228));
 sg13g2_dlygate4sd3_1 hold210 (.A(\test_integrator_a_output.bitseq[7] ),
    .X(net229));
 sg13g2_dlygate4sd3_1 hold211 (.A(_0733_),
    .X(net230));
 sg13g2_dlygate4sd3_1 hold212 (.A(\integrator_b_counter.value_output[8] ),
    .X(net231));
 sg13g2_dlygate4sd3_1 hold213 (.A(\system_integrator_a_output.input_bits[1] ),
    .X(net232));
 sg13g2_dlygate4sd3_1 hold214 (.A(_0581_),
    .X(net233));
 sg13g2_dlygate4sd3_1 hold215 (.A(\test_integrator_a_counter.value_output[0] ),
    .X(net234));
 sg13g2_dlygate4sd3_1 hold216 (.A(\test_integrator_b_output.input_bits[6] ),
    .X(net235));
 sg13g2_dlygate4sd3_1 hold217 (.A(_0488_),
    .X(net236));
 sg13g2_dlygate4sd3_1 hold218 (.A(\test_integrator_a_output.bitseq[6] ),
    .X(net237));
 sg13g2_dlygate4sd3_1 hold219 (.A(_0551_),
    .X(net238));
 sg13g2_dlygate4sd3_1 hold220 (.A(\system_integrator_a_output.input_bits[0] ),
    .X(net239));
 sg13g2_dlygate4sd3_1 hold221 (.A(_1932_),
    .X(net240));
 sg13g2_dlygate4sd3_1 hold222 (.A(\integrator_b_sng_comparator.bits_b[6] ),
    .X(net241));
 sg13g2_dlygate4sd3_1 hold223 (.A(\input_a_sng_comparator.bits_a[4] ),
    .X(net242));
 sg13g2_dlygate4sd3_1 hold224 (.A(\integrator_a_counter.value_output[8] ),
    .X(net243));
 sg13g2_dlygate4sd3_1 hold225 (.A(\test_integrator_a_output.bitseq[0] ),
    .X(net244));
 sg13g2_dlygate4sd3_1 hold226 (.A(_0545_),
    .X(net245));
 sg13g2_dlygate4sd3_1 hold227 (.A(\system_integrator_a_output.input_bits[3] ),
    .X(net246));
 sg13g2_dlygate4sd3_1 hold228 (.A(_0583_),
    .X(net247));
 sg13g2_dlygate4sd3_1 hold229 (.A(\integrator_a_output.input_bits[5] ),
    .X(net248));
 sg13g2_dlygate4sd3_1 hold230 (.A(_0558_),
    .X(net249));
 sg13g2_dlygate4sd3_1 hold231 (.A(\test_integrator_b_output.input_bits[2] ),
    .X(net250));
 sg13g2_dlygate4sd3_1 hold232 (.A(_0484_),
    .X(net251));
 sg13g2_dlygate4sd3_1 hold233 (.A(\system_integrator_a_counter.value_output[0] ),
    .X(net252));
 sg13g2_dlygate4sd3_1 hold234 (.A(\clk_counter[7] ),
    .X(net253));
 sg13g2_dlygate4sd3_1 hold235 (.A(_0069_),
    .X(net254));
 sg13g2_dlygate4sd3_1 hold236 (.A(\integrator_c_output.input_bits[7] ),
    .X(net255));
 sg13g2_dlygate4sd3_1 hold237 (.A(_0578_),
    .X(net256));
 sg13g2_dlygate4sd3_1 hold238 (.A(\system_integrator_a_counter.value_output[8] ),
    .X(net257));
 sg13g2_dlygate4sd3_1 hold239 (.A(\serial_input.output_bitcounter_2[2] ),
    .X(net258));
 sg13g2_dlygate4sd3_1 hold240 (.A(_0626_),
    .X(net259));
 sg13g2_dlygate4sd3_1 hold241 (.A(\system_integrator_b_output.input_bits[6] ),
    .X(net260));
 sg13g2_dlygate4sd3_1 hold242 (.A(_0595_),
    .X(net261));
 sg13g2_dlygate4sd3_1 hold243 (.A(\integrator_a_output.input_bits[7] ),
    .X(net262));
 sg13g2_dlygate4sd3_1 hold244 (.A(_0560_),
    .X(net263));
 sg13g2_dlygate4sd3_1 hold245 (.A(\test_integrator_a_output.input_bits[7] ),
    .X(net264));
 sg13g2_dlygate4sd3_1 hold246 (.A(_0605_),
    .X(net265));
 sg13g2_dlygate4sd3_1 hold247 (.A(\integrator_c_output.input_bits[1] ),
    .X(net266));
 sg13g2_dlygate4sd3_1 hold248 (.A(_0572_),
    .X(net267));
 sg13g2_dlygate4sd3_1 hold249 (.A(\serial_input.output_bitcounter_2[0] ),
    .X(net268));
 sg13g2_dlygate4sd3_1 hold250 (.A(_0624_),
    .X(net269));
 sg13g2_dlygate4sd3_1 hold251 (.A(\clk_counter[11] ),
    .X(net270));
 sg13g2_dlygate4sd3_1 hold252 (.A(_0056_),
    .X(net271));
 sg13g2_dlygate4sd3_1 hold253 (.A(\system_integrator_b_output.input_bits[5] ),
    .X(net272));
 sg13g2_dlygate4sd3_1 hold254 (.A(_0594_),
    .X(net273));
 sg13g2_dlygate4sd3_1 hold255 (.A(\integrator_a_output.input_bits[3] ),
    .X(net274));
 sg13g2_dlygate4sd3_1 hold256 (.A(_0556_),
    .X(net275));
 sg13g2_dlygate4sd3_1 hold257 (.A(\system_integrator_a_output.input_bits[4] ),
    .X(net276));
 sg13g2_dlygate4sd3_1 hold258 (.A(_0584_),
    .X(net277));
 sg13g2_dlygate4sd3_1 hold259 (.A(\integrator_c_output.input_bits[3] ),
    .X(net278));
 sg13g2_dlygate4sd3_1 hold260 (.A(_0574_),
    .X(net279));
 sg13g2_dlygate4sd3_1 hold261 (.A(\system_integrator_b_output.input_bits[7] ),
    .X(net280));
 sg13g2_dlygate4sd3_1 hold262 (.A(_0596_),
    .X(net281));
 sg13g2_dlygate4sd3_1 hold263 (.A(\test_integrator_a_output.input_bits[2] ),
    .X(net282));
 sg13g2_dlygate4sd3_1 hold264 (.A(_0600_),
    .X(net283));
 sg13g2_dlygate4sd3_1 hold265 (.A(\serial_input.output_bitcounter_2[1] ),
    .X(net284));
 sg13g2_dlygate4sd3_1 hold266 (.A(_0625_),
    .X(net285));
 sg13g2_dlygate4sd3_1 hold267 (.A(\system_integrator_b_output.input_bits[0] ),
    .X(net286));
 sg13g2_dlygate4sd3_1 hold268 (.A(_0589_),
    .X(net287));
 sg13g2_dlygate4sd3_1 hold269 (.A(\system_integrator_a_output.input_bits[6] ),
    .X(net288));
 sg13g2_dlygate4sd3_1 hold270 (.A(_0586_),
    .X(net289));
 sg13g2_dlygate4sd3_1 hold271 (.A(\serial_input.output_bitcounter_1[6] ),
    .X(net290));
 sg13g2_dlygate4sd3_1 hold272 (.A(_0420_),
    .X(net291));
 sg13g2_dlygate4sd3_1 hold273 (.A(\system_integrator_b_counter.value_output[8] ),
    .X(net292));
 sg13g2_dlygate4sd3_1 hold274 (.A(\system_integrator_b_output.input_bits[1] ),
    .X(net293));
 sg13g2_dlygate4sd3_1 hold275 (.A(_0590_),
    .X(net294));
 sg13g2_dlygate4sd3_1 hold276 (.A(\test_integrator_a_output.input_bits[6] ),
    .X(net295));
 sg13g2_dlygate4sd3_1 hold277 (.A(_0604_),
    .X(net296));
 sg13g2_dlygate4sd3_1 hold278 (.A(_0037_),
    .X(net297));
 sg13g2_dlygate4sd3_1 hold279 (.A(_1444_),
    .X(net298));
 sg13g2_dlygate4sd3_1 hold280 (.A(_0453_),
    .X(net299));
 sg13g2_dlygate4sd3_1 hold281 (.A(\serial_input.output_bitcounter_1[2] ),
    .X(net300));
 sg13g2_dlygate4sd3_1 hold282 (.A(\clk_counter[6] ),
    .X(net301));
 sg13g2_dlygate4sd3_1 hold283 (.A(_0068_),
    .X(net302));
 sg13g2_dlygate4sd3_1 hold284 (.A(\integrator_c_output.counter[3] ),
    .X(net303));
 sg13g2_dlygate4sd3_1 hold285 (.A(_0011_),
    .X(net304));
 sg13g2_dlygate4sd3_1 hold286 (.A(\serial_input.loop ),
    .X(net305));
 sg13g2_dlygate4sd3_1 hold287 (.A(\clk_counter[17] ),
    .X(net306));
 sg13g2_dlygate4sd3_1 hold288 (.A(_0062_),
    .X(net307));
 sg13g2_dlygate4sd3_1 hold289 (.A(\system_integrator_a_output.counter[3] ),
    .X(net308));
 sg13g2_dlygate4sd3_1 hold290 (.A(_0016_),
    .X(net309));
 sg13g2_dlygate4sd3_1 hold291 (.A(\serial_input.output_bitcounter_1[7] ),
    .X(net310));
 sg13g2_dlygate4sd3_1 hold292 (.A(_0422_),
    .X(net311));
 sg13g2_dlygate4sd3_1 hold293 (.A(\integrator_c_counter.value_output[8] ),
    .X(net312));
 sg13g2_dlygate4sd3_1 hold294 (.A(\serial_input.output_bitcounter_2[4] ),
    .X(net313));
 sg13g2_dlygate4sd3_1 hold295 (.A(_0628_),
    .X(net314));
 sg13g2_dlygate4sd3_1 hold296 (.A(\integrator_c_output.input_bits[5] ),
    .X(net315));
 sg13g2_dlygate4sd3_1 hold297 (.A(_0576_),
    .X(net316));
 sg13g2_dlygate4sd3_1 hold298 (.A(\integrator_a_sng_comparator.bits_b[1] ),
    .X(net317));
 sg13g2_dlygate4sd3_1 hold299 (.A(\test_integrator_b_output.input_bits[7] ),
    .X(net318));
 sg13g2_dlygate4sd3_1 hold300 (.A(_0489_),
    .X(net319));
 sg13g2_dlygate4sd3_1 hold301 (.A(\system_integrator_b_output.counter[3] ),
    .X(net320));
 sg13g2_dlygate4sd3_1 hold302 (.A(_0020_),
    .X(net321));
 sg13g2_dlygate4sd3_1 hold303 (.A(\integrator_c_output.input_bits[6] ),
    .X(net322));
 sg13g2_dlygate4sd3_1 hold304 (.A(_0577_),
    .X(net323));
 sg13g2_dlygate4sd3_1 hold305 (.A(\input_a_sng_comparator.bits_a[6] ),
    .X(net324));
 sg13g2_dlygate4sd3_1 hold306 (.A(\input_b_sng_comparator.bits_a[8] ),
    .X(net325));
 sg13g2_dlygate4sd3_1 hold307 (.A(_0632_),
    .X(net326));
 sg13g2_dlygate4sd3_1 hold308 (.A(\serial_input.output_bitcounter_2[7] ),
    .X(net327));
 sg13g2_dlygate4sd3_1 hold309 (.A(_0412_),
    .X(net328));
 sg13g2_dlygate4sd3_1 hold310 (.A(\test_integrator_a_output.input_bits[4] ),
    .X(net329));
 sg13g2_dlygate4sd3_1 hold311 (.A(_0602_),
    .X(net330));
 sg13g2_dlygate4sd3_1 hold312 (.A(\input_b_sng_comparator.bits_a[7] ),
    .X(net331));
 sg13g2_dlygate4sd3_1 hold313 (.A(\serial_input.output_bitcounter_1[3] ),
    .X(net332));
 sg13g2_dlygate4sd3_1 hold314 (.A(\serial_input.output_bitcounter_1[5] ),
    .X(net333));
 sg13g2_dlygate4sd3_1 hold315 (.A(\system_integrator_b_output.input_bits[4] ),
    .X(net334));
 sg13g2_dlygate4sd3_1 hold316 (.A(_0593_),
    .X(net335));
 sg13g2_dlygate4sd3_1 hold317 (.A(\serial_input.output_bitcounter_2[8] ),
    .X(net336));
 sg13g2_dlygate4sd3_1 hold318 (.A(\integrator_b_output.counter[3] ),
    .X(net337));
 sg13g2_dlygate4sd3_1 hold319 (.A(_0007_),
    .X(net338));
 sg13g2_dlygate4sd3_1 hold320 (.A(\test_integrator_a_output.input_bits[3] ),
    .X(net339));
 sg13g2_dlygate4sd3_1 hold321 (.A(_0601_),
    .X(net340));
 sg13g2_dlygate4sd3_1 hold322 (.A(\integrator_a_output.input_bits[0] ),
    .X(net341));
 sg13g2_dlygate4sd3_1 hold323 (.A(_0553_),
    .X(net342));
 sg13g2_dlygate4sd3_1 hold324 (.A(\system_integrator_b_output.input_bits[2] ),
    .X(net343));
 sg13g2_dlygate4sd3_1 hold325 (.A(_0591_),
    .X(net344));
 sg13g2_dlygate4sd3_1 hold326 (.A(\integrator_c_output.input_bits[4] ),
    .X(net345));
 sg13g2_dlygate4sd3_1 hold327 (.A(_0575_),
    .X(net346));
 sg13g2_dlygate4sd3_1 hold328 (.A(\system_integrator_b_output.counter[0] ),
    .X(net347));
 sg13g2_dlygate4sd3_1 hold329 (.A(\serial_input.output_bitcounter_2[6] ),
    .X(net348));
 sg13g2_dlygate4sd3_1 hold330 (.A(_0630_),
    .X(net349));
 sg13g2_dlygate4sd3_1 hold331 (.A(\input_a_sng_comparator.bits_a[2] ),
    .X(net350));
 sg13g2_dlygate4sd3_1 hold332 (.A(\input_a_sng_comparator.bits_a[5] ),
    .X(net351));
 sg13g2_dlygate4sd3_1 hold333 (.A(\system_integrator_a_output.counter[0] ),
    .X(net352));
 sg13g2_dlygate4sd3_1 hold334 (.A(\system_integrator_b_output.input_bits[3] ),
    .X(net353));
 sg13g2_dlygate4sd3_1 hold335 (.A(_0592_),
    .X(net354));
 sg13g2_dlygate4sd3_1 hold336 (.A(\test_integrator_a_output.counter[0] ),
    .X(net355));
 sg13g2_dlygate4sd3_1 hold337 (.A(\test_integrator_a_output.counter[3] ),
    .X(net356));
 sg13g2_dlygate4sd3_1 hold338 (.A(_0024_),
    .X(net357));
 sg13g2_dlygate4sd3_1 hold339 (.A(\serial_input.output_bitcounter_2[5] ),
    .X(net358));
 sg13g2_dlygate4sd3_1 hold340 (.A(_0629_),
    .X(net359));
 sg13g2_dlygate4sd3_1 hold341 (.A(\serial_input.output_bitcounter_2[3] ),
    .X(net360));
 sg13g2_dlygate4sd3_1 hold342 (.A(\test_integrator_a_output.input_bits[5] ),
    .X(net361));
 sg13g2_dlygate4sd3_1 hold343 (.A(_0603_),
    .X(net362));
 sg13g2_dlygate4sd3_1 hold344 (.A(\integrator_a_output.counter[0] ),
    .X(net363));
 sg13g2_dlygate4sd3_1 hold345 (.A(\integrator_a_output.counter[3] ),
    .X(net364));
 sg13g2_dlygate4sd3_1 hold346 (.A(_0003_),
    .X(net365));
 sg13g2_dlygate4sd3_1 hold347 (.A(\test_integrator_a_output.input_bits[8] ),
    .X(net366));
 sg13g2_dlygate4sd3_1 hold348 (.A(_0606_),
    .X(net367));
 sg13g2_dlygate4sd3_1 hold349 (.A(\clk_counter[10] ),
    .X(net368));
 sg13g2_dlygate4sd3_1 hold350 (.A(_0055_),
    .X(net369));
 sg13g2_dlygate4sd3_1 hold351 (.A(\input_a_sng_comparator.bits_a[3] ),
    .X(net370));
 sg13g2_dlygate4sd3_1 hold352 (.A(\clk_counter[12] ),
    .X(net371));
 sg13g2_dlygate4sd3_1 hold353 (.A(_0038_),
    .X(net372));
 sg13g2_dlygate4sd3_1 hold354 (.A(_0454_),
    .X(net373));
 sg13g2_dlygate4sd3_1 hold355 (.A(_0050_),
    .X(net374));
 sg13g2_dlygate4sd3_1 hold356 (.A(_0544_),
    .X(net375));
 sg13g2_dlygate4sd3_1 hold357 (.A(\serial_input.adjustment[4] ),
    .X(net376));
 sg13g2_dlygate4sd3_1 hold358 (.A(_0440_),
    .X(net377));
 sg13g2_dlygate4sd3_1 hold359 (.A(\clk_counter[8] ),
    .X(net378));
 sg13g2_dlygate4sd3_1 hold360 (.A(_0070_),
    .X(net379));
 sg13g2_dlygate4sd3_1 hold361 (.A(\serial_input.adjustment[1] ),
    .X(net380));
 sg13g2_dlygate4sd3_1 hold362 (.A(_0437_),
    .X(net381));
 sg13g2_dlygate4sd3_1 hold363 (.A(\integrator_c_output.counter[0] ),
    .X(net382));
 sg13g2_dlygate4sd3_1 hold364 (.A(\integrator_b_output.counter[0] ),
    .X(net383));
 sg13g2_dlygate4sd3_1 hold365 (.A(_0039_),
    .X(net384));
 sg13g2_dlygate4sd3_1 hold366 (.A(_0455_),
    .X(net385));
 sg13g2_dlygate4sd3_1 hold367 (.A(\input_b_sng_comparator.bits_a[3] ),
    .X(net386));
 sg13g2_dlygate4sd3_1 hold368 (.A(\integrator_b_counter.value_output[1] ),
    .X(net387));
 sg13g2_dlygate4sd3_1 hold369 (.A(_0501_),
    .X(net388));
 sg13g2_dlygate4sd3_1 hold370 (.A(\serial_input.output_case[2] ),
    .X(net389));
 sg13g2_dlygate4sd3_1 hold371 (.A(_1538_),
    .X(net390));
 sg13g2_dlygate4sd3_1 hold372 (.A(\integrator_c_counter.value_output[0] ),
    .X(net391));
 sg13g2_dlygate4sd3_1 hold373 (.A(\test_integrator_b_output.counter[3] ),
    .X(net392));
 sg13g2_dlygate4sd3_1 hold374 (.A(_0028_),
    .X(net393));
 sg13g2_dlygate4sd3_1 hold375 (.A(\test_integrator_b_output.counter[0] ),
    .X(net394));
 sg13g2_dlygate4sd3_1 hold376 (.A(_0035_),
    .X(net395));
 sg13g2_dlygate4sd3_1 hold377 (.A(_0451_),
    .X(net396));
 sg13g2_dlygate4sd3_1 hold378 (.A(\integrator_a_counter.value_output[1] ),
    .X(net397));
 sg13g2_dlygate4sd3_1 hold379 (.A(_0492_),
    .X(net398));
 sg13g2_dlygate4sd3_1 hold380 (.A(\test_integrator_b_counter.value_output[4] ),
    .X(net399));
 sg13g2_dlygate4sd3_1 hold381 (.A(_0452_),
    .X(net400));
 sg13g2_dlygate4sd3_1 hold382 (.A(\integrator_b_sng_comparator.bits_b[8] ),
    .X(net401));
 sg13g2_dlygate4sd3_1 hold383 (.A(_0053_),
    .X(net402));
 sg13g2_dlygate4sd3_1 hold384 (.A(\input_halfprob2_sng_comparator.bits_b[8] ),
    .X(net403));
 sg13g2_dlygate4sd3_1 hold385 (.A(\serial_input.output_bitcounter_1[8] ),
    .X(net404));
 sg13g2_dlygate4sd3_1 hold386 (.A(_0615_),
    .X(net405));
 sg13g2_dlygate4sd3_1 hold387 (.A(\clk_counter[14] ),
    .X(net406));
 sg13g2_dlygate4sd3_1 hold388 (.A(\integrator_c_counter.value_output[3] ),
    .X(net407));
 sg13g2_dlygate4sd3_1 hold389 (.A(_0512_),
    .X(net408));
 sg13g2_dlygate4sd3_1 hold390 (.A(\input_a_sng_comparator.bits_a[7] ),
    .X(net409));
 sg13g2_dlygate4sd3_1 hold391 (.A(\integrator_c_counter.value_output[5] ),
    .X(net410));
 sg13g2_dlygate4sd3_1 hold392 (.A(_0514_),
    .X(net411));
 sg13g2_dlygate4sd3_1 hold393 (.A(\input_a_sng_comparator.bits_b[0] ),
    .X(net412));
 sg13g2_dlygate4sd3_1 hold394 (.A(\serial_input.output_case[0] ),
    .X(net413));
 sg13g2_dlygate4sd3_1 hold395 (.A(_1540_),
    .X(net414));
 sg13g2_dlygate4sd3_1 hold396 (.A(\integrator_c_counter.value_output[1] ),
    .X(net415));
 sg13g2_dlygate4sd3_1 hold397 (.A(_0510_),
    .X(net416));
 sg13g2_dlygate4sd3_1 hold398 (.A(_0033_),
    .X(net417));
 sg13g2_dlygate4sd3_1 hold399 (.A(_0867_),
    .X(net418));
 sg13g2_dlygate4sd3_1 hold400 (.A(_0537_),
    .X(net419));
 sg13g2_dlygate4sd3_1 hold401 (.A(_0054_),
    .X(net420));
 sg13g2_dlygate4sd3_1 hold402 (.A(\clk_counter[3] ),
    .X(net421));
 sg13g2_dlygate4sd3_1 hold403 (.A(_0065_),
    .X(net422));
 sg13g2_dlygate4sd3_1 hold404 (.A(\clk_counter[1] ),
    .X(net423));
 sg13g2_dlygate4sd3_1 hold405 (.A(_0063_),
    .X(net424));
 sg13g2_dlygate4sd3_1 hold406 (.A(\integrator_b_output.counter[1] ),
    .X(net425));
 sg13g2_dlygate4sd3_1 hold407 (.A(\clk_counter[15] ),
    .X(net426));
 sg13g2_dlygate4sd3_1 hold408 (.A(_0061_),
    .X(net427));
 sg13g2_dlygate4sd3_1 hold409 (.A(\serial_input.output_case[3] ),
    .X(net428));
 sg13g2_dlygate4sd3_1 hold410 (.A(_0427_),
    .X(net429));
 sg13g2_dlygate4sd3_1 hold411 (.A(\serial_input.output_case[1] ),
    .X(net430));
 sg13g2_dlygate4sd3_1 hold412 (.A(_0040_),
    .X(net431));
 sg13g2_dlygate4sd3_1 hold413 (.A(_1432_),
    .X(net432));
 sg13g2_dlygate4sd3_1 hold414 (.A(\integrator_c_counter.value_output[7] ),
    .X(net433));
 sg13g2_dlygate4sd3_1 hold415 (.A(_0051_),
    .X(net434));
 sg13g2_dlygate4sd3_1 hold416 (.A(\integrator_b_counter.value_output[7] ),
    .X(net435));
 sg13g2_dlygate4sd3_1 hold417 (.A(\integrator_b_counter.value_output[4] ),
    .X(net436));
 sg13g2_dlygate4sd3_1 hold418 (.A(\integrator_b_counter.value_output[3] ),
    .X(net437));
 sg13g2_dlygate4sd3_1 hold419 (.A(_0503_),
    .X(net438));
 sg13g2_dlygate4sd3_1 hold420 (.A(\system_integrator_a_counter.init_flag ),
    .X(net439));
 sg13g2_dlygate4sd3_1 hold421 (.A(_0449_),
    .X(net440));
 sg13g2_dlygate4sd3_1 hold422 (.A(\input_halfprob2_sng_comparator.bits_b[5] ),
    .X(net441));
 sg13g2_dlygate4sd3_1 hold423 (.A(\integrator_c_counter.value_output[4] ),
    .X(net442));
 sg13g2_dlygate4sd3_1 hold424 (.A(\integrator_a_counter.value_output[7] ),
    .X(net443));
 sg13g2_dlygate4sd3_1 hold425 (.A(\integrator_c_output.counter[1] ),
    .X(net444));
 sg13g2_dlygate4sd3_1 hold426 (.A(_0029_),
    .X(net445));
 sg13g2_dlygate4sd3_1 hold427 (.A(\integrator_a_counter.value_output[4] ),
    .X(net446));
 sg13g2_dlygate4sd3_1 hold428 (.A(\integrator_a_output.counter[1] ),
    .X(net447));
 sg13g2_dlygate4sd3_1 hold429 (.A(\integrator_b_counter.value_output[5] ),
    .X(net448));
 sg13g2_dlygate4sd3_1 hold430 (.A(_0505_),
    .X(net449));
 sg13g2_dlygate4sd3_1 hold431 (.A(\system_integrator_b_output.counter[1] ),
    .X(net450));
 sg13g2_dlygate4sd3_1 hold432 (.A(\input_a_sng_comparator.bits_b[4] ),
    .X(net451));
 sg13g2_dlygate4sd3_1 hold433 (.A(\system_integrator_a_output.counter[1] ),
    .X(net452));
 sg13g2_dlygate4sd3_1 hold434 (.A(\system_integrator_a_counter.value_output[7] ),
    .X(net453));
 sg13g2_dlygate4sd3_1 hold435 (.A(\test_integrator_b_output.counter[1] ),
    .X(net454));
 sg13g2_dlygate4sd3_1 hold436 (.A(\test_integrator_a_output.counter[1] ),
    .X(net455));
 sg13g2_dlygate4sd3_1 hold437 (.A(\integrator_c_counter.value_output[2] ),
    .X(net456));
 sg13g2_dlygate4sd3_1 hold438 (.A(_0511_),
    .X(net457));
 sg13g2_dlygate4sd3_1 hold439 (.A(\clk_counter[9] ),
    .X(net458));
 sg13g2_dlygate4sd3_1 hold440 (.A(\system_integrator_a_counter.value_output[6] ),
    .X(net459));
 sg13g2_dlygate4sd3_1 hold441 (.A(\system_integrator_a_counter.value_output[5] ),
    .X(net460));
 sg13g2_dlygate4sd3_1 hold442 (.A(\system_integrator_a_counter.value_output[1] ),
    .X(net461));
 sg13g2_dlygate4sd3_1 hold443 (.A(_0519_),
    .X(net462));
 sg13g2_dlygate4sd3_1 hold444 (.A(\system_integrator_a_counter.value_output[3] ),
    .X(net463));
 sg13g2_dlygate4sd3_1 hold445 (.A(\integrator_a_counter.value_output[5] ),
    .X(net464));
 sg13g2_dlygate4sd3_1 hold446 (.A(_0496_),
    .X(net465));
 sg13g2_dlygate4sd3_1 hold447 (.A(\integrator_b_counter.value_output[2] ),
    .X(net466));
 sg13g2_dlygate4sd3_1 hold448 (.A(\test_integrator_a_counter.value_output[7] ),
    .X(net467));
 sg13g2_dlygate4sd3_1 hold449 (.A(\clk_counter[4] ),
    .X(net468));
 sg13g2_dlygate4sd3_1 hold450 (.A(\clk_counter[5] ),
    .X(net469));
 sg13g2_dlygate4sd3_1 hold451 (.A(\system_integrator_b_counter.value_output[7] ),
    .X(net470));
 sg13g2_dlygate4sd3_1 hold452 (.A(\system_integrator_a_counter.value_output[4] ),
    .X(net471));
 sg13g2_dlygate4sd3_1 hold453 (.A(\system_integrator_b_counter.value_output[3] ),
    .X(net472));
 sg13g2_dlygate4sd3_1 hold454 (.A(\integrator_c_counter.value_output[6] ),
    .X(net473));
 sg13g2_dlygate4sd3_1 hold455 (.A(\integrator_a_counter.value_output[3] ),
    .X(net474));
 sg13g2_dlygate4sd3_1 hold456 (.A(\clk_counter[2] ),
    .X(net475));
 sg13g2_dlygate4sd3_1 hold457 (.A(_1598_),
    .X(net476));
 sg13g2_dlygate4sd3_1 hold458 (.A(_0064_),
    .X(net477));
 sg13g2_dlygate4sd3_1 hold459 (.A(\system_integrator_b_counter.value_output[1] ),
    .X(net478));
 sg13g2_dlygate4sd3_1 hold460 (.A(_0528_),
    .X(net479));
 sg13g2_dlygate4sd3_1 hold461 (.A(\integrator_a_counter.value_output[2] ),
    .X(net480));
 sg13g2_dlygate4sd3_1 hold462 (.A(\integrator_c_output.counter[2] ),
    .X(net481));
 sg13g2_dlygate4sd3_1 hold463 (.A(\test_integrator_b_counter.value_output[2] ),
    .X(net482));
 sg13g2_dlygate4sd3_1 hold464 (.A(_0450_),
    .X(net483));
 sg13g2_dlygate4sd3_1 hold465 (.A(\integrator_a_output.counter[2] ),
    .X(net484));
 sg13g2_dlygate4sd3_1 hold466 (.A(\system_integrator_b_output.counter[2] ),
    .X(net485));
 sg13g2_dlygate4sd3_1 hold467 (.A(\system_integrator_b_counter.value_output[5] ),
    .X(net486));
 sg13g2_dlygate4sd3_1 hold468 (.A(\system_integrator_a_output.counter[2] ),
    .X(net487));
 sg13g2_dlygate4sd3_1 hold469 (.A(\test_integrator_a_counter.value_output[4] ),
    .X(net488));
 sg13g2_dlygate4sd3_1 hold470 (.A(\system_integrator_a_counter.value_output[2] ),
    .X(net489));
 sg13g2_dlygate4sd3_1 hold471 (.A(_1049_),
    .X(net490));
 sg13g2_dlygate4sd3_1 hold472 (.A(\test_integrator_a_counter.value_output[2] ),
    .X(net491));
 sg13g2_dlygate4sd3_1 hold473 (.A(\test_integrator_a_output.counter[2] ),
    .X(net492));
 sg13g2_dlygate4sd3_1 hold474 (.A(\integrator_b_output.counter[2] ),
    .X(net493));
 sg13g2_dlygate4sd3_1 hold475 (.A(\test_integrator_b_output.counter[2] ),
    .X(net494));
 sg13g2_dlygate4sd3_1 hold476 (.A(\test_integrator_b_counter.value_output[0] ),
    .X(net495));
 sg13g2_dlygate4sd3_1 hold477 (.A(\test_integrator_a_counter.value_output[3] ),
    .X(net496));
 sg13g2_dlygate4sd3_1 hold478 (.A(\test_integrator_a_counter.value_output[6] ),
    .X(net497));
 sg13g2_dlygate4sd3_1 hold479 (.A(\integrator_a_counter.value_output[6] ),
    .X(net498));
 sg13g2_dlygate4sd3_1 hold480 (.A(\clk_counter[16] ),
    .X(net499));
 sg13g2_dlygate4sd3_1 hold481 (.A(\system_integrator_b_counter.value_output[6] ),
    .X(net500));
 sg13g2_dlygate4sd3_1 hold482 (.A(\test_integrator_a_counter.value_output[5] ),
    .X(net501));
 sg13g2_dlygate4sd3_1 hold483 (.A(\system_integrator_b_counter.value_output[4] ),
    .X(net502));
 sg13g2_dlygate4sd3_1 hold484 (.A(\system_integrator_b_counter.value_output[2] ),
    .X(net503));
 sg13g2_dlygate4sd3_1 hold485 (.A(\integrator_b_counter.value_output[6] ),
    .X(net504));
 sg13g2_dlygate4sd3_1 hold486 (.A(\serial_input.output_case[1] ),
    .X(net505));
 sg13g2_dlygate4sd3_1 hold487 (.A(\integrator_c_counter.value_output[6] ),
    .X(net506));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_4 FILLER_9_154 ();
 sg13g2_fill_2 FILLER_9_158 ();
 sg13g2_fill_1 FILLER_9_169 ();
 sg13g2_fill_2 FILLER_9_173 ();
 sg13g2_decap_8 FILLER_9_179 ();
 sg13g2_decap_8 FILLER_9_186 ();
 sg13g2_decap_8 FILLER_9_193 ();
 sg13g2_decap_8 FILLER_9_200 ();
 sg13g2_decap_8 FILLER_9_207 ();
 sg13g2_decap_8 FILLER_9_214 ();
 sg13g2_decap_8 FILLER_9_221 ();
 sg13g2_decap_8 FILLER_9_228 ();
 sg13g2_decap_8 FILLER_9_235 ();
 sg13g2_decap_8 FILLER_9_242 ();
 sg13g2_decap_8 FILLER_9_249 ();
 sg13g2_decap_8 FILLER_9_256 ();
 sg13g2_decap_8 FILLER_9_263 ();
 sg13g2_decap_8 FILLER_9_270 ();
 sg13g2_decap_8 FILLER_9_277 ();
 sg13g2_decap_8 FILLER_9_284 ();
 sg13g2_decap_8 FILLER_9_291 ();
 sg13g2_decap_8 FILLER_9_298 ();
 sg13g2_decap_8 FILLER_9_305 ();
 sg13g2_decap_8 FILLER_9_312 ();
 sg13g2_decap_8 FILLER_9_319 ();
 sg13g2_decap_8 FILLER_9_326 ();
 sg13g2_decap_8 FILLER_9_333 ();
 sg13g2_decap_8 FILLER_9_340 ();
 sg13g2_decap_8 FILLER_9_347 ();
 sg13g2_decap_8 FILLER_9_354 ();
 sg13g2_decap_8 FILLER_9_361 ();
 sg13g2_decap_8 FILLER_9_368 ();
 sg13g2_decap_8 FILLER_9_375 ();
 sg13g2_decap_8 FILLER_9_382 ();
 sg13g2_decap_8 FILLER_9_389 ();
 sg13g2_decap_8 FILLER_9_396 ();
 sg13g2_decap_4 FILLER_9_403 ();
 sg13g2_fill_2 FILLER_9_407 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_4 FILLER_10_147 ();
 sg13g2_fill_2 FILLER_10_163 ();
 sg13g2_decap_8 FILLER_10_201 ();
 sg13g2_decap_8 FILLER_10_208 ();
 sg13g2_decap_8 FILLER_10_215 ();
 sg13g2_decap_8 FILLER_10_222 ();
 sg13g2_decap_8 FILLER_10_229 ();
 sg13g2_decap_8 FILLER_10_236 ();
 sg13g2_decap_8 FILLER_10_243 ();
 sg13g2_decap_8 FILLER_10_250 ();
 sg13g2_decap_8 FILLER_10_257 ();
 sg13g2_decap_8 FILLER_10_264 ();
 sg13g2_decap_8 FILLER_10_271 ();
 sg13g2_decap_8 FILLER_10_278 ();
 sg13g2_decap_8 FILLER_10_285 ();
 sg13g2_decap_8 FILLER_10_292 ();
 sg13g2_decap_8 FILLER_10_299 ();
 sg13g2_decap_8 FILLER_10_306 ();
 sg13g2_decap_8 FILLER_10_313 ();
 sg13g2_decap_8 FILLER_10_320 ();
 sg13g2_decap_8 FILLER_10_327 ();
 sg13g2_decap_8 FILLER_10_334 ();
 sg13g2_decap_8 FILLER_10_341 ();
 sg13g2_decap_8 FILLER_10_348 ();
 sg13g2_decap_8 FILLER_10_355 ();
 sg13g2_decap_8 FILLER_10_362 ();
 sg13g2_decap_8 FILLER_10_369 ();
 sg13g2_decap_8 FILLER_10_376 ();
 sg13g2_decap_8 FILLER_10_383 ();
 sg13g2_decap_8 FILLER_10_390 ();
 sg13g2_decap_8 FILLER_10_397 ();
 sg13g2_decap_4 FILLER_10_404 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_fill_2 FILLER_11_181 ();
 sg13g2_fill_2 FILLER_11_202 ();
 sg13g2_decap_8 FILLER_11_213 ();
 sg13g2_decap_8 FILLER_11_220 ();
 sg13g2_decap_8 FILLER_11_227 ();
 sg13g2_decap_8 FILLER_11_234 ();
 sg13g2_decap_8 FILLER_11_241 ();
 sg13g2_decap_8 FILLER_11_248 ();
 sg13g2_decap_8 FILLER_11_255 ();
 sg13g2_decap_8 FILLER_11_262 ();
 sg13g2_decap_8 FILLER_11_269 ();
 sg13g2_decap_8 FILLER_11_276 ();
 sg13g2_decap_8 FILLER_11_283 ();
 sg13g2_decap_8 FILLER_11_290 ();
 sg13g2_decap_8 FILLER_11_297 ();
 sg13g2_decap_8 FILLER_11_304 ();
 sg13g2_decap_8 FILLER_11_311 ();
 sg13g2_decap_8 FILLER_11_318 ();
 sg13g2_decap_8 FILLER_11_325 ();
 sg13g2_decap_8 FILLER_11_332 ();
 sg13g2_decap_8 FILLER_11_339 ();
 sg13g2_decap_8 FILLER_11_346 ();
 sg13g2_decap_8 FILLER_11_353 ();
 sg13g2_decap_8 FILLER_11_360 ();
 sg13g2_decap_8 FILLER_11_367 ();
 sg13g2_decap_8 FILLER_11_374 ();
 sg13g2_decap_8 FILLER_11_381 ();
 sg13g2_decap_8 FILLER_11_388 ();
 sg13g2_decap_8 FILLER_11_395 ();
 sg13g2_decap_8 FILLER_11_402 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_4 FILLER_12_126 ();
 sg13g2_fill_1 FILLER_12_162 ();
 sg13g2_decap_8 FILLER_12_215 ();
 sg13g2_decap_8 FILLER_12_222 ();
 sg13g2_decap_8 FILLER_12_229 ();
 sg13g2_decap_8 FILLER_12_236 ();
 sg13g2_fill_2 FILLER_12_243 ();
 sg13g2_fill_1 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_fill_1 FILLER_12_266 ();
 sg13g2_fill_1 FILLER_12_274 ();
 sg13g2_decap_8 FILLER_12_278 ();
 sg13g2_decap_8 FILLER_12_285 ();
 sg13g2_decap_8 FILLER_12_292 ();
 sg13g2_decap_8 FILLER_12_299 ();
 sg13g2_decap_8 FILLER_12_306 ();
 sg13g2_decap_8 FILLER_12_313 ();
 sg13g2_decap_8 FILLER_12_320 ();
 sg13g2_decap_8 FILLER_12_327 ();
 sg13g2_decap_8 FILLER_12_334 ();
 sg13g2_decap_8 FILLER_12_341 ();
 sg13g2_decap_8 FILLER_12_348 ();
 sg13g2_decap_8 FILLER_12_355 ();
 sg13g2_decap_8 FILLER_12_362 ();
 sg13g2_decap_8 FILLER_12_369 ();
 sg13g2_decap_8 FILLER_12_376 ();
 sg13g2_decap_8 FILLER_12_383 ();
 sg13g2_decap_8 FILLER_12_390 ();
 sg13g2_decap_8 FILLER_12_397 ();
 sg13g2_decap_4 FILLER_12_404 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_4 FILLER_13_126 ();
 sg13g2_fill_2 FILLER_13_130 ();
 sg13g2_fill_2 FILLER_13_158 ();
 sg13g2_fill_2 FILLER_13_169 ();
 sg13g2_fill_1 FILLER_13_171 ();
 sg13g2_decap_8 FILLER_13_226 ();
 sg13g2_decap_8 FILLER_13_233 ();
 sg13g2_decap_8 FILLER_13_285 ();
 sg13g2_decap_8 FILLER_13_292 ();
 sg13g2_decap_8 FILLER_13_299 ();
 sg13g2_decap_8 FILLER_13_306 ();
 sg13g2_decap_8 FILLER_13_313 ();
 sg13g2_decap_8 FILLER_13_320 ();
 sg13g2_decap_8 FILLER_13_327 ();
 sg13g2_decap_8 FILLER_13_334 ();
 sg13g2_decap_8 FILLER_13_341 ();
 sg13g2_decap_8 FILLER_13_348 ();
 sg13g2_decap_8 FILLER_13_355 ();
 sg13g2_decap_8 FILLER_13_362 ();
 sg13g2_decap_8 FILLER_13_369 ();
 sg13g2_decap_8 FILLER_13_376 ();
 sg13g2_decap_8 FILLER_13_383 ();
 sg13g2_decap_8 FILLER_13_390 ();
 sg13g2_decap_8 FILLER_13_397 ();
 sg13g2_decap_4 FILLER_13_404 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_fill_1 FILLER_14_133 ();
 sg13g2_fill_1 FILLER_14_161 ();
 sg13g2_decap_4 FILLER_14_228 ();
 sg13g2_decap_8 FILLER_14_296 ();
 sg13g2_decap_8 FILLER_14_303 ();
 sg13g2_decap_8 FILLER_14_310 ();
 sg13g2_decap_8 FILLER_14_317 ();
 sg13g2_decap_8 FILLER_14_324 ();
 sg13g2_decap_8 FILLER_14_331 ();
 sg13g2_decap_8 FILLER_14_338 ();
 sg13g2_decap_8 FILLER_14_345 ();
 sg13g2_decap_8 FILLER_14_352 ();
 sg13g2_decap_8 FILLER_14_359 ();
 sg13g2_decap_8 FILLER_14_366 ();
 sg13g2_decap_8 FILLER_14_373 ();
 sg13g2_decap_8 FILLER_14_380 ();
 sg13g2_decap_8 FILLER_14_387 ();
 sg13g2_decap_8 FILLER_14_394 ();
 sg13g2_decap_8 FILLER_14_401 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_4 FILLER_15_126 ();
 sg13g2_fill_1 FILLER_15_163 ();
 sg13g2_fill_1 FILLER_15_173 ();
 sg13g2_decap_8 FILLER_15_312 ();
 sg13g2_decap_8 FILLER_15_319 ();
 sg13g2_decap_8 FILLER_15_326 ();
 sg13g2_decap_8 FILLER_15_333 ();
 sg13g2_decap_8 FILLER_15_340 ();
 sg13g2_decap_8 FILLER_15_347 ();
 sg13g2_decap_8 FILLER_15_354 ();
 sg13g2_decap_8 FILLER_15_361 ();
 sg13g2_decap_8 FILLER_15_368 ();
 sg13g2_decap_8 FILLER_15_375 ();
 sg13g2_decap_8 FILLER_15_382 ();
 sg13g2_decap_8 FILLER_15_389 ();
 sg13g2_decap_8 FILLER_15_396 ();
 sg13g2_decap_4 FILLER_15_403 ();
 sg13g2_fill_2 FILLER_15_407 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_4 FILLER_16_126 ();
 sg13g2_fill_1 FILLER_16_130 ();
 sg13g2_fill_2 FILLER_16_157 ();
 sg13g2_fill_2 FILLER_16_274 ();
 sg13g2_fill_2 FILLER_16_285 ();
 sg13g2_decap_8 FILLER_16_320 ();
 sg13g2_decap_8 FILLER_16_327 ();
 sg13g2_decap_8 FILLER_16_334 ();
 sg13g2_decap_8 FILLER_16_341 ();
 sg13g2_decap_8 FILLER_16_348 ();
 sg13g2_decap_8 FILLER_16_355 ();
 sg13g2_decap_8 FILLER_16_362 ();
 sg13g2_decap_8 FILLER_16_369 ();
 sg13g2_decap_8 FILLER_16_376 ();
 sg13g2_decap_8 FILLER_16_383 ();
 sg13g2_decap_8 FILLER_16_390 ();
 sg13g2_decap_8 FILLER_16_397 ();
 sg13g2_decap_4 FILLER_16_404 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_fill_1 FILLER_17_164 ();
 sg13g2_fill_1 FILLER_17_175 ();
 sg13g2_fill_2 FILLER_17_181 ();
 sg13g2_fill_1 FILLER_17_188 ();
 sg13g2_fill_2 FILLER_17_194 ();
 sg13g2_decap_8 FILLER_17_220 ();
 sg13g2_decap_8 FILLER_17_227 ();
 sg13g2_fill_2 FILLER_17_234 ();
 sg13g2_fill_1 FILLER_17_251 ();
 sg13g2_fill_2 FILLER_17_258 ();
 sg13g2_fill_2 FILLER_17_280 ();
 sg13g2_fill_2 FILLER_17_292 ();
 sg13g2_decap_8 FILLER_17_325 ();
 sg13g2_decap_8 FILLER_17_332 ();
 sg13g2_decap_8 FILLER_17_339 ();
 sg13g2_decap_8 FILLER_17_346 ();
 sg13g2_decap_8 FILLER_17_353 ();
 sg13g2_decap_8 FILLER_17_360 ();
 sg13g2_decap_8 FILLER_17_367 ();
 sg13g2_decap_8 FILLER_17_374 ();
 sg13g2_decap_8 FILLER_17_381 ();
 sg13g2_decap_8 FILLER_17_388 ();
 sg13g2_decap_8 FILLER_17_395 ();
 sg13g2_decap_8 FILLER_17_402 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_4 FILLER_18_70 ();
 sg13g2_fill_2 FILLER_18_78 ();
 sg13g2_fill_1 FILLER_18_80 ();
 sg13g2_decap_4 FILLER_18_96 ();
 sg13g2_fill_2 FILLER_18_100 ();
 sg13g2_decap_8 FILLER_18_108 ();
 sg13g2_decap_8 FILLER_18_115 ();
 sg13g2_fill_1 FILLER_18_122 ();
 sg13g2_fill_1 FILLER_18_152 ();
 sg13g2_fill_2 FILLER_18_162 ();
 sg13g2_fill_2 FILLER_18_204 ();
 sg13g2_decap_4 FILLER_18_222 ();
 sg13g2_fill_1 FILLER_18_226 ();
 sg13g2_fill_2 FILLER_18_233 ();
 sg13g2_fill_2 FILLER_18_327 ();
 sg13g2_decap_8 FILLER_18_344 ();
 sg13g2_decap_8 FILLER_18_351 ();
 sg13g2_decap_8 FILLER_18_358 ();
 sg13g2_decap_8 FILLER_18_365 ();
 sg13g2_decap_8 FILLER_18_372 ();
 sg13g2_decap_8 FILLER_18_379 ();
 sg13g2_decap_8 FILLER_18_386 ();
 sg13g2_decap_8 FILLER_18_393 ();
 sg13g2_decap_8 FILLER_18_400 ();
 sg13g2_fill_2 FILLER_18_407 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_fill_2 FILLER_19_56 ();
 sg13g2_fill_1 FILLER_19_119 ();
 sg13g2_fill_1 FILLER_19_130 ();
 sg13g2_fill_1 FILLER_19_148 ();
 sg13g2_fill_2 FILLER_19_154 ();
 sg13g2_fill_1 FILLER_19_187 ();
 sg13g2_fill_2 FILLER_19_222 ();
 sg13g2_fill_1 FILLER_19_329 ();
 sg13g2_decap_8 FILLER_19_347 ();
 sg13g2_decap_8 FILLER_19_354 ();
 sg13g2_decap_8 FILLER_19_361 ();
 sg13g2_decap_8 FILLER_19_368 ();
 sg13g2_decap_8 FILLER_19_375 ();
 sg13g2_decap_8 FILLER_19_382 ();
 sg13g2_decap_8 FILLER_19_389 ();
 sg13g2_decap_8 FILLER_19_396 ();
 sg13g2_decap_4 FILLER_19_403 ();
 sg13g2_fill_2 FILLER_19_407 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_fill_1 FILLER_20_90 ();
 sg13g2_fill_2 FILLER_20_143 ();
 sg13g2_fill_2 FILLER_20_171 ();
 sg13g2_decap_8 FILLER_20_351 ();
 sg13g2_decap_8 FILLER_20_358 ();
 sg13g2_decap_8 FILLER_20_365 ();
 sg13g2_decap_8 FILLER_20_372 ();
 sg13g2_decap_8 FILLER_20_379 ();
 sg13g2_decap_8 FILLER_20_386 ();
 sg13g2_decap_8 FILLER_20_393 ();
 sg13g2_decap_8 FILLER_20_400 ();
 sg13g2_fill_2 FILLER_20_407 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_4 FILLER_21_42 ();
 sg13g2_fill_1 FILLER_21_46 ();
 sg13g2_fill_2 FILLER_21_144 ();
 sg13g2_fill_1 FILLER_21_185 ();
 sg13g2_fill_2 FILLER_21_271 ();
 sg13g2_fill_2 FILLER_21_312 ();
 sg13g2_decap_8 FILLER_21_361 ();
 sg13g2_decap_8 FILLER_21_368 ();
 sg13g2_decap_8 FILLER_21_375 ();
 sg13g2_decap_8 FILLER_21_382 ();
 sg13g2_decap_8 FILLER_21_389 ();
 sg13g2_decap_8 FILLER_21_396 ();
 sg13g2_decap_4 FILLER_21_403 ();
 sg13g2_fill_2 FILLER_21_407 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_4 FILLER_22_28 ();
 sg13g2_fill_2 FILLER_22_32 ();
 sg13g2_fill_2 FILLER_22_60 ();
 sg13g2_fill_2 FILLER_22_95 ();
 sg13g2_fill_2 FILLER_22_145 ();
 sg13g2_fill_1 FILLER_22_152 ();
 sg13g2_fill_1 FILLER_22_171 ();
 sg13g2_fill_1 FILLER_22_191 ();
 sg13g2_fill_2 FILLER_22_220 ();
 sg13g2_fill_2 FILLER_22_244 ();
 sg13g2_fill_2 FILLER_22_280 ();
 sg13g2_fill_2 FILLER_22_306 ();
 sg13g2_fill_2 FILLER_22_317 ();
 sg13g2_decap_8 FILLER_22_354 ();
 sg13g2_decap_8 FILLER_22_361 ();
 sg13g2_decap_8 FILLER_22_368 ();
 sg13g2_decap_8 FILLER_22_375 ();
 sg13g2_decap_8 FILLER_22_382 ();
 sg13g2_decap_8 FILLER_22_389 ();
 sg13g2_decap_8 FILLER_22_396 ();
 sg13g2_decap_4 FILLER_22_403 ();
 sg13g2_fill_2 FILLER_22_407 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_fill_1 FILLER_23_35 ();
 sg13g2_fill_1 FILLER_23_65 ();
 sg13g2_fill_1 FILLER_23_92 ();
 sg13g2_fill_1 FILLER_23_141 ();
 sg13g2_fill_1 FILLER_23_173 ();
 sg13g2_fill_1 FILLER_23_179 ();
 sg13g2_fill_2 FILLER_23_206 ();
 sg13g2_fill_1 FILLER_23_234 ();
 sg13g2_fill_2 FILLER_23_244 ();
 sg13g2_fill_1 FILLER_23_329 ();
 sg13g2_decap_8 FILLER_23_348 ();
 sg13g2_decap_8 FILLER_23_355 ();
 sg13g2_decap_8 FILLER_23_362 ();
 sg13g2_decap_8 FILLER_23_369 ();
 sg13g2_decap_8 FILLER_23_376 ();
 sg13g2_decap_8 FILLER_23_383 ();
 sg13g2_decap_8 FILLER_23_390 ();
 sg13g2_decap_8 FILLER_23_397 ();
 sg13g2_decap_4 FILLER_23_404 ();
 sg13g2_fill_1 FILLER_23_408 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_fill_1 FILLER_24_28 ();
 sg13g2_fill_1 FILLER_24_65 ();
 sg13g2_fill_1 FILLER_24_234 ();
 sg13g2_fill_2 FILLER_24_290 ();
 sg13g2_decap_8 FILLER_24_344 ();
 sg13g2_decap_8 FILLER_24_360 ();
 sg13g2_decap_8 FILLER_24_367 ();
 sg13g2_decap_8 FILLER_24_374 ();
 sg13g2_decap_8 FILLER_24_381 ();
 sg13g2_decap_8 FILLER_24_388 ();
 sg13g2_decap_8 FILLER_24_395 ();
 sg13g2_decap_8 FILLER_24_402 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_fill_1 FILLER_25_28 ();
 sg13g2_fill_1 FILLER_25_73 ();
 sg13g2_fill_1 FILLER_25_102 ();
 sg13g2_fill_1 FILLER_25_112 ();
 sg13g2_fill_1 FILLER_25_122 ();
 sg13g2_fill_1 FILLER_25_175 ();
 sg13g2_fill_1 FILLER_25_212 ();
 sg13g2_fill_1 FILLER_25_239 ();
 sg13g2_fill_2 FILLER_25_259 ();
 sg13g2_fill_2 FILLER_25_307 ();
 sg13g2_fill_1 FILLER_25_326 ();
 sg13g2_fill_2 FILLER_25_342 ();
 sg13g2_fill_1 FILLER_25_353 ();
 sg13g2_decap_8 FILLER_25_381 ();
 sg13g2_decap_8 FILLER_25_388 ();
 sg13g2_decap_8 FILLER_25_395 ();
 sg13g2_decap_8 FILLER_25_402 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_4 FILLER_26_28 ();
 sg13g2_fill_2 FILLER_26_32 ();
 sg13g2_fill_2 FILLER_26_60 ();
 sg13g2_fill_2 FILLER_26_128 ();
 sg13g2_fill_1 FILLER_26_167 ();
 sg13g2_fill_2 FILLER_26_182 ();
 sg13g2_decap_4 FILLER_26_209 ();
 sg13g2_fill_2 FILLER_26_219 ();
 sg13g2_fill_1 FILLER_26_280 ();
 sg13g2_fill_2 FILLER_26_317 ();
 sg13g2_fill_1 FILLER_26_319 ();
 sg13g2_fill_1 FILLER_26_385 ();
 sg13g2_decap_8 FILLER_26_389 ();
 sg13g2_decap_8 FILLER_26_396 ();
 sg13g2_decap_4 FILLER_26_403 ();
 sg13g2_fill_2 FILLER_26_407 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_4 FILLER_27_21 ();
 sg13g2_fill_2 FILLER_27_25 ();
 sg13g2_fill_1 FILLER_27_73 ();
 sg13g2_fill_2 FILLER_27_87 ();
 sg13g2_fill_2 FILLER_27_92 ();
 sg13g2_fill_1 FILLER_27_123 ();
 sg13g2_fill_1 FILLER_27_159 ();
 sg13g2_fill_1 FILLER_27_178 ();
 sg13g2_fill_2 FILLER_27_188 ();
 sg13g2_fill_1 FILLER_27_230 ();
 sg13g2_fill_2 FILLER_27_243 ();
 sg13g2_fill_2 FILLER_27_309 ();
 sg13g2_fill_1 FILLER_27_311 ();
 sg13g2_fill_2 FILLER_27_351 ();
 sg13g2_decap_8 FILLER_27_401 ();
 sg13g2_fill_1 FILLER_27_408 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_4 FILLER_28_28 ();
 sg13g2_fill_2 FILLER_28_81 ();
 sg13g2_fill_1 FILLER_28_83 ();
 sg13g2_decap_8 FILLER_28_138 ();
 sg13g2_fill_2 FILLER_28_148 ();
 sg13g2_fill_1 FILLER_28_150 ();
 sg13g2_fill_2 FILLER_28_192 ();
 sg13g2_fill_2 FILLER_28_240 ();
 sg13g2_fill_1 FILLER_28_306 ();
 sg13g2_fill_1 FILLER_28_354 ();
 sg13g2_fill_1 FILLER_28_398 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_4 FILLER_29_35 ();
 sg13g2_decap_4 FILLER_29_54 ();
 sg13g2_fill_1 FILLER_29_58 ();
 sg13g2_fill_2 FILLER_29_94 ();
 sg13g2_decap_4 FILLER_29_131 ();
 sg13g2_fill_2 FILLER_29_135 ();
 sg13g2_decap_4 FILLER_29_145 ();
 sg13g2_fill_1 FILLER_29_149 ();
 sg13g2_decap_8 FILLER_29_205 ();
 sg13g2_decap_8 FILLER_29_212 ();
 sg13g2_fill_1 FILLER_29_219 ();
 sg13g2_decap_4 FILLER_29_239 ();
 sg13g2_fill_1 FILLER_29_265 ();
 sg13g2_fill_1 FILLER_29_297 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_fill_2 FILLER_30_72 ();
 sg13g2_fill_1 FILLER_30_74 ();
 sg13g2_decap_4 FILLER_30_120 ();
 sg13g2_fill_2 FILLER_30_124 ();
 sg13g2_fill_1 FILLER_30_131 ();
 sg13g2_decap_4 FILLER_30_162 ();
 sg13g2_fill_1 FILLER_30_166 ();
 sg13g2_fill_2 FILLER_30_175 ();
 sg13g2_fill_1 FILLER_30_177 ();
 sg13g2_decap_4 FILLER_30_220 ();
 sg13g2_fill_2 FILLER_30_224 ();
 sg13g2_fill_1 FILLER_30_246 ();
 sg13g2_fill_2 FILLER_30_262 ();
 sg13g2_fill_2 FILLER_30_306 ();
 sg13g2_fill_1 FILLER_30_348 ();
 sg13g2_fill_1 FILLER_30_358 ();
 sg13g2_fill_1 FILLER_30_378 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_4 FILLER_31_42 ();
 sg13g2_fill_2 FILLER_31_46 ();
 sg13g2_fill_1 FILLER_31_94 ();
 sg13g2_fill_2 FILLER_31_104 ();
 sg13g2_fill_1 FILLER_31_115 ();
 sg13g2_fill_2 FILLER_31_204 ();
 sg13g2_fill_2 FILLER_31_210 ();
 sg13g2_fill_1 FILLER_31_212 ();
 sg13g2_fill_2 FILLER_31_222 ();
 sg13g2_fill_1 FILLER_31_227 ();
 sg13g2_decap_8 FILLER_31_234 ();
 sg13g2_fill_2 FILLER_31_241 ();
 sg13g2_fill_1 FILLER_31_243 ();
 sg13g2_fill_2 FILLER_31_280 ();
 sg13g2_fill_2 FILLER_31_291 ();
 sg13g2_fill_1 FILLER_31_330 ();
 sg13g2_fill_2 FILLER_31_334 ();
 sg13g2_fill_1 FILLER_31_351 ();
 sg13g2_fill_1 FILLER_31_402 ();
 sg13g2_fill_1 FILLER_31_408 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_4 FILLER_32_42 ();
 sg13g2_fill_2 FILLER_32_46 ();
 sg13g2_fill_2 FILLER_32_80 ();
 sg13g2_fill_1 FILLER_32_161 ();
 sg13g2_fill_2 FILLER_32_196 ();
 sg13g2_fill_1 FILLER_32_198 ();
 sg13g2_fill_2 FILLER_32_242 ();
 sg13g2_fill_2 FILLER_32_311 ();
 sg13g2_fill_2 FILLER_32_383 ();
 sg13g2_fill_1 FILLER_32_408 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_fill_2 FILLER_33_56 ();
 sg13g2_decap_4 FILLER_33_61 ();
 sg13g2_fill_1 FILLER_33_114 ();
 sg13g2_fill_2 FILLER_33_149 ();
 sg13g2_fill_2 FILLER_33_164 ();
 sg13g2_fill_2 FILLER_33_192 ();
 sg13g2_fill_1 FILLER_33_194 ();
 sg13g2_fill_2 FILLER_33_255 ();
 sg13g2_fill_1 FILLER_33_257 ();
 sg13g2_fill_2 FILLER_33_309 ();
 sg13g2_fill_2 FILLER_33_340 ();
 sg13g2_fill_1 FILLER_33_360 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_4 FILLER_34_49 ();
 sg13g2_fill_1 FILLER_34_53 ();
 sg13g2_fill_2 FILLER_34_74 ();
 sg13g2_decap_4 FILLER_34_142 ();
 sg13g2_fill_2 FILLER_34_149 ();
 sg13g2_fill_2 FILLER_34_190 ();
 sg13g2_fill_2 FILLER_34_203 ();
 sg13g2_fill_1 FILLER_34_205 ();
 sg13g2_fill_1 FILLER_34_219 ();
 sg13g2_fill_2 FILLER_34_265 ();
 sg13g2_fill_1 FILLER_34_314 ();
 sg13g2_fill_2 FILLER_34_341 ();
 sg13g2_fill_1 FILLER_34_343 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_fill_2 FILLER_35_79 ();
 sg13g2_fill_1 FILLER_35_109 ();
 sg13g2_fill_2 FILLER_35_148 ();
 sg13g2_fill_1 FILLER_35_150 ();
 sg13g2_fill_1 FILLER_35_176 ();
 sg13g2_fill_1 FILLER_35_215 ();
 sg13g2_fill_2 FILLER_35_238 ();
 sg13g2_fill_2 FILLER_35_250 ();
 sg13g2_fill_2 FILLER_35_291 ();
 sg13g2_decap_4 FILLER_35_315 ();
 sg13g2_decap_4 FILLER_35_337 ();
 sg13g2_fill_2 FILLER_35_341 ();
 sg13g2_fill_1 FILLER_35_374 ();
 sg13g2_fill_2 FILLER_35_389 ();
 sg13g2_fill_1 FILLER_35_408 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_4 FILLER_36_56 ();
 sg13g2_fill_2 FILLER_36_60 ();
 sg13g2_fill_2 FILLER_36_98 ();
 sg13g2_fill_1 FILLER_36_126 ();
 sg13g2_fill_1 FILLER_36_131 ();
 sg13g2_fill_1 FILLER_36_138 ();
 sg13g2_fill_2 FILLER_36_148 ();
 sg13g2_fill_1 FILLER_36_150 ();
 sg13g2_fill_1 FILLER_36_177 ();
 sg13g2_decap_8 FILLER_36_213 ();
 sg13g2_fill_2 FILLER_36_224 ();
 sg13g2_decap_4 FILLER_36_234 ();
 sg13g2_decap_8 FILLER_36_241 ();
 sg13g2_decap_8 FILLER_36_248 ();
 sg13g2_fill_2 FILLER_36_255 ();
 sg13g2_fill_2 FILLER_36_260 ();
 sg13g2_fill_1 FILLER_36_262 ();
 sg13g2_decap_8 FILLER_36_270 ();
 sg13g2_decap_4 FILLER_36_277 ();
 sg13g2_fill_1 FILLER_36_281 ();
 sg13g2_decap_8 FILLER_36_286 ();
 sg13g2_decap_8 FILLER_36_293 ();
 sg13g2_fill_2 FILLER_36_300 ();
 sg13g2_fill_1 FILLER_36_302 ();
 sg13g2_fill_1 FILLER_36_306 ();
 sg13g2_decap_4 FILLER_36_312 ();
 sg13g2_fill_1 FILLER_36_337 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_fill_1 FILLER_37_75 ();
 sg13g2_fill_1 FILLER_37_94 ();
 sg13g2_decap_4 FILLER_37_127 ();
 sg13g2_fill_1 FILLER_37_131 ();
 sg13g2_decap_8 FILLER_37_141 ();
 sg13g2_decap_8 FILLER_37_148 ();
 sg13g2_fill_2 FILLER_37_155 ();
 sg13g2_fill_2 FILLER_37_182 ();
 sg13g2_decap_4 FILLER_37_223 ();
 sg13g2_fill_2 FILLER_37_227 ();
 sg13g2_fill_2 FILLER_37_264 ();
 sg13g2_fill_2 FILLER_37_271 ();
 sg13g2_fill_1 FILLER_37_273 ();
 sg13g2_decap_8 FILLER_37_303 ();
 sg13g2_fill_2 FILLER_37_381 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_4 FILLER_38_42 ();
 sg13g2_fill_2 FILLER_38_96 ();
 sg13g2_fill_1 FILLER_38_107 ();
 sg13g2_fill_2 FILLER_38_136 ();
 sg13g2_decap_8 FILLER_38_152 ();
 sg13g2_decap_8 FILLER_38_159 ();
 sg13g2_decap_4 FILLER_38_166 ();
 sg13g2_fill_2 FILLER_38_170 ();
 sg13g2_fill_1 FILLER_38_180 ();
 sg13g2_decap_4 FILLER_38_186 ();
 sg13g2_fill_1 FILLER_38_196 ();
 sg13g2_decap_8 FILLER_38_202 ();
 sg13g2_decap_8 FILLER_38_209 ();
 sg13g2_decap_8 FILLER_38_216 ();
 sg13g2_decap_8 FILLER_38_223 ();
 sg13g2_fill_1 FILLER_38_230 ();
 sg13g2_decap_8 FILLER_38_234 ();
 sg13g2_fill_2 FILLER_38_241 ();
 sg13g2_fill_2 FILLER_38_248 ();
 sg13g2_fill_2 FILLER_38_265 ();
 sg13g2_fill_2 FILLER_38_293 ();
 sg13g2_fill_1 FILLER_38_295 ();
 sg13g2_fill_1 FILLER_38_308 ();
 sg13g2_fill_2 FILLER_38_322 ();
 sg13g2_fill_1 FILLER_38_333 ();
 sg13g2_fill_1 FILLER_38_343 ();
 sg13g2_fill_2 FILLER_38_372 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_14 ();
 sg13g2_decap_8 FILLER_39_21 ();
 sg13g2_decap_8 FILLER_39_28 ();
 sg13g2_decap_8 FILLER_39_35 ();
 sg13g2_decap_8 FILLER_39_42 ();
 sg13g2_fill_2 FILLER_39_49 ();
 sg13g2_fill_1 FILLER_39_51 ();
 sg13g2_fill_2 FILLER_39_109 ();
 sg13g2_fill_1 FILLER_39_126 ();
 sg13g2_fill_1 FILLER_39_169 ();
 sg13g2_decap_8 FILLER_39_175 ();
 sg13g2_decap_4 FILLER_39_182 ();
 sg13g2_fill_1 FILLER_39_186 ();
 sg13g2_decap_4 FILLER_39_202 ();
 sg13g2_fill_1 FILLER_39_206 ();
 sg13g2_fill_2 FILLER_39_265 ();
 sg13g2_fill_1 FILLER_39_267 ();
 sg13g2_decap_4 FILLER_39_274 ();
 sg13g2_fill_2 FILLER_39_278 ();
 sg13g2_fill_2 FILLER_39_305 ();
 sg13g2_fill_2 FILLER_39_318 ();
 sg13g2_fill_1 FILLER_39_351 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_14 ();
 sg13g2_decap_8 FILLER_40_21 ();
 sg13g2_decap_8 FILLER_40_28 ();
 sg13g2_decap_8 FILLER_40_35 ();
 sg13g2_decap_8 FILLER_40_42 ();
 sg13g2_decap_8 FILLER_40_49 ();
 sg13g2_decap_4 FILLER_40_56 ();
 sg13g2_fill_1 FILLER_40_64 ();
 sg13g2_fill_1 FILLER_40_77 ();
 sg13g2_fill_1 FILLER_40_125 ();
 sg13g2_fill_2 FILLER_40_133 ();
 sg13g2_fill_1 FILLER_40_135 ();
 sg13g2_fill_2 FILLER_40_182 ();
 sg13g2_fill_2 FILLER_40_205 ();
 sg13g2_fill_1 FILLER_40_207 ();
 sg13g2_fill_2 FILLER_40_277 ();
 sg13g2_fill_1 FILLER_40_279 ();
 sg13g2_fill_2 FILLER_40_300 ();
 sg13g2_fill_1 FILLER_40_307 ();
 sg13g2_fill_1 FILLER_40_313 ();
 sg13g2_fill_1 FILLER_40_398 ();
 sg13g2_fill_1 FILLER_40_408 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_8 FILLER_41_14 ();
 sg13g2_decap_8 FILLER_41_21 ();
 sg13g2_decap_8 FILLER_41_28 ();
 sg13g2_decap_8 FILLER_41_35 ();
 sg13g2_decap_8 FILLER_41_42 ();
 sg13g2_decap_8 FILLER_41_49 ();
 sg13g2_decap_8 FILLER_41_56 ();
 sg13g2_decap_8 FILLER_41_63 ();
 sg13g2_decap_8 FILLER_41_70 ();
 sg13g2_fill_2 FILLER_41_77 ();
 sg13g2_fill_2 FILLER_41_87 ();
 sg13g2_fill_1 FILLER_41_89 ();
 sg13g2_fill_2 FILLER_41_93 ();
 sg13g2_fill_1 FILLER_41_126 ();
 sg13g2_fill_2 FILLER_41_156 ();
 sg13g2_decap_8 FILLER_41_164 ();
 sg13g2_decap_8 FILLER_41_197 ();
 sg13g2_decap_8 FILLER_41_204 ();
 sg13g2_fill_1 FILLER_41_211 ();
 sg13g2_fill_1 FILLER_41_312 ();
 sg13g2_fill_2 FILLER_41_345 ();
 sg13g2_fill_1 FILLER_41_347 ();
 sg13g2_fill_1 FILLER_41_353 ();
 sg13g2_fill_1 FILLER_41_359 ();
 sg13g2_fill_2 FILLER_41_375 ();
 sg13g2_fill_1 FILLER_41_377 ();
 sg13g2_fill_2 FILLER_41_383 ();
 sg13g2_fill_1 FILLER_41_408 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_decap_8 FILLER_42_14 ();
 sg13g2_decap_8 FILLER_42_21 ();
 sg13g2_decap_8 FILLER_42_28 ();
 sg13g2_decap_8 FILLER_42_35 ();
 sg13g2_decap_8 FILLER_42_42 ();
 sg13g2_decap_8 FILLER_42_49 ();
 sg13g2_decap_8 FILLER_42_56 ();
 sg13g2_decap_8 FILLER_42_63 ();
 sg13g2_decap_4 FILLER_42_70 ();
 sg13g2_decap_8 FILLER_42_77 ();
 sg13g2_decap_8 FILLER_42_84 ();
 sg13g2_decap_8 FILLER_42_91 ();
 sg13g2_decap_4 FILLER_42_98 ();
 sg13g2_fill_1 FILLER_42_102 ();
 sg13g2_fill_2 FILLER_42_116 ();
 sg13g2_fill_2 FILLER_42_134 ();
 sg13g2_fill_2 FILLER_42_164 ();
 sg13g2_fill_1 FILLER_42_166 ();
 sg13g2_fill_1 FILLER_42_210 ();
 sg13g2_decap_8 FILLER_42_226 ();
 sg13g2_fill_2 FILLER_42_233 ();
 sg13g2_fill_1 FILLER_42_250 ();
 sg13g2_decap_4 FILLER_42_270 ();
 sg13g2_decap_4 FILLER_42_340 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_decap_8 FILLER_43_14 ();
 sg13g2_decap_8 FILLER_43_21 ();
 sg13g2_decap_8 FILLER_43_28 ();
 sg13g2_decap_8 FILLER_43_35 ();
 sg13g2_decap_8 FILLER_43_42 ();
 sg13g2_decap_8 FILLER_43_49 ();
 sg13g2_decap_8 FILLER_43_56 ();
 sg13g2_fill_1 FILLER_43_63 ();
 sg13g2_fill_1 FILLER_43_90 ();
 sg13g2_decap_4 FILLER_43_97 ();
 sg13g2_fill_2 FILLER_43_101 ();
 sg13g2_decap_4 FILLER_43_106 ();
 sg13g2_fill_2 FILLER_43_110 ();
 sg13g2_fill_2 FILLER_43_121 ();
 sg13g2_fill_1 FILLER_43_123 ();
 sg13g2_decap_4 FILLER_43_143 ();
 sg13g2_decap_8 FILLER_43_152 ();
 sg13g2_fill_2 FILLER_43_159 ();
 sg13g2_fill_1 FILLER_43_161 ();
 sg13g2_fill_1 FILLER_43_177 ();
 sg13g2_fill_1 FILLER_43_187 ();
 sg13g2_fill_1 FILLER_43_193 ();
 sg13g2_decap_8 FILLER_43_225 ();
 sg13g2_decap_8 FILLER_43_232 ();
 sg13g2_decap_8 FILLER_43_239 ();
 sg13g2_decap_4 FILLER_43_246 ();
 sg13g2_decap_8 FILLER_43_253 ();
 sg13g2_fill_2 FILLER_43_260 ();
 sg13g2_decap_4 FILLER_43_268 ();
 sg13g2_fill_1 FILLER_43_272 ();
 sg13g2_decap_8 FILLER_43_278 ();
 sg13g2_fill_2 FILLER_43_285 ();
 sg13g2_fill_1 FILLER_43_302 ();
 sg13g2_fill_1 FILLER_43_340 ();
 sg13g2_fill_1 FILLER_43_382 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_decap_8 FILLER_44_14 ();
 sg13g2_decap_8 FILLER_44_21 ();
 sg13g2_decap_8 FILLER_44_28 ();
 sg13g2_decap_8 FILLER_44_35 ();
 sg13g2_decap_8 FILLER_44_42 ();
 sg13g2_decap_4 FILLER_44_49 ();
 sg13g2_fill_2 FILLER_44_74 ();
 sg13g2_fill_1 FILLER_44_84 ();
 sg13g2_fill_2 FILLER_44_96 ();
 sg13g2_decap_8 FILLER_44_136 ();
 sg13g2_decap_8 FILLER_44_143 ();
 sg13g2_decap_8 FILLER_44_150 ();
 sg13g2_fill_1 FILLER_44_157 ();
 sg13g2_decap_8 FILLER_44_229 ();
 sg13g2_decap_8 FILLER_44_236 ();
 sg13g2_decap_8 FILLER_44_246 ();
 sg13g2_fill_2 FILLER_44_253 ();
 sg13g2_decap_8 FILLER_44_290 ();
 sg13g2_fill_1 FILLER_44_297 ();
 sg13g2_fill_2 FILLER_44_306 ();
 sg13g2_fill_2 FILLER_44_313 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_7 ();
 sg13g2_decap_8 FILLER_45_14 ();
 sg13g2_decap_8 FILLER_45_21 ();
 sg13g2_decap_8 FILLER_45_28 ();
 sg13g2_decap_4 FILLER_45_35 ();
 sg13g2_fill_1 FILLER_45_39 ();
 sg13g2_fill_2 FILLER_45_100 ();
 sg13g2_fill_2 FILLER_45_105 ();
 sg13g2_decap_8 FILLER_45_117 ();
 sg13g2_decap_8 FILLER_45_127 ();
 sg13g2_decap_8 FILLER_45_134 ();
 sg13g2_decap_8 FILLER_45_141 ();
 sg13g2_fill_1 FILLER_45_148 ();
 sg13g2_fill_2 FILLER_45_154 ();
 sg13g2_fill_1 FILLER_45_156 ();
 sg13g2_decap_4 FILLER_45_160 ();
 sg13g2_decap_4 FILLER_45_178 ();
 sg13g2_fill_1 FILLER_45_182 ();
 sg13g2_decap_4 FILLER_45_188 ();
 sg13g2_fill_1 FILLER_45_192 ();
 sg13g2_decap_8 FILLER_45_218 ();
 sg13g2_fill_2 FILLER_45_225 ();
 sg13g2_decap_4 FILLER_45_279 ();
 sg13g2_fill_2 FILLER_45_283 ();
 sg13g2_decap_4 FILLER_45_299 ();
 sg13g2_fill_1 FILLER_45_303 ();
 sg13g2_decap_4 FILLER_45_309 ();
 sg13g2_fill_1 FILLER_45_313 ();
 sg13g2_fill_1 FILLER_45_318 ();
 sg13g2_decap_4 FILLER_45_337 ();
 sg13g2_fill_2 FILLER_45_341 ();
 sg13g2_fill_1 FILLER_45_352 ();
 sg13g2_fill_2 FILLER_45_379 ();
 sg13g2_decap_4 FILLER_45_403 ();
 sg13g2_fill_2 FILLER_45_407 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_7 ();
 sg13g2_decap_8 FILLER_46_14 ();
 sg13g2_decap_8 FILLER_46_21 ();
 sg13g2_decap_8 FILLER_46_28 ();
 sg13g2_fill_1 FILLER_46_35 ();
 sg13g2_fill_1 FILLER_46_76 ();
 sg13g2_fill_1 FILLER_46_110 ();
 sg13g2_fill_1 FILLER_46_116 ();
 sg13g2_decap_8 FILLER_46_122 ();
 sg13g2_decap_8 FILLER_46_129 ();
 sg13g2_fill_1 FILLER_46_136 ();
 sg13g2_decap_8 FILLER_46_174 ();
 sg13g2_decap_8 FILLER_46_181 ();
 sg13g2_decap_8 FILLER_46_188 ();
 sg13g2_decap_8 FILLER_46_195 ();
 sg13g2_decap_8 FILLER_46_202 ();
 sg13g2_fill_2 FILLER_46_209 ();
 sg13g2_fill_1 FILLER_46_263 ();
 sg13g2_fill_2 FILLER_46_267 ();
 sg13g2_fill_1 FILLER_46_269 ();
 sg13g2_decap_8 FILLER_46_309 ();
 sg13g2_decap_8 FILLER_46_316 ();
 sg13g2_decap_8 FILLER_46_323 ();
 sg13g2_fill_2 FILLER_46_330 ();
 sg13g2_fill_1 FILLER_46_332 ();
 sg13g2_fill_2 FILLER_46_362 ();
 sg13g2_fill_2 FILLER_46_376 ();
 sg13g2_fill_1 FILLER_46_384 ();
 sg13g2_fill_1 FILLER_46_389 ();
 sg13g2_decap_4 FILLER_46_393 ();
 sg13g2_fill_1 FILLER_46_397 ();
 sg13g2_fill_2 FILLER_46_406 ();
 sg13g2_fill_1 FILLER_46_408 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_7 ();
 sg13g2_decap_8 FILLER_47_14 ();
 sg13g2_decap_8 FILLER_47_21 ();
 sg13g2_fill_1 FILLER_47_28 ();
 sg13g2_fill_1 FILLER_47_55 ();
 sg13g2_fill_2 FILLER_47_61 ();
 sg13g2_fill_1 FILLER_47_63 ();
 sg13g2_fill_2 FILLER_47_103 ();
 sg13g2_fill_2 FILLER_47_186 ();
 sg13g2_fill_1 FILLER_47_191 ();
 sg13g2_decap_8 FILLER_47_195 ();
 sg13g2_decap_8 FILLER_47_202 ();
 sg13g2_fill_1 FILLER_47_252 ();
 sg13g2_decap_4 FILLER_47_321 ();
 sg13g2_fill_1 FILLER_47_345 ();
 sg13g2_fill_2 FILLER_47_372 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_decap_8 FILLER_48_14 ();
 sg13g2_decap_8 FILLER_48_21 ();
 sg13g2_fill_2 FILLER_48_28 ();
 sg13g2_fill_1 FILLER_48_30 ();
 sg13g2_decap_8 FILLER_48_46 ();
 sg13g2_fill_2 FILLER_48_53 ();
 sg13g2_fill_2 FILLER_48_68 ();
 sg13g2_fill_1 FILLER_48_70 ();
 sg13g2_fill_1 FILLER_48_97 ();
 sg13g2_fill_1 FILLER_48_157 ();
 sg13g2_decap_4 FILLER_48_242 ();
 sg13g2_fill_2 FILLER_48_253 ();
 sg13g2_fill_1 FILLER_48_255 ();
 sg13g2_fill_2 FILLER_48_270 ();
 sg13g2_fill_2 FILLER_48_309 ();
 sg13g2_fill_1 FILLER_48_311 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_7 ();
 sg13g2_decap_8 FILLER_49_14 ();
 sg13g2_fill_2 FILLER_49_21 ();
 sg13g2_fill_1 FILLER_49_68 ();
 sg13g2_decap_8 FILLER_49_83 ();
 sg13g2_fill_1 FILLER_49_90 ();
 sg13g2_fill_2 FILLER_49_100 ();
 sg13g2_fill_1 FILLER_49_102 ();
 sg13g2_fill_2 FILLER_49_114 ();
 sg13g2_fill_1 FILLER_49_116 ();
 sg13g2_fill_2 FILLER_49_145 ();
 sg13g2_fill_1 FILLER_49_181 ();
 sg13g2_decap_8 FILLER_49_246 ();
 sg13g2_decap_8 FILLER_49_253 ();
 sg13g2_decap_4 FILLER_49_263 ();
 sg13g2_fill_2 FILLER_49_281 ();
 sg13g2_fill_1 FILLER_49_301 ();
 sg13g2_fill_1 FILLER_49_325 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_8 FILLER_50_7 ();
 sg13g2_decap_4 FILLER_50_14 ();
 sg13g2_fill_1 FILLER_50_18 ();
 sg13g2_fill_1 FILLER_50_100 ();
 sg13g2_decap_8 FILLER_50_129 ();
 sg13g2_fill_1 FILLER_50_136 ();
 sg13g2_decap_4 FILLER_50_211 ();
 sg13g2_decap_4 FILLER_50_226 ();
 sg13g2_fill_1 FILLER_50_230 ();
 sg13g2_fill_2 FILLER_50_298 ();
 sg13g2_fill_1 FILLER_50_300 ();
 sg13g2_fill_1 FILLER_50_340 ();
 sg13g2_fill_1 FILLER_50_408 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_decap_8 FILLER_51_7 ();
 sg13g2_decap_8 FILLER_51_14 ();
 sg13g2_fill_2 FILLER_51_21 ();
 sg13g2_fill_1 FILLER_51_23 ();
 sg13g2_fill_1 FILLER_51_65 ();
 sg13g2_fill_2 FILLER_51_79 ();
 sg13g2_fill_1 FILLER_51_81 ();
 sg13g2_fill_1 FILLER_51_127 ();
 sg13g2_fill_1 FILLER_51_133 ();
 sg13g2_decap_4 FILLER_51_139 ();
 sg13g2_decap_4 FILLER_51_191 ();
 sg13g2_fill_1 FILLER_51_195 ();
 sg13g2_decap_8 FILLER_51_275 ();
 sg13g2_fill_2 FILLER_51_282 ();
 sg13g2_fill_1 FILLER_51_284 ();
 sg13g2_fill_2 FILLER_51_290 ();
 sg13g2_fill_1 FILLER_51_326 ();
 sg13g2_fill_1 FILLER_51_408 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_decap_8 FILLER_52_7 ();
 sg13g2_decap_8 FILLER_52_14 ();
 sg13g2_decap_8 FILLER_52_21 ();
 sg13g2_fill_2 FILLER_52_28 ();
 sg13g2_fill_2 FILLER_52_38 ();
 sg13g2_fill_1 FILLER_52_49 ();
 sg13g2_fill_2 FILLER_52_77 ();
 sg13g2_fill_1 FILLER_52_118 ();
 sg13g2_fill_1 FILLER_52_164 ();
 sg13g2_decap_8 FILLER_52_170 ();
 sg13g2_fill_2 FILLER_52_177 ();
 sg13g2_fill_1 FILLER_52_179 ();
 sg13g2_decap_4 FILLER_52_183 ();
 sg13g2_fill_1 FILLER_52_213 ();
 sg13g2_fill_1 FILLER_52_229 ();
 sg13g2_decap_8 FILLER_52_233 ();
 sg13g2_fill_2 FILLER_52_264 ();
 sg13g2_fill_1 FILLER_52_266 ();
 sg13g2_fill_2 FILLER_52_290 ();
 sg13g2_fill_1 FILLER_52_292 ();
 sg13g2_fill_2 FILLER_52_319 ();
 sg13g2_fill_2 FILLER_52_372 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_decap_8 FILLER_53_7 ();
 sg13g2_decap_8 FILLER_53_14 ();
 sg13g2_decap_4 FILLER_53_21 ();
 sg13g2_fill_1 FILLER_53_25 ();
 sg13g2_fill_1 FILLER_53_78 ();
 sg13g2_fill_2 FILLER_53_117 ();
 sg13g2_fill_1 FILLER_53_141 ();
 sg13g2_fill_2 FILLER_53_148 ();
 sg13g2_decap_8 FILLER_53_160 ();
 sg13g2_decap_4 FILLER_53_167 ();
 sg13g2_fill_2 FILLER_53_171 ();
 sg13g2_decap_4 FILLER_53_239 ();
 sg13g2_fill_2 FILLER_53_251 ();
 sg13g2_fill_1 FILLER_53_330 ();
 sg13g2_fill_1 FILLER_53_362 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_decap_8 FILLER_54_7 ();
 sg13g2_fill_2 FILLER_54_14 ();
 sg13g2_fill_1 FILLER_54_16 ();
 sg13g2_fill_1 FILLER_54_52 ();
 sg13g2_fill_2 FILLER_54_68 ();
 sg13g2_fill_1 FILLER_54_70 ();
 sg13g2_fill_2 FILLER_54_89 ();
 sg13g2_fill_2 FILLER_54_100 ();
 sg13g2_fill_1 FILLER_54_126 ();
 sg13g2_fill_2 FILLER_54_131 ();
 sg13g2_fill_2 FILLER_54_144 ();
 sg13g2_fill_2 FILLER_54_160 ();
 sg13g2_fill_1 FILLER_54_195 ();
 sg13g2_decap_4 FILLER_54_209 ();
 sg13g2_decap_8 FILLER_54_260 ();
 sg13g2_decap_8 FILLER_54_267 ();
 sg13g2_fill_1 FILLER_54_279 ();
 sg13g2_fill_2 FILLER_54_298 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_decap_8 FILLER_55_7 ();
 sg13g2_decap_8 FILLER_55_14 ();
 sg13g2_fill_1 FILLER_55_21 ();
 sg13g2_fill_1 FILLER_55_48 ();
 sg13g2_fill_2 FILLER_55_148 ();
 sg13g2_fill_2 FILLER_55_162 ();
 sg13g2_fill_1 FILLER_55_169 ();
 sg13g2_fill_1 FILLER_55_192 ();
 sg13g2_fill_1 FILLER_55_202 ();
 sg13g2_decap_8 FILLER_55_268 ();
 sg13g2_decap_8 FILLER_55_275 ();
 sg13g2_fill_1 FILLER_55_292 ();
 sg13g2_fill_2 FILLER_55_298 ();
 sg13g2_decap_4 FILLER_55_314 ();
 sg13g2_fill_1 FILLER_55_318 ();
 sg13g2_fill_2 FILLER_55_339 ();
 sg13g2_fill_1 FILLER_55_386 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_decap_8 FILLER_56_7 ();
 sg13g2_decap_8 FILLER_56_14 ();
 sg13g2_fill_2 FILLER_56_21 ();
 sg13g2_fill_1 FILLER_56_23 ();
 sg13g2_fill_2 FILLER_56_65 ();
 sg13g2_fill_1 FILLER_56_67 ();
 sg13g2_fill_2 FILLER_56_73 ();
 sg13g2_fill_1 FILLER_56_75 ();
 sg13g2_fill_1 FILLER_56_150 ();
 sg13g2_fill_2 FILLER_56_157 ();
 sg13g2_fill_2 FILLER_56_213 ();
 sg13g2_fill_2 FILLER_56_222 ();
 sg13g2_fill_1 FILLER_56_292 ();
 sg13g2_fill_2 FILLER_56_321 ();
 sg13g2_fill_1 FILLER_56_323 ();
 sg13g2_fill_1 FILLER_56_371 ();
 sg13g2_fill_2 FILLER_56_385 ();
 sg13g2_fill_1 FILLER_56_396 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_decap_8 FILLER_57_7 ();
 sg13g2_decap_4 FILLER_57_14 ();
 sg13g2_fill_2 FILLER_57_18 ();
 sg13g2_fill_1 FILLER_57_42 ();
 sg13g2_fill_2 FILLER_57_66 ();
 sg13g2_decap_4 FILLER_57_77 ();
 sg13g2_fill_2 FILLER_57_81 ();
 sg13g2_fill_1 FILLER_57_86 ();
 sg13g2_fill_1 FILLER_57_92 ();
 sg13g2_decap_8 FILLER_57_96 ();
 sg13g2_fill_2 FILLER_57_131 ();
 sg13g2_fill_2 FILLER_57_164 ();
 sg13g2_fill_2 FILLER_57_169 ();
 sg13g2_fill_1 FILLER_57_171 ();
 sg13g2_fill_2 FILLER_57_200 ();
 sg13g2_fill_2 FILLER_57_215 ();
 sg13g2_fill_1 FILLER_57_217 ();
 sg13g2_fill_2 FILLER_57_295 ();
 sg13g2_fill_1 FILLER_57_297 ();
 sg13g2_fill_1 FILLER_57_315 ();
 sg13g2_fill_1 FILLER_57_368 ();
 sg13g2_fill_1 FILLER_57_375 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_decap_8 FILLER_58_7 ();
 sg13g2_decap_8 FILLER_58_14 ();
 sg13g2_fill_2 FILLER_58_21 ();
 sg13g2_fill_1 FILLER_58_140 ();
 sg13g2_fill_2 FILLER_58_202 ();
 sg13g2_fill_1 FILLER_58_204 ();
 sg13g2_decap_8 FILLER_58_219 ();
 sg13g2_fill_1 FILLER_58_226 ();
 sg13g2_fill_2 FILLER_58_231 ();
 sg13g2_decap_8 FILLER_58_241 ();
 sg13g2_decap_4 FILLER_58_248 ();
 sg13g2_fill_2 FILLER_58_252 ();
 sg13g2_fill_1 FILLER_58_355 ();
 sg13g2_fill_1 FILLER_58_408 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_decap_8 FILLER_59_7 ();
 sg13g2_decap_8 FILLER_59_14 ();
 sg13g2_fill_2 FILLER_59_21 ();
 sg13g2_fill_1 FILLER_59_49 ();
 sg13g2_fill_1 FILLER_59_72 ();
 sg13g2_decap_8 FILLER_59_95 ();
 sg13g2_decap_8 FILLER_59_102 ();
 sg13g2_fill_1 FILLER_59_109 ();
 sg13g2_fill_1 FILLER_59_139 ();
 sg13g2_fill_1 FILLER_59_168 ();
 sg13g2_decap_4 FILLER_59_172 ();
 sg13g2_fill_2 FILLER_59_176 ();
 sg13g2_fill_1 FILLER_59_200 ();
 sg13g2_fill_1 FILLER_59_231 ();
 sg13g2_decap_8 FILLER_59_242 ();
 sg13g2_decap_4 FILLER_59_249 ();
 sg13g2_fill_2 FILLER_59_253 ();
 sg13g2_fill_1 FILLER_59_260 ();
 sg13g2_fill_1 FILLER_59_264 ();
 sg13g2_fill_2 FILLER_59_308 ();
 sg13g2_fill_2 FILLER_59_319 ();
 sg13g2_fill_1 FILLER_59_331 ();
 sg13g2_fill_1 FILLER_59_351 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_decap_8 FILLER_60_7 ();
 sg13g2_decap_8 FILLER_60_14 ();
 sg13g2_decap_4 FILLER_60_21 ();
 sg13g2_fill_2 FILLER_60_42 ();
 sg13g2_fill_1 FILLER_60_44 ();
 sg13g2_decap_8 FILLER_60_109 ();
 sg13g2_decap_8 FILLER_60_116 ();
 sg13g2_fill_1 FILLER_60_123 ();
 sg13g2_decap_4 FILLER_60_129 ();
 sg13g2_decap_8 FILLER_60_138 ();
 sg13g2_decap_8 FILLER_60_145 ();
 sg13g2_decap_8 FILLER_60_152 ();
 sg13g2_fill_2 FILLER_60_188 ();
 sg13g2_fill_1 FILLER_60_190 ();
 sg13g2_decap_4 FILLER_60_264 ();
 sg13g2_fill_2 FILLER_60_284 ();
 sg13g2_fill_2 FILLER_60_296 ();
 sg13g2_fill_1 FILLER_60_329 ();
 sg13g2_fill_1 FILLER_60_385 ();
 sg13g2_decap_4 FILLER_60_404 ();
 sg13g2_fill_1 FILLER_60_408 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_decap_8 FILLER_61_7 ();
 sg13g2_decap_8 FILLER_61_14 ();
 sg13g2_decap_8 FILLER_61_21 ();
 sg13g2_decap_4 FILLER_61_28 ();
 sg13g2_fill_1 FILLER_61_32 ();
 sg13g2_fill_1 FILLER_61_116 ();
 sg13g2_decap_4 FILLER_61_122 ();
 sg13g2_fill_1 FILLER_61_126 ();
 sg13g2_fill_2 FILLER_61_140 ();
 sg13g2_fill_1 FILLER_61_207 ();
 sg13g2_fill_1 FILLER_61_218 ();
 sg13g2_fill_2 FILLER_61_284 ();
 sg13g2_fill_1 FILLER_61_286 ();
 sg13g2_fill_1 FILLER_61_319 ();
 sg13g2_fill_2 FILLER_61_367 ();
 sg13g2_fill_1 FILLER_61_386 ();
 sg13g2_fill_1 FILLER_61_390 ();
 sg13g2_fill_2 FILLER_61_394 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_decap_8 FILLER_62_7 ();
 sg13g2_decap_8 FILLER_62_14 ();
 sg13g2_decap_8 FILLER_62_21 ();
 sg13g2_fill_2 FILLER_62_28 ();
 sg13g2_fill_1 FILLER_62_30 ();
 sg13g2_fill_1 FILLER_62_83 ();
 sg13g2_fill_2 FILLER_62_184 ();
 sg13g2_fill_2 FILLER_62_235 ();
 sg13g2_fill_1 FILLER_62_339 ();
 sg13g2_fill_1 FILLER_62_383 ();
 sg13g2_fill_1 FILLER_62_399 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_decap_8 FILLER_63_7 ();
 sg13g2_decap_8 FILLER_63_14 ();
 sg13g2_decap_8 FILLER_63_21 ();
 sg13g2_fill_1 FILLER_63_58 ();
 sg13g2_fill_2 FILLER_63_144 ();
 sg13g2_fill_1 FILLER_63_163 ();
 sg13g2_fill_2 FILLER_63_247 ();
 sg13g2_fill_1 FILLER_63_278 ();
 sg13g2_fill_1 FILLER_63_372 ();
 sg13g2_fill_1 FILLER_63_382 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_8 FILLER_64_7 ();
 sg13g2_decap_8 FILLER_64_14 ();
 sg13g2_fill_1 FILLER_64_48 ();
 sg13g2_fill_1 FILLER_64_96 ();
 sg13g2_fill_2 FILLER_64_111 ();
 sg13g2_fill_1 FILLER_64_123 ();
 sg13g2_fill_1 FILLER_64_132 ();
 sg13g2_fill_2 FILLER_64_137 ();
 sg13g2_fill_2 FILLER_64_180 ();
 sg13g2_fill_1 FILLER_64_258 ();
 sg13g2_fill_1 FILLER_64_408 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_8 FILLER_65_7 ();
 sg13g2_decap_8 FILLER_65_14 ();
 sg13g2_fill_1 FILLER_65_21 ();
 sg13g2_fill_1 FILLER_65_43 ();
 sg13g2_fill_2 FILLER_65_120 ();
 sg13g2_fill_2 FILLER_65_145 ();
 sg13g2_fill_1 FILLER_65_201 ();
 sg13g2_fill_1 FILLER_65_211 ();
 sg13g2_decap_8 FILLER_65_277 ();
 sg13g2_decap_4 FILLER_65_284 ();
 sg13g2_fill_2 FILLER_65_288 ();
 sg13g2_fill_2 FILLER_65_314 ();
 sg13g2_fill_2 FILLER_65_331 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_8 FILLER_66_7 ();
 sg13g2_decap_8 FILLER_66_14 ();
 sg13g2_fill_2 FILLER_66_21 ();
 sg13g2_fill_1 FILLER_66_80 ();
 sg13g2_fill_1 FILLER_66_133 ();
 sg13g2_fill_1 FILLER_66_142 ();
 sg13g2_fill_2 FILLER_66_155 ();
 sg13g2_fill_2 FILLER_66_193 ();
 sg13g2_decap_8 FILLER_66_223 ();
 sg13g2_fill_2 FILLER_66_230 ();
 sg13g2_decap_8 FILLER_66_286 ();
 sg13g2_fill_1 FILLER_66_293 ();
 sg13g2_fill_1 FILLER_66_300 ();
 sg13g2_fill_2 FILLER_66_314 ();
 sg13g2_decap_8 FILLER_66_328 ();
 sg13g2_decap_4 FILLER_66_335 ();
 sg13g2_fill_2 FILLER_66_339 ();
 sg13g2_fill_1 FILLER_66_349 ();
 sg13g2_fill_1 FILLER_66_377 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_8 FILLER_67_7 ();
 sg13g2_decap_8 FILLER_67_14 ();
 sg13g2_decap_8 FILLER_67_21 ();
 sg13g2_decap_4 FILLER_67_28 ();
 sg13g2_fill_2 FILLER_67_118 ();
 sg13g2_fill_2 FILLER_67_126 ();
 sg13g2_fill_2 FILLER_67_151 ();
 sg13g2_fill_1 FILLER_67_162 ();
 sg13g2_fill_2 FILLER_67_177 ();
 sg13g2_decap_4 FILLER_67_218 ();
 sg13g2_fill_1 FILLER_67_222 ();
 sg13g2_fill_2 FILLER_67_244 ();
 sg13g2_fill_1 FILLER_67_298 ();
 sg13g2_fill_1 FILLER_67_397 ();
 sg13g2_fill_2 FILLER_67_407 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_8 FILLER_68_7 ();
 sg13g2_decap_8 FILLER_68_14 ();
 sg13g2_decap_4 FILLER_68_21 ();
 sg13g2_fill_1 FILLER_68_60 ();
 sg13g2_fill_1 FILLER_68_87 ();
 sg13g2_decap_4 FILLER_68_198 ();
 sg13g2_fill_1 FILLER_68_202 ();
 sg13g2_fill_1 FILLER_68_206 ();
 sg13g2_decap_8 FILLER_68_210 ();
 sg13g2_decap_4 FILLER_68_217 ();
 sg13g2_fill_1 FILLER_68_260 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_8 FILLER_69_7 ();
 sg13g2_decap_4 FILLER_69_14 ();
 sg13g2_fill_2 FILLER_69_18 ();
 sg13g2_fill_1 FILLER_69_62 ();
 sg13g2_fill_2 FILLER_69_145 ();
 sg13g2_decap_4 FILLER_69_164 ();
 sg13g2_fill_1 FILLER_69_168 ();
 sg13g2_fill_1 FILLER_69_206 ();
 sg13g2_fill_1 FILLER_69_212 ();
 sg13g2_fill_1 FILLER_69_257 ();
 sg13g2_fill_2 FILLER_69_347 ();
 sg13g2_fill_1 FILLER_69_349 ();
 sg13g2_fill_1 FILLER_69_366 ();
 sg13g2_fill_2 FILLER_69_372 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_decap_8 FILLER_70_14 ();
 sg13g2_decap_4 FILLER_70_21 ();
 sg13g2_fill_2 FILLER_70_93 ();
 sg13g2_fill_1 FILLER_70_100 ();
 sg13g2_fill_1 FILLER_70_124 ();
 sg13g2_decap_4 FILLER_70_158 ();
 sg13g2_fill_1 FILLER_70_162 ();
 sg13g2_decap_4 FILLER_70_170 ();
 sg13g2_fill_2 FILLER_70_174 ();
 sg13g2_fill_2 FILLER_70_216 ();
 sg13g2_fill_2 FILLER_70_296 ();
 sg13g2_decap_8 FILLER_70_338 ();
 sg13g2_decap_4 FILLER_70_345 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_decap_8 FILLER_71_7 ();
 sg13g2_decap_8 FILLER_71_14 ();
 sg13g2_fill_2 FILLER_71_21 ();
 sg13g2_fill_1 FILLER_71_72 ();
 sg13g2_fill_1 FILLER_71_181 ();
 sg13g2_fill_1 FILLER_71_324 ();
 sg13g2_fill_2 FILLER_71_334 ();
 sg13g2_fill_2 FILLER_71_346 ();
 sg13g2_fill_1 FILLER_71_348 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_decap_8 FILLER_72_14 ();
 sg13g2_decap_8 FILLER_72_21 ();
 sg13g2_fill_1 FILLER_72_28 ();
 sg13g2_fill_2 FILLER_72_128 ();
 sg13g2_fill_2 FILLER_72_210 ();
 sg13g2_fill_1 FILLER_72_396 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_decap_8 FILLER_73_14 ();
 sg13g2_decap_8 FILLER_73_21 ();
 sg13g2_decap_4 FILLER_73_28 ();
 sg13g2_fill_2 FILLER_73_75 ();
 sg13g2_fill_2 FILLER_73_97 ();
 sg13g2_fill_1 FILLER_73_182 ();
 sg13g2_fill_1 FILLER_73_247 ();
 sg13g2_fill_2 FILLER_73_329 ();
 sg13g2_fill_2 FILLER_73_335 ();
 sg13g2_fill_2 FILLER_73_354 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_decap_8 FILLER_74_14 ();
 sg13g2_decap_8 FILLER_74_21 ();
 sg13g2_decap_8 FILLER_74_28 ();
 sg13g2_decap_8 FILLER_74_35 ();
 sg13g2_fill_1 FILLER_74_68 ();
 sg13g2_fill_2 FILLER_74_78 ();
 sg13g2_fill_2 FILLER_74_110 ();
 sg13g2_fill_1 FILLER_74_194 ();
 sg13g2_decap_4 FILLER_74_199 ();
 sg13g2_fill_2 FILLER_74_203 ();
 sg13g2_decap_8 FILLER_74_209 ();
 sg13g2_decap_8 FILLER_74_220 ();
 sg13g2_fill_1 FILLER_74_230 ();
 sg13g2_fill_2 FILLER_74_261 ();
 sg13g2_fill_1 FILLER_74_330 ();
 sg13g2_fill_1 FILLER_74_382 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_14 ();
 sg13g2_decap_8 FILLER_75_21 ();
 sg13g2_decap_8 FILLER_75_28 ();
 sg13g2_decap_8 FILLER_75_35 ();
 sg13g2_decap_8 FILLER_75_42 ();
 sg13g2_decap_4 FILLER_75_49 ();
 sg13g2_fill_2 FILLER_75_53 ();
 sg13g2_fill_2 FILLER_75_65 ();
 sg13g2_fill_1 FILLER_75_67 ();
 sg13g2_fill_2 FILLER_75_110 ();
 sg13g2_fill_2 FILLER_75_136 ();
 sg13g2_fill_2 FILLER_75_152 ();
 sg13g2_decap_8 FILLER_75_190 ();
 sg13g2_decap_4 FILLER_75_197 ();
 sg13g2_fill_1 FILLER_75_220 ();
 sg13g2_fill_1 FILLER_75_251 ();
 sg13g2_fill_1 FILLER_75_355 ();
 sg13g2_fill_2 FILLER_75_363 ();
 sg13g2_fill_1 FILLER_75_374 ();
 sg13g2_fill_1 FILLER_75_396 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_8 FILLER_76_21 ();
 sg13g2_decap_8 FILLER_76_28 ();
 sg13g2_decap_8 FILLER_76_35 ();
 sg13g2_decap_8 FILLER_76_42 ();
 sg13g2_decap_8 FILLER_76_49 ();
 sg13g2_decap_8 FILLER_76_56 ();
 sg13g2_decap_8 FILLER_76_63 ();
 sg13g2_fill_2 FILLER_76_70 ();
 sg13g2_fill_1 FILLER_76_72 ();
 sg13g2_fill_1 FILLER_76_108 ();
 sg13g2_fill_1 FILLER_76_179 ();
 sg13g2_fill_1 FILLER_76_194 ();
 sg13g2_fill_1 FILLER_76_199 ();
 sg13g2_fill_2 FILLER_76_270 ();
 sg13g2_decap_8 FILLER_76_308 ();
 sg13g2_fill_2 FILLER_76_315 ();
 sg13g2_fill_1 FILLER_76_323 ();
 sg13g2_fill_1 FILLER_76_386 ();
 sg13g2_fill_1 FILLER_76_399 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_decap_8 FILLER_77_28 ();
 sg13g2_decap_8 FILLER_77_35 ();
 sg13g2_decap_8 FILLER_77_42 ();
 sg13g2_decap_8 FILLER_77_49 ();
 sg13g2_decap_8 FILLER_77_56 ();
 sg13g2_decap_8 FILLER_77_63 ();
 sg13g2_decap_8 FILLER_77_70 ();
 sg13g2_fill_1 FILLER_77_151 ();
 sg13g2_fill_1 FILLER_77_161 ();
 sg13g2_fill_2 FILLER_77_197 ();
 sg13g2_fill_1 FILLER_77_199 ();
 sg13g2_fill_2 FILLER_77_206 ();
 sg13g2_fill_1 FILLER_77_208 ();
 sg13g2_fill_1 FILLER_77_226 ();
 sg13g2_fill_2 FILLER_77_307 ();
 sg13g2_fill_1 FILLER_77_335 ();
 sg13g2_fill_1 FILLER_77_408 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_decap_8 FILLER_78_28 ();
 sg13g2_decap_8 FILLER_78_35 ();
 sg13g2_decap_8 FILLER_78_42 ();
 sg13g2_decap_8 FILLER_78_49 ();
 sg13g2_decap_8 FILLER_78_56 ();
 sg13g2_decap_8 FILLER_78_63 ();
 sg13g2_fill_1 FILLER_78_70 ();
 sg13g2_fill_1 FILLER_78_97 ();
 sg13g2_fill_2 FILLER_78_210 ();
 sg13g2_fill_1 FILLER_78_252 ();
 sg13g2_fill_1 FILLER_78_296 ();
 sg13g2_decap_4 FILLER_78_306 ();
 sg13g2_fill_2 FILLER_78_390 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_decap_8 FILLER_79_35 ();
 sg13g2_decap_8 FILLER_79_42 ();
 sg13g2_decap_8 FILLER_79_49 ();
 sg13g2_decap_8 FILLER_79_56 ();
 sg13g2_fill_1 FILLER_79_63 ();
 sg13g2_fill_2 FILLER_79_125 ();
 sg13g2_fill_1 FILLER_79_188 ();
 sg13g2_fill_2 FILLER_79_247 ();
 sg13g2_fill_1 FILLER_79_275 ();
 sg13g2_decap_8 FILLER_79_301 ();
 sg13g2_decap_8 FILLER_79_308 ();
 sg13g2_decap_8 FILLER_79_315 ();
 sg13g2_fill_2 FILLER_79_322 ();
 sg13g2_fill_2 FILLER_79_407 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_42 ();
 sg13g2_decap_8 FILLER_80_49 ();
 sg13g2_decap_4 FILLER_80_60 ();
 sg13g2_fill_2 FILLER_80_108 ();
 sg13g2_fill_2 FILLER_80_174 ();
 sg13g2_decap_4 FILLER_80_192 ();
 sg13g2_fill_1 FILLER_80_217 ();
 sg13g2_fill_2 FILLER_80_231 ();
 sg13g2_fill_1 FILLER_80_237 ();
 sg13g2_decap_8 FILLER_80_293 ();
 sg13g2_decap_8 FILLER_80_300 ();
 sg13g2_decap_8 FILLER_80_307 ();
 sg13g2_decap_8 FILLER_80_314 ();
 sg13g2_decap_4 FILLER_80_321 ();
 sg13g2_fill_1 FILLER_80_325 ();
 sg13g2_fill_2 FILLER_80_341 ();
 sg13g2_fill_1 FILLER_80_343 ();
 sg13g2_decap_4 FILLER_80_405 ();
 assign uio_oe[0] = net3;
 assign uio_oe[1] = net4;
 assign uio_oe[2] = net5;
 assign uio_oe[3] = net6;
 assign uio_oe[4] = net7;
 assign uio_oe[5] = net8;
 assign uio_oe[6] = net9;
 assign uio_oe[7] = net10;
 assign uio_out[0] = net11;
 assign uio_out[1] = net12;
 assign uio_out[2] = net13;
 assign uio_out[3] = net14;
 assign uio_out[4] = net15;
 assign uio_out[5] = net16;
 assign uio_out[6] = net17;
 assign uio_out[7] = net18;
endmodule

module tt_um_kentrane_tinyspectrum (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire _297_;
 wire _298_;
 wire _299_;
 wire _300_;
 wire _301_;
 wire _302_;
 wire _303_;
 wire _304_;
 wire _305_;
 wire _306_;
 wire _307_;
 wire _308_;
 wire _309_;
 wire \counter[0] ;
 wire \counter[10] ;
 wire \counter[11] ;
 wire \counter[12] ;
 wire \counter[13] ;
 wire \counter[14] ;
 wire \counter[15] ;
 wire \counter[16] ;
 wire \counter[17] ;
 wire \counter[18] ;
 wire \counter[19] ;
 wire \counter[1] ;
 wire \counter[2] ;
 wire \counter[3] ;
 wire \counter[4] ;
 wire \counter[5] ;
 wire \counter[6] ;
 wire \counter[7] ;
 wire \counter[8] ;
 wire \counter[9] ;
 wire tone_out;
 wire \tremolo_counter[0] ;
 wire \tremolo_counter[1] ;
 wire \tremolo_counter[2] ;
 wire \tremolo_counter[3] ;
 wire \tremolo_counter[4] ;
 wire \tremolo_counter[5] ;
 wire \tremolo_counter[6] ;
 wire \tremolo_counter[7] ;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire clknet_0_clk;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;

 sg13g2_inv_1 _310_ (.Y(_287_),
    .A(net102));
 sg13g2_inv_1 _311_ (.Y(_288_),
    .A(net103));
 sg13g2_inv_2 _312_ (.Y(_289_),
    .A(net96));
 sg13g2_inv_1 _313_ (.Y(_290_),
    .A(net57));
 sg13g2_inv_1 _314_ (.Y(_291_),
    .A(_005_));
 sg13g2_inv_2 _315_ (.Y(_292_),
    .A(net43));
 sg13g2_inv_1 _316_ (.Y(_293_),
    .A(_013_));
 sg13g2_inv_1 _317_ (.Y(_294_),
    .A(net41));
 sg13g2_and2_2 _318_ (.A(net100),
    .B(net98),
    .X(_295_));
 sg13g2_nand2_1 _319_ (.Y(_044_),
    .A(net101),
    .B(net98));
 sg13g2_nor2b_2 _320_ (.A(net104),
    .B_N(net105),
    .Y(_045_));
 sg13g2_nand2b_2 _321_ (.Y(_046_),
    .B(net106),
    .A_N(net103));
 sg13g2_nor2b_2 _322_ (.A(net101),
    .B_N(net98),
    .Y(_047_));
 sg13g2_and2_1 _323_ (.A(net105),
    .B(net103),
    .X(_048_));
 sg13g2_nand2_2 _324_ (.Y(_049_),
    .A(net106),
    .B(net103));
 sg13g2_a22oi_1 _325_ (.Y(_050_),
    .B1(_047_),
    .B2(_048_),
    .A2(_045_),
    .A1(_295_));
 sg13g2_nor2_1 _326_ (.A(net105),
    .B(net103),
    .Y(_051_));
 sg13g2_nor3_2 _327_ (.A(net99),
    .B(net106),
    .C(net104),
    .Y(_052_));
 sg13g2_nor2_1 _328_ (.A(net100),
    .B(net97),
    .Y(_053_));
 sg13g2_or2_2 _329_ (.X(_054_),
    .B(net97),
    .A(net100));
 sg13g2_o21ai_1 _330_ (.B1(net93),
    .Y(_055_),
    .A1(_046_),
    .A2(_054_));
 sg13g2_a21oi_1 _331_ (.A1(net100),
    .A2(_052_),
    .Y(_056_),
    .B1(_055_));
 sg13g2_and2_1 _332_ (.A(_050_),
    .B(_056_),
    .X(uo_out[0]));
 sg13g2_nor2_1 _333_ (.A(net100),
    .B(net105),
    .Y(_057_));
 sg13g2_nor2_1 _334_ (.A(_045_),
    .B(_057_),
    .Y(_058_));
 sg13g2_nor2b_2 _335_ (.A(net97),
    .B_N(net100),
    .Y(_059_));
 sg13g2_nand2b_1 _336_ (.Y(_060_),
    .B(net100),
    .A_N(net97));
 sg13g2_nor2b_2 _337_ (.A(net105),
    .B_N(net103),
    .Y(_061_));
 sg13g2_nand2b_1 _338_ (.Y(_062_),
    .B(net104),
    .A_N(net106));
 sg13g2_o21ai_1 _339_ (.B1(_059_),
    .Y(_063_),
    .A1(_045_),
    .A2(_061_));
 sg13g2_nand2_1 _340_ (.Y(_064_),
    .A(net93),
    .B(_063_));
 sg13g2_a21oi_1 _341_ (.A1(net97),
    .A2(_058_),
    .Y(uo_out[1]),
    .B1(_064_));
 sg13g2_o21ai_1 _342_ (.B1(net93),
    .Y(_065_),
    .A1(_054_),
    .A2(_062_));
 sg13g2_a21oi_1 _343_ (.A1(_295_),
    .A2(_046_),
    .Y(uo_out[2]),
    .B1(_065_));
 sg13g2_xnor2_1 _344_ (.Y(_066_),
    .A(net102),
    .B(net106));
 sg13g2_and3_2 _345_ (.X(_067_),
    .A(net2),
    .B(net104),
    .C(_066_));
 sg13g2_nor3_1 _346_ (.A(_045_),
    .B(_060_),
    .C(_061_),
    .Y(_068_));
 sg13g2_nor3_1 _347_ (.A(_055_),
    .B(_067_),
    .C(_068_),
    .Y(uo_out[3]));
 sg13g2_nor2_1 _348_ (.A(net98),
    .B(_057_),
    .Y(_069_));
 sg13g2_or3_1 _349_ (.A(net98),
    .B(_057_),
    .C(_061_),
    .X(_070_));
 sg13g2_nand2_1 _350_ (.Y(_071_),
    .A(net93),
    .B(_070_));
 sg13g2_a21oi_1 _351_ (.A1(_045_),
    .A2(_047_),
    .Y(uo_out[4]),
    .B1(_071_));
 sg13g2_nand2_1 _352_ (.Y(_072_),
    .A(net101),
    .B(_049_));
 sg13g2_nor2_1 _353_ (.A(net97),
    .B(_051_),
    .Y(_073_));
 sg13g2_o21ai_1 _354_ (.B1(net93),
    .Y(_074_),
    .A1(_044_),
    .A2(_046_));
 sg13g2_a21oi_1 _355_ (.A1(_072_),
    .A2(_073_),
    .Y(uo_out[5]),
    .B1(_074_));
 sg13g2_nor3_2 _356_ (.A(net102),
    .B(net99),
    .C(net104),
    .Y(_075_));
 sg13g2_a21oi_1 _357_ (.A1(net92),
    .A2(_059_),
    .Y(_076_),
    .B1(_075_));
 sg13g2_nand2_1 _358_ (.Y(_077_),
    .A(net93),
    .B(_076_));
 sg13g2_a21oi_2 _359_ (.B1(_077_),
    .Y(uo_out[6]),
    .A2(_051_),
    .A1(_295_));
 sg13g2_nand2b_1 _360_ (.Y(_078_),
    .B(net6),
    .A_N(\tremolo_counter[7] ));
 sg13g2_and3_1 _361_ (.X(uo_out[7]),
    .A(net93),
    .B(tone_out),
    .C(_078_));
 sg13g2_nand2_1 _362_ (.Y(_079_),
    .A(net93),
    .B(net1));
 sg13g2_nor2b_1 _363_ (.A(\counter[18] ),
    .B_N(_000_),
    .Y(_080_));
 sg13g2_nand2_1 _364_ (.Y(_081_),
    .A(_001_),
    .B(_002_));
 sg13g2_nand3_1 _365_ (.B(_002_),
    .C(_080_),
    .A(_001_),
    .Y(_082_));
 sg13g2_and2_1 _366_ (.A(net94),
    .B(net96),
    .X(_083_));
 sg13g2_o21ai_1 _367_ (.B1(_047_),
    .Y(_084_),
    .A1(_045_),
    .A2(_061_));
 sg13g2_nand2_1 _368_ (.Y(_085_),
    .A(net100),
    .B(_046_));
 sg13g2_nand3_1 _369_ (.B(_084_),
    .C(_085_),
    .A(_070_),
    .Y(_086_));
 sg13g2_nor2b_2 _370_ (.A(net96),
    .B_N(net95),
    .Y(_087_));
 sg13g2_nor3_1 _371_ (.A(_045_),
    .B(_067_),
    .C(_075_),
    .Y(_088_));
 sg13g2_or3_1 _372_ (.A(_045_),
    .B(_067_),
    .C(_075_),
    .X(_089_));
 sg13g2_nor2_2 _373_ (.A(net94),
    .B(_289_),
    .Y(_090_));
 sg13g2_nand2b_1 _374_ (.Y(_091_),
    .B(net96),
    .A_N(net95));
 sg13g2_o21ai_1 _375_ (.B1(_076_),
    .Y(_092_),
    .A1(net103),
    .A2(_044_));
 sg13g2_nor2_1 _376_ (.A(net94),
    .B(net96),
    .Y(_093_));
 sg13g2_nand2_2 _377_ (.Y(_094_),
    .A(_050_),
    .B(_063_));
 sg13g2_mux4_1 _378_ (.S0(net3),
    .A0(_094_),
    .A1(_092_),
    .A2(_089_),
    .A3(_086_),
    .S1(net95),
    .X(_095_));
 sg13g2_a21o_1 _379_ (.A2(_051_),
    .A1(_295_),
    .B1(_047_),
    .X(_096_));
 sg13g2_a21o_1 _380_ (.A2(_085_),
    .A1(_069_),
    .B1(_096_),
    .X(_097_));
 sg13g2_mux4_1 _381_ (.S0(net3),
    .A0(_097_),
    .A1(_094_),
    .A2(_092_),
    .A3(_089_),
    .S1(net95),
    .X(_098_));
 sg13g2_and3_1 _382_ (.X(_099_),
    .A(net99),
    .B(_062_),
    .C(_066_));
 sg13g2_nand2_1 _383_ (.Y(_100_),
    .A(net105),
    .B(_053_));
 sg13g2_a22oi_1 _384_ (.Y(_101_),
    .B1(_059_),
    .B2(net92),
    .A2(_053_),
    .A1(net105));
 sg13g2_a21oi_1 _385_ (.A1(_295_),
    .A2(_061_),
    .Y(_102_),
    .B1(_052_));
 sg13g2_nand3b_1 _386_ (.B(_101_),
    .C(_102_),
    .Y(_103_),
    .A_N(_099_));
 sg13g2_a21o_1 _387_ (.A2(_066_),
    .A1(net99),
    .B1(_073_),
    .X(_104_));
 sg13g2_mux4_1 _388_ (.S0(net96),
    .A0(_103_),
    .A1(_104_),
    .A2(_097_),
    .A3(_094_),
    .S1(net95),
    .X(_105_));
 sg13g2_mux4_1 _389_ (.S0(net96),
    .A0(_104_),
    .A1(_097_),
    .A2(_094_),
    .A3(_092_),
    .S1(net95),
    .X(_106_));
 sg13g2_or3_1 _390_ (.A(_098_),
    .B(_105_),
    .C(_106_),
    .X(_107_));
 sg13g2_nor4_2 _391_ (.A(_095_),
    .B(_098_),
    .C(_105_),
    .Y(_108_),
    .D(_106_));
 sg13g2_nand2b_1 _392_ (.Y(_109_),
    .B(_090_),
    .A_N(_086_));
 sg13g2_a22oi_1 _393_ (.Y(_110_),
    .B1(_062_),
    .B2(net102),
    .A2(_046_),
    .A1(net99));
 sg13g2_a21oi_1 _394_ (.A1(net101),
    .A2(net105),
    .Y(_111_),
    .B1(net103));
 sg13g2_nor2_1 _395_ (.A(_295_),
    .B(_111_),
    .Y(_112_));
 sg13g2_a21oi_2 _396_ (.B1(_112_),
    .Y(_113_),
    .A2(_052_),
    .A1(_287_));
 sg13g2_a21o_1 _397_ (.A2(_052_),
    .A1(_287_),
    .B1(_112_),
    .X(_114_));
 sg13g2_nand2_1 _398_ (.Y(_115_),
    .A(_087_),
    .B(_113_));
 sg13g2_a22oi_1 _399_ (.Y(_116_),
    .B1(_110_),
    .B2(_083_),
    .A2(_093_),
    .A1(_088_));
 sg13g2_nand3_1 _400_ (.B(_115_),
    .C(_116_),
    .A(_109_),
    .Y(_117_));
 sg13g2_o21ai_1 _401_ (.B1(\counter[5] ),
    .Y(_118_),
    .A1(_108_),
    .A2(_117_));
 sg13g2_nand2_1 _402_ (.Y(_119_),
    .A(_089_),
    .B(_090_));
 sg13g2_nand2_1 _403_ (.Y(_120_),
    .A(_086_),
    .B(_087_));
 sg13g2_a22oi_1 _404_ (.Y(_121_),
    .B1(_114_),
    .B2(_083_),
    .A2(net87),
    .A1(_092_));
 sg13g2_nand3_1 _405_ (.B(_120_),
    .C(_121_),
    .A(_119_),
    .Y(_122_));
 sg13g2_xor2_1 _406_ (.B(_122_),
    .A(_108_),
    .X(_123_));
 sg13g2_o21ai_1 _407_ (.B1(_118_),
    .Y(_124_),
    .A1(_006_),
    .A2(_123_));
 sg13g2_nor3_1 _408_ (.A(\counter[5] ),
    .B(_108_),
    .C(_117_),
    .Y(_125_));
 sg13g2_o21ai_1 _409_ (.B1(net97),
    .Y(_126_),
    .A1(net92),
    .A2(_111_));
 sg13g2_and3_1 _410_ (.X(_127_),
    .A(_063_),
    .B(_100_),
    .C(_126_));
 sg13g2_a22oi_1 _411_ (.Y(_128_),
    .B1(_049_),
    .B2(net99),
    .A2(net104),
    .A1(net102));
 sg13g2_nor2_2 _412_ (.A(_099_),
    .B(_128_),
    .Y(_129_));
 sg13g2_mux4_1 _413_ (.S0(_289_),
    .A0(_110_),
    .A1(_113_),
    .A2(_127_),
    .A3(_129_),
    .S1(net4),
    .X(_130_));
 sg13g2_and2_1 _414_ (.A(_291_),
    .B(_130_),
    .X(_131_));
 sg13g2_nor2_1 _415_ (.A(_291_),
    .B(_130_),
    .Y(_132_));
 sg13g2_nor3_1 _416_ (.A(_087_),
    .B(_099_),
    .C(_128_),
    .Y(_133_));
 sg13g2_a21oi_1 _417_ (.A1(_087_),
    .A2(_110_),
    .Y(_134_),
    .B1(_133_));
 sg13g2_nor2_1 _418_ (.A(_091_),
    .B(_113_),
    .Y(_135_));
 sg13g2_a221oi_1 _419_ (.B2(net94),
    .C1(_135_),
    .B1(_134_),
    .A1(_086_),
    .Y(_136_),
    .A2(net87));
 sg13g2_xnor2_1 _420_ (.Y(_137_),
    .A(\counter[6] ),
    .B(_136_));
 sg13g2_nor4_1 _421_ (.A(_125_),
    .B(_131_),
    .C(_132_),
    .D(_137_),
    .Y(_138_));
 sg13g2_nand2_1 _422_ (.Y(_139_),
    .A(_006_),
    .B(_123_));
 sg13g2_nand3b_1 _423_ (.B(_138_),
    .C(_139_),
    .Y(_140_),
    .A_N(_124_));
 sg13g2_inv_1 _424_ (.Y(_141_),
    .A(_140_));
 sg13g2_xor2_1 _425_ (.B(_106_),
    .A(_105_),
    .X(_142_));
 sg13g2_nand2_1 _426_ (.Y(_143_),
    .A(\counter[1] ),
    .B(_142_));
 sg13g2_nor2_1 _427_ (.A(\counter[0] ),
    .B(_105_),
    .Y(_144_));
 sg13g2_xnor2_1 _428_ (.Y(_145_),
    .A(\counter[1] ),
    .B(_142_));
 sg13g2_o21ai_1 _429_ (.B1(_143_),
    .Y(_146_),
    .A1(_144_),
    .A2(_145_));
 sg13g2_xnor2_1 _430_ (.Y(_147_),
    .A(_095_),
    .B(_107_));
 sg13g2_nand2_1 _431_ (.Y(_148_),
    .A(_292_),
    .B(_147_));
 sg13g2_o21ai_1 _432_ (.B1(_098_),
    .Y(_149_),
    .A1(_105_),
    .A2(_106_));
 sg13g2_nand3_1 _433_ (.B(_107_),
    .C(_149_),
    .A(_007_),
    .Y(_150_));
 sg13g2_a21o_1 _434_ (.A2(_149_),
    .A1(_107_),
    .B1(_007_),
    .X(_151_));
 sg13g2_a22oi_1 _435_ (.Y(_152_),
    .B1(_150_),
    .B2(_151_),
    .A2(_147_),
    .A1(_292_));
 sg13g2_nor2_1 _436_ (.A(_292_),
    .B(_147_),
    .Y(_153_));
 sg13g2_and3_1 _437_ (.X(_154_),
    .A(\counter[2] ),
    .B(_107_),
    .C(_149_));
 sg13g2_a221oi_1 _438_ (.B2(_148_),
    .C1(_153_),
    .B1(_154_),
    .A1(_146_),
    .Y(_155_),
    .A2(_152_));
 sg13g2_a22oi_1 _439_ (.Y(_156_),
    .B1(_136_),
    .B2(_293_),
    .A2(_130_),
    .A1(_291_));
 sg13g2_nor2_1 _440_ (.A(_132_),
    .B(_156_),
    .Y(_157_));
 sg13g2_a21oi_1 _441_ (.A1(_124_),
    .A2(_138_),
    .Y(_158_),
    .B1(_157_));
 sg13g2_o21ai_1 _442_ (.B1(_158_),
    .Y(_159_),
    .A1(_140_),
    .A2(_155_));
 sg13g2_nor2_2 _443_ (.A(net92),
    .B(_054_),
    .Y(_160_));
 sg13g2_a21oi_1 _444_ (.A1(_295_),
    .A2(net92),
    .Y(_161_),
    .B1(_160_));
 sg13g2_a21o_1 _445_ (.A2(net92),
    .A1(_295_),
    .B1(_160_),
    .X(_162_));
 sg13g2_o21ai_1 _446_ (.B1(_091_),
    .Y(_163_),
    .A1(_134_),
    .A2(_161_));
 sg13g2_nand2b_1 _447_ (.Y(_164_),
    .B(_162_),
    .A_N(net94));
 sg13g2_nor2_1 _448_ (.A(_047_),
    .B(_049_),
    .Y(_165_));
 sg13g2_nor2_1 _449_ (.A(_059_),
    .B(_165_),
    .Y(_166_));
 sg13g2_o21ai_1 _450_ (.B1(_060_),
    .Y(_167_),
    .A1(_047_),
    .A2(_049_));
 sg13g2_a22oi_1 _451_ (.Y(_168_),
    .B1(_167_),
    .B2(net87),
    .A2(_164_),
    .A1(_163_));
 sg13g2_xnor2_1 _452_ (.Y(_169_),
    .A(\counter[12] ),
    .B(_168_));
 sg13g2_a22oi_1 _453_ (.Y(_170_),
    .B1(_161_),
    .B2(net87),
    .A2(_160_),
    .A1(_090_));
 sg13g2_and2_1 _454_ (.A(\counter[13] ),
    .B(_170_),
    .X(_171_));
 sg13g2_nor2_1 _455_ (.A(\counter[13] ),
    .B(_170_),
    .Y(_172_));
 sg13g2_nand2_1 _456_ (.Y(_173_),
    .A(net87),
    .B(_160_));
 sg13g2_xor2_1 _457_ (.B(_173_),
    .A(\counter[14] ),
    .X(_174_));
 sg13g2_nand2_1 _458_ (.Y(_175_),
    .A(_003_),
    .B(_174_));
 sg13g2_nor4_2 _459_ (.A(_169_),
    .B(_171_),
    .C(_172_),
    .Y(_176_),
    .D(_175_));
 sg13g2_a221oi_1 _460_ (.B2(_053_),
    .C1(_052_),
    .B1(net92),
    .A1(_288_),
    .Y(_177_),
    .A2(_047_));
 sg13g2_nor2b_2 _461_ (.A(_067_),
    .B_N(_177_),
    .Y(_178_));
 sg13g2_nand2b_1 _462_ (.Y(_179_),
    .B(net97),
    .A_N(_087_));
 sg13g2_o21ai_1 _463_ (.B1(net94),
    .Y(_180_),
    .A1(_165_),
    .A2(_179_));
 sg13g2_a21oi_1 _464_ (.A1(_167_),
    .A2(_179_),
    .Y(_181_),
    .B1(_180_));
 sg13g2_a221oi_1 _465_ (.B2(_090_),
    .C1(_181_),
    .B1(_178_),
    .A1(net87),
    .Y(_182_),
    .A2(_127_));
 sg13g2_xor2_1 _466_ (.B(_182_),
    .A(\counter[10] ),
    .X(_183_));
 sg13g2_mux4_1 _467_ (.S0(_289_),
    .A0(_127_),
    .A1(_129_),
    .A2(_166_),
    .A3(_178_),
    .S1(net94),
    .X(_184_));
 sg13g2_nor2_1 _468_ (.A(\counter[9] ),
    .B(_184_),
    .Y(_185_));
 sg13g2_nand2_1 _469_ (.Y(_186_),
    .A(net87),
    .B(_178_));
 sg13g2_o21ai_1 _470_ (.B1(_083_),
    .Y(_187_),
    .A1(net92),
    .A2(_054_));
 sg13g2_o21ai_1 _471_ (.B1(_187_),
    .Y(_188_),
    .A1(_091_),
    .A2(_167_));
 sg13g2_a21oi_1 _472_ (.A1(_087_),
    .A2(_162_),
    .Y(_189_),
    .B1(_188_));
 sg13g2_nand3_1 _473_ (.B(_186_),
    .C(_189_),
    .A(_004_),
    .Y(_190_));
 sg13g2_a21o_1 _474_ (.A2(_189_),
    .A1(_186_),
    .B1(_004_),
    .X(_191_));
 sg13g2_nand2_1 _475_ (.Y(_192_),
    .A(_190_),
    .B(_191_));
 sg13g2_nor3_1 _476_ (.A(_183_),
    .B(_185_),
    .C(_192_),
    .Y(_193_));
 sg13g2_nand2_1 _477_ (.Y(_194_),
    .A(\counter[9] ),
    .B(_184_));
 sg13g2_a21oi_1 _478_ (.A1(net95),
    .A2(_127_),
    .Y(_195_),
    .B1(net96));
 sg13g2_nor2_1 _479_ (.A(net94),
    .B(_129_),
    .Y(_196_));
 sg13g2_nor2b_1 _480_ (.A(_178_),
    .B_N(_083_),
    .Y(_197_));
 sg13g2_nor3_1 _481_ (.A(_195_),
    .B(_196_),
    .C(_197_),
    .Y(_198_));
 sg13g2_a21oi_1 _482_ (.A1(net87),
    .A2(_110_),
    .Y(_199_),
    .B1(_198_));
 sg13g2_xnor2_1 _483_ (.Y(_200_),
    .A(\counter[8] ),
    .B(_199_));
 sg13g2_and3_1 _484_ (.X(_201_),
    .A(_193_),
    .B(_194_),
    .C(_200_));
 sg13g2_and2_1 _485_ (.A(_176_),
    .B(_201_),
    .X(_202_));
 sg13g2_nor2_1 _486_ (.A(_010_),
    .B(_172_),
    .Y(_203_));
 sg13g2_a21oi_1 _487_ (.A1(_168_),
    .A2(_203_),
    .Y(_204_),
    .B1(_171_));
 sg13g2_nor2b_1 _488_ (.A(_204_),
    .B_N(_174_),
    .Y(_205_));
 sg13g2_nand2b_1 _489_ (.Y(_206_),
    .B(_173_),
    .A_N(_009_));
 sg13g2_nand3b_1 _490_ (.B(_206_),
    .C(_003_),
    .Y(_207_),
    .A_N(_205_));
 sg13g2_o21ai_1 _491_ (.B1(_194_),
    .Y(_208_),
    .A1(_012_),
    .A2(_199_));
 sg13g2_o21ai_1 _492_ (.B1(_191_),
    .Y(_209_),
    .A1(_011_),
    .A2(_182_));
 sg13g2_a22oi_1 _493_ (.Y(_210_),
    .B1(_209_),
    .B2(_190_),
    .A2(_208_),
    .A1(_193_));
 sg13g2_inv_1 _494_ (.Y(_211_),
    .A(_210_));
 sg13g2_a221oi_1 _495_ (.B2(_176_),
    .C1(_207_),
    .B1(_211_),
    .A1(_159_),
    .Y(_212_),
    .A2(_202_));
 sg13g2_a21oi_1 _496_ (.A1(_080_),
    .A2(_081_),
    .Y(_213_),
    .B1(net89));
 sg13g2_nand3_1 _497_ (.B(_008_),
    .C(_213_),
    .A(_000_),
    .Y(_214_));
 sg13g2_and2_1 _498_ (.A(\counter[0] ),
    .B(_105_),
    .X(_215_));
 sg13g2_nor2_1 _499_ (.A(_082_),
    .B(_153_),
    .Y(_216_));
 sg13g2_nor3_1 _500_ (.A(_144_),
    .B(_145_),
    .C(_215_),
    .Y(_217_));
 sg13g2_and2_1 _501_ (.A(_152_),
    .B(_217_),
    .X(_218_));
 sg13g2_and4_1 _502_ (.A(_176_),
    .B(_201_),
    .C(_216_),
    .D(_218_),
    .X(_219_));
 sg13g2_a21oi_1 _503_ (.A1(_141_),
    .A2(_219_),
    .Y(_220_),
    .B1(_214_));
 sg13g2_o21ai_1 _504_ (.B1(_220_),
    .Y(_221_),
    .A1(_082_),
    .A2(_212_));
 sg13g2_nand2_1 _505_ (.Y(_222_),
    .A(net71),
    .B(net89));
 sg13g2_o21ai_1 _506_ (.B1(_222_),
    .Y(_015_),
    .A1(net71),
    .A2(net86));
 sg13g2_nand2_1 _507_ (.Y(_223_),
    .A(net73),
    .B(net90));
 sg13g2_nand2_1 _508_ (.Y(_224_),
    .A(\counter[1] ),
    .B(\counter[0] ));
 sg13g2_xnor2_1 _509_ (.Y(_225_),
    .A(net73),
    .B(net71));
 sg13g2_o21ai_1 _510_ (.B1(_223_),
    .Y(_016_),
    .A1(net85),
    .A2(_225_));
 sg13g2_nand2_1 _511_ (.Y(_226_),
    .A(net59),
    .B(net90));
 sg13g2_xnor2_1 _512_ (.Y(_227_),
    .A(_007_),
    .B(_224_));
 sg13g2_o21ai_1 _513_ (.B1(_226_),
    .Y(_017_),
    .A1(net85),
    .A2(_227_));
 sg13g2_nand2_1 _514_ (.Y(_228_),
    .A(net43),
    .B(net89));
 sg13g2_nand3_1 _515_ (.B(\counter[1] ),
    .C(\counter[0] ),
    .A(\counter[2] ),
    .Y(_229_));
 sg13g2_nor2_1 _516_ (.A(_292_),
    .B(_229_),
    .Y(_230_));
 sg13g2_xnor2_1 _517_ (.Y(_231_),
    .A(_292_),
    .B(_229_));
 sg13g2_o21ai_1 _518_ (.B1(_228_),
    .Y(_018_),
    .A1(net85),
    .A2(_231_));
 sg13g2_nand2_1 _519_ (.Y(_232_),
    .A(net51),
    .B(net90));
 sg13g2_xor2_1 _520_ (.B(_230_),
    .A(_006_),
    .X(_233_));
 sg13g2_o21ai_1 _521_ (.B1(_232_),
    .Y(_019_),
    .A1(net86),
    .A2(_233_));
 sg13g2_nand2_1 _522_ (.Y(_234_),
    .A(net69),
    .B(net90));
 sg13g2_nand3_1 _523_ (.B(net51),
    .C(_230_),
    .A(\counter[5] ),
    .Y(_235_));
 sg13g2_a21o_1 _524_ (.A2(_230_),
    .A1(net51),
    .B1(net69),
    .X(_236_));
 sg13g2_nand2_1 _525_ (.Y(_237_),
    .A(_235_),
    .B(_236_));
 sg13g2_o21ai_1 _526_ (.B1(_234_),
    .Y(_020_),
    .A1(net85),
    .A2(_237_));
 sg13g2_nand2_1 _527_ (.Y(_238_),
    .A(net61),
    .B(net91));
 sg13g2_nor2_1 _528_ (.A(_013_),
    .B(_235_),
    .Y(_239_));
 sg13g2_xnor2_1 _529_ (.Y(_240_),
    .A(_013_),
    .B(_235_));
 sg13g2_o21ai_1 _530_ (.B1(_238_),
    .Y(_021_),
    .A1(net86),
    .A2(_240_));
 sg13g2_nand2_1 _531_ (.Y(_241_),
    .A(net29),
    .B(net89));
 sg13g2_xnor2_1 _532_ (.Y(_242_),
    .A(_291_),
    .B(_239_));
 sg13g2_o21ai_1 _533_ (.B1(_241_),
    .Y(_022_),
    .A1(net85),
    .A2(_242_));
 sg13g2_nand2_1 _534_ (.Y(_243_),
    .A(net57),
    .B(net88));
 sg13g2_nand2_1 _535_ (.Y(_244_),
    .A(net29),
    .B(\counter[6] ));
 sg13g2_or2_1 _536_ (.X(_245_),
    .B(_244_),
    .A(_235_));
 sg13g2_xnor2_1 _537_ (.Y(_246_),
    .A(_012_),
    .B(_245_));
 sg13g2_o21ai_1 _538_ (.B1(_243_),
    .Y(_023_),
    .A1(net84),
    .A2(_246_));
 sg13g2_nand2_1 _539_ (.Y(_247_),
    .A(net70),
    .B(net88));
 sg13g2_nor2_2 _540_ (.A(_290_),
    .B(_245_),
    .Y(_248_));
 sg13g2_nand2_1 _541_ (.Y(_249_),
    .A(\counter[9] ),
    .B(_248_));
 sg13g2_xnor2_1 _542_ (.Y(_250_),
    .A(net70),
    .B(_248_));
 sg13g2_o21ai_1 _543_ (.B1(_247_),
    .Y(_024_),
    .A1(net84),
    .A2(_250_));
 sg13g2_nand2_1 _544_ (.Y(_251_),
    .A(net55),
    .B(net88));
 sg13g2_nor2_1 _545_ (.A(_011_),
    .B(_249_),
    .Y(_252_));
 sg13g2_xnor2_1 _546_ (.Y(_253_),
    .A(_011_),
    .B(_249_));
 sg13g2_o21ai_1 _547_ (.B1(_251_),
    .Y(_025_),
    .A1(net84),
    .A2(_253_));
 sg13g2_nand2_1 _548_ (.Y(_254_),
    .A(net37),
    .B(net88));
 sg13g2_xor2_1 _549_ (.B(_252_),
    .A(_004_),
    .X(_255_));
 sg13g2_o21ai_1 _550_ (.B1(_254_),
    .Y(_026_),
    .A1(net84),
    .A2(_255_));
 sg13g2_nand2_1 _551_ (.Y(_256_),
    .A(net65),
    .B(net88));
 sg13g2_and4_1 _552_ (.A(net37),
    .B(net55),
    .C(\counter[9] ),
    .D(_248_),
    .X(_257_));
 sg13g2_xor2_1 _553_ (.B(_257_),
    .A(_010_),
    .X(_258_));
 sg13g2_o21ai_1 _554_ (.B1(_256_),
    .Y(_027_),
    .A1(net84),
    .A2(_258_));
 sg13g2_nand2_1 _555_ (.Y(_259_),
    .A(net67),
    .B(net88));
 sg13g2_a21oi_1 _556_ (.A1(net65),
    .A2(_257_),
    .Y(_260_),
    .B1(net67));
 sg13g2_nand3_1 _557_ (.B(\counter[12] ),
    .C(_257_),
    .A(\counter[13] ),
    .Y(_261_));
 sg13g2_inv_1 _558_ (.Y(_262_),
    .A(_261_));
 sg13g2_nand2b_1 _559_ (.Y(_263_),
    .B(_261_),
    .A_N(_260_));
 sg13g2_o21ai_1 _560_ (.B1(_259_),
    .Y(_028_),
    .A1(net84),
    .A2(_263_));
 sg13g2_nand2_1 _561_ (.Y(_264_),
    .A(net63),
    .B(net88));
 sg13g2_nor2_1 _562_ (.A(_009_),
    .B(_261_),
    .Y(_265_));
 sg13g2_xnor2_1 _563_ (.Y(_266_),
    .A(_009_),
    .B(_261_));
 sg13g2_o21ai_1 _564_ (.B1(_264_),
    .Y(_029_),
    .A1(net84),
    .A2(_266_));
 sg13g2_nand2_1 _565_ (.Y(_267_),
    .A(net47),
    .B(net88));
 sg13g2_xor2_1 _566_ (.B(_265_),
    .A(_003_),
    .X(_268_));
 sg13g2_o21ai_1 _567_ (.B1(_267_),
    .Y(_030_),
    .A1(net86),
    .A2(_268_));
 sg13g2_nand2_1 _568_ (.Y(_269_),
    .A(net33),
    .B(net89));
 sg13g2_nand3_1 _569_ (.B(\counter[14] ),
    .C(_262_),
    .A(\counter[15] ),
    .Y(_270_));
 sg13g2_nor2_1 _570_ (.A(_002_),
    .B(_270_),
    .Y(_271_));
 sg13g2_xnor2_1 _571_ (.Y(_272_),
    .A(_002_),
    .B(_270_));
 sg13g2_o21ai_1 _572_ (.B1(_269_),
    .Y(_031_),
    .A1(net85),
    .A2(_272_));
 sg13g2_nand2_1 _573_ (.Y(_273_),
    .A(net35),
    .B(net89));
 sg13g2_xor2_1 _574_ (.B(_271_),
    .A(_001_),
    .X(_274_));
 sg13g2_o21ai_1 _575_ (.B1(_273_),
    .Y(_032_),
    .A1(net85),
    .A2(_274_));
 sg13g2_nand2_1 _576_ (.Y(_275_),
    .A(net45),
    .B(net89));
 sg13g2_nand2_1 _577_ (.Y(_276_),
    .A(net35),
    .B(net33));
 sg13g2_nor2_1 _578_ (.A(_270_),
    .B(_276_),
    .Y(_277_));
 sg13g2_xor2_1 _579_ (.B(_277_),
    .A(_008_),
    .X(_278_));
 sg13g2_o21ai_1 _580_ (.B1(_275_),
    .Y(_033_),
    .A1(net85),
    .A2(_278_));
 sg13g2_and2_1 _581_ (.A(net25),
    .B(net89),
    .X(_034_));
 sg13g2_nor2_1 _582_ (.A(net68),
    .B(net91),
    .Y(_279_));
 sg13g2_mux2_1 _583_ (.A0(net68),
    .A1(_279_),
    .S(net84),
    .X(_035_));
 sg13g2_mux2_1 _584_ (.A0(net23),
    .A1(\tremolo_counter[0] ),
    .S(net90),
    .X(_036_));
 sg13g2_nand3_1 _585_ (.B(net1),
    .C(\tremolo_counter[0] ),
    .A(net5),
    .Y(_280_));
 sg13g2_nand4_1 _586_ (.B(net1),
    .C(\tremolo_counter[0] ),
    .A(net5),
    .Y(_281_),
    .D(net39));
 sg13g2_xnor2_1 _587_ (.Y(_037_),
    .A(net39),
    .B(_280_));
 sg13g2_nor2_1 _588_ (.A(_294_),
    .B(_281_),
    .Y(_282_));
 sg13g2_xnor2_1 _589_ (.Y(_038_),
    .A(net41),
    .B(_281_));
 sg13g2_xor2_1 _590_ (.B(_282_),
    .A(net53),
    .X(_039_));
 sg13g2_and3_1 _591_ (.X(_283_),
    .A(\tremolo_counter[3] ),
    .B(net26),
    .C(_282_));
 sg13g2_a21oi_1 _592_ (.A1(\tremolo_counter[3] ),
    .A2(_282_),
    .Y(_284_),
    .B1(net26));
 sg13g2_nor2_1 _593_ (.A(_283_),
    .B(net27),
    .Y(_040_));
 sg13g2_xor2_1 _594_ (.B(_283_),
    .A(net49),
    .X(_041_));
 sg13g2_nand3_1 _595_ (.B(net74),
    .C(_283_),
    .A(net49),
    .Y(_285_));
 sg13g2_a21o_1 _596_ (.A2(_283_),
    .A1(net49),
    .B1(net74),
    .X(_286_));
 sg13g2_and2_1 _597_ (.A(_285_),
    .B(_286_),
    .X(_042_));
 sg13g2_xnor2_1 _598_ (.Y(_043_),
    .A(net31),
    .B(_285_));
 sg13g2_dfrbp_1 _599_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net110),
    .D(net72),
    .Q_N(_309_),
    .Q(\counter[0] ));
 sg13g2_dfrbp_1 _600_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net111),
    .D(_016_),
    .Q_N(_308_),
    .Q(\counter[1] ));
 sg13g2_dfrbp_1 _601_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net111),
    .D(net60),
    .Q_N(_007_),
    .Q(\counter[2] ));
 sg13g2_dfrbp_1 _602_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net110),
    .D(net44),
    .Q_N(_307_),
    .Q(\counter[3] ));
 sg13g2_dfrbp_1 _603_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net110),
    .D(net52),
    .Q_N(_006_),
    .Q(\counter[4] ));
 sg13g2_dfrbp_1 _604_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net110),
    .D(_020_),
    .Q_N(_306_),
    .Q(\counter[5] ));
 sg13g2_dfrbp_1 _605_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net107),
    .D(net62),
    .Q_N(_013_),
    .Q(\counter[6] ));
 sg13g2_dfrbp_1 _606_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net107),
    .D(net30),
    .Q_N(_005_),
    .Q(\counter[7] ));
 sg13g2_dfrbp_1 _607_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net107),
    .D(net58),
    .Q_N(_012_),
    .Q(\counter[8] ));
 sg13g2_dfrbp_1 _608_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net107),
    .D(_024_),
    .Q_N(_305_),
    .Q(\counter[9] ));
 sg13g2_dfrbp_1 _609_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net107),
    .D(net56),
    .Q_N(_011_),
    .Q(\counter[10] ));
 sg13g2_dfrbp_1 _610_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net108),
    .D(net38),
    .Q_N(_004_),
    .Q(\counter[11] ));
 sg13g2_dfrbp_1 _611_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net107),
    .D(net66),
    .Q_N(_010_),
    .Q(\counter[12] ));
 sg13g2_dfrbp_1 _612_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net107),
    .D(_028_),
    .Q_N(_304_),
    .Q(\counter[13] ));
 sg13g2_dfrbp_1 _613_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net108),
    .D(net64),
    .Q_N(_009_),
    .Q(\counter[14] ));
 sg13g2_dfrbp_1 _614_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net107),
    .D(net48),
    .Q_N(_003_),
    .Q(\counter[15] ));
 sg13g2_dfrbp_1 _615_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net110),
    .D(net34),
    .Q_N(_002_),
    .Q(\counter[16] ));
 sg13g2_dfrbp_1 _616_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net110),
    .D(net36),
    .Q_N(_001_),
    .Q(\counter[17] ));
 sg13g2_dfrbp_1 _617_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net110),
    .D(net46),
    .Q_N(_008_),
    .Q(\counter[18] ));
 sg13g2_dfrbp_1 _618_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net110),
    .D(_034_),
    .Q_N(_000_),
    .Q(\counter[19] ));
 sg13g2_dfrbp_1 _619_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net108),
    .D(_035_),
    .Q_N(_303_),
    .Q(tone_out));
 sg13g2_dfrbp_1 _620_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net109),
    .D(net24),
    .Q_N(_014_),
    .Q(\tremolo_counter[0] ));
 sg13g2_dfrbp_1 _621_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net109),
    .D(net40),
    .Q_N(_302_),
    .Q(\tremolo_counter[1] ));
 sg13g2_dfrbp_1 _622_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net109),
    .D(net42),
    .Q_N(_301_),
    .Q(\tremolo_counter[2] ));
 sg13g2_dfrbp_1 _623_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net109),
    .D(net54),
    .Q_N(_300_),
    .Q(\tremolo_counter[3] ));
 sg13g2_dfrbp_1 _624_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net109),
    .D(net28),
    .Q_N(_299_),
    .Q(\tremolo_counter[4] ));
 sg13g2_dfrbp_1 _625_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net109),
    .D(net50),
    .Q_N(_298_),
    .Q(\tremolo_counter[5] ));
 sg13g2_dfrbp_1 _626_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net109),
    .D(_042_),
    .Q_N(_297_),
    .Q(\tremolo_counter[6] ));
 sg13g2_dfrbp_1 _627_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net109),
    .D(net32),
    .Q_N(_296_),
    .Q(\tremolo_counter[7] ));
 sg13g2_tielo tt_um_kentrane_tinyspectrum_8 (.L_LO(net8));
 sg13g2_tielo tt_um_kentrane_tinyspectrum_9 (.L_LO(net9));
 sg13g2_tielo tt_um_kentrane_tinyspectrum_10 (.L_LO(net10));
 sg13g2_tielo tt_um_kentrane_tinyspectrum_11 (.L_LO(net11));
 sg13g2_tielo tt_um_kentrane_tinyspectrum_12 (.L_LO(net12));
 sg13g2_tielo tt_um_kentrane_tinyspectrum_13 (.L_LO(net13));
 sg13g2_tielo tt_um_kentrane_tinyspectrum_14 (.L_LO(net14));
 sg13g2_tielo tt_um_kentrane_tinyspectrum_15 (.L_LO(net15));
 sg13g2_tielo tt_um_kentrane_tinyspectrum_16 (.L_LO(net16));
 sg13g2_tielo tt_um_kentrane_tinyspectrum_17 (.L_LO(net17));
 sg13g2_tielo tt_um_kentrane_tinyspectrum_18 (.L_LO(net18));
 sg13g2_tielo tt_um_kentrane_tinyspectrum_19 (.L_LO(net19));
 sg13g2_tielo tt_um_kentrane_tinyspectrum_20 (.L_LO(net20));
 sg13g2_tielo tt_um_kentrane_tinyspectrum_21 (.L_LO(net21));
 sg13g2_tielo tt_um_kentrane_tinyspectrum_22 (.L_LO(net22));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_4 fanout84 (.X(net84),
    .A(net86));
 sg13g2_buf_2 fanout85 (.A(net86),
    .X(net85));
 sg13g2_buf_2 fanout86 (.A(_221_),
    .X(net86));
 sg13g2_buf_2 fanout87 (.A(_093_),
    .X(net87));
 sg13g2_buf_2 fanout88 (.A(net91),
    .X(net88));
 sg13g2_buf_2 fanout89 (.A(net90),
    .X(net89));
 sg13g2_buf_2 fanout90 (.A(net91),
    .X(net90));
 sg13g2_buf_2 fanout91 (.A(_079_),
    .X(net91));
 sg13g2_buf_2 fanout92 (.A(_048_),
    .X(net92));
 sg13g2_buf_2 fanout93 (.A(net5),
    .X(net93));
 sg13g2_buf_2 fanout94 (.A(net95),
    .X(net94));
 sg13g2_buf_2 fanout95 (.A(net4),
    .X(net95));
 sg13g2_buf_4 fanout96 (.X(net96),
    .A(net3));
 sg13g2_buf_2 fanout97 (.A(net99),
    .X(net97));
 sg13g2_buf_1 fanout98 (.A(net99),
    .X(net98));
 sg13g2_buf_2 fanout99 (.A(net2),
    .X(net99));
 sg13g2_buf_2 fanout100 (.A(net101),
    .X(net100));
 sg13g2_buf_1 fanout101 (.A(net102),
    .X(net101));
 sg13g2_buf_2 fanout102 (.A(ui_in[2]),
    .X(net102));
 sg13g2_buf_2 fanout103 (.A(ui_in[1]),
    .X(net103));
 sg13g2_buf_2 fanout104 (.A(ui_in[1]),
    .X(net104));
 sg13g2_buf_2 fanout105 (.A(ui_in[0]),
    .X(net105));
 sg13g2_buf_2 fanout106 (.A(ui_in[0]),
    .X(net106));
 sg13g2_buf_4 fanout107 (.X(net107),
    .A(net108));
 sg13g2_buf_4 fanout108 (.X(net108),
    .A(net111));
 sg13g2_buf_4 fanout109 (.X(net109),
    .A(net111));
 sg13g2_buf_4 fanout110 (.X(net110),
    .A(net111));
 sg13g2_buf_2 fanout111 (.A(rst_n),
    .X(net111));
 sg13g2_buf_1 input1 (.A(ena),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[3]),
    .X(net2));
 sg13g2_buf_2 input3 (.A(ui_in[4]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[5]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[6]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[7]),
    .X(net6));
 sg13g2_tielo tt_um_kentrane_tinyspectrum_7 (.L_LO(net7));
 sg13g2_buf_2 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sg13g2_buf_2 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sg13g2_buf_2 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sg13g2_buf_2 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sg13g2_buf_2 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sg13g2_buf_2 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sg13g2_buf_2 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sg13g2_buf_2 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_3_3__leaf_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_3_5__leaf_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_3_7__leaf_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(_014_),
    .X(net23));
 sg13g2_dlygate4sd3_1 hold2 (.A(_036_),
    .X(net24));
 sg13g2_dlygate4sd3_1 hold3 (.A(\counter[19] ),
    .X(net25));
 sg13g2_dlygate4sd3_1 hold4 (.A(\tremolo_counter[4] ),
    .X(net26));
 sg13g2_dlygate4sd3_1 hold5 (.A(_284_),
    .X(net27));
 sg13g2_dlygate4sd3_1 hold6 (.A(_040_),
    .X(net28));
 sg13g2_dlygate4sd3_1 hold7 (.A(\counter[7] ),
    .X(net29));
 sg13g2_dlygate4sd3_1 hold8 (.A(_022_),
    .X(net30));
 sg13g2_dlygate4sd3_1 hold9 (.A(\tremolo_counter[7] ),
    .X(net31));
 sg13g2_dlygate4sd3_1 hold10 (.A(_043_),
    .X(net32));
 sg13g2_dlygate4sd3_1 hold11 (.A(\counter[16] ),
    .X(net33));
 sg13g2_dlygate4sd3_1 hold12 (.A(_031_),
    .X(net34));
 sg13g2_dlygate4sd3_1 hold13 (.A(\counter[17] ),
    .X(net35));
 sg13g2_dlygate4sd3_1 hold14 (.A(_032_),
    .X(net36));
 sg13g2_dlygate4sd3_1 hold15 (.A(\counter[11] ),
    .X(net37));
 sg13g2_dlygate4sd3_1 hold16 (.A(_026_),
    .X(net38));
 sg13g2_dlygate4sd3_1 hold17 (.A(\tremolo_counter[1] ),
    .X(net39));
 sg13g2_dlygate4sd3_1 hold18 (.A(_037_),
    .X(net40));
 sg13g2_dlygate4sd3_1 hold19 (.A(\tremolo_counter[2] ),
    .X(net41));
 sg13g2_dlygate4sd3_1 hold20 (.A(_038_),
    .X(net42));
 sg13g2_dlygate4sd3_1 hold21 (.A(\counter[3] ),
    .X(net43));
 sg13g2_dlygate4sd3_1 hold22 (.A(_018_),
    .X(net44));
 sg13g2_dlygate4sd3_1 hold23 (.A(\counter[18] ),
    .X(net45));
 sg13g2_dlygate4sd3_1 hold24 (.A(_033_),
    .X(net46));
 sg13g2_dlygate4sd3_1 hold25 (.A(\counter[15] ),
    .X(net47));
 sg13g2_dlygate4sd3_1 hold26 (.A(_030_),
    .X(net48));
 sg13g2_dlygate4sd3_1 hold27 (.A(\tremolo_counter[5] ),
    .X(net49));
 sg13g2_dlygate4sd3_1 hold28 (.A(_041_),
    .X(net50));
 sg13g2_dlygate4sd3_1 hold29 (.A(\counter[4] ),
    .X(net51));
 sg13g2_dlygate4sd3_1 hold30 (.A(_019_),
    .X(net52));
 sg13g2_dlygate4sd3_1 hold31 (.A(\tremolo_counter[3] ),
    .X(net53));
 sg13g2_dlygate4sd3_1 hold32 (.A(_039_),
    .X(net54));
 sg13g2_dlygate4sd3_1 hold33 (.A(\counter[10] ),
    .X(net55));
 sg13g2_dlygate4sd3_1 hold34 (.A(_025_),
    .X(net56));
 sg13g2_dlygate4sd3_1 hold35 (.A(\counter[8] ),
    .X(net57));
 sg13g2_dlygate4sd3_1 hold36 (.A(_023_),
    .X(net58));
 sg13g2_dlygate4sd3_1 hold37 (.A(\counter[2] ),
    .X(net59));
 sg13g2_dlygate4sd3_1 hold38 (.A(_017_),
    .X(net60));
 sg13g2_dlygate4sd3_1 hold39 (.A(\counter[6] ),
    .X(net61));
 sg13g2_dlygate4sd3_1 hold40 (.A(_021_),
    .X(net62));
 sg13g2_dlygate4sd3_1 hold41 (.A(\counter[14] ),
    .X(net63));
 sg13g2_dlygate4sd3_1 hold42 (.A(_029_),
    .X(net64));
 sg13g2_dlygate4sd3_1 hold43 (.A(\counter[12] ),
    .X(net65));
 sg13g2_dlygate4sd3_1 hold44 (.A(_027_),
    .X(net66));
 sg13g2_dlygate4sd3_1 hold45 (.A(\counter[13] ),
    .X(net67));
 sg13g2_dlygate4sd3_1 hold46 (.A(tone_out),
    .X(net68));
 sg13g2_dlygate4sd3_1 hold47 (.A(\counter[5] ),
    .X(net69));
 sg13g2_dlygate4sd3_1 hold48 (.A(\counter[9] ),
    .X(net70));
 sg13g2_dlygate4sd3_1 hold49 (.A(\counter[0] ),
    .X(net71));
 sg13g2_dlygate4sd3_1 hold50 (.A(_015_),
    .X(net72));
 sg13g2_dlygate4sd3_1 hold51 (.A(\counter[1] ),
    .X(net73));
 sg13g2_dlygate4sd3_1 hold52 (.A(\tremolo_counter[6] ),
    .X(net74));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_fill_2 FILLER_14_406 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_252 ();
 sg13g2_decap_8 FILLER_15_259 ();
 sg13g2_decap_8 FILLER_15_266 ();
 sg13g2_decap_8 FILLER_15_273 ();
 sg13g2_decap_8 FILLER_15_280 ();
 sg13g2_decap_8 FILLER_15_287 ();
 sg13g2_decap_8 FILLER_15_294 ();
 sg13g2_decap_8 FILLER_15_301 ();
 sg13g2_decap_8 FILLER_15_308 ();
 sg13g2_decap_8 FILLER_15_315 ();
 sg13g2_decap_8 FILLER_15_322 ();
 sg13g2_decap_8 FILLER_15_329 ();
 sg13g2_decap_8 FILLER_15_336 ();
 sg13g2_decap_8 FILLER_15_343 ();
 sg13g2_decap_8 FILLER_15_350 ();
 sg13g2_decap_8 FILLER_15_357 ();
 sg13g2_decap_8 FILLER_15_364 ();
 sg13g2_decap_8 FILLER_15_371 ();
 sg13g2_decap_8 FILLER_15_378 ();
 sg13g2_decap_8 FILLER_15_385 ();
 sg13g2_decap_8 FILLER_15_392 ();
 sg13g2_decap_8 FILLER_15_399 ();
 sg13g2_fill_2 FILLER_15_406 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_decap_8 FILLER_16_217 ();
 sg13g2_decap_8 FILLER_16_224 ();
 sg13g2_decap_8 FILLER_16_231 ();
 sg13g2_decap_8 FILLER_16_238 ();
 sg13g2_decap_8 FILLER_16_245 ();
 sg13g2_decap_8 FILLER_16_252 ();
 sg13g2_decap_8 FILLER_16_259 ();
 sg13g2_decap_8 FILLER_16_266 ();
 sg13g2_decap_8 FILLER_16_273 ();
 sg13g2_decap_8 FILLER_16_280 ();
 sg13g2_decap_8 FILLER_16_287 ();
 sg13g2_decap_8 FILLER_16_294 ();
 sg13g2_decap_8 FILLER_16_301 ();
 sg13g2_decap_8 FILLER_16_308 ();
 sg13g2_decap_8 FILLER_16_315 ();
 sg13g2_decap_8 FILLER_16_322 ();
 sg13g2_decap_8 FILLER_16_329 ();
 sg13g2_decap_8 FILLER_16_336 ();
 sg13g2_decap_8 FILLER_16_343 ();
 sg13g2_decap_8 FILLER_16_350 ();
 sg13g2_decap_8 FILLER_16_357 ();
 sg13g2_decap_8 FILLER_16_364 ();
 sg13g2_decap_8 FILLER_16_371 ();
 sg13g2_decap_8 FILLER_16_378 ();
 sg13g2_decap_8 FILLER_16_385 ();
 sg13g2_decap_8 FILLER_16_392 ();
 sg13g2_decap_8 FILLER_16_399 ();
 sg13g2_fill_2 FILLER_16_406 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_decap_8 FILLER_17_168 ();
 sg13g2_decap_8 FILLER_17_175 ();
 sg13g2_decap_8 FILLER_17_182 ();
 sg13g2_decap_8 FILLER_17_189 ();
 sg13g2_decap_8 FILLER_17_196 ();
 sg13g2_decap_8 FILLER_17_203 ();
 sg13g2_decap_8 FILLER_17_210 ();
 sg13g2_decap_8 FILLER_17_217 ();
 sg13g2_decap_8 FILLER_17_224 ();
 sg13g2_decap_8 FILLER_17_231 ();
 sg13g2_decap_8 FILLER_17_238 ();
 sg13g2_decap_8 FILLER_17_245 ();
 sg13g2_decap_8 FILLER_17_252 ();
 sg13g2_decap_8 FILLER_17_259 ();
 sg13g2_decap_8 FILLER_17_266 ();
 sg13g2_decap_8 FILLER_17_273 ();
 sg13g2_decap_8 FILLER_17_280 ();
 sg13g2_decap_8 FILLER_17_287 ();
 sg13g2_decap_8 FILLER_17_294 ();
 sg13g2_decap_8 FILLER_17_301 ();
 sg13g2_decap_8 FILLER_17_308 ();
 sg13g2_decap_8 FILLER_17_315 ();
 sg13g2_decap_8 FILLER_17_322 ();
 sg13g2_decap_8 FILLER_17_329 ();
 sg13g2_decap_8 FILLER_17_336 ();
 sg13g2_decap_8 FILLER_17_343 ();
 sg13g2_decap_8 FILLER_17_350 ();
 sg13g2_decap_8 FILLER_17_357 ();
 sg13g2_decap_8 FILLER_17_364 ();
 sg13g2_decap_8 FILLER_17_371 ();
 sg13g2_decap_8 FILLER_17_378 ();
 sg13g2_decap_8 FILLER_17_385 ();
 sg13g2_decap_8 FILLER_17_392 ();
 sg13g2_decap_8 FILLER_17_399 ();
 sg13g2_fill_2 FILLER_17_406 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_decap_8 FILLER_18_147 ();
 sg13g2_decap_8 FILLER_18_154 ();
 sg13g2_decap_8 FILLER_18_161 ();
 sg13g2_decap_8 FILLER_18_168 ();
 sg13g2_decap_8 FILLER_18_175 ();
 sg13g2_decap_8 FILLER_18_182 ();
 sg13g2_decap_8 FILLER_18_189 ();
 sg13g2_decap_8 FILLER_18_196 ();
 sg13g2_decap_8 FILLER_18_203 ();
 sg13g2_decap_8 FILLER_18_210 ();
 sg13g2_decap_8 FILLER_18_217 ();
 sg13g2_decap_8 FILLER_18_224 ();
 sg13g2_decap_8 FILLER_18_231 ();
 sg13g2_decap_8 FILLER_18_238 ();
 sg13g2_decap_8 FILLER_18_245 ();
 sg13g2_decap_8 FILLER_18_252 ();
 sg13g2_decap_8 FILLER_18_259 ();
 sg13g2_decap_8 FILLER_18_266 ();
 sg13g2_decap_8 FILLER_18_273 ();
 sg13g2_decap_8 FILLER_18_280 ();
 sg13g2_decap_8 FILLER_18_287 ();
 sg13g2_decap_8 FILLER_18_294 ();
 sg13g2_decap_8 FILLER_18_301 ();
 sg13g2_decap_8 FILLER_18_308 ();
 sg13g2_decap_8 FILLER_18_315 ();
 sg13g2_decap_8 FILLER_18_322 ();
 sg13g2_decap_8 FILLER_18_329 ();
 sg13g2_decap_8 FILLER_18_336 ();
 sg13g2_decap_8 FILLER_18_343 ();
 sg13g2_decap_8 FILLER_18_350 ();
 sg13g2_decap_8 FILLER_18_357 ();
 sg13g2_decap_8 FILLER_18_364 ();
 sg13g2_decap_8 FILLER_18_371 ();
 sg13g2_decap_8 FILLER_18_378 ();
 sg13g2_decap_8 FILLER_18_385 ();
 sg13g2_decap_8 FILLER_18_392 ();
 sg13g2_decap_8 FILLER_18_399 ();
 sg13g2_fill_2 FILLER_18_406 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_decap_8 FILLER_19_140 ();
 sg13g2_decap_8 FILLER_19_147 ();
 sg13g2_decap_8 FILLER_19_154 ();
 sg13g2_decap_8 FILLER_19_161 ();
 sg13g2_decap_8 FILLER_19_168 ();
 sg13g2_decap_8 FILLER_19_175 ();
 sg13g2_decap_8 FILLER_19_182 ();
 sg13g2_decap_8 FILLER_19_189 ();
 sg13g2_decap_8 FILLER_19_196 ();
 sg13g2_decap_8 FILLER_19_203 ();
 sg13g2_decap_8 FILLER_19_210 ();
 sg13g2_decap_8 FILLER_19_217 ();
 sg13g2_decap_8 FILLER_19_224 ();
 sg13g2_decap_8 FILLER_19_231 ();
 sg13g2_decap_8 FILLER_19_238 ();
 sg13g2_decap_8 FILLER_19_245 ();
 sg13g2_decap_8 FILLER_19_252 ();
 sg13g2_decap_8 FILLER_19_259 ();
 sg13g2_decap_8 FILLER_19_266 ();
 sg13g2_decap_8 FILLER_19_273 ();
 sg13g2_decap_8 FILLER_19_280 ();
 sg13g2_decap_8 FILLER_19_287 ();
 sg13g2_decap_8 FILLER_19_294 ();
 sg13g2_decap_8 FILLER_19_301 ();
 sg13g2_decap_8 FILLER_19_308 ();
 sg13g2_decap_8 FILLER_19_315 ();
 sg13g2_decap_8 FILLER_19_322 ();
 sg13g2_decap_8 FILLER_19_329 ();
 sg13g2_decap_8 FILLER_19_336 ();
 sg13g2_decap_8 FILLER_19_343 ();
 sg13g2_decap_8 FILLER_19_350 ();
 sg13g2_decap_8 FILLER_19_357 ();
 sg13g2_decap_8 FILLER_19_364 ();
 sg13g2_decap_8 FILLER_19_371 ();
 sg13g2_decap_8 FILLER_19_378 ();
 sg13g2_decap_8 FILLER_19_385 ();
 sg13g2_decap_8 FILLER_19_392 ();
 sg13g2_decap_8 FILLER_19_399 ();
 sg13g2_fill_2 FILLER_19_406 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_decap_8 FILLER_20_126 ();
 sg13g2_decap_8 FILLER_20_133 ();
 sg13g2_decap_8 FILLER_20_140 ();
 sg13g2_decap_8 FILLER_20_147 ();
 sg13g2_decap_8 FILLER_20_154 ();
 sg13g2_decap_8 FILLER_20_161 ();
 sg13g2_decap_8 FILLER_20_168 ();
 sg13g2_decap_8 FILLER_20_175 ();
 sg13g2_decap_8 FILLER_20_182 ();
 sg13g2_decap_8 FILLER_20_189 ();
 sg13g2_decap_8 FILLER_20_196 ();
 sg13g2_decap_8 FILLER_20_203 ();
 sg13g2_decap_8 FILLER_20_210 ();
 sg13g2_decap_8 FILLER_20_217 ();
 sg13g2_decap_8 FILLER_20_224 ();
 sg13g2_decap_8 FILLER_20_231 ();
 sg13g2_decap_8 FILLER_20_238 ();
 sg13g2_decap_8 FILLER_20_245 ();
 sg13g2_decap_8 FILLER_20_252 ();
 sg13g2_decap_8 FILLER_20_259 ();
 sg13g2_decap_8 FILLER_20_266 ();
 sg13g2_decap_8 FILLER_20_273 ();
 sg13g2_decap_8 FILLER_20_280 ();
 sg13g2_decap_8 FILLER_20_287 ();
 sg13g2_decap_8 FILLER_20_294 ();
 sg13g2_decap_8 FILLER_20_301 ();
 sg13g2_decap_8 FILLER_20_308 ();
 sg13g2_decap_8 FILLER_20_315 ();
 sg13g2_decap_8 FILLER_20_322 ();
 sg13g2_decap_8 FILLER_20_329 ();
 sg13g2_decap_8 FILLER_20_336 ();
 sg13g2_decap_8 FILLER_20_343 ();
 sg13g2_decap_8 FILLER_20_350 ();
 sg13g2_decap_8 FILLER_20_357 ();
 sg13g2_decap_8 FILLER_20_364 ();
 sg13g2_decap_8 FILLER_20_371 ();
 sg13g2_decap_8 FILLER_20_378 ();
 sg13g2_decap_8 FILLER_20_385 ();
 sg13g2_decap_8 FILLER_20_392 ();
 sg13g2_decap_8 FILLER_20_399 ();
 sg13g2_fill_2 FILLER_20_406 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_decap_8 FILLER_21_119 ();
 sg13g2_decap_8 FILLER_21_126 ();
 sg13g2_decap_8 FILLER_21_133 ();
 sg13g2_decap_8 FILLER_21_140 ();
 sg13g2_decap_8 FILLER_21_147 ();
 sg13g2_decap_8 FILLER_21_154 ();
 sg13g2_decap_8 FILLER_21_161 ();
 sg13g2_decap_8 FILLER_21_168 ();
 sg13g2_decap_8 FILLER_21_175 ();
 sg13g2_decap_8 FILLER_21_182 ();
 sg13g2_decap_8 FILLER_21_189 ();
 sg13g2_decap_8 FILLER_21_196 ();
 sg13g2_decap_8 FILLER_21_203 ();
 sg13g2_decap_8 FILLER_21_210 ();
 sg13g2_decap_4 FILLER_21_217 ();
 sg13g2_fill_1 FILLER_21_221 ();
 sg13g2_decap_8 FILLER_21_226 ();
 sg13g2_decap_4 FILLER_21_233 ();
 sg13g2_fill_2 FILLER_21_263 ();
 sg13g2_decap_8 FILLER_21_292 ();
 sg13g2_decap_8 FILLER_21_299 ();
 sg13g2_decap_8 FILLER_21_306 ();
 sg13g2_decap_8 FILLER_21_313 ();
 sg13g2_decap_8 FILLER_21_320 ();
 sg13g2_decap_8 FILLER_21_327 ();
 sg13g2_decap_8 FILLER_21_334 ();
 sg13g2_decap_8 FILLER_21_341 ();
 sg13g2_decap_8 FILLER_21_348 ();
 sg13g2_decap_8 FILLER_21_355 ();
 sg13g2_decap_8 FILLER_21_362 ();
 sg13g2_decap_8 FILLER_21_369 ();
 sg13g2_decap_8 FILLER_21_376 ();
 sg13g2_decap_8 FILLER_21_383 ();
 sg13g2_decap_8 FILLER_21_390 ();
 sg13g2_decap_8 FILLER_21_397 ();
 sg13g2_decap_4 FILLER_21_404 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_8 FILLER_22_105 ();
 sg13g2_decap_8 FILLER_22_112 ();
 sg13g2_decap_8 FILLER_22_119 ();
 sg13g2_decap_8 FILLER_22_126 ();
 sg13g2_decap_8 FILLER_22_133 ();
 sg13g2_decap_8 FILLER_22_140 ();
 sg13g2_decap_8 FILLER_22_147 ();
 sg13g2_decap_8 FILLER_22_154 ();
 sg13g2_decap_8 FILLER_22_161 ();
 sg13g2_decap_8 FILLER_22_168 ();
 sg13g2_decap_8 FILLER_22_175 ();
 sg13g2_decap_8 FILLER_22_182 ();
 sg13g2_decap_8 FILLER_22_189 ();
 sg13g2_decap_4 FILLER_22_196 ();
 sg13g2_fill_1 FILLER_22_200 ();
 sg13g2_fill_2 FILLER_22_294 ();
 sg13g2_decap_8 FILLER_22_304 ();
 sg13g2_decap_4 FILLER_22_311 ();
 sg13g2_fill_2 FILLER_22_315 ();
 sg13g2_decap_8 FILLER_22_325 ();
 sg13g2_decap_8 FILLER_22_379 ();
 sg13g2_fill_1 FILLER_22_386 ();
 sg13g2_decap_8 FILLER_22_396 ();
 sg13g2_decap_4 FILLER_22_403 ();
 sg13g2_fill_2 FILLER_22_407 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_98 ();
 sg13g2_decap_8 FILLER_23_105 ();
 sg13g2_decap_8 FILLER_23_112 ();
 sg13g2_decap_8 FILLER_23_119 ();
 sg13g2_decap_8 FILLER_23_126 ();
 sg13g2_decap_8 FILLER_23_133 ();
 sg13g2_decap_8 FILLER_23_140 ();
 sg13g2_decap_8 FILLER_23_147 ();
 sg13g2_decap_8 FILLER_23_154 ();
 sg13g2_decap_8 FILLER_23_161 ();
 sg13g2_decap_8 FILLER_23_168 ();
 sg13g2_decap_8 FILLER_23_175 ();
 sg13g2_decap_8 FILLER_23_182 ();
 sg13g2_fill_1 FILLER_23_189 ();
 sg13g2_fill_2 FILLER_23_233 ();
 sg13g2_fill_1 FILLER_23_265 ();
 sg13g2_fill_1 FILLER_23_313 ();
 sg13g2_fill_2 FILLER_23_340 ();
 sg13g2_fill_2 FILLER_23_355 ();
 sg13g2_fill_1 FILLER_23_357 ();
 sg13g2_fill_2 FILLER_23_371 ();
 sg13g2_fill_1 FILLER_23_373 ();
 sg13g2_decap_8 FILLER_23_400 ();
 sg13g2_fill_2 FILLER_23_407 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_decap_8 FILLER_24_98 ();
 sg13g2_decap_8 FILLER_24_105 ();
 sg13g2_decap_8 FILLER_24_112 ();
 sg13g2_decap_8 FILLER_24_119 ();
 sg13g2_decap_8 FILLER_24_126 ();
 sg13g2_decap_8 FILLER_24_133 ();
 sg13g2_decap_8 FILLER_24_140 ();
 sg13g2_decap_8 FILLER_24_147 ();
 sg13g2_decap_8 FILLER_24_154 ();
 sg13g2_decap_8 FILLER_24_161 ();
 sg13g2_decap_8 FILLER_24_168 ();
 sg13g2_decap_8 FILLER_24_175 ();
 sg13g2_decap_4 FILLER_24_182 ();
 sg13g2_fill_1 FILLER_24_186 ();
 sg13g2_decap_4 FILLER_24_204 ();
 sg13g2_fill_1 FILLER_24_230 ();
 sg13g2_fill_1 FILLER_24_250 ();
 sg13g2_fill_1 FILLER_24_263 ();
 sg13g2_fill_1 FILLER_24_277 ();
 sg13g2_fill_2 FILLER_24_312 ();
 sg13g2_fill_2 FILLER_24_346 ();
 sg13g2_fill_1 FILLER_24_348 ();
 sg13g2_fill_2 FILLER_24_362 ();
 sg13g2_decap_8 FILLER_24_396 ();
 sg13g2_decap_4 FILLER_24_403 ();
 sg13g2_fill_2 FILLER_24_407 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_8 FILLER_25_91 ();
 sg13g2_decap_8 FILLER_25_98 ();
 sg13g2_decap_8 FILLER_25_105 ();
 sg13g2_decap_8 FILLER_25_112 ();
 sg13g2_decap_8 FILLER_25_119 ();
 sg13g2_decap_8 FILLER_25_126 ();
 sg13g2_decap_8 FILLER_25_133 ();
 sg13g2_decap_8 FILLER_25_140 ();
 sg13g2_decap_8 FILLER_25_147 ();
 sg13g2_decap_8 FILLER_25_154 ();
 sg13g2_decap_8 FILLER_25_161 ();
 sg13g2_decap_8 FILLER_25_168 ();
 sg13g2_decap_8 FILLER_25_175 ();
 sg13g2_decap_8 FILLER_25_182 ();
 sg13g2_fill_1 FILLER_25_189 ();
 sg13g2_decap_8 FILLER_25_251 ();
 sg13g2_decap_8 FILLER_25_261 ();
 sg13g2_fill_2 FILLER_25_268 ();
 sg13g2_decap_4 FILLER_25_278 ();
 sg13g2_fill_1 FILLER_25_282 ();
 sg13g2_fill_1 FILLER_25_318 ();
 sg13g2_fill_2 FILLER_25_352 ();
 sg13g2_fill_1 FILLER_25_354 ();
 sg13g2_fill_2 FILLER_25_374 ();
 sg13g2_decap_8 FILLER_25_402 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_decap_8 FILLER_26_91 ();
 sg13g2_decap_8 FILLER_26_98 ();
 sg13g2_decap_8 FILLER_26_105 ();
 sg13g2_decap_8 FILLER_26_112 ();
 sg13g2_decap_8 FILLER_26_119 ();
 sg13g2_decap_8 FILLER_26_126 ();
 sg13g2_decap_8 FILLER_26_133 ();
 sg13g2_decap_8 FILLER_26_140 ();
 sg13g2_decap_8 FILLER_26_147 ();
 sg13g2_decap_8 FILLER_26_154 ();
 sg13g2_decap_8 FILLER_26_161 ();
 sg13g2_decap_8 FILLER_26_168 ();
 sg13g2_decap_8 FILLER_26_175 ();
 sg13g2_fill_1 FILLER_26_182 ();
 sg13g2_fill_1 FILLER_26_209 ();
 sg13g2_decap_4 FILLER_26_219 ();
 sg13g2_fill_2 FILLER_26_231 ();
 sg13g2_fill_1 FILLER_26_233 ();
 sg13g2_fill_1 FILLER_26_260 ();
 sg13g2_fill_1 FILLER_26_301 ();
 sg13g2_fill_1 FILLER_26_311 ();
 sg13g2_fill_2 FILLER_26_325 ();
 sg13g2_fill_1 FILLER_26_327 ();
 sg13g2_fill_2 FILLER_26_340 ();
 sg13g2_decap_8 FILLER_26_393 ();
 sg13g2_decap_8 FILLER_26_400 ();
 sg13g2_fill_2 FILLER_26_407 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_decap_8 FILLER_27_84 ();
 sg13g2_decap_8 FILLER_27_91 ();
 sg13g2_decap_8 FILLER_27_98 ();
 sg13g2_decap_8 FILLER_27_105 ();
 sg13g2_decap_8 FILLER_27_112 ();
 sg13g2_decap_8 FILLER_27_119 ();
 sg13g2_decap_8 FILLER_27_126 ();
 sg13g2_decap_8 FILLER_27_133 ();
 sg13g2_decap_8 FILLER_27_140 ();
 sg13g2_decap_8 FILLER_27_147 ();
 sg13g2_decap_8 FILLER_27_154 ();
 sg13g2_decap_8 FILLER_27_161 ();
 sg13g2_decap_8 FILLER_27_168 ();
 sg13g2_decap_4 FILLER_27_175 ();
 sg13g2_fill_2 FILLER_27_179 ();
 sg13g2_fill_2 FILLER_27_215 ();
 sg13g2_decap_8 FILLER_27_260 ();
 sg13g2_fill_2 FILLER_27_267 ();
 sg13g2_fill_1 FILLER_27_269 ();
 sg13g2_fill_2 FILLER_27_331 ();
 sg13g2_fill_1 FILLER_27_360 ();
 sg13g2_fill_1 FILLER_27_378 ();
 sg13g2_decap_4 FILLER_27_405 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_decap_8 FILLER_28_84 ();
 sg13g2_decap_8 FILLER_28_91 ();
 sg13g2_decap_8 FILLER_28_98 ();
 sg13g2_decap_8 FILLER_28_105 ();
 sg13g2_decap_8 FILLER_28_112 ();
 sg13g2_decap_8 FILLER_28_119 ();
 sg13g2_decap_8 FILLER_28_126 ();
 sg13g2_decap_8 FILLER_28_133 ();
 sg13g2_decap_8 FILLER_28_140 ();
 sg13g2_decap_8 FILLER_28_147 ();
 sg13g2_decap_8 FILLER_28_154 ();
 sg13g2_decap_8 FILLER_28_161 ();
 sg13g2_decap_8 FILLER_28_168 ();
 sg13g2_decap_8 FILLER_28_175 ();
 sg13g2_fill_2 FILLER_28_182 ();
 sg13g2_fill_2 FILLER_28_224 ();
 sg13g2_fill_1 FILLER_28_226 ();
 sg13g2_decap_4 FILLER_28_239 ();
 sg13g2_fill_1 FILLER_28_243 ();
 sg13g2_fill_1 FILLER_28_249 ();
 sg13g2_fill_2 FILLER_28_259 ();
 sg13g2_fill_2 FILLER_28_266 ();
 sg13g2_decap_4 FILLER_28_273 ();
 sg13g2_fill_2 FILLER_28_324 ();
 sg13g2_fill_1 FILLER_28_326 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_decap_8 FILLER_29_84 ();
 sg13g2_decap_8 FILLER_29_91 ();
 sg13g2_decap_8 FILLER_29_98 ();
 sg13g2_decap_8 FILLER_29_105 ();
 sg13g2_decap_8 FILLER_29_112 ();
 sg13g2_decap_8 FILLER_29_119 ();
 sg13g2_decap_8 FILLER_29_126 ();
 sg13g2_decap_8 FILLER_29_133 ();
 sg13g2_decap_8 FILLER_29_140 ();
 sg13g2_decap_8 FILLER_29_147 ();
 sg13g2_decap_8 FILLER_29_154 ();
 sg13g2_decap_8 FILLER_29_161 ();
 sg13g2_decap_8 FILLER_29_168 ();
 sg13g2_decap_8 FILLER_29_175 ();
 sg13g2_decap_8 FILLER_29_182 ();
 sg13g2_fill_2 FILLER_29_189 ();
 sg13g2_fill_1 FILLER_29_191 ();
 sg13g2_decap_4 FILLER_29_202 ();
 sg13g2_decap_4 FILLER_29_239 ();
 sg13g2_decap_4 FILLER_29_289 ();
 sg13g2_fill_2 FILLER_29_293 ();
 sg13g2_fill_2 FILLER_29_302 ();
 sg13g2_decap_8 FILLER_29_322 ();
 sg13g2_decap_4 FILLER_29_329 ();
 sg13g2_decap_8 FILLER_29_337 ();
 sg13g2_fill_1 FILLER_29_354 ();
 sg13g2_fill_1 FILLER_29_390 ();
 sg13g2_fill_1 FILLER_29_408 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_77 ();
 sg13g2_decap_8 FILLER_30_84 ();
 sg13g2_decap_8 FILLER_30_91 ();
 sg13g2_decap_8 FILLER_30_98 ();
 sg13g2_decap_8 FILLER_30_105 ();
 sg13g2_decap_8 FILLER_30_112 ();
 sg13g2_decap_8 FILLER_30_119 ();
 sg13g2_decap_8 FILLER_30_126 ();
 sg13g2_decap_8 FILLER_30_133 ();
 sg13g2_decap_8 FILLER_30_140 ();
 sg13g2_decap_8 FILLER_30_147 ();
 sg13g2_decap_8 FILLER_30_154 ();
 sg13g2_decap_8 FILLER_30_161 ();
 sg13g2_decap_8 FILLER_30_168 ();
 sg13g2_decap_4 FILLER_30_175 ();
 sg13g2_fill_2 FILLER_30_179 ();
 sg13g2_decap_8 FILLER_30_211 ();
 sg13g2_decap_4 FILLER_30_218 ();
 sg13g2_fill_2 FILLER_30_222 ();
 sg13g2_decap_8 FILLER_30_230 ();
 sg13g2_fill_2 FILLER_30_237 ();
 sg13g2_fill_1 FILLER_30_239 ();
 sg13g2_fill_1 FILLER_30_246 ();
 sg13g2_fill_2 FILLER_30_251 ();
 sg13g2_fill_1 FILLER_30_253 ();
 sg13g2_decap_8 FILLER_30_259 ();
 sg13g2_fill_2 FILLER_30_266 ();
 sg13g2_fill_2 FILLER_30_280 ();
 sg13g2_fill_1 FILLER_30_282 ();
 sg13g2_fill_2 FILLER_30_309 ();
 sg13g2_decap_4 FILLER_30_324 ();
 sg13g2_fill_1 FILLER_30_328 ();
 sg13g2_fill_2 FILLER_30_346 ();
 sg13g2_fill_1 FILLER_30_348 ();
 sg13g2_fill_1 FILLER_30_361 ();
 sg13g2_fill_2 FILLER_30_380 ();
 sg13g2_fill_1 FILLER_30_408 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_decap_8 FILLER_31_84 ();
 sg13g2_decap_8 FILLER_31_91 ();
 sg13g2_decap_8 FILLER_31_98 ();
 sg13g2_decap_8 FILLER_31_105 ();
 sg13g2_decap_8 FILLER_31_112 ();
 sg13g2_decap_8 FILLER_31_119 ();
 sg13g2_decap_8 FILLER_31_126 ();
 sg13g2_decap_8 FILLER_31_133 ();
 sg13g2_decap_8 FILLER_31_140 ();
 sg13g2_decap_8 FILLER_31_147 ();
 sg13g2_decap_8 FILLER_31_154 ();
 sg13g2_decap_8 FILLER_31_161 ();
 sg13g2_decap_8 FILLER_31_168 ();
 sg13g2_decap_8 FILLER_31_175 ();
 sg13g2_decap_8 FILLER_31_182 ();
 sg13g2_decap_8 FILLER_31_198 ();
 sg13g2_decap_8 FILLER_31_205 ();
 sg13g2_fill_2 FILLER_31_216 ();
 sg13g2_fill_1 FILLER_31_218 ();
 sg13g2_fill_2 FILLER_31_234 ();
 sg13g2_fill_2 FILLER_31_256 ();
 sg13g2_fill_2 FILLER_31_268 ();
 sg13g2_fill_1 FILLER_31_270 ();
 sg13g2_decap_8 FILLER_31_288 ();
 sg13g2_decap_8 FILLER_31_299 ();
 sg13g2_decap_8 FILLER_31_306 ();
 sg13g2_fill_1 FILLER_31_313 ();
 sg13g2_decap_8 FILLER_31_319 ();
 sg13g2_fill_1 FILLER_31_326 ();
 sg13g2_fill_1 FILLER_31_350 ();
 sg13g2_decap_8 FILLER_31_355 ();
 sg13g2_fill_2 FILLER_31_392 ();
 sg13g2_fill_1 FILLER_31_408 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_8 FILLER_32_84 ();
 sg13g2_decap_8 FILLER_32_91 ();
 sg13g2_decap_8 FILLER_32_98 ();
 sg13g2_decap_8 FILLER_32_105 ();
 sg13g2_decap_8 FILLER_32_112 ();
 sg13g2_decap_8 FILLER_32_119 ();
 sg13g2_decap_8 FILLER_32_126 ();
 sg13g2_decap_8 FILLER_32_133 ();
 sg13g2_decap_8 FILLER_32_140 ();
 sg13g2_decap_8 FILLER_32_147 ();
 sg13g2_decap_8 FILLER_32_154 ();
 sg13g2_decap_8 FILLER_32_161 ();
 sg13g2_decap_8 FILLER_32_168 ();
 sg13g2_decap_8 FILLER_32_175 ();
 sg13g2_decap_8 FILLER_32_182 ();
 sg13g2_fill_2 FILLER_32_189 ();
 sg13g2_fill_1 FILLER_32_191 ();
 sg13g2_fill_2 FILLER_32_203 ();
 sg13g2_fill_2 FILLER_32_220 ();
 sg13g2_fill_2 FILLER_32_231 ();
 sg13g2_fill_1 FILLER_32_233 ();
 sg13g2_decap_4 FILLER_32_252 ();
 sg13g2_fill_2 FILLER_32_256 ();
 sg13g2_fill_1 FILLER_32_269 ();
 sg13g2_decap_8 FILLER_32_279 ();
 sg13g2_fill_2 FILLER_32_286 ();
 sg13g2_fill_1 FILLER_32_288 ();
 sg13g2_fill_1 FILLER_32_318 ();
 sg13g2_decap_4 FILLER_32_339 ();
 sg13g2_decap_8 FILLER_32_394 ();
 sg13g2_decap_8 FILLER_32_401 ();
 sg13g2_fill_1 FILLER_32_408 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_decap_8 FILLER_33_91 ();
 sg13g2_decap_8 FILLER_33_98 ();
 sg13g2_decap_8 FILLER_33_105 ();
 sg13g2_decap_8 FILLER_33_112 ();
 sg13g2_decap_8 FILLER_33_119 ();
 sg13g2_decap_8 FILLER_33_126 ();
 sg13g2_decap_8 FILLER_33_133 ();
 sg13g2_decap_8 FILLER_33_140 ();
 sg13g2_decap_8 FILLER_33_147 ();
 sg13g2_decap_8 FILLER_33_154 ();
 sg13g2_decap_8 FILLER_33_161 ();
 sg13g2_decap_8 FILLER_33_168 ();
 sg13g2_decap_8 FILLER_33_175 ();
 sg13g2_decap_4 FILLER_33_182 ();
 sg13g2_fill_1 FILLER_33_186 ();
 sg13g2_decap_8 FILLER_33_212 ();
 sg13g2_fill_1 FILLER_33_219 ();
 sg13g2_decap_4 FILLER_33_225 ();
 sg13g2_decap_8 FILLER_33_235 ();
 sg13g2_fill_2 FILLER_33_251 ();
 sg13g2_fill_1 FILLER_33_260 ();
 sg13g2_fill_1 FILLER_33_286 ();
 sg13g2_fill_2 FILLER_33_295 ();
 sg13g2_decap_8 FILLER_33_318 ();
 sg13g2_decap_4 FILLER_33_325 ();
 sg13g2_fill_1 FILLER_33_329 ();
 sg13g2_fill_2 FILLER_33_344 ();
 sg13g2_fill_1 FILLER_33_346 ();
 sg13g2_fill_2 FILLER_33_356 ();
 sg13g2_decap_8 FILLER_33_397 ();
 sg13g2_decap_4 FILLER_33_404 ();
 sg13g2_fill_1 FILLER_33_408 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_decap_8 FILLER_34_91 ();
 sg13g2_decap_8 FILLER_34_98 ();
 sg13g2_decap_8 FILLER_34_105 ();
 sg13g2_decap_8 FILLER_34_112 ();
 sg13g2_decap_8 FILLER_34_119 ();
 sg13g2_decap_8 FILLER_34_126 ();
 sg13g2_decap_8 FILLER_34_133 ();
 sg13g2_decap_8 FILLER_34_140 ();
 sg13g2_decap_8 FILLER_34_147 ();
 sg13g2_decap_8 FILLER_34_154 ();
 sg13g2_decap_8 FILLER_34_161 ();
 sg13g2_decap_8 FILLER_34_168 ();
 sg13g2_decap_8 FILLER_34_175 ();
 sg13g2_decap_8 FILLER_34_182 ();
 sg13g2_fill_2 FILLER_34_189 ();
 sg13g2_decap_4 FILLER_34_206 ();
 sg13g2_fill_2 FILLER_34_237 ();
 sg13g2_fill_2 FILLER_34_254 ();
 sg13g2_fill_1 FILLER_34_256 ();
 sg13g2_decap_8 FILLER_34_263 ();
 sg13g2_fill_1 FILLER_34_270 ();
 sg13g2_decap_4 FILLER_34_280 ();
 sg13g2_fill_2 FILLER_34_326 ();
 sg13g2_fill_1 FILLER_34_328 ();
 sg13g2_decap_8 FILLER_34_399 ();
 sg13g2_fill_2 FILLER_34_406 ();
 sg13g2_fill_1 FILLER_34_408 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_decap_8 FILLER_35_98 ();
 sg13g2_decap_8 FILLER_35_105 ();
 sg13g2_decap_8 FILLER_35_112 ();
 sg13g2_decap_8 FILLER_35_119 ();
 sg13g2_decap_8 FILLER_35_126 ();
 sg13g2_decap_8 FILLER_35_133 ();
 sg13g2_decap_8 FILLER_35_140 ();
 sg13g2_decap_8 FILLER_35_147 ();
 sg13g2_decap_8 FILLER_35_154 ();
 sg13g2_decap_8 FILLER_35_161 ();
 sg13g2_decap_8 FILLER_35_168 ();
 sg13g2_decap_8 FILLER_35_175 ();
 sg13g2_decap_8 FILLER_35_182 ();
 sg13g2_decap_8 FILLER_35_189 ();
 sg13g2_fill_2 FILLER_35_196 ();
 sg13g2_decap_8 FILLER_35_206 ();
 sg13g2_fill_2 FILLER_35_213 ();
 sg13g2_fill_2 FILLER_35_220 ();
 sg13g2_fill_2 FILLER_35_232 ();
 sg13g2_fill_1 FILLER_35_234 ();
 sg13g2_fill_1 FILLER_35_252 ();
 sg13g2_fill_1 FILLER_35_259 ();
 sg13g2_decap_4 FILLER_35_267 ();
 sg13g2_fill_1 FILLER_35_271 ();
 sg13g2_decap_8 FILLER_35_284 ();
 sg13g2_decap_4 FILLER_35_296 ();
 sg13g2_fill_2 FILLER_35_300 ();
 sg13g2_decap_8 FILLER_35_387 ();
 sg13g2_decap_8 FILLER_35_394 ();
 sg13g2_decap_8 FILLER_35_401 ();
 sg13g2_fill_1 FILLER_35_408 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_decap_8 FILLER_36_112 ();
 sg13g2_decap_8 FILLER_36_119 ();
 sg13g2_decap_8 FILLER_36_126 ();
 sg13g2_decap_8 FILLER_36_133 ();
 sg13g2_decap_8 FILLER_36_140 ();
 sg13g2_decap_8 FILLER_36_147 ();
 sg13g2_decap_8 FILLER_36_154 ();
 sg13g2_decap_8 FILLER_36_161 ();
 sg13g2_decap_8 FILLER_36_168 ();
 sg13g2_decap_8 FILLER_36_175 ();
 sg13g2_decap_8 FILLER_36_182 ();
 sg13g2_decap_8 FILLER_36_189 ();
 sg13g2_fill_2 FILLER_36_208 ();
 sg13g2_fill_2 FILLER_36_230 ();
 sg13g2_fill_1 FILLER_36_232 ();
 sg13g2_fill_2 FILLER_36_237 ();
 sg13g2_decap_8 FILLER_36_252 ();
 sg13g2_fill_2 FILLER_36_281 ();
 sg13g2_fill_1 FILLER_36_283 ();
 sg13g2_fill_2 FILLER_36_323 ();
 sg13g2_fill_1 FILLER_36_325 ();
 sg13g2_decap_8 FILLER_36_391 ();
 sg13g2_decap_8 FILLER_36_398 ();
 sg13g2_decap_4 FILLER_36_405 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_8 FILLER_37_112 ();
 sg13g2_decap_8 FILLER_37_119 ();
 sg13g2_decap_8 FILLER_37_126 ();
 sg13g2_decap_8 FILLER_37_133 ();
 sg13g2_decap_8 FILLER_37_140 ();
 sg13g2_decap_8 FILLER_37_147 ();
 sg13g2_decap_8 FILLER_37_154 ();
 sg13g2_decap_8 FILLER_37_161 ();
 sg13g2_decap_8 FILLER_37_168 ();
 sg13g2_decap_8 FILLER_37_175 ();
 sg13g2_decap_8 FILLER_37_182 ();
 sg13g2_decap_4 FILLER_37_189 ();
 sg13g2_fill_1 FILLER_37_193 ();
 sg13g2_fill_2 FILLER_37_230 ();
 sg13g2_fill_1 FILLER_37_241 ();
 sg13g2_fill_1 FILLER_37_270 ();
 sg13g2_fill_2 FILLER_37_285 ();
 sg13g2_decap_8 FILLER_37_402 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_4 FILLER_38_60 ();
 sg13g2_decap_4 FILLER_38_68 ();
 sg13g2_decap_4 FILLER_38_76 ();
 sg13g2_decap_4 FILLER_38_84 ();
 sg13g2_decap_4 FILLER_38_92 ();
 sg13g2_decap_4 FILLER_38_100 ();
 sg13g2_decap_4 FILLER_38_108 ();
 sg13g2_decap_4 FILLER_38_116 ();
 sg13g2_decap_4 FILLER_38_124 ();
 sg13g2_decap_4 FILLER_38_132 ();
 sg13g2_decap_4 FILLER_38_140 ();
 sg13g2_decap_4 FILLER_38_148 ();
 sg13g2_decap_4 FILLER_38_156 ();
 sg13g2_decap_4 FILLER_38_164 ();
 sg13g2_decap_4 FILLER_38_172 ();
 sg13g2_decap_8 FILLER_38_180 ();
 sg13g2_decap_8 FILLER_38_187 ();
 sg13g2_decap_8 FILLER_38_194 ();
 sg13g2_decap_4 FILLER_38_201 ();
 sg13g2_fill_1 FILLER_38_205 ();
 sg13g2_fill_1 FILLER_38_210 ();
 sg13g2_decap_8 FILLER_38_216 ();
 sg13g2_fill_2 FILLER_38_223 ();
 sg13g2_decap_8 FILLER_38_237 ();
 sg13g2_decap_8 FILLER_38_244 ();
 sg13g2_fill_2 FILLER_38_255 ();
 sg13g2_fill_1 FILLER_38_257 ();
 sg13g2_fill_1 FILLER_38_268 ();
 sg13g2_decap_4 FILLER_38_284 ();
 sg13g2_fill_2 FILLER_38_288 ();
 sg13g2_fill_1 FILLER_38_343 ();
 sg13g2_fill_2 FILLER_38_360 ();
 sg13g2_fill_2 FILLER_38_407 ();
 assign uio_oe[0] = net7;
 assign uio_oe[1] = net8;
 assign uio_oe[2] = net9;
 assign uio_oe[3] = net10;
 assign uio_oe[4] = net11;
 assign uio_oe[5] = net12;
 assign uio_oe[6] = net13;
 assign uio_oe[7] = net14;
 assign uio_out[0] = net15;
 assign uio_out[1] = net16;
 assign uio_out[2] = net17;
 assign uio_out[3] = net18;
 assign uio_out[4] = net19;
 assign uio_out[5] = net20;
 assign uio_out[6] = net21;
 assign uio_out[7] = net22;
endmodule

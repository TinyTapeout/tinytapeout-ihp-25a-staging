module tt_um_neural_navigators (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire clk_regs;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire \u_toplayer.delay_counter_layer1[0] ;
 wire \u_toplayer.delay_counter_layer1[1] ;
 wire \u_toplayer.delay_counter_layer2[0] ;
 wire \u_toplayer.delay_counter_layer2[1] ;
 wire \u_toplayer.delay_counter_layer3[0] ;
 wire \u_toplayer.delay_counter_layer3[1] ;
 wire \u_toplayer.delayed_done_layer1 ;
 wire \u_toplayer.delayed_done_layer2 ;
 wire \u_toplayer.delayed_done_layer3 ;
 wire \u_toplayer.done_layer1 ;
 wire \u_toplayer.done_layer2 ;
 wire \u_toplayer.done_layer3 ;
 wire \u_toplayer.outreg[0] ;
 wire \u_toplayer.outreg[10] ;
 wire \u_toplayer.outreg[11] ;
 wire \u_toplayer.outreg[12] ;
 wire \u_toplayer.outreg[13] ;
 wire \u_toplayer.outreg[14] ;
 wire \u_toplayer.outreg[15] ;
 wire \u_toplayer.outreg[16] ;
 wire \u_toplayer.outreg[17] ;
 wire \u_toplayer.outreg[18] ;
 wire \u_toplayer.outreg[19] ;
 wire \u_toplayer.outreg[1] ;
 wire \u_toplayer.outreg[20] ;
 wire \u_toplayer.outreg[21] ;
 wire \u_toplayer.outreg[22] ;
 wire \u_toplayer.outreg[23] ;
 wire \u_toplayer.outreg[24] ;
 wire \u_toplayer.outreg[25] ;
 wire \u_toplayer.outreg[26] ;
 wire \u_toplayer.outreg[27] ;
 wire \u_toplayer.outreg[28] ;
 wire \u_toplayer.outreg[29] ;
 wire \u_toplayer.outreg[2] ;
 wire \u_toplayer.outreg[30] ;
 wire \u_toplayer.outreg[31] ;
 wire \u_toplayer.outreg[32] ;
 wire \u_toplayer.outreg[33] ;
 wire \u_toplayer.outreg[34] ;
 wire \u_toplayer.outreg[35] ;
 wire \u_toplayer.outreg[36] ;
 wire \u_toplayer.outreg[37] ;
 wire \u_toplayer.outreg[38] ;
 wire \u_toplayer.outreg[39] ;
 wire \u_toplayer.outreg[3] ;
 wire \u_toplayer.outreg[40] ;
 wire \u_toplayer.outreg[41] ;
 wire \u_toplayer.outreg[42] ;
 wire \u_toplayer.outreg[43] ;
 wire \u_toplayer.outreg[44] ;
 wire \u_toplayer.outreg[45] ;
 wire \u_toplayer.outreg[46] ;
 wire \u_toplayer.outreg[47] ;
 wire \u_toplayer.outreg[48] ;
 wire \u_toplayer.outreg[49] ;
 wire \u_toplayer.outreg[4] ;
 wire \u_toplayer.outreg[50] ;
 wire \u_toplayer.outreg[51] ;
 wire \u_toplayer.outreg[52] ;
 wire \u_toplayer.outreg[53] ;
 wire \u_toplayer.outreg[54] ;
 wire \u_toplayer.outreg[55] ;
 wire \u_toplayer.outreg[56] ;
 wire \u_toplayer.outreg[57] ;
 wire \u_toplayer.outreg[58] ;
 wire \u_toplayer.outreg[59] ;
 wire \u_toplayer.outreg[5] ;
 wire \u_toplayer.outreg[60] ;
 wire \u_toplayer.outreg[61] ;
 wire \u_toplayer.outreg[62] ;
 wire \u_toplayer.outreg[63] ;
 wire \u_toplayer.outreg[64] ;
 wire \u_toplayer.outreg[65] ;
 wire \u_toplayer.outreg[66] ;
 wire \u_toplayer.outreg[67] ;
 wire \u_toplayer.outreg[68] ;
 wire \u_toplayer.outreg[69] ;
 wire \u_toplayer.outreg[6] ;
 wire \u_toplayer.outreg[70] ;
 wire \u_toplayer.outreg[71] ;
 wire \u_toplayer.outreg[72] ;
 wire \u_toplayer.outreg[73] ;
 wire \u_toplayer.outreg[74] ;
 wire \u_toplayer.outreg[75] ;
 wire \u_toplayer.outreg[76] ;
 wire \u_toplayer.outreg[77] ;
 wire \u_toplayer.outreg[78] ;
 wire \u_toplayer.outreg[79] ;
 wire \u_toplayer.outreg[7] ;
 wire \u_toplayer.outreg[8] ;
 wire \u_toplayer.outreg[9] ;
 wire \u_toplayer.reg_layer1[0] ;
 wire \u_toplayer.reg_layer1[100] ;
 wire \u_toplayer.reg_layer1[101] ;
 wire \u_toplayer.reg_layer1[102] ;
 wire \u_toplayer.reg_layer1[103] ;
 wire \u_toplayer.reg_layer1[104] ;
 wire \u_toplayer.reg_layer1[105] ;
 wire \u_toplayer.reg_layer1[106] ;
 wire \u_toplayer.reg_layer1[107] ;
 wire \u_toplayer.reg_layer1[108] ;
 wire \u_toplayer.reg_layer1[109] ;
 wire \u_toplayer.reg_layer1[10] ;
 wire \u_toplayer.reg_layer1[110] ;
 wire \u_toplayer.reg_layer1[111] ;
 wire \u_toplayer.reg_layer1[112] ;
 wire \u_toplayer.reg_layer1[113] ;
 wire \u_toplayer.reg_layer1[114] ;
 wire \u_toplayer.reg_layer1[115] ;
 wire \u_toplayer.reg_layer1[116] ;
 wire \u_toplayer.reg_layer1[117] ;
 wire \u_toplayer.reg_layer1[118] ;
 wire \u_toplayer.reg_layer1[119] ;
 wire \u_toplayer.reg_layer1[11] ;
 wire \u_toplayer.reg_layer1[120] ;
 wire \u_toplayer.reg_layer1[121] ;
 wire \u_toplayer.reg_layer1[122] ;
 wire \u_toplayer.reg_layer1[123] ;
 wire \u_toplayer.reg_layer1[124] ;
 wire \u_toplayer.reg_layer1[125] ;
 wire \u_toplayer.reg_layer1[126] ;
 wire \u_toplayer.reg_layer1[127] ;
 wire \u_toplayer.reg_layer1[128] ;
 wire \u_toplayer.reg_layer1[129] ;
 wire \u_toplayer.reg_layer1[12] ;
 wire \u_toplayer.reg_layer1[130] ;
 wire \u_toplayer.reg_layer1[131] ;
 wire \u_toplayer.reg_layer1[132] ;
 wire \u_toplayer.reg_layer1[133] ;
 wire \u_toplayer.reg_layer1[134] ;
 wire \u_toplayer.reg_layer1[135] ;
 wire \u_toplayer.reg_layer1[136] ;
 wire \u_toplayer.reg_layer1[137] ;
 wire \u_toplayer.reg_layer1[138] ;
 wire \u_toplayer.reg_layer1[139] ;
 wire \u_toplayer.reg_layer1[13] ;
 wire \u_toplayer.reg_layer1[140] ;
 wire \u_toplayer.reg_layer1[141] ;
 wire \u_toplayer.reg_layer1[142] ;
 wire \u_toplayer.reg_layer1[143] ;
 wire \u_toplayer.reg_layer1[144] ;
 wire \u_toplayer.reg_layer1[145] ;
 wire \u_toplayer.reg_layer1[146] ;
 wire \u_toplayer.reg_layer1[147] ;
 wire \u_toplayer.reg_layer1[148] ;
 wire \u_toplayer.reg_layer1[149] ;
 wire \u_toplayer.reg_layer1[14] ;
 wire \u_toplayer.reg_layer1[150] ;
 wire \u_toplayer.reg_layer1[151] ;
 wire \u_toplayer.reg_layer1[152] ;
 wire \u_toplayer.reg_layer1[153] ;
 wire \u_toplayer.reg_layer1[154] ;
 wire \u_toplayer.reg_layer1[155] ;
 wire \u_toplayer.reg_layer1[156] ;
 wire \u_toplayer.reg_layer1[157] ;
 wire \u_toplayer.reg_layer1[158] ;
 wire \u_toplayer.reg_layer1[159] ;
 wire \u_toplayer.reg_layer1[15] ;
 wire \u_toplayer.reg_layer1[160] ;
 wire \u_toplayer.reg_layer1[161] ;
 wire \u_toplayer.reg_layer1[162] ;
 wire \u_toplayer.reg_layer1[163] ;
 wire \u_toplayer.reg_layer1[164] ;
 wire \u_toplayer.reg_layer1[165] ;
 wire \u_toplayer.reg_layer1[166] ;
 wire \u_toplayer.reg_layer1[167] ;
 wire \u_toplayer.reg_layer1[168] ;
 wire \u_toplayer.reg_layer1[169] ;
 wire \u_toplayer.reg_layer1[16] ;
 wire \u_toplayer.reg_layer1[170] ;
 wire \u_toplayer.reg_layer1[171] ;
 wire \u_toplayer.reg_layer1[172] ;
 wire \u_toplayer.reg_layer1[173] ;
 wire \u_toplayer.reg_layer1[174] ;
 wire \u_toplayer.reg_layer1[175] ;
 wire \u_toplayer.reg_layer1[176] ;
 wire \u_toplayer.reg_layer1[177] ;
 wire \u_toplayer.reg_layer1[178] ;
 wire \u_toplayer.reg_layer1[179] ;
 wire \u_toplayer.reg_layer1[17] ;
 wire \u_toplayer.reg_layer1[180] ;
 wire \u_toplayer.reg_layer1[181] ;
 wire \u_toplayer.reg_layer1[182] ;
 wire \u_toplayer.reg_layer1[183] ;
 wire \u_toplayer.reg_layer1[184] ;
 wire \u_toplayer.reg_layer1[185] ;
 wire \u_toplayer.reg_layer1[186] ;
 wire \u_toplayer.reg_layer1[187] ;
 wire \u_toplayer.reg_layer1[188] ;
 wire \u_toplayer.reg_layer1[189] ;
 wire \u_toplayer.reg_layer1[18] ;
 wire \u_toplayer.reg_layer1[190] ;
 wire \u_toplayer.reg_layer1[191] ;
 wire \u_toplayer.reg_layer1[192] ;
 wire \u_toplayer.reg_layer1[193] ;
 wire \u_toplayer.reg_layer1[194] ;
 wire \u_toplayer.reg_layer1[195] ;
 wire \u_toplayer.reg_layer1[196] ;
 wire \u_toplayer.reg_layer1[197] ;
 wire \u_toplayer.reg_layer1[198] ;
 wire \u_toplayer.reg_layer1[199] ;
 wire \u_toplayer.reg_layer1[19] ;
 wire \u_toplayer.reg_layer1[1] ;
 wire \u_toplayer.reg_layer1[200] ;
 wire \u_toplayer.reg_layer1[201] ;
 wire \u_toplayer.reg_layer1[202] ;
 wire \u_toplayer.reg_layer1[203] ;
 wire \u_toplayer.reg_layer1[204] ;
 wire \u_toplayer.reg_layer1[205] ;
 wire \u_toplayer.reg_layer1[206] ;
 wire \u_toplayer.reg_layer1[207] ;
 wire \u_toplayer.reg_layer1[208] ;
 wire \u_toplayer.reg_layer1[209] ;
 wire \u_toplayer.reg_layer1[20] ;
 wire \u_toplayer.reg_layer1[210] ;
 wire \u_toplayer.reg_layer1[211] ;
 wire \u_toplayer.reg_layer1[212] ;
 wire \u_toplayer.reg_layer1[213] ;
 wire \u_toplayer.reg_layer1[214] ;
 wire \u_toplayer.reg_layer1[215] ;
 wire \u_toplayer.reg_layer1[216] ;
 wire \u_toplayer.reg_layer1[217] ;
 wire \u_toplayer.reg_layer1[218] ;
 wire \u_toplayer.reg_layer1[219] ;
 wire \u_toplayer.reg_layer1[21] ;
 wire \u_toplayer.reg_layer1[220] ;
 wire \u_toplayer.reg_layer1[221] ;
 wire \u_toplayer.reg_layer1[222] ;
 wire \u_toplayer.reg_layer1[223] ;
 wire \u_toplayer.reg_layer1[224] ;
 wire \u_toplayer.reg_layer1[225] ;
 wire \u_toplayer.reg_layer1[226] ;
 wire \u_toplayer.reg_layer1[227] ;
 wire \u_toplayer.reg_layer1[228] ;
 wire \u_toplayer.reg_layer1[229] ;
 wire \u_toplayer.reg_layer1[22] ;
 wire \u_toplayer.reg_layer1[230] ;
 wire \u_toplayer.reg_layer1[231] ;
 wire \u_toplayer.reg_layer1[232] ;
 wire \u_toplayer.reg_layer1[233] ;
 wire \u_toplayer.reg_layer1[234] ;
 wire \u_toplayer.reg_layer1[235] ;
 wire \u_toplayer.reg_layer1[236] ;
 wire \u_toplayer.reg_layer1[237] ;
 wire \u_toplayer.reg_layer1[238] ;
 wire \u_toplayer.reg_layer1[239] ;
 wire \u_toplayer.reg_layer1[23] ;
 wire \u_toplayer.reg_layer1[240] ;
 wire \u_toplayer.reg_layer1[241] ;
 wire \u_toplayer.reg_layer1[242] ;
 wire \u_toplayer.reg_layer1[243] ;
 wire \u_toplayer.reg_layer1[244] ;
 wire \u_toplayer.reg_layer1[245] ;
 wire \u_toplayer.reg_layer1[246] ;
 wire \u_toplayer.reg_layer1[247] ;
 wire \u_toplayer.reg_layer1[248] ;
 wire \u_toplayer.reg_layer1[249] ;
 wire \u_toplayer.reg_layer1[24] ;
 wire \u_toplayer.reg_layer1[250] ;
 wire \u_toplayer.reg_layer1[251] ;
 wire \u_toplayer.reg_layer1[252] ;
 wire \u_toplayer.reg_layer1[253] ;
 wire \u_toplayer.reg_layer1[254] ;
 wire \u_toplayer.reg_layer1[255] ;
 wire \u_toplayer.reg_layer1[25] ;
 wire \u_toplayer.reg_layer1[26] ;
 wire \u_toplayer.reg_layer1[27] ;
 wire \u_toplayer.reg_layer1[28] ;
 wire \u_toplayer.reg_layer1[29] ;
 wire \u_toplayer.reg_layer1[2] ;
 wire \u_toplayer.reg_layer1[30] ;
 wire \u_toplayer.reg_layer1[31] ;
 wire \u_toplayer.reg_layer1[32] ;
 wire \u_toplayer.reg_layer1[33] ;
 wire \u_toplayer.reg_layer1[34] ;
 wire \u_toplayer.reg_layer1[35] ;
 wire \u_toplayer.reg_layer1[36] ;
 wire \u_toplayer.reg_layer1[37] ;
 wire \u_toplayer.reg_layer1[38] ;
 wire \u_toplayer.reg_layer1[39] ;
 wire \u_toplayer.reg_layer1[3] ;
 wire \u_toplayer.reg_layer1[40] ;
 wire \u_toplayer.reg_layer1[41] ;
 wire \u_toplayer.reg_layer1[42] ;
 wire \u_toplayer.reg_layer1[43] ;
 wire \u_toplayer.reg_layer1[44] ;
 wire \u_toplayer.reg_layer1[45] ;
 wire \u_toplayer.reg_layer1[46] ;
 wire \u_toplayer.reg_layer1[47] ;
 wire \u_toplayer.reg_layer1[48] ;
 wire \u_toplayer.reg_layer1[49] ;
 wire \u_toplayer.reg_layer1[4] ;
 wire \u_toplayer.reg_layer1[50] ;
 wire \u_toplayer.reg_layer1[51] ;
 wire \u_toplayer.reg_layer1[52] ;
 wire \u_toplayer.reg_layer1[53] ;
 wire \u_toplayer.reg_layer1[54] ;
 wire \u_toplayer.reg_layer1[55] ;
 wire \u_toplayer.reg_layer1[56] ;
 wire \u_toplayer.reg_layer1[57] ;
 wire \u_toplayer.reg_layer1[58] ;
 wire \u_toplayer.reg_layer1[59] ;
 wire \u_toplayer.reg_layer1[5] ;
 wire \u_toplayer.reg_layer1[60] ;
 wire \u_toplayer.reg_layer1[61] ;
 wire \u_toplayer.reg_layer1[62] ;
 wire \u_toplayer.reg_layer1[63] ;
 wire \u_toplayer.reg_layer1[64] ;
 wire \u_toplayer.reg_layer1[65] ;
 wire \u_toplayer.reg_layer1[66] ;
 wire \u_toplayer.reg_layer1[67] ;
 wire \u_toplayer.reg_layer1[68] ;
 wire \u_toplayer.reg_layer1[69] ;
 wire \u_toplayer.reg_layer1[6] ;
 wire \u_toplayer.reg_layer1[70] ;
 wire \u_toplayer.reg_layer1[71] ;
 wire \u_toplayer.reg_layer1[72] ;
 wire \u_toplayer.reg_layer1[73] ;
 wire \u_toplayer.reg_layer1[74] ;
 wire \u_toplayer.reg_layer1[75] ;
 wire \u_toplayer.reg_layer1[76] ;
 wire \u_toplayer.reg_layer1[77] ;
 wire \u_toplayer.reg_layer1[78] ;
 wire \u_toplayer.reg_layer1[79] ;
 wire \u_toplayer.reg_layer1[7] ;
 wire \u_toplayer.reg_layer1[80] ;
 wire \u_toplayer.reg_layer1[81] ;
 wire \u_toplayer.reg_layer1[82] ;
 wire \u_toplayer.reg_layer1[83] ;
 wire \u_toplayer.reg_layer1[84] ;
 wire \u_toplayer.reg_layer1[85] ;
 wire \u_toplayer.reg_layer1[86] ;
 wire \u_toplayer.reg_layer1[87] ;
 wire \u_toplayer.reg_layer1[88] ;
 wire \u_toplayer.reg_layer1[89] ;
 wire \u_toplayer.reg_layer1[8] ;
 wire \u_toplayer.reg_layer1[90] ;
 wire \u_toplayer.reg_layer1[91] ;
 wire \u_toplayer.reg_layer1[92] ;
 wire \u_toplayer.reg_layer1[93] ;
 wire \u_toplayer.reg_layer1[94] ;
 wire \u_toplayer.reg_layer1[95] ;
 wire \u_toplayer.reg_layer1[96] ;
 wire \u_toplayer.reg_layer1[97] ;
 wire \u_toplayer.reg_layer1[98] ;
 wire \u_toplayer.reg_layer1[99] ;
 wire \u_toplayer.reg_layer1[9] ;
 wire \u_toplayer.reg_layer2[0] ;
 wire \u_toplayer.reg_layer2[100] ;
 wire \u_toplayer.reg_layer2[101] ;
 wire \u_toplayer.reg_layer2[102] ;
 wire \u_toplayer.reg_layer2[103] ;
 wire \u_toplayer.reg_layer2[104] ;
 wire \u_toplayer.reg_layer2[105] ;
 wire \u_toplayer.reg_layer2[106] ;
 wire \u_toplayer.reg_layer2[107] ;
 wire \u_toplayer.reg_layer2[108] ;
 wire \u_toplayer.reg_layer2[109] ;
 wire \u_toplayer.reg_layer2[10] ;
 wire \u_toplayer.reg_layer2[110] ;
 wire \u_toplayer.reg_layer2[111] ;
 wire \u_toplayer.reg_layer2[112] ;
 wire \u_toplayer.reg_layer2[113] ;
 wire \u_toplayer.reg_layer2[114] ;
 wire \u_toplayer.reg_layer2[115] ;
 wire \u_toplayer.reg_layer2[116] ;
 wire \u_toplayer.reg_layer2[117] ;
 wire \u_toplayer.reg_layer2[118] ;
 wire \u_toplayer.reg_layer2[119] ;
 wire \u_toplayer.reg_layer2[11] ;
 wire \u_toplayer.reg_layer2[120] ;
 wire \u_toplayer.reg_layer2[121] ;
 wire \u_toplayer.reg_layer2[122] ;
 wire \u_toplayer.reg_layer2[123] ;
 wire \u_toplayer.reg_layer2[124] ;
 wire \u_toplayer.reg_layer2[125] ;
 wire \u_toplayer.reg_layer2[126] ;
 wire \u_toplayer.reg_layer2[127] ;
 wire \u_toplayer.reg_layer2[128] ;
 wire \u_toplayer.reg_layer2[129] ;
 wire \u_toplayer.reg_layer2[12] ;
 wire \u_toplayer.reg_layer2[130] ;
 wire \u_toplayer.reg_layer2[131] ;
 wire \u_toplayer.reg_layer2[132] ;
 wire \u_toplayer.reg_layer2[133] ;
 wire \u_toplayer.reg_layer2[134] ;
 wire \u_toplayer.reg_layer2[135] ;
 wire \u_toplayer.reg_layer2[136] ;
 wire \u_toplayer.reg_layer2[137] ;
 wire \u_toplayer.reg_layer2[138] ;
 wire \u_toplayer.reg_layer2[139] ;
 wire \u_toplayer.reg_layer2[13] ;
 wire \u_toplayer.reg_layer2[140] ;
 wire \u_toplayer.reg_layer2[141] ;
 wire \u_toplayer.reg_layer2[142] ;
 wire \u_toplayer.reg_layer2[143] ;
 wire \u_toplayer.reg_layer2[144] ;
 wire \u_toplayer.reg_layer2[145] ;
 wire \u_toplayer.reg_layer2[146] ;
 wire \u_toplayer.reg_layer2[147] ;
 wire \u_toplayer.reg_layer2[148] ;
 wire \u_toplayer.reg_layer2[149] ;
 wire \u_toplayer.reg_layer2[14] ;
 wire \u_toplayer.reg_layer2[150] ;
 wire \u_toplayer.reg_layer2[151] ;
 wire \u_toplayer.reg_layer2[152] ;
 wire \u_toplayer.reg_layer2[153] ;
 wire \u_toplayer.reg_layer2[154] ;
 wire \u_toplayer.reg_layer2[155] ;
 wire \u_toplayer.reg_layer2[156] ;
 wire \u_toplayer.reg_layer2[157] ;
 wire \u_toplayer.reg_layer2[158] ;
 wire \u_toplayer.reg_layer2[159] ;
 wire \u_toplayer.reg_layer2[15] ;
 wire \u_toplayer.reg_layer2[160] ;
 wire \u_toplayer.reg_layer2[161] ;
 wire \u_toplayer.reg_layer2[162] ;
 wire \u_toplayer.reg_layer2[163] ;
 wire \u_toplayer.reg_layer2[164] ;
 wire \u_toplayer.reg_layer2[165] ;
 wire \u_toplayer.reg_layer2[166] ;
 wire \u_toplayer.reg_layer2[167] ;
 wire \u_toplayer.reg_layer2[168] ;
 wire \u_toplayer.reg_layer2[169] ;
 wire \u_toplayer.reg_layer2[16] ;
 wire \u_toplayer.reg_layer2[170] ;
 wire \u_toplayer.reg_layer2[171] ;
 wire \u_toplayer.reg_layer2[172] ;
 wire \u_toplayer.reg_layer2[173] ;
 wire \u_toplayer.reg_layer2[174] ;
 wire \u_toplayer.reg_layer2[175] ;
 wire \u_toplayer.reg_layer2[176] ;
 wire \u_toplayer.reg_layer2[177] ;
 wire \u_toplayer.reg_layer2[178] ;
 wire \u_toplayer.reg_layer2[179] ;
 wire \u_toplayer.reg_layer2[17] ;
 wire \u_toplayer.reg_layer2[180] ;
 wire \u_toplayer.reg_layer2[181] ;
 wire \u_toplayer.reg_layer2[182] ;
 wire \u_toplayer.reg_layer2[183] ;
 wire \u_toplayer.reg_layer2[184] ;
 wire \u_toplayer.reg_layer2[185] ;
 wire \u_toplayer.reg_layer2[186] ;
 wire \u_toplayer.reg_layer2[187] ;
 wire \u_toplayer.reg_layer2[188] ;
 wire \u_toplayer.reg_layer2[189] ;
 wire \u_toplayer.reg_layer2[18] ;
 wire \u_toplayer.reg_layer2[190] ;
 wire \u_toplayer.reg_layer2[191] ;
 wire \u_toplayer.reg_layer2[192] ;
 wire \u_toplayer.reg_layer2[193] ;
 wire \u_toplayer.reg_layer2[194] ;
 wire \u_toplayer.reg_layer2[195] ;
 wire \u_toplayer.reg_layer2[196] ;
 wire \u_toplayer.reg_layer2[197] ;
 wire \u_toplayer.reg_layer2[198] ;
 wire \u_toplayer.reg_layer2[199] ;
 wire \u_toplayer.reg_layer2[19] ;
 wire \u_toplayer.reg_layer2[1] ;
 wire \u_toplayer.reg_layer2[200] ;
 wire \u_toplayer.reg_layer2[201] ;
 wire \u_toplayer.reg_layer2[202] ;
 wire \u_toplayer.reg_layer2[203] ;
 wire \u_toplayer.reg_layer2[204] ;
 wire \u_toplayer.reg_layer2[205] ;
 wire \u_toplayer.reg_layer2[206] ;
 wire \u_toplayer.reg_layer2[207] ;
 wire \u_toplayer.reg_layer2[208] ;
 wire \u_toplayer.reg_layer2[209] ;
 wire \u_toplayer.reg_layer2[20] ;
 wire \u_toplayer.reg_layer2[210] ;
 wire \u_toplayer.reg_layer2[211] ;
 wire \u_toplayer.reg_layer2[212] ;
 wire \u_toplayer.reg_layer2[213] ;
 wire \u_toplayer.reg_layer2[214] ;
 wire \u_toplayer.reg_layer2[215] ;
 wire \u_toplayer.reg_layer2[216] ;
 wire \u_toplayer.reg_layer2[217] ;
 wire \u_toplayer.reg_layer2[218] ;
 wire \u_toplayer.reg_layer2[219] ;
 wire \u_toplayer.reg_layer2[21] ;
 wire \u_toplayer.reg_layer2[220] ;
 wire \u_toplayer.reg_layer2[221] ;
 wire \u_toplayer.reg_layer2[222] ;
 wire \u_toplayer.reg_layer2[223] ;
 wire \u_toplayer.reg_layer2[224] ;
 wire \u_toplayer.reg_layer2[225] ;
 wire \u_toplayer.reg_layer2[226] ;
 wire \u_toplayer.reg_layer2[227] ;
 wire \u_toplayer.reg_layer2[228] ;
 wire \u_toplayer.reg_layer2[229] ;
 wire \u_toplayer.reg_layer2[22] ;
 wire \u_toplayer.reg_layer2[230] ;
 wire \u_toplayer.reg_layer2[231] ;
 wire \u_toplayer.reg_layer2[232] ;
 wire \u_toplayer.reg_layer2[233] ;
 wire \u_toplayer.reg_layer2[234] ;
 wire \u_toplayer.reg_layer2[235] ;
 wire \u_toplayer.reg_layer2[236] ;
 wire \u_toplayer.reg_layer2[237] ;
 wire \u_toplayer.reg_layer2[238] ;
 wire \u_toplayer.reg_layer2[239] ;
 wire \u_toplayer.reg_layer2[23] ;
 wire \u_toplayer.reg_layer2[240] ;
 wire \u_toplayer.reg_layer2[241] ;
 wire \u_toplayer.reg_layer2[242] ;
 wire \u_toplayer.reg_layer2[243] ;
 wire \u_toplayer.reg_layer2[244] ;
 wire \u_toplayer.reg_layer2[245] ;
 wire \u_toplayer.reg_layer2[246] ;
 wire \u_toplayer.reg_layer2[247] ;
 wire \u_toplayer.reg_layer2[248] ;
 wire \u_toplayer.reg_layer2[249] ;
 wire \u_toplayer.reg_layer2[24] ;
 wire \u_toplayer.reg_layer2[250] ;
 wire \u_toplayer.reg_layer2[251] ;
 wire \u_toplayer.reg_layer2[252] ;
 wire \u_toplayer.reg_layer2[253] ;
 wire \u_toplayer.reg_layer2[254] ;
 wire \u_toplayer.reg_layer2[255] ;
 wire \u_toplayer.reg_layer2[25] ;
 wire \u_toplayer.reg_layer2[26] ;
 wire \u_toplayer.reg_layer2[27] ;
 wire \u_toplayer.reg_layer2[28] ;
 wire \u_toplayer.reg_layer2[29] ;
 wire \u_toplayer.reg_layer2[2] ;
 wire \u_toplayer.reg_layer2[30] ;
 wire \u_toplayer.reg_layer2[31] ;
 wire \u_toplayer.reg_layer2[32] ;
 wire \u_toplayer.reg_layer2[33] ;
 wire \u_toplayer.reg_layer2[34] ;
 wire \u_toplayer.reg_layer2[35] ;
 wire \u_toplayer.reg_layer2[36] ;
 wire \u_toplayer.reg_layer2[37] ;
 wire \u_toplayer.reg_layer2[38] ;
 wire \u_toplayer.reg_layer2[39] ;
 wire \u_toplayer.reg_layer2[3] ;
 wire \u_toplayer.reg_layer2[40] ;
 wire \u_toplayer.reg_layer2[41] ;
 wire \u_toplayer.reg_layer2[42] ;
 wire \u_toplayer.reg_layer2[43] ;
 wire \u_toplayer.reg_layer2[44] ;
 wire \u_toplayer.reg_layer2[45] ;
 wire \u_toplayer.reg_layer2[46] ;
 wire \u_toplayer.reg_layer2[47] ;
 wire \u_toplayer.reg_layer2[48] ;
 wire \u_toplayer.reg_layer2[49] ;
 wire \u_toplayer.reg_layer2[4] ;
 wire \u_toplayer.reg_layer2[50] ;
 wire \u_toplayer.reg_layer2[51] ;
 wire \u_toplayer.reg_layer2[52] ;
 wire \u_toplayer.reg_layer2[53] ;
 wire \u_toplayer.reg_layer2[54] ;
 wire \u_toplayer.reg_layer2[55] ;
 wire \u_toplayer.reg_layer2[56] ;
 wire \u_toplayer.reg_layer2[57] ;
 wire \u_toplayer.reg_layer2[58] ;
 wire \u_toplayer.reg_layer2[59] ;
 wire \u_toplayer.reg_layer2[5] ;
 wire \u_toplayer.reg_layer2[60] ;
 wire \u_toplayer.reg_layer2[61] ;
 wire \u_toplayer.reg_layer2[62] ;
 wire \u_toplayer.reg_layer2[63] ;
 wire \u_toplayer.reg_layer2[64] ;
 wire \u_toplayer.reg_layer2[65] ;
 wire \u_toplayer.reg_layer2[66] ;
 wire \u_toplayer.reg_layer2[67] ;
 wire \u_toplayer.reg_layer2[68] ;
 wire \u_toplayer.reg_layer2[69] ;
 wire \u_toplayer.reg_layer2[6] ;
 wire \u_toplayer.reg_layer2[70] ;
 wire \u_toplayer.reg_layer2[71] ;
 wire \u_toplayer.reg_layer2[72] ;
 wire \u_toplayer.reg_layer2[73] ;
 wire \u_toplayer.reg_layer2[74] ;
 wire \u_toplayer.reg_layer2[75] ;
 wire \u_toplayer.reg_layer2[76] ;
 wire \u_toplayer.reg_layer2[77] ;
 wire \u_toplayer.reg_layer2[78] ;
 wire \u_toplayer.reg_layer2[79] ;
 wire \u_toplayer.reg_layer2[7] ;
 wire \u_toplayer.reg_layer2[80] ;
 wire \u_toplayer.reg_layer2[81] ;
 wire \u_toplayer.reg_layer2[82] ;
 wire \u_toplayer.reg_layer2[83] ;
 wire \u_toplayer.reg_layer2[84] ;
 wire \u_toplayer.reg_layer2[85] ;
 wire \u_toplayer.reg_layer2[86] ;
 wire \u_toplayer.reg_layer2[87] ;
 wire \u_toplayer.reg_layer2[88] ;
 wire \u_toplayer.reg_layer2[89] ;
 wire \u_toplayer.reg_layer2[8] ;
 wire \u_toplayer.reg_layer2[90] ;
 wire \u_toplayer.reg_layer2[91] ;
 wire \u_toplayer.reg_layer2[92] ;
 wire \u_toplayer.reg_layer2[93] ;
 wire \u_toplayer.reg_layer2[94] ;
 wire \u_toplayer.reg_layer2[95] ;
 wire \u_toplayer.reg_layer2[96] ;
 wire \u_toplayer.reg_layer2[97] ;
 wire \u_toplayer.reg_layer2[98] ;
 wire \u_toplayer.reg_layer2[99] ;
 wire \u_toplayer.reg_layer2[9] ;
 wire \u_toplayer.u_layer1.neuron_index[0] ;
 wire \u_toplayer.u_layer1.neuron_index[1] ;
 wire \u_toplayer.u_layer1.neuron_index[2] ;
 wire \u_toplayer.u_layer1.neuron_index[3] ;
 wire \u_toplayer.u_layer1.neuron_index[4] ;
 wire \u_toplayer.u_layer1.neuron_index[5] ;
 wire \u_toplayer.u_layer1.statel1[0] ;
 wire \u_toplayer.u_layer1.statel1[1] ;
 wire \u_toplayer.u_layer1.statel1[2] ;
 wire \u_toplayer.u_layer1.statel1[3] ;
 wire \u_toplayer.u_layer1.statel1[4] ;
 wire \u_toplayer.u_layer1.statel1[5] ;
 wire \u_toplayer.u_layer1.statel1[6] ;
 wire \u_toplayer.u_layer1.statel1[7] ;
 wire \u_toplayer.u_layer1.statel1[8] ;
 wire \u_toplayer.u_layer1.sum[0] ;
 wire \u_toplayer.u_layer1.sum[1] ;
 wire \u_toplayer.u_layer1.sum[2] ;
 wire \u_toplayer.u_layer1.sum[3] ;
 wire \u_toplayer.u_layer1.sum[4] ;
 wire \u_toplayer.u_layer1.sum[5] ;
 wire \u_toplayer.u_layer1.sum[6] ;
 wire \u_toplayer.u_layer1.sum[7] ;
 wire \u_toplayer.u_layer1.u_neuron.acc[0] ;
 wire \u_toplayer.u_layer1.u_neuron.acc[10] ;
 wire \u_toplayer.u_layer1.u_neuron.acc[11] ;
 wire \u_toplayer.u_layer1.u_neuron.acc[12] ;
 wire \u_toplayer.u_layer1.u_neuron.acc[13] ;
 wire \u_toplayer.u_layer1.u_neuron.acc[14] ;
 wire \u_toplayer.u_layer1.u_neuron.acc[15] ;
 wire \u_toplayer.u_layer1.u_neuron.acc[16] ;
 wire \u_toplayer.u_layer1.u_neuron.acc[17] ;
 wire \u_toplayer.u_layer1.u_neuron.acc[18] ;
 wire \u_toplayer.u_layer1.u_neuron.acc[19] ;
 wire \u_toplayer.u_layer1.u_neuron.acc[1] ;
 wire \u_toplayer.u_layer1.u_neuron.acc[20] ;
 wire \u_toplayer.u_layer1.u_neuron.acc[21] ;
 wire \u_toplayer.u_layer1.u_neuron.acc[22] ;
 wire \u_toplayer.u_layer1.u_neuron.acc[23] ;
 wire \u_toplayer.u_layer1.u_neuron.acc[2] ;
 wire \u_toplayer.u_layer1.u_neuron.acc[3] ;
 wire \u_toplayer.u_layer1.u_neuron.acc[4] ;
 wire \u_toplayer.u_layer1.u_neuron.acc[5] ;
 wire \u_toplayer.u_layer1.u_neuron.acc[6] ;
 wire \u_toplayer.u_layer1.u_neuron.acc[7] ;
 wire \u_toplayer.u_layer1.u_neuron.acc[8] ;
 wire \u_toplayer.u_layer1.u_neuron.acc[9] ;
 wire \u_toplayer.u_layer1.u_neuron.b[0] ;
 wire \u_toplayer.u_layer1.u_neuron.b[1] ;
 wire \u_toplayer.u_layer1.u_neuron.b[2] ;
 wire \u_toplayer.u_layer1.u_neuron.b[3] ;
 wire \u_toplayer.u_layer1.u_neuron.b[4] ;
 wire \u_toplayer.u_layer1.u_neuron.b[5] ;
 wire \u_toplayer.u_layer1.u_neuron.b[6] ;
 wire \u_toplayer.u_layer1.u_neuron.b[7] ;
 wire \u_toplayer.u_layer1.u_neuron.instCtrl.state[0] ;
 wire \u_toplayer.u_layer1.u_neuron.instCtrl.state[1] ;
 wire \u_toplayer.u_layer1.u_neuron.instCtrl.state[2] ;
 wire \u_toplayer.u_layer1.u_neuron.instCtrl.state[3] ;
 wire \u_toplayer.u_layer1.u_neuron.instCtrl.state[4] ;
 wire \u_toplayer.u_layer1.u_neuron.instCtrl.state[5] ;
 wire \u_toplayer.u_layer1.u_neuron.instCtrl.state[6] ;
 wire \u_toplayer.u_layer1.u_neuron.instCtrl.state[7] ;
 wire \u_toplayer.u_layer1.u_neuron.instCtrl.state[8] ;
 wire \u_toplayer.u_layer1.u_neuron.mult[0] ;
 wire \u_toplayer.u_layer1.u_neuron.mult[10] ;
 wire \u_toplayer.u_layer1.u_neuron.mult[11] ;
 wire \u_toplayer.u_layer1.u_neuron.mult[12] ;
 wire \u_toplayer.u_layer1.u_neuron.mult[13] ;
 wire \u_toplayer.u_layer1.u_neuron.mult[14] ;
 wire \u_toplayer.u_layer1.u_neuron.mult[15] ;
 wire \u_toplayer.u_layer1.u_neuron.mult[1] ;
 wire \u_toplayer.u_layer1.u_neuron.mult[2] ;
 wire \u_toplayer.u_layer1.u_neuron.mult[3] ;
 wire \u_toplayer.u_layer1.u_neuron.mult[4] ;
 wire \u_toplayer.u_layer1.u_neuron.mult[5] ;
 wire \u_toplayer.u_layer1.u_neuron.mult[6] ;
 wire \u_toplayer.u_layer1.u_neuron.mult[7] ;
 wire \u_toplayer.u_layer1.u_neuron.mult[8] ;
 wire \u_toplayer.u_layer1.u_neuron.mult[9] ;
 wire \u_toplayer.u_layer2.neuron_index[0] ;
 wire \u_toplayer.u_layer2.neuron_index[1] ;
 wire \u_toplayer.u_layer2.neuron_index[2] ;
 wire \u_toplayer.u_layer2.neuron_index[3] ;
 wire \u_toplayer.u_layer2.neuron_index[4] ;
 wire \u_toplayer.u_layer2.neuron_index[5] ;
 wire \u_toplayer.u_layer2.statel2[0] ;
 wire \u_toplayer.u_layer2.statel2[1] ;
 wire \u_toplayer.u_layer2.statel2[2] ;
 wire \u_toplayer.u_layer2.statel2[3] ;
 wire \u_toplayer.u_layer2.statel2[4] ;
 wire \u_toplayer.u_layer2.statel2[5] ;
 wire \u_toplayer.u_layer2.statel2[6] ;
 wire \u_toplayer.u_layer2.statel2[7] ;
 wire \u_toplayer.u_layer2.statel2[8] ;
 wire \u_toplayer.u_layer2.sum[0] ;
 wire \u_toplayer.u_layer2.sum[1] ;
 wire \u_toplayer.u_layer2.sum[2] ;
 wire \u_toplayer.u_layer2.sum[3] ;
 wire \u_toplayer.u_layer2.sum[4] ;
 wire \u_toplayer.u_layer2.sum[5] ;
 wire \u_toplayer.u_layer2.sum[6] ;
 wire \u_toplayer.u_layer2.sum[7] ;
 wire \u_toplayer.u_layer2.u_neuron.acc[0] ;
 wire \u_toplayer.u_layer2.u_neuron.acc[10] ;
 wire \u_toplayer.u_layer2.u_neuron.acc[11] ;
 wire \u_toplayer.u_layer2.u_neuron.acc[12] ;
 wire \u_toplayer.u_layer2.u_neuron.acc[13] ;
 wire \u_toplayer.u_layer2.u_neuron.acc[14] ;
 wire \u_toplayer.u_layer2.u_neuron.acc[15] ;
 wire \u_toplayer.u_layer2.u_neuron.acc[16] ;
 wire \u_toplayer.u_layer2.u_neuron.acc[17] ;
 wire \u_toplayer.u_layer2.u_neuron.acc[18] ;
 wire \u_toplayer.u_layer2.u_neuron.acc[19] ;
 wire \u_toplayer.u_layer2.u_neuron.acc[1] ;
 wire \u_toplayer.u_layer2.u_neuron.acc[20] ;
 wire \u_toplayer.u_layer2.u_neuron.acc[21] ;
 wire \u_toplayer.u_layer2.u_neuron.acc[22] ;
 wire \u_toplayer.u_layer2.u_neuron.acc[23] ;
 wire \u_toplayer.u_layer2.u_neuron.acc[2] ;
 wire \u_toplayer.u_layer2.u_neuron.acc[3] ;
 wire \u_toplayer.u_layer2.u_neuron.acc[4] ;
 wire \u_toplayer.u_layer2.u_neuron.acc[5] ;
 wire \u_toplayer.u_layer2.u_neuron.acc[6] ;
 wire \u_toplayer.u_layer2.u_neuron.acc[7] ;
 wire \u_toplayer.u_layer2.u_neuron.acc[8] ;
 wire \u_toplayer.u_layer2.u_neuron.acc[9] ;
 wire \u_toplayer.u_layer2.u_neuron.din[0] ;
 wire \u_toplayer.u_layer2.u_neuron.din[1] ;
 wire \u_toplayer.u_layer2.u_neuron.din[2] ;
 wire \u_toplayer.u_layer2.u_neuron.din[3] ;
 wire \u_toplayer.u_layer2.u_neuron.din[4] ;
 wire \u_toplayer.u_layer2.u_neuron.din[5] ;
 wire \u_toplayer.u_layer2.u_neuron.din[6] ;
 wire \u_toplayer.u_layer2.u_neuron.din[7] ;
 wire \u_toplayer.u_layer2.u_neuron.instCtrl.state[0] ;
 wire \u_toplayer.u_layer2.u_neuron.instCtrl.state[1] ;
 wire \u_toplayer.u_layer2.u_neuron.instCtrl.state[2] ;
 wire \u_toplayer.u_layer2.u_neuron.instCtrl.state[3] ;
 wire \u_toplayer.u_layer2.u_neuron.instCtrl.state[4] ;
 wire \u_toplayer.u_layer2.u_neuron.instCtrl.state[5] ;
 wire \u_toplayer.u_layer2.u_neuron.mult[0] ;
 wire \u_toplayer.u_layer2.u_neuron.mult[10] ;
 wire \u_toplayer.u_layer2.u_neuron.mult[11] ;
 wire \u_toplayer.u_layer2.u_neuron.mult[12] ;
 wire \u_toplayer.u_layer2.u_neuron.mult[13] ;
 wire \u_toplayer.u_layer2.u_neuron.mult[14] ;
 wire \u_toplayer.u_layer2.u_neuron.mult[15] ;
 wire \u_toplayer.u_layer2.u_neuron.mult[1] ;
 wire \u_toplayer.u_layer2.u_neuron.mult[2] ;
 wire \u_toplayer.u_layer2.u_neuron.mult[3] ;
 wire \u_toplayer.u_layer2.u_neuron.mult[4] ;
 wire \u_toplayer.u_layer2.u_neuron.mult[5] ;
 wire \u_toplayer.u_layer2.u_neuron.mult[6] ;
 wire \u_toplayer.u_layer2.u_neuron.mult[7] ;
 wire \u_toplayer.u_layer2.u_neuron.mult[8] ;
 wire \u_toplayer.u_layer2.u_neuron.mult[9] ;
 wire \u_toplayer.u_layer3.neuron_index[0] ;
 wire \u_toplayer.u_layer3.neuron_index[1] ;
 wire \u_toplayer.u_layer3.neuron_index[2] ;
 wire \u_toplayer.u_layer3.neuron_index[3] ;
 wire \u_toplayer.u_layer3.neuron_index[4] ;
 wire \u_toplayer.u_layer3.neuron_index[5] ;
 wire \u_toplayer.u_layer3.stateout[0] ;
 wire \u_toplayer.u_layer3.stateout[1] ;
 wire \u_toplayer.u_layer3.stateout[2] ;
 wire \u_toplayer.u_layer3.stateout[3] ;
 wire \u_toplayer.u_layer3.stateout[4] ;
 wire \u_toplayer.u_layer3.stateout[5] ;
 wire \u_toplayer.u_layer3.stateout[6] ;
 wire \u_toplayer.u_layer3.stateout[7] ;
 wire \u_toplayer.u_layer3.stateout[8] ;
 wire \u_toplayer.u_layer3.sum[0] ;
 wire \u_toplayer.u_layer3.sum[1] ;
 wire \u_toplayer.u_layer3.sum[2] ;
 wire \u_toplayer.u_layer3.sum[3] ;
 wire \u_toplayer.u_layer3.sum[4] ;
 wire \u_toplayer.u_layer3.sum[5] ;
 wire \u_toplayer.u_layer3.sum[6] ;
 wire \u_toplayer.u_layer3.sum[7] ;
 wire \u_toplayer.u_layer3.u_neuron.acc[0] ;
 wire \u_toplayer.u_layer3.u_neuron.acc[10] ;
 wire \u_toplayer.u_layer3.u_neuron.acc[11] ;
 wire \u_toplayer.u_layer3.u_neuron.acc[12] ;
 wire \u_toplayer.u_layer3.u_neuron.acc[13] ;
 wire \u_toplayer.u_layer3.u_neuron.acc[14] ;
 wire \u_toplayer.u_layer3.u_neuron.acc[15] ;
 wire \u_toplayer.u_layer3.u_neuron.acc[16] ;
 wire \u_toplayer.u_layer3.u_neuron.acc[17] ;
 wire \u_toplayer.u_layer3.u_neuron.acc[18] ;
 wire \u_toplayer.u_layer3.u_neuron.acc[19] ;
 wire \u_toplayer.u_layer3.u_neuron.acc[1] ;
 wire \u_toplayer.u_layer3.u_neuron.acc[20] ;
 wire \u_toplayer.u_layer3.u_neuron.acc[21] ;
 wire \u_toplayer.u_layer3.u_neuron.acc[22] ;
 wire \u_toplayer.u_layer3.u_neuron.acc[23] ;
 wire \u_toplayer.u_layer3.u_neuron.acc[2] ;
 wire \u_toplayer.u_layer3.u_neuron.acc[3] ;
 wire \u_toplayer.u_layer3.u_neuron.acc[4] ;
 wire \u_toplayer.u_layer3.u_neuron.acc[5] ;
 wire \u_toplayer.u_layer3.u_neuron.acc[6] ;
 wire \u_toplayer.u_layer3.u_neuron.acc[7] ;
 wire \u_toplayer.u_layer3.u_neuron.acc[8] ;
 wire \u_toplayer.u_layer3.u_neuron.acc[9] ;
 wire \u_toplayer.u_layer3.u_neuron.din[0] ;
 wire \u_toplayer.u_layer3.u_neuron.din[1] ;
 wire \u_toplayer.u_layer3.u_neuron.din[2] ;
 wire \u_toplayer.u_layer3.u_neuron.din[3] ;
 wire \u_toplayer.u_layer3.u_neuron.din[4] ;
 wire \u_toplayer.u_layer3.u_neuron.din[5] ;
 wire \u_toplayer.u_layer3.u_neuron.din[6] ;
 wire \u_toplayer.u_layer3.u_neuron.din[7] ;
 wire \u_toplayer.u_layer3.u_neuron.instCtrl.state[0] ;
 wire \u_toplayer.u_layer3.u_neuron.instCtrl.state[1] ;
 wire \u_toplayer.u_layer3.u_neuron.instCtrl.state[2] ;
 wire \u_toplayer.u_layer3.u_neuron.instCtrl.state[3] ;
 wire \u_toplayer.u_layer3.u_neuron.instCtrl.state[4] ;
 wire \u_toplayer.u_layer3.u_neuron.instCtrl.state[5] ;
 wire \u_toplayer.u_layer3.u_neuron.mult[0] ;
 wire \u_toplayer.u_layer3.u_neuron.mult[10] ;
 wire \u_toplayer.u_layer3.u_neuron.mult[11] ;
 wire \u_toplayer.u_layer3.u_neuron.mult[12] ;
 wire \u_toplayer.u_layer3.u_neuron.mult[13] ;
 wire \u_toplayer.u_layer3.u_neuron.mult[14] ;
 wire \u_toplayer.u_layer3.u_neuron.mult[15] ;
 wire \u_toplayer.u_layer3.u_neuron.mult[1] ;
 wire \u_toplayer.u_layer3.u_neuron.mult[2] ;
 wire \u_toplayer.u_layer3.u_neuron.mult[3] ;
 wire \u_toplayer.u_layer3.u_neuron.mult[4] ;
 wire \u_toplayer.u_layer3.u_neuron.mult[5] ;
 wire \u_toplayer.u_layer3.u_neuron.mult[6] ;
 wire \u_toplayer.u_layer3.u_neuron.mult[7] ;
 wire \u_toplayer.u_layer3.u_neuron.mult[8] ;
 wire \u_toplayer.u_layer3.u_neuron.mult[9] ;
 wire \u_toplayer.u_outlayer.u_neuron.acc[0] ;
 wire \u_toplayer.u_outlayer.u_neuron.acc[10] ;
 wire \u_toplayer.u_outlayer.u_neuron.acc[11] ;
 wire \u_toplayer.u_outlayer.u_neuron.acc[12] ;
 wire \u_toplayer.u_outlayer.u_neuron.acc[13] ;
 wire \u_toplayer.u_outlayer.u_neuron.acc[14] ;
 wire \u_toplayer.u_outlayer.u_neuron.acc[15] ;
 wire \u_toplayer.u_outlayer.u_neuron.acc[16] ;
 wire \u_toplayer.u_outlayer.u_neuron.acc[17] ;
 wire \u_toplayer.u_outlayer.u_neuron.acc[18] ;
 wire \u_toplayer.u_outlayer.u_neuron.acc[19] ;
 wire \u_toplayer.u_outlayer.u_neuron.acc[1] ;
 wire \u_toplayer.u_outlayer.u_neuron.acc[20] ;
 wire \u_toplayer.u_outlayer.u_neuron.acc[21] ;
 wire \u_toplayer.u_outlayer.u_neuron.acc[22] ;
 wire \u_toplayer.u_outlayer.u_neuron.acc[23] ;
 wire \u_toplayer.u_outlayer.u_neuron.acc[2] ;
 wire \u_toplayer.u_outlayer.u_neuron.acc[3] ;
 wire \u_toplayer.u_outlayer.u_neuron.acc[4] ;
 wire \u_toplayer.u_outlayer.u_neuron.acc[5] ;
 wire \u_toplayer.u_outlayer.u_neuron.acc[6] ;
 wire \u_toplayer.u_outlayer.u_neuron.acc[7] ;
 wire \u_toplayer.u_outlayer.u_neuron.acc[8] ;
 wire \u_toplayer.u_outlayer.u_neuron.acc[9] ;
 wire \u_toplayer.u_outlayer.u_neuron.din[0] ;
 wire \u_toplayer.u_outlayer.u_neuron.din[1] ;
 wire \u_toplayer.u_outlayer.u_neuron.din[2] ;
 wire \u_toplayer.u_outlayer.u_neuron.din[3] ;
 wire \u_toplayer.u_outlayer.u_neuron.din[4] ;
 wire \u_toplayer.u_outlayer.u_neuron.din[5] ;
 wire \u_toplayer.u_outlayer.u_neuron.din[6] ;
 wire \u_toplayer.u_outlayer.u_neuron.din[7] ;
 wire \u_toplayer.u_outlayer.u_neuron.instCtrl.state[0] ;
 wire \u_toplayer.u_outlayer.u_neuron.instCtrl.state[1] ;
 wire \u_toplayer.u_outlayer.u_neuron.instCtrl.state[2] ;
 wire \u_toplayer.u_outlayer.u_neuron.instCtrl.state[3] ;
 wire \u_toplayer.u_outlayer.u_neuron.mult[0] ;
 wire \u_toplayer.u_outlayer.u_neuron.mult[10] ;
 wire \u_toplayer.u_outlayer.u_neuron.mult[11] ;
 wire \u_toplayer.u_outlayer.u_neuron.mult[12] ;
 wire \u_toplayer.u_outlayer.u_neuron.mult[13] ;
 wire \u_toplayer.u_outlayer.u_neuron.mult[14] ;
 wire \u_toplayer.u_outlayer.u_neuron.mult[15] ;
 wire \u_toplayer.u_outlayer.u_neuron.mult[1] ;
 wire \u_toplayer.u_outlayer.u_neuron.mult[2] ;
 wire \u_toplayer.u_outlayer.u_neuron.mult[3] ;
 wire \u_toplayer.u_outlayer.u_neuron.mult[4] ;
 wire \u_toplayer.u_outlayer.u_neuron.mult[5] ;
 wire \u_toplayer.u_outlayer.u_neuron.mult[6] ;
 wire \u_toplayer.u_outlayer.u_neuron.mult[7] ;
 wire \u_toplayer.u_outlayer.u_neuron.mult[8] ;
 wire \u_toplayer.u_outlayer.u_neuron.mult[9] ;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net2692;
 wire net2693;
 wire net2694;
 wire net2695;
 wire net2696;
 wire net2697;
 wire net2698;
 wire net2699;
 wire net2700;
 wire net2701;
 wire net2702;
 wire net2703;
 wire net2704;
 wire net2705;
 wire net2706;
 wire net2707;
 wire net2708;
 wire net2709;
 wire net2710;
 wire net2711;
 wire net2712;
 wire net2713;
 wire net2714;
 wire net2715;
 wire net2716;
 wire net2717;
 wire net2718;
 wire net2719;
 wire net2720;
 wire net2721;
 wire net2722;
 wire net2723;
 wire net2724;
 wire net2725;
 wire net2726;
 wire net2727;
 wire net2728;
 wire net2729;
 wire net2730;
 wire net2731;
 wire net2732;
 wire net2733;
 wire net2734;
 wire net2735;
 wire net2736;
 wire net2737;
 wire net2738;
 wire net2739;
 wire net2740;
 wire net2741;
 wire net2742;
 wire net2743;
 wire net2744;
 wire net2745;
 wire net2746;
 wire net2747;
 wire net2748;
 wire net2749;
 wire net2750;
 wire net2751;
 wire net2752;
 wire net2753;
 wire net2754;
 wire net2755;
 wire net2756;
 wire net2757;
 wire net2758;
 wire net2759;
 wire net2760;
 wire net2761;
 wire net2762;
 wire net2763;
 wire net2764;
 wire net2765;
 wire net2766;
 wire net2767;
 wire net2768;
 wire net2769;
 wire net2770;
 wire net2771;
 wire net2772;
 wire net2773;
 wire net2774;
 wire net2775;
 wire net2776;
 wire net2777;
 wire net2778;
 wire net2779;
 wire net2780;
 wire net2781;
 wire net2782;
 wire net2783;
 wire net2784;
 wire net2785;
 wire net2786;
 wire net2787;
 wire net2788;
 wire net2789;
 wire net2790;
 wire net2791;
 wire net2792;
 wire net2793;
 wire net2794;
 wire net2795;
 wire net2796;
 wire net2797;
 wire net2798;
 wire net2799;
 wire net2800;
 wire net2801;
 wire net2802;
 wire net2803;
 wire net2804;
 wire net2805;
 wire net2806;
 wire net2807;
 wire net2808;
 wire net2809;
 wire net2810;
 wire net2811;
 wire net2812;
 wire net2813;
 wire net2814;
 wire net2815;
 wire net2816;
 wire net2817;
 wire net2818;
 wire net2819;
 wire net2820;
 wire net2821;
 wire net2822;
 wire net2823;
 wire net2824;
 wire net2825;
 wire net2826;
 wire net2827;
 wire net2828;
 wire net2829;
 wire net2830;
 wire net2831;
 wire net2832;
 wire net2833;
 wire net2834;
 wire net2835;
 wire net2836;
 wire net2837;
 wire net2838;
 wire net2839;
 wire net2840;
 wire net2841;
 wire net2842;
 wire net2843;
 wire net2844;
 wire net2845;
 wire net2846;
 wire net2847;
 wire net2848;
 wire net2849;
 wire net2850;
 wire net2851;
 wire net2852;
 wire net2853;
 wire net2854;
 wire net2855;
 wire net2856;
 wire net2857;
 wire net2858;
 wire net2859;
 wire net2860;
 wire net2861;
 wire net2862;
 wire net2863;
 wire net2864;
 wire net2865;
 wire net2866;
 wire net2867;
 wire net2868;
 wire net2869;
 wire net2870;
 wire net2871;
 wire net2872;
 wire net2873;
 wire net2874;
 wire net2875;
 wire net2876;
 wire net2877;
 wire net2878;
 wire net2879;
 wire net2880;
 wire net2881;
 wire net2882;
 wire net2883;
 wire net2884;
 wire net2885;
 wire net2886;
 wire net2887;
 wire net2888;
 wire net2889;
 wire net2890;
 wire net2891;
 wire net2892;
 wire net2893;
 wire net2894;
 wire net2895;
 wire net2896;
 wire net2897;
 wire net2898;
 wire net2899;
 wire net2900;
 wire net2901;
 wire net2902;
 wire net2903;
 wire net2904;
 wire net2905;
 wire net2906;
 wire net2907;
 wire net2908;
 wire net2909;
 wire net2910;
 wire net2911;
 wire net2912;
 wire net2913;
 wire net2914;
 wire net2915;
 wire net2916;
 wire net2917;
 wire net2918;
 wire net2919;
 wire net2920;
 wire net2921;
 wire net2922;
 wire net2923;
 wire net2924;
 wire net2925;
 wire net2926;
 wire net2927;
 wire net2928;
 wire net2929;
 wire net2930;
 wire net2931;
 wire net2932;
 wire net2933;
 wire net2934;
 wire net2935;
 wire net2936;
 wire net2937;
 wire net2938;
 wire net2939;
 wire net2940;
 wire net2941;
 wire net2942;
 wire net2943;
 wire net2944;
 wire net2945;
 wire net2946;
 wire net2947;
 wire net2948;
 wire net2949;
 wire net2950;
 wire net2951;
 wire net2952;
 wire net2953;
 wire net2954;
 wire net2955;
 wire net2956;
 wire net2957;
 wire net2958;
 wire net2959;
 wire net2960;
 wire net2961;
 wire net2962;
 wire net2963;
 wire net2964;
 wire net2965;
 wire net2966;
 wire net2967;
 wire net2968;
 wire net2969;
 wire net2970;
 wire net2971;
 wire net2972;
 wire net2973;
 wire net2974;
 wire net2975;
 wire net2976;
 wire net2977;
 wire net2978;
 wire net2979;
 wire net2980;
 wire net2981;
 wire net2982;
 wire net2983;
 wire net2984;
 wire net2985;
 wire net2986;
 wire net2987;
 wire net2988;
 wire net2989;
 wire net2990;
 wire net2991;
 wire net2992;
 wire net2993;
 wire net2994;
 wire net2995;
 wire net2996;
 wire net2997;
 wire net2998;
 wire net2999;
 wire net3000;
 wire net3001;
 wire net3002;
 wire net3003;
 wire net3004;
 wire net3005;
 wire net3006;
 wire net3007;
 wire net3008;
 wire net3009;
 wire net3010;
 wire net3011;
 wire net3012;
 wire net3013;
 wire net3014;
 wire net3015;
 wire net3016;
 wire net3017;
 wire net3018;
 wire net3019;
 wire net3020;
 wire net3021;
 wire net3022;
 wire net3023;
 wire net3024;
 wire net3025;
 wire net3026;
 wire net3027;
 wire net3028;
 wire net3029;
 wire net3030;
 wire net3031;
 wire net3032;
 wire net3033;
 wire net3034;
 wire net3035;
 wire net3036;
 wire net3037;
 wire net3038;
 wire net3039;
 wire net3040;
 wire net3041;
 wire net3042;
 wire net3043;
 wire net3044;
 wire net3045;
 wire net3046;
 wire net3047;
 wire net3048;
 wire net3049;
 wire net3050;
 wire net3051;
 wire net3052;
 wire net3053;
 wire net3054;
 wire net3055;
 wire net3056;
 wire net3057;
 wire net3058;
 wire net3059;
 wire net3060;
 wire net3061;
 wire net3062;
 wire net3063;
 wire net3064;
 wire net3065;
 wire net3066;
 wire net3067;
 wire net3068;
 wire net3069;
 wire net3070;
 wire net3071;
 wire net3072;
 wire net3073;
 wire net3074;
 wire net3075;
 wire net3076;
 wire net3077;
 wire net3078;
 wire net3079;
 wire net3080;
 wire net3081;
 wire net3082;
 wire net3083;
 wire net3084;
 wire net3085;
 wire net3086;
 wire net3087;
 wire net3088;
 wire net3089;
 wire net3090;
 wire net3091;
 wire net3092;
 wire net3093;
 wire net3094;
 wire net3095;
 wire net3096;
 wire net3097;
 wire net3098;
 wire net3099;
 wire net3100;
 wire net3101;
 wire net3102;
 wire net3103;
 wire net3104;
 wire net3105;
 wire net3106;
 wire net3107;
 wire net3108;
 wire net3109;
 wire net3110;
 wire net3111;
 wire net3112;
 wire net3113;
 wire net3114;
 wire net3115;
 wire net3116;
 wire net3117;
 wire net3118;
 wire net3119;
 wire net3120;
 wire net3121;
 wire net3122;
 wire net3123;
 wire net3124;
 wire net3125;
 wire net3126;
 wire net3127;
 wire net3128;
 wire net3129;
 wire net3130;
 wire net3131;
 wire net3132;
 wire net3133;
 wire net3134;
 wire net3135;
 wire net3136;
 wire net3137;
 wire net3138;
 wire net3139;
 wire net3140;
 wire net3141;
 wire net3142;
 wire net3143;
 wire net3144;
 wire net3145;
 wire net3146;
 wire net3147;
 wire net3148;
 wire net3149;
 wire net3150;
 wire net3151;
 wire net3152;
 wire net3153;
 wire net3154;
 wire net3155;
 wire net3156;
 wire net3157;
 wire net3158;
 wire net3159;
 wire net3160;
 wire net3161;
 wire net3162;
 wire net3163;
 wire net3164;
 wire net3165;
 wire net3166;
 wire net3167;
 wire net3168;
 wire net3169;
 wire net3170;
 wire net3171;
 wire net3172;
 wire net3173;
 wire net3174;
 wire net3175;
 wire net3176;
 wire net3177;
 wire net3178;
 wire net3179;
 wire net3180;
 wire net3181;
 wire net3182;
 wire net3183;
 wire net3184;
 wire net3185;
 wire net3186;
 wire net3187;
 wire net3188;
 wire net3189;
 wire net3190;
 wire net3191;
 wire net3192;
 wire net3193;
 wire net3194;
 wire net3195;
 wire net3196;
 wire net3197;
 wire net3198;
 wire net3199;
 wire net3200;
 wire net3201;
 wire net3202;
 wire net3203;
 wire net3204;
 wire net3205;
 wire net3206;
 wire net3207;
 wire net3208;
 wire net3209;
 wire net3210;
 wire net3211;
 wire net3212;
 wire net3213;
 wire net3214;
 wire net3215;
 wire net3216;
 wire net3217;
 wire net3218;
 wire net3219;
 wire net3220;
 wire net3221;
 wire net3222;
 wire net3223;
 wire net3224;
 wire net3225;
 wire net3226;
 wire net3227;
 wire net3228;
 wire net3229;
 wire net3230;
 wire net3231;
 wire net3232;
 wire net3233;
 wire net3234;
 wire net3235;
 wire net3236;
 wire net3237;
 wire net3238;
 wire net3239;
 wire net3240;
 wire net3241;
 wire net3242;
 wire net3243;
 wire net3244;
 wire net3245;
 wire net3246;
 wire net3247;
 wire net3248;
 wire net3249;
 wire net3250;
 wire net3251;
 wire net3252;
 wire net3253;
 wire net3254;
 wire net3255;
 wire net3256;
 wire net3257;
 wire net3258;
 wire net3259;
 wire net3260;
 wire net3261;
 wire net3262;
 wire net3263;
 wire net3264;
 wire net3265;
 wire net3266;
 wire net3267;
 wire net3268;
 wire net3269;
 wire net3270;
 wire net3271;
 wire net3272;
 wire net3273;
 wire net3274;
 wire net3275;
 wire net3276;
 wire net3277;
 wire net3278;
 wire net3279;
 wire net3280;
 wire net3281;
 wire net3282;
 wire net3283;
 wire net3284;
 wire net3285;
 wire net3286;
 wire net3287;
 wire net3288;
 wire net3289;
 wire net3290;
 wire net3291;
 wire net3292;
 wire net3293;
 wire net3294;
 wire net3295;
 wire net3296;
 wire net3297;
 wire net3298;
 wire net3299;
 wire net3300;
 wire net3301;
 wire net3302;
 wire net3303;
 wire net3304;
 wire net3305;
 wire net3306;
 wire net3307;
 wire net3308;
 wire net3309;
 wire net3310;
 wire net3311;
 wire net3312;
 wire net3313;
 wire net3314;
 wire net3315;
 wire net3316;
 wire net3317;
 wire net3318;
 wire net3319;
 wire net3320;
 wire net3321;
 wire net3322;
 wire net3323;
 wire net3324;
 wire net3325;
 wire net3326;
 wire net3327;
 wire net3328;
 wire net3329;
 wire net3330;
 wire net3331;
 wire net3332;
 wire net3333;
 wire net3334;
 wire net3335;
 wire net3336;
 wire net3337;
 wire net3338;
 wire net3339;
 wire net3340;
 wire net3341;
 wire net3342;
 wire net3343;
 wire net3344;
 wire net3345;
 wire net3346;
 wire net3347;
 wire net3348;
 wire net3349;
 wire net3350;
 wire net3351;
 wire net3352;
 wire net3353;
 wire net3354;
 wire net3355;
 wire net3356;
 wire net3357;
 wire net3358;
 wire net3359;
 wire net3360;
 wire net3361;
 wire net3362;
 wire net3363;
 wire net3364;
 wire net3365;
 wire net3366;
 wire net3367;
 wire net3368;
 wire net3369;
 wire net3370;
 wire net3371;
 wire net3372;
 wire net3373;
 wire net3374;
 wire net3375;
 wire net3376;
 wire net3377;
 wire net3378;
 wire net3379;
 wire net3380;
 wire net3381;
 wire net3382;
 wire net3383;
 wire net3384;
 wire net3385;
 wire net3386;
 wire net3387;
 wire net3388;
 wire net3389;
 wire net3390;
 wire net3391;
 wire net3392;
 wire net3393;
 wire net3394;
 wire net3395;
 wire net3396;
 wire net3397;
 wire net3398;
 wire net3399;
 wire net3400;
 wire net3401;
 wire net3402;
 wire net3403;
 wire net3404;
 wire net3405;
 wire net3406;
 wire net3407;
 wire net3408;
 wire net3409;
 wire net3410;
 wire net3411;
 wire net3412;
 wire net3413;
 wire net3414;
 wire net3415;
 wire net3416;
 wire net3417;
 wire net3418;
 wire net3419;
 wire net3420;
 wire net3421;
 wire net3422;
 wire net3423;
 wire net3424;
 wire net3425;
 wire net3426;
 wire net3427;
 wire net3428;
 wire net3429;
 wire net3430;
 wire net3431;
 wire net3432;
 wire net3433;
 wire net3434;
 wire net3435;
 wire net3436;
 wire net3437;
 wire net3438;
 wire net3439;
 wire net3440;
 wire net3441;
 wire net3442;
 wire net3443;
 wire net3444;
 wire net3445;
 wire net3446;
 wire net3447;
 wire net3448;
 wire net3449;
 wire net3450;
 wire net3451;
 wire net3452;
 wire net3453;
 wire net3454;
 wire net3455;
 wire net3456;
 wire net3457;
 wire net3458;
 wire net3459;
 wire net3460;
 wire net3461;
 wire net3462;
 wire net3463;
 wire net3464;
 wire net3465;
 wire net3466;
 wire net3467;
 wire net3468;
 wire net3469;
 wire net3470;
 wire net3471;
 wire net3472;
 wire net3473;
 wire net3474;
 wire net3475;
 wire net3476;
 wire net3477;
 wire net3478;
 wire net3479;
 wire net3480;
 wire net3481;
 wire net3482;
 wire net3483;
 wire net3484;
 wire net3485;
 wire net3486;
 wire net3487;
 wire net3488;
 wire net3489;
 wire net3490;
 wire net3491;
 wire net3492;
 wire net3493;
 wire net3494;
 wire net3495;
 wire net3496;
 wire net3497;
 wire net3498;
 wire net3499;
 wire net3500;
 wire net3501;
 wire net3502;
 wire net3503;
 wire net3504;
 wire net3505;
 wire net3506;
 wire net3507;
 wire net3508;
 wire net3509;
 wire net3510;
 wire net3511;
 wire net3512;
 wire net3513;
 wire net3514;
 wire net3515;
 wire net3516;
 wire net3517;
 wire net3518;
 wire net3519;
 wire net3520;
 wire net3521;
 wire net3522;
 wire net3523;
 wire net3524;
 wire net3525;
 wire net3526;
 wire net3527;
 wire net3528;
 wire net3529;
 wire net3530;
 wire net3531;
 wire net3532;
 wire net3533;
 wire net3534;
 wire net3535;
 wire net3536;
 wire net3537;
 wire net3538;
 wire net3539;
 wire net3540;
 wire net3541;
 wire net3542;
 wire net3543;
 wire net3544;
 wire net3545;
 wire net3546;
 wire net3547;
 wire net3548;
 wire net3549;
 wire net3550;
 wire net3551;
 wire net3552;
 wire net3553;
 wire net3554;
 wire net3555;
 wire net3556;
 wire net3557;
 wire net3558;
 wire net3559;
 wire net3560;
 wire net3561;
 wire net3562;
 wire net3563;
 wire net3564;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_leaf_0_clk_regs;
 wire clknet_leaf_1_clk_regs;
 wire clknet_leaf_2_clk_regs;
 wire clknet_leaf_3_clk_regs;
 wire clknet_leaf_4_clk_regs;
 wire clknet_leaf_5_clk_regs;
 wire clknet_leaf_6_clk_regs;
 wire clknet_leaf_7_clk_regs;
 wire clknet_leaf_8_clk_regs;
 wire clknet_leaf_9_clk_regs;
 wire clknet_leaf_10_clk_regs;
 wire clknet_leaf_11_clk_regs;
 wire clknet_leaf_12_clk_regs;
 wire clknet_leaf_13_clk_regs;
 wire clknet_leaf_14_clk_regs;
 wire clknet_leaf_15_clk_regs;
 wire clknet_leaf_16_clk_regs;
 wire clknet_leaf_17_clk_regs;
 wire clknet_leaf_18_clk_regs;
 wire clknet_leaf_19_clk_regs;
 wire clknet_leaf_20_clk_regs;
 wire clknet_leaf_21_clk_regs;
 wire clknet_leaf_22_clk_regs;
 wire clknet_leaf_23_clk_regs;
 wire clknet_leaf_24_clk_regs;
 wire clknet_leaf_25_clk_regs;
 wire clknet_leaf_26_clk_regs;
 wire clknet_leaf_27_clk_regs;
 wire clknet_leaf_28_clk_regs;
 wire clknet_leaf_29_clk_regs;
 wire clknet_leaf_30_clk_regs;
 wire clknet_leaf_31_clk_regs;
 wire clknet_leaf_32_clk_regs;
 wire clknet_leaf_33_clk_regs;
 wire clknet_leaf_34_clk_regs;
 wire clknet_leaf_35_clk_regs;
 wire clknet_leaf_36_clk_regs;
 wire clknet_leaf_37_clk_regs;
 wire clknet_leaf_38_clk_regs;
 wire clknet_leaf_39_clk_regs;
 wire clknet_leaf_40_clk_regs;
 wire clknet_leaf_41_clk_regs;
 wire clknet_leaf_42_clk_regs;
 wire clknet_leaf_43_clk_regs;
 wire clknet_leaf_44_clk_regs;
 wire clknet_leaf_45_clk_regs;
 wire clknet_leaf_46_clk_regs;
 wire clknet_leaf_47_clk_regs;
 wire clknet_leaf_48_clk_regs;
 wire clknet_leaf_49_clk_regs;
 wire clknet_leaf_50_clk_regs;
 wire clknet_leaf_51_clk_regs;
 wire clknet_leaf_52_clk_regs;
 wire clknet_leaf_53_clk_regs;
 wire clknet_leaf_54_clk_regs;
 wire clknet_leaf_55_clk_regs;
 wire clknet_leaf_56_clk_regs;
 wire clknet_leaf_57_clk_regs;
 wire clknet_leaf_58_clk_regs;
 wire clknet_leaf_59_clk_regs;
 wire clknet_leaf_60_clk_regs;
 wire clknet_leaf_61_clk_regs;
 wire clknet_leaf_62_clk_regs;
 wire clknet_leaf_63_clk_regs;
 wire clknet_leaf_64_clk_regs;
 wire clknet_leaf_65_clk_regs;
 wire clknet_leaf_66_clk_regs;
 wire clknet_leaf_67_clk_regs;
 wire clknet_leaf_68_clk_regs;
 wire clknet_leaf_69_clk_regs;
 wire clknet_leaf_70_clk_regs;
 wire clknet_leaf_71_clk_regs;
 wire clknet_leaf_72_clk_regs;
 wire clknet_leaf_73_clk_regs;
 wire clknet_leaf_74_clk_regs;
 wire clknet_leaf_75_clk_regs;
 wire clknet_leaf_76_clk_regs;
 wire clknet_leaf_77_clk_regs;
 wire clknet_leaf_78_clk_regs;
 wire clknet_leaf_79_clk_regs;
 wire clknet_leaf_80_clk_regs;
 wire clknet_leaf_81_clk_regs;
 wire clknet_leaf_82_clk_regs;
 wire clknet_leaf_83_clk_regs;
 wire clknet_leaf_84_clk_regs;
 wire clknet_leaf_85_clk_regs;
 wire clknet_leaf_86_clk_regs;
 wire clknet_leaf_87_clk_regs;
 wire clknet_leaf_88_clk_regs;
 wire clknet_leaf_90_clk_regs;
 wire clknet_leaf_91_clk_regs;
 wire clknet_leaf_92_clk_regs;
 wire clknet_leaf_93_clk_regs;
 wire clknet_leaf_94_clk_regs;
 wire clknet_leaf_95_clk_regs;
 wire clknet_leaf_96_clk_regs;
 wire clknet_leaf_97_clk_regs;
 wire clknet_leaf_98_clk_regs;
 wire clknet_leaf_99_clk_regs;
 wire clknet_leaf_100_clk_regs;
 wire clknet_leaf_101_clk_regs;
 wire clknet_leaf_102_clk_regs;
 wire clknet_leaf_103_clk_regs;
 wire clknet_leaf_104_clk_regs;
 wire clknet_leaf_105_clk_regs;
 wire clknet_leaf_106_clk_regs;
 wire clknet_leaf_107_clk_regs;
 wire clknet_leaf_108_clk_regs;
 wire clknet_leaf_109_clk_regs;
 wire clknet_leaf_110_clk_regs;
 wire clknet_leaf_111_clk_regs;
 wire clknet_0_clk_regs;
 wire clknet_4_0_0_clk_regs;
 wire clknet_4_1_0_clk_regs;
 wire clknet_4_2_0_clk_regs;
 wire clknet_4_3_0_clk_regs;
 wire clknet_4_4_0_clk_regs;
 wire clknet_4_5_0_clk_regs;
 wire clknet_4_6_0_clk_regs;
 wire clknet_4_7_0_clk_regs;
 wire clknet_4_8_0_clk_regs;
 wire clknet_4_9_0_clk_regs;
 wire clknet_4_10_0_clk_regs;
 wire clknet_4_11_0_clk_regs;
 wire clknet_4_12_0_clk_regs;
 wire clknet_4_13_0_clk_regs;
 wire clknet_4_14_0_clk_regs;
 wire clknet_4_15_0_clk_regs;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net1210;
 wire net1211;
 wire net1212;

 sg13g2_inv_1 _06888_ (.Y(_01018_),
    .A(\u_toplayer.u_layer3.stateout[8] ));
 sg13g2_inv_1 _06889_ (.Y(_01019_),
    .A(net895));
 sg13g2_inv_1 _06890_ (.Y(_01020_),
    .A(net892));
 sg13g2_inv_1 _06891_ (.Y(_01021_),
    .A(net831));
 sg13g2_inv_1 _06892_ (.Y(_01022_),
    .A(\u_toplayer.delay_counter_layer1[1] ));
 sg13g2_inv_1 _06893_ (.Y(_01023_),
    .A(\u_toplayer.delay_counter_layer2[1] ));
 sg13g2_inv_1 _06894_ (.Y(_01024_),
    .A(net980));
 sg13g2_inv_1 _06895_ (.Y(_01025_),
    .A(\u_toplayer.delay_counter_layer3[1] ));
 sg13g2_inv_1 _06896_ (.Y(_01026_),
    .A(\u_toplayer.u_layer1.statel1[8] ));
 sg13g2_inv_1 _06897_ (.Y(_01027_),
    .A(net1015));
 sg13g2_inv_1 _06898_ (.Y(_01028_),
    .A(net972));
 sg13g2_inv_1 _06899_ (.Y(_01029_),
    .A(net3230));
 sg13g2_inv_1 _06900_ (.Y(_01030_),
    .A(\u_toplayer.u_layer1.u_neuron.instCtrl.state[1] ));
 sg13g2_inv_2 _06901_ (.Y(_01031_),
    .A(\u_toplayer.delayed_done_layer1 ));
 sg13g2_inv_1 _06902_ (.Y(_01032_),
    .A(net1149));
 sg13g2_inv_2 _06903_ (.Y(_01033_),
    .A(net3149));
 sg13g2_inv_1 _06904_ (.Y(_01034_),
    .A(net937));
 sg13g2_inv_1 _06905_ (.Y(_01035_),
    .A(net3242));
 sg13g2_inv_1 _06906_ (.Y(_01036_),
    .A(net3102));
 sg13g2_inv_1 _06907_ (.Y(_01037_),
    .A(net1161));
 sg13g2_inv_1 _06908_ (.Y(_01038_),
    .A(net1118));
 sg13g2_inv_1 _06909_ (.Y(_01039_),
    .A(net1170));
 sg13g2_inv_1 _06910_ (.Y(_01040_),
    .A(net1155));
 sg13g2_inv_1 _06911_ (.Y(_01041_),
    .A(net1158));
 sg13g2_inv_1 _06912_ (.Y(_01042_),
    .A(net1083));
 sg13g2_inv_1 _06913_ (.Y(_01043_),
    .A(net1110));
 sg13g2_inv_1 _06914_ (.Y(_01044_),
    .A(net1051));
 sg13g2_inv_1 _06915_ (.Y(_01045_),
    .A(net3195));
 sg13g2_inv_4 _06916_ (.A(net3390),
    .Y(_01046_));
 sg13g2_inv_1 _06917_ (.Y(_01047_),
    .A(net3359));
 sg13g2_inv_1 _06918_ (.Y(_01048_),
    .A(\u_toplayer.u_outlayer.u_neuron.mult[12] ));
 sg13g2_inv_2 _06919_ (.Y(_01049_),
    .A(net3285));
 sg13g2_inv_1 _06920_ (.Y(_01050_),
    .A(net1206));
 sg13g2_inv_1 _06921_ (.Y(_01051_),
    .A(net1130));
 sg13g2_inv_1 _06922_ (.Y(_01052_),
    .A(net1122));
 sg13g2_inv_1 _06923_ (.Y(_01053_),
    .A(net1111));
 sg13g2_inv_1 _06924_ (.Y(_01054_),
    .A(net3157));
 sg13g2_inv_1 _06925_ (.Y(_01055_),
    .A(net1088));
 sg13g2_inv_1 _06926_ (.Y(_01056_),
    .A(net1095));
 sg13g2_inv_1 _06927_ (.Y(_01057_),
    .A(net1144));
 sg13g2_inv_1 _06928_ (.Y(_01058_),
    .A(net1151));
 sg13g2_inv_1 _06929_ (.Y(_01059_),
    .A(net924));
 sg13g2_inv_1 _06930_ (.Y(_01060_),
    .A(net1109));
 sg13g2_inv_1 _06931_ (.Y(_01061_),
    .A(net1032));
 sg13g2_inv_1 _06932_ (.Y(_01062_),
    .A(net1121));
 sg13g2_inv_1 _06933_ (.Y(_01063_),
    .A(net898));
 sg13g2_inv_1 _06934_ (.Y(_01064_),
    .A(net3155));
 sg13g2_inv_1 _06935_ (.Y(_01065_),
    .A(net681));
 sg13g2_inv_1 _06936_ (.Y(_01066_),
    .A(\u_toplayer.reg_layer2[72] ));
 sg13g2_inv_1 _06937_ (.Y(_01067_),
    .A(\u_toplayer.reg_layer2[104] ));
 sg13g2_inv_1 _06938_ (.Y(_01068_),
    .A(\u_toplayer.reg_layer2[200] ));
 sg13g2_inv_1 _06939_ (.Y(_01069_),
    .A(\u_toplayer.reg_layer2[232] ));
 sg13g2_inv_1 _06940_ (.Y(_01070_),
    .A(\u_toplayer.reg_layer2[73] ));
 sg13g2_inv_1 _06941_ (.Y(_01071_),
    .A(\u_toplayer.reg_layer2[105] ));
 sg13g2_inv_1 _06942_ (.Y(_01072_),
    .A(\u_toplayer.reg_layer2[201] ));
 sg13g2_inv_1 _06943_ (.Y(_01073_),
    .A(\u_toplayer.reg_layer2[233] ));
 sg13g2_inv_1 _06944_ (.Y(_01074_),
    .A(\u_toplayer.reg_layer2[74] ));
 sg13g2_inv_1 _06945_ (.Y(_01075_),
    .A(\u_toplayer.reg_layer2[106] ));
 sg13g2_inv_1 _06946_ (.Y(_01076_),
    .A(\u_toplayer.reg_layer2[202] ));
 sg13g2_inv_1 _06947_ (.Y(_01077_),
    .A(\u_toplayer.reg_layer2[234] ));
 sg13g2_inv_1 _06948_ (.Y(_01078_),
    .A(\u_toplayer.reg_layer2[75] ));
 sg13g2_inv_1 _06949_ (.Y(_01079_),
    .A(\u_toplayer.reg_layer2[107] ));
 sg13g2_inv_1 _06950_ (.Y(_01080_),
    .A(\u_toplayer.reg_layer2[203] ));
 sg13g2_inv_1 _06951_ (.Y(_01081_),
    .A(\u_toplayer.reg_layer2[235] ));
 sg13g2_inv_1 _06952_ (.Y(_01082_),
    .A(\u_toplayer.reg_layer2[76] ));
 sg13g2_inv_1 _06953_ (.Y(_01083_),
    .A(\u_toplayer.reg_layer2[108] ));
 sg13g2_inv_1 _06954_ (.Y(_01084_),
    .A(\u_toplayer.reg_layer2[204] ));
 sg13g2_inv_1 _06955_ (.Y(_01085_),
    .A(\u_toplayer.reg_layer2[77] ));
 sg13g2_inv_1 _06956_ (.Y(_01086_),
    .A(\u_toplayer.reg_layer2[109] ));
 sg13g2_inv_1 _06957_ (.Y(_01087_),
    .A(\u_toplayer.reg_layer2[205] ));
 sg13g2_inv_1 _06958_ (.Y(_01088_),
    .A(\u_toplayer.reg_layer2[237] ));
 sg13g2_inv_1 _06959_ (.Y(_01089_),
    .A(\u_toplayer.reg_layer2[78] ));
 sg13g2_inv_1 _06960_ (.Y(_01090_),
    .A(\u_toplayer.reg_layer2[110] ));
 sg13g2_inv_1 _06961_ (.Y(_01091_),
    .A(\u_toplayer.reg_layer2[206] ));
 sg13g2_inv_1 _06962_ (.Y(_01092_),
    .A(\u_toplayer.reg_layer2[79] ));
 sg13g2_inv_1 _06963_ (.Y(_01093_),
    .A(\u_toplayer.reg_layer2[111] ));
 sg13g2_inv_1 _06964_ (.Y(_01094_),
    .A(\u_toplayer.reg_layer2[207] ));
 sg13g2_inv_1 _06965_ (.Y(_01095_),
    .A(net3172));
 sg13g2_inv_1 _06966_ (.Y(_01096_),
    .A(net3169));
 sg13g2_inv_1 _06967_ (.Y(_01097_),
    .A(net1136));
 sg13g2_inv_1 _06968_ (.Y(_01098_),
    .A(net1055));
 sg13g2_inv_1 _06969_ (.Y(_01099_),
    .A(net821));
 sg13g2_inv_1 _06970_ (.Y(_01100_),
    .A(net1137));
 sg13g2_inv_1 _06971_ (.Y(_01101_),
    .A(net1157));
 sg13g2_inv_1 _06972_ (.Y(_01102_),
    .A(net785));
 sg13g2_inv_1 _06973_ (.Y(_01103_),
    .A(net1037));
 sg13g2_inv_1 _06974_ (.Y(_01104_),
    .A(net1173));
 sg13g2_inv_1 _06975_ (.Y(_01105_),
    .A(net3060));
 sg13g2_inv_1 _06976_ (.Y(_01106_),
    .A(net1114));
 sg13g2_inv_1 _06977_ (.Y(_01107_),
    .A(net3062));
 sg13g2_inv_1 _06978_ (.Y(_01108_),
    .A(net1070));
 sg13g2_inv_1 _06979_ (.Y(_01109_),
    .A(net1132));
 sg13g2_inv_1 _06980_ (.Y(_01110_),
    .A(net1119));
 sg13g2_inv_1 _06981_ (.Y(_01111_),
    .A(net1050));
 sg13g2_inv_1 _06982_ (.Y(_01112_),
    .A(net1124));
 sg13g2_inv_1 _06983_ (.Y(_01113_),
    .A(net1081));
 sg13g2_inv_1 _06984_ (.Y(_01114_),
    .A(net1168));
 sg13g2_inv_1 _06985_ (.Y(_01115_),
    .A(net1104));
 sg13g2_inv_1 _06986_ (.Y(_01116_),
    .A(net3059));
 sg13g2_inv_1 _06987_ (.Y(_01117_),
    .A(net871));
 sg13g2_inv_1 _06988_ (.Y(_01118_),
    .A(\u_toplayer.reg_layer1[72] ));
 sg13g2_inv_1 _06989_ (.Y(_01119_),
    .A(\u_toplayer.reg_layer1[104] ));
 sg13g2_inv_1 _06990_ (.Y(_01120_),
    .A(\u_toplayer.reg_layer1[200] ));
 sg13g2_inv_1 _06991_ (.Y(_01121_),
    .A(\u_toplayer.reg_layer1[73] ));
 sg13g2_inv_1 _06992_ (.Y(_01122_),
    .A(\u_toplayer.reg_layer1[105] ));
 sg13g2_inv_1 _06993_ (.Y(_01123_),
    .A(\u_toplayer.reg_layer1[201] ));
 sg13g2_inv_1 _06994_ (.Y(_01124_),
    .A(\u_toplayer.reg_layer1[233] ));
 sg13g2_inv_1 _06995_ (.Y(_01125_),
    .A(\u_toplayer.reg_layer1[74] ));
 sg13g2_inv_1 _06996_ (.Y(_01126_),
    .A(\u_toplayer.reg_layer1[106] ));
 sg13g2_inv_1 _06997_ (.Y(_01127_),
    .A(\u_toplayer.reg_layer1[202] ));
 sg13g2_inv_1 _06998_ (.Y(_01128_),
    .A(\u_toplayer.reg_layer1[234] ));
 sg13g2_inv_1 _06999_ (.Y(_01129_),
    .A(\u_toplayer.reg_layer1[75] ));
 sg13g2_inv_1 _07000_ (.Y(_01130_),
    .A(\u_toplayer.reg_layer1[107] ));
 sg13g2_inv_1 _07001_ (.Y(_01131_),
    .A(\u_toplayer.reg_layer1[203] ));
 sg13g2_inv_1 _07002_ (.Y(_01132_),
    .A(\u_toplayer.reg_layer1[235] ));
 sg13g2_inv_1 _07003_ (.Y(_01133_),
    .A(\u_toplayer.reg_layer1[76] ));
 sg13g2_inv_1 _07004_ (.Y(_01134_),
    .A(\u_toplayer.reg_layer1[204] ));
 sg13g2_inv_1 _07005_ (.Y(_01135_),
    .A(\u_toplayer.reg_layer1[77] ));
 sg13g2_inv_1 _07006_ (.Y(_01136_),
    .A(\u_toplayer.reg_layer1[109] ));
 sg13g2_inv_1 _07007_ (.Y(_01137_),
    .A(\u_toplayer.reg_layer1[205] ));
 sg13g2_inv_1 _07008_ (.Y(_01138_),
    .A(\u_toplayer.reg_layer1[237] ));
 sg13g2_inv_1 _07009_ (.Y(_01139_),
    .A(\u_toplayer.reg_layer1[78] ));
 sg13g2_inv_1 _07010_ (.Y(_01140_),
    .A(\u_toplayer.reg_layer1[110] ));
 sg13g2_inv_1 _07011_ (.Y(_01141_),
    .A(\u_toplayer.reg_layer1[206] ));
 sg13g2_inv_1 _07012_ (.Y(_01142_),
    .A(\u_toplayer.reg_layer1[238] ));
 sg13g2_inv_1 _07013_ (.Y(_01143_),
    .A(\u_toplayer.reg_layer1[79] ));
 sg13g2_inv_1 _07014_ (.Y(_01144_),
    .A(\u_toplayer.reg_layer1[111] ));
 sg13g2_inv_1 _07015_ (.Y(_01145_),
    .A(\u_toplayer.reg_layer1[207] ));
 sg13g2_inv_1 _07016_ (.Y(_01146_),
    .A(\u_toplayer.reg_layer1[239] ));
 sg13g2_inv_1 _07017_ (.Y(_01147_),
    .A(_00049_));
 sg13g2_inv_1 _07018_ (.Y(_01148_),
    .A(\u_toplayer.u_layer2.u_neuron.mult[11] ));
 sg13g2_inv_2 _07019_ (.Y(_01149_),
    .A(net3193));
 sg13g2_inv_1 _07020_ (.Y(_01150_),
    .A(net3084));
 sg13g2_inv_1 _07021_ (.Y(_01151_),
    .A(net3083));
 sg13g2_inv_1 _07022_ (.Y(_01152_),
    .A(net1181));
 sg13g2_inv_1 _07023_ (.Y(_01153_),
    .A(net1143));
 sg13g2_inv_1 _07024_ (.Y(_01154_),
    .A(net3030));
 sg13g2_inv_1 _07025_ (.Y(_01155_),
    .A(net1172));
 sg13g2_inv_1 _07026_ (.Y(_01156_),
    .A(net1153));
 sg13g2_inv_1 _07027_ (.Y(_01157_),
    .A(net1084));
 sg13g2_inv_1 _07028_ (.Y(_01158_),
    .A(net1069));
 sg13g2_inv_1 _07029_ (.Y(_01159_),
    .A(net1049));
 sg13g2_inv_1 _07030_ (.Y(_01160_),
    .A(net1117));
 sg13g2_inv_1 _07031_ (.Y(_01161_),
    .A(net3027));
 sg13g2_inv_1 _07032_ (.Y(_01162_),
    .A(net3029));
 sg13g2_inv_1 _07033_ (.Y(_01163_),
    .A(net1112));
 sg13g2_inv_1 _07034_ (.Y(_01164_),
    .A(net1180));
 sg13g2_inv_1 _07035_ (.Y(_01165_),
    .A(net1154));
 sg13g2_inv_2 _07036_ (.Y(_01166_),
    .A(net1064));
 sg13g2_inv_1 _07037_ (.Y(_01167_),
    .A(net1074));
 sg13g2_inv_1 _07038_ (.Y(_01168_),
    .A(net1062));
 sg13g2_inv_1 _07039_ (.Y(_01169_),
    .A(net1185));
 sg13g2_inv_1 _07040_ (.Y(_01170_),
    .A(net3025));
 sg13g2_inv_1 _07041_ (.Y(_01171_),
    .A(net1120));
 sg13g2_inv_1 _07042_ (.Y(_01172_),
    .A(net886));
 sg13g2_inv_1 _07043_ (.Y(_01173_),
    .A(net1063));
 sg13g2_inv_1 _07044_ (.Y(_01174_),
    .A(net825));
 sg13g2_inv_1 _07045_ (.Y(_01175_),
    .A(net945));
 sg13g2_inv_2 _07046_ (.Y(_01176_),
    .A(net3050));
 sg13g2_inv_1 _07047_ (.Y(_01177_),
    .A(net910));
 sg13g2_inv_1 _07048_ (.Y(_01178_),
    .A(net3046));
 sg13g2_inv_1 _07049_ (.Y(_01179_),
    .A(net3045));
 sg13g2_inv_1 _07050_ (.Y(_01180_),
    .A(net3043));
 sg13g2_inv_1 _07051_ (.Y(_01181_),
    .A(net3040));
 sg13g2_inv_1 _07052_ (.Y(_01182_),
    .A(net3039));
 sg13g2_inv_1 _07053_ (.Y(_01183_),
    .A(net3037));
 sg13g2_inv_1 _07054_ (.Y(_01184_),
    .A(net3034));
 sg13g2_inv_1 _12781__2 (.Y(net21),
    .A(clknet_4_3_0_clk));
 sg13g2_nor2_1 _07056_ (.A(net120),
    .B(net121),
    .Y(_01185_));
 sg13g2_nand3_1 _07057_ (.B(\u_toplayer.delayed_done_layer2 ),
    .C(_01185_),
    .A(_01020_),
    .Y(_01186_));
 sg13g2_nand2_1 _07058_ (.Y(_01187_),
    .A(net840),
    .B(net116));
 sg13g2_nor2_1 _07059_ (.A(\u_toplayer.u_layer3.stateout[4] ),
    .B(net863),
    .Y(_01188_));
 sg13g2_nand3_1 _07060_ (.B(net939),
    .C(_01188_),
    .A(net895),
    .Y(_01189_));
 sg13g2_nor4_2 _07061_ (.A(net978),
    .B(_01186_),
    .C(_01187_),
    .Y(_01190_),
    .D(_01189_));
 sg13g2_nand2_1 _07062_ (.Y(_01191_),
    .A(\u_toplayer.u_layer3.stateout[2] ),
    .B(\u_toplayer.u_layer3.stateout[1] ));
 sg13g2_a21oi_1 _07063_ (.A1(_01188_),
    .A2(_01191_),
    .Y(_01192_),
    .B1(_01019_));
 sg13g2_nor3_1 _07064_ (.A(\u_toplayer.u_layer3.stateout[8] ),
    .B(_01186_),
    .C(_01192_),
    .Y(_01193_));
 sg13g2_nor2_2 _07065_ (.A(_01190_),
    .B(_01193_),
    .Y(_01194_));
 sg13g2_nand2_1 _07066_ (.Y(_01195_),
    .A(\u_toplayer.u_layer3.stateout[8] ),
    .B(_01194_));
 sg13g2_o21ai_1 _07067_ (.B1(_01195_),
    .Y(_00348_),
    .A1(net116),
    .A2(_01194_));
 sg13g2_nor2b_1 _07068_ (.A(_01194_),
    .B_N(net840),
    .Y(_01196_));
 sg13g2_and2_1 _07069_ (.A(net978),
    .B(_01196_),
    .X(_01197_));
 sg13g2_and2_1 _07070_ (.A(net939),
    .B(_01197_),
    .X(_01198_));
 sg13g2_nand3_1 _07071_ (.B(net863),
    .C(_01198_),
    .A(net1036),
    .Y(_01199_));
 sg13g2_a21oi_1 _07072_ (.A1(_01019_),
    .A2(_01199_),
    .Y(_00345_),
    .B1(_01190_));
 sg13g2_a21o_1 _07073_ (.A2(_01198_),
    .A1(net863),
    .B1(net1036),
    .X(_01200_));
 sg13g2_and2_1 _07074_ (.A(_01199_),
    .B(_01200_),
    .X(_00344_));
 sg13g2_xor2_1 _07075_ (.B(_01198_),
    .A(net863),
    .X(_00343_));
 sg13g2_nor2_1 _07076_ (.A(net939),
    .B(_01197_),
    .Y(_01201_));
 sg13g2_nor3_1 _07077_ (.A(_01190_),
    .B(_01198_),
    .C(net940),
    .Y(_00342_));
 sg13g2_nor2_1 _07078_ (.A(net978),
    .B(_01196_),
    .Y(_01202_));
 sg13g2_nor3_1 _07079_ (.A(_01190_),
    .B(_01197_),
    .C(_01202_),
    .Y(_00341_));
 sg13g2_xnor2_1 _07080_ (.Y(_00340_),
    .A(net840),
    .B(_01194_));
 sg13g2_nand2b_1 _07081_ (.Y(_01203_),
    .B(net1211),
    .A_N(\u_toplayer.u_layer3.neuron_index[0] ));
 sg13g2_nor3_1 _07082_ (.A(\u_toplayer.u_layer3.neuron_index[5] ),
    .B(\u_toplayer.u_layer3.neuron_index[4] ),
    .C(_01203_),
    .Y(_01204_));
 sg13g2_nand3_1 _07083_ (.B(\u_toplayer.delayed_done_layer2 ),
    .C(_01204_),
    .A(\u_toplayer.u_layer3.neuron_index[3] ),
    .Y(_01205_));
 sg13g2_o21ai_1 _07084_ (.B1(_01020_),
    .Y(_00323_),
    .A1(\u_toplayer.u_layer3.neuron_index[2] ),
    .A2(_01205_));
 sg13g2_nor3_2 _07085_ (.A(\u_toplayer.u_layer3.neuron_index[2] ),
    .B(\u_toplayer.u_layer3.neuron_index[1] ),
    .C(_01021_),
    .Y(_01206_));
 sg13g2_nor2b_1 _07086_ (.A(\u_toplayer.u_layer3.neuron_index[3] ),
    .B_N(_01206_),
    .Y(_01207_));
 sg13g2_nor2b_2 _07087_ (.A(\u_toplayer.u_layer3.neuron_index[4] ),
    .B_N(_01207_),
    .Y(_01208_));
 sg13g2_inv_1 _07088_ (.Y(_01209_),
    .A(_01208_));
 sg13g2_xnor2_1 _07089_ (.Y(_01210_),
    .A(\u_toplayer.u_layer3.neuron_index[5] ),
    .B(_01208_));
 sg13g2_nor2_2 _07090_ (.A(\u_toplayer.u_layer3.neuron_index[1] ),
    .B(\u_toplayer.u_layer3.neuron_index[0] ),
    .Y(_01211_));
 sg13g2_nand2_1 _07091_ (.Y(_01212_),
    .A(net993),
    .B(\u_toplayer.u_layer3.neuron_index[0] ));
 sg13g2_nor2b_1 _07092_ (.A(_01211_),
    .B_N(_01212_),
    .Y(_01213_));
 sg13g2_inv_1 _07093_ (.Y(_01214_),
    .A(_01213_));
 sg13g2_nor3_1 _07094_ (.A(\u_toplayer.u_layer3.neuron_index[5] ),
    .B(_00052_),
    .C(_01214_),
    .Y(_01215_));
 sg13g2_xnor2_1 _07095_ (.Y(_01216_),
    .A(\u_toplayer.u_layer3.neuron_index[3] ),
    .B(_01206_));
 sg13g2_xor2_1 _07096_ (.B(_01206_),
    .A(\u_toplayer.u_layer3.neuron_index[3] ),
    .X(_01217_));
 sg13g2_nor2_1 _07097_ (.A(\u_toplayer.u_layer3.neuron_index[2] ),
    .B(net2867),
    .Y(_01218_));
 sg13g2_nand4_1 _07098_ (.B(net895),
    .C(_01185_),
    .A(_01018_),
    .Y(_01219_),
    .D(_01190_));
 sg13g2_nor2b_2 _07099_ (.A(_01207_),
    .B_N(\u_toplayer.u_layer3.neuron_index[4] ),
    .Y(_01220_));
 sg13g2_nor3_2 _07100_ (.A(_01208_),
    .B(net2838),
    .C(_01220_),
    .Y(_01221_));
 sg13g2_nor3_2 _07101_ (.A(_01208_),
    .B(net2838),
    .C(_01220_),
    .Y(_01222_));
 sg13g2_nand3_1 _07102_ (.B(_01218_),
    .C(_01222_),
    .A(net2840),
    .Y(_01223_));
 sg13g2_nand2_1 _07103_ (.Y(_01224_),
    .A(net148),
    .B(_01223_));
 sg13g2_nand2_1 _07104_ (.Y(_01225_),
    .A(\u_toplayer.u_layer3.sum[7] ),
    .B(net2839));
 sg13g2_xor2_1 _07105_ (.B(_01211_),
    .A(\u_toplayer.u_layer3.neuron_index[2] ),
    .X(_01226_));
 sg13g2_nor4_2 _07106_ (.A(_01208_),
    .B(net2838),
    .C(_01220_),
    .Y(_01227_),
    .D(_01226_));
 sg13g2_nand2b_1 _07107_ (.Y(_01228_),
    .B(_01227_),
    .A_N(_01225_));
 sg13g2_o21ai_1 _07108_ (.B1(_01224_),
    .Y(_00322_),
    .A1(_01216_),
    .A2(_01228_));
 sg13g2_nand2_1 _07109_ (.Y(_01229_),
    .A(net388),
    .B(_01223_));
 sg13g2_nand2_1 _07110_ (.Y(_01230_),
    .A(\u_toplayer.u_layer3.sum[6] ),
    .B(net2841));
 sg13g2_nand3_1 _07111_ (.B(net2841),
    .C(_01227_),
    .A(\u_toplayer.u_layer3.sum[6] ),
    .Y(_01231_));
 sg13g2_o21ai_1 _07112_ (.B1(_01229_),
    .Y(_00321_),
    .A1(_01216_),
    .A2(_01231_));
 sg13g2_nand2_1 _07113_ (.Y(_01232_),
    .A(net196),
    .B(_01223_));
 sg13g2_nand2_1 _07114_ (.Y(_01233_),
    .A(\u_toplayer.u_layer3.sum[5] ),
    .B(net2839));
 sg13g2_nand3_1 _07115_ (.B(net2840),
    .C(_01227_),
    .A(\u_toplayer.u_layer3.sum[5] ),
    .Y(_01234_));
 sg13g2_o21ai_1 _07116_ (.B1(_01232_),
    .Y(_00320_),
    .A1(net2867),
    .A2(_01234_));
 sg13g2_nand2_1 _07117_ (.Y(_01235_),
    .A(net224),
    .B(_01223_));
 sg13g2_nand2_1 _07118_ (.Y(_01236_),
    .A(\u_toplayer.u_layer3.sum[4] ),
    .B(net2839));
 sg13g2_nand3_1 _07119_ (.B(net2840),
    .C(_01227_),
    .A(\u_toplayer.u_layer3.sum[4] ),
    .Y(_01237_));
 sg13g2_o21ai_1 _07120_ (.B1(_01235_),
    .Y(_00319_),
    .A1(net2867),
    .A2(_01237_));
 sg13g2_nand2_1 _07121_ (.Y(_01238_),
    .A(net346),
    .B(_01223_));
 sg13g2_nand2_1 _07122_ (.Y(_01239_),
    .A(\u_toplayer.u_layer3.sum[3] ),
    .B(net2839));
 sg13g2_nand3_1 _07123_ (.B(net2840),
    .C(_01227_),
    .A(\u_toplayer.u_layer3.sum[3] ),
    .Y(_01240_));
 sg13g2_o21ai_1 _07124_ (.B1(_01238_),
    .Y(_00318_),
    .A1(net2867),
    .A2(_01240_));
 sg13g2_nand2_1 _07125_ (.Y(_01241_),
    .A(net142),
    .B(_01223_));
 sg13g2_nand2_1 _07126_ (.Y(_01242_),
    .A(\u_toplayer.u_layer3.sum[2] ),
    .B(net2839));
 sg13g2_nand3_1 _07127_ (.B(net2840),
    .C(_01227_),
    .A(\u_toplayer.u_layer3.sum[2] ),
    .Y(_01243_));
 sg13g2_o21ai_1 _07128_ (.B1(_01241_),
    .Y(_00317_),
    .A1(net2867),
    .A2(_01243_));
 sg13g2_nand2_1 _07129_ (.Y(_01244_),
    .A(net212),
    .B(_01223_));
 sg13g2_nand2_1 _07130_ (.Y(_01245_),
    .A(\u_toplayer.u_layer3.sum[1] ),
    .B(net2839));
 sg13g2_nand3_1 _07131_ (.B(net2840),
    .C(_01227_),
    .A(\u_toplayer.u_layer3.sum[1] ),
    .Y(_01246_));
 sg13g2_o21ai_1 _07132_ (.B1(_01244_),
    .Y(_00316_),
    .A1(net2867),
    .A2(_01246_));
 sg13g2_nand2_1 _07133_ (.Y(_01247_),
    .A(net158),
    .B(_01223_));
 sg13g2_nand2_1 _07134_ (.Y(_01248_),
    .A(\u_toplayer.u_layer3.sum[0] ),
    .B(net2839));
 sg13g2_nand3_1 _07135_ (.B(net2840),
    .C(_01227_),
    .A(\u_toplayer.u_layer3.sum[0] ),
    .Y(_01249_));
 sg13g2_o21ai_1 _07136_ (.B1(_01247_),
    .Y(_00315_),
    .A1(net2867),
    .A2(_01249_));
 sg13g2_nand2_1 _07137_ (.Y(_01250_),
    .A(_01210_),
    .B(_01211_));
 sg13g2_and2_1 _07138_ (.A(net2867),
    .B(_01226_),
    .X(_01251_));
 sg13g2_nand2_2 _07139_ (.Y(_01252_),
    .A(_01222_),
    .B(_01251_));
 sg13g2_or2_2 _07140_ (.X(_01253_),
    .B(net2767),
    .A(net2768));
 sg13g2_mux2_1 _07141_ (.A0(\u_toplayer.u_layer3.sum[7] ),
    .A1(net791),
    .S(_01253_),
    .X(_00314_));
 sg13g2_mux2_1 _07142_ (.A0(\u_toplayer.u_layer3.sum[6] ),
    .A1(net848),
    .S(_01253_),
    .X(_00313_));
 sg13g2_mux2_1 _07143_ (.A0(\u_toplayer.u_layer3.sum[5] ),
    .A1(net811),
    .S(_01253_),
    .X(_00312_));
 sg13g2_mux2_1 _07144_ (.A0(\u_toplayer.u_layer3.sum[4] ),
    .A1(net818),
    .S(_01253_),
    .X(_00311_));
 sg13g2_mux2_1 _07145_ (.A0(\u_toplayer.u_layer3.sum[3] ),
    .A1(net786),
    .S(_01253_),
    .X(_00310_));
 sg13g2_mux2_1 _07146_ (.A0(\u_toplayer.u_layer3.sum[2] ),
    .A1(net744),
    .S(_01253_),
    .X(_00309_));
 sg13g2_mux2_1 _07147_ (.A0(\u_toplayer.u_layer3.sum[1] ),
    .A1(net752),
    .S(_01253_),
    .X(_00308_));
 sg13g2_mux2_1 _07148_ (.A0(\u_toplayer.u_layer3.sum[0] ),
    .A1(net787),
    .S(_01253_),
    .X(_00307_));
 sg13g2_nand3_1 _07149_ (.B(_01210_),
    .C(_01214_),
    .A(_01021_),
    .Y(_01254_));
 sg13g2_or2_2 _07150_ (.X(_01255_),
    .B(_01254_),
    .A(_01252_));
 sg13g2_mux2_1 _07151_ (.A0(\u_toplayer.u_layer3.sum[7] ),
    .A1(net884),
    .S(_01255_),
    .X(_00306_));
 sg13g2_mux2_1 _07152_ (.A0(\u_toplayer.u_layer3.sum[6] ),
    .A1(net851),
    .S(_01255_),
    .X(_00305_));
 sg13g2_mux2_1 _07153_ (.A0(\u_toplayer.u_layer3.sum[5] ),
    .A1(net855),
    .S(_01255_),
    .X(_00304_));
 sg13g2_mux2_1 _07154_ (.A0(\u_toplayer.u_layer3.sum[4] ),
    .A1(net887),
    .S(_01255_),
    .X(_00303_));
 sg13g2_mux2_1 _07155_ (.A0(\u_toplayer.u_layer3.sum[3] ),
    .A1(net894),
    .S(_01255_),
    .X(_00302_));
 sg13g2_mux2_1 _07156_ (.A0(\u_toplayer.u_layer3.sum[2] ),
    .A1(net869),
    .S(_01255_),
    .X(_00301_));
 sg13g2_mux2_1 _07157_ (.A0(\u_toplayer.u_layer3.sum[1] ),
    .A1(net852),
    .S(_01255_),
    .X(_00300_));
 sg13g2_mux2_1 _07158_ (.A0(\u_toplayer.u_layer3.sum[0] ),
    .A1(net862),
    .S(_01255_),
    .X(_00299_));
 sg13g2_nand2b_2 _07159_ (.Y(_01256_),
    .B(_01210_),
    .A_N(_01203_));
 sg13g2_or2_2 _07160_ (.X(_01257_),
    .B(_01256_),
    .A(_01252_));
 sg13g2_mux2_1 _07161_ (.A0(\u_toplayer.u_layer3.sum[7] ),
    .A1(net844),
    .S(_01257_),
    .X(_00298_));
 sg13g2_mux2_1 _07162_ (.A0(\u_toplayer.u_layer3.sum[6] ),
    .A1(net859),
    .S(_01257_),
    .X(_00297_));
 sg13g2_mux2_1 _07163_ (.A0(\u_toplayer.u_layer3.sum[5] ),
    .A1(net861),
    .S(_01257_),
    .X(_00296_));
 sg13g2_mux2_1 _07164_ (.A0(\u_toplayer.u_layer3.sum[4] ),
    .A1(net826),
    .S(_01257_),
    .X(_00295_));
 sg13g2_mux2_1 _07165_ (.A0(\u_toplayer.u_layer3.sum[3] ),
    .A1(net865),
    .S(_01257_),
    .X(_00294_));
 sg13g2_mux2_1 _07166_ (.A0(\u_toplayer.u_layer3.sum[2] ),
    .A1(net816),
    .S(_01257_),
    .X(_00293_));
 sg13g2_mux2_1 _07167_ (.A0(\u_toplayer.u_layer3.sum[1] ),
    .A1(net839),
    .S(_01257_),
    .X(_00292_));
 sg13g2_mux2_1 _07168_ (.A0(\u_toplayer.u_layer3.sum[0] ),
    .A1(net868),
    .S(_01257_),
    .X(_00291_));
 sg13g2_nand3_1 _07169_ (.B(_01222_),
    .C(_01251_),
    .A(net2839),
    .Y(_01258_));
 sg13g2_nand2_1 _07170_ (.Y(_01259_),
    .A(net144),
    .B(_01258_));
 sg13g2_o21ai_1 _07171_ (.B1(_01259_),
    .Y(_00290_),
    .A1(_01225_),
    .A2(_01252_));
 sg13g2_nand2_1 _07172_ (.Y(_01260_),
    .A(net217),
    .B(_01258_));
 sg13g2_o21ai_1 _07173_ (.B1(_01260_),
    .Y(_00289_),
    .A1(_01230_),
    .A2(net2767));
 sg13g2_nand2_1 _07174_ (.Y(_01261_),
    .A(net159),
    .B(_01258_));
 sg13g2_o21ai_1 _07175_ (.B1(_01261_),
    .Y(_00288_),
    .A1(_01233_),
    .A2(net2767));
 sg13g2_nand2_1 _07176_ (.Y(_01262_),
    .A(net147),
    .B(_01258_));
 sg13g2_o21ai_1 _07177_ (.B1(_01262_),
    .Y(_00287_),
    .A1(_01236_),
    .A2(net2767));
 sg13g2_nand2_1 _07178_ (.Y(_01263_),
    .A(net139),
    .B(_01258_));
 sg13g2_o21ai_1 _07179_ (.B1(_01263_),
    .Y(_00286_),
    .A1(_01239_),
    .A2(net2767));
 sg13g2_nand2_1 _07180_ (.Y(_01264_),
    .A(net162),
    .B(_01258_));
 sg13g2_o21ai_1 _07181_ (.B1(_01264_),
    .Y(_00285_),
    .A1(_01242_),
    .A2(net2767));
 sg13g2_nand2_1 _07182_ (.Y(_01265_),
    .A(net195),
    .B(_01258_));
 sg13g2_o21ai_1 _07183_ (.B1(_01265_),
    .Y(_00284_),
    .A1(_01245_),
    .A2(net2767));
 sg13g2_nand2_1 _07184_ (.Y(_01266_),
    .A(net152),
    .B(_01258_));
 sg13g2_o21ai_1 _07185_ (.B1(_01266_),
    .Y(_00283_),
    .A1(_01248_),
    .A2(net2767));
 sg13g2_nor2_2 _07186_ (.A(net2866),
    .B(_01226_),
    .Y(_01267_));
 sg13g2_nor4_2 _07187_ (.A(\u_toplayer.u_layer3.neuron_index[4] ),
    .B(net2866),
    .C(_01219_),
    .Y(_01268_),
    .D(_01226_));
 sg13g2_nand3_1 _07188_ (.B(_01211_),
    .C(_01268_),
    .A(_01210_),
    .Y(_01269_));
 sg13g2_nand2_1 _07189_ (.Y(_01270_),
    .A(net135),
    .B(_01269_));
 sg13g2_nand3_1 _07190_ (.B(_01221_),
    .C(_01267_),
    .A(\u_toplayer.u_layer3.sum[7] ),
    .Y(_01271_));
 sg13g2_o21ai_1 _07191_ (.B1(_01270_),
    .Y(_00282_),
    .A1(_01250_),
    .A2(_01271_));
 sg13g2_nand2_1 _07192_ (.Y(_01272_),
    .A(net129),
    .B(_01269_));
 sg13g2_nand3_1 _07193_ (.B(_01221_),
    .C(_01267_),
    .A(\u_toplayer.u_layer3.sum[6] ),
    .Y(_01273_));
 sg13g2_o21ai_1 _07194_ (.B1(_01272_),
    .Y(_00281_),
    .A1(net2768),
    .A2(_01273_));
 sg13g2_nand2_1 _07195_ (.Y(_01274_),
    .A(net134),
    .B(_01269_));
 sg13g2_nand3_1 _07196_ (.B(_01221_),
    .C(_01267_),
    .A(\u_toplayer.u_layer3.sum[5] ),
    .Y(_01275_));
 sg13g2_o21ai_1 _07197_ (.B1(_01274_),
    .Y(_00280_),
    .A1(net2768),
    .A2(_01275_));
 sg13g2_nand2_1 _07198_ (.Y(_01276_),
    .A(net138),
    .B(_01269_));
 sg13g2_nand3_1 _07199_ (.B(_01221_),
    .C(_01267_),
    .A(\u_toplayer.u_layer3.sum[4] ),
    .Y(_01277_));
 sg13g2_o21ai_1 _07200_ (.B1(_01276_),
    .Y(_00279_),
    .A1(net2768),
    .A2(_01277_));
 sg13g2_nand2_1 _07201_ (.Y(_01278_),
    .A(net161),
    .B(_01269_));
 sg13g2_nand3_1 _07202_ (.B(_01221_),
    .C(_01267_),
    .A(\u_toplayer.u_layer3.sum[3] ),
    .Y(_01279_));
 sg13g2_o21ai_1 _07203_ (.B1(_01278_),
    .Y(_00278_),
    .A1(net2768),
    .A2(_01279_));
 sg13g2_nand2_1 _07204_ (.Y(_01280_),
    .A(net137),
    .B(_01269_));
 sg13g2_nand3_1 _07205_ (.B(_01221_),
    .C(_01267_),
    .A(\u_toplayer.u_layer3.sum[2] ),
    .Y(_01281_));
 sg13g2_o21ai_1 _07206_ (.B1(_01280_),
    .Y(_00277_),
    .A1(net2768),
    .A2(_01281_));
 sg13g2_nand2_1 _07207_ (.Y(_01282_),
    .A(net146),
    .B(_01269_));
 sg13g2_nand3_1 _07208_ (.B(_01221_),
    .C(_01267_),
    .A(\u_toplayer.u_layer3.sum[1] ),
    .Y(_01283_));
 sg13g2_o21ai_1 _07209_ (.B1(_01282_),
    .Y(_00276_),
    .A1(net2768),
    .A2(_01283_));
 sg13g2_nand2_1 _07210_ (.Y(_01284_),
    .A(net133),
    .B(_01269_));
 sg13g2_nand3_1 _07211_ (.B(_01221_),
    .C(_01267_),
    .A(\u_toplayer.u_layer3.sum[0] ),
    .Y(_01285_));
 sg13g2_o21ai_1 _07212_ (.B1(_01284_),
    .Y(_00275_),
    .A1(net2768),
    .A2(_01285_));
 sg13g2_nand2b_2 _07213_ (.Y(_01286_),
    .B(_01268_),
    .A_N(net2766));
 sg13g2_nand2_1 _07214_ (.Y(_01287_),
    .A(net153),
    .B(_01286_));
 sg13g2_o21ai_1 _07215_ (.B1(_01287_),
    .Y(_00274_),
    .A1(_01254_),
    .A2(_01271_));
 sg13g2_nand2_1 _07216_ (.Y(_01288_),
    .A(net252),
    .B(_01286_));
 sg13g2_o21ai_1 _07217_ (.B1(_01288_),
    .Y(_00273_),
    .A1(net2766),
    .A2(_01273_));
 sg13g2_nand2_1 _07218_ (.Y(_01289_),
    .A(net160),
    .B(_01286_));
 sg13g2_o21ai_1 _07219_ (.B1(_01289_),
    .Y(_00272_),
    .A1(net2766),
    .A2(_01275_));
 sg13g2_nand2_1 _07220_ (.Y(_01290_),
    .A(net594),
    .B(_01286_));
 sg13g2_o21ai_1 _07221_ (.B1(_01290_),
    .Y(_00271_),
    .A1(net2766),
    .A2(_01277_));
 sg13g2_nand2_1 _07222_ (.Y(_01291_),
    .A(net187),
    .B(_01286_));
 sg13g2_o21ai_1 _07223_ (.B1(_01291_),
    .Y(_00270_),
    .A1(net2766),
    .A2(_01279_));
 sg13g2_nand2_1 _07224_ (.Y(_01292_),
    .A(net380),
    .B(_01286_));
 sg13g2_o21ai_1 _07225_ (.B1(_01292_),
    .Y(_00269_),
    .A1(net2766),
    .A2(_01281_));
 sg13g2_nand2_1 _07226_ (.Y(_01293_),
    .A(net170),
    .B(_01286_));
 sg13g2_o21ai_1 _07227_ (.B1(_01293_),
    .Y(_00268_),
    .A1(net2766),
    .A2(_01283_));
 sg13g2_nand2_1 _07228_ (.Y(_01294_),
    .A(net145),
    .B(_01286_));
 sg13g2_o21ai_1 _07229_ (.B1(_01294_),
    .Y(_00267_),
    .A1(net2766),
    .A2(_01285_));
 sg13g2_nand2b_2 _07230_ (.Y(_01295_),
    .B(_01268_),
    .A_N(net2765));
 sg13g2_nand2_1 _07231_ (.Y(_01296_),
    .A(net190),
    .B(_01295_));
 sg13g2_o21ai_1 _07232_ (.B1(_01296_),
    .Y(_00266_),
    .A1(_01256_),
    .A2(_01271_));
 sg13g2_nand2_1 _07233_ (.Y(_01297_),
    .A(net192),
    .B(_01295_));
 sg13g2_o21ai_1 _07234_ (.B1(_01297_),
    .Y(_00265_),
    .A1(net2765),
    .A2(_01273_));
 sg13g2_nand2_1 _07235_ (.Y(_01298_),
    .A(net143),
    .B(_01295_));
 sg13g2_o21ai_1 _07236_ (.B1(_01298_),
    .Y(_00264_),
    .A1(net2765),
    .A2(_01275_));
 sg13g2_nand2_1 _07237_ (.Y(_01299_),
    .A(net140),
    .B(_01295_));
 sg13g2_o21ai_1 _07238_ (.B1(_01299_),
    .Y(_00263_),
    .A1(net2765),
    .A2(_01277_));
 sg13g2_nand2_1 _07239_ (.Y(_01300_),
    .A(net168),
    .B(_01295_));
 sg13g2_o21ai_1 _07240_ (.B1(_01300_),
    .Y(_00262_),
    .A1(net2765),
    .A2(_01279_));
 sg13g2_nand2_1 _07241_ (.Y(_01301_),
    .A(net171),
    .B(_01295_));
 sg13g2_o21ai_1 _07242_ (.B1(_01301_),
    .Y(_00261_),
    .A1(net2765),
    .A2(_01281_));
 sg13g2_nand2_1 _07243_ (.Y(_01302_),
    .A(net157),
    .B(_01295_));
 sg13g2_o21ai_1 _07244_ (.B1(_01302_),
    .Y(_00260_),
    .A1(net2765),
    .A2(_01283_));
 sg13g2_nand2_1 _07245_ (.Y(_01303_),
    .A(net426),
    .B(_01295_));
 sg13g2_o21ai_1 _07246_ (.B1(_01303_),
    .Y(_00259_),
    .A1(net2765),
    .A2(_01285_));
 sg13g2_nand2_2 _07247_ (.Y(_01304_),
    .A(net2840),
    .B(_01268_));
 sg13g2_nand2_1 _07248_ (.Y(_01305_),
    .A(net249),
    .B(_01304_));
 sg13g2_o21ai_1 _07249_ (.B1(_01305_),
    .Y(_00258_),
    .A1(_01217_),
    .A2(_01228_));
 sg13g2_nand2_1 _07250_ (.Y(_01306_),
    .A(net155),
    .B(_01304_));
 sg13g2_o21ai_1 _07251_ (.B1(_01306_),
    .Y(_00257_),
    .A1(net2866),
    .A2(_01231_));
 sg13g2_nand2_1 _07252_ (.Y(_01307_),
    .A(net149),
    .B(_01304_));
 sg13g2_o21ai_1 _07253_ (.B1(_01307_),
    .Y(_00256_),
    .A1(net2866),
    .A2(_01234_));
 sg13g2_nand2_1 _07254_ (.Y(_01308_),
    .A(net151),
    .B(_01304_));
 sg13g2_o21ai_1 _07255_ (.B1(_01308_),
    .Y(_00255_),
    .A1(net2866),
    .A2(_01237_));
 sg13g2_nand2_1 _07256_ (.Y(_01309_),
    .A(net141),
    .B(_01304_));
 sg13g2_o21ai_1 _07257_ (.B1(_01309_),
    .Y(_00254_),
    .A1(net2866),
    .A2(_01240_));
 sg13g2_nand2_1 _07258_ (.Y(_01310_),
    .A(net240),
    .B(_01304_));
 sg13g2_o21ai_1 _07259_ (.B1(_01310_),
    .Y(_00253_),
    .A1(net2866),
    .A2(_01243_));
 sg13g2_nand2_1 _07260_ (.Y(_01311_),
    .A(net211),
    .B(_01304_));
 sg13g2_o21ai_1 _07261_ (.B1(_01311_),
    .Y(_00252_),
    .A1(net2866),
    .A2(_01246_));
 sg13g2_nand2_1 _07262_ (.Y(_01312_),
    .A(net150),
    .B(_01304_));
 sg13g2_o21ai_1 _07263_ (.B1(_01312_),
    .Y(_00251_),
    .A1(_01217_),
    .A2(_01249_));
 sg13g2_nor4_2 _07264_ (.A(\u_toplayer.u_layer3.neuron_index[5] ),
    .B(\u_toplayer.u_layer3.neuron_index[0] ),
    .C(_01209_),
    .Y(_01313_),
    .D(net2838));
 sg13g2_mux2_1 _07265_ (.A0(net504),
    .A1(\u_toplayer.u_layer3.sum[7] ),
    .S(_01313_),
    .X(_00250_));
 sg13g2_mux2_1 _07266_ (.A0(net177),
    .A1(\u_toplayer.u_layer3.sum[6] ),
    .S(_01313_),
    .X(_00249_));
 sg13g2_mux2_1 _07267_ (.A0(net281),
    .A1(\u_toplayer.u_layer3.sum[5] ),
    .S(_01313_),
    .X(_00248_));
 sg13g2_mux2_1 _07268_ (.A0(net165),
    .A1(\u_toplayer.u_layer3.sum[4] ),
    .S(_01313_),
    .X(_00247_));
 sg13g2_mux2_1 _07269_ (.A0(net591),
    .A1(\u_toplayer.u_layer3.sum[3] ),
    .S(_01313_),
    .X(_00246_));
 sg13g2_mux2_1 _07270_ (.A0(net261),
    .A1(\u_toplayer.u_layer3.sum[2] ),
    .S(_01313_),
    .X(_00245_));
 sg13g2_mux2_1 _07271_ (.A0(net395),
    .A1(\u_toplayer.u_layer3.sum[1] ),
    .S(_01313_),
    .X(_00244_));
 sg13g2_mux2_1 _07272_ (.A0(net164),
    .A1(\u_toplayer.u_layer3.sum[0] ),
    .S(_01313_),
    .X(_00243_));
 sg13g2_nor2_2 _07273_ (.A(_01212_),
    .B(_01219_),
    .Y(_01314_));
 sg13g2_nand3_1 _07274_ (.B(\u_toplayer.u_layer3.neuron_index[2] ),
    .C(_01314_),
    .A(net1190),
    .Y(_01315_));
 sg13g2_nand4_1 _07275_ (.B(\u_toplayer.u_layer3.neuron_index[3] ),
    .C(\u_toplayer.u_layer3.neuron_index[2] ),
    .A(\u_toplayer.u_layer3.neuron_index[4] ),
    .Y(_01316_),
    .D(_01314_));
 sg13g2_xnor2_1 _07276_ (.Y(_00226_),
    .A(net1024),
    .B(_01316_));
 sg13g2_xnor2_1 _07277_ (.Y(_00225_),
    .A(net1034),
    .B(_01315_));
 sg13g2_a21o_1 _07278_ (.A2(_01314_),
    .A1(net1098),
    .B1(net1190),
    .X(_01317_));
 sg13g2_and2_1 _07279_ (.A(_01315_),
    .B(_01317_),
    .X(_00224_));
 sg13g2_xor2_1 _07280_ (.B(_01314_),
    .A(net1098),
    .X(_00223_));
 sg13g2_nand2_1 _07281_ (.Y(_01318_),
    .A(net993),
    .B(net2838));
 sg13g2_o21ai_1 _07282_ (.B1(_01318_),
    .Y(_00222_),
    .A1(_01214_),
    .A2(net2838));
 sg13g2_nand2_1 _07283_ (.Y(_01319_),
    .A(\u_toplayer.u_layer3.neuron_index[0] ),
    .B(net2838));
 sg13g2_o21ai_1 _07284_ (.B1(_01319_),
    .Y(_00221_),
    .A1(_01021_),
    .A2(net2838));
 sg13g2_or2_1 _07285_ (.X(_00010_),
    .B(net124),
    .A(net812));
 sg13g2_or2_2 _07286_ (.X(_00009_),
    .B(net130),
    .A(net925));
 sg13g2_or2_1 _07287_ (.X(_00011_),
    .B(net907),
    .A(net126));
 sg13g2_nor2b_1 _07288_ (.A(net3187),
    .B_N(net3024),
    .Y(_00025_));
 sg13g2_nor2b_2 _07289_ (.A(net3185),
    .B_N(net3187),
    .Y(_01320_));
 sg13g2_nor2b_1 _07290_ (.A(net3188),
    .B_N(net3185),
    .Y(_01321_));
 sg13g2_nand2_1 _07291_ (.Y(_01322_),
    .A(net3024),
    .B(net3016));
 sg13g2_o21ai_1 _07292_ (.B1(net3024),
    .Y(_01323_),
    .A1(_01320_),
    .A2(net3016));
 sg13g2_inv_1 _07293_ (.Y(_00026_),
    .A(_01323_));
 sg13g2_and2_1 _07294_ (.A(net3187),
    .B(net3184),
    .X(_01324_));
 sg13g2_o21ai_1 _07295_ (.B1(net3024),
    .Y(_01325_),
    .A1(net3182),
    .A2(net3012));
 sg13g2_a21oi_1 _07296_ (.A1(net3182),
    .A2(net3013),
    .Y(_00027_),
    .B1(_01325_));
 sg13g2_nor2b_1 _07297_ (.A(net958),
    .B_N(net3013),
    .Y(_01326_));
 sg13g2_o21ai_1 _07298_ (.B1(net3024),
    .Y(_01327_),
    .A1(net3180),
    .A2(_01326_));
 sg13g2_a21oi_1 _07299_ (.A1(net3180),
    .A2(_01326_),
    .Y(_00028_),
    .B1(_01327_));
 sg13g2_nand2b_2 _07300_ (.Y(_01328_),
    .B(\u_toplayer.delayed_done_layer2 ),
    .A_N(net881));
 sg13g2_nor2b_1 _07301_ (.A(net1178),
    .B_N(\u_toplayer.delayed_done_layer2 ),
    .Y(_01329_));
 sg13g2_nor2b_1 _07302_ (.A(net3100),
    .B_N(_01329_),
    .Y(_01330_));
 sg13g2_nor2_1 _07303_ (.A(net3112),
    .B(net3127),
    .Y(_01331_));
 sg13g2_o21ai_1 _07304_ (.B1(_01330_),
    .Y(_01332_),
    .A1(net3018),
    .A2(_01331_));
 sg13g2_a21oi_1 _07305_ (.A1(_01328_),
    .A2(_01332_),
    .Y(_00019_),
    .B1(net3127));
 sg13g2_nor2_2 _07306_ (.A(net3102),
    .B(net3100),
    .Y(_01333_));
 sg13g2_nand2b_1 _07307_ (.Y(_01334_),
    .B(_01333_),
    .A_N(net3098));
 sg13g2_and2_1 _07308_ (.A(net3112),
    .B(net3127),
    .X(_01335_));
 sg13g2_nand2_2 _07309_ (.Y(_01336_),
    .A(net3112),
    .B(net3127));
 sg13g2_nand3b_1 _07310_ (.B(_01336_),
    .C(\u_toplayer.delayed_done_layer2 ),
    .Y(_01337_),
    .A_N(_01331_));
 sg13g2_a21oi_1 _07311_ (.A1(net881),
    .A2(_01334_),
    .Y(_00020_),
    .B1(_01337_));
 sg13g2_xnor2_1 _07312_ (.Y(_01338_),
    .A(net3102),
    .B(net3001));
 sg13g2_a21oi_1 _07313_ (.A1(_01328_),
    .A2(_01332_),
    .Y(_00021_),
    .B1(_01338_));
 sg13g2_nor2_1 _07314_ (.A(net1005),
    .B(_01336_),
    .Y(_01339_));
 sg13g2_xnor2_1 _07315_ (.Y(_01340_),
    .A(net3100),
    .B(_01339_));
 sg13g2_nor2_1 _07316_ (.A(_01328_),
    .B(_01340_),
    .Y(_00022_));
 sg13g2_nor3_1 _07317_ (.A(_00037_),
    .B(net964),
    .C(_01336_),
    .Y(_01341_));
 sg13g2_xnor2_1 _07318_ (.Y(_01342_),
    .A(net3098),
    .B(net965));
 sg13g2_nor2_1 _07319_ (.A(_01328_),
    .B(net966),
    .Y(_00023_));
 sg13g2_a21oi_1 _07320_ (.A1(_01065_),
    .A2(_01341_),
    .Y(_01343_),
    .B1(\u_toplayer.u_layer3.u_neuron.instCtrl.state[5] ));
 sg13g2_o21ai_1 _07321_ (.B1(_01330_),
    .Y(_01344_),
    .A1(_00037_),
    .A2(_01331_));
 sg13g2_a21oi_1 _07322_ (.A1(_01328_),
    .A2(_01344_),
    .Y(_00024_),
    .B1(net682));
 sg13g2_nand2b_2 _07323_ (.Y(_01345_),
    .B(net1174),
    .A_N(net1071));
 sg13g2_nor3_1 _07324_ (.A(_01031_),
    .B(net3238),
    .C(net3234),
    .Y(_01346_));
 sg13g2_nor2_2 _07325_ (.A(net3255),
    .B(net3277),
    .Y(_01347_));
 sg13g2_o21ai_1 _07326_ (.B1(_01346_),
    .Y(_01348_),
    .A1(net3020),
    .A2(_01347_));
 sg13g2_a21oi_1 _07327_ (.A1(_01345_),
    .A2(_01348_),
    .Y(_00013_),
    .B1(net3277));
 sg13g2_nor2_1 _07328_ (.A(net3239),
    .B(net3235),
    .Y(_01349_));
 sg13g2_nor3_1 _07329_ (.A(net3242),
    .B(net3238),
    .C(net3234),
    .Y(_01350_));
 sg13g2_nor2b_1 _07330_ (.A(_01350_),
    .B_N(net1071),
    .Y(_01351_));
 sg13g2_and2_1 _07331_ (.A(net3245),
    .B(net3258),
    .X(_01352_));
 sg13g2_nand2_2 _07332_ (.Y(_01353_),
    .A(net3255),
    .B(net3277));
 sg13g2_nor4_1 _07333_ (.A(_01031_),
    .B(_01347_),
    .C(net1072),
    .D(net2993),
    .Y(_00014_));
 sg13g2_xnor2_1 _07334_ (.Y(_01354_),
    .A(net3242),
    .B(net2993));
 sg13g2_a21oi_1 _07335_ (.A1(_01345_),
    .A2(_01348_),
    .Y(_00015_),
    .B1(_01354_));
 sg13g2_nor2_1 _07336_ (.A(net999),
    .B(_01353_),
    .Y(_01355_));
 sg13g2_xnor2_1 _07337_ (.Y(_01356_),
    .A(net3238),
    .B(_01355_));
 sg13g2_nor2_1 _07338_ (.A(_01345_),
    .B(net1000),
    .Y(_00016_));
 sg13g2_nor3_1 _07339_ (.A(_00040_),
    .B(net931),
    .C(_01353_),
    .Y(_01357_));
 sg13g2_xnor2_1 _07340_ (.Y(_01358_),
    .A(net3234),
    .B(net932));
 sg13g2_nor2_1 _07341_ (.A(_01345_),
    .B(net933),
    .Y(_00017_));
 sg13g2_a21oi_1 _07342_ (.A1(_01117_),
    .A2(_01357_),
    .Y(_01359_),
    .B1(\u_toplayer.u_layer2.u_neuron.instCtrl.state[5] ));
 sg13g2_o21ai_1 _07343_ (.B1(_01346_),
    .Y(_01360_),
    .A1(_00040_),
    .A2(_01347_));
 sg13g2_a21oi_1 _07344_ (.A1(_01345_),
    .A2(_01360_),
    .Y(_00018_),
    .B1(net872));
 sg13g2_nand2_1 _07345_ (.Y(_01361_),
    .A(net3021),
    .B(net118));
 sg13g2_nor3_1 _07346_ (.A(\u_toplayer.u_layer1.u_neuron.instCtrl.state[4] ),
    .B(\u_toplayer.u_layer1.u_neuron.instCtrl.state[6] ),
    .C(\u_toplayer.u_layer1.u_neuron.instCtrl.state[5] ),
    .Y(_01362_));
 sg13g2_nor3_1 _07347_ (.A(net3021),
    .B(\u_toplayer.u_layer1.u_neuron.instCtrl.state[2] ),
    .C(\u_toplayer.u_layer1.u_neuron.instCtrl.state[3] ),
    .Y(_01363_));
 sg13g2_nand3_1 _07348_ (.B(_01362_),
    .C(_01363_),
    .A(_00044_),
    .Y(_01364_));
 sg13g2_o21ai_1 _07349_ (.B1(_01361_),
    .Y(_00000_),
    .A1(\u_toplayer.u_layer1.u_neuron.instCtrl.state[0] ),
    .A2(_01364_));
 sg13g2_nand2_1 _07350_ (.Y(_01365_),
    .A(\u_toplayer.u_layer1.u_neuron.instCtrl.state[0] ),
    .B(_01030_));
 sg13g2_xor2_1 _07351_ (.B(net1065),
    .A(\u_toplayer.u_layer1.u_neuron.instCtrl.state[0] ),
    .X(_01366_));
 sg13g2_nand2_1 _07352_ (.Y(_01367_),
    .A(\u_toplayer.u_layer1.u_neuron.instCtrl.state[0] ),
    .B(\u_toplayer.u_layer1.u_neuron.instCtrl.state[1] ));
 sg13g2_nand2b_1 _07353_ (.Y(_01368_),
    .B(_01367_),
    .A_N(net1106));
 sg13g2_nand3b_1 _07354_ (.B(_00044_),
    .C(_01362_),
    .Y(_01369_),
    .A_N(\u_toplayer.u_layer1.u_neuron.instCtrl.state[3] ));
 sg13g2_o21ai_1 _07355_ (.B1(net1039),
    .Y(_01370_),
    .A1(_01368_),
    .A2(_01369_));
 sg13g2_and2_1 _07356_ (.A(net1066),
    .B(net1040),
    .X(_00001_));
 sg13g2_nand3_1 _07357_ (.B(net1106),
    .C(net1065),
    .A(\u_toplayer.u_layer1.u_neuron.instCtrl.state[0] ),
    .Y(_01371_));
 sg13g2_and3_1 _07358_ (.X(_00002_),
    .A(net3229),
    .B(_01368_),
    .C(net1107));
 sg13g2_nor2_1 _07359_ (.A(_00045_),
    .B(_01367_),
    .Y(_01372_));
 sg13g2_o21ai_1 _07360_ (.B1(net3229),
    .Y(_01373_),
    .A1(net918),
    .A2(_01372_));
 sg13g2_a21oi_1 _07361_ (.A1(net918),
    .A2(_01372_),
    .Y(_00003_),
    .B1(_01373_));
 sg13g2_nor3_1 _07362_ (.A(_00045_),
    .B(_00046_),
    .C(_01367_),
    .Y(_01374_));
 sg13g2_o21ai_1 _07363_ (.B1(net3229),
    .Y(_01375_),
    .A1(net511),
    .A2(_01374_));
 sg13g2_a21oi_1 _07364_ (.A1(net511),
    .A2(_01374_),
    .Y(_00004_),
    .B1(_01375_));
 sg13g2_nor2b_1 _07365_ (.A(_00047_),
    .B_N(_01374_),
    .Y(_01376_));
 sg13g2_o21ai_1 _07366_ (.B1(net3229),
    .Y(_01377_),
    .A1(net569),
    .A2(_01376_));
 sg13g2_a21oi_1 _07367_ (.A1(net569),
    .A2(_01376_),
    .Y(_00005_),
    .B1(_01377_));
 sg13g2_nor2b_2 _07368_ (.A(_00048_),
    .B_N(_01376_),
    .Y(_01378_));
 sg13g2_o21ai_1 _07369_ (.B1(net3229),
    .Y(_01379_),
    .A1(net554),
    .A2(_01378_));
 sg13g2_a21oi_1 _07370_ (.A1(net554),
    .A2(_01378_),
    .Y(_00006_),
    .B1(_01379_));
 sg13g2_a21oi_1 _07371_ (.A1(_01147_),
    .A2(_01378_),
    .Y(_01380_),
    .B1(net770));
 sg13g2_nand3_1 _07372_ (.B(_01147_),
    .C(_01378_),
    .A(net770),
    .Y(_01381_));
 sg13g2_nand2_1 _07373_ (.Y(_01382_),
    .A(net3229),
    .B(_01381_));
 sg13g2_nor2_1 _07374_ (.A(net771),
    .B(_01382_),
    .Y(_00007_));
 sg13g2_nand2_1 _07375_ (.Y(_01383_),
    .A(net3021),
    .B(_01381_));
 sg13g2_and2_1 _07376_ (.A(net1040),
    .B(_01383_),
    .X(_00008_));
 sg13g2_nor2_1 _07377_ (.A(\u_toplayer.u_layer1.neuron_index[1] ),
    .B(net3055),
    .Y(_01384_));
 sg13g2_nor3_1 _07378_ (.A(net3057),
    .B(\u_toplayer.u_layer1.neuron_index[1] ),
    .C(net3055),
    .Y(_01385_));
 sg13g2_nor2b_1 _07379_ (.A(net3053),
    .B_N(net2980),
    .Y(_01386_));
 sg13g2_nor2_1 _07380_ (.A(net3053),
    .B(net1028),
    .Y(_01387_));
 sg13g2_nand3_1 _07381_ (.B(net2980),
    .C(_01387_),
    .A(net1010),
    .Y(_01388_));
 sg13g2_nand2b_1 _07382_ (.Y(_00012_),
    .B(_01388_),
    .A_N(net943));
 sg13g2_and2_1 _07383_ (.A(net3179),
    .B(net3182),
    .X(_01389_));
 sg13g2_nand2_1 _07384_ (.Y(_01390_),
    .A(net3179),
    .B(net3182));
 sg13g2_nand2_1 _07385_ (.Y(_01391_),
    .A(net3024),
    .B(net2977));
 sg13g2_o21ai_1 _07386_ (.B1(\u_toplayer.delayed_done_layer3 ),
    .Y(_01392_),
    .A1(net3016),
    .A2(net2977));
 sg13g2_nand2_1 _07387_ (.Y(_01393_),
    .A(net901),
    .B(net2941));
 sg13g2_nand2_1 _07388_ (.Y(_01394_),
    .A(net3346),
    .B(net3225));
 sg13g2_o21ai_1 _07389_ (.B1(_01393_),
    .Y(_00149_),
    .A1(net2943),
    .A2(_01394_));
 sg13g2_a22oi_1 _07390_ (.Y(_01395_),
    .B1(net3221),
    .B2(net3346),
    .A2(net3336),
    .A1(net3224));
 sg13g2_and4_1 _07391_ (.A(net3346),
    .B(net3224),
    .C(net3336),
    .D(net3221),
    .X(_01396_));
 sg13g2_nor3_1 _07392_ (.A(net2943),
    .B(_01395_),
    .C(_01396_),
    .Y(_01397_));
 sg13g2_a21o_1 _07393_ (.A2(net2941),
    .A1(net991),
    .B1(_01397_),
    .X(_00150_));
 sg13g2_and4_1 _07394_ (.A(net3224),
    .B(net3335),
    .C(net3222),
    .D(net3322),
    .X(_01398_));
 sg13g2_a22oi_1 _07395_ (.Y(_01399_),
    .B1(net3322),
    .B2(net3224),
    .A2(net3222),
    .A1(net3335));
 sg13g2_nand2_1 _07396_ (.Y(_01400_),
    .A(net3345),
    .B(net3220));
 sg13g2_nor3_1 _07397_ (.A(_01398_),
    .B(_01399_),
    .C(_01400_),
    .Y(_01401_));
 sg13g2_o21ai_1 _07398_ (.B1(_01400_),
    .Y(_01402_),
    .A1(_01398_),
    .A2(_01399_));
 sg13g2_nor2b_1 _07399_ (.A(_01401_),
    .B_N(_01402_),
    .Y(_01403_));
 sg13g2_nand2_2 _07400_ (.Y(_01404_),
    .A(_01396_),
    .B(_01403_));
 sg13g2_nor2_1 _07401_ (.A(_01396_),
    .B(_01403_),
    .Y(_01405_));
 sg13g2_nor2_1 _07402_ (.A(net2943),
    .B(_01405_),
    .Y(_01406_));
 sg13g2_a22oi_1 _07403_ (.Y(_01407_),
    .B1(_01404_),
    .B2(_01406_),
    .A2(net2941),
    .A1(net920));
 sg13g2_inv_1 _07404_ (.Y(_00151_),
    .A(_01407_));
 sg13g2_nand2_1 _07405_ (.Y(_01408_),
    .A(net836),
    .B(net2940));
 sg13g2_and2_1 _07406_ (.A(net3345),
    .B(net3217),
    .X(_01409_));
 sg13g2_nand2_1 _07407_ (.Y(_01410_),
    .A(net3345),
    .B(net3217));
 sg13g2_nand2_1 _07408_ (.Y(_01411_),
    .A(net3336),
    .B(net3220));
 sg13g2_and4_1 _07409_ (.A(net3224),
    .B(net3221),
    .C(net3322),
    .D(net3310),
    .X(_01412_));
 sg13g2_nand4_1 _07410_ (.B(net3221),
    .C(net3321),
    .A(net3225),
    .Y(_01413_),
    .D(net3310));
 sg13g2_a22oi_1 _07411_ (.Y(_01414_),
    .B1(net3310),
    .B2(net3224),
    .A2(net3322),
    .A1(net3221));
 sg13g2_or3_1 _07412_ (.A(_01411_),
    .B(_01412_),
    .C(_01414_),
    .X(_01415_));
 sg13g2_o21ai_1 _07413_ (.B1(_01411_),
    .Y(_01416_),
    .A1(_01412_),
    .A2(_01414_));
 sg13g2_nand3_1 _07414_ (.B(_01415_),
    .C(_01416_),
    .A(_01398_),
    .Y(_01417_));
 sg13g2_inv_1 _07415_ (.Y(_01418_),
    .A(_01417_));
 sg13g2_a21oi_1 _07416_ (.A1(_01415_),
    .A2(_01416_),
    .Y(_01419_),
    .B1(_01398_));
 sg13g2_nand3b_1 _07417_ (.B(_01409_),
    .C(_01417_),
    .Y(_01420_),
    .A_N(_01419_));
 sg13g2_o21ai_1 _07418_ (.B1(_01410_),
    .Y(_01421_),
    .A1(_01418_),
    .A2(_01419_));
 sg13g2_nand3_1 _07419_ (.B(_01420_),
    .C(_01421_),
    .A(_01401_),
    .Y(_01422_));
 sg13g2_a21o_1 _07420_ (.A2(_01421_),
    .A1(_01420_),
    .B1(_01401_),
    .X(_01423_));
 sg13g2_nand2_1 _07421_ (.Y(_01424_),
    .A(_01422_),
    .B(_01423_));
 sg13g2_xnor2_1 _07422_ (.Y(_01425_),
    .A(_01404_),
    .B(_01424_));
 sg13g2_o21ai_1 _07423_ (.B1(_01408_),
    .Y(_00152_),
    .A1(net2943),
    .A2(_01425_));
 sg13g2_nand2_1 _07424_ (.Y(_01426_),
    .A(net874),
    .B(net2941));
 sg13g2_nand2_1 _07425_ (.Y(_01427_),
    .A(_01417_),
    .B(_01420_));
 sg13g2_a22oi_1 _07426_ (.Y(_01428_),
    .B1(net3299),
    .B2(net3224),
    .A2(net3216),
    .A1(net3345));
 sg13g2_nand4_1 _07427_ (.B(net3224),
    .C(net3216),
    .A(net3345),
    .Y(_01429_),
    .D(net3299));
 sg13g2_nand2b_1 _07428_ (.Y(_01430_),
    .B(_01429_),
    .A_N(_01428_));
 sg13g2_o21ai_1 _07429_ (.B1(_01413_),
    .Y(_01431_),
    .A1(_01411_),
    .A2(_01414_));
 sg13g2_nand2_1 _07430_ (.Y(_01432_),
    .A(net3335),
    .B(net3217));
 sg13g2_and4_1 _07431_ (.A(net3221),
    .B(net3321),
    .C(net3219),
    .D(net3308),
    .X(_01433_));
 sg13g2_nand4_1 _07432_ (.B(net3321),
    .C(net3220),
    .A(net3221),
    .Y(_01434_),
    .D(net3308));
 sg13g2_a22oi_1 _07433_ (.Y(_01435_),
    .B1(net3308),
    .B2(net3221),
    .A2(net3219),
    .A1(net3321));
 sg13g2_or3_1 _07434_ (.A(_01432_),
    .B(_01433_),
    .C(_01435_),
    .X(_01436_));
 sg13g2_o21ai_1 _07435_ (.B1(_01432_),
    .Y(_01437_),
    .A1(_01433_),
    .A2(_01435_));
 sg13g2_and3_1 _07436_ (.X(_01438_),
    .A(_01431_),
    .B(_01436_),
    .C(_01437_));
 sg13g2_a21oi_1 _07437_ (.A1(_01436_),
    .A2(_01437_),
    .Y(_01439_),
    .B1(_01431_));
 sg13g2_o21ai_1 _07438_ (.B1(_01430_),
    .Y(_01440_),
    .A1(_01438_),
    .A2(_01439_));
 sg13g2_or3_1 _07439_ (.A(_01430_),
    .B(_01438_),
    .C(_01439_),
    .X(_01441_));
 sg13g2_and2_1 _07440_ (.A(_01440_),
    .B(_01441_),
    .X(_01442_));
 sg13g2_nand2_1 _07441_ (.Y(_01443_),
    .A(_01427_),
    .B(_01442_));
 sg13g2_xnor2_1 _07442_ (.Y(_01444_),
    .A(_01427_),
    .B(_01442_));
 sg13g2_nor2_1 _07443_ (.A(_01422_),
    .B(_01444_),
    .Y(_01445_));
 sg13g2_xnor2_1 _07444_ (.Y(_01446_),
    .A(_01422_),
    .B(_01444_));
 sg13g2_o21ai_1 _07445_ (.B1(_01446_),
    .Y(_01447_),
    .A1(_01404_),
    .A2(_01424_));
 sg13g2_or3_1 _07446_ (.A(_01404_),
    .B(_01424_),
    .C(_01444_),
    .X(_01448_));
 sg13g2_nand4_1 _07447_ (.B(net2978),
    .C(_01447_),
    .A(net3024),
    .Y(_01449_),
    .D(_01448_));
 sg13g2_nand2_1 _07448_ (.Y(_00153_),
    .A(_01426_),
    .B(_01449_));
 sg13g2_nand2_1 _07449_ (.Y(_01450_),
    .A(net955),
    .B(net2940));
 sg13g2_nand2b_1 _07450_ (.Y(_01451_),
    .B(_01441_),
    .A_N(_01438_));
 sg13g2_nand2_1 _07451_ (.Y(_01452_),
    .A(net3225),
    .B(net3294));
 sg13g2_and4_1 _07452_ (.A(net3345),
    .B(net3223),
    .C(net3299),
    .D(net3214),
    .X(_01453_));
 sg13g2_a22oi_1 _07453_ (.Y(_01454_),
    .B1(net3214),
    .B2(net3345),
    .A2(net3299),
    .A1(net3223));
 sg13g2_nor3_1 _07454_ (.A(_01452_),
    .B(_01453_),
    .C(_01454_),
    .Y(_01455_));
 sg13g2_o21ai_1 _07455_ (.B1(_01452_),
    .Y(_01456_),
    .A1(_01453_),
    .A2(_01454_));
 sg13g2_nand2b_1 _07456_ (.Y(_01457_),
    .B(_01456_),
    .A_N(_01455_));
 sg13g2_o21ai_1 _07457_ (.B1(_01434_),
    .Y(_01458_),
    .A1(_01432_),
    .A2(_01435_));
 sg13g2_nand2_1 _07458_ (.Y(_01459_),
    .A(net3335),
    .B(net3216));
 sg13g2_and4_1 _07459_ (.A(net3321),
    .B(net3219),
    .C(net3308),
    .D(net3217),
    .X(_01460_));
 sg13g2_nand4_1 _07460_ (.B(net3219),
    .C(net3308),
    .A(net3321),
    .Y(_01461_),
    .D(net3217));
 sg13g2_a22oi_1 _07461_ (.Y(_01462_),
    .B1(net3217),
    .B2(net3321),
    .A2(net3308),
    .A1(net3219));
 sg13g2_or3_1 _07462_ (.A(_01459_),
    .B(_01460_),
    .C(_01462_),
    .X(_01463_));
 sg13g2_o21ai_1 _07463_ (.B1(_01459_),
    .Y(_01464_),
    .A1(_01460_),
    .A2(_01462_));
 sg13g2_nand3_1 _07464_ (.B(_01463_),
    .C(_01464_),
    .A(_01458_),
    .Y(_01465_));
 sg13g2_a21oi_1 _07465_ (.A1(_01463_),
    .A2(_01464_),
    .Y(_01466_),
    .B1(_01458_));
 sg13g2_a21o_1 _07466_ (.A2(_01464_),
    .A1(_01463_),
    .B1(_01458_),
    .X(_01467_));
 sg13g2_nand2_1 _07467_ (.Y(_01468_),
    .A(_01465_),
    .B(_01467_));
 sg13g2_xnor2_1 _07468_ (.Y(_01469_),
    .A(_01457_),
    .B(_01468_));
 sg13g2_nand2b_1 _07469_ (.Y(_01470_),
    .B(_01451_),
    .A_N(_01469_));
 sg13g2_xor2_1 _07470_ (.B(_01469_),
    .A(_01451_),
    .X(_01471_));
 sg13g2_xor2_1 _07471_ (.B(_01471_),
    .A(_01429_),
    .X(_01472_));
 sg13g2_o21ai_1 _07472_ (.B1(_01443_),
    .Y(_01473_),
    .A1(_01422_),
    .A2(_01444_));
 sg13g2_xnor2_1 _07473_ (.Y(_01474_),
    .A(_01472_),
    .B(_01473_));
 sg13g2_nor2_1 _07474_ (.A(_01448_),
    .B(_01474_),
    .Y(_01475_));
 sg13g2_a21o_1 _07475_ (.A2(_01474_),
    .A1(_01448_),
    .B1(net2943),
    .X(_01476_));
 sg13g2_o21ai_1 _07476_ (.B1(_01450_),
    .Y(_00154_),
    .A1(_01475_),
    .A2(_01476_));
 sg13g2_nand2_1 _07477_ (.Y(_01477_),
    .A(net952),
    .B(net2940));
 sg13g2_nand2_1 _07478_ (.Y(_01478_),
    .A(_01445_),
    .B(_01472_));
 sg13g2_o21ai_1 _07479_ (.B1(_01478_),
    .Y(_01479_),
    .A1(_01448_),
    .A2(_01474_));
 sg13g2_nor2b_1 _07480_ (.A(_01443_),
    .B_N(_01472_),
    .Y(_01480_));
 sg13g2_o21ai_1 _07481_ (.B1(_01470_),
    .Y(_01481_),
    .A1(_01429_),
    .A2(_01471_));
 sg13g2_or2_1 _07482_ (.X(_01482_),
    .B(_01455_),
    .A(_01453_));
 sg13g2_nand2_1 _07483_ (.Y(_01483_),
    .A(net3225),
    .B(net3288));
 sg13g2_nand2b_1 _07484_ (.Y(_01484_),
    .B(_01482_),
    .A_N(_01483_));
 sg13g2_xor2_1 _07485_ (.B(_01483_),
    .A(_01482_),
    .X(_01485_));
 sg13g2_o21ai_1 _07486_ (.B1(_01465_),
    .Y(_01486_),
    .A1(_01457_),
    .A2(_01466_));
 sg13g2_nand2_1 _07487_ (.Y(_01487_),
    .A(net3223),
    .B(net3294));
 sg13g2_nand2_1 _07488_ (.Y(_01488_),
    .A(net3345),
    .B(net3211));
 sg13g2_nand2_1 _07489_ (.Y(_01489_),
    .A(net3219),
    .B(net3299));
 sg13g2_xor2_1 _07490_ (.B(_01489_),
    .A(_01488_),
    .X(_01490_));
 sg13g2_nand2b_1 _07491_ (.Y(_01491_),
    .B(_01490_),
    .A_N(_01487_));
 sg13g2_xnor2_1 _07492_ (.Y(_01492_),
    .A(_01487_),
    .B(_01490_));
 sg13g2_o21ai_1 _07493_ (.B1(_01461_),
    .Y(_01493_),
    .A1(_01459_),
    .A2(_01462_));
 sg13g2_nand2_1 _07494_ (.Y(_01494_),
    .A(net3335),
    .B(net3214));
 sg13g2_and4_1 _07495_ (.A(net3322),
    .B(net3308),
    .C(net3218),
    .D(net3216),
    .X(_01495_));
 sg13g2_nand4_1 _07496_ (.B(net3309),
    .C(net3218),
    .A(net3322),
    .Y(_01496_),
    .D(net3215));
 sg13g2_a22oi_1 _07497_ (.Y(_01497_),
    .B1(net3215),
    .B2(net3321),
    .A2(net3218),
    .A1(net3308));
 sg13g2_or3_1 _07498_ (.A(_01494_),
    .B(_01495_),
    .C(_01497_),
    .X(_01498_));
 sg13g2_o21ai_1 _07499_ (.B1(_01494_),
    .Y(_01499_),
    .A1(_01495_),
    .A2(_01497_));
 sg13g2_nand3_1 _07500_ (.B(_01498_),
    .C(_01499_),
    .A(_01493_),
    .Y(_01500_));
 sg13g2_a21o_1 _07501_ (.A2(_01499_),
    .A1(_01498_),
    .B1(_01493_),
    .X(_01501_));
 sg13g2_nand3_1 _07502_ (.B(_01500_),
    .C(_01501_),
    .A(_01492_),
    .Y(_01502_));
 sg13g2_a21o_1 _07503_ (.A2(_01501_),
    .A1(_01500_),
    .B1(_01492_),
    .X(_01503_));
 sg13g2_and3_1 _07504_ (.X(_01504_),
    .A(_01486_),
    .B(_01502_),
    .C(_01503_));
 sg13g2_a21oi_1 _07505_ (.A1(_01502_),
    .A2(_01503_),
    .Y(_01505_),
    .B1(_01486_));
 sg13g2_o21ai_1 _07506_ (.B1(_01485_),
    .Y(_01506_),
    .A1(_01504_),
    .A2(_01505_));
 sg13g2_or3_1 _07507_ (.A(_01485_),
    .B(_01504_),
    .C(_01505_),
    .X(_01507_));
 sg13g2_nand2_1 _07508_ (.Y(_01508_),
    .A(_01506_),
    .B(_01507_));
 sg13g2_nand2b_1 _07509_ (.Y(_01509_),
    .B(_01481_),
    .A_N(_01508_));
 sg13g2_xnor2_1 _07510_ (.Y(_01510_),
    .A(_01481_),
    .B(_01508_));
 sg13g2_and2_1 _07511_ (.A(_01480_),
    .B(_01510_),
    .X(_01511_));
 sg13g2_xor2_1 _07512_ (.B(_01510_),
    .A(_01480_),
    .X(_01512_));
 sg13g2_nor2_1 _07513_ (.A(_01479_),
    .B(_01512_),
    .Y(_01513_));
 sg13g2_a21o_1 _07514_ (.A2(_01512_),
    .A1(_01479_),
    .B1(net2943),
    .X(_01514_));
 sg13g2_o21ai_1 _07515_ (.B1(_01477_),
    .Y(_00155_),
    .A1(_01513_),
    .A2(_01514_));
 sg13g2_a21o_1 _07516_ (.A2(_01512_),
    .A1(_01479_),
    .B1(_01511_),
    .X(_01515_));
 sg13g2_nand2b_1 _07517_ (.Y(_01516_),
    .B(_01507_),
    .A_N(_01504_));
 sg13g2_o21ai_1 _07518_ (.B1(_01491_),
    .Y(_01517_),
    .A1(_01488_),
    .A2(_01489_));
 sg13g2_nor2_1 _07519_ (.A(net3225),
    .B(net3279),
    .Y(_01518_));
 sg13g2_nand2_1 _07520_ (.Y(_01519_),
    .A(net3220),
    .B(net3292));
 sg13g2_nor2_1 _07521_ (.A(_01487_),
    .B(_01519_),
    .Y(_01520_));
 sg13g2_a22oi_1 _07522_ (.Y(_01521_),
    .B1(net3292),
    .B2(net3223),
    .A2(net3294),
    .A1(net3219));
 sg13g2_nor2_1 _07523_ (.A(_01520_),
    .B(_01521_),
    .Y(_01522_));
 sg13g2_xor2_1 _07524_ (.B(_01522_),
    .A(_01518_),
    .X(_01523_));
 sg13g2_nand2_1 _07525_ (.Y(_01524_),
    .A(_01517_),
    .B(_01523_));
 sg13g2_xnor2_1 _07526_ (.Y(_01525_),
    .A(_01517_),
    .B(_01523_));
 sg13g2_nand2_1 _07527_ (.Y(_01526_),
    .A(_01500_),
    .B(_01502_));
 sg13g2_nand2_1 _07528_ (.Y(_01527_),
    .A(net3218),
    .B(net3299));
 sg13g2_and2_1 _07529_ (.A(net3335),
    .B(net3205),
    .X(_01528_));
 sg13g2_nand2_2 _07530_ (.Y(_01529_),
    .A(net3337),
    .B(net3205));
 sg13g2_and4_1 _07531_ (.A(net3346),
    .B(net3335),
    .C(net3211),
    .D(net3208),
    .X(_01530_));
 sg13g2_a22oi_1 _07532_ (.Y(_01531_),
    .B1(net3208),
    .B2(net3346),
    .A2(net3211),
    .A1(net3335));
 sg13g2_nor3_1 _07533_ (.A(_01527_),
    .B(_01530_),
    .C(_01531_),
    .Y(_01532_));
 sg13g2_o21ai_1 _07534_ (.B1(_01527_),
    .Y(_01533_),
    .A1(_01530_),
    .A2(_01531_));
 sg13g2_nor2b_1 _07535_ (.A(_01532_),
    .B_N(_01533_),
    .Y(_01534_));
 sg13g2_o21ai_1 _07536_ (.B1(_01496_),
    .Y(_01535_),
    .A1(_01494_),
    .A2(_01497_));
 sg13g2_nand2_1 _07537_ (.Y(_01536_),
    .A(net3323),
    .B(net3213));
 sg13g2_and3_1 _07538_ (.X(_01537_),
    .A(net3309),
    .B(net3215),
    .C(net3285));
 sg13g2_nand3_1 _07539_ (.B(net3215),
    .C(net3285),
    .A(net3309),
    .Y(_01538_));
 sg13g2_a21oi_1 _07540_ (.A1(net3309),
    .A2(net3215),
    .Y(_01539_),
    .B1(net3285));
 sg13g2_or3_1 _07541_ (.A(_01536_),
    .B(_01537_),
    .C(_01539_),
    .X(_01540_));
 sg13g2_o21ai_1 _07542_ (.B1(_01536_),
    .Y(_01541_),
    .A1(_01537_),
    .A2(_01539_));
 sg13g2_nand3_1 _07543_ (.B(_01540_),
    .C(_01541_),
    .A(_01535_),
    .Y(_01542_));
 sg13g2_a21o_1 _07544_ (.A2(_01541_),
    .A1(_01540_),
    .B1(_01535_),
    .X(_01543_));
 sg13g2_nand3_1 _07545_ (.B(_01542_),
    .C(_01543_),
    .A(_01534_),
    .Y(_01544_));
 sg13g2_a21o_1 _07546_ (.A2(_01543_),
    .A1(_01542_),
    .B1(_01534_),
    .X(_01545_));
 sg13g2_nand2_1 _07547_ (.Y(_01546_),
    .A(_01544_),
    .B(_01545_));
 sg13g2_nand2b_1 _07548_ (.Y(_01547_),
    .B(_01526_),
    .A_N(_01546_));
 sg13g2_nor2b_1 _07549_ (.A(_01526_),
    .B_N(_01546_),
    .Y(_01548_));
 sg13g2_xnor2_1 _07550_ (.Y(_01549_),
    .A(_01526_),
    .B(_01546_));
 sg13g2_xnor2_1 _07551_ (.Y(_01550_),
    .A(_01525_),
    .B(_01549_));
 sg13g2_nand2_1 _07552_ (.Y(_01551_),
    .A(_01516_),
    .B(_01550_));
 sg13g2_xnor2_1 _07553_ (.Y(_01552_),
    .A(_01516_),
    .B(_01550_));
 sg13g2_xor2_1 _07554_ (.B(_01552_),
    .A(_01484_),
    .X(_01553_));
 sg13g2_nor2b_1 _07555_ (.A(_01509_),
    .B_N(_01553_),
    .Y(_01554_));
 sg13g2_xnor2_1 _07556_ (.Y(_01555_),
    .A(_01509_),
    .B(_01553_));
 sg13g2_nand2_1 _07557_ (.Y(_01556_),
    .A(_01515_),
    .B(_01555_));
 sg13g2_nor2_1 _07558_ (.A(_01515_),
    .B(_01555_),
    .Y(_01557_));
 sg13g2_nor2_1 _07559_ (.A(net2943),
    .B(_01557_),
    .Y(_01558_));
 sg13g2_a22oi_1 _07560_ (.Y(_01559_),
    .B1(_01556_),
    .B2(_01558_),
    .A2(net2940),
    .A1(net988));
 sg13g2_inv_1 _07561_ (.Y(_00156_),
    .A(_01559_));
 sg13g2_o21ai_1 _07562_ (.B1(_01547_),
    .Y(_01560_),
    .A1(_01525_),
    .A2(_01548_));
 sg13g2_a21oi_1 _07563_ (.A1(_01518_),
    .A2(_01522_),
    .Y(_01561_),
    .B1(_01520_));
 sg13g2_or2_1 _07564_ (.X(_01562_),
    .B(_01532_),
    .A(_01530_));
 sg13g2_nor2_1 _07565_ (.A(net3223),
    .B(net3279),
    .Y(_01563_));
 sg13g2_nor3_1 _07566_ (.A(net3222),
    .B(net3279),
    .C(_01519_),
    .Y(_01564_));
 sg13g2_inv_1 _07567_ (.Y(_01565_),
    .A(_01564_));
 sg13g2_xnor2_1 _07568_ (.Y(_01566_),
    .A(_01519_),
    .B(_01563_));
 sg13g2_xnor2_1 _07569_ (.Y(_01567_),
    .A(_01562_),
    .B(_01566_));
 sg13g2_nor2_1 _07570_ (.A(_01561_),
    .B(_01567_),
    .Y(_01568_));
 sg13g2_xnor2_1 _07571_ (.Y(_01569_),
    .A(_01561_),
    .B(_01567_));
 sg13g2_nand2_1 _07572_ (.Y(_01570_),
    .A(_01542_),
    .B(_01544_));
 sg13g2_nand2_1 _07573_ (.Y(_01571_),
    .A(net3217),
    .B(net3294));
 sg13g2_and3_1 _07574_ (.X(_01572_),
    .A(net3),
    .B(net3300),
    .C(net3205));
 sg13g2_nand2_1 _07575_ (.Y(_01573_),
    .A(net3216),
    .B(net2975));
 sg13g2_a22oi_1 _07576_ (.Y(_01574_),
    .B1(net3208),
    .B2(net3347),
    .A2(net3299),
    .A1(net3215));
 sg13g2_a21oi_1 _07577_ (.A1(net3215),
    .A2(net2975),
    .Y(_01575_),
    .B1(_01574_));
 sg13g2_xor2_1 _07578_ (.B(_01575_),
    .A(_01571_),
    .X(_01576_));
 sg13g2_o21ai_1 _07579_ (.B1(_01538_),
    .Y(_01577_),
    .A1(_01536_),
    .A2(_01539_));
 sg13g2_and4_1 _07580_ (.A(net3323),
    .B(net3309),
    .C(net3213),
    .D(net3211),
    .X(_01578_));
 sg13g2_nand4_1 _07581_ (.B(net3309),
    .C(net3212),
    .A(net3323),
    .Y(_01579_),
    .D(net3209));
 sg13g2_a22oi_1 _07582_ (.Y(_01580_),
    .B1(net3209),
    .B2(net3323),
    .A2(net3212),
    .A1(net3309));
 sg13g2_nand3b_1 _07583_ (.B(_01528_),
    .C(_01579_),
    .Y(_01581_),
    .A_N(_01580_));
 sg13g2_o21ai_1 _07584_ (.B1(_01529_),
    .Y(_01582_),
    .A1(_01578_),
    .A2(_01580_));
 sg13g2_nand3_1 _07585_ (.B(_01581_),
    .C(_01582_),
    .A(_01577_),
    .Y(_01583_));
 sg13g2_a21oi_1 _07586_ (.A1(_01581_),
    .A2(_01582_),
    .Y(_01584_),
    .B1(_01577_));
 sg13g2_a21o_1 _07587_ (.A2(_01582_),
    .A1(_01581_),
    .B1(_01577_),
    .X(_01585_));
 sg13g2_nand2_1 _07588_ (.Y(_01586_),
    .A(_01583_),
    .B(_01585_));
 sg13g2_xnor2_1 _07589_ (.Y(_01587_),
    .A(_01576_),
    .B(_01586_));
 sg13g2_nand2b_1 _07590_ (.Y(_01588_),
    .B(_01570_),
    .A_N(_01587_));
 sg13g2_xor2_1 _07591_ (.B(_01587_),
    .A(_01570_),
    .X(_01589_));
 sg13g2_xor2_1 _07592_ (.B(_01589_),
    .A(_01569_),
    .X(_01590_));
 sg13g2_nand2_1 _07593_ (.Y(_01591_),
    .A(_01560_),
    .B(_01590_));
 sg13g2_xnor2_1 _07594_ (.Y(_01592_),
    .A(_01560_),
    .B(_01590_));
 sg13g2_xor2_1 _07595_ (.B(_01592_),
    .A(_01524_),
    .X(_01593_));
 sg13g2_o21ai_1 _07596_ (.B1(_01551_),
    .Y(_01594_),
    .A1(_01484_),
    .A2(_01552_));
 sg13g2_nand2_2 _07597_ (.Y(_01595_),
    .A(_01593_),
    .B(_01594_));
 sg13g2_xnor2_1 _07598_ (.Y(_01596_),
    .A(_01593_),
    .B(_01594_));
 sg13g2_a21oi_1 _07599_ (.A1(_01515_),
    .A2(_01555_),
    .Y(_01597_),
    .B1(_01554_));
 sg13g2_or2_2 _07600_ (.X(_01598_),
    .B(_01597_),
    .A(_01596_));
 sg13g2_a21oi_1 _07601_ (.A1(_01596_),
    .A2(_01597_),
    .Y(_01599_),
    .B1(net2942));
 sg13g2_a22oi_1 _07602_ (.Y(_01600_),
    .B1(_01598_),
    .B2(_01599_),
    .A2(net2940),
    .A1(net1008));
 sg13g2_inv_1 _07603_ (.Y(_00157_),
    .A(_01600_));
 sg13g2_o21ai_1 _07604_ (.B1(_01591_),
    .Y(_01601_),
    .A1(_01524_),
    .A2(_01592_));
 sg13g2_a21oi_1 _07605_ (.A1(_01562_),
    .A2(_01566_),
    .Y(_01602_),
    .B1(_01568_));
 sg13g2_o21ai_1 _07606_ (.B1(_01588_),
    .Y(_01603_),
    .A1(_01569_),
    .A2(_01589_));
 sg13g2_o21ai_1 _07607_ (.B1(_01573_),
    .Y(_01604_),
    .A1(_01571_),
    .A2(_01574_));
 sg13g2_nand2_1 _07608_ (.Y(_01605_),
    .A(net3218),
    .B(net3288));
 sg13g2_nor2_1 _07609_ (.A(net3220),
    .B(net3279),
    .Y(_01606_));
 sg13g2_nand2b_1 _07610_ (.Y(_01607_),
    .B(_01606_),
    .A_N(_01605_));
 sg13g2_xnor2_1 _07611_ (.Y(_01608_),
    .A(_01605_),
    .B(_01606_));
 sg13g2_nand2_1 _07612_ (.Y(_01609_),
    .A(_01604_),
    .B(_01608_));
 sg13g2_xnor2_1 _07613_ (.Y(_01610_),
    .A(_01604_),
    .B(_01608_));
 sg13g2_xnor2_1 _07614_ (.Y(_01611_),
    .A(_01565_),
    .B(_01610_));
 sg13g2_o21ai_1 _07615_ (.B1(_01583_),
    .Y(_01612_),
    .A1(_01576_),
    .A2(_01584_));
 sg13g2_nand2_1 _07616_ (.Y(_01613_),
    .A(net3216),
    .B(net3294));
 sg13g2_nand2_1 _07617_ (.Y(_01614_),
    .A(net3213),
    .B(net2975));
 sg13g2_a22oi_1 _07618_ (.Y(_01615_),
    .B1(net3207),
    .B2(net3346),
    .A2(net3212),
    .A1(net3299));
 sg13g2_a21oi_1 _07619_ (.A1(net3212),
    .A2(net2975),
    .Y(_01616_),
    .B1(_01615_));
 sg13g2_xor2_1 _07620_ (.B(_01616_),
    .A(_01613_),
    .X(_01617_));
 sg13g2_o21ai_1 _07621_ (.B1(_01579_),
    .Y(_01618_),
    .A1(_01529_),
    .A2(_01580_));
 sg13g2_and4_1 _07622_ (.A(net3323),
    .B(net3311),
    .C(net3209),
    .D(net3205),
    .X(_01619_));
 sg13g2_nand4_1 _07623_ (.B(net3311),
    .C(net3209),
    .A(net3326),
    .Y(_01620_),
    .D(net3205));
 sg13g2_a22oi_1 _07624_ (.Y(_01621_),
    .B1(net3205),
    .B2(net3326),
    .A2(net3209),
    .A1(net3311));
 sg13g2_nand3b_1 _07625_ (.B(_01528_),
    .C(_01620_),
    .Y(_01622_),
    .A_N(_01621_));
 sg13g2_o21ai_1 _07626_ (.B1(_01529_),
    .Y(_01623_),
    .A1(_01619_),
    .A2(_01621_));
 sg13g2_and3_1 _07627_ (.X(_01624_),
    .A(_01618_),
    .B(_01622_),
    .C(_01623_));
 sg13g2_nand3_1 _07628_ (.B(_01622_),
    .C(_01623_),
    .A(_01618_),
    .Y(_01625_));
 sg13g2_a21oi_1 _07629_ (.A1(_01622_),
    .A2(_01623_),
    .Y(_01626_),
    .B1(_01618_));
 sg13g2_or3_1 _07630_ (.A(_01617_),
    .B(_01624_),
    .C(_01626_),
    .X(_01627_));
 sg13g2_o21ai_1 _07631_ (.B1(_01617_),
    .Y(_01628_),
    .A1(_01624_),
    .A2(_01626_));
 sg13g2_and3_1 _07632_ (.X(_01629_),
    .A(_01612_),
    .B(_01627_),
    .C(_01628_));
 sg13g2_nand3_1 _07633_ (.B(_01627_),
    .C(_01628_),
    .A(_01612_),
    .Y(_01630_));
 sg13g2_a21oi_1 _07634_ (.A1(_01627_),
    .A2(_01628_),
    .Y(_01631_),
    .B1(_01612_));
 sg13g2_nor2_1 _07635_ (.A(_01629_),
    .B(_01631_),
    .Y(_01632_));
 sg13g2_xor2_1 _07636_ (.B(_01632_),
    .A(_01611_),
    .X(_01633_));
 sg13g2_nand2b_1 _07637_ (.Y(_01634_),
    .B(_01603_),
    .A_N(_01633_));
 sg13g2_xor2_1 _07638_ (.B(_01633_),
    .A(_01603_),
    .X(_01635_));
 sg13g2_xor2_1 _07639_ (.B(_01635_),
    .A(_01602_),
    .X(_01636_));
 sg13g2_nand2_1 _07640_ (.Y(_01637_),
    .A(_01601_),
    .B(_01636_));
 sg13g2_nor2_1 _07641_ (.A(_01601_),
    .B(_01636_),
    .Y(_01638_));
 sg13g2_xnor2_1 _07642_ (.Y(_01639_),
    .A(_01601_),
    .B(_01636_));
 sg13g2_a21oi_1 _07643_ (.A1(_01595_),
    .A2(_01598_),
    .Y(_01640_),
    .B1(_01639_));
 sg13g2_nand3_1 _07644_ (.B(_01598_),
    .C(_01639_),
    .A(_01595_),
    .Y(_01641_));
 sg13g2_nor2_1 _07645_ (.A(net2942),
    .B(_01640_),
    .Y(_01642_));
 sg13g2_a22oi_1 _07646_ (.Y(_01643_),
    .B1(_01641_),
    .B2(_01642_),
    .A2(net2940),
    .A1(net1017));
 sg13g2_inv_1 _07647_ (.Y(_00158_),
    .A(_01643_));
 sg13g2_and2_1 _07648_ (.A(net1078),
    .B(net2940),
    .X(_01644_));
 sg13g2_o21ai_1 _07649_ (.B1(_01609_),
    .Y(_01645_),
    .A1(_01565_),
    .A2(_01610_));
 sg13g2_o21ai_1 _07650_ (.B1(_01630_),
    .Y(_01646_),
    .A1(_01611_),
    .A2(_01631_));
 sg13g2_o21ai_1 _07651_ (.B1(_01614_),
    .Y(_01647_),
    .A1(_01613_),
    .A2(_01615_));
 sg13g2_nand2_2 _07652_ (.Y(_01648_),
    .A(\u_toplayer.u_outlayer.u_neuron.din[4] ),
    .B(net3288));
 sg13g2_nor2_1 _07653_ (.A(net3218),
    .B(net3279),
    .Y(_01649_));
 sg13g2_nand2b_1 _07654_ (.Y(_01650_),
    .B(_01649_),
    .A_N(_01648_));
 sg13g2_xnor2_1 _07655_ (.Y(_01651_),
    .A(_01648_),
    .B(_01649_));
 sg13g2_nand2_1 _07656_ (.Y(_01652_),
    .A(_01647_),
    .B(_01651_));
 sg13g2_xnor2_1 _07657_ (.Y(_01653_),
    .A(_01647_),
    .B(_01651_));
 sg13g2_xnor2_1 _07658_ (.Y(_01654_),
    .A(_01607_),
    .B(_01653_));
 sg13g2_o21ai_1 _07659_ (.B1(_01625_),
    .Y(_01655_),
    .A1(_01617_),
    .A2(_01626_));
 sg13g2_and2_1 _07660_ (.A(net3212),
    .B(net3294),
    .X(_01656_));
 sg13g2_a22oi_1 _07661_ (.Y(_01657_),
    .B1(net3207),
    .B2(net3346),
    .A2(net3210),
    .A1(net3300));
 sg13g2_a21oi_1 _07662_ (.A1(net3210),
    .A2(_01572_),
    .Y(_01658_),
    .B1(_01657_));
 sg13g2_xor2_1 _07663_ (.B(_01658_),
    .A(_01656_),
    .X(_01659_));
 sg13g2_o21ai_1 _07664_ (.B1(_01620_),
    .Y(_01660_),
    .A1(_01529_),
    .A2(_01621_));
 sg13g2_xor2_1 _07665_ (.B(net3312),
    .A(net3326),
    .X(_01661_));
 sg13g2_nand2b_1 _07666_ (.Y(_01662_),
    .B(net3205),
    .A_N(net3336));
 sg13g2_mux2_1 _07667_ (.A0(_01529_),
    .A1(_01662_),
    .S(_01661_),
    .X(_01663_));
 sg13g2_a21oi_2 _07668_ (.B1(_01663_),
    .Y(_01664_),
    .A2(_01622_),
    .A1(_01620_));
 sg13g2_xnor2_1 _07669_ (.Y(_01665_),
    .A(_01660_),
    .B(_01663_));
 sg13g2_xnor2_1 _07670_ (.Y(_01666_),
    .A(_01659_),
    .B(_01665_));
 sg13g2_nand2b_1 _07671_ (.Y(_01667_),
    .B(_01655_),
    .A_N(_01666_));
 sg13g2_xor2_1 _07672_ (.B(_01666_),
    .A(_01655_),
    .X(_01668_));
 sg13g2_xor2_1 _07673_ (.B(_01668_),
    .A(_01654_),
    .X(_01669_));
 sg13g2_xnor2_1 _07674_ (.Y(_01670_),
    .A(_01646_),
    .B(_01669_));
 sg13g2_nor2b_1 _07675_ (.A(_01670_),
    .B_N(_01645_),
    .Y(_01671_));
 sg13g2_xor2_1 _07676_ (.B(_01670_),
    .A(_01645_),
    .X(_01672_));
 sg13g2_o21ai_1 _07677_ (.B1(_01634_),
    .Y(_01673_),
    .A1(_01602_),
    .A2(_01635_));
 sg13g2_nor2b_1 _07678_ (.A(_01672_),
    .B_N(_01673_),
    .Y(_01674_));
 sg13g2_xor2_1 _07679_ (.B(_01673_),
    .A(_01672_),
    .X(_01675_));
 sg13g2_inv_1 _07680_ (.Y(_01676_),
    .A(_01675_));
 sg13g2_nor3_1 _07681_ (.A(_01596_),
    .B(_01597_),
    .C(_01639_),
    .Y(_01677_));
 sg13g2_o21ai_1 _07682_ (.B1(_01637_),
    .Y(_01678_),
    .A1(_01595_),
    .A2(_01638_));
 sg13g2_o21ai_1 _07683_ (.B1(_01676_),
    .Y(_01679_),
    .A1(_01677_),
    .A2(_01678_));
 sg13g2_nor3_1 _07684_ (.A(_01676_),
    .B(_01677_),
    .C(_01678_),
    .Y(_01680_));
 sg13g2_nor2_1 _07685_ (.A(net2942),
    .B(_01680_),
    .Y(_01681_));
 sg13g2_a21o_1 _07686_ (.A2(_01681_),
    .A1(_01679_),
    .B1(_01644_),
    .X(_00159_));
 sg13g2_nand2_1 _07687_ (.Y(_01682_),
    .A(net833),
    .B(net2940));
 sg13g2_nor2b_1 _07688_ (.A(_01674_),
    .B_N(_01679_),
    .Y(_01683_));
 sg13g2_a21o_1 _07689_ (.A2(_01669_),
    .A1(_01646_),
    .B1(_01671_),
    .X(_01684_));
 sg13g2_o21ai_1 _07690_ (.B1(_01652_),
    .Y(_01685_),
    .A1(_01607_),
    .A2(_01653_));
 sg13g2_o21ai_1 _07691_ (.B1(_01667_),
    .Y(_01686_),
    .A1(_01654_),
    .A2(_01668_));
 sg13g2_a22oi_1 _07692_ (.Y(_01687_),
    .B1(_01656_),
    .B2(_01658_),
    .A2(net2975),
    .A1(net3210));
 sg13g2_nand2_1 _07693_ (.Y(_01688_),
    .A(net3212),
    .B(net3288));
 sg13g2_nor2_1 _07694_ (.A(net3215),
    .B(net3280),
    .Y(_01689_));
 sg13g2_nand2b_1 _07695_ (.Y(_01690_),
    .B(_01689_),
    .A_N(_01688_));
 sg13g2_xnor2_1 _07696_ (.Y(_01691_),
    .A(_01688_),
    .B(_01689_));
 sg13g2_nand2b_1 _07697_ (.Y(_01692_),
    .B(_01691_),
    .A_N(_01687_));
 sg13g2_xor2_1 _07698_ (.B(_01691_),
    .A(_01687_),
    .X(_01693_));
 sg13g2_xnor2_1 _07699_ (.Y(_01694_),
    .A(_01650_),
    .B(_01693_));
 sg13g2_a21oi_2 _07700_ (.B1(_01664_),
    .Y(_01695_),
    .A2(_01665_),
    .A1(_01659_));
 sg13g2_o21ai_1 _07701_ (.B1(net3206),
    .Y(_01696_),
    .A1(net3347),
    .A2(net3300));
 sg13g2_nor2_2 _07702_ (.A(_01572_),
    .B(_01696_),
    .Y(_01697_));
 sg13g2_nand2_1 _07703_ (.Y(_01698_),
    .A(net3295),
    .B(net3209));
 sg13g2_nor3_1 _07704_ (.A(net2975),
    .B(_01696_),
    .C(_01698_),
    .Y(_01699_));
 sg13g2_xor2_1 _07705_ (.B(_01698_),
    .A(_01697_),
    .X(_01700_));
 sg13g2_o21ai_1 _07706_ (.B1(net3205),
    .Y(_01701_),
    .A1(net3326),
    .A2(net3312));
 sg13g2_a21oi_2 _07707_ (.B1(_01664_),
    .Y(_01702_),
    .A2(_01701_),
    .A1(_01529_));
 sg13g2_nand2b_1 _07708_ (.Y(_01703_),
    .B(_01702_),
    .A_N(_01700_));
 sg13g2_xnor2_1 _07709_ (.Y(_01704_),
    .A(_01700_),
    .B(_01702_));
 sg13g2_inv_1 _07710_ (.Y(_01705_),
    .A(_01704_));
 sg13g2_xnor2_1 _07711_ (.Y(_01706_),
    .A(_01695_),
    .B(_01704_));
 sg13g2_nand2b_1 _07712_ (.Y(_01707_),
    .B(_01706_),
    .A_N(_01694_));
 sg13g2_xnor2_1 _07713_ (.Y(_01708_),
    .A(_01694_),
    .B(_01706_));
 sg13g2_xnor2_1 _07714_ (.Y(_01709_),
    .A(_01686_),
    .B(_01708_));
 sg13g2_nor2b_1 _07715_ (.A(_01709_),
    .B_N(_01685_),
    .Y(_01710_));
 sg13g2_xnor2_1 _07716_ (.Y(_01711_),
    .A(_01685_),
    .B(_01709_));
 sg13g2_nor2_1 _07717_ (.A(_01684_),
    .B(_01711_),
    .Y(_01712_));
 sg13g2_xnor2_1 _07718_ (.Y(_01713_),
    .A(_01684_),
    .B(_01711_));
 sg13g2_a21oi_1 _07719_ (.A1(_01683_),
    .A2(_01713_),
    .Y(_01714_),
    .B1(net2943));
 sg13g2_o21ai_1 _07720_ (.B1(_01714_),
    .Y(_01715_),
    .A1(_01683_),
    .A2(_01713_));
 sg13g2_nand2_1 _07721_ (.Y(_00160_),
    .A(_01682_),
    .B(_01715_));
 sg13g2_o21ai_1 _07722_ (.B1(_01692_),
    .Y(_01716_),
    .A1(_01650_),
    .A2(_01693_));
 sg13g2_o21ai_1 _07723_ (.B1(_01707_),
    .Y(_01717_),
    .A1(_01695_),
    .A2(_01705_));
 sg13g2_nand2b_1 _07724_ (.Y(_01718_),
    .B(_01703_),
    .A_N(_01664_));
 sg13g2_and2_1 _07725_ (.A(net3294),
    .B(net3206),
    .X(_01719_));
 sg13g2_xor2_1 _07726_ (.B(_01719_),
    .A(_01697_),
    .X(_01720_));
 sg13g2_xnor2_1 _07727_ (.Y(_01721_),
    .A(_01702_),
    .B(_01720_));
 sg13g2_inv_1 _07728_ (.Y(_01722_),
    .A(_01721_));
 sg13g2_xnor2_1 _07729_ (.Y(_01723_),
    .A(_01718_),
    .B(_01722_));
 sg13g2_nor2_1 _07730_ (.A(net2975),
    .B(_01699_),
    .Y(_01724_));
 sg13g2_nand2_1 _07731_ (.Y(_01725_),
    .A(net3209),
    .B(net3288));
 sg13g2_nor2_1 _07732_ (.A(net3212),
    .B(net3279),
    .Y(_01726_));
 sg13g2_nor3_2 _07733_ (.A(net3212),
    .B(net3280),
    .C(_01725_),
    .Y(_01727_));
 sg13g2_xnor2_1 _07734_ (.Y(_01728_),
    .A(_01725_),
    .B(_01726_));
 sg13g2_nand2b_1 _07735_ (.Y(_01729_),
    .B(_01728_),
    .A_N(_01724_));
 sg13g2_xor2_1 _07736_ (.B(_01728_),
    .A(_01724_),
    .X(_01730_));
 sg13g2_xnor2_1 _07737_ (.Y(_01731_),
    .A(_01690_),
    .B(_01730_));
 sg13g2_nor2_1 _07738_ (.A(_01723_),
    .B(_01731_),
    .Y(_01732_));
 sg13g2_xor2_1 _07739_ (.B(_01731_),
    .A(_01723_),
    .X(_01733_));
 sg13g2_xnor2_1 _07740_ (.Y(_01734_),
    .A(_01717_),
    .B(_01733_));
 sg13g2_nor2b_1 _07741_ (.A(_01734_),
    .B_N(_01716_),
    .Y(_01735_));
 sg13g2_xor2_1 _07742_ (.B(_01734_),
    .A(_01716_),
    .X(_01736_));
 sg13g2_a21o_1 _07743_ (.A2(_01708_),
    .A1(_01686_),
    .B1(_01710_),
    .X(_01737_));
 sg13g2_nand2b_1 _07744_ (.Y(_01738_),
    .B(_01737_),
    .A_N(_01736_));
 sg13g2_xor2_1 _07745_ (.B(_01737_),
    .A(_01736_),
    .X(_01739_));
 sg13g2_nor2_1 _07746_ (.A(_01675_),
    .B(_01713_),
    .Y(_01740_));
 sg13g2_nor2b_1 _07747_ (.A(_01712_),
    .B_N(_01674_),
    .Y(_01741_));
 sg13g2_a221oi_1 _07748_ (.B2(_01678_),
    .C1(_01741_),
    .B1(_01740_),
    .A1(_01684_),
    .Y(_01742_),
    .A2(_01711_));
 sg13g2_nand2b_1 _07749_ (.Y(_01743_),
    .B(_01740_),
    .A_N(_01639_));
 sg13g2_o21ai_1 _07750_ (.B1(_01742_),
    .Y(_01744_),
    .A1(_01598_),
    .A2(_01743_));
 sg13g2_nand2b_2 _07751_ (.Y(_01745_),
    .B(_01744_),
    .A_N(_01739_));
 sg13g2_nor2b_1 _07752_ (.A(_01744_),
    .B_N(_01739_),
    .Y(_01746_));
 sg13g2_nor2_1 _07753_ (.A(net2944),
    .B(_01746_),
    .Y(_01747_));
 sg13g2_a22oi_1 _07754_ (.Y(_01748_),
    .B1(_01745_),
    .B2(_01747_),
    .A2(net2941),
    .A1(net1060));
 sg13g2_inv_1 _07755_ (.Y(_00161_),
    .A(_01748_));
 sg13g2_and2_1 _07756_ (.A(net1199),
    .B(net2941),
    .X(_01749_));
 sg13g2_o21ai_1 _07757_ (.B1(_01729_),
    .Y(_01750_),
    .A1(_01690_),
    .A2(_01730_));
 sg13g2_a21oi_1 _07758_ (.A1(_01718_),
    .A2(_01722_),
    .Y(_01751_),
    .B1(_01732_));
 sg13g2_nand2_1 _07759_ (.Y(_01752_),
    .A(_01664_),
    .B(_01720_));
 sg13g2_or3_1 _07760_ (.A(_01664_),
    .B(_01702_),
    .C(_01720_),
    .X(_01753_));
 sg13g2_nand2_2 _07761_ (.Y(_01754_),
    .A(_01752_),
    .B(_01753_));
 sg13g2_a21oi_2 _07762_ (.B1(net2975),
    .Y(_01755_),
    .A2(_01719_),
    .A1(_01697_));
 sg13g2_nand2_1 _07763_ (.Y(_01756_),
    .A(net3288),
    .B(net3206));
 sg13g2_nor2_1 _07764_ (.A(net3209),
    .B(net3279),
    .Y(_01757_));
 sg13g2_nand2b_1 _07765_ (.Y(_01758_),
    .B(_01757_),
    .A_N(_01756_));
 sg13g2_xnor2_1 _07766_ (.Y(_01759_),
    .A(_01756_),
    .B(_01757_));
 sg13g2_nand2b_1 _07767_ (.Y(_01760_),
    .B(_01759_),
    .A_N(_01755_));
 sg13g2_xor2_1 _07768_ (.B(_01759_),
    .A(_01755_),
    .X(_01761_));
 sg13g2_inv_1 _07769_ (.Y(_01762_),
    .A(_01761_));
 sg13g2_nand2_1 _07770_ (.Y(_01763_),
    .A(_01727_),
    .B(_01762_));
 sg13g2_xor2_1 _07771_ (.B(_01761_),
    .A(_01727_),
    .X(_01764_));
 sg13g2_nor2_1 _07772_ (.A(_01754_),
    .B(_01764_),
    .Y(_01765_));
 sg13g2_xor2_1 _07773_ (.B(_01764_),
    .A(_01754_),
    .X(_01766_));
 sg13g2_nor2b_1 _07774_ (.A(_01751_),
    .B_N(_01766_),
    .Y(_01767_));
 sg13g2_xnor2_1 _07775_ (.Y(_01768_),
    .A(_01751_),
    .B(_01766_));
 sg13g2_xnor2_1 _07776_ (.Y(_01769_),
    .A(_01750_),
    .B(_01768_));
 sg13g2_a21oi_1 _07777_ (.A1(_01717_),
    .A2(_01733_),
    .Y(_01770_),
    .B1(_01735_));
 sg13g2_nor2_1 _07778_ (.A(_01769_),
    .B(_01770_),
    .Y(_01771_));
 sg13g2_xnor2_1 _07779_ (.Y(_01772_),
    .A(_01769_),
    .B(_01770_));
 sg13g2_nor2_1 _07780_ (.A(_01745_),
    .B(_01772_),
    .Y(_01773_));
 sg13g2_nand3_1 _07781_ (.B(_01745_),
    .C(_01772_),
    .A(_01738_),
    .Y(_01774_));
 sg13g2_nor2_1 _07782_ (.A(_01738_),
    .B(_01772_),
    .Y(_01775_));
 sg13g2_nor3_1 _07783_ (.A(net2944),
    .B(_01773_),
    .C(_01775_),
    .Y(_01776_));
 sg13g2_a21o_1 _07784_ (.A2(_01776_),
    .A1(_01774_),
    .B1(_01749_),
    .X(_00162_));
 sg13g2_and2_1 _07785_ (.A(net1200),
    .B(net2941),
    .X(_01777_));
 sg13g2_nor2_1 _07786_ (.A(_01771_),
    .B(_01775_),
    .Y(_01778_));
 sg13g2_o21ai_1 _07787_ (.B1(_01778_),
    .Y(_01779_),
    .A1(_01745_),
    .A2(_01772_));
 sg13g2_nand2_1 _07788_ (.Y(_01780_),
    .A(_01760_),
    .B(_01763_));
 sg13g2_a21oi_1 _07789_ (.A1(_01664_),
    .A2(_01720_),
    .Y(_01781_),
    .B1(_01765_));
 sg13g2_o21ai_1 _07790_ (.B1(_01756_),
    .Y(_01782_),
    .A1(net3279),
    .A2(net3206));
 sg13g2_nand2b_1 _07791_ (.Y(_01783_),
    .B(_01782_),
    .A_N(_01755_));
 sg13g2_nand2_1 _07792_ (.Y(_01784_),
    .A(_01758_),
    .B(_01783_));
 sg13g2_xor2_1 _07793_ (.B(_01782_),
    .A(_01755_),
    .X(_01785_));
 sg13g2_mux2_1 _07794_ (.A0(_01755_),
    .A1(_01785_),
    .S(_01758_),
    .X(_01786_));
 sg13g2_xnor2_1 _07795_ (.Y(_01787_),
    .A(_01754_),
    .B(_01786_));
 sg13g2_xnor2_1 _07796_ (.Y(_01788_),
    .A(_01781_),
    .B(_01787_));
 sg13g2_nand2b_1 _07797_ (.Y(_01789_),
    .B(_01780_),
    .A_N(_01788_));
 sg13g2_xor2_1 _07798_ (.B(_01788_),
    .A(_01780_),
    .X(_01790_));
 sg13g2_a21oi_1 _07799_ (.A1(_01750_),
    .A2(_01768_),
    .Y(_01791_),
    .B1(_01767_));
 sg13g2_nor2_1 _07800_ (.A(_01790_),
    .B(_01791_),
    .Y(_01792_));
 sg13g2_xor2_1 _07801_ (.B(_01791_),
    .A(_01790_),
    .X(_01793_));
 sg13g2_or2_1 _07802_ (.X(_01794_),
    .B(_01793_),
    .A(_01779_));
 sg13g2_a21oi_1 _07803_ (.A1(_01779_),
    .A2(_01793_),
    .Y(_01795_),
    .B1(net2944));
 sg13g2_a21o_1 _07804_ (.A2(_01795_),
    .A1(_01794_),
    .B1(_01777_),
    .X(_00163_));
 sg13g2_and2_1 _07805_ (.A(net1115),
    .B(_01392_),
    .X(_01796_));
 sg13g2_o21ai_1 _07806_ (.B1(_01789_),
    .Y(_01797_),
    .A1(_01781_),
    .A2(_01787_));
 sg13g2_mux2_1 _07807_ (.A0(_01752_),
    .A1(_01753_),
    .S(_01785_),
    .X(_01798_));
 sg13g2_xnor2_1 _07808_ (.Y(_01799_),
    .A(_01784_),
    .B(_01798_));
 sg13g2_o21ai_1 _07809_ (.B1(_01799_),
    .Y(_01800_),
    .A1(_01754_),
    .A2(_01758_));
 sg13g2_xnor2_1 _07810_ (.Y(_01801_),
    .A(_01797_),
    .B(_01800_));
 sg13g2_nor2_1 _07811_ (.A(_01792_),
    .B(_01801_),
    .Y(_01802_));
 sg13g2_a21o_1 _07812_ (.A2(_01802_),
    .A1(_01795_),
    .B1(_01796_),
    .X(_00164_));
 sg13g2_o21ai_1 _07813_ (.B1(net3024),
    .Y(_01803_),
    .A1(_01320_),
    .A2(net2977));
 sg13g2_nand2_1 _07814_ (.Y(_01804_),
    .A(net3225),
    .B(net2939));
 sg13g2_and3_2 _07815_ (.X(_01805_),
    .A(net3180),
    .B(net958),
    .C(_00036_));
 sg13g2_mux2_1 _07816_ (.A0(\u_toplayer.outreg[64] ),
    .A1(\u_toplayer.outreg[72] ),
    .S(net3188),
    .X(_01806_));
 sg13g2_mux2_1 _07817_ (.A0(\u_toplayer.outreg[32] ),
    .A1(\u_toplayer.outreg[40] ),
    .S(net3187),
    .X(_01807_));
 sg13g2_nand2b_1 _07818_ (.Y(_01808_),
    .B(_01807_),
    .A_N(net3185));
 sg13g2_a22oi_1 _07819_ (.Y(_01809_),
    .B1(net3012),
    .B2(\u_toplayer.outreg[56] ),
    .A2(net3015),
    .A1(\u_toplayer.outreg[48] ));
 sg13g2_nand3_1 _07820_ (.B(_01808_),
    .C(_01809_),
    .A(net3183),
    .Y(_01810_));
 sg13g2_mux2_1 _07821_ (.A0(\u_toplayer.outreg[0] ),
    .A1(\u_toplayer.outreg[8] ),
    .S(net3190),
    .X(_01811_));
 sg13g2_nand2b_1 _07822_ (.Y(_01812_),
    .B(_01811_),
    .A_N(net3184));
 sg13g2_a221oi_1 _07823_ (.B2(\u_toplayer.outreg[24] ),
    .C1(net3181),
    .B1(net3011),
    .A1(\u_toplayer.outreg[16] ),
    .Y(_01813_),
    .A2(net3014));
 sg13g2_a21oi_1 _07824_ (.A1(_01812_),
    .A2(_01813_),
    .Y(_01814_),
    .B1(net3179));
 sg13g2_a22oi_1 _07825_ (.Y(_01815_),
    .B1(_01810_),
    .B2(_01814_),
    .A2(_01806_),
    .A1(_01805_));
 sg13g2_o21ai_1 _07826_ (.B1(_01804_),
    .Y(_00165_),
    .A1(net2942),
    .A2(_01815_));
 sg13g2_nand2_1 _07827_ (.Y(_01816_),
    .A(net3223),
    .B(_01803_));
 sg13g2_mux2_1 _07828_ (.A0(\u_toplayer.outreg[65] ),
    .A1(\u_toplayer.outreg[73] ),
    .S(net3189),
    .X(_01817_));
 sg13g2_nor2b_1 _07829_ (.A(net3189),
    .B_N(\u_toplayer.outreg[1] ),
    .Y(_01818_));
 sg13g2_a21oi_1 _07830_ (.A1(\u_toplayer.outreg[9] ),
    .A2(net3189),
    .Y(_01819_),
    .B1(_01818_));
 sg13g2_a221oi_1 _07831_ (.B2(\u_toplayer.outreg[25] ),
    .C1(net3181),
    .B1(net3011),
    .A1(\u_toplayer.outreg[17] ),
    .Y(_01820_),
    .A2(net3014));
 sg13g2_o21ai_1 _07832_ (.B1(_01820_),
    .Y(_01821_),
    .A1(net3184),
    .A2(_01819_));
 sg13g2_mux2_1 _07833_ (.A0(\u_toplayer.outreg[33] ),
    .A1(\u_toplayer.outreg[41] ),
    .S(net3188),
    .X(_01822_));
 sg13g2_nand2b_1 _07834_ (.Y(_01823_),
    .B(_01822_),
    .A_N(net3184));
 sg13g2_a22oi_1 _07835_ (.Y(_01824_),
    .B1(net3011),
    .B2(\u_toplayer.outreg[57] ),
    .A2(net3015),
    .A1(\u_toplayer.outreg[49] ));
 sg13g2_nand3_1 _07836_ (.B(_01823_),
    .C(_01824_),
    .A(net3183),
    .Y(_01825_));
 sg13g2_nor2b_1 _07837_ (.A(net3179),
    .B_N(_01825_),
    .Y(_01826_));
 sg13g2_a22oi_1 _07838_ (.Y(_01827_),
    .B1(_01821_),
    .B2(_01826_),
    .A2(_01817_),
    .A1(_01805_));
 sg13g2_o21ai_1 _07839_ (.B1(_01816_),
    .Y(_00166_),
    .A1(net2942),
    .A2(_01827_));
 sg13g2_nand2_1 _07840_ (.Y(_01828_),
    .A(net3219),
    .B(_01803_));
 sg13g2_mux2_1 _07841_ (.A0(\u_toplayer.outreg[66] ),
    .A1(\u_toplayer.outreg[74] ),
    .S(net3190),
    .X(_01829_));
 sg13g2_mux2_1 _07842_ (.A0(\u_toplayer.outreg[34] ),
    .A1(\u_toplayer.outreg[42] ),
    .S(net3188),
    .X(_01830_));
 sg13g2_nand2b_1 _07843_ (.Y(_01831_),
    .B(_01830_),
    .A_N(net3184));
 sg13g2_a22oi_1 _07844_ (.Y(_01832_),
    .B1(net3011),
    .B2(\u_toplayer.outreg[58] ),
    .A2(net3015),
    .A1(\u_toplayer.outreg[50] ));
 sg13g2_nand3_1 _07845_ (.B(_01831_),
    .C(_01832_),
    .A(net3181),
    .Y(_01833_));
 sg13g2_mux2_1 _07846_ (.A0(\u_toplayer.outreg[2] ),
    .A1(\u_toplayer.outreg[10] ),
    .S(net3189),
    .X(_01834_));
 sg13g2_nand2b_1 _07847_ (.Y(_01835_),
    .B(_01834_),
    .A_N(net3186));
 sg13g2_a221oi_1 _07848_ (.B2(\u_toplayer.outreg[26] ),
    .C1(net3181),
    .B1(net3011),
    .A1(\u_toplayer.outreg[18] ),
    .Y(_01836_),
    .A2(net3014));
 sg13g2_a21oi_1 _07849_ (.A1(_01835_),
    .A2(_01836_),
    .Y(_01837_),
    .B1(net3179));
 sg13g2_a22oi_1 _07850_ (.Y(_01838_),
    .B1(_01833_),
    .B2(_01837_),
    .A2(_01829_),
    .A1(_01805_));
 sg13g2_o21ai_1 _07851_ (.B1(_01828_),
    .Y(_00167_),
    .A1(net2944),
    .A2(_01838_));
 sg13g2_nand2_1 _07852_ (.Y(_01839_),
    .A(net3217),
    .B(net2939));
 sg13g2_mux2_1 _07853_ (.A0(\u_toplayer.outreg[67] ),
    .A1(\u_toplayer.outreg[75] ),
    .S(net3190),
    .X(_01840_));
 sg13g2_nor2b_1 _07854_ (.A(net3189),
    .B_N(\u_toplayer.outreg[3] ),
    .Y(_01841_));
 sg13g2_a21oi_1 _07855_ (.A1(\u_toplayer.outreg[11] ),
    .A2(net3189),
    .Y(_01842_),
    .B1(_01841_));
 sg13g2_a221oi_1 _07856_ (.B2(\u_toplayer.outreg[27] ),
    .C1(net3181),
    .B1(net3011),
    .A1(\u_toplayer.outreg[19] ),
    .Y(_01843_),
    .A2(net3014));
 sg13g2_o21ai_1 _07857_ (.B1(_01843_),
    .Y(_01844_),
    .A1(net3186),
    .A2(_01842_));
 sg13g2_nor2b_1 _07858_ (.A(net3188),
    .B_N(\u_toplayer.outreg[35] ),
    .Y(_01845_));
 sg13g2_a21oi_1 _07859_ (.A1(\u_toplayer.outreg[43] ),
    .A2(net3188),
    .Y(_01846_),
    .B1(_01845_));
 sg13g2_a22oi_1 _07860_ (.Y(_01847_),
    .B1(net3011),
    .B2(\u_toplayer.outreg[59] ),
    .A2(net3015),
    .A1(\u_toplayer.outreg[51] ));
 sg13g2_o21ai_1 _07861_ (.B1(_01847_),
    .Y(_01848_),
    .A1(net3184),
    .A2(_01846_));
 sg13g2_inv_1 _07862_ (.Y(_01849_),
    .A(_01848_));
 sg13g2_a21oi_1 _07863_ (.A1(net3183),
    .A2(_01849_),
    .Y(_01850_),
    .B1(net3179));
 sg13g2_a22oi_1 _07864_ (.Y(_01851_),
    .B1(_01844_),
    .B2(_01850_),
    .A2(_01840_),
    .A1(_01805_));
 sg13g2_o21ai_1 _07865_ (.B1(_01839_),
    .Y(_00168_),
    .A1(net2944),
    .A2(_01851_));
 sg13g2_nand2_1 _07866_ (.Y(_01852_),
    .A(net3216),
    .B(net2939));
 sg13g2_mux2_1 _07867_ (.A0(\u_toplayer.outreg[68] ),
    .A1(\u_toplayer.outreg[76] ),
    .S(net3189),
    .X(_01853_));
 sg13g2_mux2_1 _07868_ (.A0(\u_toplayer.outreg[36] ),
    .A1(\u_toplayer.outreg[44] ),
    .S(net3188),
    .X(_01854_));
 sg13g2_nand2b_1 _07869_ (.Y(_01855_),
    .B(_01854_),
    .A_N(net3184));
 sg13g2_a22oi_1 _07870_ (.Y(_01856_),
    .B1(net3013),
    .B2(\u_toplayer.outreg[60] ),
    .A2(net3015),
    .A1(\u_toplayer.outreg[52] ));
 sg13g2_nand3_1 _07871_ (.B(_01855_),
    .C(_01856_),
    .A(net3181),
    .Y(_01857_));
 sg13g2_mux2_1 _07872_ (.A0(\u_toplayer.outreg[4] ),
    .A1(\u_toplayer.outreg[12] ),
    .S(net3189),
    .X(_01858_));
 sg13g2_nand2b_1 _07873_ (.Y(_01859_),
    .B(_01858_),
    .A_N(net3186));
 sg13g2_a221oi_1 _07874_ (.B2(\u_toplayer.outreg[28] ),
    .C1(net3181),
    .B1(net3011),
    .A1(\u_toplayer.outreg[20] ),
    .Y(_01860_),
    .A2(net3014));
 sg13g2_a21oi_1 _07875_ (.A1(_01859_),
    .A2(_01860_),
    .Y(_01861_),
    .B1(net3179));
 sg13g2_a22oi_1 _07876_ (.Y(_01862_),
    .B1(_01857_),
    .B2(_01861_),
    .A2(_01853_),
    .A1(_01805_));
 sg13g2_o21ai_1 _07877_ (.B1(_01852_),
    .Y(_00169_),
    .A1(net2944),
    .A2(_01862_));
 sg13g2_nand2_1 _07878_ (.Y(_01863_),
    .A(net3214),
    .B(net2939));
 sg13g2_mux2_1 _07879_ (.A0(\u_toplayer.outreg[69] ),
    .A1(\u_toplayer.outreg[77] ),
    .S(net3190),
    .X(_01864_));
 sg13g2_mux2_1 _07880_ (.A0(\u_toplayer.outreg[37] ),
    .A1(\u_toplayer.outreg[45] ),
    .S(net3187),
    .X(_01865_));
 sg13g2_nand2b_1 _07881_ (.Y(_01866_),
    .B(_01865_),
    .A_N(net3185));
 sg13g2_a22oi_1 _07882_ (.Y(_01867_),
    .B1(net3012),
    .B2(\u_toplayer.outreg[61] ),
    .A2(_01321_),
    .A1(\u_toplayer.outreg[53] ));
 sg13g2_nand3_1 _07883_ (.B(_01866_),
    .C(_01867_),
    .A(net3182),
    .Y(_01868_));
 sg13g2_mux2_1 _07884_ (.A0(\u_toplayer.outreg[5] ),
    .A1(\u_toplayer.outreg[13] ),
    .S(net3191),
    .X(_01869_));
 sg13g2_nand2b_1 _07885_ (.Y(_01870_),
    .B(_01869_),
    .A_N(net3186));
 sg13g2_a221oi_1 _07886_ (.B2(\u_toplayer.outreg[29] ),
    .C1(net3182),
    .B1(net3012),
    .A1(\u_toplayer.outreg[21] ),
    .Y(_01871_),
    .A2(net3014));
 sg13g2_a21oi_1 _07887_ (.A1(_01870_),
    .A2(_01871_),
    .Y(_01872_),
    .B1(net3180));
 sg13g2_a22oi_1 _07888_ (.Y(_01873_),
    .B1(_01868_),
    .B2(_01872_),
    .A2(_01864_),
    .A1(_01805_));
 sg13g2_o21ai_1 _07889_ (.B1(_01863_),
    .Y(_00170_),
    .A1(net2942),
    .A2(_01873_));
 sg13g2_nand2_1 _07890_ (.Y(_01874_),
    .A(net3211),
    .B(net2939));
 sg13g2_mux2_1 _07891_ (.A0(\u_toplayer.outreg[70] ),
    .A1(\u_toplayer.outreg[78] ),
    .S(net3190),
    .X(_01875_));
 sg13g2_mux2_1 _07892_ (.A0(\u_toplayer.outreg[38] ),
    .A1(\u_toplayer.outreg[46] ),
    .S(net3187),
    .X(_01876_));
 sg13g2_nand2b_1 _07893_ (.Y(_01877_),
    .B(_01876_),
    .A_N(net3185));
 sg13g2_a22oi_1 _07894_ (.Y(_01878_),
    .B1(net3012),
    .B2(\u_toplayer.outreg[62] ),
    .A2(net3016),
    .A1(\u_toplayer.outreg[54] ));
 sg13g2_nand3_1 _07895_ (.B(_01877_),
    .C(_01878_),
    .A(net3183),
    .Y(_01879_));
 sg13g2_mux2_1 _07896_ (.A0(\u_toplayer.outreg[6] ),
    .A1(\u_toplayer.outreg[14] ),
    .S(net3190),
    .X(_01880_));
 sg13g2_nand2b_1 _07897_ (.Y(_01881_),
    .B(_01880_),
    .A_N(net3186));
 sg13g2_a221oi_1 _07898_ (.B2(\u_toplayer.outreg[30] ),
    .C1(net3181),
    .B1(net3012),
    .A1(\u_toplayer.outreg[22] ),
    .Y(_01882_),
    .A2(net3014));
 sg13g2_a21oi_1 _07899_ (.A1(_01881_),
    .A2(_01882_),
    .Y(_01883_),
    .B1(net3180));
 sg13g2_a22oi_1 _07900_ (.Y(_01884_),
    .B1(_01879_),
    .B2(_01883_),
    .A2(_01875_),
    .A1(_01805_));
 sg13g2_o21ai_1 _07901_ (.B1(_01874_),
    .Y(_00171_),
    .A1(net2942),
    .A2(_01884_));
 sg13g2_nand2_1 _07902_ (.Y(_01885_),
    .A(net3208),
    .B(net2939));
 sg13g2_mux2_1 _07903_ (.A0(\u_toplayer.outreg[71] ),
    .A1(\u_toplayer.outreg[79] ),
    .S(net3190),
    .X(_01886_));
 sg13g2_nor2b_1 _07904_ (.A(net3191),
    .B_N(\u_toplayer.outreg[7] ),
    .Y(_01887_));
 sg13g2_a21oi_1 _07905_ (.A1(\u_toplayer.outreg[15] ),
    .A2(net3191),
    .Y(_01888_),
    .B1(_01887_));
 sg13g2_a221oi_1 _07906_ (.B2(\u_toplayer.outreg[31] ),
    .C1(net3182),
    .B1(net3012),
    .A1(\u_toplayer.outreg[23] ),
    .Y(_01889_),
    .A2(net3014));
 sg13g2_o21ai_1 _07907_ (.B1(_01889_),
    .Y(_01890_),
    .A1(net3186),
    .A2(_01888_));
 sg13g2_nor2b_1 _07908_ (.A(net3187),
    .B_N(\u_toplayer.outreg[39] ),
    .Y(_01891_));
 sg13g2_a21oi_1 _07909_ (.A1(\u_toplayer.outreg[47] ),
    .A2(net3187),
    .Y(_01892_),
    .B1(_01891_));
 sg13g2_a22oi_1 _07910_ (.Y(_01893_),
    .B1(net3012),
    .B2(\u_toplayer.outreg[63] ),
    .A2(net3016),
    .A1(\u_toplayer.outreg[55] ));
 sg13g2_o21ai_1 _07911_ (.B1(_01893_),
    .Y(_01894_),
    .A1(net3184),
    .A2(_01892_));
 sg13g2_inv_1 _07912_ (.Y(_01895_),
    .A(_01894_));
 sg13g2_a21oi_1 _07913_ (.A1(net3182),
    .A2(_01895_),
    .Y(_01896_),
    .B1(net3179));
 sg13g2_a22oi_1 _07914_ (.Y(_01897_),
    .B1(_01890_),
    .B2(_01896_),
    .A2(_01886_),
    .A1(_01805_));
 sg13g2_o21ai_1 _07915_ (.B1(_01885_),
    .Y(_00172_),
    .A1(net2942),
    .A2(_01897_));
 sg13g2_nand3_1 _07916_ (.B(net3016),
    .C(_01389_),
    .A(\u_toplayer.delayed_done_layer3 ),
    .Y(_01898_));
 sg13g2_nand2_1 _07917_ (.Y(_01899_),
    .A(net903),
    .B(_01898_));
 sg13g2_nor4_1 _07918_ (.A(\u_toplayer.u_outlayer.u_neuron.acc[12] ),
    .B(\u_toplayer.u_outlayer.u_neuron.acc[11] ),
    .C(\u_toplayer.u_outlayer.u_neuron.acc[10] ),
    .D(net3199),
    .Y(_01900_));
 sg13g2_nor4_1 _07919_ (.A(\u_toplayer.u_outlayer.u_neuron.acc[7] ),
    .B(\u_toplayer.u_outlayer.u_neuron.acc[15] ),
    .C(\u_toplayer.u_outlayer.u_neuron.acc[14] ),
    .D(\u_toplayer.u_outlayer.u_neuron.acc[13] ),
    .Y(_01901_));
 sg13g2_nor4_1 _07920_ (.A(\u_toplayer.u_outlayer.u_neuron.acc[8] ),
    .B(\u_toplayer.u_outlayer.u_neuron.acc[22] ),
    .C(\u_toplayer.u_outlayer.u_neuron.acc[21] ),
    .D(net3195),
    .Y(_01902_));
 sg13g2_nor4_1 _07921_ (.A(\u_toplayer.u_outlayer.u_neuron.acc[19] ),
    .B(net3196),
    .C(\u_toplayer.u_outlayer.u_neuron.acc[17] ),
    .D(net3197),
    .Y(_01903_));
 sg13g2_and3_1 _07922_ (.X(_01904_),
    .A(_01900_),
    .B(_01901_),
    .C(_01903_));
 sg13g2_a21oi_2 _07923_ (.B1(\u_toplayer.u_outlayer.u_neuron.acc[23] ),
    .Y(_01905_),
    .A2(_01904_),
    .A1(_01902_));
 sg13g2_nor2_1 _07924_ (.A(\u_toplayer.u_outlayer.u_neuron.acc[0] ),
    .B(_01905_),
    .Y(_01906_));
 sg13g2_nor4_1 _07925_ (.A(\u_toplayer.u_outlayer.u_neuron.acc[3] ),
    .B(\u_toplayer.u_outlayer.u_neuron.acc[2] ),
    .C(net3201),
    .D(\u_toplayer.u_outlayer.u_neuron.acc[0] ),
    .Y(_01907_));
 sg13g2_nor3_1 _07926_ (.A(_01037_),
    .B(\u_toplayer.u_outlayer.u_neuron.acc[6] ),
    .C(net3200),
    .Y(_01908_));
 sg13g2_nand3_1 _07927_ (.B(_01907_),
    .C(_01908_),
    .A(_01039_),
    .Y(_01909_));
 sg13g2_nand4_1 _07928_ (.B(\u_toplayer.u_outlayer.u_neuron.acc[11] ),
    .C(\u_toplayer.u_outlayer.u_neuron.acc[10] ),
    .A(\u_toplayer.u_outlayer.u_neuron.acc[12] ),
    .Y(_01910_),
    .D(net3199));
 sg13g2_nand4_1 _07929_ (.B(\u_toplayer.u_outlayer.u_neuron.acc[15] ),
    .C(\u_toplayer.u_outlayer.u_neuron.acc[14] ),
    .A(\u_toplayer.u_outlayer.u_neuron.acc[7] ),
    .Y(_01911_),
    .D(\u_toplayer.u_outlayer.u_neuron.acc[13] ));
 sg13g2_nand4_1 _07930_ (.B(net3196),
    .C(\u_toplayer.u_outlayer.u_neuron.acc[17] ),
    .A(\u_toplayer.u_outlayer.u_neuron.acc[19] ),
    .Y(_01912_),
    .D(net3197));
 sg13g2_nand4_1 _07931_ (.B(\u_toplayer.u_outlayer.u_neuron.acc[22] ),
    .C(\u_toplayer.u_outlayer.u_neuron.acc[21] ),
    .A(\u_toplayer.u_outlayer.u_neuron.acc[8] ),
    .Y(_01913_),
    .D(net3195));
 sg13g2_nor4_1 _07932_ (.A(_01910_),
    .B(_01911_),
    .C(_01912_),
    .D(_01913_),
    .Y(_01914_));
 sg13g2_nand2_1 _07933_ (.Y(_01915_),
    .A(_01909_),
    .B(_01914_));
 sg13g2_a21o_2 _07934_ (.A2(_01915_),
    .A1(\u_toplayer.u_outlayer.u_neuron.acc[23] ),
    .B1(net2938),
    .X(_01916_));
 sg13g2_o21ai_1 _07935_ (.B1(net904),
    .Y(_00173_),
    .A1(_01906_),
    .A2(_01916_));
 sg13g2_nand2_1 _07936_ (.Y(_01917_),
    .A(net883),
    .B(net2938));
 sg13g2_nor2_1 _07937_ (.A(net3201),
    .B(_01905_),
    .Y(_01918_));
 sg13g2_o21ai_1 _07938_ (.B1(_01917_),
    .Y(_00174_),
    .A1(_01916_),
    .A2(_01918_));
 sg13g2_nand2_1 _07939_ (.Y(_01919_),
    .A(net807),
    .B(net2938));
 sg13g2_nor2_1 _07940_ (.A(\u_toplayer.u_outlayer.u_neuron.acc[2] ),
    .B(_01905_),
    .Y(_01920_));
 sg13g2_o21ai_1 _07941_ (.B1(_01919_),
    .Y(_00175_),
    .A1(_01916_),
    .A2(_01920_));
 sg13g2_nand2_1 _07942_ (.Y(_01921_),
    .A(net849),
    .B(net2938));
 sg13g2_nor2_1 _07943_ (.A(\u_toplayer.u_outlayer.u_neuron.acc[3] ),
    .B(_01905_),
    .Y(_01922_));
 sg13g2_o21ai_1 _07944_ (.B1(_01921_),
    .Y(_00176_),
    .A1(_01916_),
    .A2(_01922_));
 sg13g2_nand2_1 _07945_ (.Y(_01923_),
    .A(net899),
    .B(net2938));
 sg13g2_nor2_1 _07946_ (.A(\u_toplayer.u_outlayer.u_neuron.acc[4] ),
    .B(_01905_),
    .Y(_01924_));
 sg13g2_o21ai_1 _07947_ (.B1(_01923_),
    .Y(_00177_),
    .A1(_01916_),
    .A2(_01924_));
 sg13g2_nand2_1 _07948_ (.Y(_01925_),
    .A(net908),
    .B(net2938));
 sg13g2_nor2_1 _07949_ (.A(\u_toplayer.u_outlayer.u_neuron.acc[5] ),
    .B(_01905_),
    .Y(_01926_));
 sg13g2_o21ai_1 _07950_ (.B1(_01925_),
    .Y(_00178_),
    .A1(_01916_),
    .A2(_01926_));
 sg13g2_nand2_1 _07951_ (.Y(_01927_),
    .A(net866),
    .B(net2938));
 sg13g2_nor2_1 _07952_ (.A(\u_toplayer.u_outlayer.u_neuron.acc[6] ),
    .B(_01905_),
    .Y(_01928_));
 sg13g2_o21ai_1 _07953_ (.B1(_01927_),
    .Y(_00179_),
    .A1(_01916_),
    .A2(_01928_));
 sg13g2_mux2_1 _07954_ (.A0(\u_toplayer.u_outlayer.u_neuron.acc[23] ),
    .A1(net984),
    .S(net2938),
    .X(_00180_));
 sg13g2_nand3b_1 _07955_ (.B(_01333_),
    .C(\u_toplayer.u_layer3.u_neuron.instCtrl.state[5] ),
    .Y(_01929_),
    .A_N(net3098));
 sg13g2_nor3_2 _07956_ (.A(_00034_),
    .B(_01336_),
    .C(_01929_),
    .Y(_01930_));
 sg13g2_or3_2 _07957_ (.A(_00034_),
    .B(_01336_),
    .C(_01929_),
    .X(_01931_));
 sg13g2_nor2_1 _07958_ (.A(net3112),
    .B(_01929_),
    .Y(_01932_));
 sg13g2_o21ai_1 _07959_ (.B1(_00034_),
    .Y(_01933_),
    .A1(net3127),
    .A2(_01929_));
 sg13g2_nor2b_2 _07960_ (.A(net3127),
    .B_N(net3112),
    .Y(_01934_));
 sg13g2_nor2b_1 _07961_ (.A(_01932_),
    .B_N(_01933_),
    .Y(_01935_));
 sg13g2_nand2b_2 _07962_ (.Y(_01936_),
    .B(_01933_),
    .A_N(_01932_));
 sg13g2_o21ai_1 _07963_ (.B1(_01935_),
    .Y(_01937_),
    .A1(_01336_),
    .A2(_01929_));
 sg13g2_nand2_1 _07964_ (.Y(_01938_),
    .A(\u_toplayer.delayed_done_layer2 ),
    .B(_01937_));
 sg13g2_nor2_1 _07965_ (.A(net3018),
    .B(net3100),
    .Y(_01939_));
 sg13g2_nand4_1 _07966_ (.B(_01329_),
    .C(_01331_),
    .A(\u_toplayer.u_layer3.u_neuron.instCtrl.state[5] ),
    .Y(_01940_),
    .D(_01939_));
 sg13g2_and2_1 _07967_ (.A(net2817),
    .B(_01940_),
    .X(_01941_));
 sg13g2_nand2_1 _07968_ (.Y(_01942_),
    .A(net2817),
    .B(_01940_));
 sg13g2_nand2_1 _07969_ (.Y(_01943_),
    .A(net2895),
    .B(net2759));
 sg13g2_nand2_1 _07970_ (.Y(_01944_),
    .A(net927),
    .B(net2731));
 sg13g2_nand3_1 _07971_ (.B(net2863),
    .C(net2759),
    .A(net2895),
    .Y(_01945_));
 sg13g2_nand2_1 _07972_ (.Y(_01946_),
    .A(net3348),
    .B(net3178));
 sg13g2_o21ai_1 _07973_ (.B1(_01944_),
    .Y(_00181_),
    .A1(net2728),
    .A2(_01946_));
 sg13g2_nand4_1 _07974_ (.B(net3339),
    .C(net3178),
    .A(net3348),
    .Y(_01947_),
    .D(net3176));
 sg13g2_inv_1 _07975_ (.Y(_01948_),
    .A(_01947_));
 sg13g2_a22oi_1 _07976_ (.Y(_01949_),
    .B1(net3176),
    .B2(net3348),
    .A2(net3178),
    .A1(net3339));
 sg13g2_nor3_1 _07977_ (.A(net2728),
    .B(_01948_),
    .C(_01949_),
    .Y(_01950_));
 sg13g2_a21o_1 _07978_ (.A2(net2731),
    .A1(net995),
    .B1(_01950_),
    .X(_00182_));
 sg13g2_nand2_1 _07979_ (.Y(_01951_),
    .A(net889),
    .B(net2731));
 sg13g2_nand2_1 _07980_ (.Y(_01952_),
    .A(net3328),
    .B(net3178));
 sg13g2_and4_1 _07981_ (.A(net3348),
    .B(net3339),
    .C(net3176),
    .D(net3174),
    .X(_01953_));
 sg13g2_a22oi_1 _07982_ (.Y(_01954_),
    .B1(net3174),
    .B2(net3348),
    .A2(net3176),
    .A1(net3339));
 sg13g2_nor2_1 _07983_ (.A(_01953_),
    .B(_01954_),
    .Y(_01955_));
 sg13g2_nor3_1 _07984_ (.A(_01952_),
    .B(_01953_),
    .C(_01954_),
    .Y(_01956_));
 sg13g2_xnor2_1 _07985_ (.Y(_01957_),
    .A(_01952_),
    .B(_01955_));
 sg13g2_and2_1 _07986_ (.A(_01948_),
    .B(_01957_),
    .X(_01958_));
 sg13g2_xnor2_1 _07987_ (.Y(_01959_),
    .A(_01948_),
    .B(_01957_));
 sg13g2_o21ai_1 _07988_ (.B1(_01951_),
    .Y(_00183_),
    .A1(net2728),
    .A2(_01959_));
 sg13g2_nand2_1 _07989_ (.Y(_01960_),
    .A(net917),
    .B(net2731));
 sg13g2_nand2_2 _07990_ (.Y(_01961_),
    .A(net3315),
    .B(net3178));
 sg13g2_or2_1 _07991_ (.X(_01962_),
    .B(_01956_),
    .A(_01953_));
 sg13g2_nand2_1 _07992_ (.Y(_01963_),
    .A(net3331),
    .B(net3176));
 sg13g2_and4_1 _07993_ (.A(net3349),
    .B(net3338),
    .C(net3174),
    .D(net3171),
    .X(_01964_));
 sg13g2_nand4_1 _07994_ (.B(net3338),
    .C(net3174),
    .A(net3349),
    .Y(_01965_),
    .D(net3171));
 sg13g2_a22oi_1 _07995_ (.Y(_01966_),
    .B1(net3171),
    .B2(net3349),
    .A2(net3174),
    .A1(net3338));
 sg13g2_nor3_1 _07996_ (.A(_01963_),
    .B(_01964_),
    .C(_01966_),
    .Y(_01967_));
 sg13g2_o21ai_1 _07997_ (.B1(_01963_),
    .Y(_01968_),
    .A1(_01964_),
    .A2(_01966_));
 sg13g2_nor2b_1 _07998_ (.A(_01967_),
    .B_N(_01968_),
    .Y(_01969_));
 sg13g2_nand2_1 _07999_ (.Y(_01970_),
    .A(_01962_),
    .B(_01969_));
 sg13g2_nor2_1 _08000_ (.A(_01962_),
    .B(_01969_),
    .Y(_01971_));
 sg13g2_xor2_1 _08001_ (.B(_01969_),
    .A(_01962_),
    .X(_01972_));
 sg13g2_xnor2_1 _08002_ (.Y(_01973_),
    .A(_01961_),
    .B(_01972_));
 sg13g2_and2_1 _08003_ (.A(_01958_),
    .B(_01973_),
    .X(_01974_));
 sg13g2_xnor2_1 _08004_ (.Y(_01975_),
    .A(_01958_),
    .B(_01973_));
 sg13g2_o21ai_1 _08005_ (.B1(_01960_),
    .Y(_00184_),
    .A1(net2728),
    .A2(_01975_));
 sg13g2_nand2_1 _08006_ (.Y(_01976_),
    .A(net947),
    .B(net2731));
 sg13g2_a22oi_1 _08007_ (.Y(_01977_),
    .B1(net3176),
    .B2(net3315),
    .A2(net3178),
    .A1(net3304));
 sg13g2_nand2_2 _08008_ (.Y(_01978_),
    .A(net3304),
    .B(net3176));
 sg13g2_nor2_1 _08009_ (.A(_01961_),
    .B(_01978_),
    .Y(_01979_));
 sg13g2_or2_1 _08010_ (.X(_01980_),
    .B(_01978_),
    .A(_01961_));
 sg13g2_nand2b_1 _08011_ (.Y(_01981_),
    .B(_01980_),
    .A_N(_01977_));
 sg13g2_o21ai_1 _08012_ (.B1(_01965_),
    .Y(_01982_),
    .A1(_01963_),
    .A2(_01966_));
 sg13g2_nand2_1 _08013_ (.Y(_01983_),
    .A(net3331),
    .B(net3174));
 sg13g2_and4_1 _08014_ (.A(net3350),
    .B(net3338),
    .C(net3171),
    .D(net3168),
    .X(_01984_));
 sg13g2_nand4_1 _08015_ (.B(net3338),
    .C(net3171),
    .A(net3349),
    .Y(_01985_),
    .D(net3168));
 sg13g2_a22oi_1 _08016_ (.Y(_01986_),
    .B1(net3168),
    .B2(net3349),
    .A2(net3171),
    .A1(net3338));
 sg13g2_or3_1 _08017_ (.A(_01983_),
    .B(_01984_),
    .C(_01986_),
    .X(_01987_));
 sg13g2_o21ai_1 _08018_ (.B1(_01983_),
    .Y(_01988_),
    .A1(_01984_),
    .A2(_01986_));
 sg13g2_and3_1 _08019_ (.X(_01989_),
    .A(_01982_),
    .B(_01987_),
    .C(_01988_));
 sg13g2_nand3_1 _08020_ (.B(_01987_),
    .C(_01988_),
    .A(_01982_),
    .Y(_01990_));
 sg13g2_a21oi_1 _08021_ (.A1(_01987_),
    .A2(_01988_),
    .Y(_01991_),
    .B1(_01982_));
 sg13g2_nor2_1 _08022_ (.A(_01989_),
    .B(_01991_),
    .Y(_01992_));
 sg13g2_xnor2_1 _08023_ (.Y(_01993_),
    .A(_01981_),
    .B(_01992_));
 sg13g2_o21ai_1 _08024_ (.B1(_01970_),
    .Y(_01994_),
    .A1(_01961_),
    .A2(_01971_));
 sg13g2_and2_1 _08025_ (.A(_01993_),
    .B(_01994_),
    .X(_01995_));
 sg13g2_xor2_1 _08026_ (.B(_01994_),
    .A(_01993_),
    .X(_01996_));
 sg13g2_nand2_1 _08027_ (.Y(_01997_),
    .A(_01974_),
    .B(_01996_));
 sg13g2_xnor2_1 _08028_ (.Y(_01998_),
    .A(_01974_),
    .B(_01996_));
 sg13g2_o21ai_1 _08029_ (.B1(_01976_),
    .Y(_00185_),
    .A1(net2728),
    .A2(_01998_));
 sg13g2_nand2_1 _08030_ (.Y(_01999_),
    .A(net996),
    .B(net2731));
 sg13g2_o21ai_1 _08031_ (.B1(_01990_),
    .Y(_02000_),
    .A1(_01981_),
    .A2(_01991_));
 sg13g2_nand2_1 _08032_ (.Y(_02001_),
    .A(net3296),
    .B(net3178));
 sg13g2_nand2_1 _08033_ (.Y(_02002_),
    .A(net3315),
    .B(net3174));
 sg13g2_xor2_1 _08034_ (.B(_02002_),
    .A(_01978_),
    .X(_02003_));
 sg13g2_nand2b_1 _08035_ (.Y(_02004_),
    .B(_02003_),
    .A_N(_02001_));
 sg13g2_xnor2_1 _08036_ (.Y(_02005_),
    .A(_02001_),
    .B(_02003_));
 sg13g2_o21ai_1 _08037_ (.B1(_01985_),
    .Y(_02006_),
    .A1(_01983_),
    .A2(_01986_));
 sg13g2_nand2_1 _08038_ (.Y(_02007_),
    .A(net3332),
    .B(net3172));
 sg13g2_and4_1 _08039_ (.A(net3353),
    .B(net3340),
    .C(net3168),
    .D(net3165),
    .X(_02008_));
 sg13g2_nand4_1 _08040_ (.B(net3340),
    .C(net3168),
    .A(net3353),
    .Y(_02009_),
    .D(net3165));
 sg13g2_a22oi_1 _08041_ (.Y(_02010_),
    .B1(net3165),
    .B2(net3353),
    .A2(net3168),
    .A1(net3340));
 sg13g2_or3_1 _08042_ (.A(_02007_),
    .B(_02008_),
    .C(_02010_),
    .X(_02011_));
 sg13g2_o21ai_1 _08043_ (.B1(_02007_),
    .Y(_02012_),
    .A1(_02008_),
    .A2(_02010_));
 sg13g2_and3_1 _08044_ (.X(_02013_),
    .A(_02006_),
    .B(_02011_),
    .C(_02012_));
 sg13g2_nand3_1 _08045_ (.B(_02011_),
    .C(_02012_),
    .A(_02006_),
    .Y(_02014_));
 sg13g2_a21o_1 _08046_ (.A2(_02012_),
    .A1(_02011_),
    .B1(_02006_),
    .X(_02015_));
 sg13g2_nand3_1 _08047_ (.B(_02014_),
    .C(_02015_),
    .A(_02005_),
    .Y(_02016_));
 sg13g2_a21o_1 _08048_ (.A2(_02015_),
    .A1(_02014_),
    .B1(_02005_),
    .X(_02017_));
 sg13g2_and3_1 _08049_ (.X(_02018_),
    .A(_02000_),
    .B(_02016_),
    .C(_02017_));
 sg13g2_a21oi_1 _08050_ (.A1(_02016_),
    .A2(_02017_),
    .Y(_02019_),
    .B1(_02000_));
 sg13g2_a21o_1 _08051_ (.A2(_02017_),
    .A1(_02016_),
    .B1(_02000_),
    .X(_02020_));
 sg13g2_o21ai_1 _08052_ (.B1(_01980_),
    .Y(_02021_),
    .A1(_02018_),
    .A2(_02019_));
 sg13g2_nand3b_1 _08053_ (.B(_02020_),
    .C(_01979_),
    .Y(_02022_),
    .A_N(_02018_));
 sg13g2_and3_1 _08054_ (.X(_02023_),
    .A(_01995_),
    .B(_02021_),
    .C(_02022_));
 sg13g2_nand3_1 _08055_ (.B(_02021_),
    .C(_02022_),
    .A(_01995_),
    .Y(_02024_));
 sg13g2_a21oi_1 _08056_ (.A1(_02021_),
    .A2(_02022_),
    .Y(_02025_),
    .B1(_01995_));
 sg13g2_nor3_2 _08057_ (.A(_01997_),
    .B(_02023_),
    .C(_02025_),
    .Y(_02026_));
 sg13g2_o21ai_1 _08058_ (.B1(_01997_),
    .Y(_02027_),
    .A1(_02023_),
    .A2(_02025_));
 sg13g2_nand2b_1 _08059_ (.Y(_02028_),
    .B(_02027_),
    .A_N(net2728));
 sg13g2_o21ai_1 _08060_ (.B1(_01999_),
    .Y(_00186_),
    .A1(_02026_),
    .A2(_02028_));
 sg13g2_nand2_1 _08061_ (.Y(_02029_),
    .A(net857),
    .B(net2731));
 sg13g2_a21o_1 _08062_ (.A2(_02020_),
    .A1(_01979_),
    .B1(_02018_),
    .X(_02030_));
 sg13g2_o21ai_1 _08063_ (.B1(_02004_),
    .Y(_02031_),
    .A1(_01978_),
    .A2(_02002_));
 sg13g2_nand2_1 _08064_ (.Y(_02032_),
    .A(net3289),
    .B(net3178));
 sg13g2_nand2b_1 _08065_ (.Y(_02033_),
    .B(_02031_),
    .A_N(_02032_));
 sg13g2_xor2_1 _08066_ (.B(_02032_),
    .A(_02031_),
    .X(_02034_));
 sg13g2_a21o_1 _08067_ (.A2(_02015_),
    .A1(_02005_),
    .B1(_02013_),
    .X(_02035_));
 sg13g2_nand2_1 _08068_ (.Y(_02036_),
    .A(net3297),
    .B(net3177));
 sg13g2_nand2_1 _08069_ (.Y(_02037_),
    .A(net3302),
    .B(net3172));
 sg13g2_and4_1 _08070_ (.A(net3314),
    .B(net3303),
    .C(net3175),
    .D(net3171),
    .X(_02038_));
 sg13g2_a22oi_1 _08071_ (.Y(_02039_),
    .B1(net3171),
    .B2(net3314),
    .A2(net3175),
    .A1(net3303));
 sg13g2_nor3_1 _08072_ (.A(_02036_),
    .B(_02038_),
    .C(_02039_),
    .Y(_02040_));
 sg13g2_o21ai_1 _08073_ (.B1(_02036_),
    .Y(_02041_),
    .A1(_02038_),
    .A2(_02039_));
 sg13g2_nand2b_1 _08074_ (.Y(_02042_),
    .B(_02041_),
    .A_N(_02040_));
 sg13g2_o21ai_1 _08075_ (.B1(_02009_),
    .Y(_02043_),
    .A1(_02007_),
    .A2(_02010_));
 sg13g2_and2_1 _08076_ (.A(net3332),
    .B(net3169),
    .X(_02044_));
 sg13g2_nand2_1 _08077_ (.Y(_02045_),
    .A(net3332),
    .B(net3168));
 sg13g2_and2_1 _08078_ (.A(net3340),
    .B(net3163),
    .X(_02046_));
 sg13g2_and4_1 _08079_ (.A(net3353),
    .B(net3340),
    .C(net3165),
    .D(net3163),
    .X(_02047_));
 sg13g2_nand4_1 _08080_ (.B(net3340),
    .C(net3165),
    .A(net3353),
    .Y(_02048_),
    .D(net3163));
 sg13g2_a22oi_1 _08081_ (.Y(_02049_),
    .B1(net3163),
    .B2(net3353),
    .A2(net3165),
    .A1(net3340));
 sg13g2_nand3b_1 _08082_ (.B(_02044_),
    .C(_02048_),
    .Y(_02050_),
    .A_N(_02049_));
 sg13g2_o21ai_1 _08083_ (.B1(_02045_),
    .Y(_02051_),
    .A1(_02047_),
    .A2(_02049_));
 sg13g2_and3_1 _08084_ (.X(_02052_),
    .A(_02043_),
    .B(_02050_),
    .C(_02051_));
 sg13g2_nand3_1 _08085_ (.B(_02050_),
    .C(_02051_),
    .A(_02043_),
    .Y(_02053_));
 sg13g2_a21oi_1 _08086_ (.A1(_02050_),
    .A2(_02051_),
    .Y(_02054_),
    .B1(_02043_));
 sg13g2_or3_1 _08087_ (.A(_02042_),
    .B(_02052_),
    .C(_02054_),
    .X(_02055_));
 sg13g2_o21ai_1 _08088_ (.B1(_02042_),
    .Y(_02056_),
    .A1(_02052_),
    .A2(_02054_));
 sg13g2_and3_1 _08089_ (.X(_02057_),
    .A(_02035_),
    .B(_02055_),
    .C(_02056_));
 sg13g2_nand3_1 _08090_ (.B(_02055_),
    .C(_02056_),
    .A(_02035_),
    .Y(_02058_));
 sg13g2_a21oi_1 _08091_ (.A1(_02055_),
    .A2(_02056_),
    .Y(_02059_),
    .B1(_02035_));
 sg13g2_o21ai_1 _08092_ (.B1(_02034_),
    .Y(_02060_),
    .A1(_02057_),
    .A2(_02059_));
 sg13g2_or3_1 _08093_ (.A(_02034_),
    .B(_02057_),
    .C(_02059_),
    .X(_02061_));
 sg13g2_and3_2 _08094_ (.X(_02062_),
    .A(_02030_),
    .B(_02060_),
    .C(_02061_));
 sg13g2_a21oi_1 _08095_ (.A1(_02060_),
    .A2(_02061_),
    .Y(_02063_),
    .B1(_02030_));
 sg13g2_nor3_1 _08096_ (.A(_02024_),
    .B(_02062_),
    .C(_02063_),
    .Y(_02064_));
 sg13g2_o21ai_1 _08097_ (.B1(_02024_),
    .Y(_02065_),
    .A1(_02062_),
    .A2(_02063_));
 sg13g2_nor2b_1 _08098_ (.A(_02064_),
    .B_N(_02065_),
    .Y(_02066_));
 sg13g2_xnor2_1 _08099_ (.Y(_02067_),
    .A(_02026_),
    .B(_02066_));
 sg13g2_o21ai_1 _08100_ (.B1(_02029_),
    .Y(_00187_),
    .A1(net2728),
    .A2(_02067_));
 sg13g2_a21oi_1 _08101_ (.A1(_02026_),
    .A2(_02065_),
    .Y(_02068_),
    .B1(_02064_));
 sg13g2_o21ai_1 _08102_ (.B1(_02058_),
    .Y(_02069_),
    .A1(_02034_),
    .A2(_02059_));
 sg13g2_or2_1 _08103_ (.X(_02070_),
    .B(_02040_),
    .A(_02038_));
 sg13g2_nor2_1 _08104_ (.A(net3281),
    .B(\u_toplayer.u_layer3.u_neuron.din[0] ),
    .Y(_02071_));
 sg13g2_nand2_2 _08105_ (.Y(_02072_),
    .A(net3289),
    .B(net3175));
 sg13g2_nand2_1 _08106_ (.Y(_02073_),
    .A(net3297),
    .B(net3174));
 sg13g2_nand2_1 _08107_ (.Y(_02074_),
    .A(net3290),
    .B(net3176));
 sg13g2_nor2_1 _08108_ (.A(_02036_),
    .B(_02072_),
    .Y(_02075_));
 sg13g2_xor2_1 _08109_ (.B(_02074_),
    .A(_02073_),
    .X(_02076_));
 sg13g2_xor2_1 _08110_ (.B(_02076_),
    .A(_02071_),
    .X(_02077_));
 sg13g2_nand2_1 _08111_ (.Y(_02078_),
    .A(_02070_),
    .B(_02077_));
 sg13g2_xnor2_1 _08112_ (.Y(_02079_),
    .A(_02070_),
    .B(_02077_));
 sg13g2_inv_1 _08113_ (.Y(_02080_),
    .A(_02079_));
 sg13g2_o21ai_1 _08114_ (.B1(_02053_),
    .Y(_02081_),
    .A1(_02042_),
    .A2(_02054_));
 sg13g2_and2_1 _08115_ (.A(net3314),
    .B(net3165),
    .X(_02082_));
 sg13g2_nand2_1 _08116_ (.Y(_02083_),
    .A(_02044_),
    .B(_02082_));
 sg13g2_a22oi_1 _08117_ (.Y(_02084_),
    .B1(net3165),
    .B2(net3332),
    .A2(net3168),
    .A1(net3314));
 sg13g2_a21oi_1 _08118_ (.A1(_02044_),
    .A2(_02082_),
    .Y(_02085_),
    .B1(_02084_));
 sg13g2_xnor2_1 _08119_ (.Y(_02086_),
    .A(_02037_),
    .B(_02085_));
 sg13g2_o21ai_1 _08120_ (.B1(_02048_),
    .Y(_02087_),
    .A1(_02045_),
    .A2(_02049_));
 sg13g2_nand3_1 _08121_ (.B(net3286),
    .C(net3160),
    .A(net3353),
    .Y(_02088_));
 sg13g2_a21o_1 _08122_ (.A2(net3160),
    .A1(net3354),
    .B1(net3286),
    .X(_02089_));
 sg13g2_nand3_1 _08123_ (.B(_02088_),
    .C(_02089_),
    .A(_02046_),
    .Y(_02090_));
 sg13g2_a21o_1 _08124_ (.A2(_02089_),
    .A1(_02088_),
    .B1(_02046_),
    .X(_02091_));
 sg13g2_nand3_1 _08125_ (.B(_02090_),
    .C(_02091_),
    .A(_02087_),
    .Y(_02092_));
 sg13g2_a21o_1 _08126_ (.A2(_02091_),
    .A1(_02090_),
    .B1(_02087_),
    .X(_02093_));
 sg13g2_nand3_1 _08127_ (.B(_02092_),
    .C(_02093_),
    .A(_02086_),
    .Y(_02094_));
 sg13g2_a21o_1 _08128_ (.A2(_02093_),
    .A1(_02092_),
    .B1(_02086_),
    .X(_02095_));
 sg13g2_nand3_1 _08129_ (.B(_02094_),
    .C(_02095_),
    .A(_02081_),
    .Y(_02096_));
 sg13g2_a21o_1 _08130_ (.A2(_02095_),
    .A1(_02094_),
    .B1(_02081_),
    .X(_02097_));
 sg13g2_nand3_1 _08131_ (.B(_02096_),
    .C(_02097_),
    .A(_02080_),
    .Y(_02098_));
 sg13g2_a21o_1 _08132_ (.A2(_02097_),
    .A1(_02096_),
    .B1(_02080_),
    .X(_02099_));
 sg13g2_and3_1 _08133_ (.X(_02100_),
    .A(_02069_),
    .B(_02098_),
    .C(_02099_));
 sg13g2_a21oi_1 _08134_ (.A1(_02098_),
    .A2(_02099_),
    .Y(_02101_),
    .B1(_02069_));
 sg13g2_o21ai_1 _08135_ (.B1(_02033_),
    .Y(_02102_),
    .A1(_02100_),
    .A2(_02101_));
 sg13g2_or3_1 _08136_ (.A(_02033_),
    .B(_02100_),
    .C(_02101_),
    .X(_02103_));
 sg13g2_and2_1 _08137_ (.A(_02102_),
    .B(_02103_),
    .X(_02104_));
 sg13g2_nand3_1 _08138_ (.B(_02102_),
    .C(_02103_),
    .A(_02062_),
    .Y(_02105_));
 sg13g2_a21oi_1 _08139_ (.A1(_02102_),
    .A2(_02103_),
    .Y(_02106_),
    .B1(_02062_));
 sg13g2_xnor2_1 _08140_ (.Y(_02107_),
    .A(_02062_),
    .B(_02104_));
 sg13g2_or2_1 _08141_ (.X(_02108_),
    .B(_02107_),
    .A(_02068_));
 sg13g2_a21oi_1 _08142_ (.A1(_02068_),
    .A2(_02107_),
    .Y(_02109_),
    .B1(net2728));
 sg13g2_a22oi_1 _08143_ (.Y(_02110_),
    .B1(_02108_),
    .B2(_02109_),
    .A2(net2730),
    .A1(net942));
 sg13g2_inv_1 _08144_ (.Y(_00188_),
    .A(_02110_));
 sg13g2_nand2_1 _08145_ (.Y(_02111_),
    .A(net963),
    .B(net2730));
 sg13g2_nand2_1 _08146_ (.Y(_02112_),
    .A(_02096_),
    .B(_02098_));
 sg13g2_a21oi_1 _08147_ (.A1(_02071_),
    .A2(_02076_),
    .Y(_02113_),
    .B1(_02075_));
 sg13g2_o21ai_1 _08148_ (.B1(_02083_),
    .Y(_02114_),
    .A1(_02037_),
    .A2(_02084_));
 sg13g2_nor2_1 _08149_ (.A(net3281),
    .B(net3177),
    .Y(_02115_));
 sg13g2_nor3_2 _08150_ (.A(net3283),
    .B(net3177),
    .C(_02072_),
    .Y(_02116_));
 sg13g2_xnor2_1 _08151_ (.Y(_02117_),
    .A(_02072_),
    .B(_02115_));
 sg13g2_nand2_1 _08152_ (.Y(_02118_),
    .A(_02114_),
    .B(_02117_));
 sg13g2_xnor2_1 _08153_ (.Y(_02119_),
    .A(_02114_),
    .B(_02117_));
 sg13g2_xnor2_1 _08154_ (.Y(_02120_),
    .A(_02113_),
    .B(_02119_));
 sg13g2_nand2_1 _08155_ (.Y(_02121_),
    .A(_02092_),
    .B(_02094_));
 sg13g2_nand2_1 _08156_ (.Y(_02122_),
    .A(net3296),
    .B(net3172));
 sg13g2_and3_1 _08157_ (.X(_02123_),
    .A(net3302),
    .B(net3169),
    .C(_02082_));
 sg13g2_a21oi_1 _08158_ (.A1(net3302),
    .A2(net3169),
    .Y(_02124_),
    .B1(_02082_));
 sg13g2_nor3_1 _08159_ (.A(_02122_),
    .B(_02123_),
    .C(_02124_),
    .Y(_02125_));
 sg13g2_o21ai_1 _08160_ (.B1(_02122_),
    .Y(_02126_),
    .A1(_02123_),
    .A2(_02124_));
 sg13g2_nand2b_1 _08161_ (.Y(_02127_),
    .B(_02126_),
    .A_N(_02125_));
 sg13g2_nand2_1 _08162_ (.Y(_02128_),
    .A(_02088_),
    .B(_02090_));
 sg13g2_and3_1 _08163_ (.X(_02129_),
    .A(net3354),
    .B(net3341),
    .C(net3162));
 sg13g2_nand3_1 _08164_ (.B(net3341),
    .C(net3160),
    .A(net3354),
    .Y(_02130_));
 sg13g2_o21ai_1 _08165_ (.B1(net3160),
    .Y(_02131_),
    .A1(net3354),
    .A2(net3341));
 sg13g2_nand2_1 _08166_ (.Y(_02132_),
    .A(net3332),
    .B(net3163));
 sg13g2_or3_1 _08167_ (.A(_02129_),
    .B(_02131_),
    .C(_02132_),
    .X(_02133_));
 sg13g2_o21ai_1 _08168_ (.B1(_02132_),
    .Y(_02134_),
    .A1(_02129_),
    .A2(_02131_));
 sg13g2_nand2_1 _08169_ (.Y(_02135_),
    .A(_02133_),
    .B(_02134_));
 sg13g2_nand2b_1 _08170_ (.Y(_02136_),
    .B(_02128_),
    .A_N(_02135_));
 sg13g2_xor2_1 _08171_ (.B(_02135_),
    .A(_02128_),
    .X(_02137_));
 sg13g2_xor2_1 _08172_ (.B(_02137_),
    .A(_02127_),
    .X(_02138_));
 sg13g2_nand2_1 _08173_ (.Y(_02139_),
    .A(_02121_),
    .B(_02138_));
 sg13g2_xnor2_1 _08174_ (.Y(_02140_),
    .A(_02121_),
    .B(_02138_));
 sg13g2_xnor2_1 _08175_ (.Y(_02141_),
    .A(_02120_),
    .B(_02140_));
 sg13g2_nand2b_1 _08176_ (.Y(_02142_),
    .B(_02112_),
    .A_N(_02141_));
 sg13g2_xor2_1 _08177_ (.B(_02141_),
    .A(_02112_),
    .X(_02143_));
 sg13g2_xor2_1 _08178_ (.B(_02143_),
    .A(_02078_),
    .X(_02144_));
 sg13g2_nand2b_1 _08179_ (.Y(_02145_),
    .B(_02103_),
    .A_N(_02100_));
 sg13g2_and2_1 _08180_ (.A(_02144_),
    .B(_02145_),
    .X(_02146_));
 sg13g2_xor2_1 _08181_ (.B(_02145_),
    .A(_02144_),
    .X(_02147_));
 sg13g2_o21ai_1 _08182_ (.B1(_02105_),
    .Y(_02148_),
    .A1(_02068_),
    .A2(_02106_));
 sg13g2_a21oi_1 _08183_ (.A1(_02147_),
    .A2(_02148_),
    .Y(_02149_),
    .B1(net2729));
 sg13g2_o21ai_1 _08184_ (.B1(_02149_),
    .Y(_02150_),
    .A1(_02147_),
    .A2(_02148_));
 sg13g2_nand2_1 _08185_ (.Y(_00189_),
    .A(_02111_),
    .B(_02150_));
 sg13g2_a21oi_1 _08186_ (.A1(_02147_),
    .A2(_02148_),
    .Y(_02151_),
    .B1(_02146_));
 sg13g2_o21ai_1 _08187_ (.B1(_02118_),
    .Y(_02152_),
    .A1(_02113_),
    .A2(_02119_));
 sg13g2_o21ai_1 _08188_ (.B1(_02139_),
    .Y(_02153_),
    .A1(_02120_),
    .A2(_02140_));
 sg13g2_or2_1 _08189_ (.X(_02154_),
    .B(_02125_),
    .A(_02123_));
 sg13g2_nand2_1 _08190_ (.Y(_02155_),
    .A(net3289),
    .B(net3172));
 sg13g2_nor2_1 _08191_ (.A(net3281),
    .B(net3175),
    .Y(_02156_));
 sg13g2_nor3_1 _08192_ (.A(net3281),
    .B(net3175),
    .C(_02155_),
    .Y(_02157_));
 sg13g2_xnor2_1 _08193_ (.Y(_02158_),
    .A(_02155_),
    .B(_02156_));
 sg13g2_and2_1 _08194_ (.A(_02154_),
    .B(_02158_),
    .X(_02159_));
 sg13g2_xor2_1 _08195_ (.B(_02158_),
    .A(_02154_),
    .X(_02160_));
 sg13g2_xnor2_1 _08196_ (.Y(_02161_),
    .A(_02116_),
    .B(_02160_));
 sg13g2_o21ai_1 _08197_ (.B1(_02136_),
    .Y(_02162_),
    .A1(_02127_),
    .A2(_02137_));
 sg13g2_nand2_1 _08198_ (.Y(_02163_),
    .A(net3296),
    .B(net3170));
 sg13g2_and4_1 _08199_ (.A(net3316),
    .B(net3303),
    .C(net3167),
    .D(net3164),
    .X(_02164_));
 sg13g2_a22oi_1 _08200_ (.Y(_02165_),
    .B1(net3164),
    .B2(net3314),
    .A2(net3167),
    .A1(net3303));
 sg13g2_nor2_1 _08201_ (.A(_02164_),
    .B(_02165_),
    .Y(_02166_));
 sg13g2_nand2b_1 _08202_ (.Y(_02167_),
    .B(_02166_),
    .A_N(_02163_));
 sg13g2_xor2_1 _08203_ (.B(_02166_),
    .A(_02163_),
    .X(_02168_));
 sg13g2_and2_1 _08204_ (.A(net3332),
    .B(net3162),
    .X(_02169_));
 sg13g2_nand2_1 _08205_ (.Y(_02170_),
    .A(net3332),
    .B(net3160));
 sg13g2_or3_1 _08206_ (.A(_02129_),
    .B(_02131_),
    .C(_02169_),
    .X(_02171_));
 sg13g2_o21ai_1 _08207_ (.B1(_02169_),
    .Y(_02172_),
    .A1(_02129_),
    .A2(_02131_));
 sg13g2_and4_1 _08208_ (.A(net3354),
    .B(net3341),
    .C(net3332),
    .D(net3160),
    .X(_02173_));
 sg13g2_nand4_1 _08209_ (.B(net3340),
    .C(net3333),
    .A(net3353),
    .Y(_02174_),
    .D(net3161));
 sg13g2_and4_1 _08210_ (.A(_02130_),
    .B(_02133_),
    .C(_02171_),
    .D(_02172_),
    .X(_02175_));
 sg13g2_or3_1 _08211_ (.A(_02168_),
    .B(_02173_),
    .C(_02175_),
    .X(_02176_));
 sg13g2_o21ai_1 _08212_ (.B1(_02168_),
    .Y(_02177_),
    .A1(_02173_),
    .A2(_02175_));
 sg13g2_nand2_1 _08213_ (.Y(_02178_),
    .A(_02176_),
    .B(_02177_));
 sg13g2_nand2b_1 _08214_ (.Y(_02179_),
    .B(_02162_),
    .A_N(_02178_));
 sg13g2_nor2b_1 _08215_ (.A(_02162_),
    .B_N(_02178_),
    .Y(_02180_));
 sg13g2_xnor2_1 _08216_ (.Y(_02181_),
    .A(_02162_),
    .B(_02178_));
 sg13g2_xnor2_1 _08217_ (.Y(_02182_),
    .A(_02161_),
    .B(_02181_));
 sg13g2_nand2_1 _08218_ (.Y(_02183_),
    .A(_02153_),
    .B(_02182_));
 sg13g2_xnor2_1 _08219_ (.Y(_02184_),
    .A(_02153_),
    .B(_02182_));
 sg13g2_nand2b_1 _08220_ (.Y(_02185_),
    .B(_02152_),
    .A_N(_02184_));
 sg13g2_xor2_1 _08221_ (.B(_02184_),
    .A(_02152_),
    .X(_02186_));
 sg13g2_o21ai_1 _08222_ (.B1(_02142_),
    .Y(_02187_),
    .A1(_02078_),
    .A2(_02143_));
 sg13g2_nor2b_1 _08223_ (.A(_02186_),
    .B_N(_02187_),
    .Y(_02188_));
 sg13g2_xnor2_1 _08224_ (.Y(_02189_),
    .A(_02186_),
    .B(_02187_));
 sg13g2_nor2b_1 _08225_ (.A(_02151_),
    .B_N(_02189_),
    .Y(_02190_));
 sg13g2_nor2b_1 _08226_ (.A(_02189_),
    .B_N(_02151_),
    .Y(_02191_));
 sg13g2_nor3_1 _08227_ (.A(net2729),
    .B(_02190_),
    .C(_02191_),
    .Y(_02192_));
 sg13g2_a21o_1 _08228_ (.A2(net2730),
    .A1(net957),
    .B1(_02192_),
    .X(_00190_));
 sg13g2_a21oi_1 _08229_ (.A1(_02116_),
    .A2(_02160_),
    .Y(_02193_),
    .B1(_02159_));
 sg13g2_o21ai_1 _08230_ (.B1(_02179_),
    .Y(_02194_),
    .A1(_02161_),
    .A2(_02180_));
 sg13g2_nand2b_1 _08231_ (.Y(_02195_),
    .B(_02167_),
    .A_N(_02164_));
 sg13g2_a22oi_1 _08232_ (.Y(_02196_),
    .B1(net3169),
    .B2(net3290),
    .A2(_01095_),
    .A1(net3286));
 sg13g2_nand3_1 _08233_ (.B(net3286),
    .C(net3169),
    .A(net3289),
    .Y(_02197_));
 sg13g2_nor2_1 _08234_ (.A(net3173),
    .B(_02197_),
    .Y(_02198_));
 sg13g2_nor2_1 _08235_ (.A(_02196_),
    .B(_02198_),
    .Y(_02199_));
 sg13g2_and2_1 _08236_ (.A(_02195_),
    .B(_02199_),
    .X(_02200_));
 sg13g2_xor2_1 _08237_ (.B(_02199_),
    .A(_02195_),
    .X(_02201_));
 sg13g2_xnor2_1 _08238_ (.Y(_02202_),
    .A(_02157_),
    .B(_02201_));
 sg13g2_nand2_1 _08239_ (.Y(_02203_),
    .A(_02174_),
    .B(_02176_));
 sg13g2_a22oi_1 _08240_ (.Y(_02204_),
    .B1(net3160),
    .B2(net3316),
    .A2(net3163),
    .A1(net3302));
 sg13g2_and3_1 _08241_ (.X(_02205_),
    .A(net3314),
    .B(net3302),
    .C(net3161));
 sg13g2_nand3_1 _08242_ (.B(net3302),
    .C(net3161),
    .A(net3314),
    .Y(_02206_));
 sg13g2_nand4_1 _08243_ (.B(net3302),
    .C(net3164),
    .A(net3316),
    .Y(_02207_),
    .D(net3160));
 sg13g2_nor2b_1 _08244_ (.A(_02204_),
    .B_N(_02207_),
    .Y(_02208_));
 sg13g2_nand2_1 _08245_ (.Y(_02209_),
    .A(net3296),
    .B(net3167));
 sg13g2_xor2_1 _08246_ (.B(_02209_),
    .A(_02208_),
    .X(_02210_));
 sg13g2_a21o_2 _08247_ (.A2(_02170_),
    .A1(_02131_),
    .B1(_02173_),
    .X(_02211_));
 sg13g2_xor2_1 _08248_ (.B(_02211_),
    .A(_02210_),
    .X(_02212_));
 sg13g2_nand2_1 _08249_ (.Y(_02213_),
    .A(_02203_),
    .B(_02212_));
 sg13g2_xnor2_1 _08250_ (.Y(_02214_),
    .A(_02203_),
    .B(_02212_));
 sg13g2_xor2_1 _08251_ (.B(_02214_),
    .A(_02202_),
    .X(_02215_));
 sg13g2_nand2_1 _08252_ (.Y(_02216_),
    .A(_02194_),
    .B(_02215_));
 sg13g2_xnor2_1 _08253_ (.Y(_02217_),
    .A(_02194_),
    .B(_02215_));
 sg13g2_or2_1 _08254_ (.X(_02218_),
    .B(_02217_),
    .A(_02193_));
 sg13g2_xnor2_1 _08255_ (.Y(_02219_),
    .A(_02193_),
    .B(_02217_));
 sg13g2_a21oi_1 _08256_ (.A1(_02183_),
    .A2(_02185_),
    .Y(_02220_),
    .B1(_02219_));
 sg13g2_nand3_1 _08257_ (.B(_02185_),
    .C(_02219_),
    .A(_02183_),
    .Y(_02221_));
 sg13g2_nand2b_1 _08258_ (.Y(_02222_),
    .B(_02221_),
    .A_N(_02220_));
 sg13g2_inv_1 _08259_ (.Y(_02223_),
    .A(_02222_));
 sg13g2_nor3_1 _08260_ (.A(_02188_),
    .B(_02190_),
    .C(_02223_),
    .Y(_02224_));
 sg13g2_o21ai_1 _08261_ (.B1(_02223_),
    .Y(_02225_),
    .A1(_02188_),
    .A2(_02190_));
 sg13g2_nor2_1 _08262_ (.A(net2729),
    .B(_02224_),
    .Y(_02226_));
 sg13g2_a22oi_1 _08263_ (.Y(_02227_),
    .B1(_02225_),
    .B2(_02226_),
    .A2(net2730),
    .A1(net990));
 sg13g2_inv_1 _08264_ (.Y(_00191_),
    .A(_02227_));
 sg13g2_nand2b_1 _08265_ (.Y(_02228_),
    .B(_02225_),
    .A_N(_02220_));
 sg13g2_a21oi_1 _08266_ (.A1(_02157_),
    .A2(_02201_),
    .Y(_02229_),
    .B1(_02200_));
 sg13g2_o21ai_1 _08267_ (.B1(_02213_),
    .Y(_02230_),
    .A1(_02202_),
    .A2(_02214_));
 sg13g2_o21ai_1 _08268_ (.B1(_02207_),
    .Y(_02231_),
    .A1(_02204_),
    .A2(_02209_));
 sg13g2_a22oi_1 _08269_ (.Y(_02232_),
    .B1(net3166),
    .B2(net3289),
    .A2(_01096_),
    .A1(net3286));
 sg13g2_and4_1 _08270_ (.A(net3289),
    .B(net3286),
    .C(_01096_),
    .D(net3166),
    .X(_02233_));
 sg13g2_nor2_1 _08271_ (.A(_02232_),
    .B(_02233_),
    .Y(_02234_));
 sg13g2_xnor2_1 _08272_ (.Y(_02235_),
    .A(_02231_),
    .B(_02234_));
 sg13g2_nor3_1 _08273_ (.A(net3173),
    .B(_02197_),
    .C(_02235_),
    .Y(_02236_));
 sg13g2_xnor2_1 _08274_ (.Y(_02237_),
    .A(_02198_),
    .B(_02235_));
 sg13g2_o21ai_1 _08275_ (.B1(_02174_),
    .Y(_02238_),
    .A1(_02210_),
    .A2(_02211_));
 sg13g2_o21ai_1 _08276_ (.B1(net3161),
    .Y(_02239_),
    .A1(net3314),
    .A2(net3302));
 sg13g2_nor2_1 _08277_ (.A(_02205_),
    .B(_02239_),
    .Y(_02240_));
 sg13g2_nand2_1 _08278_ (.Y(_02241_),
    .A(net3296),
    .B(net3164));
 sg13g2_nor3_1 _08279_ (.A(_02205_),
    .B(_02239_),
    .C(_02241_),
    .Y(_02242_));
 sg13g2_xor2_1 _08280_ (.B(_02241_),
    .A(_02240_),
    .X(_02243_));
 sg13g2_xnor2_1 _08281_ (.Y(_02244_),
    .A(_02211_),
    .B(_02243_));
 sg13g2_nor2b_1 _08282_ (.A(_02244_),
    .B_N(_02238_),
    .Y(_02245_));
 sg13g2_nand2b_1 _08283_ (.Y(_02246_),
    .B(_02244_),
    .A_N(_02238_));
 sg13g2_nand2b_1 _08284_ (.Y(_02247_),
    .B(_02246_),
    .A_N(_02245_));
 sg13g2_xnor2_1 _08285_ (.Y(_02248_),
    .A(_02237_),
    .B(_02247_));
 sg13g2_nand2_1 _08286_ (.Y(_02249_),
    .A(_02230_),
    .B(_02248_));
 sg13g2_xnor2_1 _08287_ (.Y(_02250_),
    .A(_02230_),
    .B(_02248_));
 sg13g2_xnor2_1 _08288_ (.Y(_02251_),
    .A(_02229_),
    .B(_02250_));
 sg13g2_a21o_1 _08289_ (.A2(_02218_),
    .A1(_02216_),
    .B1(_02251_),
    .X(_02252_));
 sg13g2_nand3_1 _08290_ (.B(_02218_),
    .C(_02251_),
    .A(_02216_),
    .Y(_02253_));
 sg13g2_a21oi_1 _08291_ (.A1(_02252_),
    .A2(_02253_),
    .Y(_02254_),
    .B1(_02228_));
 sg13g2_and3_1 _08292_ (.X(_02255_),
    .A(_02228_),
    .B(_02252_),
    .C(_02253_));
 sg13g2_nor3_1 _08293_ (.A(net2729),
    .B(_02254_),
    .C(_02255_),
    .Y(_02256_));
 sg13g2_a21o_1 _08294_ (.A2(net2730),
    .A1(net1012),
    .B1(_02256_),
    .X(_00192_));
 sg13g2_nand2_1 _08295_ (.Y(_02257_),
    .A(net998),
    .B(net2730));
 sg13g2_a21oi_2 _08296_ (.B1(_02236_),
    .Y(_02258_),
    .A2(_02234_),
    .A1(_02231_));
 sg13g2_a21oi_1 _08297_ (.A1(_02237_),
    .A2(_02246_),
    .Y(_02259_),
    .B1(_02245_));
 sg13g2_o21ai_1 _08298_ (.B1(_02174_),
    .Y(_02260_),
    .A1(_02211_),
    .A2(_02243_));
 sg13g2_nand2_1 _08299_ (.Y(_02261_),
    .A(net3296),
    .B(net3161));
 sg13g2_xor2_1 _08300_ (.B(_02261_),
    .A(_02240_),
    .X(_02262_));
 sg13g2_xnor2_1 _08301_ (.Y(_02263_),
    .A(_02211_),
    .B(_02262_));
 sg13g2_inv_1 _08302_ (.Y(_02264_),
    .A(_02263_));
 sg13g2_xor2_1 _08303_ (.B(_02263_),
    .A(_02260_),
    .X(_02265_));
 sg13g2_nor2_1 _08304_ (.A(_02205_),
    .B(_02242_),
    .Y(_02266_));
 sg13g2_nand2_1 _08305_ (.Y(_02267_),
    .A(net3289),
    .B(net3163));
 sg13g2_nor2_1 _08306_ (.A(net3281),
    .B(net3166),
    .Y(_02268_));
 sg13g2_nor3_1 _08307_ (.A(net3281),
    .B(net3167),
    .C(_02267_),
    .Y(_02269_));
 sg13g2_xnor2_1 _08308_ (.Y(_02270_),
    .A(_02267_),
    .B(_02268_));
 sg13g2_nand2b_1 _08309_ (.Y(_02271_),
    .B(_02270_),
    .A_N(_02266_));
 sg13g2_xnor2_1 _08310_ (.Y(_02272_),
    .A(_02266_),
    .B(_02270_));
 sg13g2_nand2_1 _08311_ (.Y(_02273_),
    .A(_02233_),
    .B(_02272_));
 sg13g2_xnor2_1 _08312_ (.Y(_02274_),
    .A(_02233_),
    .B(_02272_));
 sg13g2_nor2_1 _08313_ (.A(_02265_),
    .B(_02274_),
    .Y(_02275_));
 sg13g2_xor2_1 _08314_ (.B(_02274_),
    .A(_02265_),
    .X(_02276_));
 sg13g2_nand2b_1 _08315_ (.Y(_02277_),
    .B(_02276_),
    .A_N(_02259_));
 sg13g2_xnor2_1 _08316_ (.Y(_02278_),
    .A(_02259_),
    .B(_02276_));
 sg13g2_inv_1 _08317_ (.Y(_02279_),
    .A(_02278_));
 sg13g2_xnor2_1 _08318_ (.Y(_02280_),
    .A(_02258_),
    .B(_02278_));
 sg13g2_o21ai_1 _08319_ (.B1(_02249_),
    .Y(_02281_),
    .A1(_02229_),
    .A2(_02250_));
 sg13g2_xor2_1 _08320_ (.B(_02281_),
    .A(_02280_),
    .X(_02282_));
 sg13g2_nand3_1 _08321_ (.B(_02148_),
    .C(_02189_),
    .A(_02147_),
    .Y(_02283_));
 sg13g2_nor2b_1 _08322_ (.A(_02188_),
    .B_N(_02252_),
    .Y(_02284_));
 sg13g2_a22oi_1 _08323_ (.Y(_02285_),
    .B1(_02220_),
    .B2(_02253_),
    .A2(_02189_),
    .A1(_02146_));
 sg13g2_nand3_1 _08324_ (.B(_02284_),
    .C(_02285_),
    .A(_02283_),
    .Y(_02286_));
 sg13g2_nand2_1 _08325_ (.Y(_02287_),
    .A(_02221_),
    .B(_02253_));
 sg13g2_nand2_1 _08326_ (.Y(_02288_),
    .A(_02252_),
    .B(_02287_));
 sg13g2_nand3_1 _08327_ (.B(_02286_),
    .C(_02288_),
    .A(_02282_),
    .Y(_02289_));
 sg13g2_a21oi_1 _08328_ (.A1(_02286_),
    .A2(_02288_),
    .Y(_02290_),
    .B1(_02282_));
 sg13g2_nand2b_1 _08329_ (.Y(_02291_),
    .B(_02289_),
    .A_N(net2729));
 sg13g2_o21ai_1 _08330_ (.B1(_02257_),
    .Y(_00193_),
    .A1(_02290_),
    .A2(_02291_));
 sg13g2_nand2_1 _08331_ (.Y(_02292_),
    .A(net974),
    .B(net2730));
 sg13g2_nand2_1 _08332_ (.Y(_02293_),
    .A(_02271_),
    .B(_02273_));
 sg13g2_a21oi_1 _08333_ (.A1(_02260_),
    .A2(_02264_),
    .Y(_02294_),
    .B1(_02275_));
 sg13g2_or2_1 _08334_ (.X(_02295_),
    .B(_02262_),
    .A(_02174_));
 sg13g2_nand3_1 _08335_ (.B(_02211_),
    .C(_02262_),
    .A(_02174_),
    .Y(_02296_));
 sg13g2_inv_1 _08336_ (.Y(_02297_),
    .A(_02296_));
 sg13g2_and2_1 _08337_ (.A(_02295_),
    .B(_02296_),
    .X(_02298_));
 sg13g2_o21ai_1 _08338_ (.B1(_02206_),
    .Y(_02299_),
    .A1(_02239_),
    .A2(_02261_));
 sg13g2_nand2_1 _08339_ (.Y(_02300_),
    .A(net3289),
    .B(net3161));
 sg13g2_nor2_1 _08340_ (.A(net3281),
    .B(net3163),
    .Y(_02301_));
 sg13g2_nor2_1 _08341_ (.A(_02300_),
    .B(_02301_),
    .Y(_02302_));
 sg13g2_xnor2_1 _08342_ (.Y(_02303_),
    .A(_02300_),
    .B(_02301_));
 sg13g2_xor2_1 _08343_ (.B(_02303_),
    .A(_02299_),
    .X(_02304_));
 sg13g2_and2_1 _08344_ (.A(_02269_),
    .B(_02304_),
    .X(_02305_));
 sg13g2_xnor2_1 _08345_ (.Y(_02306_),
    .A(_02269_),
    .B(_02304_));
 sg13g2_xor2_1 _08346_ (.B(_02306_),
    .A(_02298_),
    .X(_02307_));
 sg13g2_nor2_1 _08347_ (.A(_02294_),
    .B(_02307_),
    .Y(_02308_));
 sg13g2_xor2_1 _08348_ (.B(_02307_),
    .A(_02294_),
    .X(_02309_));
 sg13g2_xor2_1 _08349_ (.B(_02309_),
    .A(_02293_),
    .X(_02310_));
 sg13g2_o21ai_1 _08350_ (.B1(_02277_),
    .Y(_02311_),
    .A1(_02258_),
    .A2(_02279_));
 sg13g2_nand2_1 _08351_ (.Y(_02312_),
    .A(_02310_),
    .B(_02311_));
 sg13g2_xor2_1 _08352_ (.B(_02311_),
    .A(_02310_),
    .X(_02313_));
 sg13g2_nand2b_1 _08353_ (.Y(_02314_),
    .B(_02313_),
    .A_N(_02289_));
 sg13g2_a21oi_1 _08354_ (.A1(_02280_),
    .A2(_02281_),
    .Y(_02315_),
    .B1(_02313_));
 sg13g2_and2_1 _08355_ (.A(_02289_),
    .B(_02315_),
    .X(_02316_));
 sg13g2_nand3_1 _08356_ (.B(_02281_),
    .C(_02313_),
    .A(_02280_),
    .Y(_02317_));
 sg13g2_nand3b_1 _08357_ (.B(_02314_),
    .C(_02317_),
    .Y(_02318_),
    .A_N(net2729));
 sg13g2_o21ai_1 _08358_ (.B1(_02292_),
    .Y(_00194_),
    .A1(_02316_),
    .A2(_02318_));
 sg13g2_nand2_1 _08359_ (.Y(_02319_),
    .A(net1021),
    .B(net2730));
 sg13g2_nand3_1 _08360_ (.B(_02314_),
    .C(_02317_),
    .A(_02312_),
    .Y(_02320_));
 sg13g2_a21o_1 _08361_ (.A2(_02303_),
    .A1(_02299_),
    .B1(_02305_),
    .X(_02321_));
 sg13g2_o21ai_1 _08362_ (.B1(_02295_),
    .Y(_02322_),
    .A1(_02297_),
    .A2(_02306_));
 sg13g2_nor2_1 _08363_ (.A(net3281),
    .B(net3161),
    .Y(_02323_));
 sg13g2_nor3_1 _08364_ (.A(_02299_),
    .B(_02302_),
    .C(_02323_),
    .Y(_02324_));
 sg13g2_o21ai_1 _08365_ (.B1(_02299_),
    .Y(_02325_),
    .A1(_02302_),
    .A2(_02323_));
 sg13g2_nand2b_1 _08366_ (.Y(_02326_),
    .B(_02325_),
    .A_N(_02324_));
 sg13g2_xnor2_1 _08367_ (.Y(_02327_),
    .A(_02298_),
    .B(_02326_));
 sg13g2_xnor2_1 _08368_ (.Y(_02328_),
    .A(_02322_),
    .B(_02327_));
 sg13g2_nor2b_1 _08369_ (.A(_02328_),
    .B_N(_02321_),
    .Y(_02329_));
 sg13g2_xnor2_1 _08370_ (.Y(_02330_),
    .A(_02321_),
    .B(_02328_));
 sg13g2_a21oi_1 _08371_ (.A1(_02293_),
    .A2(_02309_),
    .Y(_02331_),
    .B1(_02308_));
 sg13g2_nand2b_1 _08372_ (.Y(_02332_),
    .B(_02330_),
    .A_N(_02331_));
 sg13g2_xnor2_1 _08373_ (.Y(_02333_),
    .A(_02330_),
    .B(_02331_));
 sg13g2_nor2_1 _08374_ (.A(_02320_),
    .B(_02333_),
    .Y(_02334_));
 sg13g2_a21o_1 _08375_ (.A2(_02333_),
    .A1(_02320_),
    .B1(net2729),
    .X(_02335_));
 sg13g2_o21ai_1 _08376_ (.B1(_02319_),
    .Y(_00195_),
    .A1(_02334_),
    .A2(_02335_));
 sg13g2_nand2_1 _08377_ (.Y(_02336_),
    .A(net3204),
    .B(net2731));
 sg13g2_a21oi_1 _08378_ (.A1(_02295_),
    .A2(_02325_),
    .Y(_02337_),
    .B1(_02324_));
 sg13g2_nand2_1 _08379_ (.Y(_02338_),
    .A(_02296_),
    .B(_02337_));
 sg13g2_a21o_1 _08380_ (.A2(_02327_),
    .A1(_02322_),
    .B1(_02329_),
    .X(_02339_));
 sg13g2_a22oi_1 _08381_ (.Y(_02340_),
    .B1(_02338_),
    .B2(_02339_),
    .A2(_02324_),
    .A1(_02297_));
 sg13g2_nand2_1 _08382_ (.Y(_02341_),
    .A(_02332_),
    .B(_02340_));
 sg13g2_o21ai_1 _08383_ (.B1(_02336_),
    .Y(_00196_),
    .A1(_02335_),
    .A2(_02341_));
 sg13g2_and2_1 _08384_ (.A(_01322_),
    .B(net2939),
    .X(_02342_));
 sg13g2_nand2_2 _08385_ (.Y(_02343_),
    .A(_01322_),
    .B(net2939));
 sg13g2_nor2_1 _08386_ (.A(net1089),
    .B(_02343_),
    .Y(_02344_));
 sg13g2_and2_1 _08387_ (.A(_01320_),
    .B(net2979),
    .X(_02345_));
 sg13g2_nand2_2 _08388_ (.Y(_02346_),
    .A(_01320_),
    .B(net2979));
 sg13g2_nand2_1 _08389_ (.Y(_02347_),
    .A(\u_toplayer.u_outlayer.u_neuron.acc[0] ),
    .B(net3404));
 sg13g2_xor2_1 _08390_ (.B(net3404),
    .A(\u_toplayer.u_outlayer.u_neuron.acc[0] ),
    .X(_02348_));
 sg13g2_nand2_1 _08391_ (.Y(_02349_),
    .A(\u_toplayer.u_outlayer.u_neuron.acc[0] ),
    .B(net1212));
 sg13g2_xor2_1 _08392_ (.B(net901),
    .A(\u_toplayer.u_outlayer.u_neuron.acc[0] ),
    .X(_02350_));
 sg13g2_a22oi_1 _08393_ (.Y(_02351_),
    .B1(_02350_),
    .B2(net2977),
    .A2(_02348_),
    .A1(net2934));
 sg13g2_a21oi_1 _08394_ (.A1(net2891),
    .A2(_02351_),
    .Y(_00197_),
    .B1(_02344_));
 sg13g2_nand2_1 _08395_ (.Y(_02352_),
    .A(net3201),
    .B(\u_toplayer.u_outlayer.u_neuron.mult[1] ));
 sg13g2_nor2_1 _08396_ (.A(net3201),
    .B(\u_toplayer.u_outlayer.u_neuron.mult[1] ),
    .Y(_02353_));
 sg13g2_xor2_1 _08397_ (.B(\u_toplayer.u_outlayer.u_neuron.mult[1] ),
    .A(net3201),
    .X(_02354_));
 sg13g2_xnor2_1 _08398_ (.Y(_02355_),
    .A(_02349_),
    .B(_02354_));
 sg13g2_nand2_1 _08399_ (.Y(_02356_),
    .A(net3201),
    .B(net3400));
 sg13g2_nor2_1 _08400_ (.A(net3201),
    .B(net3400),
    .Y(_02357_));
 sg13g2_xor2_1 _08401_ (.B(net3400),
    .A(net3201),
    .X(_02358_));
 sg13g2_xnor2_1 _08402_ (.Y(_02359_),
    .A(_02347_),
    .B(_02358_));
 sg13g2_a22oi_1 _08403_ (.Y(_02360_),
    .B1(_02359_),
    .B2(net2934),
    .A2(_02355_),
    .A1(net2977));
 sg13g2_nor2_1 _08404_ (.A(net822),
    .B(net2891),
    .Y(_02361_));
 sg13g2_a21oi_1 _08405_ (.A1(net2891),
    .A2(_02360_),
    .Y(_00198_),
    .B1(_02361_));
 sg13g2_and2_1 _08406_ (.A(\u_toplayer.u_outlayer.u_neuron.acc[2] ),
    .B(\u_toplayer.u_outlayer.u_neuron.mult[2] ),
    .X(_02362_));
 sg13g2_xor2_1 _08407_ (.B(\u_toplayer.u_outlayer.u_neuron.mult[2] ),
    .A(\u_toplayer.u_outlayer.u_neuron.acc[2] ),
    .X(_02363_));
 sg13g2_o21ai_1 _08408_ (.B1(_02352_),
    .Y(_02364_),
    .A1(_02349_),
    .A2(_02353_));
 sg13g2_nand2_1 _08409_ (.Y(_02365_),
    .A(_02363_),
    .B(_02364_));
 sg13g2_o21ai_1 _08410_ (.B1(net2977),
    .Y(_02366_),
    .A1(_02363_),
    .A2(_02364_));
 sg13g2_inv_1 _08411_ (.Y(_02367_),
    .A(_02366_));
 sg13g2_and2_1 _08412_ (.A(\u_toplayer.u_outlayer.u_neuron.acc[2] ),
    .B(net3396),
    .X(_02368_));
 sg13g2_xor2_1 _08413_ (.B(net3396),
    .A(\u_toplayer.u_outlayer.u_neuron.acc[2] ),
    .X(_02369_));
 sg13g2_o21ai_1 _08414_ (.B1(_02356_),
    .Y(_02370_),
    .A1(_02347_),
    .A2(_02357_));
 sg13g2_o21ai_1 _08415_ (.B1(net2934),
    .Y(_02371_),
    .A1(_02369_),
    .A2(_02370_));
 sg13g2_a21oi_1 _08416_ (.A1(_02369_),
    .A2(_02370_),
    .Y(_02372_),
    .B1(_02371_));
 sg13g2_a21oi_1 _08417_ (.A1(_02365_),
    .A2(_02367_),
    .Y(_02373_),
    .B1(_02372_));
 sg13g2_nor2_1 _08418_ (.A(net1116),
    .B(net2891),
    .Y(_02374_));
 sg13g2_a21oi_1 _08419_ (.A1(net2891),
    .A2(_02373_),
    .Y(_00199_),
    .B1(_02374_));
 sg13g2_nand2_1 _08420_ (.Y(_02375_),
    .A(\u_toplayer.u_outlayer.u_neuron.acc[3] ),
    .B(\u_toplayer.u_outlayer.u_neuron.mult[3] ));
 sg13g2_xnor2_1 _08421_ (.Y(_02376_),
    .A(\u_toplayer.u_outlayer.u_neuron.acc[3] ),
    .B(\u_toplayer.u_outlayer.u_neuron.mult[3] ));
 sg13g2_a21oi_1 _08422_ (.A1(_02363_),
    .A2(_02364_),
    .Y(_02377_),
    .B1(_02362_));
 sg13g2_xnor2_1 _08423_ (.Y(_02378_),
    .A(_02376_),
    .B(_02377_));
 sg13g2_nand2_1 _08424_ (.Y(_02379_),
    .A(\u_toplayer.u_outlayer.u_neuron.acc[3] ),
    .B(net3393));
 sg13g2_xnor2_1 _08425_ (.Y(_02380_),
    .A(\u_toplayer.u_outlayer.u_neuron.acc[3] ),
    .B(net3393));
 sg13g2_a21oi_2 _08426_ (.B1(_02368_),
    .Y(_02381_),
    .A2(_02370_),
    .A1(_02369_));
 sg13g2_a21oi_1 _08427_ (.A1(_02380_),
    .A2(_02381_),
    .Y(_02382_),
    .B1(_02346_));
 sg13g2_o21ai_1 _08428_ (.B1(_02382_),
    .Y(_02383_),
    .A1(_02380_),
    .A2(_02381_));
 sg13g2_o21ai_1 _08429_ (.B1(_02383_),
    .Y(_02384_),
    .A1(net2979),
    .A2(_02378_));
 sg13g2_mux2_1 _08430_ (.A0(net1100),
    .A1(_02384_),
    .S(net2891),
    .X(_00200_));
 sg13g2_and2_1 _08431_ (.A(\u_toplayer.u_outlayer.u_neuron.acc[4] ),
    .B(\u_toplayer.u_outlayer.u_neuron.mult[4] ),
    .X(_02385_));
 sg13g2_xor2_1 _08432_ (.B(\u_toplayer.u_outlayer.u_neuron.mult[4] ),
    .A(\u_toplayer.u_outlayer.u_neuron.acc[4] ),
    .X(_02386_));
 sg13g2_o21ai_1 _08433_ (.B1(_02375_),
    .Y(_02387_),
    .A1(_02376_),
    .A2(_02377_));
 sg13g2_or2_1 _08434_ (.X(_02388_),
    .B(_02387_),
    .A(_02386_));
 sg13g2_a21oi_1 _08435_ (.A1(_02386_),
    .A2(_02387_),
    .Y(_02389_),
    .B1(_01389_));
 sg13g2_nor2_1 _08436_ (.A(_01039_),
    .B(_01046_),
    .Y(_02390_));
 sg13g2_xor2_1 _08437_ (.B(net3390),
    .A(\u_toplayer.u_outlayer.u_neuron.acc[4] ),
    .X(_02391_));
 sg13g2_o21ai_1 _08438_ (.B1(_02379_),
    .Y(_02392_),
    .A1(_02380_),
    .A2(_02381_));
 sg13g2_o21ai_1 _08439_ (.B1(net2934),
    .Y(_02393_),
    .A1(_02391_),
    .A2(_02392_));
 sg13g2_a21o_1 _08440_ (.A2(_02392_),
    .A1(_02391_),
    .B1(_02393_),
    .X(_02394_));
 sg13g2_a21oi_1 _08441_ (.A1(_02388_),
    .A2(_02389_),
    .Y(_02395_),
    .B1(net2893));
 sg13g2_a22oi_1 _08442_ (.Y(_00201_),
    .B1(_02394_),
    .B2(_02395_),
    .A2(_02342_),
    .A1(_01039_));
 sg13g2_nor2_1 _08443_ (.A(net3200),
    .B(net2891),
    .Y(_02396_));
 sg13g2_a21oi_1 _08444_ (.A1(_02391_),
    .A2(_02392_),
    .Y(_02397_),
    .B1(_02390_));
 sg13g2_nor2_1 _08445_ (.A(net3200),
    .B(net3387),
    .Y(_02398_));
 sg13g2_xor2_1 _08446_ (.B(net3387),
    .A(net3200),
    .X(_02399_));
 sg13g2_xnor2_1 _08447_ (.Y(_02400_),
    .A(_02397_),
    .B(_02399_));
 sg13g2_a21oi_1 _08448_ (.A1(_02386_),
    .A2(_02387_),
    .Y(_02401_),
    .B1(_02385_));
 sg13g2_nor2_1 _08449_ (.A(net3200),
    .B(\u_toplayer.u_outlayer.u_neuron.mult[5] ),
    .Y(_02402_));
 sg13g2_xor2_1 _08450_ (.B(\u_toplayer.u_outlayer.u_neuron.mult[5] ),
    .A(net3200),
    .X(_02403_));
 sg13g2_xnor2_1 _08451_ (.Y(_02404_),
    .A(_02401_),
    .B(_02403_));
 sg13g2_a22oi_1 _08452_ (.Y(_02405_),
    .B1(_02404_),
    .B2(net2977),
    .A2(_02400_),
    .A1(net2934));
 sg13g2_a21oi_1 _08453_ (.A1(net2891),
    .A2(_02405_),
    .Y(_00202_),
    .B1(_02396_));
 sg13g2_nand2_1 _08454_ (.Y(_02406_),
    .A(\u_toplayer.u_outlayer.u_neuron.acc[6] ),
    .B(\u_toplayer.u_outlayer.u_neuron.mult[6] ));
 sg13g2_xnor2_1 _08455_ (.Y(_02407_),
    .A(\u_toplayer.u_outlayer.u_neuron.acc[6] ),
    .B(\u_toplayer.u_outlayer.u_neuron.mult[6] ));
 sg13g2_a221oi_1 _08456_ (.B2(_02387_),
    .C1(_02385_),
    .B1(_02386_),
    .A1(net3200),
    .Y(_02408_),
    .A2(\u_toplayer.u_outlayer.u_neuron.mult[5] ));
 sg13g2_o21ai_1 _08457_ (.B1(_02407_),
    .Y(_02409_),
    .A1(_02402_),
    .A2(_02408_));
 sg13g2_or3_1 _08458_ (.A(_02402_),
    .B(_02407_),
    .C(_02408_),
    .X(_02410_));
 sg13g2_nand3_1 _08459_ (.B(_02409_),
    .C(_02410_),
    .A(net2977),
    .Y(_02411_));
 sg13g2_and2_1 _08460_ (.A(\u_toplayer.u_outlayer.u_neuron.acc[6] ),
    .B(net1),
    .X(_02412_));
 sg13g2_xnor2_1 _08461_ (.Y(_02413_),
    .A(\u_toplayer.u_outlayer.u_neuron.acc[6] ),
    .B(net1));
 sg13g2_a221oi_1 _08462_ (.B2(_02392_),
    .C1(_02390_),
    .B1(_02391_),
    .A1(net3200),
    .Y(_02414_),
    .A2(net3387));
 sg13g2_o21ai_1 _08463_ (.B1(_02413_),
    .Y(_02415_),
    .A1(_02398_),
    .A2(_02414_));
 sg13g2_nor3_2 _08464_ (.A(_02398_),
    .B(_02413_),
    .C(_02414_),
    .Y(_02416_));
 sg13g2_nor2_1 _08465_ (.A(_02346_),
    .B(_02416_),
    .Y(_02417_));
 sg13g2_a21oi_1 _08466_ (.A1(_02415_),
    .A2(_02417_),
    .Y(_02418_),
    .B1(net2893));
 sg13g2_a22oi_1 _08467_ (.Y(_00203_),
    .B1(_02411_),
    .B2(_02418_),
    .A2(net2893),
    .A1(_01038_));
 sg13g2_nand2_1 _08468_ (.Y(_02419_),
    .A(\u_toplayer.u_outlayer.u_neuron.acc[7] ),
    .B(net3362));
 sg13g2_xor2_1 _08469_ (.B(net3362),
    .A(\u_toplayer.u_outlayer.u_neuron.acc[7] ),
    .X(_02420_));
 sg13g2_nor3_1 _08470_ (.A(_02412_),
    .B(_02416_),
    .C(_02420_),
    .Y(_02421_));
 sg13g2_o21ai_1 _08471_ (.B1(_02420_),
    .Y(_02422_),
    .A1(_02412_),
    .A2(_02416_));
 sg13g2_nor2_1 _08472_ (.A(_02346_),
    .B(_02421_),
    .Y(_02423_));
 sg13g2_nand2_1 _08473_ (.Y(_02424_),
    .A(\u_toplayer.u_outlayer.u_neuron.acc[7] ),
    .B(\u_toplayer.u_outlayer.u_neuron.mult[7] ));
 sg13g2_xnor2_1 _08474_ (.Y(_02425_),
    .A(\u_toplayer.u_outlayer.u_neuron.acc[7] ),
    .B(\u_toplayer.u_outlayer.u_neuron.mult[7] ));
 sg13g2_a21o_1 _08475_ (.A2(_02410_),
    .A1(_02406_),
    .B1(_02425_),
    .X(_02426_));
 sg13g2_nand3_1 _08476_ (.B(_02410_),
    .C(_02425_),
    .A(_02406_),
    .Y(_02427_));
 sg13g2_nand3_1 _08477_ (.B(_02426_),
    .C(_02427_),
    .A(net2976),
    .Y(_02428_));
 sg13g2_a21oi_1 _08478_ (.A1(_02422_),
    .A2(_02423_),
    .Y(_02429_),
    .B1(net2893));
 sg13g2_a22oi_1 _08479_ (.Y(_00204_),
    .B1(_02428_),
    .B2(_02429_),
    .A2(net2893),
    .A1(_01037_));
 sg13g2_nor2_1 _08480_ (.A(net1140),
    .B(net2888),
    .Y(_02430_));
 sg13g2_nand2_1 _08481_ (.Y(_02431_),
    .A(_02419_),
    .B(_02422_));
 sg13g2_nand2_1 _08482_ (.Y(_02432_),
    .A(\u_toplayer.u_outlayer.u_neuron.acc[8] ),
    .B(net3357));
 sg13g2_xor2_1 _08483_ (.B(net3357),
    .A(\u_toplayer.u_outlayer.u_neuron.acc[8] ),
    .X(_02433_));
 sg13g2_inv_1 _08484_ (.Y(_02434_),
    .A(_02433_));
 sg13g2_nor2_1 _08485_ (.A(_02431_),
    .B(_02433_),
    .Y(_02435_));
 sg13g2_nand2_1 _08486_ (.Y(_02436_),
    .A(_02431_),
    .B(_02433_));
 sg13g2_nor2_1 _08487_ (.A(net2932),
    .B(_02435_),
    .Y(_02437_));
 sg13g2_and2_1 _08488_ (.A(\u_toplayer.u_outlayer.u_neuron.acc[8] ),
    .B(\u_toplayer.u_outlayer.u_neuron.mult[8] ),
    .X(_02438_));
 sg13g2_xnor2_1 _08489_ (.Y(_02439_),
    .A(\u_toplayer.u_outlayer.u_neuron.acc[8] ),
    .B(\u_toplayer.u_outlayer.u_neuron.mult[8] ));
 sg13g2_a21oi_2 _08490_ (.B1(_02439_),
    .Y(_02440_),
    .A2(_02426_),
    .A1(_02424_));
 sg13g2_nand3_1 _08491_ (.B(_02426_),
    .C(_02439_),
    .A(_02424_),
    .Y(_02441_));
 sg13g2_nor2b_1 _08492_ (.A(_02440_),
    .B_N(_02441_),
    .Y(_02442_));
 sg13g2_a22oi_1 _08493_ (.Y(_02443_),
    .B1(_02442_),
    .B2(net2976),
    .A2(_02437_),
    .A1(_02436_));
 sg13g2_a21oi_1 _08494_ (.A1(net2888),
    .A2(_02443_),
    .Y(_00205_),
    .B1(_02430_));
 sg13g2_nor2_1 _08495_ (.A(net3199),
    .B(net2888),
    .Y(_02444_));
 sg13g2_nor2_1 _08496_ (.A(net3199),
    .B(\u_toplayer.u_outlayer.u_neuron.mult[9] ),
    .Y(_02445_));
 sg13g2_xnor2_1 _08497_ (.Y(_02446_),
    .A(\u_toplayer.u_outlayer.u_neuron.acc[9] ),
    .B(\u_toplayer.u_outlayer.u_neuron.mult[9] ));
 sg13g2_nor2_1 _08498_ (.A(_02438_),
    .B(_02440_),
    .Y(_02447_));
 sg13g2_xor2_1 _08499_ (.B(_02447_),
    .A(_02446_),
    .X(_02448_));
 sg13g2_xnor2_1 _08500_ (.Y(_02449_),
    .A(net3199),
    .B(net3357));
 sg13g2_and2_1 _08501_ (.A(_02432_),
    .B(_02436_),
    .X(_02450_));
 sg13g2_o21ai_1 _08502_ (.B1(net2933),
    .Y(_02451_),
    .A1(_02449_),
    .A2(_02450_));
 sg13g2_a21oi_1 _08503_ (.A1(_02449_),
    .A2(_02450_),
    .Y(_02452_),
    .B1(_02451_));
 sg13g2_a21oi_1 _08504_ (.A1(net2976),
    .A2(_02448_),
    .Y(_02453_),
    .B1(_02452_));
 sg13g2_a21oi_1 _08505_ (.A1(net2888),
    .A2(_02453_),
    .Y(_00206_),
    .B1(_02444_));
 sg13g2_nor2_1 _08506_ (.A(net1127),
    .B(net2890),
    .Y(_02454_));
 sg13g2_nand2_1 _08507_ (.Y(_02455_),
    .A(\u_toplayer.u_outlayer.u_neuron.acc[10] ),
    .B(net3357));
 sg13g2_xnor2_1 _08508_ (.Y(_02456_),
    .A(\u_toplayer.u_outlayer.u_neuron.acc[10] ),
    .B(net3357));
 sg13g2_o21ai_1 _08509_ (.B1(net3357),
    .Y(_02457_),
    .A1(net3199),
    .A2(\u_toplayer.u_outlayer.u_neuron.acc[8] ));
 sg13g2_nand2_1 _08510_ (.Y(_02458_),
    .A(_02436_),
    .B(_02457_));
 sg13g2_o21ai_1 _08511_ (.B1(_02458_),
    .Y(_02459_),
    .A1(net3199),
    .A2(net3357));
 sg13g2_or2_1 _08512_ (.X(_02460_),
    .B(_02459_),
    .A(_02456_));
 sg13g2_a21oi_1 _08513_ (.A1(_02456_),
    .A2(_02459_),
    .Y(_02461_),
    .B1(net2932));
 sg13g2_nand2_1 _08514_ (.Y(_02462_),
    .A(\u_toplayer.u_outlayer.u_neuron.acc[10] ),
    .B(\u_toplayer.u_outlayer.u_neuron.mult[10] ));
 sg13g2_xnor2_1 _08515_ (.Y(_02463_),
    .A(\u_toplayer.u_outlayer.u_neuron.acc[10] ),
    .B(\u_toplayer.u_outlayer.u_neuron.mult[10] ));
 sg13g2_a21o_1 _08516_ (.A2(\u_toplayer.u_outlayer.u_neuron.mult[9] ),
    .A1(net3199),
    .B1(_02438_),
    .X(_02464_));
 sg13g2_nor2_1 _08517_ (.A(_02440_),
    .B(_02464_),
    .Y(_02465_));
 sg13g2_or2_1 _08518_ (.X(_02466_),
    .B(_02465_),
    .A(_02445_));
 sg13g2_or2_1 _08519_ (.X(_02467_),
    .B(_02466_),
    .A(_02463_));
 sg13g2_a21oi_1 _08520_ (.A1(_02463_),
    .A2(_02466_),
    .Y(_02468_),
    .B1(net2979));
 sg13g2_a22oi_1 _08521_ (.Y(_02469_),
    .B1(_02467_),
    .B2(_02468_),
    .A2(_02461_),
    .A1(_02460_));
 sg13g2_a21oi_1 _08522_ (.A1(net2890),
    .A2(_02469_),
    .Y(_00207_),
    .B1(_02454_));
 sg13g2_xnor2_1 _08523_ (.Y(_02470_),
    .A(\u_toplayer.u_outlayer.u_neuron.acc[11] ),
    .B(net3363));
 sg13g2_and2_1 _08524_ (.A(_02455_),
    .B(_02460_),
    .X(_02471_));
 sg13g2_a21oi_1 _08525_ (.A1(_02470_),
    .A2(_02471_),
    .Y(_02472_),
    .B1(net2932));
 sg13g2_o21ai_1 _08526_ (.B1(_02472_),
    .Y(_02473_),
    .A1(_02470_),
    .A2(_02471_));
 sg13g2_nor2_1 _08527_ (.A(\u_toplayer.u_outlayer.u_neuron.acc[11] ),
    .B(\u_toplayer.u_outlayer.u_neuron.mult[11] ),
    .Y(_02474_));
 sg13g2_nand2_1 _08528_ (.Y(_02475_),
    .A(\u_toplayer.u_outlayer.u_neuron.acc[11] ),
    .B(\u_toplayer.u_outlayer.u_neuron.mult[11] ));
 sg13g2_nand2b_1 _08529_ (.Y(_02476_),
    .B(_02475_),
    .A_N(_02474_));
 sg13g2_nand3_1 _08530_ (.B(_02467_),
    .C(_02476_),
    .A(_02462_),
    .Y(_02477_));
 sg13g2_a21oi_1 _08531_ (.A1(_02462_),
    .A2(_02467_),
    .Y(_02478_),
    .B1(_02476_));
 sg13g2_nor2_1 _08532_ (.A(_01389_),
    .B(_02478_),
    .Y(_02479_));
 sg13g2_a21oi_1 _08533_ (.A1(_02477_),
    .A2(_02479_),
    .Y(_02480_),
    .B1(_02342_));
 sg13g2_a22oi_1 _08534_ (.Y(_00208_),
    .B1(_02473_),
    .B2(_02480_),
    .A2(_02342_),
    .A1(_01042_));
 sg13g2_nand2_1 _08535_ (.Y(_02481_),
    .A(\u_toplayer.u_outlayer.u_neuron.acc[12] ),
    .B(net3359));
 sg13g2_xnor2_1 _08536_ (.Y(_02482_),
    .A(\u_toplayer.u_outlayer.u_neuron.acc[12] ),
    .B(net3363));
 sg13g2_or4_1 _08537_ (.A(_02434_),
    .B(_02449_),
    .C(_02456_),
    .D(_02470_),
    .X(_02483_));
 sg13g2_a21oi_1 _08538_ (.A1(_02419_),
    .A2(_02422_),
    .Y(_02484_),
    .B1(_02483_));
 sg13g2_nand2b_1 _08539_ (.Y(_02485_),
    .B(_02431_),
    .A_N(_02483_));
 sg13g2_o21ai_1 _08540_ (.B1(net3357),
    .Y(_02486_),
    .A1(\u_toplayer.u_outlayer.u_neuron.acc[11] ),
    .A2(\u_toplayer.u_outlayer.u_neuron.acc[10] ));
 sg13g2_and2_1 _08541_ (.A(_02457_),
    .B(_02486_),
    .X(_02487_));
 sg13g2_nand3_1 _08542_ (.B(_02485_),
    .C(_02487_),
    .A(_02482_),
    .Y(_02488_));
 sg13g2_a21o_1 _08543_ (.A2(_02487_),
    .A1(_02485_),
    .B1(_02482_),
    .X(_02489_));
 sg13g2_nand3_1 _08544_ (.B(_02488_),
    .C(_02489_),
    .A(net2933),
    .Y(_02490_));
 sg13g2_nor3_1 _08545_ (.A(_02446_),
    .B(_02463_),
    .C(_02476_),
    .Y(_02491_));
 sg13g2_nor3_1 _08546_ (.A(_02445_),
    .B(_02463_),
    .C(_02476_),
    .Y(_02492_));
 sg13g2_o21ai_1 _08547_ (.B1(_02475_),
    .Y(_02493_),
    .A1(_02462_),
    .A2(_02474_));
 sg13g2_a221oi_1 _08548_ (.B2(_02464_),
    .C1(_02493_),
    .B1(_02492_),
    .A1(_02440_),
    .Y(_02494_),
    .A2(_02491_));
 sg13g2_xnor2_1 _08549_ (.Y(_02495_),
    .A(\u_toplayer.u_outlayer.u_neuron.acc[12] ),
    .B(\u_toplayer.u_outlayer.u_neuron.mult[12] ));
 sg13g2_or2_1 _08550_ (.X(_02496_),
    .B(_02495_),
    .A(_02494_));
 sg13g2_a21oi_1 _08551_ (.A1(_02494_),
    .A2(_02495_),
    .Y(_02497_),
    .B1(net2979));
 sg13g2_a21oi_1 _08552_ (.A1(_02496_),
    .A2(_02497_),
    .Y(_02498_),
    .B1(net2892));
 sg13g2_a22oi_1 _08553_ (.Y(_00209_),
    .B1(_02490_),
    .B2(_02498_),
    .A2(net2892),
    .A1(_01041_));
 sg13g2_nor2_1 _08554_ (.A(net3198),
    .B(net2888),
    .Y(_02499_));
 sg13g2_nor2_1 _08555_ (.A(net3198),
    .B(net3358),
    .Y(_02500_));
 sg13g2_xor2_1 _08556_ (.B(net3358),
    .A(net3198),
    .X(_02501_));
 sg13g2_nand2_1 _08557_ (.Y(_02502_),
    .A(_02481_),
    .B(_02489_));
 sg13g2_xor2_1 _08558_ (.B(_02502_),
    .A(_02501_),
    .X(_02503_));
 sg13g2_nor2_1 _08559_ (.A(net3198),
    .B(\u_toplayer.u_outlayer.u_neuron.mult[13] ),
    .Y(_02504_));
 sg13g2_xnor2_1 _08560_ (.Y(_02505_),
    .A(net3198),
    .B(\u_toplayer.u_outlayer.u_neuron.mult[13] ));
 sg13g2_o21ai_1 _08561_ (.B1(_02496_),
    .Y(_02506_),
    .A1(_01041_),
    .A2(_01048_));
 sg13g2_xnor2_1 _08562_ (.Y(_02507_),
    .A(_02505_),
    .B(_02506_));
 sg13g2_a22oi_1 _08563_ (.Y(_02508_),
    .B1(_02507_),
    .B2(net2976),
    .A2(_02503_),
    .A1(net2933));
 sg13g2_a21oi_1 _08564_ (.A1(net2888),
    .A2(_02508_),
    .Y(_00210_),
    .B1(_02499_));
 sg13g2_nand2_1 _08565_ (.Y(_02509_),
    .A(\u_toplayer.u_outlayer.u_neuron.acc[14] ),
    .B(net3358));
 sg13g2_xnor2_1 _08566_ (.Y(_02510_),
    .A(\u_toplayer.u_outlayer.u_neuron.acc[14] ),
    .B(net3358));
 sg13g2_a21oi_1 _08567_ (.A1(net3198),
    .A2(net3358),
    .Y(_02511_),
    .B1(_02502_));
 sg13g2_o21ai_1 _08568_ (.B1(_02510_),
    .Y(_02512_),
    .A1(_02500_),
    .A2(_02511_));
 sg13g2_or3_1 _08569_ (.A(_02500_),
    .B(_02510_),
    .C(_02511_),
    .X(_02513_));
 sg13g2_nand3_1 _08570_ (.B(_02512_),
    .C(_02513_),
    .A(net2933),
    .Y(_02514_));
 sg13g2_nand2_1 _08571_ (.Y(_02515_),
    .A(\u_toplayer.u_outlayer.u_neuron.acc[14] ),
    .B(\u_toplayer.u_outlayer.u_neuron.mult[14] ));
 sg13g2_xnor2_1 _08572_ (.Y(_02516_),
    .A(\u_toplayer.u_outlayer.u_neuron.acc[14] ),
    .B(\u_toplayer.u_outlayer.u_neuron.mult[14] ));
 sg13g2_a22oi_1 _08573_ (.Y(_02517_),
    .B1(\u_toplayer.u_outlayer.u_neuron.mult[13] ),
    .B2(net3198),
    .A2(\u_toplayer.u_outlayer.u_neuron.mult[12] ),
    .A1(\u_toplayer.u_outlayer.u_neuron.acc[12] ));
 sg13g2_a21oi_1 _08574_ (.A1(_02496_),
    .A2(_02517_),
    .Y(_02518_),
    .B1(_02504_));
 sg13g2_nand2b_1 _08575_ (.Y(_02519_),
    .B(_02518_),
    .A_N(_02516_));
 sg13g2_xnor2_1 _08576_ (.Y(_02520_),
    .A(_02516_),
    .B(_02518_));
 sg13g2_a21oi_1 _08577_ (.A1(net2976),
    .A2(_02520_),
    .Y(_02521_),
    .B1(net2892));
 sg13g2_a22oi_1 _08578_ (.Y(_00211_),
    .B1(_02514_),
    .B2(_02521_),
    .A2(net2892),
    .A1(_01040_));
 sg13g2_nor2_1 _08579_ (.A(net1058),
    .B(net2888),
    .Y(_02522_));
 sg13g2_xnor2_1 _08580_ (.Y(_02523_),
    .A(\u_toplayer.u_outlayer.u_neuron.acc[15] ),
    .B(net3358));
 sg13g2_a21oi_1 _08581_ (.A1(_02509_),
    .A2(_02513_),
    .Y(_02524_),
    .B1(_02523_));
 sg13g2_nand3_1 _08582_ (.B(_02513_),
    .C(_02523_),
    .A(_02509_),
    .Y(_02525_));
 sg13g2_nor2_1 _08583_ (.A(net2932),
    .B(_02524_),
    .Y(_02526_));
 sg13g2_nor2_1 _08584_ (.A(\u_toplayer.u_outlayer.u_neuron.acc[15] ),
    .B(net3226),
    .Y(_02527_));
 sg13g2_nand2_1 _08585_ (.Y(_02528_),
    .A(\u_toplayer.u_outlayer.u_neuron.acc[15] ),
    .B(net3226));
 sg13g2_nand2b_1 _08586_ (.Y(_02529_),
    .B(_02528_),
    .A_N(_02527_));
 sg13g2_and2_1 _08587_ (.A(_02515_),
    .B(_02519_),
    .X(_02530_));
 sg13g2_o21ai_1 _08588_ (.B1(net2976),
    .Y(_02531_),
    .A1(_02529_),
    .A2(_02530_));
 sg13g2_a21oi_1 _08589_ (.A1(_02529_),
    .A2(_02530_),
    .Y(_02532_),
    .B1(_02531_));
 sg13g2_a21oi_1 _08590_ (.A1(_02525_),
    .A2(_02526_),
    .Y(_02533_),
    .B1(_02532_));
 sg13g2_a21oi_1 _08591_ (.A1(net2888),
    .A2(_02533_),
    .Y(_00212_),
    .B1(_02522_));
 sg13g2_or4_1 _08592_ (.A(_02495_),
    .B(_02505_),
    .C(_02516_),
    .D(_02529_),
    .X(_02534_));
 sg13g2_o21ai_1 _08593_ (.B1(_02528_),
    .Y(_02535_),
    .A1(_02515_),
    .A2(_02527_));
 sg13g2_nor4_1 _08594_ (.A(_02504_),
    .B(_02516_),
    .C(_02517_),
    .D(_02529_),
    .Y(_02536_));
 sg13g2_nor2_1 _08595_ (.A(_02535_),
    .B(_02536_),
    .Y(_02537_));
 sg13g2_o21ai_1 _08596_ (.B1(_02537_),
    .Y(_02538_),
    .A1(_02494_),
    .A2(_02534_));
 sg13g2_xnor2_1 _08597_ (.Y(_02539_),
    .A(net3197),
    .B(net3227));
 sg13g2_inv_1 _08598_ (.Y(_02540_),
    .A(_02539_));
 sg13g2_and2_1 _08599_ (.A(_02538_),
    .B(_02540_),
    .X(_02541_));
 sg13g2_o21ai_1 _08600_ (.B1(net2978),
    .Y(_02542_),
    .A1(_02538_),
    .A2(_02540_));
 sg13g2_nand2b_1 _08601_ (.Y(_02543_),
    .B(_02501_),
    .A_N(_02482_));
 sg13g2_nor3_1 _08602_ (.A(_02510_),
    .B(_02523_),
    .C(_02543_),
    .Y(_02544_));
 sg13g2_o21ai_1 _08603_ (.B1(net3358),
    .Y(_02545_),
    .A1(\u_toplayer.u_outlayer.u_neuron.acc[15] ),
    .A2(\u_toplayer.u_outlayer.u_neuron.acc[14] ));
 sg13g2_nand3_1 _08604_ (.B(_02487_),
    .C(_02545_),
    .A(_02481_),
    .Y(_02546_));
 sg13g2_a221oi_1 _08605_ (.B2(_02544_),
    .C1(_02546_),
    .B1(_02484_),
    .A1(net3198),
    .Y(_02547_),
    .A2(net3358));
 sg13g2_nand2_1 _08606_ (.Y(_02548_),
    .A(net3197),
    .B(net3360));
 sg13g2_xnor2_1 _08607_ (.Y(_02549_),
    .A(net3197),
    .B(net3360));
 sg13g2_a21oi_1 _08608_ (.A1(_02547_),
    .A2(_02549_),
    .Y(_02550_),
    .B1(net2932));
 sg13g2_o21ai_1 _08609_ (.B1(_02550_),
    .Y(_02551_),
    .A1(_02547_),
    .A2(_02549_));
 sg13g2_o21ai_1 _08610_ (.B1(_02551_),
    .Y(_02552_),
    .A1(_02541_),
    .A2(_02542_));
 sg13g2_mux2_1 _08611_ (.A0(net823),
    .A1(_02552_),
    .S(net2889),
    .X(_00213_));
 sg13g2_nor2_1 _08612_ (.A(net1079),
    .B(net2889),
    .Y(_02553_));
 sg13g2_xor2_1 _08613_ (.B(net3227),
    .A(\u_toplayer.u_outlayer.u_neuron.acc[17] ),
    .X(_02554_));
 sg13g2_a21oi_1 _08614_ (.A1(net3197),
    .A2(net3227),
    .Y(_02555_),
    .B1(_02541_));
 sg13g2_xnor2_1 _08615_ (.Y(_02556_),
    .A(_02554_),
    .B(_02555_));
 sg13g2_xnor2_1 _08616_ (.Y(_02557_),
    .A(\u_toplayer.u_outlayer.u_neuron.acc[17] ),
    .B(net3360));
 sg13g2_o21ai_1 _08617_ (.B1(_02548_),
    .Y(_02558_),
    .A1(_02547_),
    .A2(_02549_));
 sg13g2_xnor2_1 _08618_ (.Y(_02559_),
    .A(_02557_),
    .B(_02558_));
 sg13g2_a22oi_1 _08619_ (.Y(_02560_),
    .B1(_02559_),
    .B2(net2933),
    .A2(_02556_),
    .A1(net2978));
 sg13g2_a21oi_1 _08620_ (.A1(net2889),
    .A2(_02560_),
    .Y(_00214_),
    .B1(_02553_));
 sg13g2_nor2_1 _08621_ (.A(net3196),
    .B(net2889),
    .Y(_02561_));
 sg13g2_nand2_1 _08622_ (.Y(_02562_),
    .A(net3196),
    .B(net3226));
 sg13g2_xnor2_1 _08623_ (.Y(_02563_),
    .A(\u_toplayer.u_outlayer.u_neuron.acc[18] ),
    .B(net3227));
 sg13g2_o21ai_1 _08624_ (.B1(net3227),
    .Y(_02564_),
    .A1(\u_toplayer.u_outlayer.u_neuron.acc[17] ),
    .A2(net3197));
 sg13g2_inv_1 _08625_ (.Y(_02565_),
    .A(_02564_));
 sg13g2_a21oi_1 _08626_ (.A1(_02541_),
    .A2(_02554_),
    .Y(_02566_),
    .B1(_02565_));
 sg13g2_or2_1 _08627_ (.X(_02567_),
    .B(_02566_),
    .A(_02563_));
 sg13g2_a21oi_1 _08628_ (.A1(_02563_),
    .A2(_02566_),
    .Y(_02568_),
    .B1(net2979));
 sg13g2_xnor2_1 _08629_ (.Y(_02569_),
    .A(net3196),
    .B(net3360));
 sg13g2_or2_1 _08630_ (.X(_02570_),
    .B(_02557_),
    .A(_02549_));
 sg13g2_or2_1 _08631_ (.X(_02571_),
    .B(_02570_),
    .A(_02547_));
 sg13g2_o21ai_1 _08632_ (.B1(net3361),
    .Y(_02572_),
    .A1(\u_toplayer.u_outlayer.u_neuron.acc[17] ),
    .A2(net3197));
 sg13g2_a21oi_1 _08633_ (.A1(_02571_),
    .A2(_02572_),
    .Y(_02573_),
    .B1(_02569_));
 sg13g2_nand3_1 _08634_ (.B(_02571_),
    .C(_02572_),
    .A(_02569_),
    .Y(_02574_));
 sg13g2_nor2_1 _08635_ (.A(net2932),
    .B(_02573_),
    .Y(_02575_));
 sg13g2_a22oi_1 _08636_ (.Y(_02576_),
    .B1(_02574_),
    .B2(_02575_),
    .A2(_02568_),
    .A1(_02567_));
 sg13g2_a21oi_1 _08637_ (.A1(net2889),
    .A2(_02576_),
    .Y(_00215_),
    .B1(_02561_));
 sg13g2_nor2_1 _08638_ (.A(net1067),
    .B(net2889),
    .Y(_02577_));
 sg13g2_xnor2_1 _08639_ (.Y(_02578_),
    .A(\u_toplayer.u_outlayer.u_neuron.acc[19] ),
    .B(net3226));
 sg13g2_nand2_1 _08640_ (.Y(_02579_),
    .A(_02562_),
    .B(_02567_));
 sg13g2_xnor2_1 _08641_ (.Y(_02580_),
    .A(_02578_),
    .B(_02579_));
 sg13g2_xnor2_1 _08642_ (.Y(_02581_),
    .A(\u_toplayer.u_outlayer.u_neuron.acc[19] ),
    .B(net3360));
 sg13g2_a21oi_1 _08643_ (.A1(net3196),
    .A2(net3360),
    .Y(_02582_),
    .B1(_02573_));
 sg13g2_o21ai_1 _08644_ (.B1(net2933),
    .Y(_02583_),
    .A1(_02581_),
    .A2(_02582_));
 sg13g2_a21oi_1 _08645_ (.A1(_02581_),
    .A2(_02582_),
    .Y(_02584_),
    .B1(_02583_));
 sg13g2_a21oi_1 _08646_ (.A1(net2978),
    .A2(_02580_),
    .Y(_02585_),
    .B1(_02584_));
 sg13g2_a21oi_1 _08647_ (.A1(net2889),
    .A2(_02585_),
    .Y(_00216_),
    .B1(_02577_));
 sg13g2_nor2_1 _08648_ (.A(_02563_),
    .B(_02578_),
    .Y(_02586_));
 sg13g2_nand4_1 _08649_ (.B(_02540_),
    .C(_02554_),
    .A(_02538_),
    .Y(_02587_),
    .D(_02586_));
 sg13g2_o21ai_1 _08650_ (.B1(net3227),
    .Y(_02588_),
    .A1(\u_toplayer.u_outlayer.u_neuron.acc[19] ),
    .A2(net3196));
 sg13g2_nand3_1 _08651_ (.B(_02587_),
    .C(_02588_),
    .A(_02564_),
    .Y(_02589_));
 sg13g2_xor2_1 _08652_ (.B(net3226),
    .A(net3195),
    .X(_02590_));
 sg13g2_xnor2_1 _08653_ (.Y(_02591_),
    .A(\u_toplayer.u_outlayer.u_neuron.acc[20] ),
    .B(net3226));
 sg13g2_and2_1 _08654_ (.A(_02589_),
    .B(_02590_),
    .X(_02592_));
 sg13g2_nor2_1 _08655_ (.A(net2979),
    .B(_02592_),
    .Y(_02593_));
 sg13g2_o21ai_1 _08656_ (.B1(_02593_),
    .Y(_02594_),
    .A1(_02589_),
    .A2(_02590_));
 sg13g2_xnor2_1 _08657_ (.Y(_02595_),
    .A(net3195),
    .B(net3360));
 sg13g2_or4_1 _08658_ (.A(_02547_),
    .B(_02569_),
    .C(_02570_),
    .D(_02581_),
    .X(_02596_));
 sg13g2_o21ai_1 _08659_ (.B1(net3360),
    .Y(_02597_),
    .A1(\u_toplayer.u_outlayer.u_neuron.acc[19] ),
    .A2(net3196));
 sg13g2_nand2_1 _08660_ (.Y(_02598_),
    .A(_02572_),
    .B(_02597_));
 sg13g2_inv_1 _08661_ (.Y(_02599_),
    .A(_02598_));
 sg13g2_a21o_1 _08662_ (.A2(_02599_),
    .A1(_02596_),
    .B1(_02595_),
    .X(_02600_));
 sg13g2_nand3_1 _08663_ (.B(_02596_),
    .C(_02599_),
    .A(_02595_),
    .Y(_02601_));
 sg13g2_and2_1 _08664_ (.A(net2933),
    .B(_02601_),
    .X(_02602_));
 sg13g2_a21oi_1 _08665_ (.A1(_02600_),
    .A2(_02602_),
    .Y(_02603_),
    .B1(net2893));
 sg13g2_a22oi_1 _08666_ (.Y(_00217_),
    .B1(_02594_),
    .B2(_02603_),
    .A2(net2893),
    .A1(_01045_));
 sg13g2_xnor2_1 _08667_ (.Y(_02604_),
    .A(\u_toplayer.u_outlayer.u_neuron.acc[21] ),
    .B(net3226));
 sg13g2_a21oi_1 _08668_ (.A1(net3195),
    .A2(net3226),
    .Y(_02605_),
    .B1(_02592_));
 sg13g2_xor2_1 _08669_ (.B(_02605_),
    .A(_02604_),
    .X(_02606_));
 sg13g2_xor2_1 _08670_ (.B(net3359),
    .A(\u_toplayer.u_outlayer.u_neuron.acc[21] ),
    .X(_02607_));
 sg13g2_inv_1 _08671_ (.Y(_02608_),
    .A(_02607_));
 sg13g2_o21ai_1 _08672_ (.B1(_02600_),
    .Y(_02609_),
    .A1(_01045_),
    .A2(_01047_));
 sg13g2_xnor2_1 _08673_ (.Y(_02610_),
    .A(_02608_),
    .B(_02609_));
 sg13g2_a221oi_1 _08674_ (.B2(net2933),
    .C1(net2892),
    .B1(_02610_),
    .A1(net2976),
    .Y(_02611_),
    .A2(_02606_));
 sg13g2_a21oi_1 _08675_ (.A1(_01044_),
    .A2(net2892),
    .Y(_00218_),
    .B1(_02611_));
 sg13g2_nand2_1 _08676_ (.Y(_02612_),
    .A(\u_toplayer.u_outlayer.u_neuron.acc[22] ),
    .B(net3361));
 sg13g2_xor2_1 _08677_ (.B(net3361),
    .A(\u_toplayer.u_outlayer.u_neuron.acc[22] ),
    .X(_02613_));
 sg13g2_o21ai_1 _08678_ (.B1(net3359),
    .Y(_02614_),
    .A1(\u_toplayer.u_outlayer.u_neuron.acc[21] ),
    .A2(net3195));
 sg13g2_o21ai_1 _08679_ (.B1(_02614_),
    .Y(_02615_),
    .A1(_02600_),
    .A2(_02608_));
 sg13g2_nor2_1 _08680_ (.A(_02613_),
    .B(_02615_),
    .Y(_02616_));
 sg13g2_nand2_1 _08681_ (.Y(_02617_),
    .A(_02613_),
    .B(_02615_));
 sg13g2_nor2_1 _08682_ (.A(net2932),
    .B(_02616_),
    .Y(_02618_));
 sg13g2_and2_1 _08683_ (.A(\u_toplayer.u_outlayer.u_neuron.acc[22] ),
    .B(net3228),
    .X(_02619_));
 sg13g2_xor2_1 _08684_ (.B(net3228),
    .A(\u_toplayer.u_outlayer.u_neuron.acc[22] ),
    .X(_02620_));
 sg13g2_nor2_1 _08685_ (.A(_02591_),
    .B(_02604_),
    .Y(_02621_));
 sg13g2_o21ai_1 _08686_ (.B1(net3228),
    .Y(_02622_),
    .A1(\u_toplayer.u_outlayer.u_neuron.acc[21] ),
    .A2(net3195));
 sg13g2_inv_1 _08687_ (.Y(_02623_),
    .A(_02622_));
 sg13g2_a21o_1 _08688_ (.A2(_02621_),
    .A1(_02589_),
    .B1(_02623_),
    .X(_02624_));
 sg13g2_a21oi_1 _08689_ (.A1(_02620_),
    .A2(_02624_),
    .Y(_02625_),
    .B1(net2979));
 sg13g2_o21ai_1 _08690_ (.B1(_02625_),
    .Y(_02626_),
    .A1(_02620_),
    .A2(_02624_));
 sg13g2_a21oi_1 _08691_ (.A1(_02617_),
    .A2(_02618_),
    .Y(_02627_),
    .B1(net2892));
 sg13g2_a22oi_1 _08692_ (.Y(_00219_),
    .B1(_02626_),
    .B2(_02627_),
    .A2(net2892),
    .A1(_01043_));
 sg13g2_nor2_1 _08693_ (.A(net1042),
    .B(net2889),
    .Y(_02628_));
 sg13g2_xnor2_1 _08694_ (.Y(_02629_),
    .A(\u_toplayer.u_outlayer.u_neuron.acc[23] ),
    .B(net3361));
 sg13g2_a21oi_1 _08695_ (.A1(_02612_),
    .A2(_02617_),
    .Y(_02630_),
    .B1(_02629_));
 sg13g2_nand3_1 _08696_ (.B(_02617_),
    .C(_02629_),
    .A(_02612_),
    .Y(_02631_));
 sg13g2_nor2_1 _08697_ (.A(net2932),
    .B(_02630_),
    .Y(_02632_));
 sg13g2_a21oi_1 _08698_ (.A1(_02620_),
    .A2(_02624_),
    .Y(_02633_),
    .B1(_02619_));
 sg13g2_xor2_1 _08699_ (.B(net3228),
    .A(\u_toplayer.u_outlayer.u_neuron.acc[23] ),
    .X(_02634_));
 sg13g2_xnor2_1 _08700_ (.Y(_02635_),
    .A(_02633_),
    .B(_02634_));
 sg13g2_a22oi_1 _08701_ (.Y(_02636_),
    .B1(_02635_),
    .B2(net2976),
    .A2(_02632_),
    .A1(_02631_));
 sg13g2_a21oi_1 _08702_ (.A1(net2890),
    .A2(_02636_),
    .Y(_00220_),
    .B1(_02628_));
 sg13g2_nand2_2 _08703_ (.Y(_02637_),
    .A(\u_toplayer.u_layer2.u_neuron.instCtrl.state[5] ),
    .B(_01350_));
 sg13g2_nor3_1 _08704_ (.A(_00032_),
    .B(_01353_),
    .C(_02637_),
    .Y(_02638_));
 sg13g2_or3_1 _08705_ (.A(_00032_),
    .B(_01353_),
    .C(_02637_),
    .X(_02639_));
 sg13g2_nor2_1 _08706_ (.A(net3255),
    .B(_02637_),
    .Y(_02640_));
 sg13g2_o21ai_1 _08707_ (.B1(_00032_),
    .Y(_02641_),
    .A1(net3277),
    .A2(_02637_));
 sg13g2_nor2b_2 _08708_ (.A(net3258),
    .B_N(net3245),
    .Y(_02642_));
 sg13g2_nor2b_1 _08709_ (.A(_02640_),
    .B_N(_02641_),
    .Y(_02643_));
 sg13g2_nand2b_1 _08710_ (.Y(_02644_),
    .B(_02641_),
    .A_N(_02640_));
 sg13g2_o21ai_1 _08711_ (.B1(net2860),
    .Y(_02645_),
    .A1(_01353_),
    .A2(_02637_));
 sg13g2_and2_1 _08712_ (.A(\u_toplayer.delayed_done_layer1 ),
    .B(_02645_),
    .X(_02646_));
 sg13g2_nand2_2 _08713_ (.Y(_02647_),
    .A(\u_toplayer.delayed_done_layer1 ),
    .B(_02645_));
 sg13g2_and4_1 _08714_ (.A(net3242),
    .B(\u_toplayer.u_layer2.u_neuron.instCtrl.state[5] ),
    .C(_01346_),
    .D(_01347_),
    .X(_02648_));
 sg13g2_nor2_1 _08715_ (.A(_02646_),
    .B(_02648_),
    .Y(_02649_));
 sg13g2_o21ai_1 _08716_ (.B1(net2884),
    .Y(_02650_),
    .A1(_02646_),
    .A2(_02648_));
 sg13g2_nand2_1 _08717_ (.Y(_02651_),
    .A(net929),
    .B(_02650_));
 sg13g2_nor2_2 _08718_ (.A(net2861),
    .B(net2748),
    .Y(_02652_));
 sg13g2_nand2b_2 _08719_ (.Y(_02653_),
    .B(net2858),
    .A_N(_02650_));
 sg13g2_nand2_2 _08720_ (.Y(_02654_),
    .A(net3349),
    .B(net3095));
 sg13g2_o21ai_1 _08721_ (.B1(_02651_),
    .Y(_00227_),
    .A1(_02653_),
    .A2(_02654_));
 sg13g2_nand2_2 _08722_ (.Y(_02655_),
    .A(net3338),
    .B(net3093));
 sg13g2_nor2_1 _08723_ (.A(_02654_),
    .B(_02655_),
    .Y(_02656_));
 sg13g2_a22oi_1 _08724_ (.Y(_02657_),
    .B1(net3093),
    .B2(net3349),
    .A2(net3095),
    .A1(net3342));
 sg13g2_nor3_1 _08725_ (.A(_02653_),
    .B(_02656_),
    .C(_02657_),
    .Y(_02658_));
 sg13g2_a21o_1 _08726_ (.A2(net2748),
    .A1(net1003),
    .B1(_02658_),
    .X(_00228_));
 sg13g2_nand2_1 _08727_ (.Y(_02659_),
    .A(net830),
    .B(net2748));
 sg13g2_nand2_1 _08728_ (.Y(_02660_),
    .A(net3328),
    .B(net3091));
 sg13g2_nor2_1 _08729_ (.A(_02654_),
    .B(_02660_),
    .Y(_02661_));
 sg13g2_a22oi_1 _08730_ (.Y(_02662_),
    .B1(net3091),
    .B2(net3349),
    .A2(net3095),
    .A1(net3328));
 sg13g2_or2_1 _08731_ (.X(_02663_),
    .B(_02662_),
    .A(_02661_));
 sg13g2_inv_1 _08732_ (.Y(_02664_),
    .A(_02663_));
 sg13g2_nand2b_1 _08733_ (.Y(_02665_),
    .B(_02654_),
    .A_N(_02655_));
 sg13g2_xnor2_1 _08734_ (.Y(_02666_),
    .A(_02663_),
    .B(_02665_));
 sg13g2_o21ai_1 _08735_ (.B1(_02659_),
    .Y(_00229_),
    .A1(_02653_),
    .A2(_02666_));
 sg13g2_nand2_1 _08736_ (.Y(_02667_),
    .A(net888),
    .B(net2748));
 sg13g2_a21oi_1 _08737_ (.A1(_02654_),
    .A2(_02662_),
    .Y(_02668_),
    .B1(_02655_));
 sg13g2_nand4_1 _08738_ (.B(net3315),
    .C(net3094),
    .A(net3339),
    .Y(_02669_),
    .D(net3090));
 sg13g2_inv_1 _08739_ (.Y(_02670_),
    .A(_02669_));
 sg13g2_a22oi_1 _08740_ (.Y(_02671_),
    .B1(net3091),
    .B2(net3338),
    .A2(net3094),
    .A1(net3315));
 sg13g2_nor2_2 _08741_ (.A(_02670_),
    .B(_02671_),
    .Y(_02672_));
 sg13g2_and4_1 _08742_ (.A(net3350),
    .B(net3328),
    .C(net3092),
    .D(net3089),
    .X(_02673_));
 sg13g2_a22oi_1 _08743_ (.Y(_02674_),
    .B1(net3089),
    .B2(net3348),
    .A2(net3093),
    .A1(net3328));
 sg13g2_nor2_1 _08744_ (.A(_02673_),
    .B(_02674_),
    .Y(_02675_));
 sg13g2_and2_1 _08745_ (.A(_02661_),
    .B(_02675_),
    .X(_02676_));
 sg13g2_xor2_1 _08746_ (.B(_02675_),
    .A(_02661_),
    .X(_02677_));
 sg13g2_xor2_1 _08747_ (.B(_02677_),
    .A(_02672_),
    .X(_02678_));
 sg13g2_xnor2_1 _08748_ (.Y(_02679_),
    .A(_02672_),
    .B(_02677_));
 sg13g2_xnor2_1 _08749_ (.Y(_02680_),
    .A(_02668_),
    .B(_02678_));
 sg13g2_o21ai_1 _08750_ (.B1(_02667_),
    .Y(_00230_),
    .A1(net2727),
    .A2(_02680_));
 sg13g2_nand2_1 _08751_ (.Y(_02681_),
    .A(net897),
    .B(net2748));
 sg13g2_nand2_1 _08752_ (.Y(_02682_),
    .A(_02656_),
    .B(_02678_));
 sg13g2_nor2_1 _08753_ (.A(_02664_),
    .B(_02682_),
    .Y(_02683_));
 sg13g2_nor3_1 _08754_ (.A(_02655_),
    .B(_02663_),
    .C(_02679_),
    .Y(_02684_));
 sg13g2_nand2_1 _08755_ (.Y(_02685_),
    .A(net3339),
    .B(net3089));
 sg13g2_nand2_1 _08756_ (.Y(_02686_),
    .A(net3315),
    .B(net3093));
 sg13g2_or2_1 _08757_ (.X(_02687_),
    .B(_02686_),
    .A(_02685_));
 sg13g2_xor2_1 _08758_ (.B(_02686_),
    .A(_02685_),
    .X(_02688_));
 sg13g2_nand2_1 _08759_ (.Y(_02689_),
    .A(_02670_),
    .B(_02688_));
 sg13g2_xnor2_1 _08760_ (.Y(_02690_),
    .A(_02669_),
    .B(_02688_));
 sg13g2_nand2_1 _08761_ (.Y(_02691_),
    .A(net3301),
    .B(net3086));
 sg13g2_and4_2 _08762_ (.A(net3348),
    .B(net3304),
    .C(net3095),
    .D(net3087),
    .X(_02692_));
 sg13g2_a22oi_1 _08763_ (.Y(_02693_),
    .B1(net3087),
    .B2(net3348),
    .A2(net3095),
    .A1(net3304));
 sg13g2_or3_1 _08764_ (.A(_02660_),
    .B(_02692_),
    .C(_02693_),
    .X(_02694_));
 sg13g2_o21ai_1 _08765_ (.B1(_02660_),
    .Y(_02695_),
    .A1(_02692_),
    .A2(_02693_));
 sg13g2_nand3_1 _08766_ (.B(_02694_),
    .C(_02695_),
    .A(_02673_),
    .Y(_02696_));
 sg13g2_inv_1 _08767_ (.Y(_02697_),
    .A(_02696_));
 sg13g2_a21o_1 _08768_ (.A2(_02695_),
    .A1(_02694_),
    .B1(_02673_),
    .X(_02698_));
 sg13g2_and2_1 _08769_ (.A(_02696_),
    .B(_02698_),
    .X(_02699_));
 sg13g2_xnor2_1 _08770_ (.Y(_02700_),
    .A(_02690_),
    .B(_02699_));
 sg13g2_a21oi_1 _08771_ (.A1(_02672_),
    .A2(_02677_),
    .Y(_02701_),
    .B1(_02676_));
 sg13g2_nor2_1 _08772_ (.A(_02700_),
    .B(_02701_),
    .Y(_02702_));
 sg13g2_xnor2_1 _08773_ (.Y(_02703_),
    .A(_02700_),
    .B(_02701_));
 sg13g2_nor4_1 _08774_ (.A(_02655_),
    .B(_02663_),
    .C(_02679_),
    .D(_02703_),
    .Y(_02704_));
 sg13g2_xnor2_1 _08775_ (.Y(_02705_),
    .A(_02684_),
    .B(_02703_));
 sg13g2_nor3_1 _08776_ (.A(_02664_),
    .B(_02682_),
    .C(_02703_),
    .Y(_02706_));
 sg13g2_o21ai_1 _08777_ (.B1(_02652_),
    .Y(_02707_),
    .A1(_02683_),
    .A2(_02705_));
 sg13g2_o21ai_1 _08778_ (.B1(_02681_),
    .Y(_00231_),
    .A1(_02706_),
    .A2(_02707_));
 sg13g2_nand2_1 _08779_ (.Y(_02708_),
    .A(net948),
    .B(net2748));
 sg13g2_nor2_1 _08780_ (.A(_02704_),
    .B(_02706_),
    .Y(_02709_));
 sg13g2_a21o_1 _08781_ (.A2(_02698_),
    .A1(_02690_),
    .B1(_02697_),
    .X(_02710_));
 sg13g2_a22oi_1 _08782_ (.Y(_02711_),
    .B1(net3087),
    .B2(net3339),
    .A2(net3091),
    .A1(net3315));
 sg13g2_nand2_1 _08783_ (.Y(_02712_),
    .A(net3313),
    .B(net3087));
 sg13g2_nand4_1 _08784_ (.B(net3315),
    .C(net3090),
    .A(net3339),
    .Y(_02713_),
    .D(net3086));
 sg13g2_nor2b_1 _08785_ (.A(_02711_),
    .B_N(_02713_),
    .Y(_02714_));
 sg13g2_xor2_1 _08786_ (.B(_02714_),
    .A(_02692_),
    .X(_02715_));
 sg13g2_nor2b_1 _08787_ (.A(_02687_),
    .B_N(_02715_),
    .Y(_02716_));
 sg13g2_xnor2_1 _08788_ (.Y(_02717_),
    .A(_02687_),
    .B(_02715_));
 sg13g2_nand2_1 _08789_ (.Y(_02718_),
    .A(net3347),
    .B(net3085));
 sg13g2_nand2_1 _08790_ (.Y(_02719_),
    .A(net3295),
    .B(net3092));
 sg13g2_and4_1 _08791_ (.A(net3304),
    .B(net3296),
    .C(net3094),
    .D(net3092),
    .X(_02720_));
 sg13g2_a22oi_1 _08792_ (.Y(_02721_),
    .B1(net3092),
    .B2(net3304),
    .A2(net3095),
    .A1(net3296));
 sg13g2_o21ai_1 _08793_ (.B1(_02718_),
    .Y(_02722_),
    .A1(_02720_),
    .A2(_02721_));
 sg13g2_or3_1 _08794_ (.A(_02718_),
    .B(_02720_),
    .C(_02721_),
    .X(_02723_));
 sg13g2_and4_1 _08795_ (.A(net3328),
    .B(net3088),
    .C(_02722_),
    .D(_02723_),
    .X(_02724_));
 sg13g2_nand4_1 _08796_ (.B(net3088),
    .C(_02722_),
    .A(net3328),
    .Y(_02725_),
    .D(_02723_));
 sg13g2_a22oi_1 _08797_ (.Y(_02726_),
    .B1(_02722_),
    .B2(_02723_),
    .A2(net3088),
    .A1(net3328));
 sg13g2_or3_1 _08798_ (.A(_02694_),
    .B(_02724_),
    .C(_02726_),
    .X(_02727_));
 sg13g2_o21ai_1 _08799_ (.B1(_02694_),
    .Y(_02728_),
    .A1(_02724_),
    .A2(_02726_));
 sg13g2_nand3_1 _08800_ (.B(_02727_),
    .C(_02728_),
    .A(_02717_),
    .Y(_02729_));
 sg13g2_a21o_1 _08801_ (.A2(_02728_),
    .A1(_02727_),
    .B1(_02717_),
    .X(_02730_));
 sg13g2_and3_1 _08802_ (.X(_02731_),
    .A(_02710_),
    .B(_02729_),
    .C(_02730_));
 sg13g2_a21oi_1 _08803_ (.A1(_02729_),
    .A2(_02730_),
    .Y(_02732_),
    .B1(_02710_));
 sg13g2_o21ai_1 _08804_ (.B1(_02689_),
    .Y(_02733_),
    .A1(_02731_),
    .A2(_02732_));
 sg13g2_or3_1 _08805_ (.A(_02689_),
    .B(_02731_),
    .C(_02732_),
    .X(_02734_));
 sg13g2_nand2_1 _08806_ (.Y(_02735_),
    .A(_02733_),
    .B(_02734_));
 sg13g2_nand3_1 _08807_ (.B(_02733_),
    .C(_02734_),
    .A(_02702_),
    .Y(_02736_));
 sg13g2_a21oi_1 _08808_ (.A1(_02733_),
    .A2(_02734_),
    .Y(_02737_),
    .B1(_02702_));
 sg13g2_xor2_1 _08809_ (.B(_02735_),
    .A(_02702_),
    .X(_02738_));
 sg13g2_xnor2_1 _08810_ (.Y(_02739_),
    .A(_02709_),
    .B(_02738_));
 sg13g2_o21ai_1 _08811_ (.B1(_02708_),
    .Y(_00232_),
    .A1(net2727),
    .A2(_02739_));
 sg13g2_a21oi_2 _08812_ (.B1(_02716_),
    .Y(_02740_),
    .A2(_02714_),
    .A1(_02692_));
 sg13g2_inv_1 _08813_ (.Y(_02741_),
    .A(_02740_));
 sg13g2_and2_1 _08814_ (.A(_02727_),
    .B(_02729_),
    .X(_02742_));
 sg13g2_nor2b_1 _08815_ (.A(_02720_),
    .B_N(_02723_),
    .Y(_02743_));
 sg13g2_a22oi_1 _08816_ (.Y(_02744_),
    .B1(net3085),
    .B2(net3334),
    .A2(net3089),
    .A1(net3307));
 sg13g2_nand4_1 _08817_ (.B(net3307),
    .C(net3089),
    .A(net3334),
    .Y(_02745_),
    .D(\u_toplayer.u_layer2.u_neuron.din[5] ));
 sg13g2_nor2b_1 _08818_ (.A(_02744_),
    .B_N(_02745_),
    .Y(_02746_));
 sg13g2_nand2b_1 _08819_ (.Y(_02747_),
    .B(_02746_),
    .A_N(_02743_));
 sg13g2_xor2_1 _08820_ (.B(_02746_),
    .A(_02743_),
    .X(_02748_));
 sg13g2_xor2_1 _08821_ (.B(_02748_),
    .A(_02713_),
    .X(_02749_));
 sg13g2_nand2_1 _08822_ (.Y(_02750_),
    .A(net3347),
    .B(\u_toplayer.u_layer2.u_neuron.din[6] ));
 sg13g2_nand2_1 _08823_ (.Y(_02751_),
    .A(net3301),
    .B(net3090));
 sg13g2_or2_1 _08824_ (.X(_02752_),
    .B(_02751_),
    .A(_02719_));
 sg13g2_and2_1 _08825_ (.A(_02719_),
    .B(_02751_),
    .X(_02753_));
 sg13g2_xor2_1 _08826_ (.B(_02751_),
    .A(_02719_),
    .X(_02754_));
 sg13g2_xnor2_1 _08827_ (.Y(_02755_),
    .A(_02750_),
    .B(_02754_));
 sg13g2_nand2_1 _08828_ (.Y(_02756_),
    .A(net3287),
    .B(net3086));
 sg13g2_nand4_1 _08829_ (.B(net3287),
    .C(net3094),
    .A(net3327),
    .Y(_02757_),
    .D(net3086));
 sg13g2_inv_1 _08830_ (.Y(_02758_),
    .A(_02757_));
 sg13g2_a22oi_1 _08831_ (.Y(_02759_),
    .B1(net3086),
    .B2(net3327),
    .A2(net3094),
    .A1(net3290));
 sg13g2_nor2_1 _08832_ (.A(_02758_),
    .B(_02759_),
    .Y(_02760_));
 sg13g2_nand2_1 _08833_ (.Y(_02761_),
    .A(_02755_),
    .B(_02760_));
 sg13g2_xnor2_1 _08834_ (.Y(_02762_),
    .A(_02755_),
    .B(_02760_));
 sg13g2_nor2_1 _08835_ (.A(_02725_),
    .B(_02762_),
    .Y(_02763_));
 sg13g2_xnor2_1 _08836_ (.Y(_02764_),
    .A(_02724_),
    .B(_02762_));
 sg13g2_xnor2_1 _08837_ (.Y(_02765_),
    .A(_02749_),
    .B(_02764_));
 sg13g2_nor2_1 _08838_ (.A(_02742_),
    .B(_02765_),
    .Y(_02766_));
 sg13g2_xor2_1 _08839_ (.B(_02765_),
    .A(_02742_),
    .X(_02767_));
 sg13g2_xnor2_1 _08840_ (.Y(_02768_),
    .A(_02740_),
    .B(_02767_));
 sg13g2_nand2b_1 _08841_ (.Y(_02769_),
    .B(_02734_),
    .A_N(_02731_));
 sg13g2_and2_1 _08842_ (.A(_02768_),
    .B(_02769_),
    .X(_02770_));
 sg13g2_xor2_1 _08843_ (.B(_02769_),
    .A(_02768_),
    .X(_02771_));
 sg13g2_o21ai_1 _08844_ (.B1(_02736_),
    .Y(_02772_),
    .A1(_02709_),
    .A2(_02737_));
 sg13g2_nor2_1 _08845_ (.A(_02771_),
    .B(_02772_),
    .Y(_02773_));
 sg13g2_nand2_1 _08846_ (.Y(_02774_),
    .A(_02771_),
    .B(_02772_));
 sg13g2_nor2_1 _08847_ (.A(net2727),
    .B(_02773_),
    .Y(_02775_));
 sg13g2_a22oi_1 _08848_ (.Y(_02776_),
    .B1(_02774_),
    .B2(_02775_),
    .A2(net2748),
    .A1(net975));
 sg13g2_inv_1 _08849_ (.Y(_00233_),
    .A(_02776_));
 sg13g2_o21ai_1 _08850_ (.B1(_02747_),
    .Y(_02777_),
    .A1(_02713_),
    .A2(_02748_));
 sg13g2_a21oi_1 _08851_ (.A1(_02749_),
    .A2(_02764_),
    .Y(_02778_),
    .B1(_02763_));
 sg13g2_o21ai_1 _08852_ (.B1(_02752_),
    .Y(_02779_),
    .A1(_02750_),
    .A2(_02753_));
 sg13g2_nand2_1 _08853_ (.Y(_02780_),
    .A(net3347),
    .B(net3082));
 sg13g2_nand2_1 _08854_ (.Y(_02781_),
    .A(net3337),
    .B(\u_toplayer.u_layer2.u_neuron.din[6] ));
 sg13g2_xor2_1 _08855_ (.B(_02781_),
    .A(net2953),
    .X(_02782_));
 sg13g2_nand2b_1 _08856_ (.Y(_02783_),
    .B(_02782_),
    .A_N(_02712_));
 sg13g2_xnor2_1 _08857_ (.Y(_02784_),
    .A(_02712_),
    .B(_02782_));
 sg13g2_nand2_1 _08858_ (.Y(_02785_),
    .A(_02779_),
    .B(_02784_));
 sg13g2_xnor2_1 _08859_ (.Y(_02786_),
    .A(_02779_),
    .B(_02784_));
 sg13g2_xor2_1 _08860_ (.B(_02786_),
    .A(_02745_),
    .X(_02787_));
 sg13g2_nand2_1 _08861_ (.Y(_02788_),
    .A(net3301),
    .B(net3088));
 sg13g2_and2_1 _08862_ (.A(net3288),
    .B(net3090),
    .X(_02789_));
 sg13g2_and4_1 _08863_ (.A(net3293),
    .B(net3287),
    .C(net3092),
    .D(net3090),
    .X(_02790_));
 sg13g2_a22oi_1 _08864_ (.Y(_02791_),
    .B1(net3090),
    .B2(net3293),
    .A2(net3092),
    .A1(net3287));
 sg13g2_nor3_1 _08865_ (.A(_02788_),
    .B(_02790_),
    .C(_02791_),
    .Y(_02792_));
 sg13g2_o21ai_1 _08866_ (.B1(_02788_),
    .Y(_02793_),
    .A1(_02790_),
    .A2(_02791_));
 sg13g2_nor2b_1 _08867_ (.A(_02792_),
    .B_N(_02793_),
    .Y(_02794_));
 sg13g2_nand2_1 _08868_ (.Y(_02795_),
    .A(net3327),
    .B(net3085));
 sg13g2_nand2_1 _08869_ (.Y(_02796_),
    .A(net3284),
    .B(net3094));
 sg13g2_xor2_1 _08870_ (.B(_02796_),
    .A(_02795_),
    .X(_02797_));
 sg13g2_xnor2_1 _08871_ (.Y(_02798_),
    .A(_02757_),
    .B(_02797_));
 sg13g2_and2_1 _08872_ (.A(_02794_),
    .B(_02798_),
    .X(_02799_));
 sg13g2_xnor2_1 _08873_ (.Y(_02800_),
    .A(_02794_),
    .B(_02798_));
 sg13g2_nor2_1 _08874_ (.A(_02761_),
    .B(_02800_),
    .Y(_02801_));
 sg13g2_xor2_1 _08875_ (.B(_02800_),
    .A(_02761_),
    .X(_02802_));
 sg13g2_xnor2_1 _08876_ (.Y(_02803_),
    .A(_02787_),
    .B(_02802_));
 sg13g2_nor2_1 _08877_ (.A(_02778_),
    .B(_02803_),
    .Y(_02804_));
 sg13g2_xor2_1 _08878_ (.B(_02803_),
    .A(_02778_),
    .X(_02805_));
 sg13g2_xnor2_1 _08879_ (.Y(_02806_),
    .A(_02777_),
    .B(_02805_));
 sg13g2_a21oi_1 _08880_ (.A1(_02741_),
    .A2(_02767_),
    .Y(_02807_),
    .B1(_02766_));
 sg13g2_nor2_1 _08881_ (.A(_02806_),
    .B(_02807_),
    .Y(_02808_));
 sg13g2_xor2_1 _08882_ (.B(_02807_),
    .A(_02806_),
    .X(_02809_));
 sg13g2_nand3_1 _08883_ (.B(_02772_),
    .C(_02809_),
    .A(_02771_),
    .Y(_02810_));
 sg13g2_nor2_1 _08884_ (.A(_02770_),
    .B(_02809_),
    .Y(_02811_));
 sg13g2_nand2_1 _08885_ (.Y(_02812_),
    .A(_02774_),
    .B(_02811_));
 sg13g2_a21oi_1 _08886_ (.A1(_02770_),
    .A2(_02809_),
    .Y(_02813_),
    .B1(net2727));
 sg13g2_and2_1 _08887_ (.A(_02810_),
    .B(_02813_),
    .X(_02814_));
 sg13g2_a22oi_1 _08888_ (.Y(_02815_),
    .B1(_02812_),
    .B2(_02814_),
    .A2(net2748),
    .A1(net944));
 sg13g2_inv_1 _08889_ (.Y(_00234_),
    .A(_02815_));
 sg13g2_nand2_1 _08890_ (.Y(_02816_),
    .A(net916),
    .B(net2749));
 sg13g2_o21ai_1 _08891_ (.B1(_02785_),
    .Y(_02817_),
    .A1(_02745_),
    .A2(_02786_));
 sg13g2_a21oi_1 _08892_ (.A1(_02787_),
    .A2(_02802_),
    .Y(_02818_),
    .B1(_02801_));
 sg13g2_o21ai_1 _08893_ (.B1(_02783_),
    .Y(_02819_),
    .A1(net2953),
    .A2(_02781_));
 sg13g2_or2_1 _08894_ (.X(_02820_),
    .B(_02792_),
    .A(_02790_));
 sg13g2_a22oi_1 _08895_ (.Y(_02821_),
    .B1(net3083),
    .B2(net3334),
    .A2(\u_toplayer.u_layer2.u_neuron.din[5] ),
    .A1(net3307));
 sg13g2_nand4_1 _08896_ (.B(net3307),
    .C(\u_toplayer.u_layer2.u_neuron.din[5] ),
    .A(net3334),
    .Y(_02822_),
    .D(net3083));
 sg13g2_nor2b_1 _08897_ (.A(_02821_),
    .B_N(_02822_),
    .Y(_02823_));
 sg13g2_xnor2_1 _08898_ (.Y(_02824_),
    .A(_02820_),
    .B(_02823_));
 sg13g2_nor2b_1 _08899_ (.A(_02824_),
    .B_N(_02819_),
    .Y(_02825_));
 sg13g2_xor2_1 _08900_ (.B(_02824_),
    .A(_02819_),
    .X(_02826_));
 sg13g2_a21o_1 _08901_ (.A2(_02797_),
    .A1(_02758_),
    .B1(_02799_),
    .X(_02827_));
 sg13g2_nand2_1 _08902_ (.Y(_02828_),
    .A(net3293),
    .B(net3088));
 sg13g2_xor2_1 _08903_ (.B(_02828_),
    .A(_02691_),
    .X(_02829_));
 sg13g2_nand2b_1 _08904_ (.Y(_02830_),
    .B(_02829_),
    .A_N(net2953));
 sg13g2_xnor2_1 _08905_ (.Y(_02831_),
    .A(net2952),
    .B(_02829_));
 sg13g2_inv_1 _08906_ (.Y(_02832_),
    .A(_02831_));
 sg13g2_a21oi_1 _08907_ (.A1(net3094),
    .A2(_02795_),
    .Y(_02833_),
    .B1(net3280));
 sg13g2_nand2_1 _08908_ (.Y(_02834_),
    .A(net3327),
    .B(net3084));
 sg13g2_nor2b_1 _08909_ (.A(net3092),
    .B_N(net3284),
    .Y(_02835_));
 sg13g2_nor2b_1 _08910_ (.A(_02834_),
    .B_N(_02835_),
    .Y(_02836_));
 sg13g2_xnor2_1 _08911_ (.Y(_02837_),
    .A(_02834_),
    .B(_02835_));
 sg13g2_xor2_1 _08912_ (.B(_02837_),
    .A(_02789_),
    .X(_02838_));
 sg13g2_nand2_1 _08913_ (.Y(_02839_),
    .A(_02833_),
    .B(_02838_));
 sg13g2_xnor2_1 _08914_ (.Y(_02840_),
    .A(_02833_),
    .B(_02838_));
 sg13g2_xnor2_1 _08915_ (.Y(_02841_),
    .A(_02832_),
    .B(_02840_));
 sg13g2_nand2b_1 _08916_ (.Y(_02842_),
    .B(_02827_),
    .A_N(_02841_));
 sg13g2_xor2_1 _08917_ (.B(_02841_),
    .A(_02827_),
    .X(_02843_));
 sg13g2_xor2_1 _08918_ (.B(_02843_),
    .A(_02826_),
    .X(_02844_));
 sg13g2_nor2b_1 _08919_ (.A(_02818_),
    .B_N(_02844_),
    .Y(_02845_));
 sg13g2_xnor2_1 _08920_ (.Y(_02846_),
    .A(_02818_),
    .B(_02844_));
 sg13g2_xor2_1 _08921_ (.B(_02846_),
    .A(_02817_),
    .X(_02847_));
 sg13g2_xnor2_1 _08922_ (.Y(_02848_),
    .A(_02817_),
    .B(_02846_));
 sg13g2_a21oi_1 _08923_ (.A1(_02777_),
    .A2(_02805_),
    .Y(_02849_),
    .B1(_02804_));
 sg13g2_a21o_1 _08924_ (.A2(_02805_),
    .A1(_02777_),
    .B1(_02804_),
    .X(_02850_));
 sg13g2_nor2_1 _08925_ (.A(_02848_),
    .B(_02849_),
    .Y(_02851_));
 sg13g2_xnor2_1 _08926_ (.Y(_02852_),
    .A(_02848_),
    .B(_02849_));
 sg13g2_a21oi_1 _08927_ (.A1(_02770_),
    .A2(_02809_),
    .Y(_02853_),
    .B1(_02808_));
 sg13g2_and2_1 _08928_ (.A(_02810_),
    .B(_02853_),
    .X(_02854_));
 sg13g2_a21oi_2 _08929_ (.B1(_02852_),
    .Y(_02855_),
    .A2(_02853_),
    .A1(_02810_));
 sg13g2_a21o_1 _08930_ (.A2(_02854_),
    .A1(_02852_),
    .B1(net2727),
    .X(_02856_));
 sg13g2_o21ai_1 _08931_ (.B1(_02816_),
    .Y(_00235_),
    .A1(_02855_),
    .A2(_02856_));
 sg13g2_a21o_1 _08932_ (.A2(_02846_),
    .A1(_02817_),
    .B1(_02845_),
    .X(_02857_));
 sg13g2_a21o_1 _08933_ (.A2(_02823_),
    .A1(_02820_),
    .B1(_02825_),
    .X(_02858_));
 sg13g2_inv_1 _08934_ (.Y(_02859_),
    .A(_02858_));
 sg13g2_o21ai_1 _08935_ (.B1(_02842_),
    .Y(_02860_),
    .A1(_02826_),
    .A2(_02843_));
 sg13g2_o21ai_1 _08936_ (.B1(_02830_),
    .Y(_02861_),
    .A1(_02691_),
    .A2(_02828_));
 sg13g2_a22oi_1 _08937_ (.Y(_02862_),
    .B1(net3083),
    .B2(net3334),
    .A2(net3084),
    .A1(net3307));
 sg13g2_nand4_1 _08938_ (.B(net3307),
    .C(net3084),
    .A(net3334),
    .Y(_02863_),
    .D(net3083));
 sg13g2_nor2b_1 _08939_ (.A(_02862_),
    .B_N(_02863_),
    .Y(_02864_));
 sg13g2_nand2_1 _08940_ (.Y(_02865_),
    .A(_02861_),
    .B(_02864_));
 sg13g2_xnor2_1 _08941_ (.Y(_02866_),
    .A(_02861_),
    .B(_02864_));
 sg13g2_xor2_1 _08942_ (.B(_02866_),
    .A(_02822_),
    .X(_02867_));
 sg13g2_o21ai_1 _08943_ (.B1(_02839_),
    .Y(_02868_),
    .A1(_02832_),
    .A2(_02840_));
 sg13g2_nand2_1 _08944_ (.Y(_02869_),
    .A(net3293),
    .B(net3085));
 sg13g2_nor2_1 _08945_ (.A(_02691_),
    .B(_02869_),
    .Y(_02870_));
 sg13g2_a22oi_1 _08946_ (.Y(_02871_),
    .B1(net3085),
    .B2(net3301),
    .A2(net3086),
    .A1(net3293));
 sg13g2_nor3_1 _08947_ (.A(net2953),
    .B(_02870_),
    .C(_02871_),
    .Y(_02872_));
 sg13g2_o21ai_1 _08948_ (.B1(net2952),
    .Y(_02873_),
    .A1(_02870_),
    .A2(_02871_));
 sg13g2_nor2b_1 _08949_ (.A(_02872_),
    .B_N(_02873_),
    .Y(_02874_));
 sg13g2_a21oi_1 _08950_ (.A1(_02789_),
    .A2(_02837_),
    .Y(_02875_),
    .B1(_02836_));
 sg13g2_nand2_1 _08951_ (.Y(_02876_),
    .A(net3287),
    .B(net3088));
 sg13g2_nand2_2 _08952_ (.Y(_02877_),
    .A(net3324),
    .B(net3083));
 sg13g2_nor2b_1 _08953_ (.A(net3090),
    .B_N(net3284),
    .Y(_02878_));
 sg13g2_nand2b_1 _08954_ (.Y(_02879_),
    .B(_02878_),
    .A_N(_02877_));
 sg13g2_a21oi_1 _08955_ (.A1(net3327),
    .A2(net3083),
    .Y(_02880_),
    .B1(_02878_));
 sg13g2_xnor2_1 _08956_ (.Y(_02881_),
    .A(net2951),
    .B(_02878_));
 sg13g2_xnor2_1 _08957_ (.Y(_02882_),
    .A(_02876_),
    .B(_02881_));
 sg13g2_nor2b_1 _08958_ (.A(_02875_),
    .B_N(_02882_),
    .Y(_02883_));
 sg13g2_xnor2_1 _08959_ (.Y(_02884_),
    .A(_02875_),
    .B(_02882_));
 sg13g2_xnor2_1 _08960_ (.Y(_02885_),
    .A(_02874_),
    .B(_02884_));
 sg13g2_nor2b_1 _08961_ (.A(_02885_),
    .B_N(_02868_),
    .Y(_02886_));
 sg13g2_nand2b_1 _08962_ (.Y(_02887_),
    .B(_02885_),
    .A_N(_02868_));
 sg13g2_xnor2_1 _08963_ (.Y(_02888_),
    .A(_02868_),
    .B(_02885_));
 sg13g2_xnor2_1 _08964_ (.Y(_02889_),
    .A(_02867_),
    .B(_02888_));
 sg13g2_nand2b_1 _08965_ (.Y(_02890_),
    .B(_02860_),
    .A_N(_02889_));
 sg13g2_xor2_1 _08966_ (.B(_02889_),
    .A(_02860_),
    .X(_02891_));
 sg13g2_xnor2_1 _08967_ (.Y(_02892_),
    .A(_02858_),
    .B(_02891_));
 sg13g2_nand2_1 _08968_ (.Y(_02893_),
    .A(_02857_),
    .B(_02892_));
 sg13g2_nor2_1 _08969_ (.A(_02857_),
    .B(_02892_),
    .Y(_02894_));
 sg13g2_xor2_1 _08970_ (.B(_02892_),
    .A(_02857_),
    .X(_02895_));
 sg13g2_o21ai_1 _08971_ (.B1(_02895_),
    .Y(_02896_),
    .A1(_02851_),
    .A2(_02855_));
 sg13g2_nor3_1 _08972_ (.A(_02851_),
    .B(_02855_),
    .C(_02895_),
    .Y(_02897_));
 sg13g2_nor2_1 _08973_ (.A(net2727),
    .B(_02897_),
    .Y(_02898_));
 sg13g2_a22oi_1 _08974_ (.Y(_02899_),
    .B1(_02896_),
    .B2(_02898_),
    .A2(net2749),
    .A1(net950));
 sg13g2_inv_1 _08975_ (.Y(_00236_),
    .A(_02899_));
 sg13g2_nand2_1 _08976_ (.Y(_02900_),
    .A(net977),
    .B(net2749));
 sg13g2_o21ai_1 _08977_ (.B1(_02865_),
    .Y(_02901_),
    .A1(_02822_),
    .A2(_02866_));
 sg13g2_a21oi_1 _08978_ (.A1(_02867_),
    .A2(_02887_),
    .Y(_02902_),
    .B1(_02886_));
 sg13g2_or2_1 _08979_ (.X(_02903_),
    .B(_02872_),
    .A(_02870_));
 sg13g2_o21ai_1 _08980_ (.B1(net3082),
    .Y(_02904_),
    .A1(net3334),
    .A2(net3307));
 sg13g2_a21oi_1 _08981_ (.A1(net3334),
    .A2(net3307),
    .Y(_02905_),
    .B1(_02904_));
 sg13g2_xor2_1 _08982_ (.B(_02905_),
    .A(_02903_),
    .X(_02906_));
 sg13g2_nor2b_1 _08983_ (.A(_02863_),
    .B_N(_02906_),
    .Y(_02907_));
 sg13g2_xnor2_1 _08984_ (.Y(_02908_),
    .A(_02863_),
    .B(_02906_));
 sg13g2_a21o_1 _08985_ (.A2(_02884_),
    .A1(_02874_),
    .B1(_02883_),
    .X(_02909_));
 sg13g2_nand2_1 _08986_ (.Y(_02910_),
    .A(net3301),
    .B(net3084));
 sg13g2_xor2_1 _08987_ (.B(_02910_),
    .A(_02869_),
    .X(_02911_));
 sg13g2_nand2b_1 _08988_ (.Y(_02912_),
    .B(_02911_),
    .A_N(net2952));
 sg13g2_xnor2_1 _08989_ (.Y(_02913_),
    .A(net2952),
    .B(_02911_));
 sg13g2_inv_1 _08990_ (.Y(_02914_),
    .A(_02913_));
 sg13g2_o21ai_1 _08991_ (.B1(_02879_),
    .Y(_02915_),
    .A1(_02876_),
    .A2(_02880_));
 sg13g2_nor2b_1 _08992_ (.A(net3088),
    .B_N(net3284),
    .Y(_02916_));
 sg13g2_nand2b_1 _08993_ (.Y(_02917_),
    .B(_02916_),
    .A_N(_02877_));
 sg13g2_a21oi_1 _08994_ (.A1(net3324),
    .A2(net3082),
    .Y(_02918_),
    .B1(_02916_));
 sg13g2_xnor2_1 _08995_ (.Y(_02919_),
    .A(_02877_),
    .B(_02916_));
 sg13g2_xnor2_1 _08996_ (.Y(_02920_),
    .A(_02756_),
    .B(_02919_));
 sg13g2_nand2_1 _08997_ (.Y(_02921_),
    .A(_02915_),
    .B(_02920_));
 sg13g2_xnor2_1 _08998_ (.Y(_02922_),
    .A(_02915_),
    .B(_02920_));
 sg13g2_xnor2_1 _08999_ (.Y(_02923_),
    .A(_02914_),
    .B(_02922_));
 sg13g2_nor2b_1 _09000_ (.A(_02923_),
    .B_N(_02909_),
    .Y(_02924_));
 sg13g2_xnor2_1 _09001_ (.Y(_02925_),
    .A(_02909_),
    .B(_02923_));
 sg13g2_xnor2_1 _09002_ (.Y(_02926_),
    .A(_02908_),
    .B(_02925_));
 sg13g2_nor2_1 _09003_ (.A(_02902_),
    .B(_02926_),
    .Y(_02927_));
 sg13g2_xor2_1 _09004_ (.B(_02926_),
    .A(_02902_),
    .X(_02928_));
 sg13g2_xnor2_1 _09005_ (.Y(_02929_),
    .A(_02901_),
    .B(_02928_));
 sg13g2_o21ai_1 _09006_ (.B1(_02890_),
    .Y(_02930_),
    .A1(_02859_),
    .A2(_02891_));
 sg13g2_nor2b_1 _09007_ (.A(_02929_),
    .B_N(_02930_),
    .Y(_02931_));
 sg13g2_xnor2_1 _09008_ (.Y(_02932_),
    .A(_02929_),
    .B(_02930_));
 sg13g2_xor2_1 _09009_ (.B(_02930_),
    .A(_02929_),
    .X(_02933_));
 sg13g2_a22oi_1 _09010_ (.Y(_02934_),
    .B1(_02857_),
    .B2(_02892_),
    .A2(_02850_),
    .A1(_02847_));
 sg13g2_nand3_1 _09011_ (.B(_02896_),
    .C(_02933_),
    .A(_02893_),
    .Y(_02935_));
 sg13g2_a21oi_1 _09012_ (.A1(_02893_),
    .A2(_02896_),
    .Y(_02936_),
    .B1(_02933_));
 sg13g2_nand2_1 _09013_ (.Y(_02937_),
    .A(_02652_),
    .B(_02935_));
 sg13g2_o21ai_1 _09014_ (.B1(_02900_),
    .Y(_00237_),
    .A1(_02936_),
    .A2(_02937_));
 sg13g2_or2_1 _09015_ (.X(_02938_),
    .B(_02936_),
    .A(_02931_));
 sg13g2_a21o_1 _09016_ (.A2(_02928_),
    .A1(_02901_),
    .B1(_02927_),
    .X(_02939_));
 sg13g2_a21o_1 _09017_ (.A2(_02905_),
    .A1(_02903_),
    .B1(_02907_),
    .X(_02940_));
 sg13g2_a21oi_1 _09018_ (.A1(_02908_),
    .A2(_02925_),
    .Y(_02941_),
    .B1(_02924_));
 sg13g2_o21ai_1 _09019_ (.B1(_02912_),
    .Y(_02942_),
    .A1(_02869_),
    .A2(_02910_));
 sg13g2_nand2b_1 _09020_ (.Y(_02943_),
    .B(_02942_),
    .A_N(_02904_));
 sg13g2_inv_1 _09021_ (.Y(_02944_),
    .A(_02943_));
 sg13g2_xnor2_1 _09022_ (.Y(_02945_),
    .A(_02904_),
    .B(_02942_));
 sg13g2_o21ai_1 _09023_ (.B1(_02921_),
    .Y(_02946_),
    .A1(_02914_),
    .A2(_02922_));
 sg13g2_a22oi_1 _09024_ (.Y(_02947_),
    .B1(net3082),
    .B2(net3301),
    .A2(net3084),
    .A1(net3293));
 sg13g2_nand3_1 _09025_ (.B(net3293),
    .C(net3082),
    .A(net3301),
    .Y(_02948_));
 sg13g2_nor2_1 _09026_ (.A(_01150_),
    .B(_02948_),
    .Y(_02949_));
 sg13g2_nor3_1 _09027_ (.A(net2952),
    .B(_02947_),
    .C(_02949_),
    .Y(_02950_));
 sg13g2_o21ai_1 _09028_ (.B1(net2952),
    .Y(_02951_),
    .A1(_02947_),
    .A2(_02949_));
 sg13g2_nand2b_1 _09029_ (.Y(_02952_),
    .B(_02951_),
    .A_N(_02950_));
 sg13g2_o21ai_1 _09030_ (.B1(_02917_),
    .Y(_02953_),
    .A1(_02756_),
    .A2(_02918_));
 sg13g2_nand2_1 _09031_ (.Y(_02954_),
    .A(net3287),
    .B(net3085));
 sg13g2_nor2b_1 _09032_ (.A(net3086),
    .B_N(net3284),
    .Y(_02955_));
 sg13g2_nand2b_1 _09033_ (.Y(_02956_),
    .B(_02955_),
    .A_N(net2951));
 sg13g2_xnor2_1 _09034_ (.Y(_02957_),
    .A(net2951),
    .B(_02955_));
 sg13g2_nand2b_1 _09035_ (.Y(_02958_),
    .B(_02957_),
    .A_N(_02954_));
 sg13g2_xnor2_1 _09036_ (.Y(_02959_),
    .A(_02954_),
    .B(_02957_));
 sg13g2_nand2_1 _09037_ (.Y(_02960_),
    .A(_02953_),
    .B(_02959_));
 sg13g2_xnor2_1 _09038_ (.Y(_02961_),
    .A(_02953_),
    .B(_02959_));
 sg13g2_xnor2_1 _09039_ (.Y(_02962_),
    .A(_02952_),
    .B(_02961_));
 sg13g2_nor2b_1 _09040_ (.A(_02962_),
    .B_N(_02946_),
    .Y(_02963_));
 sg13g2_xnor2_1 _09041_ (.Y(_02964_),
    .A(_02946_),
    .B(_02962_));
 sg13g2_xnor2_1 _09042_ (.Y(_02965_),
    .A(_02945_),
    .B(_02964_));
 sg13g2_nor2_1 _09043_ (.A(_02941_),
    .B(_02965_),
    .Y(_02966_));
 sg13g2_xor2_1 _09044_ (.B(_02965_),
    .A(_02941_),
    .X(_02967_));
 sg13g2_xor2_1 _09045_ (.B(_02967_),
    .A(_02940_),
    .X(_02968_));
 sg13g2_or2_1 _09046_ (.X(_02969_),
    .B(_02968_),
    .A(_02939_));
 sg13g2_nand2_1 _09047_ (.Y(_02970_),
    .A(_02939_),
    .B(_02968_));
 sg13g2_and2_1 _09048_ (.A(_02969_),
    .B(_02970_),
    .X(_02971_));
 sg13g2_xnor2_1 _09049_ (.Y(_02972_),
    .A(_02939_),
    .B(_02968_));
 sg13g2_o21ai_1 _09050_ (.B1(_02652_),
    .Y(_02973_),
    .A1(_02938_),
    .A2(_02971_));
 sg13g2_a21oi_1 _09051_ (.A1(_02938_),
    .A2(_02971_),
    .Y(_02974_),
    .B1(_02973_));
 sg13g2_a21o_1 _09052_ (.A2(net2749),
    .A1(net1013),
    .B1(_02974_),
    .X(_00238_));
 sg13g2_nand2_1 _09053_ (.Y(_02975_),
    .A(net949),
    .B(net2749));
 sg13g2_a21oi_1 _09054_ (.A1(_02945_),
    .A2(_02964_),
    .Y(_02976_),
    .B1(_02963_));
 sg13g2_or2_1 _09055_ (.X(_02977_),
    .B(_02950_),
    .A(_02949_));
 sg13g2_nand2b_1 _09056_ (.Y(_02978_),
    .B(_02977_),
    .A_N(_02904_));
 sg13g2_inv_1 _09057_ (.Y(_02979_),
    .A(_02978_));
 sg13g2_xor2_1 _09058_ (.B(_02977_),
    .A(_02904_),
    .X(_02980_));
 sg13g2_o21ai_1 _09059_ (.B1(_02960_),
    .Y(_02981_),
    .A1(_02952_),
    .A2(_02961_));
 sg13g2_nand2_1 _09060_ (.Y(_02982_),
    .A(_02956_),
    .B(_02958_));
 sg13g2_nand2_1 _09061_ (.Y(_02983_),
    .A(net3287),
    .B(net3084));
 sg13g2_nand2b_1 _09062_ (.Y(_02984_),
    .B(net3284),
    .A_N(net3085));
 sg13g2_xor2_1 _09063_ (.B(_02984_),
    .A(net2951),
    .X(_02985_));
 sg13g2_nand2b_1 _09064_ (.Y(_02986_),
    .B(_02985_),
    .A_N(_02983_));
 sg13g2_xnor2_1 _09065_ (.Y(_02987_),
    .A(_02983_),
    .B(_02985_));
 sg13g2_xnor2_1 _09066_ (.Y(_02988_),
    .A(_02982_),
    .B(_02987_));
 sg13g2_o21ai_1 _09067_ (.B1(net3082),
    .Y(_02989_),
    .A1(net3301),
    .A2(net3293));
 sg13g2_nor2b_1 _09068_ (.A(_02989_),
    .B_N(_02948_),
    .Y(_02990_));
 sg13g2_xnor2_1 _09069_ (.Y(_02991_),
    .A(net2952),
    .B(_02990_));
 sg13g2_inv_1 _09070_ (.Y(_02992_),
    .A(_02991_));
 sg13g2_nor2_1 _09071_ (.A(_02988_),
    .B(_02992_),
    .Y(_02993_));
 sg13g2_xnor2_1 _09072_ (.Y(_02994_),
    .A(_02988_),
    .B(_02991_));
 sg13g2_xnor2_1 _09073_ (.Y(_02995_),
    .A(_02981_),
    .B(_02994_));
 sg13g2_nor2_1 _09074_ (.A(_02980_),
    .B(_02995_),
    .Y(_02996_));
 sg13g2_xnor2_1 _09075_ (.Y(_02997_),
    .A(_02980_),
    .B(_02995_));
 sg13g2_nor2_1 _09076_ (.A(_02976_),
    .B(_02997_),
    .Y(_02998_));
 sg13g2_xor2_1 _09077_ (.B(_02997_),
    .A(_02976_),
    .X(_02999_));
 sg13g2_xnor2_1 _09078_ (.Y(_03000_),
    .A(_02943_),
    .B(_02999_));
 sg13g2_a21oi_1 _09079_ (.A1(_02940_),
    .A2(_02967_),
    .Y(_03001_),
    .B1(_02966_));
 sg13g2_nor2b_1 _09080_ (.A(_03001_),
    .B_N(_03000_),
    .Y(_03002_));
 sg13g2_inv_1 _09081_ (.Y(_03003_),
    .A(_03002_));
 sg13g2_xor2_1 _09082_ (.B(_03001_),
    .A(_03000_),
    .X(_03004_));
 sg13g2_inv_1 _09083_ (.Y(_03005_),
    .A(_03004_));
 sg13g2_nand2_1 _09084_ (.Y(_03006_),
    .A(_02931_),
    .B(_02969_));
 sg13g2_or4_1 _09085_ (.A(_02894_),
    .B(_02933_),
    .C(_02934_),
    .D(_02972_),
    .X(_03007_));
 sg13g2_nand3_1 _09086_ (.B(_03006_),
    .C(_03007_),
    .A(_02970_),
    .Y(_03008_));
 sg13g2_and4_1 _09087_ (.A(_02855_),
    .B(_02895_),
    .C(_02932_),
    .D(_02971_),
    .X(_03009_));
 sg13g2_nor3_1 _09088_ (.A(_03005_),
    .B(_03008_),
    .C(_03009_),
    .Y(_03010_));
 sg13g2_o21ai_1 _09089_ (.B1(_03005_),
    .Y(_03011_),
    .A1(_03008_),
    .A2(_03009_));
 sg13g2_nand2_1 _09090_ (.Y(_03012_),
    .A(_02652_),
    .B(_03011_));
 sg13g2_o21ai_1 _09091_ (.B1(_02975_),
    .Y(_00239_),
    .A1(_03010_),
    .A2(_03012_));
 sg13g2_a21oi_1 _09092_ (.A1(_02981_),
    .A2(_02994_),
    .Y(_03013_),
    .B1(_02996_));
 sg13g2_a21oi_1 _09093_ (.A1(_02982_),
    .A2(_02987_),
    .Y(_03014_),
    .B1(_02993_));
 sg13g2_o21ai_1 _09094_ (.B1(_02986_),
    .Y(_03015_),
    .A1(net2951),
    .A2(_02984_));
 sg13g2_and2_1 _09095_ (.A(net3287),
    .B(net3082),
    .X(_03016_));
 sg13g2_nand2_1 _09096_ (.Y(_03017_),
    .A(net3284),
    .B(_01150_));
 sg13g2_nor2_1 _09097_ (.A(net2951),
    .B(_03017_),
    .Y(_03018_));
 sg13g2_xor2_1 _09098_ (.B(_03017_),
    .A(net2951),
    .X(_03019_));
 sg13g2_xor2_1 _09099_ (.B(_03019_),
    .A(_03016_),
    .X(_03020_));
 sg13g2_nand2_1 _09100_ (.Y(_03021_),
    .A(_03015_),
    .B(_03020_));
 sg13g2_xnor2_1 _09101_ (.Y(_03022_),
    .A(_03015_),
    .B(_03020_));
 sg13g2_xnor2_1 _09102_ (.Y(_03023_),
    .A(_02992_),
    .B(_03022_));
 sg13g2_nor2_1 _09103_ (.A(_03014_),
    .B(_03023_),
    .Y(_03024_));
 sg13g2_xnor2_1 _09104_ (.Y(_03025_),
    .A(_03014_),
    .B(_03023_));
 sg13g2_o21ai_1 _09105_ (.B1(_02948_),
    .Y(_03026_),
    .A1(net2952),
    .A2(_02989_));
 sg13g2_nand2b_2 _09106_ (.Y(_03027_),
    .B(_03026_),
    .A_N(_02904_));
 sg13g2_nand2b_1 _09107_ (.Y(_03028_),
    .B(_02904_),
    .A_N(_03026_));
 sg13g2_nand2_2 _09108_ (.Y(_03029_),
    .A(_03027_),
    .B(_03028_));
 sg13g2_nor2_1 _09109_ (.A(_03025_),
    .B(_03029_),
    .Y(_03030_));
 sg13g2_xor2_1 _09110_ (.B(_03029_),
    .A(_03025_),
    .X(_03031_));
 sg13g2_nor2b_1 _09111_ (.A(_03013_),
    .B_N(_03031_),
    .Y(_03032_));
 sg13g2_xnor2_1 _09112_ (.Y(_03033_),
    .A(_03013_),
    .B(_03031_));
 sg13g2_xnor2_1 _09113_ (.Y(_03034_),
    .A(_02978_),
    .B(_03033_));
 sg13g2_a21oi_1 _09114_ (.A1(_02944_),
    .A2(_02999_),
    .Y(_03035_),
    .B1(_02998_));
 sg13g2_inv_1 _09115_ (.Y(_03036_),
    .A(_03035_));
 sg13g2_xnor2_1 _09116_ (.Y(_03037_),
    .A(_03034_),
    .B(_03036_));
 sg13g2_nand3_1 _09117_ (.B(_03011_),
    .C(_03037_),
    .A(_03003_),
    .Y(_03038_));
 sg13g2_nor2_1 _09118_ (.A(_03011_),
    .B(_03037_),
    .Y(_03039_));
 sg13g2_nor2_1 _09119_ (.A(_03003_),
    .B(_03037_),
    .Y(_03040_));
 sg13g2_nor3_1 _09120_ (.A(net2727),
    .B(_03039_),
    .C(_03040_),
    .Y(_03041_));
 sg13g2_a22oi_1 _09121_ (.Y(_03042_),
    .B1(_03038_),
    .B2(_03041_),
    .A2(net2749),
    .A1(net1004));
 sg13g2_inv_1 _09122_ (.Y(_00240_),
    .A(_03042_));
 sg13g2_nand2_1 _09123_ (.Y(_03043_),
    .A(net1002),
    .B(net2749));
 sg13g2_a21oi_1 _09124_ (.A1(_03034_),
    .A2(_03036_),
    .Y(_03044_),
    .B1(_03040_));
 sg13g2_o21ai_1 _09125_ (.B1(_03044_),
    .Y(_03045_),
    .A1(_03011_),
    .A2(_03037_));
 sg13g2_nor2_1 _09126_ (.A(_03024_),
    .B(_03030_),
    .Y(_03046_));
 sg13g2_o21ai_1 _09127_ (.B1(_03021_),
    .Y(_03047_),
    .A1(_02992_),
    .A2(_03022_));
 sg13g2_a21oi_1 _09128_ (.A1(net3284),
    .A2(_01151_),
    .Y(_03048_),
    .B1(_03016_));
 sg13g2_a221oi_1 _09129_ (.B2(net2951),
    .C1(_03018_),
    .B1(_03048_),
    .A1(_03016_),
    .Y(_03049_),
    .A2(_03019_));
 sg13g2_a21oi_2 _09130_ (.B1(_03049_),
    .Y(_03050_),
    .A2(_03016_),
    .A1(net3324));
 sg13g2_nand2_1 _09131_ (.Y(_03051_),
    .A(_02992_),
    .B(_03050_));
 sg13g2_xnor2_1 _09132_ (.Y(_03052_),
    .A(_02991_),
    .B(_03050_));
 sg13g2_nand2_1 _09133_ (.Y(_03053_),
    .A(_03047_),
    .B(_03052_));
 sg13g2_xnor2_1 _09134_ (.Y(_03054_),
    .A(_03047_),
    .B(_03052_));
 sg13g2_xnor2_1 _09135_ (.Y(_03055_),
    .A(_03029_),
    .B(_03054_));
 sg13g2_xor2_1 _09136_ (.B(_03055_),
    .A(_03046_),
    .X(_03056_));
 sg13g2_nand2b_1 _09137_ (.Y(_03057_),
    .B(_03056_),
    .A_N(_03027_));
 sg13g2_xor2_1 _09138_ (.B(_03056_),
    .A(_03027_),
    .X(_03058_));
 sg13g2_a21oi_1 _09139_ (.A1(_02979_),
    .A2(_03033_),
    .Y(_03059_),
    .B1(_03032_));
 sg13g2_xor2_1 _09140_ (.B(_03059_),
    .A(_03058_),
    .X(_03060_));
 sg13g2_nor2_1 _09141_ (.A(_03045_),
    .B(_03060_),
    .Y(_03061_));
 sg13g2_a21o_1 _09142_ (.A2(_03060_),
    .A1(_03045_),
    .B1(net2727),
    .X(_03062_));
 sg13g2_o21ai_1 _09143_ (.B1(_03043_),
    .Y(_00241_),
    .A1(_03061_),
    .A2(_03062_));
 sg13g2_nand2_1 _09144_ (.Y(_03063_),
    .A(net3194),
    .B(net2749));
 sg13g2_o21ai_1 _09145_ (.B1(_03057_),
    .Y(_03064_),
    .A1(_03046_),
    .A2(_03055_));
 sg13g2_o21ai_1 _09146_ (.B1(_03053_),
    .Y(_03065_),
    .A1(_03029_),
    .A2(_03054_));
 sg13g2_xnor2_1 _09147_ (.Y(_03066_),
    .A(_03028_),
    .B(_03051_));
 sg13g2_xor2_1 _09148_ (.B(_03066_),
    .A(_03065_),
    .X(_03067_));
 sg13g2_xnor2_1 _09149_ (.Y(_03068_),
    .A(_03064_),
    .B(_03067_));
 sg13g2_o21ai_1 _09150_ (.B1(_03068_),
    .Y(_03069_),
    .A1(_03058_),
    .A2(_03059_));
 sg13g2_o21ai_1 _09151_ (.B1(_03063_),
    .Y(_00242_),
    .A1(_03062_),
    .A2(_03069_));
 sg13g2_nand3_1 _09152_ (.B(_00034_),
    .C(_01937_),
    .A(\u_toplayer.delayed_done_layer2 ),
    .Y(_03070_));
 sg13g2_a21oi_1 _09153_ (.A1(net3136),
    .A2(_01067_),
    .Y(_03071_),
    .B1(net3114));
 sg13g2_o21ai_1 _09154_ (.B1(_03071_),
    .Y(_03072_),
    .A1(net3136),
    .A2(\u_toplayer.reg_layer2[96] ));
 sg13g2_a22oi_1 _09155_ (.Y(_03073_),
    .B1(net2973),
    .B2(\u_toplayer.reg_layer2[112] ),
    .A2(net3006),
    .A1(\u_toplayer.reg_layer2[120] ));
 sg13g2_nand3_1 _09156_ (.B(_03072_),
    .C(_03073_),
    .A(net3103),
    .Y(_03074_));
 sg13g2_a21oi_1 _09157_ (.A1(net3136),
    .A2(_01066_),
    .Y(_03075_),
    .B1(net3111));
 sg13g2_o21ai_1 _09158_ (.B1(_03075_),
    .Y(_03076_),
    .A1(net3124),
    .A2(\u_toplayer.reg_layer2[64] ));
 sg13g2_a22oi_1 _09159_ (.Y(_03077_),
    .B1(net2968),
    .B2(\u_toplayer.reg_layer2[80] ),
    .A2(net3001),
    .A1(\u_toplayer.reg_layer2[88] ));
 sg13g2_nand3_1 _09160_ (.B(_03076_),
    .C(_03077_),
    .A(net3017),
    .Y(_03078_));
 sg13g2_nand3_1 _09161_ (.B(_03074_),
    .C(_03078_),
    .A(net3101),
    .Y(_03079_));
 sg13g2_nor2b_1 _09162_ (.A(net3121),
    .B_N(\u_toplayer.reg_layer2[0] ),
    .Y(_03080_));
 sg13g2_a21oi_1 _09163_ (.A1(net3122),
    .A2(\u_toplayer.reg_layer2[8] ),
    .Y(_03081_),
    .B1(_03080_));
 sg13g2_a22oi_1 _09164_ (.Y(_03082_),
    .B1(net2966),
    .B2(\u_toplayer.reg_layer2[16] ),
    .A2(net2999),
    .A1(\u_toplayer.reg_layer2[24] ));
 sg13g2_o21ai_1 _09165_ (.B1(_03082_),
    .Y(_03083_),
    .A1(net3108),
    .A2(_03081_));
 sg13g2_nand2b_1 _09166_ (.Y(_03084_),
    .B(net3132),
    .A_N(\u_toplayer.reg_layer2[40] ));
 sg13g2_o21ai_1 _09167_ (.B1(_03084_),
    .Y(_03085_),
    .A1(net3129),
    .A2(\u_toplayer.reg_layer2[32] ));
 sg13g2_a22oi_1 _09168_ (.Y(_03086_),
    .B1(net2971),
    .B2(\u_toplayer.reg_layer2[48] ),
    .A2(net3004),
    .A1(\u_toplayer.reg_layer2[56] ));
 sg13g2_o21ai_1 _09169_ (.B1(_03086_),
    .Y(_03087_),
    .A1(net3108),
    .A2(_03085_));
 sg13g2_a221oi_1 _09170_ (.B2(net2936),
    .C1(net3096),
    .B1(_03087_),
    .A1(net3008),
    .Y(_03088_),
    .A2(_03083_));
 sg13g2_a21oi_1 _09171_ (.A1(net3136),
    .A2(_01069_),
    .Y(_03089_),
    .B1(net3114));
 sg13g2_o21ai_1 _09172_ (.B1(_03089_),
    .Y(_03090_),
    .A1(net3136),
    .A2(\u_toplayer.reg_layer2[224] ));
 sg13g2_a221oi_1 _09173_ (.B2(\u_toplayer.reg_layer2[240] ),
    .C1(net3017),
    .B1(net2973),
    .A1(\u_toplayer.reg_layer2[248] ),
    .Y(_03091_),
    .A2(net3006));
 sg13g2_a21oi_1 _09174_ (.A1(net3136),
    .A2(_01068_),
    .Y(_03092_),
    .B1(net3114));
 sg13g2_o21ai_1 _09175_ (.B1(_03092_),
    .Y(_03093_),
    .A1(net3124),
    .A2(\u_toplayer.reg_layer2[192] ));
 sg13g2_a221oi_1 _09176_ (.B2(\u_toplayer.reg_layer2[208] ),
    .C1(net3102),
    .B1(net2968),
    .A1(\u_toplayer.reg_layer2[216] ),
    .Y(_03094_),
    .A2(net3003));
 sg13g2_a22oi_1 _09177_ (.Y(_03095_),
    .B1(_03093_),
    .B2(_03094_),
    .A2(_03091_),
    .A1(_03090_));
 sg13g2_nand2_1 _09178_ (.Y(_03096_),
    .A(net3099),
    .B(_03095_));
 sg13g2_nand2b_1 _09179_ (.Y(_03097_),
    .B(net3120),
    .A_N(\u_toplayer.reg_layer2[136] ));
 sg13g2_o21ai_1 _09180_ (.B1(_03097_),
    .Y(_03098_),
    .A1(net3117),
    .A2(\u_toplayer.reg_layer2[128] ));
 sg13g2_a22oi_1 _09181_ (.Y(_03099_),
    .B1(net2966),
    .B2(\u_toplayer.reg_layer2[144] ),
    .A2(net2999),
    .A1(\u_toplayer.reg_layer2[152] ));
 sg13g2_o21ai_1 _09182_ (.B1(_03099_),
    .Y(_03100_),
    .A1(net3106),
    .A2(_03098_));
 sg13g2_nand2b_1 _09183_ (.Y(_03101_),
    .B(net3132),
    .A_N(\u_toplayer.reg_layer2[168] ));
 sg13g2_o21ai_1 _09184_ (.B1(_03101_),
    .Y(_03102_),
    .A1(net3132),
    .A2(\u_toplayer.reg_layer2[160] ));
 sg13g2_a22oi_1 _09185_ (.Y(_03103_),
    .B1(net2971),
    .B2(\u_toplayer.reg_layer2[176] ),
    .A2(net3004),
    .A1(\u_toplayer.reg_layer2[184] ));
 sg13g2_o21ai_1 _09186_ (.B1(_03103_),
    .Y(_03104_),
    .A1(net3108),
    .A2(_03102_));
 sg13g2_a22oi_1 _09187_ (.Y(_03105_),
    .B1(_03104_),
    .B2(net2936),
    .A2(_03100_),
    .A1(net3009));
 sg13g2_and2_1 _09188_ (.A(net3097),
    .B(_03105_),
    .X(_03106_));
 sg13g2_a221oi_1 _09189_ (.B2(_03106_),
    .C1(_03070_),
    .B1(_03096_),
    .A1(_03079_),
    .Y(_03107_),
    .A2(_03088_));
 sg13g2_a21o_1 _09190_ (.A2(_01938_),
    .A1(net1022),
    .B1(_03107_),
    .X(_00324_));
 sg13g2_a21oi_1 _09191_ (.A1(net3137),
    .A2(_01073_),
    .Y(_03108_),
    .B1(net3114));
 sg13g2_o21ai_1 _09192_ (.B1(_03108_),
    .Y(_03109_),
    .A1(net3136),
    .A2(\u_toplayer.reg_layer2[225] ));
 sg13g2_a22oi_1 _09193_ (.Y(_03110_),
    .B1(net2973),
    .B2(\u_toplayer.reg_layer2[241] ),
    .A2(net3005),
    .A1(\u_toplayer.reg_layer2[249] ));
 sg13g2_nand3_1 _09194_ (.B(_03109_),
    .C(_03110_),
    .A(net3103),
    .Y(_03111_));
 sg13g2_a21oi_1 _09195_ (.A1(net3125),
    .A2(_01072_),
    .Y(_03112_),
    .B1(net3112));
 sg13g2_o21ai_1 _09196_ (.B1(_03112_),
    .Y(_03113_),
    .A1(net3125),
    .A2(\u_toplayer.reg_layer2[193] ));
 sg13g2_a22oi_1 _09197_ (.Y(_03114_),
    .B1(net2968),
    .B2(\u_toplayer.reg_layer2[209] ),
    .A2(net3001),
    .A1(\u_toplayer.reg_layer2[217] ));
 sg13g2_nand3_1 _09198_ (.B(_03113_),
    .C(_03114_),
    .A(net3017),
    .Y(_03115_));
 sg13g2_nand3_1 _09199_ (.B(_03111_),
    .C(_03115_),
    .A(net3101),
    .Y(_03116_));
 sg13g2_nor2b_1 _09200_ (.A(net3130),
    .B_N(\u_toplayer.reg_layer2[161] ),
    .Y(_03117_));
 sg13g2_a21oi_1 _09201_ (.A1(net3129),
    .A2(\u_toplayer.reg_layer2[169] ),
    .Y(_03118_),
    .B1(_03117_));
 sg13g2_a22oi_1 _09202_ (.Y(_03119_),
    .B1(net2971),
    .B2(\u_toplayer.reg_layer2[177] ),
    .A2(net3004),
    .A1(\u_toplayer.reg_layer2[185] ));
 sg13g2_o21ai_1 _09203_ (.B1(_03119_),
    .Y(_03120_),
    .A1(net3109),
    .A2(_03118_));
 sg13g2_nand2b_1 _09204_ (.Y(_03121_),
    .B(net3118),
    .A_N(\u_toplayer.reg_layer2[137] ));
 sg13g2_o21ai_1 _09205_ (.B1(_03121_),
    .Y(_03122_),
    .A1(net3118),
    .A2(\u_toplayer.reg_layer2[129] ));
 sg13g2_a22oi_1 _09206_ (.Y(_03123_),
    .B1(net2965),
    .B2(\u_toplayer.reg_layer2[145] ),
    .A2(net2998),
    .A1(\u_toplayer.reg_layer2[153] ));
 sg13g2_o21ai_1 _09207_ (.B1(_03123_),
    .Y(_03124_),
    .A1(net3107),
    .A2(_03122_));
 sg13g2_a22oi_1 _09208_ (.Y(_03125_),
    .B1(_03124_),
    .B2(net3010),
    .A2(_03120_),
    .A1(net2937));
 sg13g2_nand3_1 _09209_ (.B(_03116_),
    .C(_03125_),
    .A(net3098),
    .Y(_03126_));
 sg13g2_a21oi_1 _09210_ (.A1(net3137),
    .A2(_01071_),
    .Y(_03127_),
    .B1(net3114));
 sg13g2_o21ai_1 _09211_ (.B1(_03127_),
    .Y(_03128_),
    .A1(net3136),
    .A2(\u_toplayer.reg_layer2[97] ));
 sg13g2_a22oi_1 _09212_ (.Y(_03129_),
    .B1(net2972),
    .B2(\u_toplayer.reg_layer2[113] ),
    .A2(net3005),
    .A1(\u_toplayer.reg_layer2[121] ));
 sg13g2_nand3_1 _09213_ (.B(_03128_),
    .C(_03129_),
    .A(net3103),
    .Y(_03130_));
 sg13g2_a21oi_1 _09214_ (.A1(net3126),
    .A2(_01070_),
    .Y(_03131_),
    .B1(net3116));
 sg13g2_o21ai_1 _09215_ (.B1(_03131_),
    .Y(_03132_),
    .A1(net3125),
    .A2(\u_toplayer.reg_layer2[65] ));
 sg13g2_a22oi_1 _09216_ (.Y(_03133_),
    .B1(net2968),
    .B2(\u_toplayer.reg_layer2[81] ),
    .A2(net3001),
    .A1(\u_toplayer.reg_layer2[89] ));
 sg13g2_nand3_1 _09217_ (.B(_03132_),
    .C(_03133_),
    .A(net3017),
    .Y(_03134_));
 sg13g2_nand3_1 _09218_ (.B(_03130_),
    .C(_03134_),
    .A(net3101),
    .Y(_03135_));
 sg13g2_nand2b_1 _09219_ (.Y(_03136_),
    .B(net3135),
    .A_N(\u_toplayer.reg_layer2[41] ));
 sg13g2_o21ai_1 _09220_ (.B1(_03136_),
    .Y(_03137_),
    .A1(net3135),
    .A2(\u_toplayer.reg_layer2[33] ));
 sg13g2_a22oi_1 _09221_ (.Y(_03138_),
    .B1(net2972),
    .B2(\u_toplayer.reg_layer2[49] ),
    .A2(net3005),
    .A1(\u_toplayer.reg_layer2[57] ));
 sg13g2_o21ai_1 _09222_ (.B1(_03138_),
    .Y(_03139_),
    .A1(net3109),
    .A2(_03137_));
 sg13g2_nor2b_1 _09223_ (.A(net3119),
    .B_N(\u_toplayer.reg_layer2[1] ),
    .Y(_03140_));
 sg13g2_a21oi_1 _09224_ (.A1(net3119),
    .A2(\u_toplayer.reg_layer2[9] ),
    .Y(_03141_),
    .B1(_03140_));
 sg13g2_a22oi_1 _09225_ (.Y(_03142_),
    .B1(net2965),
    .B2(\u_toplayer.reg_layer2[17] ),
    .A2(net2998),
    .A1(\u_toplayer.reg_layer2[25] ));
 sg13g2_o21ai_1 _09226_ (.B1(_03142_),
    .Y(_03143_),
    .A1(net3107),
    .A2(_03141_));
 sg13g2_a221oi_1 _09227_ (.B2(net3009),
    .C1(net3096),
    .B1(_03143_),
    .A1(net2935),
    .Y(_03144_),
    .A2(_03139_));
 sg13g2_a21oi_1 _09228_ (.A1(_03135_),
    .A2(_03144_),
    .Y(_03145_),
    .B1(_03070_));
 sg13g2_a22oi_1 _09229_ (.Y(_03146_),
    .B1(_03126_),
    .B2(_03145_),
    .A2(_01938_),
    .A1(net3177));
 sg13g2_inv_1 _09230_ (.Y(_00325_),
    .A(_03146_));
 sg13g2_a21oi_1 _09231_ (.A1(net3137),
    .A2(_01074_),
    .Y(_03147_),
    .B1(net3114));
 sg13g2_o21ai_1 _09232_ (.B1(_03147_),
    .Y(_03148_),
    .A1(net3125),
    .A2(\u_toplayer.reg_layer2[66] ));
 sg13g2_a22oi_1 _09233_ (.Y(_03149_),
    .B1(net2968),
    .B2(\u_toplayer.reg_layer2[82] ),
    .A2(net3001),
    .A1(\u_toplayer.reg_layer2[90] ));
 sg13g2_nand3_1 _09234_ (.B(_03148_),
    .C(_03149_),
    .A(_01036_),
    .Y(_03150_));
 sg13g2_a21oi_1 _09235_ (.A1(net3141),
    .A2(_01075_),
    .Y(_03151_),
    .B1(net3115));
 sg13g2_o21ai_1 _09236_ (.B1(_03151_),
    .Y(_03152_),
    .A1(net3141),
    .A2(\u_toplayer.reg_layer2[98] ));
 sg13g2_a22oi_1 _09237_ (.Y(_03153_),
    .B1(net2973),
    .B2(\u_toplayer.reg_layer2[114] ),
    .A2(net3007),
    .A1(\u_toplayer.reg_layer2[122] ));
 sg13g2_nand3_1 _09238_ (.B(_03152_),
    .C(_03153_),
    .A(net3104),
    .Y(_03154_));
 sg13g2_nand3_1 _09239_ (.B(_03150_),
    .C(_03154_),
    .A(net3100),
    .Y(_03155_));
 sg13g2_nor2b_1 _09240_ (.A(net3121),
    .B_N(\u_toplayer.reg_layer2[2] ),
    .Y(_03156_));
 sg13g2_a21oi_1 _09241_ (.A1(net3121),
    .A2(\u_toplayer.reg_layer2[10] ),
    .Y(_03157_),
    .B1(_03156_));
 sg13g2_a22oi_1 _09242_ (.Y(_03158_),
    .B1(net2966),
    .B2(\u_toplayer.reg_layer2[18] ),
    .A2(net2999),
    .A1(\u_toplayer.reg_layer2[26] ));
 sg13g2_o21ai_1 _09243_ (.B1(_03158_),
    .Y(_03159_),
    .A1(net3110),
    .A2(_03157_));
 sg13g2_nand2b_1 _09244_ (.Y(_03160_),
    .B(net3132),
    .A_N(\u_toplayer.reg_layer2[42] ));
 sg13g2_o21ai_1 _09245_ (.B1(_03160_),
    .Y(_03161_),
    .A1(net3132),
    .A2(\u_toplayer.reg_layer2[34] ));
 sg13g2_a22oi_1 _09246_ (.Y(_03162_),
    .B1(net2971),
    .B2(\u_toplayer.reg_layer2[50] ),
    .A2(net3004),
    .A1(\u_toplayer.reg_layer2[58] ));
 sg13g2_o21ai_1 _09247_ (.B1(_03162_),
    .Y(_03163_),
    .A1(net3108),
    .A2(_03161_));
 sg13g2_a221oi_1 _09248_ (.B2(net2936),
    .C1(net3096),
    .B1(_03163_),
    .A1(net3008),
    .Y(_03164_),
    .A2(_03159_));
 sg13g2_a21oi_1 _09249_ (.A1(net3137),
    .A2(_01076_),
    .Y(_03165_),
    .B1(net3114));
 sg13g2_o21ai_1 _09250_ (.B1(_03165_),
    .Y(_03166_),
    .A1(net3125),
    .A2(\u_toplayer.reg_layer2[194] ));
 sg13g2_a22oi_1 _09251_ (.Y(_03167_),
    .B1(net2968),
    .B2(\u_toplayer.reg_layer2[210] ),
    .A2(net3001),
    .A1(\u_toplayer.reg_layer2[218] ));
 sg13g2_nand3_1 _09252_ (.B(_03166_),
    .C(_03167_),
    .A(net3017),
    .Y(_03168_));
 sg13g2_a21oi_1 _09253_ (.A1(net3140),
    .A2(_01077_),
    .Y(_03169_),
    .B1(net3113));
 sg13g2_o21ai_1 _09254_ (.B1(_03169_),
    .Y(_03170_),
    .A1(net3140),
    .A2(\u_toplayer.reg_layer2[226] ));
 sg13g2_a22oi_1 _09255_ (.Y(_03171_),
    .B1(net2973),
    .B2(\u_toplayer.reg_layer2[242] ),
    .A2(net3007),
    .A1(\u_toplayer.reg_layer2[250] ));
 sg13g2_nand3_1 _09256_ (.B(_03170_),
    .C(_03171_),
    .A(net3103),
    .Y(_03172_));
 sg13g2_nand3_1 _09257_ (.B(_03168_),
    .C(_03172_),
    .A(net3100),
    .Y(_03173_));
 sg13g2_nand2b_1 _09258_ (.Y(_03174_),
    .B(net3118),
    .A_N(\u_toplayer.reg_layer2[138] ));
 sg13g2_o21ai_1 _09259_ (.B1(_03174_),
    .Y(_03175_),
    .A1(net3118),
    .A2(\u_toplayer.reg_layer2[130] ));
 sg13g2_a22oi_1 _09260_ (.Y(_03176_),
    .B1(net2965),
    .B2(\u_toplayer.reg_layer2[146] ),
    .A2(net3000),
    .A1(\u_toplayer.reg_layer2[154] ));
 sg13g2_o21ai_1 _09261_ (.B1(_03176_),
    .Y(_03177_),
    .A1(net3110),
    .A2(_03175_));
 sg13g2_nor2b_1 _09262_ (.A(net3133),
    .B_N(\u_toplayer.reg_layer2[162] ),
    .Y(_03178_));
 sg13g2_a21oi_1 _09263_ (.A1(net3133),
    .A2(\u_toplayer.reg_layer2[170] ),
    .Y(_03179_),
    .B1(_03178_));
 sg13g2_a22oi_1 _09264_ (.Y(_03180_),
    .B1(net2971),
    .B2(\u_toplayer.reg_layer2[178] ),
    .A2(net3004),
    .A1(\u_toplayer.reg_layer2[186] ));
 sg13g2_o21ai_1 _09265_ (.B1(_03180_),
    .Y(_03181_),
    .A1(net3108),
    .A2(_03179_));
 sg13g2_a22oi_1 _09266_ (.Y(_03182_),
    .B1(_03181_),
    .B2(net2935),
    .A2(_03177_),
    .A1(net3008));
 sg13g2_and2_1 _09267_ (.A(net3096),
    .B(_03182_),
    .X(_03183_));
 sg13g2_a221oi_1 _09268_ (.B2(_03183_),
    .C1(_03070_),
    .B1(_03173_),
    .A1(_03155_),
    .Y(_03184_),
    .A2(_03164_));
 sg13g2_a21o_1 _09269_ (.A2(net2817),
    .A1(net3175),
    .B1(_03184_),
    .X(_00326_));
 sg13g2_a21oi_1 _09270_ (.A1(net3140),
    .A2(_01081_),
    .Y(_03185_),
    .B1(net3113));
 sg13g2_o21ai_1 _09271_ (.B1(_03185_),
    .Y(_03186_),
    .A1(net3140),
    .A2(\u_toplayer.reg_layer2[227] ));
 sg13g2_a22oi_1 _09272_ (.Y(_03187_),
    .B1(net2973),
    .B2(\u_toplayer.reg_layer2[243] ),
    .A2(net3006),
    .A1(\u_toplayer.reg_layer2[251] ));
 sg13g2_nand3_1 _09273_ (.B(_03186_),
    .C(_03187_),
    .A(net3103),
    .Y(_03188_));
 sg13g2_a21oi_1 _09274_ (.A1(net3125),
    .A2(_01080_),
    .Y(_03189_),
    .B1(net3112));
 sg13g2_o21ai_1 _09275_ (.B1(_03189_),
    .Y(_03190_),
    .A1(net3125),
    .A2(\u_toplayer.reg_layer2[195] ));
 sg13g2_a22oi_1 _09276_ (.Y(_03191_),
    .B1(net2969),
    .B2(\u_toplayer.reg_layer2[211] ),
    .A2(net3002),
    .A1(\u_toplayer.reg_layer2[219] ));
 sg13g2_nand3_1 _09277_ (.B(_03190_),
    .C(_03191_),
    .A(net3018),
    .Y(_03192_));
 sg13g2_nand3_1 _09278_ (.B(_03188_),
    .C(_03192_),
    .A(net3100),
    .Y(_03193_));
 sg13g2_nor2b_1 _09279_ (.A(net3132),
    .B_N(\u_toplayer.reg_layer2[163] ),
    .Y(_03194_));
 sg13g2_a21oi_2 _09280_ (.B1(_03194_),
    .Y(_03195_),
    .A2(\u_toplayer.reg_layer2[171] ),
    .A1(net3134));
 sg13g2_a22oi_1 _09281_ (.Y(_03196_),
    .B1(net2972),
    .B2(\u_toplayer.reg_layer2[179] ),
    .A2(net3005),
    .A1(\u_toplayer.reg_layer2[187] ));
 sg13g2_o21ai_1 _09282_ (.B1(_03196_),
    .Y(_03197_),
    .A1(net3115),
    .A2(_03195_));
 sg13g2_nand2b_1 _09283_ (.Y(_03198_),
    .B(net3119),
    .A_N(\u_toplayer.reg_layer2[139] ));
 sg13g2_o21ai_1 _09284_ (.B1(_03198_),
    .Y(_03199_),
    .A1(net3118),
    .A2(\u_toplayer.reg_layer2[131] ));
 sg13g2_a22oi_1 _09285_ (.Y(_03200_),
    .B1(net2965),
    .B2(\u_toplayer.reg_layer2[147] ),
    .A2(net2998),
    .A1(\u_toplayer.reg_layer2[155] ));
 sg13g2_o21ai_1 _09286_ (.B1(_03200_),
    .Y(_03201_),
    .A1(net3110),
    .A2(_03199_));
 sg13g2_a22oi_1 _09287_ (.Y(_03202_),
    .B1(_03201_),
    .B2(net3010),
    .A2(_03197_),
    .A1(net2937));
 sg13g2_nand3_1 _09288_ (.B(_03193_),
    .C(_03202_),
    .A(net3098),
    .Y(_03203_));
 sg13g2_a21oi_1 _09289_ (.A1(net3126),
    .A2(_01078_),
    .Y(_03204_),
    .B1(net3111));
 sg13g2_o21ai_1 _09290_ (.B1(_03204_),
    .Y(_03205_),
    .A1(net3126),
    .A2(\u_toplayer.reg_layer2[67] ));
 sg13g2_a22oi_1 _09291_ (.Y(_03206_),
    .B1(net2970),
    .B2(\u_toplayer.reg_layer2[83] ),
    .A2(net3003),
    .A1(\u_toplayer.reg_layer2[91] ));
 sg13g2_nand3_1 _09292_ (.B(_03205_),
    .C(_03206_),
    .A(net3018),
    .Y(_03207_));
 sg13g2_a21oi_1 _09293_ (.A1(net3140),
    .A2(_01079_),
    .Y(_03208_),
    .B1(net3113));
 sg13g2_o21ai_1 _09294_ (.B1(_03208_),
    .Y(_03209_),
    .A1(net3140),
    .A2(\u_toplayer.reg_layer2[99] ));
 sg13g2_a22oi_1 _09295_ (.Y(_03210_),
    .B1(net2973),
    .B2(\u_toplayer.reg_layer2[115] ),
    .A2(net3006),
    .A1(\u_toplayer.reg_layer2[123] ));
 sg13g2_nand3_1 _09296_ (.B(_03209_),
    .C(_03210_),
    .A(net3103),
    .Y(_03211_));
 sg13g2_nand3_1 _09297_ (.B(_03207_),
    .C(_03211_),
    .A(net3100),
    .Y(_03212_));
 sg13g2_nand2b_1 _09298_ (.Y(_03213_),
    .B(net3134),
    .A_N(\u_toplayer.reg_layer2[43] ));
 sg13g2_o21ai_1 _09299_ (.B1(_03213_),
    .Y(_03214_),
    .A1(net3134),
    .A2(\u_toplayer.reg_layer2[35] ));
 sg13g2_a22oi_1 _09300_ (.Y(_03215_),
    .B1(net2971),
    .B2(\u_toplayer.reg_layer2[51] ),
    .A2(net3004),
    .A1(\u_toplayer.reg_layer2[59] ));
 sg13g2_o21ai_1 _09301_ (.B1(_03215_),
    .Y(_03216_),
    .A1(net3109),
    .A2(_03214_));
 sg13g2_nand2b_1 _09302_ (.Y(_03217_),
    .B(net3121),
    .A_N(\u_toplayer.reg_layer2[11] ));
 sg13g2_o21ai_1 _09303_ (.B1(_03217_),
    .Y(_03218_),
    .A1(net3121),
    .A2(\u_toplayer.reg_layer2[3] ));
 sg13g2_a22oi_1 _09304_ (.Y(_03219_),
    .B1(net2965),
    .B2(\u_toplayer.reg_layer2[19] ),
    .A2(net2998),
    .A1(\u_toplayer.reg_layer2[27] ));
 sg13g2_o21ai_1 _09305_ (.B1(_03219_),
    .Y(_03220_),
    .A1(net3109),
    .A2(_03218_));
 sg13g2_a221oi_1 _09306_ (.B2(net3009),
    .C1(net3096),
    .B1(_03220_),
    .A1(net2935),
    .Y(_03221_),
    .A2(_03216_));
 sg13g2_a21oi_1 _09307_ (.A1(_03212_),
    .A2(_03221_),
    .Y(_03222_),
    .B1(_03070_));
 sg13g2_a22oi_1 _09308_ (.Y(_03223_),
    .B1(_03203_),
    .B2(_03222_),
    .A2(net2817),
    .A1(net3173));
 sg13g2_inv_1 _09309_ (.Y(_00327_),
    .A(_03223_));
 sg13g2_a21oi_1 _09310_ (.A1(net3138),
    .A2(_01083_),
    .Y(_03224_),
    .B1(net3115));
 sg13g2_o21ai_1 _09311_ (.B1(_03224_),
    .Y(_03225_),
    .A1(net3138),
    .A2(\u_toplayer.reg_layer2[100] ));
 sg13g2_a22oi_1 _09312_ (.Y(_03226_),
    .B1(net2974),
    .B2(\u_toplayer.reg_layer2[116] ),
    .A2(net3006),
    .A1(\u_toplayer.reg_layer2[124] ));
 sg13g2_nand3_1 _09313_ (.B(_03225_),
    .C(_03226_),
    .A(net3104),
    .Y(_03227_));
 sg13g2_a21oi_1 _09314_ (.A1(net3123),
    .A2(_01082_),
    .Y(_03228_),
    .B1(net3111));
 sg13g2_o21ai_1 _09315_ (.B1(_03228_),
    .Y(_03229_),
    .A1(net3123),
    .A2(\u_toplayer.reg_layer2[68] ));
 sg13g2_a22oi_1 _09316_ (.Y(_03230_),
    .B1(net2969),
    .B2(\u_toplayer.reg_layer2[84] ),
    .A2(net3002),
    .A1(\u_toplayer.reg_layer2[92] ));
 sg13g2_nand3_1 _09317_ (.B(_03229_),
    .C(_03230_),
    .A(net3017),
    .Y(_03231_));
 sg13g2_nand3_1 _09318_ (.B(_03227_),
    .C(_03231_),
    .A(net3099),
    .Y(_03232_));
 sg13g2_nand2b_1 _09319_ (.Y(_03233_),
    .B(net3132),
    .A_N(\u_toplayer.reg_layer2[44] ));
 sg13g2_o21ai_1 _09320_ (.B1(_03233_),
    .Y(_03234_),
    .A1(net3132),
    .A2(\u_toplayer.reg_layer2[36] ));
 sg13g2_a22oi_1 _09321_ (.Y(_03235_),
    .B1(net2971),
    .B2(\u_toplayer.reg_layer2[52] ),
    .A2(net3004),
    .A1(\u_toplayer.reg_layer2[60] ));
 sg13g2_o21ai_1 _09322_ (.B1(_03235_),
    .Y(_03236_),
    .A1(net3108),
    .A2(_03234_));
 sg13g2_nor2b_1 _09323_ (.A(net3121),
    .B_N(\u_toplayer.reg_layer2[4] ),
    .Y(_03237_));
 sg13g2_a21oi_1 _09324_ (.A1(net3121),
    .A2(\u_toplayer.reg_layer2[12] ),
    .Y(_03238_),
    .B1(_03237_));
 sg13g2_a22oi_1 _09325_ (.Y(_03239_),
    .B1(net2965),
    .B2(\u_toplayer.reg_layer2[20] ),
    .A2(net2998),
    .A1(\u_toplayer.reg_layer2[28] ));
 sg13g2_o21ai_1 _09326_ (.B1(_03239_),
    .Y(_03240_),
    .A1(net3109),
    .A2(_03238_));
 sg13g2_a221oi_1 _09327_ (.B2(net3010),
    .C1(net3097),
    .B1(_03240_),
    .A1(net2937),
    .Y(_03241_),
    .A2(_03236_));
 sg13g2_a21oi_1 _09328_ (.A1(net3122),
    .A2(_01084_),
    .Y(_03242_),
    .B1(net3109));
 sg13g2_o21ai_1 _09329_ (.B1(_03242_),
    .Y(_03243_),
    .A1(net3122),
    .A2(\u_toplayer.reg_layer2[196] ));
 sg13g2_a221oi_1 _09330_ (.B2(\u_toplayer.reg_layer2[212] ),
    .C1(net3102),
    .B1(net2969),
    .A1(\u_toplayer.reg_layer2[220] ),
    .Y(_03244_),
    .A2(net3002));
 sg13g2_mux4_1 _09331_ (.S0(net3134),
    .A0(\u_toplayer.reg_layer2[228] ),
    .A1(\u_toplayer.reg_layer2[236] ),
    .A2(\u_toplayer.reg_layer2[244] ),
    .A3(\u_toplayer.reg_layer2[252] ),
    .S1(net3115),
    .X(_03245_));
 sg13g2_o21ai_1 _09332_ (.B1(net3099),
    .Y(_03246_),
    .A1(net3017),
    .A2(_03245_));
 sg13g2_a21oi_1 _09333_ (.A1(_03243_),
    .A2(_03244_),
    .Y(_03247_),
    .B1(_03246_));
 sg13g2_nand2b_1 _09334_ (.Y(_03248_),
    .B(net3118),
    .A_N(\u_toplayer.reg_layer2[140] ));
 sg13g2_o21ai_1 _09335_ (.B1(_03248_),
    .Y(_03249_),
    .A1(net3119),
    .A2(\u_toplayer.reg_layer2[132] ));
 sg13g2_a22oi_1 _09336_ (.Y(_03250_),
    .B1(net2970),
    .B2(\u_toplayer.reg_layer2[148] ),
    .A2(net2998),
    .A1(\u_toplayer.reg_layer2[156] ));
 sg13g2_o21ai_1 _09337_ (.B1(_03250_),
    .Y(_03251_),
    .A1(net3107),
    .A2(_03249_));
 sg13g2_nor2b_1 _09338_ (.A(net3133),
    .B_N(\u_toplayer.reg_layer2[164] ),
    .Y(_03252_));
 sg13g2_a21oi_1 _09339_ (.A1(net3133),
    .A2(\u_toplayer.reg_layer2[172] ),
    .Y(_03253_),
    .B1(_03252_));
 sg13g2_a22oi_1 _09340_ (.Y(_03254_),
    .B1(net2971),
    .B2(\u_toplayer.reg_layer2[180] ),
    .A2(net3004),
    .A1(\u_toplayer.reg_layer2[188] ));
 sg13g2_o21ai_1 _09341_ (.B1(_03254_),
    .Y(_03255_),
    .A1(net3108),
    .A2(_03253_));
 sg13g2_a221oi_1 _09342_ (.B2(net2937),
    .C1(_03247_),
    .B1(_03255_),
    .A1(net3010),
    .Y(_03256_),
    .A2(_03251_));
 sg13g2_a221oi_1 _09343_ (.B2(net3097),
    .C1(_03070_),
    .B1(_03256_),
    .A1(_03232_),
    .Y(_03257_),
    .A2(_03241_));
 sg13g2_a21o_1 _09344_ (.A2(net2817),
    .A1(net3170),
    .B1(_03257_),
    .X(_00328_));
 sg13g2_a21oi_1 _09345_ (.A1(net3124),
    .A2(_01087_),
    .Y(_03258_),
    .B1(net3111));
 sg13g2_o21ai_1 _09346_ (.B1(_03258_),
    .Y(_03259_),
    .A1(net3124),
    .A2(\u_toplayer.reg_layer2[197] ));
 sg13g2_a22oi_1 _09347_ (.Y(_03260_),
    .B1(net2968),
    .B2(\u_toplayer.reg_layer2[213] ),
    .A2(net3001),
    .A1(\u_toplayer.reg_layer2[221] ));
 sg13g2_nand3_1 _09348_ (.B(_03259_),
    .C(_03260_),
    .A(net3018),
    .Y(_03261_));
 sg13g2_a21oi_1 _09349_ (.A1(net3139),
    .A2(_01088_),
    .Y(_03262_),
    .B1(net3113));
 sg13g2_o21ai_1 _09350_ (.B1(_03262_),
    .Y(_03263_),
    .A1(net3139),
    .A2(\u_toplayer.reg_layer2[229] ));
 sg13g2_a22oi_1 _09351_ (.Y(_03264_),
    .B1(net2972),
    .B2(\u_toplayer.reg_layer2[245] ),
    .A2(net3005),
    .A1(\u_toplayer.reg_layer2[253] ));
 sg13g2_nand3_1 _09352_ (.B(_03263_),
    .C(_03264_),
    .A(net3103),
    .Y(_03265_));
 sg13g2_nand3_1 _09353_ (.B(_03261_),
    .C(_03265_),
    .A(net3099),
    .Y(_03266_));
 sg13g2_nor2b_1 _09354_ (.A(net3130),
    .B_N(\u_toplayer.reg_layer2[165] ),
    .Y(_03267_));
 sg13g2_a21oi_1 _09355_ (.A1(net3130),
    .A2(\u_toplayer.reg_layer2[173] ),
    .Y(_03268_),
    .B1(_03267_));
 sg13g2_a22oi_1 _09356_ (.Y(_03269_),
    .B1(net2967),
    .B2(\u_toplayer.reg_layer2[181] ),
    .A2(net3000),
    .A1(\u_toplayer.reg_layer2[189] ));
 sg13g2_o21ai_1 _09357_ (.B1(_03269_),
    .Y(_03270_),
    .A1(net3106),
    .A2(_03268_));
 sg13g2_nand2b_1 _09358_ (.Y(_03271_),
    .B(net3118),
    .A_N(\u_toplayer.reg_layer2[141] ));
 sg13g2_o21ai_1 _09359_ (.B1(_03271_),
    .Y(_03272_),
    .A1(net3118),
    .A2(\u_toplayer.reg_layer2[133] ));
 sg13g2_a22oi_1 _09360_ (.Y(_03273_),
    .B1(net2965),
    .B2(\u_toplayer.reg_layer2[149] ),
    .A2(net2998),
    .A1(\u_toplayer.reg_layer2[157] ));
 sg13g2_o21ai_1 _09361_ (.B1(_03273_),
    .Y(_03274_),
    .A1(net3107),
    .A2(_03272_));
 sg13g2_a22oi_1 _09362_ (.Y(_03275_),
    .B1(_03274_),
    .B2(net3008),
    .A2(_03270_),
    .A1(net2935));
 sg13g2_nand3_1 _09363_ (.B(_03266_),
    .C(_03275_),
    .A(net3098),
    .Y(_03276_));
 sg13g2_a21oi_1 _09364_ (.A1(net3139),
    .A2(_01086_),
    .Y(_03277_),
    .B1(net3113));
 sg13g2_o21ai_1 _09365_ (.B1(_03277_),
    .Y(_03278_),
    .A1(net3139),
    .A2(\u_toplayer.reg_layer2[101] ));
 sg13g2_a22oi_1 _09366_ (.Y(_03279_),
    .B1(net2972),
    .B2(\u_toplayer.reg_layer2[117] ),
    .A2(net3005),
    .A1(\u_toplayer.reg_layer2[125] ));
 sg13g2_nand3_1 _09367_ (.B(_03278_),
    .C(_03279_),
    .A(net3103),
    .Y(_03280_));
 sg13g2_a21oi_1 _09368_ (.A1(net3125),
    .A2(_01085_),
    .Y(_03281_),
    .B1(net3111));
 sg13g2_o21ai_1 _09369_ (.B1(_03281_),
    .Y(_03282_),
    .A1(net3124),
    .A2(\u_toplayer.reg_layer2[69] ));
 sg13g2_a22oi_1 _09370_ (.Y(_03283_),
    .B1(net2968),
    .B2(\u_toplayer.reg_layer2[85] ),
    .A2(net3001),
    .A1(\u_toplayer.reg_layer2[93] ));
 sg13g2_nand3_1 _09371_ (.B(_03282_),
    .C(_03283_),
    .A(net3018),
    .Y(_03284_));
 sg13g2_nand3_1 _09372_ (.B(_03280_),
    .C(_03284_),
    .A(net3099),
    .Y(_03285_));
 sg13g2_nand2b_1 _09373_ (.Y(_03286_),
    .B(net3119),
    .A_N(\u_toplayer.reg_layer2[13] ));
 sg13g2_o21ai_1 _09374_ (.B1(_03286_),
    .Y(_03287_),
    .A1(net3119),
    .A2(\u_toplayer.reg_layer2[5] ));
 sg13g2_a22oi_1 _09375_ (.Y(_03288_),
    .B1(net2965),
    .B2(\u_toplayer.reg_layer2[21] ),
    .A2(net2998),
    .A1(\u_toplayer.reg_layer2[29] ));
 sg13g2_o21ai_1 _09376_ (.B1(_03288_),
    .Y(_03289_),
    .A1(net3107),
    .A2(_03287_));
 sg13g2_nand2b_1 _09377_ (.Y(_03290_),
    .B(net3130),
    .A_N(\u_toplayer.reg_layer2[45] ));
 sg13g2_o21ai_1 _09378_ (.B1(_03290_),
    .Y(_03291_),
    .A1(net3130),
    .A2(\u_toplayer.reg_layer2[37] ));
 sg13g2_a22oi_1 _09379_ (.Y(_03292_),
    .B1(net2967),
    .B2(\u_toplayer.reg_layer2[53] ),
    .A2(net3000),
    .A1(\u_toplayer.reg_layer2[61] ));
 sg13g2_o21ai_1 _09380_ (.B1(_03292_),
    .Y(_03293_),
    .A1(net3106),
    .A2(_03291_));
 sg13g2_a221oi_1 _09381_ (.B2(net2935),
    .C1(net3096),
    .B1(_03293_),
    .A1(net3008),
    .Y(_03294_),
    .A2(_03289_));
 sg13g2_a21oi_1 _09382_ (.A1(_03285_),
    .A2(_03294_),
    .Y(_03295_),
    .B1(_03070_));
 sg13g2_a22oi_1 _09383_ (.Y(_03296_),
    .B1(_03276_),
    .B2(_03295_),
    .A2(net2817),
    .A1(net1023));
 sg13g2_inv_1 _09384_ (.Y(_00329_),
    .A(_03296_));
 sg13g2_nor2b_1 _09385_ (.A(\u_toplayer.reg_layer2[238] ),
    .B_N(net3138),
    .Y(_03297_));
 sg13g2_nor2_1 _09386_ (.A(net3138),
    .B(\u_toplayer.reg_layer2[230] ),
    .Y(_03298_));
 sg13g2_nor3_1 _09387_ (.A(net3113),
    .B(_03297_),
    .C(_03298_),
    .Y(_03299_));
 sg13g2_a221oi_1 _09388_ (.B2(\u_toplayer.reg_layer2[246] ),
    .C1(_03299_),
    .B1(net2973),
    .A1(\u_toplayer.reg_layer2[254] ),
    .Y(_03300_),
    .A2(net3006));
 sg13g2_a21oi_1 _09389_ (.A1(net3123),
    .A2(_01091_),
    .Y(_03301_),
    .B1(net3111));
 sg13g2_o21ai_1 _09390_ (.B1(_03301_),
    .Y(_03302_),
    .A1(net3123),
    .A2(\u_toplayer.reg_layer2[198] ));
 sg13g2_a221oi_1 _09391_ (.B2(\u_toplayer.reg_layer2[214] ),
    .C1(net3102),
    .B1(net2969),
    .A1(\u_toplayer.reg_layer2[222] ),
    .Y(_03303_),
    .A2(net3002));
 sg13g2_a22oi_1 _09392_ (.Y(_03304_),
    .B1(_03302_),
    .B2(_03303_),
    .A2(_03300_),
    .A1(net3102));
 sg13g2_nand2_1 _09393_ (.Y(_03305_),
    .A(net3099),
    .B(_03304_));
 sg13g2_nand2b_1 _09394_ (.Y(_03306_),
    .B(net3129),
    .A_N(\u_toplayer.reg_layer2[174] ));
 sg13g2_o21ai_1 _09395_ (.B1(_03306_),
    .Y(_03307_),
    .A1(net3131),
    .A2(\u_toplayer.reg_layer2[166] ));
 sg13g2_a22oi_1 _09396_ (.Y(_03308_),
    .B1(net2967),
    .B2(\u_toplayer.reg_layer2[182] ),
    .A2(net3000),
    .A1(\u_toplayer.reg_layer2[190] ));
 sg13g2_o21ai_1 _09397_ (.B1(_03308_),
    .Y(_03309_),
    .A1(net3106),
    .A2(_03307_));
 sg13g2_nand2b_1 _09398_ (.Y(_03310_),
    .B(net3117),
    .A_N(\u_toplayer.reg_layer2[142] ));
 sg13g2_o21ai_1 _09399_ (.B1(_03310_),
    .Y(_03311_),
    .A1(net3117),
    .A2(\u_toplayer.reg_layer2[134] ));
 sg13g2_a22oi_1 _09400_ (.Y(_03312_),
    .B1(net2966),
    .B2(\u_toplayer.reg_layer2[150] ),
    .A2(net2999),
    .A1(\u_toplayer.reg_layer2[158] ));
 sg13g2_o21ai_1 _09401_ (.B1(_03312_),
    .Y(_03313_),
    .A1(net3106),
    .A2(_03311_));
 sg13g2_a22oi_1 _09402_ (.Y(_03314_),
    .B1(_03313_),
    .B2(net3008),
    .A2(_03309_),
    .A1(net2935));
 sg13g2_nand3_1 _09403_ (.B(_03305_),
    .C(_03314_),
    .A(net3097),
    .Y(_03315_));
 sg13g2_a21oi_1 _09404_ (.A1(net3123),
    .A2(_01089_),
    .Y(_03316_),
    .B1(net3111));
 sg13g2_o21ai_1 _09405_ (.B1(_03316_),
    .Y(_03317_),
    .A1(net3123),
    .A2(\u_toplayer.reg_layer2[70] ));
 sg13g2_a22oi_1 _09406_ (.Y(_03318_),
    .B1(net2969),
    .B2(\u_toplayer.reg_layer2[86] ),
    .A2(net3002),
    .A1(\u_toplayer.reg_layer2[94] ));
 sg13g2_nand3_1 _09407_ (.B(_03317_),
    .C(_03318_),
    .A(net3018),
    .Y(_03319_));
 sg13g2_a21oi_1 _09408_ (.A1(net3138),
    .A2(_01090_),
    .Y(_03320_),
    .B1(net3113));
 sg13g2_o21ai_1 _09409_ (.B1(_03320_),
    .Y(_03321_),
    .A1(net3138),
    .A2(\u_toplayer.reg_layer2[102] ));
 sg13g2_a22oi_1 _09410_ (.Y(_03322_),
    .B1(net2974),
    .B2(\u_toplayer.reg_layer2[118] ),
    .A2(net3007),
    .A1(\u_toplayer.reg_layer2[126] ));
 sg13g2_nand3_1 _09411_ (.B(_03321_),
    .C(_03322_),
    .A(net3104),
    .Y(_03323_));
 sg13g2_nand3_1 _09412_ (.B(_03319_),
    .C(_03323_),
    .A(net3099),
    .Y(_03324_));
 sg13g2_nor2b_1 _09413_ (.A(net3131),
    .B_N(\u_toplayer.reg_layer2[38] ),
    .Y(_03325_));
 sg13g2_a21oi_2 _09414_ (.B1(_03325_),
    .Y(_03326_),
    .A2(\u_toplayer.reg_layer2[46] ),
    .A1(net3129));
 sg13g2_a22oi_1 _09415_ (.Y(_03327_),
    .B1(net2967),
    .B2(\u_toplayer.reg_layer2[54] ),
    .A2(net3000),
    .A1(\u_toplayer.reg_layer2[62] ));
 sg13g2_o21ai_1 _09416_ (.B1(_03327_),
    .Y(_03328_),
    .A1(net3106),
    .A2(_03326_));
 sg13g2_nand2b_1 _09417_ (.Y(_03329_),
    .B(net3117),
    .A_N(\u_toplayer.reg_layer2[14] ));
 sg13g2_o21ai_1 _09418_ (.B1(_03329_),
    .Y(_03330_),
    .A1(net3117),
    .A2(\u_toplayer.reg_layer2[6] ));
 sg13g2_a22oi_1 _09419_ (.Y(_03331_),
    .B1(net2966),
    .B2(\u_toplayer.reg_layer2[22] ),
    .A2(net2999),
    .A1(\u_toplayer.reg_layer2[30] ));
 sg13g2_o21ai_1 _09420_ (.B1(_03331_),
    .Y(_03332_),
    .A1(net3107),
    .A2(_03330_));
 sg13g2_a221oi_1 _09421_ (.B2(net3008),
    .C1(net3096),
    .B1(_03332_),
    .A1(net2935),
    .Y(_03333_),
    .A2(_03328_));
 sg13g2_a21oi_1 _09422_ (.A1(_03324_),
    .A2(_03333_),
    .Y(_03334_),
    .B1(_03070_));
 sg13g2_a22oi_1 _09423_ (.Y(_03335_),
    .B1(_03315_),
    .B2(_03334_),
    .A2(net2817),
    .A1(net1113));
 sg13g2_inv_1 _09424_ (.Y(_00330_),
    .A(_03335_));
 sg13g2_nor2b_1 _09425_ (.A(\u_toplayer.reg_layer2[239] ),
    .B_N(net3134),
    .Y(_03336_));
 sg13g2_nor2_1 _09426_ (.A(net3134),
    .B(\u_toplayer.reg_layer2[231] ),
    .Y(_03337_));
 sg13g2_nor3_1 _09427_ (.A(net3115),
    .B(_03336_),
    .C(_03337_),
    .Y(_03338_));
 sg13g2_a221oi_1 _09428_ (.B2(\u_toplayer.reg_layer2[247] ),
    .C1(_03338_),
    .B1(net2972),
    .A1(\u_toplayer.reg_layer2[255] ),
    .Y(_03339_),
    .A2(net3006));
 sg13g2_a21oi_1 _09429_ (.A1(net3122),
    .A2(_01094_),
    .Y(_03340_),
    .B1(net3109));
 sg13g2_o21ai_1 _09430_ (.B1(_03340_),
    .Y(_03341_),
    .A1(net3121),
    .A2(\u_toplayer.reg_layer2[199] ));
 sg13g2_a221oi_1 _09431_ (.B2(\u_toplayer.reg_layer2[215] ),
    .C1(net3102),
    .B1(net2969),
    .A1(\u_toplayer.reg_layer2[223] ),
    .Y(_03342_),
    .A2(net3002));
 sg13g2_a22oi_1 _09432_ (.Y(_03343_),
    .B1(_03341_),
    .B2(_03342_),
    .A2(_03339_),
    .A1(net3105));
 sg13g2_nand2_1 _09433_ (.Y(_03344_),
    .A(net3099),
    .B(_03343_));
 sg13g2_nor2b_1 _09434_ (.A(net3129),
    .B_N(\u_toplayer.reg_layer2[167] ),
    .Y(_03345_));
 sg13g2_a21oi_1 _09435_ (.A1(net3129),
    .A2(\u_toplayer.reg_layer2[175] ),
    .Y(_03346_),
    .B1(_03345_));
 sg13g2_a22oi_1 _09436_ (.Y(_03347_),
    .B1(net2967),
    .B2(\u_toplayer.reg_layer2[183] ),
    .A2(net3000),
    .A1(\u_toplayer.reg_layer2[191] ));
 sg13g2_o21ai_1 _09437_ (.B1(_03347_),
    .Y(_03348_),
    .A1(net3106),
    .A2(_03346_));
 sg13g2_nand2b_1 _09438_ (.Y(_03349_),
    .B(net3117),
    .A_N(\u_toplayer.reg_layer2[143] ));
 sg13g2_o21ai_1 _09439_ (.B1(_03349_),
    .Y(_03350_),
    .A1(net3117),
    .A2(\u_toplayer.reg_layer2[135] ));
 sg13g2_a22oi_1 _09440_ (.Y(_03351_),
    .B1(net2966),
    .B2(\u_toplayer.reg_layer2[151] ),
    .A2(net2999),
    .A1(\u_toplayer.reg_layer2[159] ));
 sg13g2_o21ai_1 _09441_ (.B1(_03351_),
    .Y(_03352_),
    .A1(net3106),
    .A2(_03350_));
 sg13g2_a22oi_1 _09442_ (.Y(_03353_),
    .B1(_03352_),
    .B2(net3008),
    .A2(_03348_),
    .A1(net2935));
 sg13g2_nand3_1 _09443_ (.B(_03344_),
    .C(_03353_),
    .A(net3097),
    .Y(_03354_));
 sg13g2_a21oi_1 _09444_ (.A1(net3123),
    .A2(_01092_),
    .Y(_03355_),
    .B1(net3111));
 sg13g2_o21ai_1 _09445_ (.B1(_03355_),
    .Y(_03356_),
    .A1(net3123),
    .A2(\u_toplayer.reg_layer2[71] ));
 sg13g2_a22oi_1 _09446_ (.Y(_03357_),
    .B1(net2969),
    .B2(\u_toplayer.reg_layer2[87] ),
    .A2(net3002),
    .A1(\u_toplayer.reg_layer2[95] ));
 sg13g2_nand3_1 _09447_ (.B(_03356_),
    .C(_03357_),
    .A(net3017),
    .Y(_03358_));
 sg13g2_a21oi_1 _09448_ (.A1(net3138),
    .A2(_01093_),
    .Y(_03359_),
    .B1(net3113));
 sg13g2_o21ai_1 _09449_ (.B1(_03359_),
    .Y(_03360_),
    .A1(net3138),
    .A2(\u_toplayer.reg_layer2[103] ));
 sg13g2_a22oi_1 _09450_ (.Y(_03361_),
    .B1(net2972),
    .B2(\u_toplayer.reg_layer2[119] ),
    .A2(net3005),
    .A1(\u_toplayer.reg_layer2[127] ));
 sg13g2_nand3_1 _09451_ (.B(_03360_),
    .C(_03361_),
    .A(net3104),
    .Y(_03362_));
 sg13g2_nand3_1 _09452_ (.B(_03358_),
    .C(_03362_),
    .A(net3101),
    .Y(_03363_));
 sg13g2_nand2b_1 _09453_ (.Y(_03364_),
    .B(net3129),
    .A_N(\u_toplayer.reg_layer2[47] ));
 sg13g2_o21ai_1 _09454_ (.B1(_03364_),
    .Y(_03365_),
    .A1(net3129),
    .A2(\u_toplayer.reg_layer2[39] ));
 sg13g2_a22oi_1 _09455_ (.Y(_03366_),
    .B1(net2967),
    .B2(\u_toplayer.reg_layer2[55] ),
    .A2(net3000),
    .A1(\u_toplayer.reg_layer2[63] ));
 sg13g2_o21ai_1 _09456_ (.B1(_03366_),
    .Y(_03367_),
    .A1(net3108),
    .A2(_03365_));
 sg13g2_nor2b_1 _09457_ (.A(net3120),
    .B_N(\u_toplayer.reg_layer2[7] ),
    .Y(_03368_));
 sg13g2_a21oi_1 _09458_ (.A1(net3117),
    .A2(\u_toplayer.reg_layer2[15] ),
    .Y(_03369_),
    .B1(_03368_));
 sg13g2_a22oi_1 _09459_ (.Y(_03370_),
    .B1(net2966),
    .B2(\u_toplayer.reg_layer2[23] ),
    .A2(net2999),
    .A1(\u_toplayer.reg_layer2[31] ));
 sg13g2_o21ai_1 _09460_ (.B1(_03370_),
    .Y(_03371_),
    .A1(net3107),
    .A2(_03369_));
 sg13g2_a221oi_1 _09461_ (.B2(net3009),
    .C1(net3096),
    .B1(_03371_),
    .A1(net2936),
    .Y(_03372_),
    .A2(_03367_));
 sg13g2_a21oi_1 _09462_ (.A1(_03363_),
    .A2(_03372_),
    .Y(_03373_),
    .B1(_03070_));
 sg13g2_a22oi_1 _09463_ (.Y(_03374_),
    .B1(_03354_),
    .B2(_03373_),
    .A2(net2817),
    .A1(net3162));
 sg13g2_inv_1 _09464_ (.Y(_00331_),
    .A(_03374_));
 sg13g2_or2_2 _09465_ (.X(_03375_),
    .B(_01940_),
    .A(_01937_));
 sg13g2_nand2_1 _09466_ (.Y(_03376_),
    .A(net1085),
    .B(_03375_));
 sg13g2_nor4_2 _09467_ (.A(\u_toplayer.u_layer3.u_neuron.acc[13] ),
    .B(\u_toplayer.u_layer3.u_neuron.acc[10] ),
    .C(\u_toplayer.u_layer3.u_neuron.acc[11] ),
    .Y(_03377_),
    .D(\u_toplayer.u_layer3.u_neuron.acc[9] ));
 sg13g2_nor4_1 _09468_ (.A(\u_toplayer.u_layer3.u_neuron.acc[7] ),
    .B(net3157),
    .C(\u_toplayer.u_layer3.u_neuron.acc[15] ),
    .D(\u_toplayer.u_layer3.u_neuron.acc[12] ),
    .Y(_03378_));
 sg13g2_nor4_1 _09469_ (.A(net3158),
    .B(\u_toplayer.u_layer3.u_neuron.acc[22] ),
    .C(\u_toplayer.u_layer3.u_neuron.acc[21] ),
    .D(net3154),
    .Y(_03379_));
 sg13g2_nor4_1 _09470_ (.A(\u_toplayer.u_layer3.u_neuron.acc[19] ),
    .B(net3155),
    .C(net3156),
    .D(\u_toplayer.u_layer3.u_neuron.acc[17] ),
    .Y(_03380_));
 sg13g2_and3_1 _09471_ (.X(_03381_),
    .A(_03377_),
    .B(_03378_),
    .C(_03380_));
 sg13g2_a21oi_2 _09472_ (.B1(net1068),
    .Y(_03382_),
    .A2(_03381_),
    .A1(_03379_));
 sg13g2_nor2_1 _09473_ (.A(net1047),
    .B(_03382_),
    .Y(_03383_));
 sg13g2_nand4_1 _09474_ (.B(\u_toplayer.u_layer3.u_neuron.acc[10] ),
    .C(\u_toplayer.u_layer3.u_neuron.acc[11] ),
    .A(\u_toplayer.u_layer3.u_neuron.acc[13] ),
    .Y(_03384_),
    .D(\u_toplayer.u_layer3.u_neuron.acc[9] ));
 sg13g2_nand4_1 _09475_ (.B(net3157),
    .C(\u_toplayer.u_layer3.u_neuron.acc[15] ),
    .A(\u_toplayer.u_layer3.u_neuron.acc[7] ),
    .Y(_03385_),
    .D(\u_toplayer.u_layer3.u_neuron.acc[12] ));
 sg13g2_nand4_1 _09476_ (.B(\u_toplayer.u_layer3.u_neuron.acc[22] ),
    .C(\u_toplayer.u_layer3.u_neuron.acc[21] ),
    .A(net3158),
    .Y(_03386_),
    .D(net3154));
 sg13g2_nand4_1 _09477_ (.B(net3155),
    .C(net3156),
    .A(\u_toplayer.u_layer3.u_neuron.acc[19] ),
    .Y(_03387_),
    .D(\u_toplayer.u_layer3.u_neuron.acc[17] ));
 sg13g2_nor3_1 _09478_ (.A(_01050_),
    .B(\u_toplayer.u_layer3.u_neuron.acc[6] ),
    .C(net3159),
    .Y(_03388_));
 sg13g2_nor4_1 _09479_ (.A(\u_toplayer.u_layer3.u_neuron.acc[3] ),
    .B(\u_toplayer.u_layer3.u_neuron.acc[2] ),
    .C(\u_toplayer.u_layer3.u_neuron.acc[1] ),
    .D(\u_toplayer.u_layer3.u_neuron.acc[0] ),
    .Y(_03389_));
 sg13g2_nand3_1 _09480_ (.B(_03388_),
    .C(_03389_),
    .A(_01052_),
    .Y(_03390_));
 sg13g2_nor4_1 _09481_ (.A(_03384_),
    .B(_03385_),
    .C(_03386_),
    .D(_03387_),
    .Y(_03391_));
 sg13g2_a21oi_1 _09482_ (.A1(_03390_),
    .A2(_03391_),
    .Y(_03392_),
    .B1(_01061_));
 sg13g2_or2_2 _09483_ (.X(_03393_),
    .B(_03392_),
    .A(net2816));
 sg13g2_o21ai_1 _09484_ (.B1(_03376_),
    .Y(_00332_),
    .A1(_03383_),
    .A2(_03393_));
 sg13g2_nand2_1 _09485_ (.Y(_03394_),
    .A(net1026),
    .B(net2816));
 sg13g2_nor2_1 _09486_ (.A(\u_toplayer.u_layer3.u_neuron.acc[1] ),
    .B(_03382_),
    .Y(_03395_));
 sg13g2_o21ai_1 _09487_ (.B1(_03394_),
    .Y(_00333_),
    .A1(_03393_),
    .A2(_03395_));
 sg13g2_nand2_1 _09488_ (.Y(_03396_),
    .A(net1053),
    .B(net2816));
 sg13g2_nor2_1 _09489_ (.A(\u_toplayer.u_layer3.u_neuron.acc[2] ),
    .B(_03382_),
    .Y(_03397_));
 sg13g2_o21ai_1 _09490_ (.B1(_03396_),
    .Y(_00334_),
    .A1(_03393_),
    .A2(_03397_));
 sg13g2_nand2_1 _09491_ (.Y(_03398_),
    .A(net1076),
    .B(net2816));
 sg13g2_nor2_1 _09492_ (.A(\u_toplayer.u_layer3.u_neuron.acc[3] ),
    .B(_03382_),
    .Y(_03399_));
 sg13g2_o21ai_1 _09493_ (.B1(_03398_),
    .Y(_00335_),
    .A1(_03393_),
    .A2(_03399_));
 sg13g2_nand2_1 _09494_ (.Y(_03400_),
    .A(net1030),
    .B(net2816));
 sg13g2_nor2_1 _09495_ (.A(\u_toplayer.u_layer3.u_neuron.acc[4] ),
    .B(_03382_),
    .Y(_03401_));
 sg13g2_o21ai_1 _09496_ (.B1(_03400_),
    .Y(_00336_),
    .A1(_03393_),
    .A2(_03401_));
 sg13g2_nand2_1 _09497_ (.Y(_03402_),
    .A(net1101),
    .B(net2816));
 sg13g2_nor2_1 _09498_ (.A(net3159),
    .B(_03382_),
    .Y(_03403_));
 sg13g2_o21ai_1 _09499_ (.B1(_03402_),
    .Y(_00337_),
    .A1(_03393_),
    .A2(_03403_));
 sg13g2_nand2_1 _09500_ (.Y(_03404_),
    .A(net1044),
    .B(net2816));
 sg13g2_nor2_1 _09501_ (.A(\u_toplayer.u_layer3.u_neuron.acc[6] ),
    .B(_03382_),
    .Y(_03405_));
 sg13g2_o21ai_1 _09502_ (.B1(_03404_),
    .Y(_00338_),
    .A1(_03393_),
    .A2(_03405_));
 sg13g2_mux2_1 _09503_ (.A0(net1032),
    .A1(\u_toplayer.u_layer3.sum[7] ),
    .S(net2816),
    .X(_00339_));
 sg13g2_nand2_1 _09504_ (.Y(_03406_),
    .A(\u_toplayer.u_layer3.u_neuron.acc[0] ),
    .B(\u_toplayer.u_layer3.u_neuron.mult[0] ));
 sg13g2_xor2_1 _09505_ (.B(net927),
    .A(\u_toplayer.u_layer3.u_neuron.acc[0] ),
    .X(_03407_));
 sg13g2_nand2_1 _09506_ (.Y(_03408_),
    .A(net3404),
    .B(\u_toplayer.u_layer3.u_neuron.acc[0] ));
 sg13g2_xor2_1 _09507_ (.B(\u_toplayer.u_layer3.u_neuron.acc[0] ),
    .A(net3404),
    .X(_03409_));
 sg13g2_a22oi_1 _09508_ (.Y(_03410_),
    .B1(_03409_),
    .B2(net2896),
    .A2(_03407_),
    .A1(net2862));
 sg13g2_nor2_1 _09509_ (.A(net1047),
    .B(net2757),
    .Y(_03411_));
 sg13g2_a21oi_1 _09510_ (.A1(net2757),
    .A2(_03410_),
    .Y(_00349_),
    .B1(_03411_));
 sg13g2_nand2_1 _09511_ (.Y(_03412_),
    .A(net3400),
    .B(\u_toplayer.u_layer3.u_neuron.acc[1] ));
 sg13g2_nor2_1 _09512_ (.A(net3400),
    .B(\u_toplayer.u_layer3.u_neuron.acc[1] ),
    .Y(_03413_));
 sg13g2_xor2_1 _09513_ (.B(\u_toplayer.u_layer3.u_neuron.acc[1] ),
    .A(net3400),
    .X(_03414_));
 sg13g2_xnor2_1 _09514_ (.Y(_03415_),
    .A(_03408_),
    .B(_03414_));
 sg13g2_nand2_1 _09515_ (.Y(_03416_),
    .A(\u_toplayer.u_layer3.u_neuron.acc[1] ),
    .B(\u_toplayer.u_layer3.u_neuron.mult[1] ));
 sg13g2_xnor2_1 _09516_ (.Y(_03417_),
    .A(\u_toplayer.u_layer3.u_neuron.acc[1] ),
    .B(\u_toplayer.u_layer3.u_neuron.mult[1] ));
 sg13g2_xor2_1 _09517_ (.B(_03417_),
    .A(_03406_),
    .X(_03418_));
 sg13g2_a22oi_1 _09518_ (.Y(_03419_),
    .B1(_03418_),
    .B2(net2862),
    .A2(_03415_),
    .A1(net2896));
 sg13g2_nor2_1 _09519_ (.A(net1086),
    .B(net2757),
    .Y(_03420_));
 sg13g2_a21oi_1 _09520_ (.A1(net2757),
    .A2(_03419_),
    .Y(_00350_),
    .B1(_03420_));
 sg13g2_and2_1 _09521_ (.A(net3396),
    .B(\u_toplayer.u_layer3.u_neuron.acc[2] ),
    .X(_03421_));
 sg13g2_xor2_1 _09522_ (.B(\u_toplayer.u_layer3.u_neuron.acc[2] ),
    .A(net3396),
    .X(_03422_));
 sg13g2_o21ai_1 _09523_ (.B1(_03412_),
    .Y(_03423_),
    .A1(_03408_),
    .A2(_03413_));
 sg13g2_nand2_1 _09524_ (.Y(_03424_),
    .A(_03422_),
    .B(_03423_));
 sg13g2_o21ai_1 _09525_ (.B1(net2896),
    .Y(_03425_),
    .A1(_03422_),
    .A2(_03423_));
 sg13g2_inv_1 _09526_ (.Y(_03426_),
    .A(_03425_));
 sg13g2_o21ai_1 _09527_ (.B1(_03416_),
    .Y(_03427_),
    .A1(_03406_),
    .A2(_03417_));
 sg13g2_and2_1 _09528_ (.A(\u_toplayer.u_layer3.u_neuron.acc[2] ),
    .B(\u_toplayer.u_layer3.u_neuron.mult[2] ),
    .X(_03428_));
 sg13g2_xor2_1 _09529_ (.B(\u_toplayer.u_layer3.u_neuron.mult[2] ),
    .A(\u_toplayer.u_layer3.u_neuron.acc[2] ),
    .X(_03429_));
 sg13g2_xor2_1 _09530_ (.B(_03429_),
    .A(_03427_),
    .X(_03430_));
 sg13g2_a22oi_1 _09531_ (.Y(_03431_),
    .B1(_03430_),
    .B2(net2862),
    .A2(_03426_),
    .A1(_03424_));
 sg13g2_nor2_1 _09532_ (.A(net1061),
    .B(net2757),
    .Y(_03432_));
 sg13g2_a21oi_1 _09533_ (.A1(net2757),
    .A2(_03431_),
    .Y(_00351_),
    .B1(_03432_));
 sg13g2_nand2_1 _09534_ (.Y(_03433_),
    .A(net3393),
    .B(\u_toplayer.u_layer3.u_neuron.acc[3] ));
 sg13g2_xnor2_1 _09535_ (.Y(_03434_),
    .A(net3393),
    .B(\u_toplayer.u_layer3.u_neuron.acc[3] ));
 sg13g2_a21oi_1 _09536_ (.A1(_03422_),
    .A2(_03423_),
    .Y(_03435_),
    .B1(_03421_));
 sg13g2_a21oi_1 _09537_ (.A1(_03434_),
    .A2(_03435_),
    .Y(_03436_),
    .B1(net2894));
 sg13g2_o21ai_1 _09538_ (.B1(_03436_),
    .Y(_03437_),
    .A1(_03434_),
    .A2(_03435_));
 sg13g2_nand2_1 _09539_ (.Y(_03438_),
    .A(\u_toplayer.u_layer3.u_neuron.acc[3] ),
    .B(\u_toplayer.u_layer3.u_neuron.mult[3] ));
 sg13g2_xnor2_1 _09540_ (.Y(_03439_),
    .A(\u_toplayer.u_layer3.u_neuron.acc[3] ),
    .B(\u_toplayer.u_layer3.u_neuron.mult[3] ));
 sg13g2_a21oi_1 _09541_ (.A1(_03427_),
    .A2(_03429_),
    .Y(_03440_),
    .B1(_03428_));
 sg13g2_xor2_1 _09542_ (.B(_03440_),
    .A(_03439_),
    .X(_03441_));
 sg13g2_a21oi_1 _09543_ (.A1(net2862),
    .A2(_03441_),
    .Y(_03442_),
    .B1(net2764));
 sg13g2_a22oi_1 _09544_ (.Y(_00352_),
    .B1(_03437_),
    .B2(_03442_),
    .A2(net2761),
    .A1(_01053_));
 sg13g2_and2_1 _09545_ (.A(\u_toplayer.u_layer3.u_neuron.acc[4] ),
    .B(\u_toplayer.u_layer3.u_neuron.mult[4] ),
    .X(_03443_));
 sg13g2_xnor2_1 _09546_ (.Y(_03444_),
    .A(\u_toplayer.u_layer3.u_neuron.acc[4] ),
    .B(\u_toplayer.u_layer3.u_neuron.mult[4] ));
 sg13g2_inv_1 _09547_ (.Y(_03445_),
    .A(_03444_));
 sg13g2_o21ai_1 _09548_ (.B1(_03438_),
    .Y(_03446_),
    .A1(_03439_),
    .A2(_03440_));
 sg13g2_xnor2_1 _09549_ (.Y(_03447_),
    .A(_03444_),
    .B(_03446_));
 sg13g2_nor2_1 _09550_ (.A(_01046_),
    .B(_01052_),
    .Y(_03448_));
 sg13g2_xor2_1 _09551_ (.B(\u_toplayer.u_layer3.u_neuron.acc[4] ),
    .A(net3390),
    .X(_03449_));
 sg13g2_o21ai_1 _09552_ (.B1(_03433_),
    .Y(_03450_),
    .A1(_03434_),
    .A2(_03435_));
 sg13g2_o21ai_1 _09553_ (.B1(net2896),
    .Y(_03451_),
    .A1(_03449_),
    .A2(_03450_));
 sg13g2_a21o_1 _09554_ (.A2(_03450_),
    .A1(_03449_),
    .B1(_03451_),
    .X(_03452_));
 sg13g2_a21oi_1 _09555_ (.A1(net2862),
    .A2(_03447_),
    .Y(_03453_),
    .B1(net2761));
 sg13g2_a22oi_1 _09556_ (.Y(_00353_),
    .B1(_03452_),
    .B2(_03453_),
    .A2(net2760),
    .A1(_01052_));
 sg13g2_nor2_1 _09557_ (.A(\u_toplayer.u_layer3.u_neuron.acc[5] ),
    .B(\u_toplayer.u_layer3.u_neuron.mult[5] ),
    .Y(_03454_));
 sg13g2_xnor2_1 _09558_ (.Y(_03455_),
    .A(net3159),
    .B(\u_toplayer.u_layer3.u_neuron.mult[5] ));
 sg13g2_a21o_1 _09559_ (.A2(_03446_),
    .A1(_03445_),
    .B1(_03443_),
    .X(_03456_));
 sg13g2_xnor2_1 _09560_ (.Y(_03457_),
    .A(_03455_),
    .B(_03456_));
 sg13g2_a21oi_1 _09561_ (.A1(_03449_),
    .A2(_03450_),
    .Y(_03458_),
    .B1(_03448_));
 sg13g2_and2_1 _09562_ (.A(net3386),
    .B(net3159),
    .X(_03459_));
 sg13g2_nor2_1 _09563_ (.A(net3386),
    .B(net3159),
    .Y(_03460_));
 sg13g2_nor3_1 _09564_ (.A(_03458_),
    .B(_03459_),
    .C(_03460_),
    .Y(_03461_));
 sg13g2_o21ai_1 _09565_ (.B1(_03458_),
    .Y(_03462_),
    .A1(_03459_),
    .A2(_03460_));
 sg13g2_nor2_1 _09566_ (.A(net2894),
    .B(_03461_),
    .Y(_03463_));
 sg13g2_a22oi_1 _09567_ (.Y(_03464_),
    .B1(_03462_),
    .B2(_03463_),
    .A2(_03457_),
    .A1(net2862));
 sg13g2_nor2_1 _09568_ (.A(net3159),
    .B(net2757),
    .Y(_03465_));
 sg13g2_a21oi_1 _09569_ (.A1(net2757),
    .A2(_03464_),
    .Y(_00354_),
    .B1(_03465_));
 sg13g2_and2_1 _09570_ (.A(\u_toplayer.u_layer3.u_neuron.acc[6] ),
    .B(\u_toplayer.u_layer3.u_neuron.mult[6] ),
    .X(_03466_));
 sg13g2_xnor2_1 _09571_ (.Y(_03467_),
    .A(\u_toplayer.u_layer3.u_neuron.acc[6] ),
    .B(\u_toplayer.u_layer3.u_neuron.mult[6] ));
 sg13g2_a221oi_1 _09572_ (.B2(_03446_),
    .C1(_03443_),
    .B1(_03445_),
    .A1(net3159),
    .Y(_03468_),
    .A2(\u_toplayer.u_layer3.u_neuron.mult[5] ));
 sg13g2_o21ai_1 _09573_ (.B1(_03467_),
    .Y(_03469_),
    .A1(_03454_),
    .A2(_03468_));
 sg13g2_nor3_2 _09574_ (.A(_03454_),
    .B(_03467_),
    .C(_03468_),
    .Y(_03470_));
 sg13g2_nor2_1 _09575_ (.A(net2865),
    .B(_03470_),
    .Y(_03471_));
 sg13g2_nand2_1 _09576_ (.Y(_03472_),
    .A(net3383),
    .B(\u_toplayer.u_layer3.u_neuron.acc[6] ));
 sg13g2_xnor2_1 _09577_ (.Y(_03473_),
    .A(net3383),
    .B(\u_toplayer.u_layer3.u_neuron.acc[6] ));
 sg13g2_a221oi_1 _09578_ (.B2(_03450_),
    .C1(_03448_),
    .B1(_03449_),
    .A1(net3386),
    .Y(_03474_),
    .A2(net3159));
 sg13g2_or3_1 _09579_ (.A(_03460_),
    .B(_03473_),
    .C(_03474_),
    .X(_03475_));
 sg13g2_o21ai_1 _09580_ (.B1(_03473_),
    .Y(_03476_),
    .A1(_03460_),
    .A2(_03474_));
 sg13g2_nand3_1 _09581_ (.B(_03475_),
    .C(_03476_),
    .A(net2896),
    .Y(_03477_));
 sg13g2_a21oi_1 _09582_ (.A1(_03469_),
    .A2(_03471_),
    .Y(_03478_),
    .B1(net2762));
 sg13g2_a22oi_1 _09583_ (.Y(_00355_),
    .B1(_03477_),
    .B2(_03478_),
    .A2(net2762),
    .A1(_01051_));
 sg13g2_and2_1 _09584_ (.A(net3373),
    .B(\u_toplayer.u_layer3.u_neuron.acc[7] ),
    .X(_03479_));
 sg13g2_xor2_1 _09585_ (.B(\u_toplayer.u_layer3.u_neuron.acc[7] ),
    .A(net3372),
    .X(_03480_));
 sg13g2_inv_1 _09586_ (.Y(_03481_),
    .A(_03480_));
 sg13g2_nand3_1 _09587_ (.B(_03475_),
    .C(_03481_),
    .A(_03472_),
    .Y(_03482_));
 sg13g2_a21oi_2 _09588_ (.B1(_03481_),
    .Y(_03483_),
    .A2(_03475_),
    .A1(_03472_));
 sg13g2_nand3b_1 _09589_ (.B(net2897),
    .C(_03482_),
    .Y(_03484_),
    .A_N(_03483_));
 sg13g2_nand2_1 _09590_ (.Y(_03485_),
    .A(\u_toplayer.u_layer3.u_neuron.acc[7] ),
    .B(\u_toplayer.u_layer3.u_neuron.mult[7] ));
 sg13g2_xor2_1 _09591_ (.B(\u_toplayer.u_layer3.u_neuron.mult[7] ),
    .A(\u_toplayer.u_layer3.u_neuron.acc[7] ),
    .X(_03486_));
 sg13g2_o21ai_1 _09592_ (.B1(_03486_),
    .Y(_03487_),
    .A1(_03466_),
    .A2(_03470_));
 sg13g2_or3_1 _09593_ (.A(_03466_),
    .B(_03470_),
    .C(_03486_),
    .X(_03488_));
 sg13g2_and2_1 _09594_ (.A(net2863),
    .B(_03487_),
    .X(_03489_));
 sg13g2_a21oi_1 _09595_ (.A1(_03488_),
    .A2(_03489_),
    .Y(_03490_),
    .B1(net2762));
 sg13g2_a22oi_1 _09596_ (.Y(_00356_),
    .B1(_03484_),
    .B2(_03490_),
    .A2(net2762),
    .A1(_01050_));
 sg13g2_nand2_1 _09597_ (.Y(_03491_),
    .A(net3373),
    .B(net3158));
 sg13g2_xor2_1 _09598_ (.B(net3158),
    .A(net3373),
    .X(_03492_));
 sg13g2_o21ai_1 _09599_ (.B1(_03492_),
    .Y(_03493_),
    .A1(_03479_),
    .A2(_03483_));
 sg13g2_or3_1 _09600_ (.A(_03479_),
    .B(_03483_),
    .C(_03492_),
    .X(_03494_));
 sg13g2_nand3_1 _09601_ (.B(_03493_),
    .C(_03494_),
    .A(net2897),
    .Y(_03495_));
 sg13g2_and2_1 _09602_ (.A(_03485_),
    .B(_03487_),
    .X(_03496_));
 sg13g2_nand2_1 _09603_ (.Y(_03497_),
    .A(net3158),
    .B(\u_toplayer.u_layer3.u_neuron.mult[8] ));
 sg13g2_xor2_1 _09604_ (.B(\u_toplayer.u_layer3.u_neuron.mult[8] ),
    .A(net3158),
    .X(_03498_));
 sg13g2_nor2b_1 _09605_ (.A(_03496_),
    .B_N(_03498_),
    .Y(_03499_));
 sg13g2_xnor2_1 _09606_ (.Y(_03500_),
    .A(_03496_),
    .B(_03498_));
 sg13g2_a21oi_1 _09607_ (.A1(net2863),
    .A2(_03500_),
    .Y(_03501_),
    .B1(net2762));
 sg13g2_a22oi_1 _09608_ (.Y(_00357_),
    .B1(_03495_),
    .B2(_03501_),
    .A2(net2763),
    .A1(_01059_));
 sg13g2_nor2_1 _09609_ (.A(\u_toplayer.u_layer3.u_neuron.acc[9] ),
    .B(\u_toplayer.u_layer3.u_neuron.mult[9] ),
    .Y(_03502_));
 sg13g2_or2_1 _09610_ (.X(_03503_),
    .B(\u_toplayer.u_layer3.u_neuron.mult[9] ),
    .A(\u_toplayer.u_layer3.u_neuron.acc[9] ));
 sg13g2_nand2_1 _09611_ (.Y(_03504_),
    .A(\u_toplayer.u_layer3.u_neuron.acc[9] ),
    .B(\u_toplayer.u_layer3.u_neuron.mult[9] ));
 sg13g2_nand2_1 _09612_ (.Y(_03505_),
    .A(_03503_),
    .B(_03504_));
 sg13g2_a21oi_1 _09613_ (.A1(net3158),
    .A2(\u_toplayer.u_layer3.u_neuron.mult[8] ),
    .Y(_03506_),
    .B1(_03499_));
 sg13g2_a21oi_1 _09614_ (.A1(_03505_),
    .A2(_03506_),
    .Y(_03507_),
    .B1(net2865));
 sg13g2_o21ai_1 _09615_ (.B1(_03507_),
    .Y(_03508_),
    .A1(_03505_),
    .A2(_03506_));
 sg13g2_xnor2_1 _09616_ (.Y(_03509_),
    .A(net3373),
    .B(\u_toplayer.u_layer3.u_neuron.acc[9] ));
 sg13g2_a21oi_1 _09617_ (.A1(_03491_),
    .A2(_03493_),
    .Y(_03510_),
    .B1(_03509_));
 sg13g2_nand3_1 _09618_ (.B(_03493_),
    .C(_03509_),
    .A(_03491_),
    .Y(_03511_));
 sg13g2_nor2_1 _09619_ (.A(net2895),
    .B(_03510_),
    .Y(_03512_));
 sg13g2_a21oi_1 _09620_ (.A1(_03511_),
    .A2(_03512_),
    .Y(_03513_),
    .B1(net2763));
 sg13g2_a22oi_1 _09621_ (.Y(_00358_),
    .B1(_03508_),
    .B2(_03513_),
    .A2(net2763),
    .A1(_01058_));
 sg13g2_and2_1 _09622_ (.A(net3374),
    .B(\u_toplayer.u_layer3.u_neuron.acc[10] ),
    .X(_03514_));
 sg13g2_xor2_1 _09623_ (.B(\u_toplayer.u_layer3.u_neuron.acc[10] ),
    .A(net3374),
    .X(_03515_));
 sg13g2_o21ai_1 _09624_ (.B1(net3372),
    .Y(_03516_),
    .A1(\u_toplayer.u_layer3.u_neuron.acc[9] ),
    .A2(net3158));
 sg13g2_o21ai_1 _09625_ (.B1(_03516_),
    .Y(_03517_),
    .A1(_03493_),
    .A2(_03509_));
 sg13g2_and2_1 _09626_ (.A(_03515_),
    .B(_03517_),
    .X(_03518_));
 sg13g2_nand2_1 _09627_ (.Y(_03519_),
    .A(\u_toplayer.u_layer3.u_neuron.acc[10] ),
    .B(\u_toplayer.u_layer3.u_neuron.mult[10] ));
 sg13g2_xnor2_1 _09628_ (.Y(_03520_),
    .A(\u_toplayer.u_layer3.u_neuron.acc[10] ),
    .B(\u_toplayer.u_layer3.u_neuron.mult[10] ));
 sg13g2_nand2_1 _09629_ (.Y(_03521_),
    .A(_03497_),
    .B(_03504_));
 sg13g2_o21ai_1 _09630_ (.B1(_03504_),
    .Y(_03522_),
    .A1(_03497_),
    .A2(_03502_));
 sg13g2_o21ai_1 _09631_ (.B1(_03503_),
    .Y(_03523_),
    .A1(_03499_),
    .A2(_03521_));
 sg13g2_or2_1 _09632_ (.X(_03524_),
    .B(_03523_),
    .A(_03520_));
 sg13g2_a21oi_1 _09633_ (.A1(_03520_),
    .A2(_03523_),
    .Y(_03525_),
    .B1(net2865));
 sg13g2_nand2_1 _09634_ (.Y(_03526_),
    .A(_03524_),
    .B(_03525_));
 sg13g2_o21ai_1 _09635_ (.B1(net2897),
    .Y(_03527_),
    .A1(_03515_),
    .A2(_03517_));
 sg13g2_o21ai_1 _09636_ (.B1(_03526_),
    .Y(_03528_),
    .A1(_03518_),
    .A2(_03527_));
 sg13g2_mux2_1 _09637_ (.A0(net1171),
    .A1(_03528_),
    .S(net2759),
    .X(_00359_));
 sg13g2_nor2_1 _09638_ (.A(\u_toplayer.u_layer3.u_neuron.acc[11] ),
    .B(\u_toplayer.u_layer3.u_neuron.mult[11] ),
    .Y(_03529_));
 sg13g2_xnor2_1 _09639_ (.Y(_03530_),
    .A(\u_toplayer.u_layer3.u_neuron.acc[11] ),
    .B(\u_toplayer.u_layer3.u_neuron.mult[11] ));
 sg13g2_nand3_1 _09640_ (.B(_03524_),
    .C(_03530_),
    .A(_03519_),
    .Y(_03531_));
 sg13g2_a21oi_1 _09641_ (.A1(_03519_),
    .A2(_03524_),
    .Y(_03532_),
    .B1(_03530_));
 sg13g2_nor2_1 _09642_ (.A(net2865),
    .B(_03532_),
    .Y(_03533_));
 sg13g2_xor2_1 _09643_ (.B(\u_toplayer.u_layer3.u_neuron.acc[11] ),
    .A(net3374),
    .X(_03534_));
 sg13g2_or3_1 _09644_ (.A(_03514_),
    .B(_03518_),
    .C(_03534_),
    .X(_03535_));
 sg13g2_o21ai_1 _09645_ (.B1(_03534_),
    .Y(_03536_),
    .A1(_03514_),
    .A2(_03518_));
 sg13g2_nand3_1 _09646_ (.B(_03535_),
    .C(_03536_),
    .A(net2897),
    .Y(_03537_));
 sg13g2_a21oi_1 _09647_ (.A1(_03531_),
    .A2(_03533_),
    .Y(_03538_),
    .B1(net2763));
 sg13g2_a22oi_1 _09648_ (.Y(_00360_),
    .B1(_03537_),
    .B2(_03538_),
    .A2(net2762),
    .A1(_01057_));
 sg13g2_nor2_1 _09649_ (.A(_03519_),
    .B(_03529_),
    .Y(_03539_));
 sg13g2_nor2_1 _09650_ (.A(_03520_),
    .B(_03530_),
    .Y(_03540_));
 sg13g2_a221oi_1 _09651_ (.B2(_03540_),
    .C1(_03539_),
    .B1(_03522_),
    .A1(\u_toplayer.u_layer3.u_neuron.acc[11] ),
    .Y(_03541_),
    .A2(\u_toplayer.u_layer3.u_neuron.mult[11] ));
 sg13g2_nand4_1 _09652_ (.B(_03503_),
    .C(_03504_),
    .A(_03498_),
    .Y(_03542_),
    .D(_03540_));
 sg13g2_o21ai_1 _09653_ (.B1(_03541_),
    .Y(_03543_),
    .A1(_03496_),
    .A2(_03542_));
 sg13g2_nand2_1 _09654_ (.Y(_03544_),
    .A(\u_toplayer.u_layer3.u_neuron.acc[12] ),
    .B(\u_toplayer.u_layer3.u_neuron.mult[12] ));
 sg13g2_xor2_1 _09655_ (.B(\u_toplayer.u_layer3.u_neuron.mult[12] ),
    .A(\u_toplayer.u_layer3.u_neuron.acc[12] ),
    .X(_03545_));
 sg13g2_nand2_1 _09656_ (.Y(_03546_),
    .A(_03543_),
    .B(_03545_));
 sg13g2_o21ai_1 _09657_ (.B1(net2863),
    .Y(_03547_),
    .A1(_03543_),
    .A2(_03545_));
 sg13g2_nand2b_1 _09658_ (.Y(_03548_),
    .B(_03546_),
    .A_N(_03547_));
 sg13g2_xnor2_1 _09659_ (.Y(_03549_),
    .A(net3375),
    .B(\u_toplayer.u_layer3.u_neuron.acc[12] ));
 sg13g2_nand2_1 _09660_ (.Y(_03550_),
    .A(_03515_),
    .B(_03534_));
 sg13g2_nor3_1 _09661_ (.A(_03493_),
    .B(_03509_),
    .C(_03550_),
    .Y(_03551_));
 sg13g2_o21ai_1 _09662_ (.B1(net3374),
    .Y(_03552_),
    .A1(\u_toplayer.u_layer3.u_neuron.acc[10] ),
    .A2(\u_toplayer.u_layer3.u_neuron.acc[11] ));
 sg13g2_nand2_1 _09663_ (.Y(_03553_),
    .A(_03516_),
    .B(_03552_));
 sg13g2_nor2_1 _09664_ (.A(_03551_),
    .B(_03553_),
    .Y(_03554_));
 sg13g2_nor2_1 _09665_ (.A(_03549_),
    .B(_03554_),
    .Y(_03555_));
 sg13g2_a21o_1 _09666_ (.A2(_03554_),
    .A1(_03549_),
    .B1(net2895),
    .X(_03556_));
 sg13g2_o21ai_1 _09667_ (.B1(_03548_),
    .Y(_03557_),
    .A1(_03555_),
    .A2(_03556_));
 sg13g2_mux2_1 _09668_ (.A0(net1163),
    .A1(_03557_),
    .S(net2759),
    .X(_00361_));
 sg13g2_nor2_1 _09669_ (.A(\u_toplayer.u_layer3.u_neuron.acc[13] ),
    .B(\u_toplayer.u_layer3.u_neuron.mult[13] ),
    .Y(_03558_));
 sg13g2_nand2_1 _09670_ (.Y(_03559_),
    .A(\u_toplayer.u_layer3.u_neuron.acc[13] ),
    .B(\u_toplayer.u_layer3.u_neuron.mult[13] ));
 sg13g2_nor2b_1 _09671_ (.A(_03558_),
    .B_N(_03559_),
    .Y(_03560_));
 sg13g2_nand2_1 _09672_ (.Y(_03561_),
    .A(_03544_),
    .B(_03546_));
 sg13g2_o21ai_1 _09673_ (.B1(net2862),
    .Y(_03562_),
    .A1(_03560_),
    .A2(_03561_));
 sg13g2_a21oi_1 _09674_ (.A1(_03560_),
    .A2(_03561_),
    .Y(_03563_),
    .B1(_03562_));
 sg13g2_xnor2_1 _09675_ (.Y(_03564_),
    .A(net3372),
    .B(\u_toplayer.u_layer3.u_neuron.acc[13] ));
 sg13g2_a21oi_1 _09676_ (.A1(net3374),
    .A2(\u_toplayer.u_layer3.u_neuron.acc[12] ),
    .Y(_03565_),
    .B1(_03555_));
 sg13g2_a21oi_1 _09677_ (.A1(_03564_),
    .A2(_03565_),
    .Y(_03566_),
    .B1(net2894));
 sg13g2_o21ai_1 _09678_ (.B1(_03566_),
    .Y(_03567_),
    .A1(_03564_),
    .A2(_03565_));
 sg13g2_nor2_1 _09679_ (.A(net2762),
    .B(_03563_),
    .Y(_03568_));
 sg13g2_a22oi_1 _09680_ (.Y(_00362_),
    .B1(_03567_),
    .B2(_03568_),
    .A2(net2762),
    .A1(_01056_));
 sg13g2_nand2_1 _09681_ (.Y(_03569_),
    .A(net3372),
    .B(net3157));
 sg13g2_xnor2_1 _09682_ (.Y(_03570_),
    .A(net3372),
    .B(net3157));
 sg13g2_o21ai_1 _09683_ (.B1(net3372),
    .Y(_03571_),
    .A1(\u_toplayer.u_layer3.u_neuron.acc[12] ),
    .A2(\u_toplayer.u_layer3.u_neuron.acc[13] ));
 sg13g2_nor3_1 _09684_ (.A(_03549_),
    .B(_03554_),
    .C(_03564_),
    .Y(_03572_));
 sg13g2_nor2b_1 _09685_ (.A(_03572_),
    .B_N(_03571_),
    .Y(_03573_));
 sg13g2_or2_1 _09686_ (.X(_03574_),
    .B(_03573_),
    .A(_03570_));
 sg13g2_a21oi_1 _09687_ (.A1(_03570_),
    .A2(_03573_),
    .Y(_03575_),
    .B1(net2894));
 sg13g2_nand2_1 _09688_ (.Y(_03576_),
    .A(net3157),
    .B(\u_toplayer.u_layer3.u_neuron.mult[14] ));
 sg13g2_xor2_1 _09689_ (.B(\u_toplayer.u_layer3.u_neuron.mult[14] ),
    .A(net3157),
    .X(_03577_));
 sg13g2_inv_1 _09690_ (.Y(_03578_),
    .A(_03577_));
 sg13g2_and2_1 _09691_ (.A(_03545_),
    .B(_03560_),
    .X(_03579_));
 sg13g2_o21ai_1 _09692_ (.B1(_03559_),
    .Y(_03580_),
    .A1(_03544_),
    .A2(_03558_));
 sg13g2_a21o_1 _09693_ (.A2(_03579_),
    .A1(_03543_),
    .B1(_03580_),
    .X(_03581_));
 sg13g2_and2_1 _09694_ (.A(_03577_),
    .B(_03581_),
    .X(_03582_));
 sg13g2_o21ai_1 _09695_ (.B1(net2862),
    .Y(_03583_),
    .A1(_03577_),
    .A2(_03581_));
 sg13g2_o21ai_1 _09696_ (.B1(net2758),
    .Y(_03584_),
    .A1(_03582_),
    .A2(_03583_));
 sg13g2_a21oi_1 _09697_ (.A1(_03574_),
    .A2(_03575_),
    .Y(_03585_),
    .B1(_03584_));
 sg13g2_a21oi_1 _09698_ (.A1(_01054_),
    .A2(net2761),
    .Y(_00363_),
    .B1(_03585_));
 sg13g2_nor2_1 _09699_ (.A(\u_toplayer.u_layer3.u_neuron.acc[15] ),
    .B(net3203),
    .Y(_03586_));
 sg13g2_nand2_1 _09700_ (.Y(_03587_),
    .A(\u_toplayer.u_layer3.u_neuron.acc[15] ),
    .B(net3203));
 sg13g2_nand2b_1 _09701_ (.Y(_03588_),
    .B(_03587_),
    .A_N(_03586_));
 sg13g2_a21oi_1 _09702_ (.A1(net3157),
    .A2(\u_toplayer.u_layer3.u_neuron.mult[14] ),
    .Y(_03589_),
    .B1(_03582_));
 sg13g2_a21oi_1 _09703_ (.A1(_03588_),
    .A2(_03589_),
    .Y(_03590_),
    .B1(net2864));
 sg13g2_o21ai_1 _09704_ (.B1(_03590_),
    .Y(_03591_),
    .A1(_03588_),
    .A2(_03589_));
 sg13g2_xnor2_1 _09705_ (.Y(_03592_),
    .A(net3372),
    .B(\u_toplayer.u_layer3.u_neuron.acc[15] ));
 sg13g2_nand3_1 _09706_ (.B(_03574_),
    .C(_03592_),
    .A(_03569_),
    .Y(_03593_));
 sg13g2_a21oi_1 _09707_ (.A1(_03569_),
    .A2(_03574_),
    .Y(_03594_),
    .B1(_03592_));
 sg13g2_nor2_1 _09708_ (.A(net2894),
    .B(_03594_),
    .Y(_03595_));
 sg13g2_a21oi_1 _09709_ (.A1(_03593_),
    .A2(_03595_),
    .Y(_03596_),
    .B1(net2761));
 sg13g2_a22oi_1 _09710_ (.Y(_00364_),
    .B1(_03591_),
    .B2(_03596_),
    .A2(net2761),
    .A1(_01055_));
 sg13g2_nor2_1 _09711_ (.A(net721),
    .B(net2758),
    .Y(_03597_));
 sg13g2_nand2_1 _09712_ (.Y(_03598_),
    .A(net3156),
    .B(net3204));
 sg13g2_xnor2_1 _09713_ (.Y(_03599_),
    .A(net3156),
    .B(net3204));
 sg13g2_o21ai_1 _09714_ (.B1(_03587_),
    .Y(_03600_),
    .A1(_03576_),
    .A2(_03586_));
 sg13g2_nor2_1 _09715_ (.A(_03578_),
    .B(_03588_),
    .Y(_03601_));
 sg13g2_and2_1 _09716_ (.A(_03579_),
    .B(_03601_),
    .X(_03602_));
 sg13g2_a221oi_1 _09717_ (.B2(_03543_),
    .C1(_03600_),
    .B1(_03602_),
    .A1(_03580_),
    .Y(_03603_),
    .A2(_03601_));
 sg13g2_or2_1 _09718_ (.X(_03604_),
    .B(_03603_),
    .A(_03599_));
 sg13g2_a21oi_1 _09719_ (.A1(_03599_),
    .A2(_03603_),
    .Y(_03605_),
    .B1(net2864));
 sg13g2_nor4_1 _09720_ (.A(_03549_),
    .B(_03564_),
    .C(_03570_),
    .D(_03592_),
    .Y(_03606_));
 sg13g2_inv_1 _09721_ (.Y(_03607_),
    .A(_03606_));
 sg13g2_nor4_2 _09722_ (.A(_03493_),
    .B(_03509_),
    .C(_03550_),
    .Y(_03608_),
    .D(_03607_));
 sg13g2_o21ai_1 _09723_ (.B1(net3372),
    .Y(_03609_),
    .A1(\u_toplayer.u_layer3.u_neuron.acc[14] ),
    .A2(\u_toplayer.u_layer3.u_neuron.acc[15] ));
 sg13g2_nand4_1 _09724_ (.B(_03552_),
    .C(_03571_),
    .A(_03516_),
    .Y(_03610_),
    .D(_03609_));
 sg13g2_xnor2_1 _09725_ (.Y(_03611_),
    .A(net3374),
    .B(net3156));
 sg13g2_inv_1 _09726_ (.Y(_03612_),
    .A(_03611_));
 sg13g2_o21ai_1 _09727_ (.B1(_03612_),
    .Y(_03613_),
    .A1(_03608_),
    .A2(_03610_));
 sg13g2_inv_1 _09728_ (.Y(_03614_),
    .A(_03613_));
 sg13g2_nor3_1 _09729_ (.A(_03608_),
    .B(_03610_),
    .C(_03612_),
    .Y(_03615_));
 sg13g2_nor2_1 _09730_ (.A(net2895),
    .B(_03615_),
    .Y(_03616_));
 sg13g2_a22oi_1 _09731_ (.Y(_03617_),
    .B1(_03613_),
    .B2(_03616_),
    .A2(_03605_),
    .A1(_03604_));
 sg13g2_a21oi_1 _09732_ (.A1(net2758),
    .A2(_03617_),
    .Y(_00365_),
    .B1(_03597_));
 sg13g2_nor2_1 _09733_ (.A(net1046),
    .B(net2758),
    .Y(_03618_));
 sg13g2_xnor2_1 _09734_ (.Y(_03619_),
    .A(\u_toplayer.u_layer3.u_neuron.acc[17] ),
    .B(net3203));
 sg13g2_a21oi_1 _09735_ (.A1(_03598_),
    .A2(_03604_),
    .Y(_03620_),
    .B1(_03619_));
 sg13g2_nand3_1 _09736_ (.B(_03604_),
    .C(_03619_),
    .A(_03598_),
    .Y(_03621_));
 sg13g2_nor2_1 _09737_ (.A(net2864),
    .B(_03620_),
    .Y(_03622_));
 sg13g2_xnor2_1 _09738_ (.Y(_03623_),
    .A(net3371),
    .B(\u_toplayer.u_layer3.u_neuron.acc[17] ));
 sg13g2_a21oi_1 _09739_ (.A1(net3375),
    .A2(net3156),
    .Y(_03624_),
    .B1(_03614_));
 sg13g2_o21ai_1 _09740_ (.B1(net2897),
    .Y(_03625_),
    .A1(_03623_),
    .A2(_03624_));
 sg13g2_a21oi_1 _09741_ (.A1(_03623_),
    .A2(_03624_),
    .Y(_03626_),
    .B1(_03625_));
 sg13g2_a21oi_1 _09742_ (.A1(_03621_),
    .A2(_03622_),
    .Y(_03627_),
    .B1(_03626_));
 sg13g2_a21oi_1 _09743_ (.A1(net2758),
    .A2(_03627_),
    .Y(_00366_),
    .B1(_03618_));
 sg13g2_nand2_1 _09744_ (.Y(_03628_),
    .A(net3155),
    .B(net3203));
 sg13g2_xnor2_1 _09745_ (.Y(_03629_),
    .A(\u_toplayer.u_layer3.u_neuron.acc[18] ),
    .B(net3203));
 sg13g2_or3_1 _09746_ (.A(_03599_),
    .B(_03603_),
    .C(_03619_),
    .X(_03630_));
 sg13g2_o21ai_1 _09747_ (.B1(net3203),
    .Y(_03631_),
    .A1(net3156),
    .A2(\u_toplayer.u_layer3.u_neuron.acc[17] ));
 sg13g2_and2_1 _09748_ (.A(_03630_),
    .B(_03631_),
    .X(_03632_));
 sg13g2_or2_1 _09749_ (.X(_03633_),
    .B(_03632_),
    .A(_03629_));
 sg13g2_a21oi_1 _09750_ (.A1(_03629_),
    .A2(_03632_),
    .Y(_03634_),
    .B1(net2865));
 sg13g2_xor2_1 _09751_ (.B(net3155),
    .A(net3371),
    .X(_03635_));
 sg13g2_nor2_1 _09752_ (.A(_03611_),
    .B(_03623_),
    .Y(_03636_));
 sg13g2_o21ai_1 _09753_ (.B1(_03636_),
    .Y(_03637_),
    .A1(_03608_),
    .A2(_03610_));
 sg13g2_o21ai_1 _09754_ (.B1(net3371),
    .Y(_03638_),
    .A1(net3156),
    .A2(\u_toplayer.u_layer3.u_neuron.acc[17] ));
 sg13g2_nand2_1 _09755_ (.Y(_03639_),
    .A(_03637_),
    .B(_03638_));
 sg13g2_and2_1 _09756_ (.A(_03635_),
    .B(_03639_),
    .X(_03640_));
 sg13g2_o21ai_1 _09757_ (.B1(net2896),
    .Y(_03641_),
    .A1(_03635_),
    .A2(_03639_));
 sg13g2_o21ai_1 _09758_ (.B1(net2758),
    .Y(_03642_),
    .A1(_03640_),
    .A2(_03641_));
 sg13g2_a21oi_1 _09759_ (.A1(_03633_),
    .A2(_03634_),
    .Y(_03643_),
    .B1(_03642_));
 sg13g2_a21oi_1 _09760_ (.A1(_01064_),
    .A2(net2761),
    .Y(_00367_),
    .B1(_03643_));
 sg13g2_nor2_1 _09761_ (.A(net1052),
    .B(net2758),
    .Y(_03644_));
 sg13g2_xnor2_1 _09762_ (.Y(_03645_),
    .A(\u_toplayer.u_layer3.u_neuron.acc[19] ),
    .B(net3203));
 sg13g2_a21oi_1 _09763_ (.A1(_03628_),
    .A2(_03633_),
    .Y(_03646_),
    .B1(_03645_));
 sg13g2_nand3_1 _09764_ (.B(_03633_),
    .C(_03645_),
    .A(_03628_),
    .Y(_03647_));
 sg13g2_nor2_1 _09765_ (.A(net2864),
    .B(_03646_),
    .Y(_03648_));
 sg13g2_xnor2_1 _09766_ (.Y(_03649_),
    .A(net3370),
    .B(\u_toplayer.u_layer3.u_neuron.acc[19] ));
 sg13g2_inv_1 _09767_ (.Y(_03650_),
    .A(_03649_));
 sg13g2_a21oi_1 _09768_ (.A1(net3370),
    .A2(net3155),
    .Y(_03651_),
    .B1(_03640_));
 sg13g2_o21ai_1 _09769_ (.B1(net2896),
    .Y(_03652_),
    .A1(_03649_),
    .A2(_03651_));
 sg13g2_a21oi_1 _09770_ (.A1(_03649_),
    .A2(_03651_),
    .Y(_03653_),
    .B1(_03652_));
 sg13g2_a21oi_1 _09771_ (.A1(_03647_),
    .A2(_03648_),
    .Y(_03654_),
    .B1(_03653_));
 sg13g2_a21oi_1 _09772_ (.A1(net2758),
    .A2(_03654_),
    .Y(_00368_),
    .B1(_03644_));
 sg13g2_or2_1 _09773_ (.X(_03655_),
    .B(_03645_),
    .A(_03629_));
 sg13g2_nor4_1 _09774_ (.A(_03599_),
    .B(_03603_),
    .C(_03619_),
    .D(_03655_),
    .Y(_03656_));
 sg13g2_o21ai_1 _09775_ (.B1(net3202),
    .Y(_03657_),
    .A1(\u_toplayer.u_layer3.u_neuron.acc[19] ),
    .A2(net3155));
 sg13g2_nand2_1 _09776_ (.Y(_03658_),
    .A(_03631_),
    .B(_03657_));
 sg13g2_nor2_2 _09777_ (.A(_03656_),
    .B(_03658_),
    .Y(_03659_));
 sg13g2_nand2_1 _09778_ (.Y(_03660_),
    .A(net3154),
    .B(net3202));
 sg13g2_xor2_1 _09779_ (.B(net3202),
    .A(net3154),
    .X(_03661_));
 sg13g2_inv_1 _09780_ (.Y(_03662_),
    .A(_03661_));
 sg13g2_a21oi_1 _09781_ (.A1(_03659_),
    .A2(_03662_),
    .Y(_03663_),
    .B1(net2864));
 sg13g2_o21ai_1 _09782_ (.B1(_03663_),
    .Y(_03664_),
    .A1(_03659_),
    .A2(_03662_));
 sg13g2_nand2_1 _09783_ (.Y(_03665_),
    .A(net3370),
    .B(net3154));
 sg13g2_xor2_1 _09784_ (.B(net3154),
    .A(net3370),
    .X(_03666_));
 sg13g2_inv_1 _09785_ (.Y(_03667_),
    .A(_03666_));
 sg13g2_nand2_1 _09786_ (.Y(_03668_),
    .A(_03635_),
    .B(_03650_));
 sg13g2_nor2_1 _09787_ (.A(_03637_),
    .B(_03668_),
    .Y(_03669_));
 sg13g2_o21ai_1 _09788_ (.B1(net3371),
    .Y(_03670_),
    .A1(\u_toplayer.u_layer3.u_neuron.acc[19] ),
    .A2(net3155));
 sg13g2_and2_1 _09789_ (.A(_03638_),
    .B(_03670_),
    .X(_03671_));
 sg13g2_nor2b_1 _09790_ (.A(_03669_),
    .B_N(_03671_),
    .Y(_03672_));
 sg13g2_o21ai_1 _09791_ (.B1(_03671_),
    .Y(_03673_),
    .A1(_03637_),
    .A2(_03668_));
 sg13g2_nand2_1 _09792_ (.Y(_03674_),
    .A(_03666_),
    .B(_03673_));
 sg13g2_a21oi_1 _09793_ (.A1(_03667_),
    .A2(_03672_),
    .Y(_03675_),
    .B1(net2894));
 sg13g2_a21oi_1 _09794_ (.A1(_03674_),
    .A2(_03675_),
    .Y(_03676_),
    .B1(net2760));
 sg13g2_a22oi_1 _09795_ (.Y(_00369_),
    .B1(_03664_),
    .B2(_03676_),
    .A2(net2760),
    .A1(_01063_));
 sg13g2_xor2_1 _09796_ (.B(net3202),
    .A(\u_toplayer.u_layer3.u_neuron.acc[21] ),
    .X(_03677_));
 sg13g2_o21ai_1 _09797_ (.B1(_03660_),
    .Y(_03678_),
    .A1(_03659_),
    .A2(_03662_));
 sg13g2_a21oi_1 _09798_ (.A1(_03677_),
    .A2(_03678_),
    .Y(_03679_),
    .B1(net2864));
 sg13g2_o21ai_1 _09799_ (.B1(_03679_),
    .Y(_03680_),
    .A1(_03677_),
    .A2(_03678_));
 sg13g2_xnor2_1 _09800_ (.Y(_03681_),
    .A(net2),
    .B(\u_toplayer.u_layer3.u_neuron.acc[21] ));
 sg13g2_inv_1 _09801_ (.Y(_03682_),
    .A(_03681_));
 sg13g2_nand3_1 _09802_ (.B(_03674_),
    .C(_03681_),
    .A(_03665_),
    .Y(_03683_));
 sg13g2_a21oi_1 _09803_ (.A1(_03665_),
    .A2(_03674_),
    .Y(_03684_),
    .B1(_03681_));
 sg13g2_nor2_1 _09804_ (.A(net2894),
    .B(_03684_),
    .Y(_03685_));
 sg13g2_a21oi_1 _09805_ (.A1(_03683_),
    .A2(_03685_),
    .Y(_03686_),
    .B1(net2760));
 sg13g2_a22oi_1 _09806_ (.Y(_00370_),
    .B1(_03680_),
    .B2(_03686_),
    .A2(net2760),
    .A1(_01062_));
 sg13g2_and2_1 _09807_ (.A(\u_toplayer.u_layer3.u_neuron.acc[22] ),
    .B(net3202),
    .X(_03687_));
 sg13g2_xor2_1 _09808_ (.B(net3202),
    .A(\u_toplayer.u_layer3.u_neuron.acc[22] ),
    .X(_03688_));
 sg13g2_nand2_1 _09809_ (.Y(_03689_),
    .A(_03661_),
    .B(_03677_));
 sg13g2_o21ai_1 _09810_ (.B1(net3202),
    .Y(_03690_),
    .A1(\u_toplayer.u_layer3.u_neuron.acc[21] ),
    .A2(net3154));
 sg13g2_o21ai_1 _09811_ (.B1(_03690_),
    .Y(_03691_),
    .A1(_03659_),
    .A2(_03689_));
 sg13g2_nor2_1 _09812_ (.A(_03688_),
    .B(_03691_),
    .Y(_03692_));
 sg13g2_nand2_1 _09813_ (.Y(_03693_),
    .A(_03688_),
    .B(_03691_));
 sg13g2_nor2_1 _09814_ (.A(net2864),
    .B(_03692_),
    .Y(_03694_));
 sg13g2_nand3_1 _09815_ (.B(_03673_),
    .C(_03682_),
    .A(_03666_),
    .Y(_03695_));
 sg13g2_o21ai_1 _09816_ (.B1(net3370),
    .Y(_03696_),
    .A1(\u_toplayer.u_layer3.u_neuron.acc[21] ),
    .A2(net3154));
 sg13g2_nand2_1 _09817_ (.Y(_03697_),
    .A(net3370),
    .B(\u_toplayer.u_layer3.u_neuron.acc[22] ));
 sg13g2_xnor2_1 _09818_ (.Y(_03698_),
    .A(net3370),
    .B(\u_toplayer.u_layer3.u_neuron.acc[22] ));
 sg13g2_a21o_1 _09819_ (.A2(_03696_),
    .A1(_03695_),
    .B1(_03698_),
    .X(_03699_));
 sg13g2_nand3_1 _09820_ (.B(_03696_),
    .C(_03698_),
    .A(_03695_),
    .Y(_03700_));
 sg13g2_nand3_1 _09821_ (.B(_03699_),
    .C(_03700_),
    .A(net2896),
    .Y(_03701_));
 sg13g2_a21oi_1 _09822_ (.A1(_03693_),
    .A2(_03694_),
    .Y(_03702_),
    .B1(net2761));
 sg13g2_a22oi_1 _09823_ (.Y(_00371_),
    .B1(_03701_),
    .B2(_03702_),
    .A2(net2760),
    .A1(_01060_));
 sg13g2_a21oi_1 _09824_ (.A1(_03688_),
    .A2(_03691_),
    .Y(_03703_),
    .B1(_03687_));
 sg13g2_xnor2_1 _09825_ (.Y(_03704_),
    .A(\u_toplayer.u_layer3.u_neuron.acc[23] ),
    .B(net3202));
 sg13g2_a21oi_1 _09826_ (.A1(_03703_),
    .A2(_03704_),
    .Y(_03705_),
    .B1(net2864));
 sg13g2_o21ai_1 _09827_ (.B1(_03705_),
    .Y(_03706_),
    .A1(_03703_),
    .A2(_03704_));
 sg13g2_xnor2_1 _09828_ (.Y(_03707_),
    .A(net3370),
    .B(\u_toplayer.u_layer3.u_neuron.acc[23] ));
 sg13g2_a21oi_1 _09829_ (.A1(_03697_),
    .A2(_03699_),
    .Y(_03708_),
    .B1(_03707_));
 sg13g2_nand3_1 _09830_ (.B(_03699_),
    .C(_03707_),
    .A(_03697_),
    .Y(_03709_));
 sg13g2_nor2_1 _09831_ (.A(net2894),
    .B(_03708_),
    .Y(_03710_));
 sg13g2_a21oi_1 _09832_ (.A1(_03709_),
    .A2(_03710_),
    .Y(_03711_),
    .B1(net2760));
 sg13g2_a22oi_1 _09833_ (.Y(_00372_),
    .B1(_03706_),
    .B2(_03711_),
    .A2(net2760),
    .A1(_01061_));
 sg13g2_nor2_1 _09834_ (.A(\u_toplayer.u_layer2.statel2[3] ),
    .B(\u_toplayer.u_layer2.statel2[1] ),
    .Y(_03712_));
 sg13g2_nand3_1 _09835_ (.B(\u_toplayer.u_layer2.statel2[2] ),
    .C(_03712_),
    .A(net860),
    .Y(_03713_));
 sg13g2_nand3b_1 _09836_ (.B(net122),
    .C(net937),
    .Y(_03714_),
    .A_N(\u_toplayer.u_layer2.statel2[4] ));
 sg13g2_or2_2 _09837_ (.X(_03715_),
    .B(net128),
    .A(net132));
 sg13g2_nand2_1 _09838_ (.Y(_03716_),
    .A(_01024_),
    .B(\u_toplayer.delayed_done_layer1 ));
 sg13g2_nor4_2 _09839_ (.A(_03713_),
    .B(_03714_),
    .C(_03715_),
    .Y(_03717_),
    .D(_03716_));
 sg13g2_and2_1 _09840_ (.A(\u_toplayer.u_layer2.statel2[1] ),
    .B(\u_toplayer.u_layer2.statel2[2] ),
    .X(_03718_));
 sg13g2_or2_1 _09841_ (.X(_03719_),
    .B(\u_toplayer.u_layer2.statel2[3] ),
    .A(\u_toplayer.u_layer2.statel2[4] ));
 sg13g2_o21ai_1 _09842_ (.B1(\u_toplayer.u_layer2.statel2[5] ),
    .Y(_03720_),
    .A1(_03718_),
    .A2(_03719_));
 sg13g2_nor2_1 _09843_ (.A(\u_toplayer.u_layer2.statel2[8] ),
    .B(_03715_),
    .Y(_03721_));
 sg13g2_nand4_1 _09844_ (.B(\u_toplayer.delayed_done_layer1 ),
    .C(_03720_),
    .A(_01024_),
    .Y(_03722_),
    .D(_03721_));
 sg13g2_or2_1 _09845_ (.X(_03723_),
    .B(_03716_),
    .A(\u_toplayer.u_layer2.statel2[4] ));
 sg13g2_nand2_1 _09846_ (.Y(_03724_),
    .A(\u_toplayer.u_layer2.statel2[5] ),
    .B(_00031_));
 sg13g2_nor4_1 _09847_ (.A(_03713_),
    .B(_03715_),
    .C(_03723_),
    .D(_03724_),
    .Y(_03725_));
 sg13g2_nand2b_2 _09848_ (.Y(_03726_),
    .B(_03722_),
    .A_N(_03717_));
 sg13g2_and2_1 _09849_ (.A(net860),
    .B(_03726_),
    .X(_03727_));
 sg13g2_and2_1 _09850_ (.A(net954),
    .B(_03727_),
    .X(_03728_));
 sg13g2_nor2_1 _09851_ (.A(net1009),
    .B(_03728_),
    .Y(_03729_));
 sg13g2_and2_1 _09852_ (.A(_03718_),
    .B(_03727_),
    .X(_03730_));
 sg13g2_nor3_1 _09853_ (.A(_03717_),
    .B(_03729_),
    .C(_03730_),
    .Y(_00670_));
 sg13g2_nor4_2 _09854_ (.A(\u_toplayer.u_layer2.statel2[8] ),
    .B(_03713_),
    .C(_03715_),
    .Y(_03731_),
    .D(_00670_));
 sg13g2_and2_2 _09855_ (.A(_03721_),
    .B(_03725_),
    .X(_03732_));
 sg13g2_mux2_1 _09856_ (.A0(\u_toplayer.u_layer2.neuron_index[0] ),
    .A1(net734),
    .S(_03732_),
    .X(_00373_));
 sg13g2_nor2b_2 _09857_ (.A(\u_toplayer.u_layer2.neuron_index[1] ),
    .B_N(\u_toplayer.u_layer2.neuron_index[0] ),
    .Y(_03733_));
 sg13g2_nor2_2 _09858_ (.A(_01032_),
    .B(\u_toplayer.u_layer2.neuron_index[0] ),
    .Y(_03734_));
 sg13g2_o21ai_1 _09859_ (.B1(_03732_),
    .Y(_03735_),
    .A1(_03733_),
    .A2(net2931));
 sg13g2_o21ai_1 _09860_ (.B1(_03735_),
    .Y(_00374_),
    .A1(_01032_),
    .A2(_03732_));
 sg13g2_nand2_2 _09861_ (.Y(_03736_),
    .A(\u_toplayer.u_layer2.neuron_index[1] ),
    .B(\u_toplayer.u_layer2.neuron_index[0] ));
 sg13g2_nand3_1 _09862_ (.B(\u_toplayer.u_layer2.neuron_index[0] ),
    .C(_03732_),
    .A(net1149),
    .Y(_03737_));
 sg13g2_nor2_1 _09863_ (.A(_01033_),
    .B(_03736_),
    .Y(_03738_));
 sg13g2_xnor2_1 _09864_ (.Y(_00375_),
    .A(net3149),
    .B(net1150));
 sg13g2_and3_2 _09865_ (.X(_03739_),
    .A(net3145),
    .B(_03732_),
    .C(net2926));
 sg13g2_a21oi_1 _09866_ (.A1(_03732_),
    .A2(net2926),
    .Y(_03740_),
    .B1(net3145));
 sg13g2_nor2_1 _09867_ (.A(_03739_),
    .B(_03740_),
    .Y(_00376_));
 sg13g2_nand2_1 _09868_ (.Y(_03741_),
    .A(\u_toplayer.u_layer2.neuron_index[4] ),
    .B(_03739_));
 sg13g2_xor2_1 _09869_ (.B(_03739_),
    .A(net1075),
    .X(_00377_));
 sg13g2_or2_2 _09870_ (.X(_03742_),
    .B(_03741_),
    .A(\u_toplayer.u_layer2.neuron_index[5] ));
 sg13g2_xnor2_1 _09871_ (.Y(_00378_),
    .A(net982),
    .B(_03741_));
 sg13g2_nor2b_1 _09872_ (.A(net770),
    .B_N(_01362_),
    .Y(_03743_));
 sg13g2_nor4_1 _09873_ (.A(\u_toplayer.u_layer1.u_neuron.instCtrl.state[0] ),
    .B(\u_toplayer.u_layer1.u_neuron.instCtrl.state[2] ),
    .C(\u_toplayer.u_layer1.u_neuron.instCtrl.state[1] ),
    .D(\u_toplayer.u_layer1.u_neuron.instCtrl.state[3] ),
    .Y(_03744_));
 sg13g2_and2_1 _09874_ (.A(_03743_),
    .B(_03744_),
    .X(_03745_));
 sg13g2_nand2_2 _09875_ (.Y(_03746_),
    .A(net3230),
    .B(_03745_));
 sg13g2_or2_1 _09876_ (.X(_03747_),
    .B(_03745_),
    .A(net3229));
 sg13g2_nand2_2 _09877_ (.Y(_03748_),
    .A(_01363_),
    .B(_03743_));
 sg13g2_nor2b_1 _09878_ (.A(_03748_),
    .B_N(_01366_),
    .Y(_03749_));
 sg13g2_o21ai_1 _09879_ (.B1(net2857),
    .Y(_03750_),
    .A1(_03747_),
    .A2(_03749_));
 sg13g2_nor2_1 _09880_ (.A(_01365_),
    .B(_03748_),
    .Y(_03751_));
 sg13g2_or2_1 _09881_ (.X(_03752_),
    .B(_03748_),
    .A(_01365_));
 sg13g2_nor2_2 _09882_ (.A(net2832),
    .B(net2855),
    .Y(_03753_));
 sg13g2_nand2b_1 _09883_ (.Y(_03754_),
    .B(net2853),
    .A_N(net2831));
 sg13g2_nand2_1 _09884_ (.Y(_03755_),
    .A(net825),
    .B(net2815));
 sg13g2_nand2_1 _09885_ (.Y(_03756_),
    .A(net3229),
    .B(_03753_));
 sg13g2_nand2_1 _09886_ (.Y(_03757_),
    .A(net3403),
    .B(net3355));
 sg13g2_o21ai_1 _09887_ (.B1(_03755_),
    .Y(_00379_),
    .A1(net2747),
    .A2(_03757_));
 sg13g2_nand4_1 _09888_ (.B(net3398),
    .C(net3352),
    .A(net3402),
    .Y(_03758_),
    .D(net3343));
 sg13g2_a22oi_1 _09889_ (.Y(_03759_),
    .B1(net3343),
    .B2(net3401),
    .A2(net3351),
    .A1(net3398));
 sg13g2_nor2_1 _09890_ (.A(net2745),
    .B(_03759_),
    .Y(_03760_));
 sg13g2_a22oi_1 _09891_ (.Y(_03761_),
    .B1(_03758_),
    .B2(_03760_),
    .A2(net2814),
    .A1(net986));
 sg13g2_inv_1 _09892_ (.Y(_00380_),
    .A(_03761_));
 sg13g2_nand2_1 _09893_ (.Y(_03762_),
    .A(net769),
    .B(net2814));
 sg13g2_and4_2 _09894_ (.A(net3401),
    .B(net3397),
    .C(net3343),
    .D(net3329),
    .X(_03763_));
 sg13g2_a22oi_1 _09895_ (.Y(_03764_),
    .B1(net3329),
    .B2(net3401),
    .A2(net3343),
    .A1(net3397));
 sg13g2_nand2_1 _09896_ (.Y(_03765_),
    .A(net3394),
    .B(net3351));
 sg13g2_nor3_2 _09897_ (.A(_03763_),
    .B(_03764_),
    .C(_03765_),
    .Y(_03766_));
 sg13g2_o21ai_1 _09898_ (.B1(_03765_),
    .Y(_03767_),
    .A1(_03763_),
    .A2(_03764_));
 sg13g2_nand2b_1 _09899_ (.Y(_03768_),
    .B(_03767_),
    .A_N(_03766_));
 sg13g2_or2_1 _09900_ (.X(_03769_),
    .B(_03768_),
    .A(_03758_));
 sg13g2_xnor2_1 _09901_ (.Y(_03770_),
    .A(_03758_),
    .B(_03768_));
 sg13g2_o21ai_1 _09902_ (.B1(_03762_),
    .Y(_00381_),
    .A1(net2745),
    .A2(_03770_));
 sg13g2_nand2_1 _09903_ (.Y(_03771_),
    .A(net3391),
    .B(net3351));
 sg13g2_nand2_1 _09904_ (.Y(_03772_),
    .A(net3394),
    .B(net3343));
 sg13g2_and4_1 _09905_ (.A(net3401),
    .B(net3397),
    .C(net3329),
    .D(net3318),
    .X(_03773_));
 sg13g2_nand4_1 _09906_ (.B(net3397),
    .C(net3325),
    .A(net3401),
    .Y(_03774_),
    .D(net3318));
 sg13g2_a22oi_1 _09907_ (.Y(_03775_),
    .B1(net3318),
    .B2(net3401),
    .A2(net3329),
    .A1(net3397));
 sg13g2_or3_1 _09908_ (.A(_03772_),
    .B(_03773_),
    .C(_03775_),
    .X(_03776_));
 sg13g2_o21ai_1 _09909_ (.B1(_03772_),
    .Y(_03777_),
    .A1(_03773_),
    .A2(_03775_));
 sg13g2_and3_1 _09910_ (.X(_03778_),
    .A(_03763_),
    .B(_03776_),
    .C(_03777_));
 sg13g2_nand3_1 _09911_ (.B(_03776_),
    .C(_03777_),
    .A(_03763_),
    .Y(_03779_));
 sg13g2_a21oi_1 _09912_ (.A1(_03776_),
    .A2(_03777_),
    .Y(_03780_),
    .B1(_03763_));
 sg13g2_nor2_1 _09913_ (.A(_03778_),
    .B(_03780_),
    .Y(_03781_));
 sg13g2_xnor2_1 _09914_ (.Y(_03782_),
    .A(_03771_),
    .B(_03781_));
 sg13g2_and2_1 _09915_ (.A(_03766_),
    .B(_03782_),
    .X(_03783_));
 sg13g2_xnor2_1 _09916_ (.Y(_03784_),
    .A(_03766_),
    .B(_03782_));
 sg13g2_or2_1 _09917_ (.X(_03785_),
    .B(_03784_),
    .A(_03769_));
 sg13g2_nand2b_1 _09918_ (.Y(_03786_),
    .B(_03785_),
    .A_N(net2745));
 sg13g2_a21oi_1 _09919_ (.A1(_03769_),
    .A2(_03784_),
    .Y(_03787_),
    .B1(_03786_));
 sg13g2_a21o_1 _09920_ (.A2(net2814),
    .A1(net953),
    .B1(_03787_),
    .X(_00382_));
 sg13g2_o21ai_1 _09921_ (.B1(_03779_),
    .Y(_03788_),
    .A1(_03771_),
    .A2(_03780_));
 sg13g2_a22oi_1 _09922_ (.Y(_03789_),
    .B1(net3305),
    .B2(net3401),
    .A2(net3351),
    .A1(net3388));
 sg13g2_nand4_1 _09923_ (.B(net3388),
    .C(net3351),
    .A(net3401),
    .Y(_03790_),
    .D(net3305));
 sg13g2_nor2b_1 _09924_ (.A(_03789_),
    .B_N(_03790_),
    .Y(_03791_));
 sg13g2_o21ai_1 _09925_ (.B1(_03774_),
    .Y(_03792_),
    .A1(_03772_),
    .A2(_03775_));
 sg13g2_nand2_1 _09926_ (.Y(_03793_),
    .A(net3391),
    .B(net3336));
 sg13g2_and4_1 _09927_ (.A(net3397),
    .B(net3394),
    .C(net3325),
    .D(net3311),
    .X(_03794_));
 sg13g2_nand4_1 _09928_ (.B(net3394),
    .C(net3325),
    .A(net3397),
    .Y(_03795_),
    .D(net3311));
 sg13g2_a22oi_1 _09929_ (.Y(_03796_),
    .B1(net3311),
    .B2(net3397),
    .A2(net3325),
    .A1(net3394));
 sg13g2_or3_1 _09930_ (.A(_03793_),
    .B(_03794_),
    .C(_03796_),
    .X(_03797_));
 sg13g2_o21ai_1 _09931_ (.B1(_03793_),
    .Y(_03798_),
    .A1(_03794_),
    .A2(_03796_));
 sg13g2_nand3_1 _09932_ (.B(_03797_),
    .C(_03798_),
    .A(_03792_),
    .Y(_03799_));
 sg13g2_a21o_1 _09933_ (.A2(_03798_),
    .A1(_03797_),
    .B1(_03792_),
    .X(_03800_));
 sg13g2_a21oi_1 _09934_ (.A1(_03799_),
    .A2(_03800_),
    .Y(_03801_),
    .B1(_03791_));
 sg13g2_nand3_1 _09935_ (.B(_03799_),
    .C(_03800_),
    .A(_03791_),
    .Y(_03802_));
 sg13g2_nand2b_1 _09936_ (.Y(_03803_),
    .B(_03802_),
    .A_N(_03801_));
 sg13g2_nor2b_1 _09937_ (.A(_03803_),
    .B_N(_03788_),
    .Y(_03804_));
 sg13g2_xnor2_1 _09938_ (.Y(_03805_),
    .A(_03788_),
    .B(_03803_));
 sg13g2_xnor2_1 _09939_ (.Y(_03806_),
    .A(_03783_),
    .B(_03805_));
 sg13g2_nand2b_1 _09940_ (.Y(_03807_),
    .B(_03805_),
    .A_N(_03785_));
 sg13g2_nand2b_1 _09941_ (.Y(_03808_),
    .B(_03807_),
    .A_N(net2745));
 sg13g2_a21oi_1 _09942_ (.A1(_03785_),
    .A2(_03806_),
    .Y(_03809_),
    .B1(_03808_));
 sg13g2_a21o_1 _09943_ (.A2(net2814),
    .A1(net976),
    .B1(_03809_),
    .X(_00383_));
 sg13g2_nand2_1 _09944_ (.Y(_03810_),
    .A(net923),
    .B(net2814));
 sg13g2_nand2_1 _09945_ (.Y(_03811_),
    .A(_03799_),
    .B(_03802_));
 sg13g2_nand2_1 _09946_ (.Y(_03812_),
    .A(net3404),
    .B(net3294));
 sg13g2_and4_1 _09947_ (.A(net3400),
    .B(net3385),
    .C(net3347),
    .D(net3300),
    .X(_03813_));
 sg13g2_a22oi_1 _09948_ (.Y(_03814_),
    .B1(net3300),
    .B2(net3398),
    .A2(net3347),
    .A1(net3385));
 sg13g2_nor3_1 _09949_ (.A(_03812_),
    .B(_03813_),
    .C(_03814_),
    .Y(_03815_));
 sg13g2_o21ai_1 _09950_ (.B1(_03812_),
    .Y(_03816_),
    .A1(_03813_),
    .A2(_03814_));
 sg13g2_nand2b_1 _09951_ (.Y(_03817_),
    .B(_03816_),
    .A_N(_03815_));
 sg13g2_o21ai_1 _09952_ (.B1(_03795_),
    .Y(_03818_),
    .A1(_03793_),
    .A2(_03796_));
 sg13g2_nand2_1 _09953_ (.Y(_03819_),
    .A(net3389),
    .B(net3336));
 sg13g2_and4_1 _09954_ (.A(net3395),
    .B(net3391),
    .C(net3326),
    .D(net3311),
    .X(_03820_));
 sg13g2_nand4_1 _09955_ (.B(net3391),
    .C(net3326),
    .A(net3395),
    .Y(_03821_),
    .D(net3312));
 sg13g2_a22oi_1 _09956_ (.Y(_03822_),
    .B1(net3311),
    .B2(net3395),
    .A2(net3325),
    .A1(net3391));
 sg13g2_or3_1 _09957_ (.A(_03819_),
    .B(_03820_),
    .C(_03822_),
    .X(_03823_));
 sg13g2_o21ai_1 _09958_ (.B1(_03819_),
    .Y(_03824_),
    .A1(_03820_),
    .A2(_03822_));
 sg13g2_nand3_1 _09959_ (.B(_03823_),
    .C(_03824_),
    .A(_03818_),
    .Y(_03825_));
 sg13g2_a21oi_1 _09960_ (.A1(_03823_),
    .A2(_03824_),
    .Y(_03826_),
    .B1(_03818_));
 sg13g2_a21o_1 _09961_ (.A2(_03824_),
    .A1(_03823_),
    .B1(_03818_),
    .X(_03827_));
 sg13g2_nand2_1 _09962_ (.Y(_03828_),
    .A(_03825_),
    .B(_03827_));
 sg13g2_xnor2_1 _09963_ (.Y(_03829_),
    .A(_03817_),
    .B(_03828_));
 sg13g2_nand2b_1 _09964_ (.Y(_03830_),
    .B(_03811_),
    .A_N(_03829_));
 sg13g2_xor2_1 _09965_ (.B(_03829_),
    .A(_03811_),
    .X(_03831_));
 sg13g2_xor2_1 _09966_ (.B(_03831_),
    .A(_03790_),
    .X(_03832_));
 sg13g2_and2_1 _09967_ (.A(_03804_),
    .B(_03832_),
    .X(_03833_));
 sg13g2_a21oi_1 _09968_ (.A1(_03783_),
    .A2(_03805_),
    .Y(_03834_),
    .B1(_03804_));
 sg13g2_nand3_1 _09969_ (.B(_03805_),
    .C(_03832_),
    .A(_03783_),
    .Y(_03835_));
 sg13g2_xor2_1 _09970_ (.B(_03834_),
    .A(_03832_),
    .X(_03836_));
 sg13g2_xnor2_1 _09971_ (.Y(_03837_),
    .A(_03807_),
    .B(_03836_));
 sg13g2_o21ai_1 _09972_ (.B1(_03810_),
    .Y(_00384_),
    .A1(net2745),
    .A2(_03837_));
 sg13g2_o21ai_1 _09973_ (.B1(_03835_),
    .Y(_03838_),
    .A1(_03807_),
    .A2(_03836_));
 sg13g2_o21ai_1 _09974_ (.B1(_03830_),
    .Y(_03839_),
    .A1(_03790_),
    .A2(_03831_));
 sg13g2_or2_1 _09975_ (.X(_03840_),
    .B(_03815_),
    .A(_03813_));
 sg13g2_nand2_1 _09976_ (.Y(_03841_),
    .A(net3402),
    .B(net3291));
 sg13g2_nand2b_1 _09977_ (.Y(_03842_),
    .B(_03840_),
    .A_N(_03841_));
 sg13g2_xnor2_1 _09978_ (.Y(_03843_),
    .A(_03840_),
    .B(_03841_));
 sg13g2_o21ai_1 _09979_ (.B1(_03825_),
    .Y(_03844_),
    .A1(_03817_),
    .A2(_03826_));
 sg13g2_nand2_1 _09980_ (.Y(_03845_),
    .A(net3398),
    .B(net3297));
 sg13g2_and2_1 _09981_ (.A(net3382),
    .B(net3351),
    .X(_03846_));
 sg13g2_nand2_1 _09982_ (.Y(_03847_),
    .A(net3382),
    .B(net3351));
 sg13g2_nand2_1 _09983_ (.Y(_03848_),
    .A(net3394),
    .B(net3305));
 sg13g2_xnor2_1 _09984_ (.Y(_03849_),
    .A(_03846_),
    .B(_03848_));
 sg13g2_nand2b_1 _09985_ (.Y(_03850_),
    .B(_03849_),
    .A_N(_03845_));
 sg13g2_xnor2_1 _09986_ (.Y(_03851_),
    .A(_03845_),
    .B(_03849_));
 sg13g2_o21ai_1 _09987_ (.B1(_03821_),
    .Y(_03852_),
    .A1(_03819_),
    .A2(_03822_));
 sg13g2_nand2_1 _09988_ (.Y(_03853_),
    .A(net3385),
    .B(net3336));
 sg13g2_and4_1 _09989_ (.A(net3391),
    .B(net3388),
    .C(net3325),
    .D(net3312),
    .X(_03854_));
 sg13g2_nand4_1 _09990_ (.B(net3388),
    .C(net3325),
    .A(net3392),
    .Y(_03855_),
    .D(net3317));
 sg13g2_a22oi_1 _09991_ (.Y(_03856_),
    .B1(net3312),
    .B2(net3391),
    .A2(net3325),
    .A1(net3388));
 sg13g2_or3_1 _09992_ (.A(_03853_),
    .B(_03854_),
    .C(_03856_),
    .X(_03857_));
 sg13g2_o21ai_1 _09993_ (.B1(_03853_),
    .Y(_03858_),
    .A1(_03854_),
    .A2(_03856_));
 sg13g2_nand3_1 _09994_ (.B(_03857_),
    .C(_03858_),
    .A(_03852_),
    .Y(_03859_));
 sg13g2_a21o_1 _09995_ (.A2(_03858_),
    .A1(_03857_),
    .B1(_03852_),
    .X(_03860_));
 sg13g2_nand3_1 _09996_ (.B(_03859_),
    .C(_03860_),
    .A(_03851_),
    .Y(_03861_));
 sg13g2_a21o_1 _09997_ (.A2(_03860_),
    .A1(_03859_),
    .B1(_03851_),
    .X(_03862_));
 sg13g2_nand3_1 _09998_ (.B(_03861_),
    .C(_03862_),
    .A(_03844_),
    .Y(_03863_));
 sg13g2_a21o_1 _09999_ (.A2(_03862_),
    .A1(_03861_),
    .B1(_03844_),
    .X(_03864_));
 sg13g2_a21oi_1 _10000_ (.A1(_03863_),
    .A2(_03864_),
    .Y(_03865_),
    .B1(_03843_));
 sg13g2_nand3_1 _10001_ (.B(_03863_),
    .C(_03864_),
    .A(_03843_),
    .Y(_03866_));
 sg13g2_nor2b_1 _10002_ (.A(_03865_),
    .B_N(_03866_),
    .Y(_03867_));
 sg13g2_nand2_1 _10003_ (.Y(_03868_),
    .A(_03839_),
    .B(_03867_));
 sg13g2_xor2_1 _10004_ (.B(_03867_),
    .A(_03839_),
    .X(_03869_));
 sg13g2_and2_1 _10005_ (.A(_03833_),
    .B(_03869_),
    .X(_03870_));
 sg13g2_xor2_1 _10006_ (.B(_03869_),
    .A(_03833_),
    .X(_03871_));
 sg13g2_a21oi_1 _10007_ (.A1(_03838_),
    .A2(_03871_),
    .Y(_03872_),
    .B1(net2745));
 sg13g2_o21ai_1 _10008_ (.B1(_03872_),
    .Y(_03873_),
    .A1(_03838_),
    .A2(_03871_));
 sg13g2_o21ai_1 _10009_ (.B1(_03873_),
    .Y(_00385_),
    .A1(_01175_),
    .A2(_03753_));
 sg13g2_a21o_1 _10010_ (.A2(_03871_),
    .A1(_03838_),
    .B1(_03870_),
    .X(_03874_));
 sg13g2_nand2_1 _10011_ (.Y(_03875_),
    .A(_03863_),
    .B(_03866_));
 sg13g2_o21ai_1 _10012_ (.B1(_03850_),
    .Y(_03876_),
    .A1(_03847_),
    .A2(_03848_));
 sg13g2_nor2_1 _10013_ (.A(net3402),
    .B(net3282),
    .Y(_03877_));
 sg13g2_nand2_2 _10014_ (.Y(_03878_),
    .A(net3394),
    .B(net3291));
 sg13g2_nor2_1 _10015_ (.A(_03845_),
    .B(_03878_),
    .Y(_03879_));
 sg13g2_a22oi_1 _10016_ (.Y(_03880_),
    .B1(net3292),
    .B2(net3398),
    .A2(net3298),
    .A1(net3394));
 sg13g2_nor2_1 _10017_ (.A(_03879_),
    .B(_03880_),
    .Y(_03881_));
 sg13g2_xor2_1 _10018_ (.B(_03881_),
    .A(_03877_),
    .X(_03882_));
 sg13g2_nand2_1 _10019_ (.Y(_03883_),
    .A(_03876_),
    .B(_03882_));
 sg13g2_xnor2_1 _10020_ (.Y(_03884_),
    .A(_03876_),
    .B(_03882_));
 sg13g2_nand2_1 _10021_ (.Y(_03885_),
    .A(_03859_),
    .B(_03861_));
 sg13g2_nand2_1 _10022_ (.Y(_03886_),
    .A(net3391),
    .B(net3305));
 sg13g2_and2_1 _10023_ (.A(net3376),
    .B(net3343),
    .X(_03887_));
 sg13g2_nand2_2 _10024_ (.Y(_03888_),
    .A(net3378),
    .B(net3344));
 sg13g2_nand2_1 _10025_ (.Y(_03889_),
    .A(_03846_),
    .B(_03887_));
 sg13g2_a22oi_1 _10026_ (.Y(_03890_),
    .B1(net3343),
    .B2(net3382),
    .A2(net3351),
    .A1(net3376));
 sg13g2_a21oi_1 _10027_ (.A1(_03846_),
    .A2(_03887_),
    .Y(_03891_),
    .B1(_03890_));
 sg13g2_xor2_1 _10028_ (.B(_03891_),
    .A(_03886_),
    .X(_03892_));
 sg13g2_o21ai_1 _10029_ (.B1(_03855_),
    .Y(_03893_),
    .A1(_03853_),
    .A2(_03856_));
 sg13g2_nand2_1 _10030_ (.Y(_03894_),
    .A(net3385),
    .B(net3330));
 sg13g2_and3_1 _10031_ (.X(_03895_),
    .A(net3388),
    .B(net3317),
    .C(net3285));
 sg13g2_nand3_1 _10032_ (.B(net3317),
    .C(net3285),
    .A(net3388),
    .Y(_03896_));
 sg13g2_a21oi_1 _10033_ (.A1(net3388),
    .A2(net3317),
    .Y(_03897_),
    .B1(net3285));
 sg13g2_or3_1 _10034_ (.A(_03894_),
    .B(_03895_),
    .C(_03897_),
    .X(_03898_));
 sg13g2_o21ai_1 _10035_ (.B1(_03894_),
    .Y(_03899_),
    .A1(_03895_),
    .A2(_03897_));
 sg13g2_nand3_1 _10036_ (.B(_03898_),
    .C(_03899_),
    .A(_03893_),
    .Y(_03900_));
 sg13g2_a21oi_1 _10037_ (.A1(_03898_),
    .A2(_03899_),
    .Y(_03901_),
    .B1(_03893_));
 sg13g2_a21o_1 _10038_ (.A2(_03899_),
    .A1(_03898_),
    .B1(_03893_),
    .X(_03902_));
 sg13g2_nand2_1 _10039_ (.Y(_03903_),
    .A(_03900_),
    .B(_03902_));
 sg13g2_xnor2_1 _10040_ (.Y(_03904_),
    .A(_03892_),
    .B(_03903_));
 sg13g2_nand2b_1 _10041_ (.Y(_03905_),
    .B(_03885_),
    .A_N(_03904_));
 sg13g2_nor2b_1 _10042_ (.A(_03885_),
    .B_N(_03904_),
    .Y(_03906_));
 sg13g2_xnor2_1 _10043_ (.Y(_03907_),
    .A(_03885_),
    .B(_03904_));
 sg13g2_xnor2_1 _10044_ (.Y(_03908_),
    .A(_03884_),
    .B(_03907_));
 sg13g2_nand2_1 _10045_ (.Y(_03909_),
    .A(_03875_),
    .B(_03908_));
 sg13g2_xnor2_1 _10046_ (.Y(_03910_),
    .A(_03875_),
    .B(_03908_));
 sg13g2_xor2_1 _10047_ (.B(_03910_),
    .A(_03842_),
    .X(_03911_));
 sg13g2_nor2b_1 _10048_ (.A(_03868_),
    .B_N(_03911_),
    .Y(_03912_));
 sg13g2_xnor2_1 _10049_ (.Y(_03913_),
    .A(_03868_),
    .B(_03911_));
 sg13g2_nor2_1 _10050_ (.A(_03874_),
    .B(_03913_),
    .Y(_03914_));
 sg13g2_a21oi_1 _10051_ (.A1(_03874_),
    .A2(_03913_),
    .Y(_03915_),
    .B1(net2745));
 sg13g2_nor2b_1 _10052_ (.A(_03914_),
    .B_N(_03915_),
    .Y(_03916_));
 sg13g2_a21o_1 _10053_ (.A2(net2814),
    .A1(net962),
    .B1(_03916_),
    .X(_00386_));
 sg13g2_nand2_1 _10054_ (.Y(_03917_),
    .A(net890),
    .B(net2814));
 sg13g2_o21ai_1 _10055_ (.B1(_03905_),
    .Y(_03918_),
    .A1(_03884_),
    .A2(_03906_));
 sg13g2_a21oi_2 _10056_ (.B1(_03879_),
    .Y(_03919_),
    .A2(_03881_),
    .A1(_03877_));
 sg13g2_o21ai_1 _10057_ (.B1(_03889_),
    .Y(_03920_),
    .A1(_03886_),
    .A2(_03890_));
 sg13g2_nor2_1 _10058_ (.A(net3398),
    .B(net3282),
    .Y(_03921_));
 sg13g2_nor3_1 _10059_ (.A(net3398),
    .B(net3282),
    .C(_03878_),
    .Y(_03922_));
 sg13g2_inv_1 _10060_ (.Y(_03923_),
    .A(_03922_));
 sg13g2_xnor2_1 _10061_ (.Y(_03924_),
    .A(_03878_),
    .B(_03921_));
 sg13g2_xnor2_1 _10062_ (.Y(_03925_),
    .A(_03920_),
    .B(_03924_));
 sg13g2_nor2_1 _10063_ (.A(_03919_),
    .B(_03925_),
    .Y(_03926_));
 sg13g2_xnor2_1 _10064_ (.Y(_03927_),
    .A(_03919_),
    .B(_03925_));
 sg13g2_o21ai_1 _10065_ (.B1(_03900_),
    .Y(_03928_),
    .A1(_03892_),
    .A2(_03901_));
 sg13g2_nand2_1 _10066_ (.Y(_03929_),
    .A(net3392),
    .B(net3298));
 sg13g2_and3_1 _10067_ (.X(_03930_),
    .A(net3377),
    .B(net3352),
    .C(net3305));
 sg13g2_nand2_1 _10068_ (.Y(_03931_),
    .A(net3389),
    .B(net3278));
 sg13g2_a22oi_1 _10069_ (.Y(_03932_),
    .B1(net3305),
    .B2(net3389),
    .A2(net3352),
    .A1(net3377));
 sg13g2_a21oi_1 _10070_ (.A1(net3389),
    .A2(net3278),
    .Y(_03933_),
    .B1(_03932_));
 sg13g2_xor2_1 _10071_ (.B(_03933_),
    .A(_03929_),
    .X(_03934_));
 sg13g2_o21ai_1 _10072_ (.B1(_03896_),
    .Y(_03935_),
    .A1(_03894_),
    .A2(_03897_));
 sg13g2_and4_1 _10073_ (.A(net3385),
    .B(net3382),
    .C(net3330),
    .D(net3318),
    .X(_03936_));
 sg13g2_nand4_1 _10074_ (.B(net3382),
    .C(net3329),
    .A(net3384),
    .Y(_03937_),
    .D(net3318));
 sg13g2_a22oi_1 _10075_ (.Y(_03938_),
    .B1(net3317),
    .B2(net3384),
    .A2(net3329),
    .A1(net3382));
 sg13g2_nand3b_1 _10076_ (.B(_03887_),
    .C(_03937_),
    .Y(_03939_),
    .A_N(_03938_));
 sg13g2_o21ai_1 _10077_ (.B1(_03888_),
    .Y(_03940_),
    .A1(_03936_),
    .A2(_03938_));
 sg13g2_and3_1 _10078_ (.X(_03941_),
    .A(_03935_),
    .B(_03939_),
    .C(_03940_));
 sg13g2_nand3_1 _10079_ (.B(_03939_),
    .C(_03940_),
    .A(_03935_),
    .Y(_03942_));
 sg13g2_a21oi_1 _10080_ (.A1(_03939_),
    .A2(_03940_),
    .Y(_03943_),
    .B1(_03935_));
 sg13g2_or3_1 _10081_ (.A(_03934_),
    .B(_03941_),
    .C(_03943_),
    .X(_03944_));
 sg13g2_o21ai_1 _10082_ (.B1(_03934_),
    .Y(_03945_),
    .A1(_03941_),
    .A2(_03943_));
 sg13g2_and3_1 _10083_ (.X(_03946_),
    .A(_03928_),
    .B(_03944_),
    .C(_03945_));
 sg13g2_nand3_1 _10084_ (.B(_03944_),
    .C(_03945_),
    .A(_03928_),
    .Y(_03947_));
 sg13g2_a21oi_1 _10085_ (.A1(_03944_),
    .A2(_03945_),
    .Y(_03948_),
    .B1(_03928_));
 sg13g2_nor2_1 _10086_ (.A(_03946_),
    .B(_03948_),
    .Y(_03949_));
 sg13g2_xnor2_1 _10087_ (.Y(_03950_),
    .A(_03927_),
    .B(_03949_));
 sg13g2_nand2_1 _10088_ (.Y(_03951_),
    .A(_03918_),
    .B(_03950_));
 sg13g2_xnor2_1 _10089_ (.Y(_03952_),
    .A(_03918_),
    .B(_03950_));
 sg13g2_xnor2_1 _10090_ (.Y(_03953_),
    .A(_03883_),
    .B(_03952_));
 sg13g2_o21ai_1 _10091_ (.B1(_03909_),
    .Y(_03954_),
    .A1(_03842_),
    .A2(_03910_));
 sg13g2_nor2b_1 _10092_ (.A(_03953_),
    .B_N(_03954_),
    .Y(_03955_));
 sg13g2_xor2_1 _10093_ (.B(_03954_),
    .A(_03953_),
    .X(_03956_));
 sg13g2_a21oi_2 _10094_ (.B1(_03912_),
    .Y(_03957_),
    .A2(_03913_),
    .A1(_03874_));
 sg13g2_nor2_1 _10095_ (.A(_03956_),
    .B(_03957_),
    .Y(_03958_));
 sg13g2_a21o_1 _10096_ (.A2(_03957_),
    .A1(_03956_),
    .B1(net2746),
    .X(_03959_));
 sg13g2_o21ai_1 _10097_ (.B1(_03917_),
    .Y(_00387_),
    .A1(_03958_),
    .A2(_03959_));
 sg13g2_o21ai_1 _10098_ (.B1(_03951_),
    .Y(_03960_),
    .A1(_03883_),
    .A2(_03952_));
 sg13g2_a21oi_1 _10099_ (.A1(_03920_),
    .A2(_03924_),
    .Y(_03961_),
    .B1(_03926_));
 sg13g2_o21ai_1 _10100_ (.B1(_03947_),
    .Y(_03962_),
    .A1(_03927_),
    .A2(_03948_));
 sg13g2_o21ai_1 _10101_ (.B1(_03931_),
    .Y(_03963_),
    .A1(_03929_),
    .A2(_03932_));
 sg13g2_nand2_1 _10102_ (.Y(_03964_),
    .A(net3392),
    .B(net3291));
 sg13g2_nor2_1 _10103_ (.A(net3395),
    .B(net3282),
    .Y(_03965_));
 sg13g2_nand2b_1 _10104_ (.Y(_03966_),
    .B(_03965_),
    .A_N(_03964_));
 sg13g2_xnor2_1 _10105_ (.Y(_03967_),
    .A(_03964_),
    .B(_03965_));
 sg13g2_nand2_1 _10106_ (.Y(_03968_),
    .A(_03963_),
    .B(_03967_));
 sg13g2_xnor2_1 _10107_ (.Y(_03969_),
    .A(_03963_),
    .B(_03967_));
 sg13g2_xnor2_1 _10108_ (.Y(_03970_),
    .A(_03923_),
    .B(_03969_));
 sg13g2_o21ai_1 _10109_ (.B1(_03942_),
    .Y(_03971_),
    .A1(_03934_),
    .A2(_03943_));
 sg13g2_nand2_1 _10110_ (.Y(_03972_),
    .A(net3389),
    .B(net3297));
 sg13g2_nand2_1 _10111_ (.Y(_03973_),
    .A(net3384),
    .B(net3278));
 sg13g2_a22oi_1 _10112_ (.Y(_03974_),
    .B1(net3305),
    .B2(net3384),
    .A2(net3352),
    .A1(net3378));
 sg13g2_a21oi_1 _10113_ (.A1(net3384),
    .A2(net3278),
    .Y(_03975_),
    .B1(_03974_));
 sg13g2_xor2_1 _10114_ (.B(_03975_),
    .A(_03972_),
    .X(_03976_));
 sg13g2_o21ai_1 _10115_ (.B1(_03937_),
    .Y(_03977_),
    .A1(_03888_),
    .A2(_03938_));
 sg13g2_and4_1 _10116_ (.A(net3382),
    .B(net3377),
    .C(net3330),
    .D(net3317),
    .X(_03978_));
 sg13g2_nand4_1 _10117_ (.B(net3377),
    .C(net3329),
    .A(net3380),
    .Y(_03979_),
    .D(net3317));
 sg13g2_a22oi_1 _10118_ (.Y(_03980_),
    .B1(net3317),
    .B2(net3380),
    .A2(net3329),
    .A1(net3377));
 sg13g2_nand3b_1 _10119_ (.B(_03887_),
    .C(_03979_),
    .Y(_03981_),
    .A_N(_03980_));
 sg13g2_o21ai_1 _10120_ (.B1(_03888_),
    .Y(_03982_),
    .A1(_03978_),
    .A2(_03980_));
 sg13g2_and3_1 _10121_ (.X(_03983_),
    .A(_03977_),
    .B(_03981_),
    .C(_03982_));
 sg13g2_nand3_1 _10122_ (.B(_03981_),
    .C(_03982_),
    .A(_03977_),
    .Y(_03984_));
 sg13g2_a21oi_1 _10123_ (.A1(_03981_),
    .A2(_03982_),
    .Y(_03985_),
    .B1(_03977_));
 sg13g2_or3_1 _10124_ (.A(_03976_),
    .B(_03983_),
    .C(_03985_),
    .X(_03986_));
 sg13g2_o21ai_1 _10125_ (.B1(_03976_),
    .Y(_03987_),
    .A1(_03983_),
    .A2(_03985_));
 sg13g2_and3_1 _10126_ (.X(_03988_),
    .A(_03971_),
    .B(_03986_),
    .C(_03987_));
 sg13g2_nand3_1 _10127_ (.B(_03986_),
    .C(_03987_),
    .A(_03971_),
    .Y(_03989_));
 sg13g2_a21oi_1 _10128_ (.A1(_03986_),
    .A2(_03987_),
    .Y(_03990_),
    .B1(_03971_));
 sg13g2_or3_1 _10129_ (.A(_03970_),
    .B(_03988_),
    .C(_03990_),
    .X(_03991_));
 sg13g2_o21ai_1 _10130_ (.B1(_03970_),
    .Y(_03992_),
    .A1(_03988_),
    .A2(_03990_));
 sg13g2_nand3_1 _10131_ (.B(_03991_),
    .C(_03992_),
    .A(_03962_),
    .Y(_03993_));
 sg13g2_a21oi_1 _10132_ (.A1(_03991_),
    .A2(_03992_),
    .Y(_03994_),
    .B1(_03962_));
 sg13g2_a21o_1 _10133_ (.A2(_03992_),
    .A1(_03991_),
    .B1(_03962_),
    .X(_03995_));
 sg13g2_nand2_1 _10134_ (.Y(_03996_),
    .A(_03993_),
    .B(_03995_));
 sg13g2_xnor2_1 _10135_ (.Y(_03997_),
    .A(_03961_),
    .B(_03996_));
 sg13g2_nor2b_1 _10136_ (.A(_03997_),
    .B_N(_03960_),
    .Y(_03998_));
 sg13g2_nand2b_1 _10137_ (.Y(_03999_),
    .B(_03997_),
    .A_N(_03960_));
 sg13g2_nand2b_1 _10138_ (.Y(_04000_),
    .B(_03999_),
    .A_N(_03998_));
 sg13g2_nor2_1 _10139_ (.A(_03955_),
    .B(_03958_),
    .Y(_04001_));
 sg13g2_a21oi_1 _10140_ (.A1(_04000_),
    .A2(_04001_),
    .Y(_04002_),
    .B1(net2745));
 sg13g2_o21ai_1 _10141_ (.B1(_04002_),
    .Y(_04003_),
    .A1(_04000_),
    .A2(_04001_));
 sg13g2_o21ai_1 _10142_ (.B1(_04003_),
    .Y(_00388_),
    .A1(_01177_),
    .A2(_03753_));
 sg13g2_nand2_1 _10143_ (.Y(_04004_),
    .A(net856),
    .B(net2815));
 sg13g2_o21ai_1 _10144_ (.B1(_03968_),
    .Y(_04005_),
    .A1(_03923_),
    .A2(_03969_));
 sg13g2_inv_1 _10145_ (.Y(_04006_),
    .A(_04005_));
 sg13g2_o21ai_1 _10146_ (.B1(_03989_),
    .Y(_04007_),
    .A1(_03970_),
    .A2(_03990_));
 sg13g2_o21ai_1 _10147_ (.B1(_03973_),
    .Y(_04008_),
    .A1(_03972_),
    .A2(_03974_));
 sg13g2_nand2_1 _10148_ (.Y(_04009_),
    .A(net3389),
    .B(net3291));
 sg13g2_nor2_1 _10149_ (.A(net3392),
    .B(net3283),
    .Y(_04010_));
 sg13g2_nand2b_1 _10150_ (.Y(_04011_),
    .B(_04010_),
    .A_N(_04009_));
 sg13g2_xnor2_1 _10151_ (.Y(_04012_),
    .A(_04009_),
    .B(_04010_));
 sg13g2_nand2_1 _10152_ (.Y(_04013_),
    .A(_04008_),
    .B(_04012_));
 sg13g2_xnor2_1 _10153_ (.Y(_04014_),
    .A(_04008_),
    .B(_04012_));
 sg13g2_xnor2_1 _10154_ (.Y(_04015_),
    .A(_03966_),
    .B(_04014_));
 sg13g2_o21ai_1 _10155_ (.B1(_03984_),
    .Y(_04016_),
    .A1(_03976_),
    .A2(_03985_));
 sg13g2_and2_1 _10156_ (.A(net3385),
    .B(net3298),
    .X(_04017_));
 sg13g2_a22oi_1 _10157_ (.Y(_04018_),
    .B1(net3305),
    .B2(net3380),
    .A2(net3352),
    .A1(net3377));
 sg13g2_a21oi_1 _10158_ (.A1(net3381),
    .A2(net3278),
    .Y(_04019_),
    .B1(_04018_));
 sg13g2_xor2_1 _10159_ (.B(_04019_),
    .A(_04017_),
    .X(_04020_));
 sg13g2_o21ai_1 _10160_ (.B1(_03979_),
    .Y(_04021_),
    .A1(_03888_),
    .A2(_03980_));
 sg13g2_nand2b_1 _10161_ (.Y(_04022_),
    .B(net3376),
    .A_N(net3344));
 sg13g2_mux2_1 _10162_ (.A0(_03888_),
    .A1(_04022_),
    .S(_01661_),
    .X(_04023_));
 sg13g2_and4_2 _10163_ (.A(net3377),
    .B(net3343),
    .C(net3330),
    .D(net3319),
    .X(_04024_));
 sg13g2_nand4_1 _10164_ (.B(net3344),
    .C(net3333),
    .A(net3378),
    .Y(_04025_),
    .D(net3319));
 sg13g2_xnor2_1 _10165_ (.Y(_04026_),
    .A(_04021_),
    .B(_04023_));
 sg13g2_xnor2_1 _10166_ (.Y(_04027_),
    .A(_04020_),
    .B(_04026_));
 sg13g2_nand2b_1 _10167_ (.Y(_04028_),
    .B(_04016_),
    .A_N(_04027_));
 sg13g2_xor2_1 _10168_ (.B(_04027_),
    .A(_04016_),
    .X(_04029_));
 sg13g2_xor2_1 _10169_ (.B(_04029_),
    .A(_04015_),
    .X(_04030_));
 sg13g2_nand2_1 _10170_ (.Y(_04031_),
    .A(_04007_),
    .B(_04030_));
 sg13g2_xnor2_1 _10171_ (.Y(_04032_),
    .A(_04007_),
    .B(_04030_));
 sg13g2_xnor2_1 _10172_ (.Y(_04033_),
    .A(_04006_),
    .B(_04032_));
 sg13g2_o21ai_1 _10173_ (.B1(_03993_),
    .Y(_04034_),
    .A1(_03961_),
    .A2(_03994_));
 sg13g2_nor2b_1 _10174_ (.A(_04033_),
    .B_N(_04034_),
    .Y(_04035_));
 sg13g2_xor2_1 _10175_ (.B(_04034_),
    .A(_04033_),
    .X(_04036_));
 sg13g2_nor3_1 _10176_ (.A(_03956_),
    .B(_03957_),
    .C(_04000_),
    .Y(_04037_));
 sg13g2_a21o_1 _10177_ (.A2(_03999_),
    .A1(_03955_),
    .B1(_03998_),
    .X(_04038_));
 sg13g2_nor2_1 _10178_ (.A(_04037_),
    .B(_04038_),
    .Y(_04039_));
 sg13g2_nor2_1 _10179_ (.A(_04036_),
    .B(_04039_),
    .Y(_04040_));
 sg13g2_a21o_1 _10180_ (.A2(_04039_),
    .A1(_04036_),
    .B1(net2746),
    .X(_04041_));
 sg13g2_o21ai_1 _10181_ (.B1(_04004_),
    .Y(_00389_),
    .A1(_04040_),
    .A2(_04041_));
 sg13g2_nand2_1 _10182_ (.Y(_04042_),
    .A(net951),
    .B(net2814));
 sg13g2_o21ai_1 _10183_ (.B1(_04031_),
    .Y(_04043_),
    .A1(_04006_),
    .A2(_04032_));
 sg13g2_o21ai_1 _10184_ (.B1(_04013_),
    .Y(_04044_),
    .A1(_03966_),
    .A2(_04014_));
 sg13g2_o21ai_1 _10185_ (.B1(_04028_),
    .Y(_04045_),
    .A1(_04015_),
    .A2(_04029_));
 sg13g2_a22oi_1 _10186_ (.Y(_04046_),
    .B1(_04017_),
    .B2(_04019_),
    .A2(net3278),
    .A1(net3380));
 sg13g2_nand2_1 _10187_ (.Y(_04047_),
    .A(net3384),
    .B(net3291));
 sg13g2_nor2_1 _10188_ (.A(net3389),
    .B(net3282),
    .Y(_04048_));
 sg13g2_nand2b_1 _10189_ (.Y(_04049_),
    .B(_04048_),
    .A_N(_04047_));
 sg13g2_xnor2_1 _10190_ (.Y(_04050_),
    .A(_04047_),
    .B(_04048_));
 sg13g2_nand2b_1 _10191_ (.Y(_04051_),
    .B(_04050_),
    .A_N(_04046_));
 sg13g2_xor2_1 _10192_ (.B(_04050_),
    .A(_04046_),
    .X(_04052_));
 sg13g2_xnor2_1 _10193_ (.Y(_04053_),
    .A(_04011_),
    .B(_04052_));
 sg13g2_a21oi_2 _10194_ (.B1(_04024_),
    .Y(_04054_),
    .A2(_04026_),
    .A1(_04020_));
 sg13g2_o21ai_1 _10195_ (.B1(net3379),
    .Y(_04055_),
    .A1(net3355),
    .A2(net3306));
 sg13g2_nor2_1 _10196_ (.A(_03930_),
    .B(_04055_),
    .Y(_04056_));
 sg13g2_nand2_1 _10197_ (.Y(_04057_),
    .A(net3380),
    .B(net3297));
 sg13g2_and2_1 _10198_ (.A(net3297),
    .B(_04056_),
    .X(_04058_));
 sg13g2_xor2_1 _10199_ (.B(_04057_),
    .A(_04056_),
    .X(_04059_));
 sg13g2_o21ai_1 _10200_ (.B1(net3377),
    .Y(_04060_),
    .A1(net3330),
    .A2(net3319));
 sg13g2_a21oi_1 _10201_ (.A1(_03888_),
    .A2(_04060_),
    .Y(_04061_),
    .B1(_04024_));
 sg13g2_inv_1 _10202_ (.Y(_04062_),
    .A(_04061_));
 sg13g2_xnor2_1 _10203_ (.Y(_04063_),
    .A(_04059_),
    .B(_04061_));
 sg13g2_nand2b_1 _10204_ (.Y(_04064_),
    .B(_04063_),
    .A_N(_04054_));
 sg13g2_xnor2_1 _10205_ (.Y(_04065_),
    .A(_04054_),
    .B(_04063_));
 sg13g2_inv_1 _10206_ (.Y(_04066_),
    .A(_04065_));
 sg13g2_xnor2_1 _10207_ (.Y(_04067_),
    .A(_04053_),
    .B(_04065_));
 sg13g2_xnor2_1 _10208_ (.Y(_04068_),
    .A(_04045_),
    .B(_04067_));
 sg13g2_nor2b_1 _10209_ (.A(_04068_),
    .B_N(_04044_),
    .Y(_04069_));
 sg13g2_xnor2_1 _10210_ (.Y(_04070_),
    .A(_04044_),
    .B(_04068_));
 sg13g2_nor2_1 _10211_ (.A(_04043_),
    .B(_04070_),
    .Y(_04071_));
 sg13g2_xor2_1 _10212_ (.B(_04070_),
    .A(_04043_),
    .X(_04072_));
 sg13g2_nor3_1 _10213_ (.A(_04035_),
    .B(_04040_),
    .C(_04072_),
    .Y(_04073_));
 sg13g2_o21ai_1 _10214_ (.B1(_04072_),
    .Y(_04074_),
    .A1(_04035_),
    .A2(_04040_));
 sg13g2_nand2b_1 _10215_ (.Y(_04075_),
    .B(_04074_),
    .A_N(net2746));
 sg13g2_o21ai_1 _10216_ (.B1(_04042_),
    .Y(_00390_),
    .A1(_04073_),
    .A2(_04075_));
 sg13g2_o21ai_1 _10217_ (.B1(_04051_),
    .Y(_04076_),
    .A1(_04011_),
    .A2(_04052_));
 sg13g2_o21ai_1 _10218_ (.B1(_04064_),
    .Y(_04077_),
    .A1(_04053_),
    .A2(_04066_));
 sg13g2_o21ai_1 _10219_ (.B1(_04025_),
    .Y(_04078_),
    .A1(_04059_),
    .A2(_04062_));
 sg13g2_a21oi_1 _10220_ (.A1(net3378),
    .A2(net3297),
    .Y(_04079_),
    .B1(_04056_));
 sg13g2_or2_1 _10221_ (.X(_04080_),
    .B(_04079_),
    .A(_04058_));
 sg13g2_xnor2_1 _10222_ (.Y(_04081_),
    .A(_04062_),
    .B(_04080_));
 sg13g2_inv_1 _10223_ (.Y(_04082_),
    .A(_04081_));
 sg13g2_xor2_1 _10224_ (.B(_04081_),
    .A(_04078_),
    .X(_04083_));
 sg13g2_a21oi_1 _10225_ (.A1(net3380),
    .A2(_04058_),
    .Y(_04084_),
    .B1(net3278));
 sg13g2_nand2_1 _10226_ (.Y(_04085_),
    .A(net3380),
    .B(net3291));
 sg13g2_nor2_1 _10227_ (.A(net3384),
    .B(net3282),
    .Y(_04086_));
 sg13g2_nor3_1 _10228_ (.A(net3384),
    .B(net3283),
    .C(_04085_),
    .Y(_04087_));
 sg13g2_xnor2_1 _10229_ (.Y(_04088_),
    .A(_04085_),
    .B(_04086_));
 sg13g2_nand2b_1 _10230_ (.Y(_04089_),
    .B(_04088_),
    .A_N(_04084_));
 sg13g2_xor2_1 _10231_ (.B(_04088_),
    .A(_04084_),
    .X(_04090_));
 sg13g2_xnor2_1 _10232_ (.Y(_04091_),
    .A(_04049_),
    .B(_04090_));
 sg13g2_nor2_1 _10233_ (.A(_04083_),
    .B(_04091_),
    .Y(_04092_));
 sg13g2_xor2_1 _10234_ (.B(_04091_),
    .A(_04083_),
    .X(_04093_));
 sg13g2_xnor2_1 _10235_ (.Y(_04094_),
    .A(_04077_),
    .B(_04093_));
 sg13g2_nor2b_1 _10236_ (.A(_04094_),
    .B_N(_04076_),
    .Y(_04095_));
 sg13g2_xor2_1 _10237_ (.B(_04094_),
    .A(_04076_),
    .X(_04096_));
 sg13g2_a21o_1 _10238_ (.A2(_04067_),
    .A1(_04045_),
    .B1(_04069_),
    .X(_04097_));
 sg13g2_nor2b_1 _10239_ (.A(_04096_),
    .B_N(_04097_),
    .Y(_04098_));
 sg13g2_xor2_1 _10240_ (.B(_04097_),
    .A(_04096_),
    .X(_04099_));
 sg13g2_nor2b_1 _10241_ (.A(_04036_),
    .B_N(_04072_),
    .Y(_04100_));
 sg13g2_inv_1 _10242_ (.Y(_04101_),
    .A(_04100_));
 sg13g2_nor2b_1 _10243_ (.A(_04071_),
    .B_N(_04035_),
    .Y(_04102_));
 sg13g2_a221oi_1 _10244_ (.B2(_04038_),
    .C1(_04102_),
    .B1(_04100_),
    .A1(_04043_),
    .Y(_04103_),
    .A2(_04070_));
 sg13g2_or4_1 _10245_ (.A(_03956_),
    .B(_03957_),
    .C(_04000_),
    .D(_04101_),
    .X(_04104_));
 sg13g2_and3_1 _10246_ (.X(_04105_),
    .A(_04099_),
    .B(_04103_),
    .C(_04104_));
 sg13g2_a21oi_1 _10247_ (.A1(_04103_),
    .A2(_04104_),
    .Y(_04106_),
    .B1(_04099_));
 sg13g2_nor3_1 _10248_ (.A(net2747),
    .B(_04105_),
    .C(_04106_),
    .Y(_04107_));
 sg13g2_a21oi_1 _10249_ (.A1(net989),
    .A2(net2815),
    .Y(_04108_),
    .B1(_04107_));
 sg13g2_inv_1 _10250_ (.Y(_00391_),
    .A(_04108_));
 sg13g2_o21ai_1 _10251_ (.B1(_04089_),
    .Y(_04109_),
    .A1(_04049_),
    .A2(_04090_));
 sg13g2_a21oi_1 _10252_ (.A1(_04078_),
    .A2(_04082_),
    .Y(_04110_),
    .B1(_04092_));
 sg13g2_nand2_1 _10253_ (.Y(_04111_),
    .A(_04024_),
    .B(_04082_));
 sg13g2_nand3_1 _10254_ (.B(_04062_),
    .C(_04080_),
    .A(_04025_),
    .Y(_04112_));
 sg13g2_and2_1 _10255_ (.A(_04111_),
    .B(_04112_),
    .X(_04113_));
 sg13g2_inv_1 _10256_ (.Y(_04114_),
    .A(_04113_));
 sg13g2_nor2_2 _10257_ (.A(net3278),
    .B(_04058_),
    .Y(_04115_));
 sg13g2_nand2_2 _10258_ (.Y(_04116_),
    .A(net3378),
    .B(net3291));
 sg13g2_nor2_1 _10259_ (.A(net3380),
    .B(net3282),
    .Y(_04117_));
 sg13g2_nor3_2 _10260_ (.A(net3381),
    .B(net3282),
    .C(_04116_),
    .Y(_04118_));
 sg13g2_xnor2_1 _10261_ (.Y(_04119_),
    .A(_04116_),
    .B(_04117_));
 sg13g2_o21ai_1 _10262_ (.B1(_04119_),
    .Y(_04120_),
    .A1(_03930_),
    .A2(_04058_));
 sg13g2_xor2_1 _10263_ (.B(_04119_),
    .A(_04115_),
    .X(_04121_));
 sg13g2_inv_1 _10264_ (.Y(_04122_),
    .A(_04121_));
 sg13g2_nand2_1 _10265_ (.Y(_04123_),
    .A(_04087_),
    .B(_04122_));
 sg13g2_xor2_1 _10266_ (.B(_04121_),
    .A(_04087_),
    .X(_04124_));
 sg13g2_xor2_1 _10267_ (.B(_04124_),
    .A(_04113_),
    .X(_04125_));
 sg13g2_nor2_1 _10268_ (.A(_04110_),
    .B(_04125_),
    .Y(_04126_));
 sg13g2_xor2_1 _10269_ (.B(_04125_),
    .A(_04110_),
    .X(_04127_));
 sg13g2_xnor2_1 _10270_ (.Y(_04128_),
    .A(_04109_),
    .B(_04127_));
 sg13g2_a21oi_1 _10271_ (.A1(_04077_),
    .A2(_04093_),
    .Y(_04129_),
    .B1(_04095_));
 sg13g2_nor2_1 _10272_ (.A(_04128_),
    .B(_04129_),
    .Y(_04130_));
 sg13g2_xor2_1 _10273_ (.B(_04129_),
    .A(_04128_),
    .X(_04131_));
 sg13g2_nor3_1 _10274_ (.A(_04098_),
    .B(_04106_),
    .C(_04131_),
    .Y(_04132_));
 sg13g2_and2_1 _10275_ (.A(_04106_),
    .B(_04131_),
    .X(_04133_));
 sg13g2_and2_1 _10276_ (.A(_04098_),
    .B(_04131_),
    .X(_04134_));
 sg13g2_nor4_1 _10277_ (.A(net2747),
    .B(_04132_),
    .C(_04133_),
    .D(_04134_),
    .Y(_04135_));
 sg13g2_a21o_1 _10278_ (.A2(net2815),
    .A1(net1007),
    .B1(_04135_),
    .X(_00392_));
 sg13g2_and2_1 _10279_ (.A(net1082),
    .B(net2815),
    .X(_04136_));
 sg13g2_or3_1 _10280_ (.A(_04130_),
    .B(_04133_),
    .C(_04134_),
    .X(_04137_));
 sg13g2_nand2_1 _10281_ (.Y(_04138_),
    .A(_04120_),
    .B(_04123_));
 sg13g2_o21ai_1 _10282_ (.B1(_04111_),
    .Y(_04139_),
    .A1(_04114_),
    .A2(_04124_));
 sg13g2_o21ai_1 _10283_ (.B1(_04116_),
    .Y(_04140_),
    .A1(net3378),
    .A2(net3283));
 sg13g2_nor2b_1 _10284_ (.A(_04115_),
    .B_N(_04140_),
    .Y(_04141_));
 sg13g2_xor2_1 _10285_ (.B(_04140_),
    .A(_04115_),
    .X(_04142_));
 sg13g2_mux2_1 _10286_ (.A0(_04142_),
    .A1(_04115_),
    .S(_04118_),
    .X(_04143_));
 sg13g2_xnor2_1 _10287_ (.Y(_04144_),
    .A(_04113_),
    .B(_04143_));
 sg13g2_xnor2_1 _10288_ (.Y(_04145_),
    .A(_04139_),
    .B(_04144_));
 sg13g2_nor2b_1 _10289_ (.A(_04145_),
    .B_N(_04138_),
    .Y(_04146_));
 sg13g2_xor2_1 _10290_ (.B(_04145_),
    .A(_04138_),
    .X(_04147_));
 sg13g2_a21oi_1 _10291_ (.A1(_04109_),
    .A2(_04127_),
    .Y(_04148_),
    .B1(_04126_));
 sg13g2_nor2_1 _10292_ (.A(_04147_),
    .B(_04148_),
    .Y(_04149_));
 sg13g2_xor2_1 _10293_ (.B(_04148_),
    .A(_04147_),
    .X(_04150_));
 sg13g2_or2_1 _10294_ (.X(_04151_),
    .B(_04150_),
    .A(_04137_));
 sg13g2_a21oi_1 _10295_ (.A1(_04137_),
    .A2(_04150_),
    .Y(_04152_),
    .B1(net2747));
 sg13g2_a21o_1 _10296_ (.A2(_04152_),
    .A1(_04151_),
    .B1(_04136_),
    .X(_00393_));
 sg13g2_and2_1 _10297_ (.A(net3144),
    .B(net2815),
    .X(_04153_));
 sg13g2_a21oi_1 _10298_ (.A1(_04139_),
    .A2(_04144_),
    .Y(_04154_),
    .B1(_04146_));
 sg13g2_nor2_1 _10299_ (.A(_04118_),
    .B(_04141_),
    .Y(_04155_));
 sg13g2_mux2_1 _10300_ (.A0(_04111_),
    .A1(_04112_),
    .S(_04142_),
    .X(_04156_));
 sg13g2_xnor2_1 _10301_ (.Y(_04157_),
    .A(_04155_),
    .B(_04156_));
 sg13g2_a21oi_1 _10302_ (.A1(_04113_),
    .A2(_04118_),
    .Y(_04158_),
    .B1(_04157_));
 sg13g2_xnor2_1 _10303_ (.Y(_04159_),
    .A(_04154_),
    .B(_04158_));
 sg13g2_nor2_1 _10304_ (.A(_04149_),
    .B(_04159_),
    .Y(_04160_));
 sg13g2_a21o_1 _10305_ (.A2(_04160_),
    .A1(_04152_),
    .B1(_04153_),
    .X(_00394_));
 sg13g2_nor3_1 _10306_ (.A(\u_toplayer.u_layer2.neuron_index[1] ),
    .B(net3145),
    .C(net3149),
    .Y(_04161_));
 sg13g2_nand2_1 _10307_ (.Y(_04162_),
    .A(_00051_),
    .B(_04161_));
 sg13g2_or3_1 _10308_ (.A(\u_toplayer.u_layer2.neuron_index[4] ),
    .B(\u_toplayer.u_layer2.neuron_index[5] ),
    .C(_04162_),
    .X(_04163_));
 sg13g2_nor3_2 _10309_ (.A(\u_toplayer.u_layer2.neuron_index[1] ),
    .B(\u_toplayer.u_layer2.neuron_index[0] ),
    .C(net3149),
    .Y(_04164_));
 sg13g2_nor2b_1 _10310_ (.A(net3145),
    .B_N(net2950),
    .Y(_04165_));
 sg13g2_xnor2_1 _10311_ (.Y(_04166_),
    .A(\u_toplayer.u_layer2.neuron_index[4] ),
    .B(_04165_));
 sg13g2_nand2b_1 _10312_ (.Y(_04167_),
    .B(_03731_),
    .A_N(_04166_));
 sg13g2_nand2b_1 _10313_ (.Y(_04168_),
    .B(_03732_),
    .A_N(_04166_));
 sg13g2_or2_2 _10314_ (.X(_04169_),
    .B(net2809),
    .A(net2883));
 sg13g2_mux2_1 _10315_ (.A0(net3080),
    .A1(net911),
    .S(_04169_),
    .X(_00395_));
 sg13g2_mux2_1 _10316_ (.A0(net3079),
    .A1(net913),
    .S(_04169_),
    .X(_00396_));
 sg13g2_mux2_1 _10317_ (.A0(net3076),
    .A1(net912),
    .S(_04169_),
    .X(_00397_));
 sg13g2_mux2_1 _10318_ (.A0(net3074),
    .A1(net936),
    .S(_04169_),
    .X(_00398_));
 sg13g2_mux2_1 _10319_ (.A0(net3071),
    .A1(net914),
    .S(_04169_),
    .X(_00399_));
 sg13g2_mux2_1 _10320_ (.A0(net3069),
    .A1(net935),
    .S(_04169_),
    .X(_00400_));
 sg13g2_mux2_1 _10321_ (.A0(net3067),
    .A1(net946),
    .S(_04169_),
    .X(_00401_));
 sg13g2_mux2_1 _10322_ (.A0(net3066),
    .A1(net956),
    .S(_04169_),
    .X(_00402_));
 sg13g2_and2_2 _10323_ (.A(_01033_),
    .B(_03733_),
    .X(_04170_));
 sg13g2_and2_1 _10324_ (.A(\u_toplayer.u_layer2.neuron_index[0] ),
    .B(_04161_),
    .X(_04171_));
 sg13g2_o21ai_1 _10325_ (.B1(\u_toplayer.u_layer2.neuron_index[5] ),
    .Y(_04172_),
    .A1(\u_toplayer.u_layer2.neuron_index[4] ),
    .A2(_04162_));
 sg13g2_nand2_2 _10326_ (.Y(_04173_),
    .A(net2879),
    .B(_04172_));
 sg13g2_nand2_2 _10327_ (.Y(_04174_),
    .A(_03731_),
    .B(_04166_));
 sg13g2_nor2_2 _10328_ (.A(_04173_),
    .B(net2716),
    .Y(_04175_));
 sg13g2_nand2_2 _10329_ (.Y(_04176_),
    .A(_04171_),
    .B(net2714));
 sg13g2_nand2_1 _10330_ (.Y(_04177_),
    .A(net731),
    .B(_04176_));
 sg13g2_xor2_1 _10331_ (.B(net2950),
    .A(net3145),
    .X(_04178_));
 sg13g2_nor2_2 _10332_ (.A(_04173_),
    .B(_04178_),
    .Y(_04179_));
 sg13g2_nand2_1 _10333_ (.Y(_04180_),
    .A(\u_toplayer.u_layer2.sum[0] ),
    .B(net2924));
 sg13g2_nand3_1 _10334_ (.B(net2925),
    .C(net2823),
    .A(net3081),
    .Y(_04181_));
 sg13g2_nand2_2 _10335_ (.Y(_04182_),
    .A(_03732_),
    .B(_04166_));
 sg13g2_o21ai_1 _10336_ (.B1(_04177_),
    .Y(_00403_),
    .A1(_04181_),
    .A2(net2794));
 sg13g2_nand2_1 _10337_ (.Y(_04183_),
    .A(net383),
    .B(_04176_));
 sg13g2_nand2_1 _10338_ (.Y(_04184_),
    .A(\u_toplayer.u_layer2.sum[1] ),
    .B(_04170_));
 sg13g2_nand3_1 _10339_ (.B(net2925),
    .C(net2824),
    .A(net3079),
    .Y(_04185_));
 sg13g2_o21ai_1 _10340_ (.B1(_04183_),
    .Y(_00404_),
    .A1(net2794),
    .A2(_04185_));
 sg13g2_nand2_1 _10341_ (.Y(_04186_),
    .A(net486),
    .B(_04176_));
 sg13g2_nand2_1 _10342_ (.Y(_04187_),
    .A(\u_toplayer.u_layer2.sum[2] ),
    .B(net2924));
 sg13g2_nand3_1 _10343_ (.B(net2925),
    .C(net2823),
    .A(net3076),
    .Y(_04188_));
 sg13g2_o21ai_1 _10344_ (.B1(_04186_),
    .Y(_00405_),
    .A1(net2794),
    .A2(_04188_));
 sg13g2_nand2_1 _10345_ (.Y(_04189_),
    .A(net494),
    .B(_04176_));
 sg13g2_nand2_1 _10346_ (.Y(_04190_),
    .A(net3074),
    .B(net2924));
 sg13g2_nand3_1 _10347_ (.B(net2925),
    .C(net2824),
    .A(net3075),
    .Y(_04191_));
 sg13g2_o21ai_1 _10348_ (.B1(_04189_),
    .Y(_00406_),
    .A1(net2793),
    .A2(_04191_));
 sg13g2_nand2_1 _10349_ (.Y(_04192_),
    .A(net846),
    .B(_04176_));
 sg13g2_nand2_1 _10350_ (.Y(_04193_),
    .A(net3072),
    .B(net2924));
 sg13g2_nand3_1 _10351_ (.B(net2925),
    .C(net2824),
    .A(net3073),
    .Y(_04194_));
 sg13g2_o21ai_1 _10352_ (.B1(_04192_),
    .Y(_00407_),
    .A1(net2796),
    .A2(_04194_));
 sg13g2_nand2_1 _10353_ (.Y(_04195_),
    .A(net244),
    .B(_04176_));
 sg13g2_nand2_1 _10354_ (.Y(_04196_),
    .A(\u_toplayer.u_layer2.sum[5] ),
    .B(_04170_));
 sg13g2_nand3_1 _10355_ (.B(net2925),
    .C(net2822),
    .A(net3069),
    .Y(_04197_));
 sg13g2_o21ai_1 _10356_ (.B1(_04195_),
    .Y(_00408_),
    .A1(net2794),
    .A2(_04197_));
 sg13g2_nand2_1 _10357_ (.Y(_04198_),
    .A(net578),
    .B(_04176_));
 sg13g2_nand2_1 _10358_ (.Y(_04199_),
    .A(\u_toplayer.u_layer2.sum[6] ),
    .B(net2924));
 sg13g2_nand3_1 _10359_ (.B(net2925),
    .C(net2823),
    .A(net3067),
    .Y(_04200_));
 sg13g2_o21ai_1 _10360_ (.B1(_04198_),
    .Y(_00409_),
    .A1(net2794),
    .A2(_04200_));
 sg13g2_nand2_1 _10361_ (.Y(_04201_),
    .A(net243),
    .B(_04176_));
 sg13g2_nand2_1 _10362_ (.Y(_04202_),
    .A(\u_toplayer.u_layer2.sum[7] ),
    .B(net2924));
 sg13g2_nand3_1 _10363_ (.B(net2925),
    .C(net2822),
    .A(net3066),
    .Y(_04203_));
 sg13g2_o21ai_1 _10364_ (.B1(_04201_),
    .Y(_00410_),
    .A1(net2793),
    .A2(_04203_));
 sg13g2_and2_1 _10365_ (.A(_01033_),
    .B(net2931),
    .X(_04204_));
 sg13g2_nor2b_1 _10366_ (.A(net3145),
    .B_N(net2875),
    .Y(_04205_));
 sg13g2_nand2_2 _10367_ (.Y(_04206_),
    .A(net2714),
    .B(_04205_));
 sg13g2_nand2_1 _10368_ (.Y(_04207_),
    .A(net746),
    .B(_04206_));
 sg13g2_nand3_1 _10369_ (.B(net2881),
    .C(net2877),
    .A(net3081),
    .Y(_04208_));
 sg13g2_nand4_1 _10370_ (.B(net2878),
    .C(net2820),
    .A(net3081),
    .Y(_04209_),
    .D(net2875));
 sg13g2_o21ai_1 _10371_ (.B1(_04207_),
    .Y(_00411_),
    .A1(net2795),
    .A2(_04209_));
 sg13g2_nand2_1 _10372_ (.Y(_04210_),
    .A(net349),
    .B(_04206_));
 sg13g2_nand3_1 _10373_ (.B(net2880),
    .C(net2877),
    .A(net3079),
    .Y(_04211_));
 sg13g2_nand4_1 _10374_ (.B(net2878),
    .C(net2824),
    .A(net3079),
    .Y(_04212_),
    .D(net2877));
 sg13g2_o21ai_1 _10375_ (.B1(_04210_),
    .Y(_00412_),
    .A1(net2796),
    .A2(_04212_));
 sg13g2_nand2_1 _10376_ (.Y(_04213_),
    .A(net412),
    .B(_04206_));
 sg13g2_nand3_1 _10377_ (.B(net2881),
    .C(net2876),
    .A(net3077),
    .Y(_04214_));
 sg13g2_nand4_1 _10378_ (.B(net2878),
    .C(net2821),
    .A(net3076),
    .Y(_04215_),
    .D(net2875));
 sg13g2_o21ai_1 _10379_ (.B1(_04213_),
    .Y(_00413_),
    .A1(net2795),
    .A2(_04215_));
 sg13g2_nand2_1 _10380_ (.Y(_04216_),
    .A(net605),
    .B(_04206_));
 sg13g2_nand3_1 _10381_ (.B(net2881),
    .C(net2876),
    .A(net3075),
    .Y(_04217_));
 sg13g2_nand4_1 _10382_ (.B(net2878),
    .C(net2824),
    .A(net3075),
    .Y(_04218_),
    .D(net2875));
 sg13g2_o21ai_1 _10383_ (.B1(_04216_),
    .Y(_00414_),
    .A1(net2795),
    .A2(_04218_));
 sg13g2_nand2_1 _10384_ (.Y(_04219_),
    .A(net409),
    .B(_04206_));
 sg13g2_nand3_1 _10385_ (.B(net2881),
    .C(net2876),
    .A(net3071),
    .Y(_04220_));
 sg13g2_nand4_1 _10386_ (.B(net2878),
    .C(net2824),
    .A(net3071),
    .Y(_04221_),
    .D(net2875));
 sg13g2_o21ai_1 _10387_ (.B1(_04219_),
    .Y(_00415_),
    .A1(net2796),
    .A2(_04221_));
 sg13g2_nand2_1 _10388_ (.Y(_04222_),
    .A(net420),
    .B(_04206_));
 sg13g2_nand3_1 _10389_ (.B(net2880),
    .C(net2876),
    .A(net3070),
    .Y(_04223_));
 sg13g2_nand4_1 _10390_ (.B(net2878),
    .C(net2821),
    .A(net3069),
    .Y(_04224_),
    .D(net2875));
 sg13g2_o21ai_1 _10391_ (.B1(_04222_),
    .Y(_00416_),
    .A1(net2795),
    .A2(_04224_));
 sg13g2_nand2_1 _10392_ (.Y(_04225_),
    .A(net592),
    .B(_04206_));
 sg13g2_nand3_1 _10393_ (.B(net2880),
    .C(net2876),
    .A(net3068),
    .Y(_04226_));
 sg13g2_nand4_1 _10394_ (.B(net2878),
    .C(net2820),
    .A(net3067),
    .Y(_04227_),
    .D(net2875));
 sg13g2_o21ai_1 _10395_ (.B1(_04225_),
    .Y(_00417_),
    .A1(net2795),
    .A2(_04227_));
 sg13g2_nand2_1 _10396_ (.Y(_04228_),
    .A(net654),
    .B(_04206_));
 sg13g2_nand3_1 _10397_ (.B(net2881),
    .C(net2876),
    .A(net3065),
    .Y(_04229_));
 sg13g2_nand4_1 _10398_ (.B(net2878),
    .C(net2820),
    .A(net3065),
    .Y(_04230_),
    .D(net2875));
 sg13g2_o21ai_1 _10399_ (.B1(_04228_),
    .Y(_00418_),
    .A1(net2795),
    .A2(_04230_));
 sg13g2_nor2_2 _10400_ (.A(net3149),
    .B(_03736_),
    .Y(_04231_));
 sg13g2_nor3_2 _10401_ (.A(net3145),
    .B(net3149),
    .C(_03736_),
    .Y(_04232_));
 sg13g2_nand2_2 _10402_ (.Y(_04233_),
    .A(net2714),
    .B(_04232_));
 sg13g2_nand2_1 _10403_ (.Y(_04234_),
    .A(net489),
    .B(_04233_));
 sg13g2_nand2_1 _10404_ (.Y(_04235_),
    .A(net3081),
    .B(_04231_));
 sg13g2_nand3_1 _10405_ (.B(net2820),
    .C(net2923),
    .A(net3081),
    .Y(_04236_));
 sg13g2_o21ai_1 _10406_ (.B1(_04234_),
    .Y(_00419_),
    .A1(net2716),
    .A2(_04236_));
 sg13g2_nand2_1 _10407_ (.Y(_04237_),
    .A(net480),
    .B(_04233_));
 sg13g2_nand2_1 _10408_ (.Y(_04238_),
    .A(net3079),
    .B(_04231_));
 sg13g2_nand3_1 _10409_ (.B(net2821),
    .C(net2923),
    .A(net3079),
    .Y(_04239_));
 sg13g2_o21ai_1 _10410_ (.B1(_04237_),
    .Y(_00420_),
    .A1(_04174_),
    .A2(_04239_));
 sg13g2_nand2_1 _10411_ (.Y(_04240_),
    .A(net210),
    .B(_04233_));
 sg13g2_nand2_1 _10412_ (.Y(_04241_),
    .A(net3076),
    .B(net2922));
 sg13g2_nand3_1 _10413_ (.B(net2821),
    .C(net2923),
    .A(net3076),
    .Y(_04242_));
 sg13g2_o21ai_1 _10414_ (.B1(_04240_),
    .Y(_00421_),
    .A1(net2716),
    .A2(_04242_));
 sg13g2_nand2_1 _10415_ (.Y(_04243_),
    .A(net587),
    .B(_04233_));
 sg13g2_nand2_1 _10416_ (.Y(_04244_),
    .A(net3075),
    .B(net2922));
 sg13g2_nand3_1 _10417_ (.B(net2820),
    .C(net2923),
    .A(net3075),
    .Y(_04245_));
 sg13g2_o21ai_1 _10418_ (.B1(_04243_),
    .Y(_00422_),
    .A1(net2716),
    .A2(_04245_));
 sg13g2_nand2_1 _10419_ (.Y(_04246_),
    .A(net364),
    .B(_04233_));
 sg13g2_nand2_1 _10420_ (.Y(_04247_),
    .A(net3071),
    .B(net2922));
 sg13g2_nand3_1 _10421_ (.B(net2820),
    .C(net2923),
    .A(net3071),
    .Y(_04248_));
 sg13g2_o21ai_1 _10422_ (.B1(_04246_),
    .Y(_00423_),
    .A1(net2716),
    .A2(_04248_));
 sg13g2_nand2_1 _10423_ (.Y(_04249_),
    .A(net537),
    .B(_04233_));
 sg13g2_nand2_1 _10424_ (.Y(_04250_),
    .A(net3069),
    .B(net2922));
 sg13g2_nand3_1 _10425_ (.B(net2821),
    .C(net2923),
    .A(net3069),
    .Y(_04251_));
 sg13g2_o21ai_1 _10426_ (.B1(_04249_),
    .Y(_00424_),
    .A1(net2716),
    .A2(_04251_));
 sg13g2_nand2_1 _10427_ (.Y(_04252_),
    .A(net741),
    .B(_04233_));
 sg13g2_nand2_1 _10428_ (.Y(_04253_),
    .A(net3067),
    .B(net2922));
 sg13g2_nand3_1 _10429_ (.B(net2820),
    .C(net2923),
    .A(net3067),
    .Y(_04254_));
 sg13g2_o21ai_1 _10430_ (.B1(_04252_),
    .Y(_00425_),
    .A1(net2716),
    .A2(_04254_));
 sg13g2_nand2_1 _10431_ (.Y(_04255_),
    .A(net758),
    .B(_04233_));
 sg13g2_nand2_1 _10432_ (.Y(_04256_),
    .A(net3065),
    .B(net2922));
 sg13g2_nand3_1 _10433_ (.B(net2820),
    .C(net2923),
    .A(net3065),
    .Y(_04257_));
 sg13g2_o21ai_1 _10434_ (.B1(_04255_),
    .Y(_00426_),
    .A1(net2716),
    .A2(_04257_));
 sg13g2_nor3_2 _10435_ (.A(\u_toplayer.u_layer2.neuron_index[1] ),
    .B(\u_toplayer.u_layer2.neuron_index[0] ),
    .C(_01033_),
    .Y(_04258_));
 sg13g2_nor2b_1 _10436_ (.A(net3148),
    .B_N(net2919),
    .Y(_04259_));
 sg13g2_nand2_2 _10437_ (.Y(_04260_),
    .A(net2715),
    .B(_04259_));
 sg13g2_nand2_1 _10438_ (.Y(_04261_),
    .A(net603),
    .B(_04260_));
 sg13g2_nand2_1 _10439_ (.Y(_04262_),
    .A(\u_toplayer.u_layer2.sum[0] ),
    .B(net2920));
 sg13g2_nand3_1 _10440_ (.B(net2826),
    .C(net2919),
    .A(net3080),
    .Y(_04263_));
 sg13g2_o21ai_1 _10441_ (.B1(_04261_),
    .Y(_00427_),
    .A1(net2799),
    .A2(_04263_));
 sg13g2_nand2_1 _10442_ (.Y(_04264_),
    .A(net616),
    .B(_04260_));
 sg13g2_nand2_1 _10443_ (.Y(_04265_),
    .A(\u_toplayer.u_layer2.sum[1] ),
    .B(net2920));
 sg13g2_nand3_1 _10444_ (.B(net2827),
    .C(net2919),
    .A(net3078),
    .Y(_04266_));
 sg13g2_o21ai_1 _10445_ (.B1(_04264_),
    .Y(_00428_),
    .A1(net2800),
    .A2(_04266_));
 sg13g2_nand2_1 _10446_ (.Y(_04267_),
    .A(net837),
    .B(_04260_));
 sg13g2_nand2_1 _10447_ (.Y(_04268_),
    .A(net3077),
    .B(net2920));
 sg13g2_nand3_1 _10448_ (.B(net2827),
    .C(net2921),
    .A(\u_toplayer.u_layer2.sum[2] ),
    .Y(_04269_));
 sg13g2_o21ai_1 _10449_ (.B1(_04267_),
    .Y(_00429_),
    .A1(net2799),
    .A2(_04269_));
 sg13g2_nand2_1 _10450_ (.Y(_04270_),
    .A(net685),
    .B(_04260_));
 sg13g2_nand2_1 _10451_ (.Y(_04271_),
    .A(net3074),
    .B(net2920));
 sg13g2_nand3_1 _10452_ (.B(net2827),
    .C(net2919),
    .A(\u_toplayer.u_layer2.sum[3] ),
    .Y(_04272_));
 sg13g2_o21ai_1 _10453_ (.B1(_04270_),
    .Y(_00430_),
    .A1(net2800),
    .A2(_04272_));
 sg13g2_nand2_1 _10454_ (.Y(_04273_),
    .A(net609),
    .B(_04260_));
 sg13g2_nand2_1 _10455_ (.Y(_04274_),
    .A(net3072),
    .B(net2921));
 sg13g2_nand3_1 _10456_ (.B(net2826),
    .C(net2919),
    .A(net3072),
    .Y(_04275_));
 sg13g2_o21ai_1 _10457_ (.B1(_04273_),
    .Y(_00431_),
    .A1(net2798),
    .A2(_04275_));
 sg13g2_nand2_1 _10458_ (.Y(_04276_),
    .A(net526),
    .B(_04260_));
 sg13g2_nand2_1 _10459_ (.Y(_04277_),
    .A(net3070),
    .B(net2920));
 sg13g2_nand3_1 _10460_ (.B(net2826),
    .C(net2919),
    .A(\u_toplayer.u_layer2.sum[5] ),
    .Y(_04278_));
 sg13g2_o21ai_1 _10461_ (.B1(_04276_),
    .Y(_00432_),
    .A1(net2798),
    .A2(_04278_));
 sg13g2_nand2_1 _10462_ (.Y(_04279_),
    .A(net172),
    .B(_04260_));
 sg13g2_nand2_1 _10463_ (.Y(_04280_),
    .A(net3068),
    .B(net2920));
 sg13g2_nand3_1 _10464_ (.B(net2825),
    .C(net2919),
    .A(\u_toplayer.u_layer2.sum[6] ),
    .Y(_04281_));
 sg13g2_o21ai_1 _10465_ (.B1(_04279_),
    .Y(_00433_),
    .A1(net2798),
    .A2(_04281_));
 sg13g2_nand2_1 _10466_ (.Y(_04282_),
    .A(net742),
    .B(_04260_));
 sg13g2_nand2_1 _10467_ (.Y(_04283_),
    .A(net3066),
    .B(net2921));
 sg13g2_nand3_1 _10468_ (.B(net2826),
    .C(net2919),
    .A(\u_toplayer.u_layer2.sum[7] ),
    .Y(_04284_));
 sg13g2_o21ai_1 _10469_ (.B1(_04282_),
    .Y(_00434_),
    .A1(net2798),
    .A2(_04284_));
 sg13g2_and2_1 _10470_ (.A(net3153),
    .B(_03733_),
    .X(_04285_));
 sg13g2_nor2b_1 _10471_ (.A(net3148),
    .B_N(net2916),
    .Y(_04286_));
 sg13g2_nand2_2 _10472_ (.Y(_04287_),
    .A(net2715),
    .B(_04286_));
 sg13g2_nand2_1 _10473_ (.Y(_04288_),
    .A(net461),
    .B(_04287_));
 sg13g2_nand2_1 _10474_ (.Y(_04289_),
    .A(\u_toplayer.u_layer2.sum[0] ),
    .B(net2918));
 sg13g2_nand3_1 _10475_ (.B(net2827),
    .C(net2916),
    .A(net3080),
    .Y(_04290_));
 sg13g2_o21ai_1 _10476_ (.B1(_04288_),
    .Y(_00435_),
    .A1(net2799),
    .A2(_04290_));
 sg13g2_nand2_1 _10477_ (.Y(_04291_),
    .A(net702),
    .B(_04287_));
 sg13g2_nand2_1 _10478_ (.Y(_04292_),
    .A(net3078),
    .B(net2917));
 sg13g2_nand3_1 _10479_ (.B(net2827),
    .C(net2918),
    .A(net3078),
    .Y(_04293_));
 sg13g2_o21ai_1 _10480_ (.B1(_04291_),
    .Y(_00436_),
    .A1(net2800),
    .A2(_04293_));
 sg13g2_nand2_1 _10481_ (.Y(_04294_),
    .A(net842),
    .B(_04287_));
 sg13g2_nand2_1 _10482_ (.Y(_04295_),
    .A(net3077),
    .B(net2917));
 sg13g2_nand3_1 _10483_ (.B(net2827),
    .C(net2916),
    .A(\u_toplayer.u_layer2.sum[2] ),
    .Y(_04296_));
 sg13g2_o21ai_1 _10484_ (.B1(_04294_),
    .Y(_00437_),
    .A1(net2799),
    .A2(_04296_));
 sg13g2_nand2_1 _10485_ (.Y(_04297_),
    .A(net455),
    .B(_04287_));
 sg13g2_nand2_1 _10486_ (.Y(_04298_),
    .A(\u_toplayer.u_layer2.sum[3] ),
    .B(net2917));
 sg13g2_nand3_1 _10487_ (.B(net2827),
    .C(net2916),
    .A(\u_toplayer.u_layer2.sum[3] ),
    .Y(_04299_));
 sg13g2_o21ai_1 _10488_ (.B1(_04297_),
    .Y(_00438_),
    .A1(net2800),
    .A2(_04299_));
 sg13g2_nand2_1 _10489_ (.Y(_04300_),
    .A(net282),
    .B(_04287_));
 sg13g2_nand2_1 _10490_ (.Y(_04301_),
    .A(net3073),
    .B(net2917));
 sg13g2_nand3_1 _10491_ (.B(net2826),
    .C(net2916),
    .A(net3072),
    .Y(_04302_));
 sg13g2_o21ai_1 _10492_ (.B1(_04300_),
    .Y(_00439_),
    .A1(net2798),
    .A2(_04302_));
 sg13g2_nand2_1 _10493_ (.Y(_04303_),
    .A(net453),
    .B(_04287_));
 sg13g2_nand2_1 _10494_ (.Y(_04304_),
    .A(net3070),
    .B(net2917));
 sg13g2_nand3_1 _10495_ (.B(net2826),
    .C(net2916),
    .A(\u_toplayer.u_layer2.sum[5] ),
    .Y(_04305_));
 sg13g2_o21ai_1 _10496_ (.B1(_04303_),
    .Y(_00440_),
    .A1(net2798),
    .A2(_04305_));
 sg13g2_nand2_1 _10497_ (.Y(_04306_),
    .A(net789),
    .B(_04287_));
 sg13g2_nand2_1 _10498_ (.Y(_04307_),
    .A(net3068),
    .B(net2918));
 sg13g2_nand3_1 _10499_ (.B(net2826),
    .C(net2916),
    .A(\u_toplayer.u_layer2.sum[6] ),
    .Y(_04308_));
 sg13g2_o21ai_1 _10500_ (.B1(_04306_),
    .Y(_00441_),
    .A1(net2798),
    .A2(_04308_));
 sg13g2_nand2_1 _10501_ (.Y(_04309_),
    .A(net188),
    .B(_04287_));
 sg13g2_nand2_1 _10502_ (.Y(_04310_),
    .A(net3066),
    .B(net2917));
 sg13g2_nand3_1 _10503_ (.B(net2826),
    .C(net2916),
    .A(\u_toplayer.u_layer2.sum[7] ),
    .Y(_04311_));
 sg13g2_o21ai_1 _10504_ (.B1(_04309_),
    .Y(_00442_),
    .A1(net2798),
    .A2(_04311_));
 sg13g2_nand2_1 _10505_ (.Y(_04312_),
    .A(net3150),
    .B(net2931));
 sg13g2_nor2_1 _10506_ (.A(net3146),
    .B(_04312_),
    .Y(_04313_));
 sg13g2_nand2_2 _10507_ (.Y(_04314_),
    .A(net2715),
    .B(_04313_));
 sg13g2_nand2_1 _10508_ (.Y(_04315_),
    .A(net524),
    .B(_04314_));
 sg13g2_nand3_1 _10509_ (.B(net3080),
    .C(net2930),
    .A(net3151),
    .Y(_04316_));
 sg13g2_nand4_1 _10510_ (.B(net3080),
    .C(_03734_),
    .A(net3153),
    .Y(_04317_),
    .D(net2825));
 sg13g2_o21ai_1 _10511_ (.B1(_04315_),
    .Y(_00443_),
    .A1(net2797),
    .A2(_04317_));
 sg13g2_nand2_1 _10512_ (.Y(_04318_),
    .A(net651),
    .B(_04314_));
 sg13g2_nand3_1 _10513_ (.B(net3078),
    .C(net2930),
    .A(net3151),
    .Y(_04319_));
 sg13g2_nand4_1 _10514_ (.B(net3078),
    .C(net2931),
    .A(net3153),
    .Y(_04320_),
    .D(net2828));
 sg13g2_o21ai_1 _10515_ (.B1(_04318_),
    .Y(_00444_),
    .A1(net2801),
    .A2(_04320_));
 sg13g2_nand2_1 _10516_ (.Y(_04321_),
    .A(net231),
    .B(_04314_));
 sg13g2_nand3_1 _10517_ (.B(net3077),
    .C(net2929),
    .A(net3152),
    .Y(_04322_));
 sg13g2_nand4_1 _10518_ (.B(net3076),
    .C(net2931),
    .A(net3150),
    .Y(_04323_),
    .D(net2825));
 sg13g2_o21ai_1 _10519_ (.B1(_04321_),
    .Y(_00445_),
    .A1(net2797),
    .A2(_04323_));
 sg13g2_nand2_1 _10520_ (.Y(_04324_),
    .A(net676),
    .B(_04314_));
 sg13g2_nand3_1 _10521_ (.B(net3074),
    .C(net2929),
    .A(net3151),
    .Y(_04325_));
 sg13g2_nand4_1 _10522_ (.B(net3074),
    .C(net2930),
    .A(net3152),
    .Y(_04326_),
    .D(net2828));
 sg13g2_o21ai_1 _10523_ (.B1(_04324_),
    .Y(_00446_),
    .A1(net2801),
    .A2(_04326_));
 sg13g2_nand2_1 _10524_ (.Y(_04327_),
    .A(net628),
    .B(_04314_));
 sg13g2_nand3_1 _10525_ (.B(net3072),
    .C(net2929),
    .A(net3151),
    .Y(_04328_));
 sg13g2_nand4_1 _10526_ (.B(net3072),
    .C(_03734_),
    .A(net3153),
    .Y(_04329_),
    .D(net2825));
 sg13g2_o21ai_1 _10527_ (.B1(_04327_),
    .Y(_00447_),
    .A1(net2797),
    .A2(_04329_));
 sg13g2_nand2_1 _10528_ (.Y(_04330_),
    .A(net565),
    .B(_04314_));
 sg13g2_nand3_1 _10529_ (.B(net3070),
    .C(net2929),
    .A(net3151),
    .Y(_04331_));
 sg13g2_nand4_1 _10530_ (.B(net3069),
    .C(net2931),
    .A(net3150),
    .Y(_04332_),
    .D(net2822));
 sg13g2_o21ai_1 _10531_ (.B1(_04330_),
    .Y(_00448_),
    .A1(net2793),
    .A2(_04332_));
 sg13g2_nand2_1 _10532_ (.Y(_04333_),
    .A(net803),
    .B(_04314_));
 sg13g2_nand3_1 _10533_ (.B(net3068),
    .C(net2929),
    .A(net3151),
    .Y(_04334_));
 sg13g2_nand4_1 _10534_ (.B(net3067),
    .C(net2931),
    .A(net3149),
    .Y(_04335_),
    .D(net2822));
 sg13g2_o21ai_1 _10535_ (.B1(_04333_),
    .Y(_00449_),
    .A1(net2793),
    .A2(_04335_));
 sg13g2_nand2_1 _10536_ (.Y(_04336_),
    .A(net613),
    .B(_04314_));
 sg13g2_nand3_1 _10537_ (.B(net3066),
    .C(net2929),
    .A(net3152),
    .Y(_04337_));
 sg13g2_nand4_1 _10538_ (.B(net3065),
    .C(net2931),
    .A(net3149),
    .Y(_04338_),
    .D(net2822));
 sg13g2_o21ai_1 _10539_ (.B1(_04336_),
    .Y(_00450_),
    .A1(net2793),
    .A2(_04338_));
 sg13g2_nor3_2 _10540_ (.A(net3145),
    .B(_01033_),
    .C(_03736_),
    .Y(_04339_));
 sg13g2_nand2_2 _10541_ (.Y(_04340_),
    .A(net2714),
    .B(_04339_));
 sg13g2_nand2_1 _10542_ (.Y(_04341_),
    .A(net612),
    .B(_04340_));
 sg13g2_nand2_1 _10543_ (.Y(_04342_),
    .A(net3080),
    .B(net2928));
 sg13g2_nand3_1 _10544_ (.B(net2926),
    .C(net2825),
    .A(net3080),
    .Y(_04343_));
 sg13g2_o21ai_1 _10545_ (.B1(_04341_),
    .Y(_00451_),
    .A1(net2797),
    .A2(_04343_));
 sg13g2_nand2_1 _10546_ (.Y(_04344_),
    .A(net590),
    .B(_04340_));
 sg13g2_nand2_1 _10547_ (.Y(_04345_),
    .A(net3078),
    .B(net2927));
 sg13g2_nand3_1 _10548_ (.B(net2928),
    .C(net2828),
    .A(net3078),
    .Y(_04346_));
 sg13g2_o21ai_1 _10549_ (.B1(_04344_),
    .Y(_00452_),
    .A1(net2797),
    .A2(_04346_));
 sg13g2_nand2_1 _10550_ (.Y(_04347_),
    .A(net638),
    .B(_04340_));
 sg13g2_nand2_1 _10551_ (.Y(_04348_),
    .A(net3077),
    .B(net2927));
 sg13g2_nand3_1 _10552_ (.B(net2926),
    .C(net2825),
    .A(net3076),
    .Y(_04349_));
 sg13g2_o21ai_1 _10553_ (.B1(_04347_),
    .Y(_00453_),
    .A1(net2797),
    .A2(_04349_));
 sg13g2_nand2_1 _10554_ (.Y(_04350_),
    .A(net194),
    .B(_04340_));
 sg13g2_nand2_1 _10555_ (.Y(_04351_),
    .A(net3074),
    .B(net2927));
 sg13g2_nand3_1 _10556_ (.B(net2927),
    .C(net2825),
    .A(net3074),
    .Y(_04352_));
 sg13g2_o21ai_1 _10557_ (.B1(_04350_),
    .Y(_00454_),
    .A1(net2797),
    .A2(_04352_));
 sg13g2_nand2_1 _10558_ (.Y(_04353_),
    .A(net559),
    .B(_04340_));
 sg13g2_nand2_1 _10559_ (.Y(_04354_),
    .A(net3072),
    .B(net2927));
 sg13g2_nand3_1 _10560_ (.B(net2926),
    .C(net2825),
    .A(net3072),
    .Y(_04355_));
 sg13g2_o21ai_1 _10561_ (.B1(_04353_),
    .Y(_00455_),
    .A1(net2797),
    .A2(_04355_));
 sg13g2_nand2_1 _10562_ (.Y(_04356_),
    .A(net269),
    .B(_04340_));
 sg13g2_nand2_1 _10563_ (.Y(_04357_),
    .A(net3070),
    .B(net2927));
 sg13g2_nand3_1 _10564_ (.B(net2926),
    .C(net2822),
    .A(net3069),
    .Y(_04358_));
 sg13g2_o21ai_1 _10565_ (.B1(_04356_),
    .Y(_00456_),
    .A1(net2793),
    .A2(_04358_));
 sg13g2_nand2_1 _10566_ (.Y(_04359_),
    .A(net433),
    .B(_04340_));
 sg13g2_nand2_1 _10567_ (.Y(_04360_),
    .A(net3068),
    .B(net2927));
 sg13g2_nand3_1 _10568_ (.B(net2926),
    .C(net2822),
    .A(net3067),
    .Y(_04361_));
 sg13g2_o21ai_1 _10569_ (.B1(_04359_),
    .Y(_00457_),
    .A1(net2793),
    .A2(_04361_));
 sg13g2_nand2_1 _10570_ (.Y(_04362_),
    .A(net404),
    .B(_04340_));
 sg13g2_nand2_1 _10571_ (.Y(_04363_),
    .A(net3066),
    .B(net2927));
 sg13g2_nand3_1 _10572_ (.B(net2926),
    .C(net2822),
    .A(net3065),
    .Y(_04364_));
 sg13g2_o21ai_1 _10573_ (.B1(_04362_),
    .Y(_00458_),
    .A1(net2793),
    .A2(_04364_));
 sg13g2_nand3_1 _10574_ (.B(net2948),
    .C(_04175_),
    .A(net3147),
    .Y(_04365_));
 sg13g2_nand2_1 _10575_ (.Y(_04366_),
    .A(net580),
    .B(_04365_));
 sg13g2_nand3_1 _10576_ (.B(net2879),
    .C(net2950),
    .A(net3081),
    .Y(_04367_));
 sg13g2_nand4_1 _10577_ (.B(net2882),
    .C(net2948),
    .A(net3080),
    .Y(_04368_),
    .D(net2829));
 sg13g2_o21ai_1 _10578_ (.B1(_04366_),
    .Y(_00459_),
    .A1(net2802),
    .A2(_04368_));
 sg13g2_nand2_1 _10579_ (.Y(_04369_),
    .A(net538),
    .B(_04365_));
 sg13g2_nand3_1 _10580_ (.B(net2880),
    .C(net2949),
    .A(net3079),
    .Y(_04370_));
 sg13g2_nand4_1 _10581_ (.B(net2882),
    .C(net2949),
    .A(net3078),
    .Y(_04371_),
    .D(net2829));
 sg13g2_o21ai_1 _10582_ (.B1(_04369_),
    .Y(_00460_),
    .A1(net2802),
    .A2(_04371_));
 sg13g2_nand2_1 _10583_ (.Y(_04372_),
    .A(net399),
    .B(_04365_));
 sg13g2_nand3_1 _10584_ (.B(net2879),
    .C(net2950),
    .A(net3076),
    .Y(_04373_));
 sg13g2_nand4_1 _10585_ (.B(net2881),
    .C(net2948),
    .A(net3077),
    .Y(_04374_),
    .D(net2829));
 sg13g2_o21ai_1 _10586_ (.B1(_04372_),
    .Y(_00461_),
    .A1(net2802),
    .A2(_04374_));
 sg13g2_nand2_1 _10587_ (.Y(_04375_),
    .A(net709),
    .B(_04365_));
 sg13g2_nand3_1 _10588_ (.B(net2879),
    .C(net2950),
    .A(net3075),
    .Y(_04376_));
 sg13g2_nand4_1 _10589_ (.B(net2881),
    .C(net2948),
    .A(net3074),
    .Y(_04377_),
    .D(net2829));
 sg13g2_o21ai_1 _10590_ (.B1(_04375_),
    .Y(_00462_),
    .A1(net2802),
    .A2(_04377_));
 sg13g2_nand2_1 _10591_ (.Y(_04378_),
    .A(net437),
    .B(_04365_));
 sg13g2_nand3_1 _10592_ (.B(net2880),
    .C(net2949),
    .A(net3071),
    .Y(_04379_));
 sg13g2_nand4_1 _10593_ (.B(net2882),
    .C(net2948),
    .A(net3071),
    .Y(_04380_),
    .D(net2829));
 sg13g2_o21ai_1 _10594_ (.B1(_04378_),
    .Y(_00463_),
    .A1(net2802),
    .A2(_04380_));
 sg13g2_nand2_1 _10595_ (.Y(_04381_),
    .A(net443),
    .B(_04365_));
 sg13g2_nand3_1 _10596_ (.B(net2879),
    .C(net2950),
    .A(net3069),
    .Y(_04382_));
 sg13g2_nand4_1 _10597_ (.B(net2882),
    .C(net2949),
    .A(net3070),
    .Y(_04383_),
    .D(_04179_));
 sg13g2_o21ai_1 _10598_ (.B1(_04381_),
    .Y(_00464_),
    .A1(_04182_),
    .A2(_04383_));
 sg13g2_nand2_1 _10599_ (.Y(_04384_),
    .A(net429),
    .B(_04365_));
 sg13g2_nand3_1 _10600_ (.B(net2879),
    .C(net2950),
    .A(net3067),
    .Y(_04385_));
 sg13g2_nand4_1 _10601_ (.B(net2881),
    .C(net2948),
    .A(net3068),
    .Y(_04386_),
    .D(net2829));
 sg13g2_o21ai_1 _10602_ (.B1(_04384_),
    .Y(_00465_),
    .A1(net2802),
    .A2(_04386_));
 sg13g2_nand2_1 _10603_ (.Y(_04387_),
    .A(net760),
    .B(_04365_));
 sg13g2_nand3_1 _10604_ (.B(net2879),
    .C(net2950),
    .A(net3065),
    .Y(_04388_));
 sg13g2_nand4_1 _10605_ (.B(net2883),
    .C(net2948),
    .A(net3066),
    .Y(_04389_),
    .D(net2829));
 sg13g2_o21ai_1 _10606_ (.B1(_04387_),
    .Y(_00466_),
    .A1(net2802),
    .A2(_04389_));
 sg13g2_nand3_1 _10607_ (.B(net2924),
    .C(net2715),
    .A(net3147),
    .Y(_04390_));
 sg13g2_nand2_1 _10608_ (.Y(_04391_),
    .A(net438),
    .B(_04390_));
 sg13g2_nand2_2 _10609_ (.Y(_04392_),
    .A(net2714),
    .B(_04178_));
 sg13g2_o21ai_1 _10610_ (.B1(_04391_),
    .Y(_00467_),
    .A1(_04180_),
    .A2(net2708));
 sg13g2_nand2_1 _10611_ (.Y(_04393_),
    .A(net753),
    .B(_04390_));
 sg13g2_o21ai_1 _10612_ (.B1(_04393_),
    .Y(_00468_),
    .A1(_04184_),
    .A2(net2710));
 sg13g2_nand2_1 _10613_ (.Y(_04394_),
    .A(net496),
    .B(_04390_));
 sg13g2_o21ai_1 _10614_ (.B1(_04394_),
    .Y(_00469_),
    .A1(_04187_),
    .A2(net2710));
 sg13g2_nand2_1 _10615_ (.Y(_04395_),
    .A(net556),
    .B(_04390_));
 sg13g2_o21ai_1 _10616_ (.B1(_04395_),
    .Y(_00470_),
    .A1(_04190_),
    .A2(net2710));
 sg13g2_nand2_1 _10617_ (.Y(_04396_),
    .A(net465),
    .B(_04390_));
 sg13g2_o21ai_1 _10618_ (.B1(_04396_),
    .Y(_00471_),
    .A1(_04193_),
    .A2(net2707));
 sg13g2_nand2_1 _10619_ (.Y(_04397_),
    .A(net665),
    .B(_04390_));
 sg13g2_o21ai_1 _10620_ (.B1(_04397_),
    .Y(_00472_),
    .A1(_04196_),
    .A2(net2708));
 sg13g2_nand2_1 _10621_ (.Y(_04398_),
    .A(net339),
    .B(_04390_));
 sg13g2_o21ai_1 _10622_ (.B1(_04398_),
    .Y(_00473_),
    .A1(_04199_),
    .A2(net2708));
 sg13g2_nand2_1 _10623_ (.Y(_04399_),
    .A(net704),
    .B(_04390_));
 sg13g2_o21ai_1 _10624_ (.B1(_04399_),
    .Y(_00474_),
    .A1(_04202_),
    .A2(net2707));
 sg13g2_nand3_1 _10625_ (.B(net2714),
    .C(net2876),
    .A(net3146),
    .Y(_04400_));
 sg13g2_nand2_1 _10626_ (.Y(_04401_),
    .A(net317),
    .B(_04400_));
 sg13g2_o21ai_1 _10627_ (.B1(_04401_),
    .Y(_00475_),
    .A1(_04208_),
    .A2(net2702));
 sg13g2_nand2_1 _10628_ (.Y(_04402_),
    .A(net750),
    .B(_04400_));
 sg13g2_o21ai_1 _10629_ (.B1(_04402_),
    .Y(_00476_),
    .A1(_04211_),
    .A2(net2702));
 sg13g2_nand2_1 _10630_ (.Y(_04403_),
    .A(net275),
    .B(_04400_));
 sg13g2_o21ai_1 _10631_ (.B1(_04403_),
    .Y(_00477_),
    .A1(_04214_),
    .A2(net2704));
 sg13g2_nand2_1 _10632_ (.Y(_04404_),
    .A(net606),
    .B(_04400_));
 sg13g2_o21ai_1 _10633_ (.B1(_04404_),
    .Y(_00478_),
    .A1(_04217_),
    .A2(net2703));
 sg13g2_nand2_1 _10634_ (.Y(_04405_),
    .A(net343),
    .B(_04400_));
 sg13g2_o21ai_1 _10635_ (.B1(_04405_),
    .Y(_00479_),
    .A1(_04220_),
    .A2(net2704));
 sg13g2_nand2_1 _10636_ (.Y(_04406_),
    .A(net233),
    .B(_04400_));
 sg13g2_o21ai_1 _10637_ (.B1(_04406_),
    .Y(_00480_),
    .A1(_04223_),
    .A2(net2703));
 sg13g2_nand2_1 _10638_ (.Y(_04407_),
    .A(net747),
    .B(_04400_));
 sg13g2_o21ai_1 _10639_ (.B1(_04407_),
    .Y(_00481_),
    .A1(_04226_),
    .A2(net2702));
 sg13g2_nand2_1 _10640_ (.Y(_04408_),
    .A(net338),
    .B(_04400_));
 sg13g2_o21ai_1 _10641_ (.B1(_04408_),
    .Y(_00482_),
    .A1(_04229_),
    .A2(net2702));
 sg13g2_nand3_1 _10642_ (.B(net2714),
    .C(net2922),
    .A(net3146),
    .Y(_04409_));
 sg13g2_nand2_1 _10643_ (.Y(_04410_),
    .A(net655),
    .B(_04409_));
 sg13g2_o21ai_1 _10644_ (.B1(_04410_),
    .Y(_00483_),
    .A1(_04235_),
    .A2(net2702));
 sg13g2_nand2_1 _10645_ (.Y(_04411_),
    .A(net201),
    .B(_04409_));
 sg13g2_o21ai_1 _10646_ (.B1(_04411_),
    .Y(_00484_),
    .A1(_04238_),
    .A2(net2703));
 sg13g2_nand2_1 _10647_ (.Y(_04412_),
    .A(net185),
    .B(_04409_));
 sg13g2_o21ai_1 _10648_ (.B1(_04412_),
    .Y(_00485_),
    .A1(_04241_),
    .A2(net2704));
 sg13g2_nand2_1 _10649_ (.Y(_04413_),
    .A(net202),
    .B(_04409_));
 sg13g2_o21ai_1 _10650_ (.B1(_04413_),
    .Y(_00486_),
    .A1(_04244_),
    .A2(net2703));
 sg13g2_nand2_1 _10651_ (.Y(_04414_),
    .A(net166),
    .B(_04409_));
 sg13g2_o21ai_1 _10652_ (.B1(_04414_),
    .Y(_00487_),
    .A1(_04247_),
    .A2(net2704));
 sg13g2_nand2_1 _10653_ (.Y(_04415_),
    .A(net250),
    .B(_04409_));
 sg13g2_o21ai_1 _10654_ (.B1(_04415_),
    .Y(_00488_),
    .A1(_04250_),
    .A2(net2702));
 sg13g2_nand2_1 _10655_ (.Y(_04416_),
    .A(net260),
    .B(_04409_));
 sg13g2_o21ai_1 _10656_ (.B1(_04416_),
    .Y(_00489_),
    .A1(_04253_),
    .A2(net2702));
 sg13g2_nand2_1 _10657_ (.Y(_04417_),
    .A(net214),
    .B(_04409_));
 sg13g2_o21ai_1 _10658_ (.B1(_04417_),
    .Y(_00490_),
    .A1(_04256_),
    .A2(net2702));
 sg13g2_nand3_1 _10659_ (.B(net2715),
    .C(net2920),
    .A(net3147),
    .Y(_04418_));
 sg13g2_nand2_1 _10660_ (.Y(_04419_),
    .A(net381),
    .B(_04418_));
 sg13g2_o21ai_1 _10661_ (.B1(_04419_),
    .Y(_00491_),
    .A1(_04262_),
    .A2(net2708));
 sg13g2_nand2_1 _10662_ (.Y(_04420_),
    .A(net397),
    .B(_04418_));
 sg13g2_o21ai_1 _10663_ (.B1(_04420_),
    .Y(_00492_),
    .A1(_04265_),
    .A2(net2708));
 sg13g2_nand2_1 _10664_ (.Y(_04421_),
    .A(net635),
    .B(_04418_));
 sg13g2_o21ai_1 _10665_ (.B1(_04421_),
    .Y(_00493_),
    .A1(_04268_),
    .A2(net2709));
 sg13g2_nand2_1 _10666_ (.Y(_04422_),
    .A(net387),
    .B(_04418_));
 sg13g2_o21ai_1 _10667_ (.B1(_04422_),
    .Y(_00494_),
    .A1(_04271_),
    .A2(net2709));
 sg13g2_nand2_1 _10668_ (.Y(_04423_),
    .A(net347),
    .B(_04418_));
 sg13g2_o21ai_1 _10669_ (.B1(_04423_),
    .Y(_00495_),
    .A1(_04274_),
    .A2(net2706));
 sg13g2_nand2_1 _10670_ (.Y(_04424_),
    .A(net588),
    .B(_04418_));
 sg13g2_o21ai_1 _10671_ (.B1(_04424_),
    .Y(_00496_),
    .A1(_04277_),
    .A2(net2709));
 sg13g2_nand2_1 _10672_ (.Y(_04425_),
    .A(net632),
    .B(_04418_));
 sg13g2_o21ai_1 _10673_ (.B1(_04425_),
    .Y(_00497_),
    .A1(_04280_),
    .A2(net2709));
 sg13g2_nand2_1 _10674_ (.Y(_04426_),
    .A(net396),
    .B(_04418_));
 sg13g2_o21ai_1 _10675_ (.B1(_04426_),
    .Y(_00498_),
    .A1(_04283_),
    .A2(net2706));
 sg13g2_nand3_1 _10676_ (.B(net2715),
    .C(net2917),
    .A(net3147),
    .Y(_04427_));
 sg13g2_nand2_1 _10677_ (.Y(_04428_),
    .A(net207),
    .B(_04427_));
 sg13g2_o21ai_1 _10678_ (.B1(_04428_),
    .Y(_00499_),
    .A1(_04289_),
    .A2(net2708));
 sg13g2_nand2_1 _10679_ (.Y(_04429_),
    .A(net483),
    .B(_04427_));
 sg13g2_o21ai_1 _10680_ (.B1(_04429_),
    .Y(_00500_),
    .A1(_04292_),
    .A2(net2708));
 sg13g2_nand2_1 _10681_ (.Y(_04430_),
    .A(net428),
    .B(_04427_));
 sg13g2_o21ai_1 _10682_ (.B1(_04430_),
    .Y(_00501_),
    .A1(_04295_),
    .A2(net2710));
 sg13g2_nand2_1 _10683_ (.Y(_04431_),
    .A(net226),
    .B(_04427_));
 sg13g2_o21ai_1 _10684_ (.B1(_04431_),
    .Y(_00502_),
    .A1(_04298_),
    .A2(net2710));
 sg13g2_nand2_1 _10685_ (.Y(_04432_),
    .A(net228),
    .B(_04427_));
 sg13g2_o21ai_1 _10686_ (.B1(_04432_),
    .Y(_00503_),
    .A1(_04301_),
    .A2(net2706));
 sg13g2_nand2_1 _10687_ (.Y(_04433_),
    .A(net644),
    .B(_04427_));
 sg13g2_o21ai_1 _10688_ (.B1(_04433_),
    .Y(_00504_),
    .A1(_04304_),
    .A2(net2710));
 sg13g2_nand2_1 _10689_ (.Y(_04434_),
    .A(net471),
    .B(_04427_));
 sg13g2_o21ai_1 _10690_ (.B1(_04434_),
    .Y(_00505_),
    .A1(_04307_),
    .A2(net2709));
 sg13g2_nand2_1 _10691_ (.Y(_04435_),
    .A(net295),
    .B(_04427_));
 sg13g2_o21ai_1 _10692_ (.B1(_04435_),
    .Y(_00506_),
    .A1(_04310_),
    .A2(net2709));
 sg13g2_nand4_1 _10693_ (.B(net3151),
    .C(net2929),
    .A(net3148),
    .Y(_04436_),
    .D(net2715));
 sg13g2_nand2_1 _10694_ (.Y(_04437_),
    .A(net619),
    .B(_04436_));
 sg13g2_o21ai_1 _10695_ (.B1(_04437_),
    .Y(_00507_),
    .A1(_04316_),
    .A2(net2707));
 sg13g2_nand2_1 _10696_ (.Y(_04438_),
    .A(net506),
    .B(_04436_));
 sg13g2_o21ai_1 _10697_ (.B1(_04438_),
    .Y(_00508_),
    .A1(_04319_),
    .A2(net2707));
 sg13g2_nand2_1 _10698_ (.Y(_04439_),
    .A(net390),
    .B(_04436_));
 sg13g2_o21ai_1 _10699_ (.B1(_04439_),
    .Y(_00509_),
    .A1(_04322_),
    .A2(net2706));
 sg13g2_nand2_1 _10700_ (.Y(_04440_),
    .A(net294),
    .B(_04436_));
 sg13g2_o21ai_1 _10701_ (.B1(_04440_),
    .Y(_00510_),
    .A1(_04325_),
    .A2(net2708));
 sg13g2_nand2_1 _10702_ (.Y(_04441_),
    .A(net271),
    .B(_04436_));
 sg13g2_o21ai_1 _10703_ (.B1(_04441_),
    .Y(_00511_),
    .A1(_04328_),
    .A2(net2706));
 sg13g2_nand2_1 _10704_ (.Y(_04442_),
    .A(net304),
    .B(_04436_));
 sg13g2_o21ai_1 _10705_ (.B1(_04442_),
    .Y(_00512_),
    .A1(_04331_),
    .A2(net2707));
 sg13g2_nand2_1 _10706_ (.Y(_04443_),
    .A(net267),
    .B(_04436_));
 sg13g2_o21ai_1 _10707_ (.B1(_04443_),
    .Y(_00513_),
    .A1(_04334_),
    .A2(net2706));
 sg13g2_nand2_1 _10708_ (.Y(_04444_),
    .A(net251),
    .B(_04436_));
 sg13g2_o21ai_1 _10709_ (.B1(_04444_),
    .Y(_00514_),
    .A1(_04337_),
    .A2(net2711));
 sg13g2_nor2_1 _10710_ (.A(\u_toplayer.u_layer2.neuron_index[4] ),
    .B(_04173_),
    .Y(_04445_));
 sg13g2_nand2_2 _10711_ (.Y(_04446_),
    .A(_03739_),
    .B(_04445_));
 sg13g2_nand2_1 _10712_ (.Y(_04447_),
    .A(net810),
    .B(_04446_));
 sg13g2_o21ai_1 _10713_ (.B1(_04447_),
    .Y(_00515_),
    .A1(_04342_),
    .A2(net2707));
 sg13g2_nand2_1 _10714_ (.Y(_04448_),
    .A(net579),
    .B(_04446_));
 sg13g2_o21ai_1 _10715_ (.B1(_04448_),
    .Y(_00516_),
    .A1(_04345_),
    .A2(net2707));
 sg13g2_nand2_1 _10716_ (.Y(_04449_),
    .A(net664),
    .B(_04446_));
 sg13g2_o21ai_1 _10717_ (.B1(_04449_),
    .Y(_00517_),
    .A1(_04348_),
    .A2(net2709));
 sg13g2_nand2_1 _10718_ (.Y(_04450_),
    .A(net273),
    .B(_04446_));
 sg13g2_o21ai_1 _10719_ (.B1(_04450_),
    .Y(_00518_),
    .A1(_04351_),
    .A2(net2709));
 sg13g2_nand2_1 _10720_ (.Y(_04451_),
    .A(net819),
    .B(_04446_));
 sg13g2_o21ai_1 _10721_ (.B1(_04451_),
    .Y(_00519_),
    .A1(_04354_),
    .A2(net2706));
 sg13g2_nand2_1 _10722_ (.Y(_04452_),
    .A(net256),
    .B(_04446_));
 sg13g2_o21ai_1 _10723_ (.B1(_04452_),
    .Y(_00520_),
    .A1(_04357_),
    .A2(net2707));
 sg13g2_nand2_1 _10724_ (.Y(_04453_),
    .A(net230),
    .B(_04446_));
 sg13g2_o21ai_1 _10725_ (.B1(_04453_),
    .Y(_00521_),
    .A1(_04360_),
    .A2(net2711));
 sg13g2_nand2_1 _10726_ (.Y(_04454_),
    .A(net225),
    .B(_04446_));
 sg13g2_o21ai_1 _10727_ (.B1(_04454_),
    .Y(_00522_),
    .A1(_04363_),
    .A2(net2706));
 sg13g2_nand2_2 _10728_ (.Y(_04455_),
    .A(\u_toplayer.u_layer2.neuron_index[4] ),
    .B(net2714));
 sg13g2_nand2_1 _10729_ (.Y(_04456_),
    .A(net334),
    .B(_04455_));
 sg13g2_o21ai_1 _10730_ (.B1(_04456_),
    .Y(_00523_),
    .A1(_04367_),
    .A2(net2705));
 sg13g2_nand2_1 _10731_ (.Y(_04457_),
    .A(net870),
    .B(_04455_));
 sg13g2_o21ai_1 _10732_ (.B1(_04457_),
    .Y(_00524_),
    .A1(_04370_),
    .A2(net2705));
 sg13g2_nand2_1 _10733_ (.Y(_04458_),
    .A(net661),
    .B(_04455_));
 sg13g2_o21ai_1 _10734_ (.B1(_04458_),
    .Y(_00525_),
    .A1(_04373_),
    .A2(net2705));
 sg13g2_nand2_1 _10735_ (.Y(_04459_),
    .A(net620),
    .B(_04455_));
 sg13g2_o21ai_1 _10736_ (.B1(_04459_),
    .Y(_00526_),
    .A1(_04376_),
    .A2(net2705));
 sg13g2_nand2_1 _10737_ (.Y(_04460_),
    .A(net663),
    .B(_04455_));
 sg13g2_o21ai_1 _10738_ (.B1(_04460_),
    .Y(_00527_),
    .A1(_04379_),
    .A2(net2705));
 sg13g2_nand2_1 _10739_ (.Y(_04461_),
    .A(net706),
    .B(_04455_));
 sg13g2_o21ai_1 _10740_ (.B1(_04461_),
    .Y(_00528_),
    .A1(_04382_),
    .A2(net2705));
 sg13g2_nand2_1 _10741_ (.Y(_04462_),
    .A(net814),
    .B(_04455_));
 sg13g2_o21ai_1 _10742_ (.B1(_04462_),
    .Y(_00529_),
    .A1(_04385_),
    .A2(net2705));
 sg13g2_nand2_1 _10743_ (.Y(_04463_),
    .A(net407),
    .B(_04455_));
 sg13g2_o21ai_1 _10744_ (.B1(_04463_),
    .Y(_00530_),
    .A1(_04388_),
    .A2(net2705));
 sg13g2_nor2_2 _10745_ (.A(_04167_),
    .B(_04173_),
    .Y(_04464_));
 sg13g2_nand2_2 _10746_ (.Y(_04465_),
    .A(_04171_),
    .B(net2712));
 sg13g2_nand2_1 _10747_ (.Y(_04466_),
    .A(net532),
    .B(_04465_));
 sg13g2_o21ai_1 _10748_ (.B1(_04466_),
    .Y(_00531_),
    .A1(net2806),
    .A2(_04181_));
 sg13g2_nand2_1 _10749_ (.Y(_04467_),
    .A(net523),
    .B(_04465_));
 sg13g2_o21ai_1 _10750_ (.B1(_04467_),
    .Y(_00532_),
    .A1(net2807),
    .A2(_04185_));
 sg13g2_nand2_1 _10751_ (.Y(_04468_),
    .A(net368),
    .B(_04465_));
 sg13g2_o21ai_1 _10752_ (.B1(_04468_),
    .Y(_00533_),
    .A1(net2805),
    .A2(_04188_));
 sg13g2_nand2_1 _10753_ (.Y(_04469_),
    .A(net637),
    .B(_04465_));
 sg13g2_o21ai_1 _10754_ (.B1(_04469_),
    .Y(_00534_),
    .A1(net2807),
    .A2(_04191_));
 sg13g2_nand2_1 _10755_ (.Y(_04470_),
    .A(net647),
    .B(_04465_));
 sg13g2_o21ai_1 _10756_ (.B1(_04470_),
    .Y(_00535_),
    .A1(net2807),
    .A2(_04194_));
 sg13g2_nand2_1 _10757_ (.Y(_04471_),
    .A(net560),
    .B(_04465_));
 sg13g2_o21ai_1 _10758_ (.B1(_04471_),
    .Y(_00536_),
    .A1(net2806),
    .A2(_04197_));
 sg13g2_nand2_1 _10759_ (.Y(_04472_),
    .A(net533),
    .B(_04465_));
 sg13g2_o21ai_1 _10760_ (.B1(_04472_),
    .Y(_00537_),
    .A1(net2806),
    .A2(_04200_));
 sg13g2_nand2_1 _10761_ (.Y(_04473_),
    .A(net703),
    .B(_04465_));
 sg13g2_o21ai_1 _10762_ (.B1(_04473_),
    .Y(_00538_),
    .A1(net2805),
    .A2(_04203_));
 sg13g2_nand2_2 _10763_ (.Y(_04474_),
    .A(_04205_),
    .B(net2712));
 sg13g2_nand2_1 _10764_ (.Y(_04475_),
    .A(net858),
    .B(_04474_));
 sg13g2_o21ai_1 _10765_ (.B1(_04475_),
    .Y(_00539_),
    .A1(net2803),
    .A2(_04209_));
 sg13g2_nand2_1 _10766_ (.Y(_04476_),
    .A(net472),
    .B(_04474_));
 sg13g2_o21ai_1 _10767_ (.B1(_04476_),
    .Y(_00540_),
    .A1(net2807),
    .A2(_04212_));
 sg13g2_nand2_1 _10768_ (.Y(_04477_),
    .A(net372),
    .B(_04474_));
 sg13g2_o21ai_1 _10769_ (.B1(_04477_),
    .Y(_00541_),
    .A1(net2804),
    .A2(_04215_));
 sg13g2_nand2_1 _10770_ (.Y(_04478_),
    .A(net614),
    .B(_04474_));
 sg13g2_o21ai_1 _10771_ (.B1(_04478_),
    .Y(_00542_),
    .A1(net2807),
    .A2(_04218_));
 sg13g2_nand2_1 _10772_ (.Y(_04479_),
    .A(net643),
    .B(_04474_));
 sg13g2_o21ai_1 _10773_ (.B1(_04479_),
    .Y(_00543_),
    .A1(net2807),
    .A2(_04221_));
 sg13g2_nand2_1 _10774_ (.Y(_04480_),
    .A(net684),
    .B(_04474_));
 sg13g2_o21ai_1 _10775_ (.B1(_04480_),
    .Y(_00544_),
    .A1(net2804),
    .A2(_04224_));
 sg13g2_nand2_1 _10776_ (.Y(_04481_),
    .A(net356),
    .B(_04474_));
 sg13g2_o21ai_1 _10777_ (.B1(_04481_),
    .Y(_00545_),
    .A1(net2803),
    .A2(_04227_));
 sg13g2_nand2_1 _10778_ (.Y(_04482_),
    .A(net641),
    .B(_04474_));
 sg13g2_o21ai_1 _10779_ (.B1(_04482_),
    .Y(_00546_),
    .A1(net2803),
    .A2(_04230_));
 sg13g2_nand2_2 _10780_ (.Y(_04483_),
    .A(_04232_),
    .B(net2712));
 sg13g2_nand2_1 _10781_ (.Y(_04484_),
    .A(net880),
    .B(_04483_));
 sg13g2_o21ai_1 _10782_ (.B1(_04484_),
    .Y(_00547_),
    .A1(net2803),
    .A2(_04236_));
 sg13g2_nand2_1 _10783_ (.Y(_04485_),
    .A(net360),
    .B(_04483_));
 sg13g2_o21ai_1 _10784_ (.B1(_04485_),
    .Y(_00548_),
    .A1(net2803),
    .A2(_04239_));
 sg13g2_nand2_1 _10785_ (.Y(_04486_),
    .A(net176),
    .B(_04483_));
 sg13g2_o21ai_1 _10786_ (.B1(_04486_),
    .Y(_00549_),
    .A1(net2804),
    .A2(_04242_));
 sg13g2_nand2_1 _10787_ (.Y(_04487_),
    .A(net221),
    .B(_04483_));
 sg13g2_o21ai_1 _10788_ (.B1(_04487_),
    .Y(_00550_),
    .A1(net2804),
    .A2(_04245_));
 sg13g2_nand2_1 _10789_ (.Y(_04488_),
    .A(net604),
    .B(_04483_));
 sg13g2_o21ai_1 _10790_ (.B1(_04488_),
    .Y(_00551_),
    .A1(net2803),
    .A2(_04248_));
 sg13g2_nand2_1 _10791_ (.Y(_04489_),
    .A(net773),
    .B(_04483_));
 sg13g2_o21ai_1 _10792_ (.B1(_04489_),
    .Y(_00552_),
    .A1(net2804),
    .A2(_04251_));
 sg13g2_nand2_1 _10793_ (.Y(_04490_),
    .A(net751),
    .B(_04483_));
 sg13g2_o21ai_1 _10794_ (.B1(_04490_),
    .Y(_00553_),
    .A1(net2803),
    .A2(_04254_));
 sg13g2_nand2_1 _10795_ (.Y(_04491_),
    .A(net593),
    .B(_04483_));
 sg13g2_o21ai_1 _10796_ (.B1(_04491_),
    .Y(_00554_),
    .A1(net2803),
    .A2(_04257_));
 sg13g2_nand2_2 _10797_ (.Y(_04492_),
    .A(_04259_),
    .B(net2713));
 sg13g2_nand2_1 _10798_ (.Y(_04493_),
    .A(net767),
    .B(_04492_));
 sg13g2_o21ai_1 _10799_ (.B1(_04493_),
    .Y(_00555_),
    .A1(net2810),
    .A2(_04263_));
 sg13g2_nand2_1 _10800_ (.Y(_04494_),
    .A(net636),
    .B(_04492_));
 sg13g2_o21ai_1 _10801_ (.B1(_04494_),
    .Y(_00556_),
    .A1(net2811),
    .A2(_04266_));
 sg13g2_nand2_1 _10802_ (.Y(_04495_),
    .A(net435),
    .B(_04492_));
 sg13g2_o21ai_1 _10803_ (.B1(_04495_),
    .Y(_00557_),
    .A1(net2811),
    .A2(_04269_));
 sg13g2_nand2_1 _10804_ (.Y(_04496_),
    .A(net600),
    .B(_04492_));
 sg13g2_o21ai_1 _10805_ (.B1(_04496_),
    .Y(_00558_),
    .A1(net2811),
    .A2(_04272_));
 sg13g2_nand2_1 _10806_ (.Y(_04497_),
    .A(net310),
    .B(_04492_));
 sg13g2_o21ai_1 _10807_ (.B1(_04497_),
    .Y(_00559_),
    .A1(net2811),
    .A2(_04275_));
 sg13g2_nand2_1 _10808_ (.Y(_04498_),
    .A(net314),
    .B(_04492_));
 sg13g2_o21ai_1 _10809_ (.B1(_04498_),
    .Y(_00560_),
    .A1(net2810),
    .A2(_04278_));
 sg13g2_nand2_1 _10810_ (.Y(_04499_),
    .A(net336),
    .B(_04492_));
 sg13g2_o21ai_1 _10811_ (.B1(_04499_),
    .Y(_00561_),
    .A1(net2808),
    .A2(_04281_));
 sg13g2_nand2_1 _10812_ (.Y(_04500_),
    .A(net528),
    .B(_04492_));
 sg13g2_o21ai_1 _10813_ (.B1(_04500_),
    .Y(_00562_),
    .A1(net2810),
    .A2(_04284_));
 sg13g2_nand2_2 _10814_ (.Y(_04501_),
    .A(_04286_),
    .B(net2713));
 sg13g2_nand2_1 _10815_ (.Y(_04502_),
    .A(net174),
    .B(_04501_));
 sg13g2_o21ai_1 _10816_ (.B1(_04502_),
    .Y(_00563_),
    .A1(net2810),
    .A2(_04290_));
 sg13g2_nand2_1 _10817_ (.Y(_04503_),
    .A(net653),
    .B(_04501_));
 sg13g2_o21ai_1 _10818_ (.B1(_04503_),
    .Y(_00564_),
    .A1(net2811),
    .A2(_04293_));
 sg13g2_nand2_1 _10819_ (.Y(_04504_),
    .A(net828),
    .B(_04501_));
 sg13g2_o21ai_1 _10820_ (.B1(_04504_),
    .Y(_00565_),
    .A1(net2810),
    .A2(_04296_));
 sg13g2_nand2_1 _10821_ (.Y(_04505_),
    .A(net776),
    .B(_04501_));
 sg13g2_o21ai_1 _10822_ (.B1(_04505_),
    .Y(_00566_),
    .A1(net2811),
    .A2(_04299_));
 sg13g2_nand2_1 _10823_ (.Y(_04506_),
    .A(net696),
    .B(_04501_));
 sg13g2_o21ai_1 _10824_ (.B1(_04506_),
    .Y(_00567_),
    .A1(net2811),
    .A2(_04302_));
 sg13g2_nand2_1 _10825_ (.Y(_04507_),
    .A(net507),
    .B(_04501_));
 sg13g2_o21ai_1 _10826_ (.B1(_04507_),
    .Y(_00568_),
    .A1(net2810),
    .A2(_04305_));
 sg13g2_nand2_1 _10827_ (.Y(_04508_),
    .A(net484),
    .B(_04501_));
 sg13g2_o21ai_1 _10828_ (.B1(_04508_),
    .Y(_00569_),
    .A1(net2810),
    .A2(_04308_));
 sg13g2_nand2_1 _10829_ (.Y(_04509_),
    .A(net621),
    .B(_04501_));
 sg13g2_o21ai_1 _10830_ (.B1(_04509_),
    .Y(_00570_),
    .A1(net2810),
    .A2(_04311_));
 sg13g2_nand2_2 _10831_ (.Y(_04510_),
    .A(_04313_),
    .B(net2712));
 sg13g2_nand2_1 _10832_ (.Y(_04511_),
    .A(net630),
    .B(_04510_));
 sg13g2_o21ai_1 _10833_ (.B1(_04511_),
    .Y(_00571_),
    .A1(net2808),
    .A2(_04317_));
 sg13g2_nand2_1 _10834_ (.Y(_04512_),
    .A(net796),
    .B(_04510_));
 sg13g2_o21ai_1 _10835_ (.B1(_04512_),
    .Y(_00572_),
    .A1(net2809),
    .A2(_04320_));
 sg13g2_nand2_1 _10836_ (.Y(_04513_),
    .A(net247),
    .B(_04510_));
 sg13g2_o21ai_1 _10837_ (.B1(_04513_),
    .Y(_00573_),
    .A1(net2808),
    .A2(_04323_));
 sg13g2_nand2_1 _10838_ (.Y(_04514_),
    .A(net595),
    .B(_04510_));
 sg13g2_o21ai_1 _10839_ (.B1(_04514_),
    .Y(_00574_),
    .A1(net2809),
    .A2(_04326_));
 sg13g2_nand2_1 _10840_ (.Y(_04515_),
    .A(net585),
    .B(_04510_));
 sg13g2_o21ai_1 _10841_ (.B1(_04515_),
    .Y(_00575_),
    .A1(net2808),
    .A2(_04329_));
 sg13g2_nand2_1 _10842_ (.Y(_04516_),
    .A(net764),
    .B(_04510_));
 sg13g2_o21ai_1 _10843_ (.B1(_04516_),
    .Y(_00576_),
    .A1(net2805),
    .A2(_04332_));
 sg13g2_nand2_1 _10844_ (.Y(_04517_),
    .A(net642),
    .B(_04510_));
 sg13g2_o21ai_1 _10845_ (.B1(_04517_),
    .Y(_00577_),
    .A1(net2805),
    .A2(_04335_));
 sg13g2_nand2_1 _10846_ (.Y(_04518_),
    .A(net410),
    .B(_04510_));
 sg13g2_o21ai_1 _10847_ (.B1(_04518_),
    .Y(_00578_),
    .A1(net2805),
    .A2(_04338_));
 sg13g2_nand2_2 _10848_ (.Y(_04519_),
    .A(_04339_),
    .B(net2712));
 sg13g2_nand2_1 _10849_ (.Y(_04520_),
    .A(net203),
    .B(_04519_));
 sg13g2_o21ai_1 _10850_ (.B1(_04520_),
    .Y(_00579_),
    .A1(net2808),
    .A2(_04343_));
 sg13g2_nand2_1 _10851_ (.Y(_04521_),
    .A(net191),
    .B(_04519_));
 sg13g2_o21ai_1 _10852_ (.B1(_04521_),
    .Y(_00580_),
    .A1(net2808),
    .A2(_04346_));
 sg13g2_nand2_1 _10853_ (.Y(_04522_),
    .A(net362),
    .B(_04519_));
 sg13g2_o21ai_1 _10854_ (.B1(_04522_),
    .Y(_00581_),
    .A1(net2808),
    .A2(_04349_));
 sg13g2_nand2_1 _10855_ (.Y(_04523_),
    .A(net277),
    .B(_04519_));
 sg13g2_o21ai_1 _10856_ (.B1(_04523_),
    .Y(_00582_),
    .A1(net2809),
    .A2(_04352_));
 sg13g2_nand2_1 _10857_ (.Y(_04524_),
    .A(net405),
    .B(_04519_));
 sg13g2_o21ai_1 _10858_ (.B1(_04524_),
    .Y(_00583_),
    .A1(net2808),
    .A2(_04355_));
 sg13g2_nand2_1 _10859_ (.Y(_04525_),
    .A(net257),
    .B(_04519_));
 sg13g2_o21ai_1 _10860_ (.B1(_04525_),
    .Y(_00584_),
    .A1(net2805),
    .A2(_04358_));
 sg13g2_nand2_1 _10861_ (.Y(_04526_),
    .A(net353),
    .B(_04519_));
 sg13g2_o21ai_1 _10862_ (.B1(_04526_),
    .Y(_00585_),
    .A1(net2805),
    .A2(_04361_));
 sg13g2_nand2_1 _10863_ (.Y(_04527_),
    .A(net535),
    .B(_04519_));
 sg13g2_o21ai_1 _10864_ (.B1(_04527_),
    .Y(_00586_),
    .A1(net2805),
    .A2(_04364_));
 sg13g2_nand3_1 _10865_ (.B(net2948),
    .C(net2713),
    .A(net3147),
    .Y(_04528_));
 sg13g2_nand2_1 _10866_ (.Y(_04529_),
    .A(net697),
    .B(_04528_));
 sg13g2_o21ai_1 _10867_ (.B1(_04529_),
    .Y(_00587_),
    .A1(net2812),
    .A2(_04368_));
 sg13g2_nand2_1 _10868_ (.Y(_04530_),
    .A(net434),
    .B(_04528_));
 sg13g2_o21ai_1 _10869_ (.B1(_04530_),
    .Y(_00588_),
    .A1(net2813),
    .A2(_04371_));
 sg13g2_nand2_1 _10870_ (.Y(_04531_),
    .A(net674),
    .B(_04528_));
 sg13g2_o21ai_1 _10871_ (.B1(_04531_),
    .Y(_00589_),
    .A1(net2813),
    .A2(_04374_));
 sg13g2_nand2_1 _10872_ (.Y(_04532_),
    .A(net710),
    .B(_04528_));
 sg13g2_o21ai_1 _10873_ (.B1(_04532_),
    .Y(_00590_),
    .A1(net2813),
    .A2(_04377_));
 sg13g2_nand2_1 _10874_ (.Y(_04533_),
    .A(net547),
    .B(_04528_));
 sg13g2_o21ai_1 _10875_ (.B1(_04533_),
    .Y(_00591_),
    .A1(net2812),
    .A2(_04380_));
 sg13g2_nand2_1 _10876_ (.Y(_04534_),
    .A(net503),
    .B(_04528_));
 sg13g2_o21ai_1 _10877_ (.B1(_04534_),
    .Y(_00592_),
    .A1(net2812),
    .A2(_04383_));
 sg13g2_nand2_1 _10878_ (.Y(_04535_),
    .A(net316),
    .B(_04528_));
 sg13g2_o21ai_1 _10879_ (.B1(_04535_),
    .Y(_00593_),
    .A1(net2812),
    .A2(_04386_));
 sg13g2_nand2_1 _10880_ (.Y(_04536_),
    .A(net563),
    .B(_04528_));
 sg13g2_o21ai_1 _10881_ (.B1(_04536_),
    .Y(_00594_),
    .A1(net2812),
    .A2(_04389_));
 sg13g2_nand3_1 _10882_ (.B(net2924),
    .C(net2713),
    .A(net3147),
    .Y(_04537_));
 sg13g2_nand2_1 _10883_ (.Y(_04538_),
    .A(net236),
    .B(_04537_));
 sg13g2_nand2_1 _10884_ (.Y(_04539_),
    .A(_04178_),
    .B(net2712));
 sg13g2_o21ai_1 _10885_ (.B1(_04538_),
    .Y(_00595_),
    .A1(_04180_),
    .A2(net2695));
 sg13g2_nand2_1 _10886_ (.Y(_04540_),
    .A(net444),
    .B(_04537_));
 sg13g2_o21ai_1 _10887_ (.B1(_04540_),
    .Y(_00596_),
    .A1(_04184_),
    .A2(net2695));
 sg13g2_nand2_1 _10888_ (.Y(_04541_),
    .A(net204),
    .B(_04537_));
 sg13g2_o21ai_1 _10889_ (.B1(_04541_),
    .Y(_00597_),
    .A1(_04187_),
    .A2(net2695));
 sg13g2_nand2_1 _10890_ (.Y(_04542_),
    .A(net716),
    .B(_04537_));
 sg13g2_o21ai_1 _10891_ (.B1(_04542_),
    .Y(_00598_),
    .A1(_04190_),
    .A2(net2695));
 sg13g2_nand2_1 _10892_ (.Y(_04543_),
    .A(net757),
    .B(_04537_));
 sg13g2_o21ai_1 _10893_ (.B1(_04543_),
    .Y(_00599_),
    .A1(_04193_),
    .A2(net2694));
 sg13g2_nand2_1 _10894_ (.Y(_04544_),
    .A(net393),
    .B(_04537_));
 sg13g2_o21ai_1 _10895_ (.B1(_04544_),
    .Y(_00600_),
    .A1(_04196_),
    .A2(net2695));
 sg13g2_nand2_1 _10896_ (.Y(_04545_),
    .A(net318),
    .B(_04537_));
 sg13g2_o21ai_1 _10897_ (.B1(_04545_),
    .Y(_00601_),
    .A1(_04199_),
    .A2(net2694));
 sg13g2_nand2_1 _10898_ (.Y(_04546_),
    .A(net707),
    .B(_04537_));
 sg13g2_o21ai_1 _10899_ (.B1(_04546_),
    .Y(_00602_),
    .A1(_04202_),
    .A2(net2701));
 sg13g2_nand3_1 _10900_ (.B(net2876),
    .C(net2712),
    .A(net3146),
    .Y(_04547_));
 sg13g2_nand2_1 _10901_ (.Y(_04548_),
    .A(net722),
    .B(_04547_));
 sg13g2_o21ai_1 _10902_ (.B1(_04548_),
    .Y(_00603_),
    .A1(_04208_),
    .A2(net2692));
 sg13g2_nand2_1 _10903_ (.Y(_04549_),
    .A(net650),
    .B(_04547_));
 sg13g2_o21ai_1 _10904_ (.B1(_04549_),
    .Y(_00604_),
    .A1(_04211_),
    .A2(net2692));
 sg13g2_nand2_1 _10905_ (.Y(_04550_),
    .A(net301),
    .B(_04547_));
 sg13g2_o21ai_1 _10906_ (.B1(_04550_),
    .Y(_00605_),
    .A1(_04214_),
    .A2(net2701));
 sg13g2_nand2_1 _10907_ (.Y(_04551_),
    .A(net740),
    .B(_04547_));
 sg13g2_o21ai_1 _10908_ (.B1(_04551_),
    .Y(_00606_),
    .A1(_04217_),
    .A2(net2692));
 sg13g2_nand2_1 _10909_ (.Y(_04552_),
    .A(net350),
    .B(_04547_));
 sg13g2_o21ai_1 _10910_ (.B1(_04552_),
    .Y(_00607_),
    .A1(_04220_),
    .A2(net2693));
 sg13g2_nand2_1 _10911_ (.Y(_04553_),
    .A(net487),
    .B(_04547_));
 sg13g2_o21ai_1 _10912_ (.B1(_04553_),
    .Y(_00608_),
    .A1(_04223_),
    .A2(net2692));
 sg13g2_nand2_1 _10913_ (.Y(_04554_),
    .A(net834),
    .B(_04547_));
 sg13g2_o21ai_1 _10914_ (.B1(_04554_),
    .Y(_00609_),
    .A1(_04226_),
    .A2(net2693));
 sg13g2_nand2_1 _10915_ (.Y(_04555_),
    .A(net768),
    .B(_04547_));
 sg13g2_o21ai_1 _10916_ (.B1(_04555_),
    .Y(_00610_),
    .A1(_04229_),
    .A2(net2693));
 sg13g2_nand3_1 _10917_ (.B(net2922),
    .C(net2712),
    .A(net3146),
    .Y(_04556_));
 sg13g2_nand2_1 _10918_ (.Y(_04557_),
    .A(net391),
    .B(_04556_));
 sg13g2_o21ai_1 _10919_ (.B1(_04557_),
    .Y(_00611_),
    .A1(_04235_),
    .A2(net2692));
 sg13g2_nand2_1 _10920_ (.Y(_04558_),
    .A(net268),
    .B(_04556_));
 sg13g2_o21ai_1 _10921_ (.B1(_04558_),
    .Y(_00612_),
    .A1(_04238_),
    .A2(net2692));
 sg13g2_nand2_1 _10922_ (.Y(_04559_),
    .A(net163),
    .B(_04556_));
 sg13g2_o21ai_1 _10923_ (.B1(_04559_),
    .Y(_00613_),
    .A1(_04241_),
    .A2(net2692));
 sg13g2_nand2_1 _10924_ (.Y(_04560_),
    .A(net662),
    .B(_04556_));
 sg13g2_o21ai_1 _10925_ (.B1(_04560_),
    .Y(_00614_),
    .A1(_04244_),
    .A2(net2693));
 sg13g2_nand2_1 _10926_ (.Y(_04561_),
    .A(net384),
    .B(_04556_));
 sg13g2_o21ai_1 _10927_ (.B1(_04561_),
    .Y(_00615_),
    .A1(_04247_),
    .A2(net2693));
 sg13g2_nand2_1 _10928_ (.Y(_04562_),
    .A(net223),
    .B(_04556_));
 sg13g2_o21ai_1 _10929_ (.B1(_04562_),
    .Y(_00616_),
    .A1(_04250_),
    .A2(net2692));
 sg13g2_nand2_1 _10930_ (.Y(_04563_),
    .A(net805),
    .B(_04556_));
 sg13g2_o21ai_1 _10931_ (.B1(_04563_),
    .Y(_00617_),
    .A1(_04253_),
    .A2(net2693));
 sg13g2_nand2_1 _10932_ (.Y(_04564_),
    .A(net411),
    .B(_04556_));
 sg13g2_o21ai_1 _10933_ (.B1(_04564_),
    .Y(_00618_),
    .A1(_04256_),
    .A2(net2693));
 sg13g2_nand3_1 _10934_ (.B(net2920),
    .C(net2713),
    .A(net3147),
    .Y(_04565_));
 sg13g2_nand2_1 _10935_ (.Y(_04566_),
    .A(net509),
    .B(_04565_));
 sg13g2_o21ai_1 _10936_ (.B1(_04566_),
    .Y(_00619_),
    .A1(_04262_),
    .A2(net2695));
 sg13g2_nand2_1 _10937_ (.Y(_04567_),
    .A(net550),
    .B(_04565_));
 sg13g2_o21ai_1 _10938_ (.B1(_04567_),
    .Y(_00620_),
    .A1(_04265_),
    .A2(net2696));
 sg13g2_nand2_1 _10939_ (.Y(_04568_),
    .A(net332),
    .B(_04565_));
 sg13g2_o21ai_1 _10940_ (.B1(_04568_),
    .Y(_00621_),
    .A1(_04268_),
    .A2(net2699));
 sg13g2_nand2_1 _10941_ (.Y(_04569_),
    .A(net693),
    .B(_04565_));
 sg13g2_o21ai_1 _10942_ (.B1(_04569_),
    .Y(_00622_),
    .A1(_04271_),
    .A2(net2699));
 sg13g2_nand2_1 _10943_ (.Y(_04570_),
    .A(net656),
    .B(_04565_));
 sg13g2_o21ai_1 _10944_ (.B1(_04570_),
    .Y(_00623_),
    .A1(_04274_),
    .A2(net2697));
 sg13g2_nand2_1 _10945_ (.Y(_04571_),
    .A(net522),
    .B(_04565_));
 sg13g2_o21ai_1 _10946_ (.B1(_04571_),
    .Y(_00624_),
    .A1(_04277_),
    .A2(net2700));
 sg13g2_nand2_1 _10947_ (.Y(_04572_),
    .A(net357),
    .B(_04565_));
 sg13g2_o21ai_1 _10948_ (.B1(_04572_),
    .Y(_00625_),
    .A1(_04280_),
    .A2(net2699));
 sg13g2_nand2_1 _10949_ (.Y(_04573_),
    .A(net520),
    .B(_04565_));
 sg13g2_o21ai_1 _10950_ (.B1(_04573_),
    .Y(_00626_),
    .A1(_04283_),
    .A2(net2698));
 sg13g2_nand3_1 _10951_ (.B(net2917),
    .C(net2713),
    .A(net3147),
    .Y(_04574_));
 sg13g2_nand2_1 _10952_ (.Y(_04575_),
    .A(net657),
    .B(_04574_));
 sg13g2_o21ai_1 _10953_ (.B1(_04575_),
    .Y(_00627_),
    .A1(_04289_),
    .A2(net2695));
 sg13g2_nand2_1 _10954_ (.Y(_04576_),
    .A(net479),
    .B(_04574_));
 sg13g2_o21ai_1 _10955_ (.B1(_04576_),
    .Y(_00628_),
    .A1(_04292_),
    .A2(net2695));
 sg13g2_nand2_1 _10956_ (.Y(_04577_),
    .A(net671),
    .B(_04574_));
 sg13g2_o21ai_1 _10957_ (.B1(_04577_),
    .Y(_00629_),
    .A1(_04295_),
    .A2(net2699));
 sg13g2_nand2_1 _10958_ (.Y(_04578_),
    .A(net440),
    .B(_04574_));
 sg13g2_o21ai_1 _10959_ (.B1(_04578_),
    .Y(_00630_),
    .A1(_04298_),
    .A2(net2699));
 sg13g2_nand2_1 _10960_ (.Y(_04579_),
    .A(net302),
    .B(_04574_));
 sg13g2_o21ai_1 _10961_ (.B1(_04579_),
    .Y(_00631_),
    .A1(_04301_),
    .A2(net2697));
 sg13g2_nand2_1 _10962_ (.Y(_04580_),
    .A(net618),
    .B(_04574_));
 sg13g2_o21ai_1 _10963_ (.B1(_04580_),
    .Y(_00632_),
    .A1(_04304_),
    .A2(net2699));
 sg13g2_nand2_1 _10964_ (.Y(_04581_),
    .A(net300),
    .B(_04574_));
 sg13g2_o21ai_1 _10965_ (.B1(_04581_),
    .Y(_00633_),
    .A1(_04307_),
    .A2(net2700));
 sg13g2_nand2_1 _10966_ (.Y(_04582_),
    .A(net323),
    .B(_04574_));
 sg13g2_o21ai_1 _10967_ (.B1(_04582_),
    .Y(_00634_),
    .A1(_04310_),
    .A2(net2697));
 sg13g2_nand4_1 _10968_ (.B(net3151),
    .C(net2929),
    .A(net3148),
    .Y(_04583_),
    .D(net2713));
 sg13g2_nand2_1 _10969_ (.Y(_04584_),
    .A(net728),
    .B(_04583_));
 sg13g2_o21ai_1 _10970_ (.B1(_04584_),
    .Y(_00635_),
    .A1(_04316_),
    .A2(net2694));
 sg13g2_nand2_1 _10971_ (.Y(_04585_),
    .A(net309),
    .B(_04583_));
 sg13g2_o21ai_1 _10972_ (.B1(_04585_),
    .Y(_00636_),
    .A1(_04319_),
    .A2(net2696));
 sg13g2_nand2_1 _10973_ (.Y(_04586_),
    .A(net589),
    .B(_04583_));
 sg13g2_o21ai_1 _10974_ (.B1(_04586_),
    .Y(_00637_),
    .A1(_04322_),
    .A2(net2697));
 sg13g2_nand2_1 _10975_ (.Y(_04587_),
    .A(net583),
    .B(_04583_));
 sg13g2_o21ai_1 _10976_ (.B1(_04587_),
    .Y(_00638_),
    .A1(_04325_),
    .A2(net2694));
 sg13g2_nand2_1 _10977_ (.Y(_04588_),
    .A(net536),
    .B(_04583_));
 sg13g2_o21ai_1 _10978_ (.B1(_04588_),
    .Y(_00639_),
    .A1(_04328_),
    .A2(net2698));
 sg13g2_nand2_1 _10979_ (.Y(_04589_),
    .A(net344),
    .B(_04583_));
 sg13g2_o21ai_1 _10980_ (.B1(_04589_),
    .Y(_00640_),
    .A1(_04331_),
    .A2(net2694));
 sg13g2_nand2_1 _10981_ (.Y(_04590_),
    .A(net459),
    .B(_04583_));
 sg13g2_o21ai_1 _10982_ (.B1(_04590_),
    .Y(_00641_),
    .A1(_04334_),
    .A2(net2697));
 sg13g2_nand2_1 _10983_ (.Y(_04591_),
    .A(net290),
    .B(_04583_));
 sg13g2_o21ai_1 _10984_ (.B1(_04591_),
    .Y(_00642_),
    .A1(_04337_),
    .A2(net2697));
 sg13g2_nand2_1 _10985_ (.Y(_04592_),
    .A(net835),
    .B(_03742_));
 sg13g2_o21ai_1 _10986_ (.B1(_04592_),
    .Y(_00643_),
    .A1(_04342_),
    .A2(net2694));
 sg13g2_nand2_1 _10987_ (.Y(_04593_),
    .A(net475),
    .B(_03742_));
 sg13g2_o21ai_1 _10988_ (.B1(_04593_),
    .Y(_00644_),
    .A1(_04345_),
    .A2(net2694));
 sg13g2_nand2_1 _10989_ (.Y(_04594_),
    .A(net266),
    .B(_03742_));
 sg13g2_o21ai_1 _10990_ (.B1(_04594_),
    .Y(_00645_),
    .A1(_04348_),
    .A2(net2697));
 sg13g2_nand2_1 _10991_ (.Y(_04595_),
    .A(net430),
    .B(_03742_));
 sg13g2_o21ai_1 _10992_ (.B1(_04595_),
    .Y(_00646_),
    .A1(_04351_),
    .A2(net2697));
 sg13g2_nand2_1 _10993_ (.Y(_04596_),
    .A(net324),
    .B(_03742_));
 sg13g2_o21ai_1 _10994_ (.B1(_04596_),
    .Y(_00647_),
    .A1(_04354_),
    .A2(net2698));
 sg13g2_nand2_1 _10995_ (.Y(_04597_),
    .A(net403),
    .B(_03742_));
 sg13g2_o21ai_1 _10996_ (.B1(_04597_),
    .Y(_00648_),
    .A1(_04357_),
    .A2(net2694));
 sg13g2_nand2_1 _10997_ (.Y(_04598_),
    .A(net470),
    .B(_03742_));
 sg13g2_o21ai_1 _10998_ (.B1(_04598_),
    .Y(_00649_),
    .A1(_04360_),
    .A2(net2698));
 sg13g2_nand2_1 _10999_ (.Y(_04599_),
    .A(net660),
    .B(_03742_));
 sg13g2_o21ai_1 _11000_ (.B1(_04599_),
    .Y(_00650_),
    .A1(_04363_),
    .A2(net2698));
 sg13g2_nand3b_1 _11001_ (.B(\u_toplayer.u_layer2.neuron_index[5] ),
    .C(_04165_),
    .Y(_04600_),
    .A_N(\u_toplayer.u_layer2.neuron_index[4] ));
 sg13g2_o21ai_1 _11002_ (.B1(_01024_),
    .Y(_00651_),
    .A1(_01031_),
    .A2(_04600_));
 sg13g2_nand2_2 _11003_ (.Y(_04601_),
    .A(net1156),
    .B(_02646_));
 sg13g2_a21oi_1 _11004_ (.A1(net3268),
    .A2(_01120_),
    .Y(_04602_),
    .B1(net3250));
 sg13g2_o21ai_1 _11005_ (.B1(_04602_),
    .Y(_04603_),
    .A1(net3267),
    .A2(\u_toplayer.reg_layer1[192] ));
 sg13g2_a221oi_1 _11006_ (.B2(\u_toplayer.reg_layer1[208] ),
    .C1(net3239),
    .B1(net2962),
    .A1(\u_toplayer.reg_layer1[216] ),
    .Y(_04604_),
    .A2(net2991));
 sg13g2_nor2b_1 _11007_ (.A(\u_toplayer.reg_layer1[232] ),
    .B_N(net3267),
    .Y(_04605_));
 sg13g2_nor2_1 _11008_ (.A(net3269),
    .B(\u_toplayer.reg_layer1[224] ),
    .Y(_04606_));
 sg13g2_nor3_1 _11009_ (.A(net3251),
    .B(_04605_),
    .C(_04606_),
    .Y(_04607_));
 sg13g2_a221oi_1 _11010_ (.B2(\u_toplayer.reg_layer1[240] ),
    .C1(_04607_),
    .B1(net2961),
    .A1(\u_toplayer.reg_layer1[248] ),
    .Y(_04608_),
    .A2(net2990));
 sg13g2_a22oi_1 _11011_ (.Y(_04609_),
    .B1(_04608_),
    .B2(net3239),
    .A2(_04604_),
    .A1(_04603_));
 sg13g2_nand2_1 _11012_ (.Y(_04610_),
    .A(net3236),
    .B(_04609_));
 sg13g2_nor2b_1 _11013_ (.A(net3262),
    .B_N(\u_toplayer.reg_layer1[128] ),
    .Y(_04611_));
 sg13g2_a21oi_1 _11014_ (.A1(net3260),
    .A2(\u_toplayer.reg_layer1[136] ),
    .Y(_04612_),
    .B1(_04611_));
 sg13g2_a22oi_1 _11015_ (.Y(_04613_),
    .B1(net2956),
    .B2(\u_toplayer.reg_layer1[144] ),
    .A2(net2986),
    .A1(\u_toplayer.reg_layer1[152] ));
 sg13g2_o21ai_1 _11016_ (.B1(_04613_),
    .Y(_04614_),
    .A1(net3248),
    .A2(_04612_));
 sg13g2_nor2_1 _11017_ (.A(net3019),
    .B(net3235),
    .Y(_04615_));
 sg13g2_nand2b_1 _11018_ (.Y(_04616_),
    .B(net3256),
    .A_N(\u_toplayer.reg_layer1[168] ));
 sg13g2_o21ai_1 _11019_ (.B1(_04616_),
    .Y(_04617_),
    .A1(net3256),
    .A2(\u_toplayer.reg_layer1[160] ));
 sg13g2_a22oi_1 _11020_ (.Y(_04618_),
    .B1(net2955),
    .B2(\u_toplayer.reg_layer1[176] ),
    .A2(net2984),
    .A1(\u_toplayer.reg_layer1[184] ));
 sg13g2_o21ai_1 _11021_ (.B1(_04618_),
    .Y(_04619_),
    .A1(net3243),
    .A2(_04617_));
 sg13g2_a22oi_1 _11022_ (.Y(_04620_),
    .B1(net2914),
    .B2(_04619_),
    .A2(_04614_),
    .A1(net2996));
 sg13g2_nand3_1 _11023_ (.B(_04610_),
    .C(_04620_),
    .A(net3234),
    .Y(_04621_));
 sg13g2_a21oi_1 _11024_ (.A1(net3267),
    .A2(_01119_),
    .Y(_04622_),
    .B1(net3250));
 sg13g2_o21ai_1 _11025_ (.B1(_04622_),
    .Y(_04623_),
    .A1(net3267),
    .A2(\u_toplayer.reg_layer1[96] ));
 sg13g2_a22oi_1 _11026_ (.Y(_04624_),
    .B1(net2960),
    .B2(\u_toplayer.reg_layer1[112] ),
    .A2(net2990),
    .A1(\u_toplayer.reg_layer1[120] ));
 sg13g2_nand3_1 _11027_ (.B(_04623_),
    .C(_04624_),
    .A(net3241),
    .Y(_04625_));
 sg13g2_a21oi_1 _11028_ (.A1(net3267),
    .A2(_01118_),
    .Y(_04626_),
    .B1(net3250));
 sg13g2_o21ai_1 _11029_ (.B1(_04626_),
    .Y(_04627_),
    .A1(net3267),
    .A2(\u_toplayer.reg_layer1[64] ));
 sg13g2_a22oi_1 _11030_ (.Y(_04628_),
    .B1(net2962),
    .B2(\u_toplayer.reg_layer1[80] ),
    .A2(net2991),
    .A1(\u_toplayer.reg_layer1[88] ));
 sg13g2_nand3_1 _11031_ (.B(_04627_),
    .C(_04628_),
    .A(net3019),
    .Y(_04629_));
 sg13g2_nand3_1 _11032_ (.B(_04625_),
    .C(_04629_),
    .A(net3237),
    .Y(_04630_));
 sg13g2_nor2b_1 _11033_ (.A(net3270),
    .B_N(\u_toplayer.reg_layer1[0] ),
    .Y(_04631_));
 sg13g2_a21oi_1 _11034_ (.A1(net3270),
    .A2(\u_toplayer.reg_layer1[8] ),
    .Y(_04632_),
    .B1(_04631_));
 sg13g2_a22oi_1 _11035_ (.Y(_04633_),
    .B1(net2954),
    .B2(\u_toplayer.reg_layer1[16] ),
    .A2(net2984),
    .A1(\u_toplayer.reg_layer1[24] ));
 sg13g2_o21ai_1 _11036_ (.B1(_04633_),
    .Y(_04634_),
    .A1(net3246),
    .A2(_04632_));
 sg13g2_nand2b_1 _11037_ (.Y(_04635_),
    .B(net3258),
    .A_N(\u_toplayer.reg_layer1[40] ));
 sg13g2_o21ai_1 _11038_ (.B1(_04635_),
    .Y(_04636_),
    .A1(net3256),
    .A2(\u_toplayer.reg_layer1[32] ));
 sg13g2_a22oi_1 _11039_ (.Y(_04637_),
    .B1(net2956),
    .B2(\u_toplayer.reg_layer1[48] ),
    .A2(net2995),
    .A1(\u_toplayer.reg_layer1[56] ));
 sg13g2_o21ai_1 _11040_ (.B1(_04637_),
    .Y(_04638_),
    .A1(net3243),
    .A2(_04636_));
 sg13g2_a221oi_1 _11041_ (.B2(net2915),
    .C1(net3232),
    .B1(_04638_),
    .A1(net2997),
    .Y(_04639_),
    .A2(_04634_));
 sg13g2_a21oi_1 _11042_ (.A1(_04630_),
    .A2(_04639_),
    .Y(_04640_),
    .B1(_04601_));
 sg13g2_a22oi_1 _11043_ (.Y(_04641_),
    .B1(_04621_),
    .B2(_04640_),
    .A2(_02647_),
    .A1(net3094));
 sg13g2_inv_1 _11044_ (.Y(_00652_),
    .A(_04641_));
 sg13g2_a21oi_1 _11045_ (.A1(net3274),
    .A2(_01122_),
    .Y(_04642_),
    .B1(net3249));
 sg13g2_o21ai_1 _11046_ (.B1(_04642_),
    .Y(_04643_),
    .A1(net3266),
    .A2(\u_toplayer.reg_layer1[97] ));
 sg13g2_a22oi_1 _11047_ (.Y(_04644_),
    .B1(net2960),
    .B2(\u_toplayer.reg_layer1[113] ),
    .A2(net2990),
    .A1(\u_toplayer.reg_layer1[121] ));
 sg13g2_nand3_1 _11048_ (.B(_04643_),
    .C(_04644_),
    .A(net3241),
    .Y(_04645_));
 sg13g2_a21oi_1 _11049_ (.A1(net3275),
    .A2(_01121_),
    .Y(_04646_),
    .B1(net3254));
 sg13g2_o21ai_1 _11050_ (.B1(_04646_),
    .Y(_04647_),
    .A1(net3275),
    .A2(\u_toplayer.reg_layer1[65] ));
 sg13g2_a22oi_1 _11051_ (.Y(_04648_),
    .B1(net2964),
    .B2(\u_toplayer.reg_layer1[81] ),
    .A2(net2992),
    .A1(\u_toplayer.reg_layer1[89] ));
 sg13g2_nand3_1 _11052_ (.B(_04647_),
    .C(_04648_),
    .A(net3020),
    .Y(_04649_));
 sg13g2_nand3_1 _11053_ (.B(_04645_),
    .C(_04649_),
    .A(net3237),
    .Y(_04650_));
 sg13g2_nand2b_1 _11054_ (.Y(_04651_),
    .B(net3258),
    .A_N(\u_toplayer.reg_layer1[41] ));
 sg13g2_o21ai_1 _11055_ (.B1(_04651_),
    .Y(_04652_),
    .A1(net3257),
    .A2(\u_toplayer.reg_layer1[33] ));
 sg13g2_a22oi_1 _11056_ (.Y(_04653_),
    .B1(net2955),
    .B2(\u_toplayer.reg_layer1[49] ),
    .A2(net2984),
    .A1(\u_toplayer.reg_layer1[57] ));
 sg13g2_o21ai_1 _11057_ (.B1(_04653_),
    .Y(_04654_),
    .A1(net3243),
    .A2(_04652_));
 sg13g2_nand2b_1 _11058_ (.Y(_04655_),
    .B(net3270),
    .A_N(\u_toplayer.reg_layer1[9] ));
 sg13g2_o21ai_1 _11059_ (.B1(_04655_),
    .Y(_04656_),
    .A1(net3270),
    .A2(\u_toplayer.reg_layer1[1] ));
 sg13g2_a22oi_1 _11060_ (.Y(_04657_),
    .B1(net2958),
    .B2(\u_toplayer.reg_layer1[17] ),
    .A2(net2988),
    .A1(\u_toplayer.reg_layer1[25] ));
 sg13g2_o21ai_1 _11061_ (.B1(_04657_),
    .Y(_04658_),
    .A1(net3246),
    .A2(_04656_));
 sg13g2_a221oi_1 _11062_ (.B2(net2997),
    .C1(net3232),
    .B1(_04658_),
    .A1(_04615_),
    .Y(_04659_),
    .A2(_04654_));
 sg13g2_a21oi_1 _11063_ (.A1(net3274),
    .A2(_01124_),
    .Y(_04660_),
    .B1(net3253));
 sg13g2_o21ai_1 _11064_ (.B1(_04660_),
    .Y(_04661_),
    .A1(net3274),
    .A2(\u_toplayer.reg_layer1[225] ));
 sg13g2_a221oi_1 _11065_ (.B2(\u_toplayer.reg_layer1[241] ),
    .C1(net3019),
    .B1(net2961),
    .A1(\u_toplayer.reg_layer1[249] ),
    .Y(_04662_),
    .A2(net2990));
 sg13g2_a21oi_1 _11066_ (.A1(net3275),
    .A2(_01123_),
    .Y(_04663_),
    .B1(net3254));
 sg13g2_o21ai_1 _11067_ (.B1(_04663_),
    .Y(_04664_),
    .A1(net3275),
    .A2(\u_toplayer.reg_layer1[193] ));
 sg13g2_a221oi_1 _11068_ (.B2(\u_toplayer.reg_layer1[209] ),
    .C1(net3242),
    .B1(net2964),
    .A1(\u_toplayer.reg_layer1[217] ),
    .Y(_04665_),
    .A2(net2992));
 sg13g2_a22oi_1 _11069_ (.Y(_04666_),
    .B1(_04664_),
    .B2(_04665_),
    .A2(_04662_),
    .A1(_04661_));
 sg13g2_nand2_1 _11070_ (.Y(_04667_),
    .A(net3237),
    .B(_04666_));
 sg13g2_nand2b_1 _11071_ (.Y(_04668_),
    .B(net3257),
    .A_N(\u_toplayer.reg_layer1[169] ));
 sg13g2_o21ai_1 _11072_ (.B1(_04668_),
    .Y(_04669_),
    .A1(net3257),
    .A2(\u_toplayer.reg_layer1[161] ));
 sg13g2_a22oi_1 _11073_ (.Y(_04670_),
    .B1(net2955),
    .B2(\u_toplayer.reg_layer1[177] ),
    .A2(net2984),
    .A1(\u_toplayer.reg_layer1[185] ));
 sg13g2_o21ai_1 _11074_ (.B1(_04670_),
    .Y(_04671_),
    .A1(net3243),
    .A2(_04669_));
 sg13g2_nor2b_1 _11075_ (.A(net3260),
    .B_N(\u_toplayer.reg_layer1[129] ),
    .Y(_04672_));
 sg13g2_a21oi_1 _11076_ (.A1(net3260),
    .A2(\u_toplayer.reg_layer1[137] ),
    .Y(_04673_),
    .B1(_04672_));
 sg13g2_a22oi_1 _11077_ (.Y(_04674_),
    .B1(net2958),
    .B2(\u_toplayer.reg_layer1[145] ),
    .A2(net2988),
    .A1(\u_toplayer.reg_layer1[153] ));
 sg13g2_o21ai_1 _11078_ (.B1(_04674_),
    .Y(_04675_),
    .A1(net3247),
    .A2(_04673_));
 sg13g2_a22oi_1 _11079_ (.Y(_04676_),
    .B1(_04675_),
    .B2(net2996),
    .A2(_04671_),
    .A1(net2914));
 sg13g2_and2_1 _11080_ (.A(net3231),
    .B(_04676_),
    .X(_04677_));
 sg13g2_a221oi_1 _11081_ (.B2(_04677_),
    .C1(_04601_),
    .B1(_04667_),
    .A1(_04650_),
    .Y(_04678_),
    .A2(_04659_));
 sg13g2_a21o_1 _11082_ (.A2(_02647_),
    .A1(net3092),
    .B1(_04678_),
    .X(_00653_));
 sg13g2_a21oi_1 _11083_ (.A1(net3266),
    .A2(_01126_),
    .Y(_04679_),
    .B1(net3249));
 sg13g2_o21ai_1 _11084_ (.B1(_04679_),
    .Y(_04680_),
    .A1(net3265),
    .A2(\u_toplayer.reg_layer1[98] ));
 sg13g2_a22oi_1 _11085_ (.Y(_04681_),
    .B1(net2960),
    .B2(\u_toplayer.reg_layer1[114] ),
    .A2(net2987),
    .A1(\u_toplayer.reg_layer1[122] ));
 sg13g2_nand3_1 _11086_ (.B(_04680_),
    .C(_04681_),
    .A(net3240),
    .Y(_04682_));
 sg13g2_a21oi_1 _11087_ (.A1(net3275),
    .A2(_01125_),
    .Y(_04683_),
    .B1(net3254));
 sg13g2_o21ai_1 _11088_ (.B1(_04683_),
    .Y(_04684_),
    .A1(net3275),
    .A2(\u_toplayer.reg_layer1[66] ));
 sg13g2_a22oi_1 _11089_ (.Y(_04685_),
    .B1(net2963),
    .B2(\u_toplayer.reg_layer1[82] ),
    .A2(net2992),
    .A1(\u_toplayer.reg_layer1[90] ));
 sg13g2_nand3_1 _11090_ (.B(_04684_),
    .C(_04685_),
    .A(net3020),
    .Y(_04686_));
 sg13g2_nand3_1 _11091_ (.B(_04682_),
    .C(_04686_),
    .A(net3236),
    .Y(_04687_));
 sg13g2_nand2b_1 _11092_ (.Y(_04688_),
    .B(net3271),
    .A_N(\u_toplayer.reg_layer1[10] ));
 sg13g2_o21ai_1 _11093_ (.B1(_04688_),
    .Y(_04689_),
    .A1(net3271),
    .A2(\u_toplayer.reg_layer1[2] ));
 sg13g2_a22oi_1 _11094_ (.Y(_04690_),
    .B1(net2954),
    .B2(\u_toplayer.reg_layer1[18] ),
    .A2(net2985),
    .A1(\u_toplayer.reg_layer1[26] ));
 sg13g2_o21ai_1 _11095_ (.B1(_04690_),
    .Y(_04691_),
    .A1(net3252),
    .A2(_04689_));
 sg13g2_nand2b_1 _11096_ (.Y(_04692_),
    .B(net3259),
    .A_N(\u_toplayer.reg_layer1[42] ));
 sg13g2_o21ai_1 _11097_ (.B1(_04692_),
    .Y(_04693_),
    .A1(net3259),
    .A2(\u_toplayer.reg_layer1[34] ));
 sg13g2_a22oi_1 _11098_ (.Y(_04694_),
    .B1(net2954),
    .B2(\u_toplayer.reg_layer1[50] ),
    .A2(net2985),
    .A1(\u_toplayer.reg_layer1[58] ));
 sg13g2_o21ai_1 _11099_ (.B1(_04694_),
    .Y(_04695_),
    .A1(net3244),
    .A2(_04693_));
 sg13g2_a221oi_1 _11100_ (.B2(net2915),
    .C1(net3233),
    .B1(_04695_),
    .A1(net2997),
    .Y(_04696_),
    .A2(_04691_));
 sg13g2_a21oi_1 _11101_ (.A1(net3275),
    .A2(_01127_),
    .Y(_04697_),
    .B1(net3254));
 sg13g2_o21ai_1 _11102_ (.B1(_04697_),
    .Y(_04698_),
    .A1(net3275),
    .A2(\u_toplayer.reg_layer1[194] ));
 sg13g2_a22oi_1 _11103_ (.Y(_04699_),
    .B1(net2963),
    .B2(\u_toplayer.reg_layer1[210] ),
    .A2(net2992),
    .A1(\u_toplayer.reg_layer1[218] ));
 sg13g2_nand3_1 _11104_ (.B(_04698_),
    .C(_04699_),
    .A(net3020),
    .Y(_04700_));
 sg13g2_a21oi_1 _11105_ (.A1(net3266),
    .A2(_01128_),
    .Y(_04701_),
    .B1(net3249));
 sg13g2_o21ai_1 _11106_ (.B1(_04701_),
    .Y(_04702_),
    .A1(net3265),
    .A2(\u_toplayer.reg_layer1[226] ));
 sg13g2_a22oi_1 _11107_ (.Y(_04703_),
    .B1(net2959),
    .B2(\u_toplayer.reg_layer1[242] ),
    .A2(net2987),
    .A1(\u_toplayer.reg_layer1[250] ));
 sg13g2_nand3_1 _11108_ (.B(_04702_),
    .C(_04703_),
    .A(net3240),
    .Y(_04704_));
 sg13g2_nand3_1 _11109_ (.B(_04700_),
    .C(_04704_),
    .A(net3236),
    .Y(_04705_));
 sg13g2_nor2b_1 _11110_ (.A(net3259),
    .B_N(\u_toplayer.reg_layer1[162] ),
    .Y(_04706_));
 sg13g2_a21oi_1 _11111_ (.A1(net3259),
    .A2(\u_toplayer.reg_layer1[170] ),
    .Y(_04707_),
    .B1(_04706_));
 sg13g2_a22oi_1 _11112_ (.Y(_04708_),
    .B1(net2954),
    .B2(\u_toplayer.reg_layer1[178] ),
    .A2(net2985),
    .A1(\u_toplayer.reg_layer1[186] ));
 sg13g2_o21ai_1 _11113_ (.B1(_04708_),
    .Y(_04709_),
    .A1(net3244),
    .A2(_04707_));
 sg13g2_nand2b_1 _11114_ (.Y(_04710_),
    .B(net3262),
    .A_N(\u_toplayer.reg_layer1[138] ));
 sg13g2_o21ai_1 _11115_ (.B1(_04710_),
    .Y(_04711_),
    .A1(net3262),
    .A2(\u_toplayer.reg_layer1[130] ));
 sg13g2_a22oi_1 _11116_ (.Y(_04712_),
    .B1(net2954),
    .B2(\u_toplayer.reg_layer1[146] ),
    .A2(net2985),
    .A1(\u_toplayer.reg_layer1[154] ));
 sg13g2_o21ai_1 _11117_ (.B1(_04712_),
    .Y(_04713_),
    .A1(net3246),
    .A2(_04711_));
 sg13g2_a22oi_1 _11118_ (.Y(_04714_),
    .B1(_04713_),
    .B2(net2996),
    .A2(_04709_),
    .A1(net2914));
 sg13g2_and2_1 _11119_ (.A(net3233),
    .B(_04714_),
    .X(_04715_));
 sg13g2_a221oi_1 _11120_ (.B2(_04715_),
    .C1(_04601_),
    .B1(_04705_),
    .A1(_04687_),
    .Y(_04716_),
    .A2(_04696_));
 sg13g2_a21o_1 _11121_ (.A2(_02647_),
    .A1(net3090),
    .B1(_04716_),
    .X(_00654_));
 sg13g2_a21oi_1 _11122_ (.A1(net3266),
    .A2(_01130_),
    .Y(_04717_),
    .B1(net3249));
 sg13g2_o21ai_1 _11123_ (.B1(_04717_),
    .Y(_04718_),
    .A1(net3265),
    .A2(\u_toplayer.reg_layer1[99] ));
 sg13g2_a22oi_1 _11124_ (.Y(_04719_),
    .B1(net2960),
    .B2(\u_toplayer.reg_layer1[115] ),
    .A2(net2990),
    .A1(\u_toplayer.reg_layer1[123] ));
 sg13g2_nand3_1 _11125_ (.B(_04718_),
    .C(_04719_),
    .A(net3240),
    .Y(_04720_));
 sg13g2_a21oi_1 _11126_ (.A1(net3276),
    .A2(_01129_),
    .Y(_04721_),
    .B1(net3254));
 sg13g2_o21ai_1 _11127_ (.B1(_04721_),
    .Y(_04722_),
    .A1(net3276),
    .A2(\u_toplayer.reg_layer1[67] ));
 sg13g2_a22oi_1 _11128_ (.Y(_04723_),
    .B1(net2963),
    .B2(\u_toplayer.reg_layer1[83] ),
    .A2(net2992),
    .A1(\u_toplayer.reg_layer1[91] ));
 sg13g2_nand3_1 _11129_ (.B(_04722_),
    .C(_04723_),
    .A(net3019),
    .Y(_04724_));
 sg13g2_nand3_1 _11130_ (.B(_04720_),
    .C(_04724_),
    .A(net3235),
    .Y(_04725_));
 sg13g2_nand2b_1 _11131_ (.Y(_04726_),
    .B(net3271),
    .A_N(\u_toplayer.reg_layer1[11] ));
 sg13g2_o21ai_1 _11132_ (.B1(_04726_),
    .Y(_04727_),
    .A1(net3271),
    .A2(\u_toplayer.reg_layer1[3] ));
 sg13g2_a22oi_1 _11133_ (.Y(_04728_),
    .B1(net2958),
    .B2(\u_toplayer.reg_layer1[19] ),
    .A2(net2988),
    .A1(\u_toplayer.reg_layer1[27] ));
 sg13g2_o21ai_1 _11134_ (.B1(_04728_),
    .Y(_04729_),
    .A1(net3252),
    .A2(_04727_));
 sg13g2_nand2b_1 _11135_ (.Y(_04730_),
    .B(net3264),
    .A_N(\u_toplayer.reg_layer1[43] ));
 sg13g2_o21ai_1 _11136_ (.B1(_04730_),
    .Y(_04731_),
    .A1(net3259),
    .A2(\u_toplayer.reg_layer1[35] ));
 sg13g2_a22oi_1 _11137_ (.Y(_04732_),
    .B1(net2954),
    .B2(\u_toplayer.reg_layer1[51] ),
    .A2(net2985),
    .A1(\u_toplayer.reg_layer1[59] ));
 sg13g2_o21ai_1 _11138_ (.B1(_04732_),
    .Y(_04733_),
    .A1(net3244),
    .A2(_04731_));
 sg13g2_a221oi_1 _11139_ (.B2(net2915),
    .C1(net3232),
    .B1(_04733_),
    .A1(net2997),
    .Y(_04734_),
    .A2(_04729_));
 sg13g2_a21oi_1 _11140_ (.A1(net3274),
    .A2(_01132_),
    .Y(_04735_),
    .B1(net3250));
 sg13g2_o21ai_1 _11141_ (.B1(_04735_),
    .Y(_04736_),
    .A1(net3266),
    .A2(\u_toplayer.reg_layer1[227] ));
 sg13g2_a22oi_1 _11142_ (.Y(_04737_),
    .B1(net2960),
    .B2(\u_toplayer.reg_layer1[243] ),
    .A2(net2990),
    .A1(\u_toplayer.reg_layer1[251] ));
 sg13g2_nand3_1 _11143_ (.B(_04736_),
    .C(_04737_),
    .A(net3240),
    .Y(_04738_));
 sg13g2_a21oi_1 _11144_ (.A1(net3276),
    .A2(_01131_),
    .Y(_04739_),
    .B1(net3254));
 sg13g2_o21ai_1 _11145_ (.B1(_04739_),
    .Y(_04740_),
    .A1(net3276),
    .A2(\u_toplayer.reg_layer1[195] ));
 sg13g2_a22oi_1 _11146_ (.Y(_04741_),
    .B1(net2963),
    .B2(\u_toplayer.reg_layer1[211] ),
    .A2(net2992),
    .A1(\u_toplayer.reg_layer1[219] ));
 sg13g2_nand3_1 _11147_ (.B(_04740_),
    .C(_04741_),
    .A(net3019),
    .Y(_04742_));
 sg13g2_nand3_1 _11148_ (.B(_04738_),
    .C(_04742_),
    .A(net3235),
    .Y(_04743_));
 sg13g2_nor2b_1 _11149_ (.A(net3261),
    .B_N(\u_toplayer.reg_layer1[131] ),
    .Y(_04744_));
 sg13g2_a21oi_1 _11150_ (.A1(net3261),
    .A2(\u_toplayer.reg_layer1[139] ),
    .Y(_04745_),
    .B1(_04744_));
 sg13g2_a22oi_1 _11151_ (.Y(_04746_),
    .B1(net2957),
    .B2(\u_toplayer.reg_layer1[147] ),
    .A2(net2989),
    .A1(\u_toplayer.reg_layer1[155] ));
 sg13g2_o21ai_1 _11152_ (.B1(_04746_),
    .Y(_04747_),
    .A1(net3246),
    .A2(_04745_));
 sg13g2_nand2b_1 _11153_ (.Y(_04748_),
    .B(net3259),
    .A_N(\u_toplayer.reg_layer1[171] ));
 sg13g2_o21ai_1 _11154_ (.B1(_04748_),
    .Y(_04749_),
    .A1(net3259),
    .A2(\u_toplayer.reg_layer1[163] ));
 sg13g2_a22oi_1 _11155_ (.Y(_04750_),
    .B1(net2954),
    .B2(\u_toplayer.reg_layer1[179] ),
    .A2(net2985),
    .A1(\u_toplayer.reg_layer1[187] ));
 sg13g2_o21ai_1 _11156_ (.B1(_04750_),
    .Y(_04751_),
    .A1(net3244),
    .A2(_04749_));
 sg13g2_a22oi_1 _11157_ (.Y(_04752_),
    .B1(_04751_),
    .B2(net2915),
    .A2(_04747_),
    .A1(net2996));
 sg13g2_and2_1 _11158_ (.A(net3232),
    .B(_04752_),
    .X(_04753_));
 sg13g2_a221oi_1 _11159_ (.B2(_04753_),
    .C1(_04601_),
    .B1(_04743_),
    .A1(_04725_),
    .Y(_04754_),
    .A2(_04734_));
 sg13g2_a21o_1 _11160_ (.A2(_02647_),
    .A1(net3088),
    .B1(_04754_),
    .X(_00655_));
 sg13g2_a21oi_1 _11161_ (.A1(net3274),
    .A2(_01133_),
    .Y(_04755_),
    .B1(net3253));
 sg13g2_o21ai_1 _11162_ (.B1(_04755_),
    .Y(_04756_),
    .A1(net3273),
    .A2(\u_toplayer.reg_layer1[68] ));
 sg13g2_a221oi_1 _11163_ (.B2(\u_toplayer.reg_layer1[84] ),
    .C1(net3239),
    .B1(net2962),
    .A1(\u_toplayer.reg_layer1[92] ),
    .Y(_04757_),
    .A2(net2991));
 sg13g2_nor2b_1 _11164_ (.A(\u_toplayer.reg_layer1[108] ),
    .B_N(net3265),
    .Y(_04758_));
 sg13g2_nor2_1 _11165_ (.A(net3269),
    .B(\u_toplayer.reg_layer1[100] ),
    .Y(_04759_));
 sg13g2_nor3_1 _11166_ (.A(net3251),
    .B(_04758_),
    .C(_04759_),
    .Y(_04760_));
 sg13g2_a221oi_1 _11167_ (.B2(\u_toplayer.reg_layer1[116] ),
    .C1(_04760_),
    .B1(net2961),
    .A1(\u_toplayer.reg_layer1[124] ),
    .Y(_04761_),
    .A2(net2990));
 sg13g2_a22oi_1 _11168_ (.Y(_04762_),
    .B1(_04761_),
    .B2(net3239),
    .A2(_04757_),
    .A1(_04756_));
 sg13g2_nor2b_1 _11169_ (.A(net3270),
    .B_N(\u_toplayer.reg_layer1[4] ),
    .Y(_04763_));
 sg13g2_a21oi_1 _11170_ (.A1(net3270),
    .A2(\u_toplayer.reg_layer1[12] ),
    .Y(_04764_),
    .B1(_04763_));
 sg13g2_a22oi_1 _11171_ (.Y(_04765_),
    .B1(net2957),
    .B2(\u_toplayer.reg_layer1[20] ),
    .A2(net2985),
    .A1(\u_toplayer.reg_layer1[28] ));
 sg13g2_o21ai_1 _11172_ (.B1(_04765_),
    .Y(_04766_),
    .A1(net3252),
    .A2(_04764_));
 sg13g2_nand2b_1 _11173_ (.Y(_04767_),
    .B(net3263),
    .A_N(\u_toplayer.reg_layer1[44] ));
 sg13g2_o21ai_1 _11174_ (.B1(_04767_),
    .Y(_04768_),
    .A1(net3263),
    .A2(\u_toplayer.reg_layer1[36] ));
 sg13g2_a22oi_1 _11175_ (.Y(_04769_),
    .B1(net2959),
    .B2(\u_toplayer.reg_layer1[52] ),
    .A2(net2987),
    .A1(\u_toplayer.reg_layer1[60] ));
 sg13g2_o21ai_1 _11176_ (.B1(_04769_),
    .Y(_04770_),
    .A1(net3248),
    .A2(_04768_));
 sg13g2_a21o_1 _11177_ (.A2(_04766_),
    .A1(net2997),
    .B1(net3233),
    .X(_04771_));
 sg13g2_a221oi_1 _11178_ (.B2(net2915),
    .C1(_04771_),
    .B1(_04770_),
    .A1(net3235),
    .Y(_04772_),
    .A2(_04762_));
 sg13g2_nor2b_1 _11179_ (.A(\u_toplayer.reg_layer1[236] ),
    .B_N(net3265),
    .Y(_04773_));
 sg13g2_nor2_1 _11180_ (.A(net3269),
    .B(\u_toplayer.reg_layer1[228] ),
    .Y(_04774_));
 sg13g2_nor3_1 _11181_ (.A(net3251),
    .B(_04773_),
    .C(_04774_),
    .Y(_04775_));
 sg13g2_a221oi_1 _11182_ (.B2(\u_toplayer.reg_layer1[244] ),
    .C1(_04775_),
    .B1(net2961),
    .A1(\u_toplayer.reg_layer1[252] ),
    .Y(_04776_),
    .A2(net2990));
 sg13g2_a21oi_1 _11183_ (.A1(net3274),
    .A2(_01134_),
    .Y(_04777_),
    .B1(net3253));
 sg13g2_o21ai_1 _11184_ (.B1(_04777_),
    .Y(_04778_),
    .A1(net3274),
    .A2(\u_toplayer.reg_layer1[196] ));
 sg13g2_a221oi_1 _11185_ (.B2(\u_toplayer.reg_layer1[212] ),
    .C1(net3241),
    .B1(net2962),
    .A1(\u_toplayer.reg_layer1[220] ),
    .Y(_04779_),
    .A2(net2991));
 sg13g2_a22oi_1 _11186_ (.Y(_04780_),
    .B1(_04778_),
    .B2(_04779_),
    .A2(_04776_),
    .A1(net3239));
 sg13g2_nor2b_1 _11187_ (.A(net3262),
    .B_N(\u_toplayer.reg_layer1[132] ),
    .Y(_04781_));
 sg13g2_a21oi_1 _11188_ (.A1(net3262),
    .A2(\u_toplayer.reg_layer1[140] ),
    .Y(_04782_),
    .B1(_04781_));
 sg13g2_a22oi_1 _11189_ (.Y(_04783_),
    .B1(net2957),
    .B2(\u_toplayer.reg_layer1[148] ),
    .A2(net2988),
    .A1(\u_toplayer.reg_layer1[156] ));
 sg13g2_o21ai_1 _11190_ (.B1(_04783_),
    .Y(_04784_),
    .A1(net3246),
    .A2(_04782_));
 sg13g2_nand2b_1 _11191_ (.Y(_04785_),
    .B(net3263),
    .A_N(\u_toplayer.reg_layer1[172] ));
 sg13g2_o21ai_1 _11192_ (.B1(_04785_),
    .Y(_04786_),
    .A1(net3263),
    .A2(\u_toplayer.reg_layer1[164] ));
 sg13g2_a22oi_1 _11193_ (.Y(_04787_),
    .B1(net2957),
    .B2(\u_toplayer.reg_layer1[180] ),
    .A2(net2988),
    .A1(\u_toplayer.reg_layer1[188] ));
 sg13g2_o21ai_1 _11194_ (.B1(_04787_),
    .Y(_04788_),
    .A1(net3247),
    .A2(_04786_));
 sg13g2_a22oi_1 _11195_ (.Y(_04789_),
    .B1(_04788_),
    .B2(net2914),
    .A2(_04784_),
    .A1(net2996));
 sg13g2_nand2_1 _11196_ (.Y(_04790_),
    .A(net3231),
    .B(_04789_));
 sg13g2_a21oi_1 _11197_ (.A1(net3235),
    .A2(_04780_),
    .Y(_04791_),
    .B1(_04790_));
 sg13g2_nor3_2 _11198_ (.A(_04601_),
    .B(_04772_),
    .C(_04791_),
    .Y(_04792_));
 sg13g2_a21o_1 _11199_ (.A2(_02647_),
    .A1(net3086),
    .B1(_04792_),
    .X(_00656_));
 sg13g2_a21oi_1 _11200_ (.A1(net3266),
    .A2(_01138_),
    .Y(_04793_),
    .B1(net3249));
 sg13g2_o21ai_1 _11201_ (.B1(_04793_),
    .Y(_04794_),
    .A1(net3265),
    .A2(\u_toplayer.reg_layer1[229] ));
 sg13g2_a22oi_1 _11202_ (.Y(_04795_),
    .B1(net2959),
    .B2(\u_toplayer.reg_layer1[245] ),
    .A2(net2987),
    .A1(\u_toplayer.reg_layer1[253] ));
 sg13g2_nand3_1 _11203_ (.B(_04794_),
    .C(_04795_),
    .A(net3241),
    .Y(_04796_));
 sg13g2_a21oi_1 _11204_ (.A1(net3273),
    .A2(_01137_),
    .Y(_04797_),
    .B1(net3250));
 sg13g2_o21ai_1 _11205_ (.B1(_04797_),
    .Y(_04798_),
    .A1(net3268),
    .A2(\u_toplayer.reg_layer1[197] ));
 sg13g2_a221oi_1 _11206_ (.B2(\u_toplayer.reg_layer1[213] ),
    .C1(net3241),
    .B1(net2963),
    .A1(\u_toplayer.reg_layer1[221] ),
    .Y(_04799_),
    .A2(net2992));
 sg13g2_nand2_1 _11207_ (.Y(_04800_),
    .A(net3237),
    .B(_04796_));
 sg13g2_a21oi_2 _11208_ (.B1(_04800_),
    .Y(_04801_),
    .A2(_04799_),
    .A1(_04798_));
 sg13g2_nor2b_1 _11209_ (.A(net3262),
    .B_N(\u_toplayer.reg_layer1[133] ),
    .Y(_04802_));
 sg13g2_a21oi_1 _11210_ (.A1(net3262),
    .A2(\u_toplayer.reg_layer1[141] ),
    .Y(_04803_),
    .B1(_04802_));
 sg13g2_a22oi_1 _11211_ (.Y(_04804_),
    .B1(net2957),
    .B2(\u_toplayer.reg_layer1[149] ),
    .A2(net2989),
    .A1(\u_toplayer.reg_layer1[157] ));
 sg13g2_o21ai_1 _11212_ (.B1(_04804_),
    .Y(_04805_),
    .A1(net3246),
    .A2(_04803_));
 sg13g2_nand2b_1 _11213_ (.Y(_04806_),
    .B(net3263),
    .A_N(\u_toplayer.reg_layer1[173] ));
 sg13g2_o21ai_1 _11214_ (.B1(_04806_),
    .Y(_04807_),
    .A1(net3263),
    .A2(\u_toplayer.reg_layer1[165] ));
 sg13g2_a22oi_1 _11215_ (.Y(_04808_),
    .B1(net2957),
    .B2(\u_toplayer.reg_layer1[181] ),
    .A2(net2988),
    .A1(\u_toplayer.reg_layer1[189] ));
 sg13g2_o21ai_1 _11216_ (.B1(_04808_),
    .Y(_04809_),
    .A1(net3247),
    .A2(_04807_));
 sg13g2_a221oi_1 _11217_ (.B2(net2915),
    .C1(_04801_),
    .B1(_04809_),
    .A1(net2997),
    .Y(_04810_),
    .A2(_04805_));
 sg13g2_a21oi_1 _11218_ (.A1(net3273),
    .A2(_01135_),
    .Y(_04811_),
    .B1(net3253));
 sg13g2_o21ai_1 _11219_ (.B1(_04811_),
    .Y(_04812_),
    .A1(net3273),
    .A2(\u_toplayer.reg_layer1[69] ));
 sg13g2_a22oi_1 _11220_ (.Y(_04813_),
    .B1(net2963),
    .B2(\u_toplayer.reg_layer1[85] ),
    .A2(net2992),
    .A1(\u_toplayer.reg_layer1[93] ));
 sg13g2_nand3_1 _11221_ (.B(_04812_),
    .C(_04813_),
    .A(net3019),
    .Y(_04814_));
 sg13g2_a21oi_1 _11222_ (.A1(net3266),
    .A2(_01136_),
    .Y(_04815_),
    .B1(net3249));
 sg13g2_o21ai_1 _11223_ (.B1(_04815_),
    .Y(_04816_),
    .A1(net3269),
    .A2(\u_toplayer.reg_layer1[101] ));
 sg13g2_a22oi_1 _11224_ (.Y(_04817_),
    .B1(net2960),
    .B2(\u_toplayer.reg_layer1[117] ),
    .A2(net2987),
    .A1(\u_toplayer.reg_layer1[125] ));
 sg13g2_nand3_1 _11225_ (.B(_04816_),
    .C(_04817_),
    .A(net3240),
    .Y(_04818_));
 sg13g2_nand3_1 _11226_ (.B(_04814_),
    .C(_04818_),
    .A(net3236),
    .Y(_04819_));
 sg13g2_nor2b_1 _11227_ (.A(net3263),
    .B_N(\u_toplayer.reg_layer1[37] ),
    .Y(_04820_));
 sg13g2_a21oi_1 _11228_ (.A1(net3263),
    .A2(\u_toplayer.reg_layer1[45] ),
    .Y(_04821_),
    .B1(_04820_));
 sg13g2_a22oi_1 _11229_ (.Y(_04822_),
    .B1(net2957),
    .B2(\u_toplayer.reg_layer1[53] ),
    .A2(net2988),
    .A1(\u_toplayer.reg_layer1[61] ));
 sg13g2_o21ai_1 _11230_ (.B1(_04822_),
    .Y(_04823_),
    .A1(net3247),
    .A2(_04821_));
 sg13g2_nand2b_1 _11231_ (.Y(_04824_),
    .B(net3270),
    .A_N(\u_toplayer.reg_layer1[13] ));
 sg13g2_o21ai_1 _11232_ (.B1(_04824_),
    .Y(_04825_),
    .A1(net3270),
    .A2(\u_toplayer.reg_layer1[5] ));
 sg13g2_a22oi_1 _11233_ (.Y(_04826_),
    .B1(net2957),
    .B2(\u_toplayer.reg_layer1[21] ),
    .A2(net2988),
    .A1(\u_toplayer.reg_layer1[29] ));
 sg13g2_o21ai_1 _11234_ (.B1(_04826_),
    .Y(_04827_),
    .A1(net3246),
    .A2(_04825_));
 sg13g2_a221oi_1 _11235_ (.B2(_01349_),
    .C1(net3231),
    .B1(_04827_),
    .A1(net2915),
    .Y(_04828_),
    .A2(_04823_));
 sg13g2_a221oi_1 _11236_ (.B2(_04828_),
    .C1(_04601_),
    .B1(_04819_),
    .A1(net3231),
    .Y(_04829_),
    .A2(_04810_));
 sg13g2_a21oi_1 _11237_ (.A1(net3085),
    .A2(_02647_),
    .Y(_04830_),
    .B1(_04829_));
 sg13g2_inv_1 _11238_ (.Y(_00657_),
    .A(_04830_));
 sg13g2_a21oi_1 _11239_ (.A1(net3273),
    .A2(_01139_),
    .Y(_04831_),
    .B1(net3253));
 sg13g2_o21ai_1 _11240_ (.B1(_04831_),
    .Y(_04832_),
    .A1(net3273),
    .A2(\u_toplayer.reg_layer1[70] ));
 sg13g2_a22oi_1 _11241_ (.Y(_04833_),
    .B1(net2962),
    .B2(\u_toplayer.reg_layer1[86] ),
    .A2(net2991),
    .A1(\u_toplayer.reg_layer1[94] ));
 sg13g2_nand3_1 _11242_ (.B(_04832_),
    .C(_04833_),
    .A(net3019),
    .Y(_04834_));
 sg13g2_a21oi_1 _11243_ (.A1(net3267),
    .A2(_01140_),
    .Y(_04835_),
    .B1(net3251));
 sg13g2_o21ai_1 _11244_ (.B1(_04835_),
    .Y(_04836_),
    .A1(net3269),
    .A2(\u_toplayer.reg_layer1[102] ));
 sg13g2_a22oi_1 _11245_ (.Y(_04837_),
    .B1(net2960),
    .B2(\u_toplayer.reg_layer1[118] ),
    .A2(net2987),
    .A1(\u_toplayer.reg_layer1[126] ));
 sg13g2_nand3_1 _11246_ (.B(_04836_),
    .C(_04837_),
    .A(net3239),
    .Y(_04838_));
 sg13g2_nand3_1 _11247_ (.B(_04834_),
    .C(_04838_),
    .A(net3236),
    .Y(_04839_));
 sg13g2_nand2b_1 _11248_ (.Y(_04840_),
    .B(net3261),
    .A_N(\u_toplayer.reg_layer1[14] ));
 sg13g2_o21ai_1 _11249_ (.B1(_04840_),
    .Y(_04841_),
    .A1(net3261),
    .A2(\u_toplayer.reg_layer1[6] ));
 sg13g2_a22oi_1 _11250_ (.Y(_04842_),
    .B1(net2958),
    .B2(\u_toplayer.reg_layer1[22] ),
    .A2(net2986),
    .A1(\u_toplayer.reg_layer1[30] ));
 sg13g2_o21ai_1 _11251_ (.B1(_04842_),
    .Y(_04843_),
    .A1(net3246),
    .A2(_04841_));
 sg13g2_nor2b_1 _11252_ (.A(net3256),
    .B_N(\u_toplayer.reg_layer1[38] ),
    .Y(_04844_));
 sg13g2_a21oi_1 _11253_ (.A1(net3256),
    .A2(\u_toplayer.reg_layer1[46] ),
    .Y(_04845_),
    .B1(_04844_));
 sg13g2_a22oi_1 _11254_ (.Y(_04846_),
    .B1(net2955),
    .B2(\u_toplayer.reg_layer1[54] ),
    .A2(net2984),
    .A1(\u_toplayer.reg_layer1[62] ));
 sg13g2_o21ai_1 _11255_ (.B1(_04846_),
    .Y(_04847_),
    .A1(net3243),
    .A2(_04845_));
 sg13g2_a221oi_1 _11256_ (.B2(net2914),
    .C1(net3231),
    .B1(_04847_),
    .A1(net2996),
    .Y(_04848_),
    .A2(_04843_));
 sg13g2_a21oi_1 _11257_ (.A1(net3267),
    .A2(_01142_),
    .Y(_04849_),
    .B1(net3250));
 sg13g2_o21ai_1 _11258_ (.B1(_04849_),
    .Y(_04850_),
    .A1(net3269),
    .A2(\u_toplayer.reg_layer1[230] ));
 sg13g2_a22oi_1 _11259_ (.Y(_04851_),
    .B1(net2959),
    .B2(\u_toplayer.reg_layer1[246] ),
    .A2(net2987),
    .A1(\u_toplayer.reg_layer1[254] ));
 sg13g2_nand3_1 _11260_ (.B(_04850_),
    .C(_04851_),
    .A(net3239),
    .Y(_04852_));
 sg13g2_a21oi_1 _11261_ (.A1(net3273),
    .A2(_01141_),
    .Y(_04853_),
    .B1(net3253));
 sg13g2_o21ai_1 _11262_ (.B1(_04853_),
    .Y(_04854_),
    .A1(net3273),
    .A2(\u_toplayer.reg_layer1[198] ));
 sg13g2_a22oi_1 _11263_ (.Y(_04855_),
    .B1(net2962),
    .B2(\u_toplayer.reg_layer1[214] ),
    .A2(net2991),
    .A1(\u_toplayer.reg_layer1[222] ));
 sg13g2_nand3_1 _11264_ (.B(_04854_),
    .C(_04855_),
    .A(net3019),
    .Y(_04856_));
 sg13g2_nand3_1 _11265_ (.B(_04852_),
    .C(_04856_),
    .A(net3236),
    .Y(_04857_));
 sg13g2_nand2b_1 _11266_ (.Y(_04858_),
    .B(net3260),
    .A_N(\u_toplayer.reg_layer1[142] ));
 sg13g2_o21ai_1 _11267_ (.B1(_04858_),
    .Y(_04859_),
    .A1(net3260),
    .A2(\u_toplayer.reg_layer1[134] ));
 sg13g2_a22oi_1 _11268_ (.Y(_04860_),
    .B1(net2958),
    .B2(\u_toplayer.reg_layer1[150] ),
    .A2(net2986),
    .A1(\u_toplayer.reg_layer1[158] ));
 sg13g2_o21ai_1 _11269_ (.B1(_04860_),
    .Y(_04861_),
    .A1(net3247),
    .A2(_04859_));
 sg13g2_nor2b_1 _11270_ (.A(net3257),
    .B_N(\u_toplayer.reg_layer1[166] ),
    .Y(_04862_));
 sg13g2_a21oi_1 _11271_ (.A1(net3256),
    .A2(\u_toplayer.reg_layer1[174] ),
    .Y(_04863_),
    .B1(_04862_));
 sg13g2_a22oi_1 _11272_ (.Y(_04864_),
    .B1(net2955),
    .B2(\u_toplayer.reg_layer1[182] ),
    .A2(net2984),
    .A1(\u_toplayer.reg_layer1[190] ));
 sg13g2_o21ai_1 _11273_ (.B1(_04864_),
    .Y(_04865_),
    .A1(net3243),
    .A2(_04863_));
 sg13g2_a22oi_1 _11274_ (.Y(_04866_),
    .B1(_04865_),
    .B2(net2914),
    .A2(_04861_),
    .A1(net2996));
 sg13g2_and2_1 _11275_ (.A(net3231),
    .B(_04866_),
    .X(_04867_));
 sg13g2_a221oi_1 _11276_ (.B2(_04867_),
    .C1(_04601_),
    .B1(_04857_),
    .A1(_04839_),
    .Y(_04868_),
    .A2(_04848_));
 sg13g2_a21o_1 _11277_ (.A2(_02647_),
    .A1(net3084),
    .B1(_04868_),
    .X(_00658_));
 sg13g2_a21oi_1 _11278_ (.A1(net3265),
    .A2(_01144_),
    .Y(_04869_),
    .B1(net3249));
 sg13g2_o21ai_1 _11279_ (.B1(_04869_),
    .Y(_04870_),
    .A1(net3269),
    .A2(\u_toplayer.reg_layer1[103] ));
 sg13g2_a22oi_1 _11280_ (.Y(_04871_),
    .B1(net2960),
    .B2(\u_toplayer.reg_layer1[119] ),
    .A2(net2989),
    .A1(\u_toplayer.reg_layer1[127] ));
 sg13g2_nand3_1 _11281_ (.B(_04870_),
    .C(_04871_),
    .A(net3240),
    .Y(_04872_));
 sg13g2_a21oi_1 _11282_ (.A1(net3276),
    .A2(_01143_),
    .Y(_04873_),
    .B1(net3253));
 sg13g2_o21ai_1 _11283_ (.B1(_04873_),
    .Y(_04874_),
    .A1(net3276),
    .A2(\u_toplayer.reg_layer1[71] ));
 sg13g2_a22oi_1 _11284_ (.Y(_04875_),
    .B1(net2963),
    .B2(\u_toplayer.reg_layer1[87] ),
    .A2(net2993),
    .A1(\u_toplayer.reg_layer1[95] ));
 sg13g2_nand3_1 _11285_ (.B(_04874_),
    .C(_04875_),
    .A(net3020),
    .Y(_04876_));
 sg13g2_nand3_1 _11286_ (.B(_04872_),
    .C(_04876_),
    .A(net3235),
    .Y(_04877_));
 sg13g2_nand2b_1 _11287_ (.Y(_04878_),
    .B(net3257),
    .A_N(\u_toplayer.reg_layer1[47] ));
 sg13g2_o21ai_1 _11288_ (.B1(_04878_),
    .Y(_04879_),
    .A1(net3256),
    .A2(\u_toplayer.reg_layer1[39] ));
 sg13g2_a22oi_1 _11289_ (.Y(_04880_),
    .B1(net2955),
    .B2(\u_toplayer.reg_layer1[55] ),
    .A2(net2984),
    .A1(\u_toplayer.reg_layer1[63] ));
 sg13g2_o21ai_1 _11290_ (.B1(_04880_),
    .Y(_04881_),
    .A1(net3243),
    .A2(_04879_));
 sg13g2_nand2b_1 _11291_ (.Y(_04882_),
    .B(net3260),
    .A_N(\u_toplayer.reg_layer1[15] ));
 sg13g2_o21ai_1 _11292_ (.B1(_04882_),
    .Y(_04883_),
    .A1(net3261),
    .A2(\u_toplayer.reg_layer1[7] ));
 sg13g2_a22oi_1 _11293_ (.Y(_04884_),
    .B1(net2956),
    .B2(\u_toplayer.reg_layer1[23] ),
    .A2(net2986),
    .A1(\u_toplayer.reg_layer1[31] ));
 sg13g2_o21ai_1 _11294_ (.B1(_04884_),
    .Y(_04885_),
    .A1(net3247),
    .A2(_04883_));
 sg13g2_a221oi_1 _11295_ (.B2(net2997),
    .C1(net3231),
    .B1(_04885_),
    .A1(net2914),
    .Y(_04886_),
    .A2(_04881_));
 sg13g2_a21oi_1 _11296_ (.A1(net3265),
    .A2(_01146_),
    .Y(_04887_),
    .B1(net3249));
 sg13g2_o21ai_1 _11297_ (.B1(_04887_),
    .Y(_04888_),
    .A1(net3269),
    .A2(\u_toplayer.reg_layer1[231] ));
 sg13g2_a22oi_1 _11298_ (.Y(_04889_),
    .B1(net2959),
    .B2(\u_toplayer.reg_layer1[247] ),
    .A2(net2987),
    .A1(\u_toplayer.reg_layer1[255] ));
 sg13g2_nand3_1 _11299_ (.B(_04888_),
    .C(_04889_),
    .A(net3240),
    .Y(_04890_));
 sg13g2_a21oi_1 _11300_ (.A1(net3276),
    .A2(_01145_),
    .Y(_04891_),
    .B1(net3253));
 sg13g2_o21ai_1 _11301_ (.B1(_04891_),
    .Y(_04892_),
    .A1(net3276),
    .A2(\u_toplayer.reg_layer1[199] ));
 sg13g2_a22oi_1 _11302_ (.Y(_04893_),
    .B1(net2963),
    .B2(\u_toplayer.reg_layer1[215] ),
    .A2(net2993),
    .A1(\u_toplayer.reg_layer1[223] ));
 sg13g2_nand3_1 _11303_ (.B(_04892_),
    .C(_04893_),
    .A(net3020),
    .Y(_04894_));
 sg13g2_nand3_1 _11304_ (.B(_04890_),
    .C(_04894_),
    .A(net3235),
    .Y(_04895_));
 sg13g2_nand2b_1 _11305_ (.Y(_04896_),
    .B(net3257),
    .A_N(\u_toplayer.reg_layer1[175] ));
 sg13g2_o21ai_1 _11306_ (.B1(_04896_),
    .Y(_04897_),
    .A1(net3256),
    .A2(\u_toplayer.reg_layer1[167] ));
 sg13g2_a22oi_1 _11307_ (.Y(_04898_),
    .B1(net2955),
    .B2(\u_toplayer.reg_layer1[183] ),
    .A2(net2984),
    .A1(\u_toplayer.reg_layer1[191] ));
 sg13g2_o21ai_1 _11308_ (.B1(_04898_),
    .Y(_04899_),
    .A1(net3243),
    .A2(_04897_));
 sg13g2_nor2b_1 _11309_ (.A(net3260),
    .B_N(\u_toplayer.reg_layer1[135] ),
    .Y(_04900_));
 sg13g2_a21oi_1 _11310_ (.A1(net3260),
    .A2(\u_toplayer.reg_layer1[143] ),
    .Y(_04901_),
    .B1(_04900_));
 sg13g2_a22oi_1 _11311_ (.Y(_04902_),
    .B1(net2954),
    .B2(\u_toplayer.reg_layer1[151] ),
    .A2(net2985),
    .A1(\u_toplayer.reg_layer1[159] ));
 sg13g2_o21ai_1 _11312_ (.B1(_04902_),
    .Y(_04903_),
    .A1(net3247),
    .A2(_04901_));
 sg13g2_a22oi_1 _11313_ (.Y(_04904_),
    .B1(_04903_),
    .B2(net2996),
    .A2(_04899_),
    .A1(net2914));
 sg13g2_and2_1 _11314_ (.A(net3231),
    .B(_04904_),
    .X(_04905_));
 sg13g2_a221oi_1 _11315_ (.B2(_04905_),
    .C1(_04601_),
    .B1(_04895_),
    .A1(_04877_),
    .Y(_04906_),
    .A2(_04886_));
 sg13g2_a21o_1 _11316_ (.A2(_02647_),
    .A1(net3082),
    .B1(_04906_),
    .X(_00659_));
 sg13g2_nand2_1 _11317_ (.Y(_04907_),
    .A(net2861),
    .B(_02648_));
 sg13g2_nand2_1 _11318_ (.Y(_04908_),
    .A(net3081),
    .B(net2819));
 sg13g2_nor4_1 _11319_ (.A(net3061),
    .B(\u_toplayer.u_layer2.u_neuron.acc[11] ),
    .C(\u_toplayer.u_layer2.u_neuron.acc[10] ),
    .D(\u_toplayer.u_layer2.u_neuron.acc[9] ),
    .Y(_04909_));
 sg13g2_nor4_1 _11320_ (.A(\u_toplayer.u_layer2.u_neuron.acc[7] ),
    .B(\u_toplayer.u_layer2.u_neuron.acc[15] ),
    .C(net3060),
    .D(\u_toplayer.u_layer2.u_neuron.acc[13] ),
    .Y(_04910_));
 sg13g2_nor4_1 _11321_ (.A(\u_toplayer.u_layer2.u_neuron.acc[8] ),
    .B(\u_toplayer.u_layer2.u_neuron.acc[22] ),
    .C(\u_toplayer.u_layer2.u_neuron.acc[21] ),
    .D(net3058),
    .Y(_04911_));
 sg13g2_nor4_1 _11322_ (.A(\u_toplayer.u_layer2.u_neuron.acc[19] ),
    .B(\u_toplayer.u_layer2.u_neuron.acc[18] ),
    .C(\u_toplayer.u_layer2.u_neuron.acc[17] ),
    .D(net3059),
    .Y(_04912_));
 sg13g2_and3_1 _11323_ (.X(_04913_),
    .A(_04909_),
    .B(_04910_),
    .C(_04912_));
 sg13g2_a21oi_2 _11324_ (.B1(net1164),
    .Y(_04914_),
    .A2(_04913_),
    .A1(_04911_));
 sg13g2_nor2_1 _11325_ (.A(net1037),
    .B(_04914_),
    .Y(_04915_));
 sg13g2_nand4_1 _11326_ (.B(\u_toplayer.u_layer2.u_neuron.acc[11] ),
    .C(net3062),
    .A(net3061),
    .Y(_04916_),
    .D(\u_toplayer.u_layer2.u_neuron.acc[9] ));
 sg13g2_nand4_1 _11327_ (.B(\u_toplayer.u_layer2.u_neuron.acc[15] ),
    .C(net3060),
    .A(\u_toplayer.u_layer2.u_neuron.acc[7] ),
    .Y(_04917_),
    .D(\u_toplayer.u_layer2.u_neuron.acc[13] ));
 sg13g2_nand4_1 _11328_ (.B(\u_toplayer.u_layer2.u_neuron.acc[22] ),
    .C(\u_toplayer.u_layer2.u_neuron.acc[21] ),
    .A(\u_toplayer.u_layer2.u_neuron.acc[8] ),
    .Y(_04918_),
    .D(net3058));
 sg13g2_nand4_1 _11329_ (.B(\u_toplayer.u_layer2.u_neuron.acc[18] ),
    .C(\u_toplayer.u_layer2.u_neuron.acc[17] ),
    .A(\u_toplayer.u_layer2.u_neuron.acc[19] ),
    .Y(_04919_),
    .D(net3059));
 sg13g2_nor3_1 _11330_ (.A(_01097_),
    .B(\u_toplayer.u_layer2.u_neuron.acc[6] ),
    .C(net3063),
    .Y(_04920_));
 sg13g2_nor4_1 _11331_ (.A(\u_toplayer.u_layer2.u_neuron.acc[3] ),
    .B(\u_toplayer.u_layer2.u_neuron.acc[2] ),
    .C(net3064),
    .D(\u_toplayer.u_layer2.u_neuron.acc[0] ),
    .Y(_04921_));
 sg13g2_nand3_1 _11332_ (.B(_04920_),
    .C(_04921_),
    .A(_01100_),
    .Y(_04922_));
 sg13g2_nor4_1 _11333_ (.A(_04916_),
    .B(_04917_),
    .C(_04918_),
    .D(_04919_),
    .Y(_04923_));
 sg13g2_a21oi_1 _11334_ (.A1(_04922_),
    .A2(_04923_),
    .Y(_04924_),
    .B1(_01110_));
 sg13g2_or2_2 _11335_ (.X(_04925_),
    .B(_04924_),
    .A(_04907_));
 sg13g2_o21ai_1 _11336_ (.B1(_04908_),
    .Y(_00660_),
    .A1(_04915_),
    .A2(_04925_));
 sg13g2_nand2_1 _11337_ (.Y(_04926_),
    .A(net3079),
    .B(net2819));
 sg13g2_nor2_1 _11338_ (.A(net3064),
    .B(_04914_),
    .Y(_04927_));
 sg13g2_o21ai_1 _11339_ (.B1(_04926_),
    .Y(_00661_),
    .A1(_04925_),
    .A2(_04927_));
 sg13g2_nand2_1 _11340_ (.Y(_04928_),
    .A(net3077),
    .B(net2819));
 sg13g2_nor2_1 _11341_ (.A(net1176),
    .B(_04914_),
    .Y(_04929_));
 sg13g2_o21ai_1 _11342_ (.B1(_04928_),
    .Y(_00662_),
    .A1(_04925_),
    .A2(_04929_));
 sg13g2_nand2_1 _11343_ (.Y(_04930_),
    .A(net3075),
    .B(net2819));
 sg13g2_nor2_1 _11344_ (.A(net1157),
    .B(_04914_),
    .Y(_04931_));
 sg13g2_o21ai_1 _11345_ (.B1(_04930_),
    .Y(_00663_),
    .A1(_04925_),
    .A2(_04931_));
 sg13g2_nand2_1 _11346_ (.Y(_04932_),
    .A(net3071),
    .B(net2819));
 sg13g2_nor2_1 _11347_ (.A(net1137),
    .B(_04914_),
    .Y(_04933_));
 sg13g2_o21ai_1 _11348_ (.B1(_04932_),
    .Y(_00664_),
    .A1(_04925_),
    .A2(_04933_));
 sg13g2_nand2_1 _11349_ (.Y(_04934_),
    .A(net3070),
    .B(net2819));
 sg13g2_nor2_1 _11350_ (.A(net3063),
    .B(_04914_),
    .Y(_04935_));
 sg13g2_o21ai_1 _11351_ (.B1(_04934_),
    .Y(_00665_),
    .A1(_04925_),
    .A2(_04935_));
 sg13g2_nand2_1 _11352_ (.Y(_04936_),
    .A(net3068),
    .B(net2819));
 sg13g2_nor2_1 _11353_ (.A(net1055),
    .B(_04914_),
    .Y(_04937_));
 sg13g2_o21ai_1 _11354_ (.B1(_04936_),
    .Y(_00666_),
    .A1(_04925_),
    .A2(_04937_));
 sg13g2_mux2_1 _11355_ (.A0(net1119),
    .A1(net3065),
    .S(net2819),
    .X(_00667_));
 sg13g2_xor2_1 _11356_ (.B(_03726_),
    .A(net860),
    .X(_00668_));
 sg13g2_nor2_1 _11357_ (.A(net954),
    .B(_03727_),
    .Y(_04938_));
 sg13g2_nor3_1 _11358_ (.A(_03717_),
    .B(_03728_),
    .C(_04938_),
    .Y(_00669_));
 sg13g2_xor2_1 _11359_ (.B(_03730_),
    .A(net979),
    .X(_00671_));
 sg13g2_nand3_1 _11360_ (.B(net979),
    .C(_03730_),
    .A(net1129),
    .Y(_04939_));
 sg13g2_a21o_1 _11361_ (.A2(_03730_),
    .A1(net979),
    .B1(net1129),
    .X(_04940_));
 sg13g2_and2_1 _11362_ (.A(_04939_),
    .B(_04940_),
    .X(_00672_));
 sg13g2_a21oi_1 _11363_ (.A1(_01034_),
    .A2(_04939_),
    .Y(_00673_),
    .B1(_03717_));
 sg13g2_nor2_1 _11364_ (.A(\u_toplayer.u_layer2.statel2[8] ),
    .B(_03726_),
    .Y(_04941_));
 sg13g2_a21oi_1 _11365_ (.A1(net122),
    .A2(_03726_),
    .Y(_00676_),
    .B1(_04941_));
 sg13g2_nand2_1 _11366_ (.Y(_04942_),
    .A(\u_toplayer.u_layer2.u_neuron.acc[0] ),
    .B(\u_toplayer.u_layer2.u_neuron.mult[0] ));
 sg13g2_xor2_1 _11367_ (.B(net929),
    .A(\u_toplayer.u_layer2.u_neuron.acc[0] ),
    .X(_04943_));
 sg13g2_nand2_1 _11368_ (.Y(_04944_),
    .A(net3403),
    .B(\u_toplayer.u_layer2.u_neuron.acc[0] ));
 sg13g2_xor2_1 _11369_ (.B(\u_toplayer.u_layer2.u_neuron.acc[0] ),
    .A(net3403),
    .X(_04945_));
 sg13g2_a221oi_1 _11370_ (.B2(net2887),
    .C1(net2755),
    .B1(_04945_),
    .A1(net2859),
    .Y(_04946_),
    .A2(_04943_));
 sg13g2_a21oi_1 _11371_ (.A1(_01103_),
    .A2(net2754),
    .Y(_00677_),
    .B1(_04946_));
 sg13g2_nand2_1 _11372_ (.Y(_04947_),
    .A(net3399),
    .B(net3064));
 sg13g2_nor2_1 _11373_ (.A(net3399),
    .B(net3064),
    .Y(_04948_));
 sg13g2_xor2_1 _11374_ (.B(net3064),
    .A(net3399),
    .X(_04949_));
 sg13g2_xnor2_1 _11375_ (.Y(_04950_),
    .A(_04944_),
    .B(_04949_));
 sg13g2_nand2_1 _11376_ (.Y(_04951_),
    .A(net3064),
    .B(\u_toplayer.u_layer2.u_neuron.mult[1] ));
 sg13g2_nor2_1 _11377_ (.A(net3064),
    .B(\u_toplayer.u_layer2.u_neuron.mult[1] ),
    .Y(_04952_));
 sg13g2_xor2_1 _11378_ (.B(\u_toplayer.u_layer2.u_neuron.mult[1] ),
    .A(net3064),
    .X(_04953_));
 sg13g2_xnor2_1 _11379_ (.Y(_04954_),
    .A(_04942_),
    .B(_04953_));
 sg13g2_a221oi_1 _11380_ (.B2(net2859),
    .C1(net2754),
    .B1(_04954_),
    .A1(net2887),
    .Y(_04955_),
    .A2(_04950_));
 sg13g2_a21oi_1 _11381_ (.A1(_01102_),
    .A2(net2754),
    .Y(_00678_),
    .B1(_04955_));
 sg13g2_o21ai_1 _11382_ (.B1(_04951_),
    .Y(_04956_),
    .A1(_04942_),
    .A2(_04952_));
 sg13g2_and2_1 _11383_ (.A(\u_toplayer.u_layer2.u_neuron.acc[2] ),
    .B(\u_toplayer.u_layer2.u_neuron.mult[2] ),
    .X(_04957_));
 sg13g2_xor2_1 _11384_ (.B(\u_toplayer.u_layer2.u_neuron.mult[2] ),
    .A(\u_toplayer.u_layer2.u_neuron.acc[2] ),
    .X(_04958_));
 sg13g2_xnor2_1 _11385_ (.Y(_04959_),
    .A(_04956_),
    .B(_04958_));
 sg13g2_and2_1 _11386_ (.A(net3396),
    .B(\u_toplayer.u_layer2.u_neuron.acc[2] ),
    .X(_04960_));
 sg13g2_xor2_1 _11387_ (.B(\u_toplayer.u_layer2.u_neuron.acc[2] ),
    .A(net3396),
    .X(_04961_));
 sg13g2_o21ai_1 _11388_ (.B1(_04947_),
    .Y(_04962_),
    .A1(_04944_),
    .A2(_04948_));
 sg13g2_a21oi_1 _11389_ (.A1(_04961_),
    .A2(_04962_),
    .Y(_04963_),
    .B1(net2885));
 sg13g2_o21ai_1 _11390_ (.B1(_04963_),
    .Y(_04964_),
    .A1(_04961_),
    .A2(_04962_));
 sg13g2_o21ai_1 _11391_ (.B1(_04964_),
    .Y(_04965_),
    .A1(net2861),
    .A2(_04959_));
 sg13g2_mux2_1 _11392_ (.A0(_04965_),
    .A1(net1176),
    .S(net2755),
    .X(_00679_));
 sg13g2_nand2_1 _11393_ (.Y(_04966_),
    .A(net3393),
    .B(\u_toplayer.u_layer2.u_neuron.acc[3] ));
 sg13g2_xnor2_1 _11394_ (.Y(_04967_),
    .A(net3393),
    .B(\u_toplayer.u_layer2.u_neuron.acc[3] ));
 sg13g2_a21oi_1 _11395_ (.A1(_04961_),
    .A2(_04962_),
    .Y(_04968_),
    .B1(_04960_));
 sg13g2_nand2_1 _11396_ (.Y(_04969_),
    .A(\u_toplayer.u_layer2.u_neuron.acc[3] ),
    .B(\u_toplayer.u_layer2.u_neuron.mult[3] ));
 sg13g2_xnor2_1 _11397_ (.Y(_04970_),
    .A(\u_toplayer.u_layer2.u_neuron.acc[3] ),
    .B(\u_toplayer.u_layer2.u_neuron.mult[3] ));
 sg13g2_a21oi_1 _11398_ (.A1(_04956_),
    .A2(_04958_),
    .Y(_04971_),
    .B1(_04957_));
 sg13g2_a21oi_1 _11399_ (.A1(_04970_),
    .A2(_04971_),
    .Y(_04972_),
    .B1(net2861));
 sg13g2_o21ai_1 _11400_ (.B1(_04972_),
    .Y(_04973_),
    .A1(_04970_),
    .A2(_04971_));
 sg13g2_a21oi_1 _11401_ (.A1(_04967_),
    .A2(_04968_),
    .Y(_04974_),
    .B1(net2885));
 sg13g2_o21ai_1 _11402_ (.B1(_04974_),
    .Y(_04975_),
    .A1(_04967_),
    .A2(_04968_));
 sg13g2_nor2b_1 _11403_ (.A(net2754),
    .B_N(_04975_),
    .Y(_04976_));
 sg13g2_a22oi_1 _11404_ (.Y(_00680_),
    .B1(_04973_),
    .B2(_04976_),
    .A2(net2754),
    .A1(_01101_));
 sg13g2_and2_1 _11405_ (.A(\u_toplayer.u_layer2.u_neuron.acc[4] ),
    .B(\u_toplayer.u_layer2.u_neuron.mult[4] ),
    .X(_04977_));
 sg13g2_xor2_1 _11406_ (.B(\u_toplayer.u_layer2.u_neuron.mult[4] ),
    .A(\u_toplayer.u_layer2.u_neuron.acc[4] ),
    .X(_04978_));
 sg13g2_o21ai_1 _11407_ (.B1(_04969_),
    .Y(_04979_),
    .A1(_04970_),
    .A2(_04971_));
 sg13g2_xor2_1 _11408_ (.B(_04979_),
    .A(_04978_),
    .X(_04980_));
 sg13g2_a21oi_1 _11409_ (.A1(net2858),
    .A2(_04980_),
    .Y(_04981_),
    .B1(net2754));
 sg13g2_nor2_1 _11410_ (.A(_01046_),
    .B(_01100_),
    .Y(_04982_));
 sg13g2_xor2_1 _11411_ (.B(\u_toplayer.u_layer2.u_neuron.acc[4] ),
    .A(net3390),
    .X(_04983_));
 sg13g2_o21ai_1 _11412_ (.B1(_04966_),
    .Y(_04984_),
    .A1(_04967_),
    .A2(_04968_));
 sg13g2_o21ai_1 _11413_ (.B1(net2887),
    .Y(_04985_),
    .A1(_04983_),
    .A2(_04984_));
 sg13g2_a21o_1 _11414_ (.A2(_04984_),
    .A1(_04983_),
    .B1(_04985_),
    .X(_04986_));
 sg13g2_a22oi_1 _11415_ (.Y(_00681_),
    .B1(_04981_),
    .B2(_04986_),
    .A2(net2754),
    .A1(_01100_));
 sg13g2_nor2_1 _11416_ (.A(net3063),
    .B(\u_toplayer.u_layer2.u_neuron.mult[5] ),
    .Y(_04987_));
 sg13g2_xor2_1 _11417_ (.B(\u_toplayer.u_layer2.u_neuron.mult[5] ),
    .A(net3063),
    .X(_04988_));
 sg13g2_a21oi_1 _11418_ (.A1(_04978_),
    .A2(_04979_),
    .Y(_04989_),
    .B1(_04977_));
 sg13g2_xnor2_1 _11419_ (.Y(_04990_),
    .A(_04988_),
    .B(_04989_));
 sg13g2_a21oi_1 _11420_ (.A1(_04983_),
    .A2(_04984_),
    .Y(_04991_),
    .B1(_04982_));
 sg13g2_and2_1 _11421_ (.A(net3386),
    .B(net3063),
    .X(_04992_));
 sg13g2_nor2_2 _11422_ (.A(net3386),
    .B(net3063),
    .Y(_04993_));
 sg13g2_nor3_1 _11423_ (.A(_04991_),
    .B(_04992_),
    .C(_04993_),
    .Y(_04994_));
 sg13g2_o21ai_1 _11424_ (.B1(_04991_),
    .Y(_04995_),
    .A1(_04992_),
    .A2(_04993_));
 sg13g2_nor2_1 _11425_ (.A(net2885),
    .B(_04994_),
    .Y(_04996_));
 sg13g2_a221oi_1 _11426_ (.B2(_04996_),
    .C1(net2755),
    .B1(_04995_),
    .A1(net2858),
    .Y(_04997_),
    .A2(_04990_));
 sg13g2_a21oi_1 _11427_ (.A1(_01099_),
    .A2(net2754),
    .Y(_00682_),
    .B1(_04997_));
 sg13g2_nand2_1 _11428_ (.Y(_04998_),
    .A(\u_toplayer.u_layer2.u_neuron.acc[6] ),
    .B(\u_toplayer.u_layer2.u_neuron.mult[6] ));
 sg13g2_xnor2_1 _11429_ (.Y(_04999_),
    .A(\u_toplayer.u_layer2.u_neuron.acc[6] ),
    .B(\u_toplayer.u_layer2.u_neuron.mult[6] ));
 sg13g2_a221oi_1 _11430_ (.B2(_04979_),
    .C1(_04977_),
    .B1(_04978_),
    .A1(net3063),
    .Y(_05000_),
    .A2(\u_toplayer.u_layer2.u_neuron.mult[5] ));
 sg13g2_or3_1 _11431_ (.A(_04987_),
    .B(_04999_),
    .C(_05000_),
    .X(_05001_));
 sg13g2_o21ai_1 _11432_ (.B1(_04999_),
    .Y(_05002_),
    .A1(_04987_),
    .A2(_05000_));
 sg13g2_and2_1 _11433_ (.A(_05001_),
    .B(_05002_),
    .X(_05003_));
 sg13g2_and2_1 _11434_ (.A(net3383),
    .B(\u_toplayer.u_layer2.u_neuron.acc[6] ),
    .X(_05004_));
 sg13g2_xnor2_1 _11435_ (.Y(_05005_),
    .A(net3383),
    .B(\u_toplayer.u_layer2.u_neuron.acc[6] ));
 sg13g2_a221oi_1 _11436_ (.B2(_04984_),
    .C1(_04982_),
    .B1(_04983_),
    .A1(net3386),
    .Y(_05006_),
    .A2(net3063));
 sg13g2_o21ai_1 _11437_ (.B1(_05005_),
    .Y(_05007_),
    .A1(_04993_),
    .A2(_05006_));
 sg13g2_nor3_2 _11438_ (.A(_04993_),
    .B(_05005_),
    .C(_05006_),
    .Y(_05008_));
 sg13g2_nor2_1 _11439_ (.A(net2885),
    .B(_05008_),
    .Y(_05009_));
 sg13g2_a221oi_1 _11440_ (.B2(_05009_),
    .C1(net2755),
    .B1(_05007_),
    .A1(net2858),
    .Y(_05010_),
    .A2(_05003_));
 sg13g2_a21oi_1 _11441_ (.A1(_01098_),
    .A2(net2755),
    .Y(_00683_),
    .B1(_05010_));
 sg13g2_nand2_1 _11442_ (.Y(_05011_),
    .A(net3366),
    .B(\u_toplayer.u_layer2.u_neuron.acc[7] ));
 sg13g2_xor2_1 _11443_ (.B(\u_toplayer.u_layer2.u_neuron.acc[7] ),
    .A(net3369),
    .X(_05012_));
 sg13g2_nor3_1 _11444_ (.A(_05004_),
    .B(_05008_),
    .C(_05012_),
    .Y(_05013_));
 sg13g2_o21ai_1 _11445_ (.B1(_05012_),
    .Y(_05014_),
    .A1(_05004_),
    .A2(_05008_));
 sg13g2_nand2_1 _11446_ (.Y(_05015_),
    .A(net2887),
    .B(_05014_));
 sg13g2_nor2_1 _11447_ (.A(_05013_),
    .B(_05015_),
    .Y(_05016_));
 sg13g2_and2_1 _11448_ (.A(\u_toplayer.u_layer2.u_neuron.acc[7] ),
    .B(\u_toplayer.u_layer2.u_neuron.mult[7] ),
    .X(_05017_));
 sg13g2_xnor2_1 _11449_ (.Y(_05018_),
    .A(\u_toplayer.u_layer2.u_neuron.acc[7] ),
    .B(\u_toplayer.u_layer2.u_neuron.mult[7] ));
 sg13g2_and3_1 _11450_ (.X(_05019_),
    .A(_04998_),
    .B(_05001_),
    .C(_05018_));
 sg13g2_a21oi_2 _11451_ (.B1(_05018_),
    .Y(_05020_),
    .A2(_05001_),
    .A1(_04998_));
 sg13g2_nor3_1 _11452_ (.A(net2861),
    .B(_05019_),
    .C(_05020_),
    .Y(_05021_));
 sg13g2_nor3_1 _11453_ (.A(net2755),
    .B(_05016_),
    .C(_05021_),
    .Y(_05022_));
 sg13g2_a21oi_1 _11454_ (.A1(_01097_),
    .A2(net2755),
    .Y(_00684_),
    .B1(_05022_));
 sg13g2_nand2_1 _11455_ (.Y(_05023_),
    .A(\u_toplayer.u_layer2.u_neuron.acc[8] ),
    .B(\u_toplayer.u_layer2.u_neuron.mult[8] ));
 sg13g2_xor2_1 _11456_ (.B(\u_toplayer.u_layer2.u_neuron.mult[8] ),
    .A(\u_toplayer.u_layer2.u_neuron.acc[8] ),
    .X(_05024_));
 sg13g2_inv_1 _11457_ (.Y(_05025_),
    .A(_05024_));
 sg13g2_nor3_1 _11458_ (.A(_05017_),
    .B(_05020_),
    .C(_05024_),
    .Y(_05026_));
 sg13g2_o21ai_1 _11459_ (.B1(_05024_),
    .Y(_05027_),
    .A1(_05017_),
    .A2(_05020_));
 sg13g2_nor2b_1 _11460_ (.A(_05026_),
    .B_N(_05027_),
    .Y(_05028_));
 sg13g2_and2_1 _11461_ (.A(_05011_),
    .B(_05014_),
    .X(_05029_));
 sg13g2_nand2_1 _11462_ (.Y(_05030_),
    .A(net3366),
    .B(\u_toplayer.u_layer2.u_neuron.acc[8] ));
 sg13g2_xnor2_1 _11463_ (.Y(_05031_),
    .A(net3366),
    .B(\u_toplayer.u_layer2.u_neuron.acc[8] ));
 sg13g2_or2_1 _11464_ (.X(_05032_),
    .B(_05031_),
    .A(_05029_));
 sg13g2_a21oi_1 _11465_ (.A1(_05029_),
    .A2(_05031_),
    .Y(_05033_),
    .B1(net2884));
 sg13g2_a221oi_1 _11466_ (.B2(_05033_),
    .C1(net2751),
    .B1(_05032_),
    .A1(net2858),
    .Y(_05034_),
    .A2(_05028_));
 sg13g2_a21oi_1 _11467_ (.A1(_01109_),
    .A2(net2755),
    .Y(_00685_),
    .B1(_05034_));
 sg13g2_nor2_1 _11468_ (.A(\u_toplayer.u_layer2.u_neuron.acc[9] ),
    .B(\u_toplayer.u_layer2.u_neuron.mult[9] ),
    .Y(_05035_));
 sg13g2_nand2_1 _11469_ (.Y(_05036_),
    .A(\u_toplayer.u_layer2.u_neuron.acc[9] ),
    .B(\u_toplayer.u_layer2.u_neuron.mult[9] ));
 sg13g2_nand2b_1 _11470_ (.Y(_05037_),
    .B(_05036_),
    .A_N(_05035_));
 sg13g2_and2_1 _11471_ (.A(_05023_),
    .B(_05027_),
    .X(_05038_));
 sg13g2_a21oi_1 _11472_ (.A1(_05037_),
    .A2(_05038_),
    .Y(_05039_),
    .B1(net2861));
 sg13g2_o21ai_1 _11473_ (.B1(_05039_),
    .Y(_05040_),
    .A1(_05037_),
    .A2(_05038_));
 sg13g2_xor2_1 _11474_ (.B(\u_toplayer.u_layer2.u_neuron.acc[9] ),
    .A(net3366),
    .X(_05041_));
 sg13g2_inv_1 _11475_ (.Y(_05042_),
    .A(_05041_));
 sg13g2_a21oi_1 _11476_ (.A1(_05030_),
    .A2(_05032_),
    .Y(_05043_),
    .B1(_05042_));
 sg13g2_nand3_1 _11477_ (.B(_05032_),
    .C(_05042_),
    .A(_05030_),
    .Y(_05044_));
 sg13g2_nor2_1 _11478_ (.A(net2884),
    .B(_05043_),
    .Y(_05045_));
 sg13g2_a21oi_1 _11479_ (.A1(_05044_),
    .A2(_05045_),
    .Y(_05046_),
    .B1(net2751));
 sg13g2_a22oi_1 _11480_ (.Y(_00686_),
    .B1(_05040_),
    .B2(_05046_),
    .A2(net2751),
    .A1(_01108_));
 sg13g2_xor2_1 _11481_ (.B(\u_toplayer.u_layer2.u_neuron.mult[10] ),
    .A(net3062),
    .X(_05047_));
 sg13g2_inv_1 _11482_ (.Y(_05048_),
    .A(_05047_));
 sg13g2_nor2_1 _11483_ (.A(_05025_),
    .B(_05037_),
    .Y(_05049_));
 sg13g2_o21ai_1 _11484_ (.B1(_05049_),
    .Y(_05050_),
    .A1(_05017_),
    .A2(_05020_));
 sg13g2_o21ai_1 _11485_ (.B1(_05036_),
    .Y(_05051_),
    .A1(_05023_),
    .A2(_05035_));
 sg13g2_nand2b_1 _11486_ (.Y(_05052_),
    .B(_05050_),
    .A_N(_05051_));
 sg13g2_and2_1 _11487_ (.A(_05047_),
    .B(_05052_),
    .X(_05053_));
 sg13g2_nor2_1 _11488_ (.A(net2861),
    .B(_05053_),
    .Y(_05054_));
 sg13g2_o21ai_1 _11489_ (.B1(_05054_),
    .Y(_05055_),
    .A1(_05047_),
    .A2(_05052_));
 sg13g2_xnor2_1 _11490_ (.Y(_05056_),
    .A(net3366),
    .B(net3062));
 sg13g2_o21ai_1 _11491_ (.B1(net3364),
    .Y(_05057_),
    .A1(\u_toplayer.u_layer2.u_neuron.acc[9] ),
    .A2(\u_toplayer.u_layer2.u_neuron.acc[8] ));
 sg13g2_nand2b_1 _11492_ (.Y(_05058_),
    .B(_05041_),
    .A_N(_05031_));
 sg13g2_o21ai_1 _11493_ (.B1(_05057_),
    .Y(_05059_),
    .A1(_05029_),
    .A2(_05058_));
 sg13g2_nor2b_1 _11494_ (.A(_05056_),
    .B_N(_05059_),
    .Y(_05060_));
 sg13g2_xnor2_1 _11495_ (.Y(_05061_),
    .A(_05056_),
    .B(_05059_));
 sg13g2_a21oi_1 _11496_ (.A1(net2886),
    .A2(_05061_),
    .Y(_05062_),
    .B1(net2750));
 sg13g2_a22oi_1 _11497_ (.Y(_00687_),
    .B1(_05055_),
    .B2(_05062_),
    .A2(net2751),
    .A1(_01107_));
 sg13g2_xnor2_1 _11498_ (.Y(_05063_),
    .A(\u_toplayer.u_layer2.u_neuron.acc[11] ),
    .B(\u_toplayer.u_layer2.u_neuron.mult[11] ));
 sg13g2_a21oi_1 _11499_ (.A1(net3062),
    .A2(\u_toplayer.u_layer2.u_neuron.mult[10] ),
    .Y(_05064_),
    .B1(_05053_));
 sg13g2_o21ai_1 _11500_ (.B1(net2858),
    .Y(_05065_),
    .A1(_05063_),
    .A2(_05064_));
 sg13g2_a21oi_1 _11501_ (.A1(_05063_),
    .A2(_05064_),
    .Y(_05066_),
    .B1(_05065_));
 sg13g2_xnor2_1 _11502_ (.Y(_05067_),
    .A(net3364),
    .B(\u_toplayer.u_layer2.u_neuron.acc[11] ));
 sg13g2_a21oi_1 _11503_ (.A1(net3366),
    .A2(net3062),
    .Y(_05068_),
    .B1(_05060_));
 sg13g2_o21ai_1 _11504_ (.B1(net2886),
    .Y(_05069_),
    .A1(_05067_),
    .A2(_05068_));
 sg13g2_a21oi_1 _11505_ (.A1(_05067_),
    .A2(_05068_),
    .Y(_05070_),
    .B1(_05069_));
 sg13g2_nor3_1 _11506_ (.A(net2750),
    .B(_05066_),
    .C(_05070_),
    .Y(_05071_));
 sg13g2_a21oi_1 _11507_ (.A1(_01106_),
    .A2(net2750),
    .Y(_00688_),
    .B1(_05071_));
 sg13g2_nand2_1 _11508_ (.Y(_05072_),
    .A(net3061),
    .B(\u_toplayer.u_layer2.u_neuron.mult[12] ));
 sg13g2_xnor2_1 _11509_ (.Y(_05073_),
    .A(net3061),
    .B(\u_toplayer.u_layer2.u_neuron.mult[12] ));
 sg13g2_a22oi_1 _11510_ (.Y(_05074_),
    .B1(\u_toplayer.u_layer2.u_neuron.mult[11] ),
    .B2(\u_toplayer.u_layer2.u_neuron.acc[11] ),
    .A2(\u_toplayer.u_layer2.u_neuron.mult[10] ),
    .A1(net3062));
 sg13g2_a21oi_1 _11511_ (.A1(_01106_),
    .A2(_01148_),
    .Y(_05075_),
    .B1(_05074_));
 sg13g2_nor2_1 _11512_ (.A(_05048_),
    .B(_05063_),
    .Y(_05076_));
 sg13g2_nor2_1 _11513_ (.A(_05051_),
    .B(_05075_),
    .Y(_05077_));
 sg13g2_nor2_1 _11514_ (.A(_05075_),
    .B(_05076_),
    .Y(_05078_));
 sg13g2_a21oi_2 _11515_ (.B1(_05078_),
    .Y(_05079_),
    .A2(_05077_),
    .A1(_05050_));
 sg13g2_nand2b_1 _11516_ (.Y(_05080_),
    .B(_05079_),
    .A_N(_05073_));
 sg13g2_nand2b_1 _11517_ (.Y(_05081_),
    .B(_05073_),
    .A_N(_05079_));
 sg13g2_nand3_1 _11518_ (.B(_05080_),
    .C(_05081_),
    .A(net2858),
    .Y(_05082_));
 sg13g2_xor2_1 _11519_ (.B(\u_toplayer.u_layer2.u_neuron.acc[12] ),
    .A(net3365),
    .X(_05083_));
 sg13g2_or3_1 _11520_ (.A(_05056_),
    .B(_05058_),
    .C(_05067_),
    .X(_05084_));
 sg13g2_a21oi_1 _11521_ (.A1(_05011_),
    .A2(_05014_),
    .Y(_05085_),
    .B1(_05084_));
 sg13g2_o21ai_1 _11522_ (.B1(net3364),
    .Y(_05086_),
    .A1(\u_toplayer.u_layer2.u_neuron.acc[11] ),
    .A2(net3062));
 sg13g2_nand3b_1 _11523_ (.B(_05086_),
    .C(_05057_),
    .Y(_05087_),
    .A_N(_05085_));
 sg13g2_and2_1 _11524_ (.A(_05083_),
    .B(_05087_),
    .X(_05088_));
 sg13g2_o21ai_1 _11525_ (.B1(net2886),
    .Y(_05089_),
    .A1(_05083_),
    .A2(_05087_));
 sg13g2_o21ai_1 _11526_ (.B1(_05082_),
    .Y(_05090_),
    .A1(_05088_),
    .A2(_05089_));
 sg13g2_mux2_1 _11527_ (.A0(_05090_),
    .A1(net3061),
    .S(net2750),
    .X(_00689_));
 sg13g2_nor2_1 _11528_ (.A(\u_toplayer.u_layer2.u_neuron.acc[13] ),
    .B(\u_toplayer.u_layer2.u_neuron.mult[13] ),
    .Y(_05091_));
 sg13g2_xnor2_1 _11529_ (.Y(_05092_),
    .A(\u_toplayer.u_layer2.u_neuron.acc[13] ),
    .B(\u_toplayer.u_layer2.u_neuron.mult[13] ));
 sg13g2_a21oi_1 _11530_ (.A1(_05072_),
    .A2(_05080_),
    .Y(_05093_),
    .B1(_05092_));
 sg13g2_nand3_1 _11531_ (.B(_05080_),
    .C(_05092_),
    .A(_05072_),
    .Y(_05094_));
 sg13g2_nand2_1 _11532_ (.Y(_05095_),
    .A(net2858),
    .B(_05094_));
 sg13g2_xor2_1 _11533_ (.B(\u_toplayer.u_layer2.u_neuron.acc[13] ),
    .A(net3364),
    .X(_05096_));
 sg13g2_a21o_1 _11534_ (.A2(net3061),
    .A1(net3365),
    .B1(_05088_),
    .X(_05097_));
 sg13g2_a21oi_1 _11535_ (.A1(_05096_),
    .A2(_05097_),
    .Y(_05098_),
    .B1(net2884));
 sg13g2_o21ai_1 _11536_ (.B1(_05098_),
    .Y(_05099_),
    .A1(_05096_),
    .A2(_05097_));
 sg13g2_o21ai_1 _11537_ (.B1(_05099_),
    .Y(_05100_),
    .A1(_05093_),
    .A2(_05095_));
 sg13g2_mux2_1 _11538_ (.A0(_05100_),
    .A1(net1159),
    .S(net2750),
    .X(_00690_));
 sg13g2_xnor2_1 _11539_ (.Y(_05101_),
    .A(net3060),
    .B(\u_toplayer.u_layer2.u_neuron.mult[14] ));
 sg13g2_a22oi_1 _11540_ (.Y(_05102_),
    .B1(\u_toplayer.u_layer2.u_neuron.mult[13] ),
    .B2(\u_toplayer.u_layer2.u_neuron.acc[13] ),
    .A2(\u_toplayer.u_layer2.u_neuron.mult[12] ),
    .A1(net3061));
 sg13g2_a21o_1 _11541_ (.A2(_05102_),
    .A1(_05080_),
    .B1(_05091_),
    .X(_05103_));
 sg13g2_nor2_1 _11542_ (.A(_05101_),
    .B(_05103_),
    .Y(_05104_));
 sg13g2_a21oi_1 _11543_ (.A1(_05101_),
    .A2(_05103_),
    .Y(_05105_),
    .B1(net2860));
 sg13g2_nand2b_1 _11544_ (.Y(_05106_),
    .B(_05105_),
    .A_N(_05104_));
 sg13g2_xnor2_1 _11545_ (.Y(_05107_),
    .A(net3364),
    .B(\u_toplayer.u_layer2.u_neuron.acc[14] ));
 sg13g2_o21ai_1 _11546_ (.B1(net3365),
    .Y(_05108_),
    .A1(\u_toplayer.u_layer2.u_neuron.acc[13] ),
    .A2(net3061));
 sg13g2_nand2_1 _11547_ (.Y(_05109_),
    .A(_05083_),
    .B(_05096_));
 sg13g2_nand2_1 _11548_ (.Y(_05110_),
    .A(_05088_),
    .B(_05096_));
 sg13g2_a21oi_1 _11549_ (.A1(_05108_),
    .A2(_05110_),
    .Y(_05111_),
    .B1(_05107_));
 sg13g2_and3_1 _11550_ (.X(_05112_),
    .A(_05107_),
    .B(_05108_),
    .C(_05110_));
 sg13g2_nor3_1 _11551_ (.A(net2884),
    .B(_05111_),
    .C(_05112_),
    .Y(_05113_));
 sg13g2_nor2_1 _11552_ (.A(net2750),
    .B(_05113_),
    .Y(_05114_));
 sg13g2_a22oi_1 _11553_ (.Y(_00691_),
    .B1(_05106_),
    .B2(_05114_),
    .A2(net2750),
    .A1(_01105_));
 sg13g2_nand2_1 _11554_ (.Y(_05115_),
    .A(_01104_),
    .B(_01149_));
 sg13g2_xnor2_1 _11555_ (.Y(_05116_),
    .A(\u_toplayer.u_layer2.u_neuron.acc[15] ),
    .B(net3194));
 sg13g2_a21oi_1 _11556_ (.A1(net3060),
    .A2(\u_toplayer.u_layer2.u_neuron.mult[14] ),
    .Y(_05117_),
    .B1(_05104_));
 sg13g2_a21oi_1 _11557_ (.A1(_05116_),
    .A2(_05117_),
    .Y(_05118_),
    .B1(net2860));
 sg13g2_o21ai_1 _11558_ (.B1(_05118_),
    .Y(_05119_),
    .A1(_05116_),
    .A2(_05117_));
 sg13g2_xnor2_1 _11559_ (.Y(_05120_),
    .A(net3364),
    .B(\u_toplayer.u_layer2.u_neuron.acc[15] ));
 sg13g2_a21oi_1 _11560_ (.A1(net3364),
    .A2(net3060),
    .Y(_05121_),
    .B1(_05111_));
 sg13g2_o21ai_1 _11561_ (.B1(net2886),
    .Y(_05122_),
    .A1(_05120_),
    .A2(_05121_));
 sg13g2_a21oi_1 _11562_ (.A1(_05120_),
    .A2(_05121_),
    .Y(_05123_),
    .B1(_05122_));
 sg13g2_nor2_1 _11563_ (.A(net2751),
    .B(_05123_),
    .Y(_05124_));
 sg13g2_a22oi_1 _11564_ (.Y(_00692_),
    .B1(_05119_),
    .B2(_05124_),
    .A2(net2750),
    .A1(_01104_));
 sg13g2_nor4_1 _11565_ (.A(_05073_),
    .B(_05092_),
    .C(_05101_),
    .D(_05116_),
    .Y(_05125_));
 sg13g2_nor4_1 _11566_ (.A(_05091_),
    .B(_05101_),
    .C(_05102_),
    .D(_05116_),
    .Y(_05126_));
 sg13g2_a22oi_1 _11567_ (.Y(_05127_),
    .B1(net3194),
    .B2(\u_toplayer.u_layer2.u_neuron.acc[15] ),
    .A2(\u_toplayer.u_layer2.u_neuron.mult[14] ),
    .A1(net3060));
 sg13g2_inv_1 _11568_ (.Y(_05128_),
    .A(_05127_));
 sg13g2_a221oi_1 _11569_ (.B2(_05115_),
    .C1(_05126_),
    .B1(_05128_),
    .A1(_05079_),
    .Y(_05129_),
    .A2(_05125_));
 sg13g2_xnor2_1 _11570_ (.Y(_05130_),
    .A(net3059),
    .B(net3193));
 sg13g2_nor2_1 _11571_ (.A(_05129_),
    .B(_05130_),
    .Y(_05131_));
 sg13g2_a21oi_1 _11572_ (.A1(_05129_),
    .A2(_05130_),
    .Y(_05132_),
    .B1(net2860));
 sg13g2_nand2b_1 _11573_ (.Y(_05133_),
    .B(_05132_),
    .A_N(_05131_));
 sg13g2_nor3_1 _11574_ (.A(_05107_),
    .B(_05109_),
    .C(_05120_),
    .Y(_05134_));
 sg13g2_o21ai_1 _11575_ (.B1(net3364),
    .Y(_05135_),
    .A1(\u_toplayer.u_layer2.u_neuron.acc[15] ),
    .A2(net3060));
 sg13g2_nand4_1 _11576_ (.B(_05086_),
    .C(_05108_),
    .A(_05057_),
    .Y(_05136_),
    .D(_05135_));
 sg13g2_a21oi_2 _11577_ (.B1(_05136_),
    .Y(_05137_),
    .A2(_05134_),
    .A1(_05085_));
 sg13g2_xnor2_1 _11578_ (.Y(_05138_),
    .A(net3367),
    .B(net3059));
 sg13g2_nor2_1 _11579_ (.A(_05137_),
    .B(_05138_),
    .Y(_05139_));
 sg13g2_nand2_1 _11580_ (.Y(_05140_),
    .A(_05137_),
    .B(_05138_));
 sg13g2_nor2_1 _11581_ (.A(net2884),
    .B(_05139_),
    .Y(_05141_));
 sg13g2_a21oi_1 _11582_ (.A1(_05140_),
    .A2(_05141_),
    .Y(_05142_),
    .B1(net2753));
 sg13g2_a22oi_1 _11583_ (.Y(_00693_),
    .B1(_05133_),
    .B2(_05142_),
    .A2(net2753),
    .A1(_01116_));
 sg13g2_xnor2_1 _11584_ (.Y(_05143_),
    .A(\u_toplayer.u_layer2.u_neuron.acc[17] ),
    .B(net3193));
 sg13g2_a21oi_1 _11585_ (.A1(net3059),
    .A2(net3193),
    .Y(_05144_),
    .B1(_05131_));
 sg13g2_a21oi_1 _11586_ (.A1(_05143_),
    .A2(_05144_),
    .Y(_05145_),
    .B1(net2860));
 sg13g2_o21ai_1 _11587_ (.B1(_05145_),
    .Y(_05146_),
    .A1(_05143_),
    .A2(_05144_));
 sg13g2_xor2_1 _11588_ (.B(\u_toplayer.u_layer2.u_neuron.acc[17] ),
    .A(net3367),
    .X(_05147_));
 sg13g2_a21o_1 _11589_ (.A2(net3059),
    .A1(net3367),
    .B1(_05139_),
    .X(_05148_));
 sg13g2_o21ai_1 _11590_ (.B1(net2886),
    .Y(_05149_),
    .A1(_05147_),
    .A2(_05148_));
 sg13g2_a21oi_1 _11591_ (.A1(_05147_),
    .A2(_05148_),
    .Y(_05150_),
    .B1(_05149_));
 sg13g2_nor2_1 _11592_ (.A(net2753),
    .B(_05150_),
    .Y(_05151_));
 sg13g2_a22oi_1 _11593_ (.Y(_00694_),
    .B1(_05146_),
    .B2(_05151_),
    .A2(net2753),
    .A1(_01115_));
 sg13g2_xor2_1 _11594_ (.B(net3192),
    .A(\u_toplayer.u_layer2.u_neuron.acc[18] ),
    .X(_05152_));
 sg13g2_nor3_2 _11595_ (.A(_05129_),
    .B(_05130_),
    .C(_05143_),
    .Y(_05153_));
 sg13g2_o21ai_1 _11596_ (.B1(net3193),
    .Y(_05154_),
    .A1(\u_toplayer.u_layer2.u_neuron.acc[17] ),
    .A2(\u_toplayer.u_layer2.u_neuron.acc[16] ));
 sg13g2_inv_1 _11597_ (.Y(_05155_),
    .A(_05154_));
 sg13g2_o21ai_1 _11598_ (.B1(_05152_),
    .Y(_05156_),
    .A1(_05153_),
    .A2(_05155_));
 sg13g2_nor3_1 _11599_ (.A(_05152_),
    .B(_05153_),
    .C(_05155_),
    .Y(_05157_));
 sg13g2_nor2_1 _11600_ (.A(net2860),
    .B(_05157_),
    .Y(_05158_));
 sg13g2_xnor2_1 _11601_ (.Y(_05159_),
    .A(net3367),
    .B(\u_toplayer.u_layer2.u_neuron.acc[18] ));
 sg13g2_nand2b_1 _11602_ (.Y(_05160_),
    .B(_05147_),
    .A_N(_05138_));
 sg13g2_nand2_1 _11603_ (.Y(_05161_),
    .A(_05139_),
    .B(_05147_));
 sg13g2_o21ai_1 _11604_ (.B1(net3367),
    .Y(_05162_),
    .A1(\u_toplayer.u_layer2.u_neuron.acc[17] ),
    .A2(net3059));
 sg13g2_a21oi_1 _11605_ (.A1(_05161_),
    .A2(_05162_),
    .Y(_05163_),
    .B1(_05159_));
 sg13g2_nand3_1 _11606_ (.B(_05161_),
    .C(_05162_),
    .A(_05159_),
    .Y(_05164_));
 sg13g2_nor2_1 _11607_ (.A(net2884),
    .B(_05163_),
    .Y(_05165_));
 sg13g2_a221oi_1 _11608_ (.B2(_05165_),
    .C1(net2753),
    .B1(_05164_),
    .A1(_05156_),
    .Y(_05166_),
    .A2(_05158_));
 sg13g2_a21oi_1 _11609_ (.A1(_01114_),
    .A2(net2752),
    .Y(_00695_),
    .B1(_05166_));
 sg13g2_xor2_1 _11610_ (.B(net3192),
    .A(\u_toplayer.u_layer2.u_neuron.acc[19] ),
    .X(_05167_));
 sg13g2_o21ai_1 _11611_ (.B1(_05156_),
    .Y(_05168_),
    .A1(_01114_),
    .A2(_01149_));
 sg13g2_a21oi_1 _11612_ (.A1(_05167_),
    .A2(_05168_),
    .Y(_05169_),
    .B1(net2860));
 sg13g2_o21ai_1 _11613_ (.B1(_05169_),
    .Y(_05170_),
    .A1(_05167_),
    .A2(_05168_));
 sg13g2_xnor2_1 _11614_ (.Y(_05171_),
    .A(net3367),
    .B(\u_toplayer.u_layer2.u_neuron.acc[19] ));
 sg13g2_a21oi_1 _11615_ (.A1(net3367),
    .A2(\u_toplayer.u_layer2.u_neuron.acc[18] ),
    .Y(_05172_),
    .B1(_05163_));
 sg13g2_o21ai_1 _11616_ (.B1(net2887),
    .Y(_05173_),
    .A1(_05171_),
    .A2(_05172_));
 sg13g2_a21oi_1 _11617_ (.A1(_05171_),
    .A2(_05172_),
    .Y(_05174_),
    .B1(_05173_));
 sg13g2_nor2_1 _11618_ (.A(net2753),
    .B(_05174_),
    .Y(_05175_));
 sg13g2_a22oi_1 _11619_ (.Y(_00696_),
    .B1(_05170_),
    .B2(_05175_),
    .A2(net2752),
    .A1(_01113_));
 sg13g2_and2_1 _11620_ (.A(_05152_),
    .B(_05167_),
    .X(_05176_));
 sg13g2_o21ai_1 _11621_ (.B1(net3192),
    .Y(_05177_),
    .A1(\u_toplayer.u_layer2.u_neuron.acc[19] ),
    .A2(\u_toplayer.u_layer2.u_neuron.acc[18] ));
 sg13g2_nand2_1 _11622_ (.Y(_05178_),
    .A(_05154_),
    .B(_05177_));
 sg13g2_a21o_1 _11623_ (.A2(_05176_),
    .A1(_05153_),
    .B1(_05178_),
    .X(_05179_));
 sg13g2_xor2_1 _11624_ (.B(net3192),
    .A(net3058),
    .X(_05180_));
 sg13g2_and2_1 _11625_ (.A(_05179_),
    .B(_05180_),
    .X(_05181_));
 sg13g2_o21ai_1 _11626_ (.B1(net2859),
    .Y(_05182_),
    .A1(_05179_),
    .A2(_05180_));
 sg13g2_nor2_1 _11627_ (.A(_05181_),
    .B(_05182_),
    .Y(_05183_));
 sg13g2_xor2_1 _11628_ (.B(net3058),
    .A(net3368),
    .X(_05184_));
 sg13g2_nor4_1 _11629_ (.A(_05137_),
    .B(_05159_),
    .C(_05160_),
    .D(_05171_),
    .Y(_05185_));
 sg13g2_o21ai_1 _11630_ (.B1(net3367),
    .Y(_05186_),
    .A1(\u_toplayer.u_layer2.u_neuron.acc[19] ),
    .A2(\u_toplayer.u_layer2.u_neuron.acc[18] ));
 sg13g2_nand2_1 _11631_ (.Y(_05187_),
    .A(_05162_),
    .B(_05186_));
 sg13g2_nor2_1 _11632_ (.A(_05185_),
    .B(_05187_),
    .Y(_05188_));
 sg13g2_nor2b_1 _11633_ (.A(_05188_),
    .B_N(_05184_),
    .Y(_05189_));
 sg13g2_o21ai_1 _11634_ (.B1(_05184_),
    .Y(_05190_),
    .A1(_05185_),
    .A2(_05187_));
 sg13g2_nand2b_1 _11635_ (.Y(_05191_),
    .B(_05188_),
    .A_N(_05184_));
 sg13g2_nor2_1 _11636_ (.A(net2884),
    .B(_05189_),
    .Y(_05192_));
 sg13g2_a21o_1 _11637_ (.A2(_05192_),
    .A1(_05191_),
    .B1(_05183_),
    .X(_05193_));
 sg13g2_mux2_1 _11638_ (.A0(_05193_),
    .A1(net3058),
    .S(net2752),
    .X(_00697_));
 sg13g2_xor2_1 _11639_ (.B(net3192),
    .A(\u_toplayer.u_layer2.u_neuron.acc[21] ),
    .X(_05194_));
 sg13g2_a21oi_1 _11640_ (.A1(net3058),
    .A2(net3192),
    .Y(_05195_),
    .B1(_05181_));
 sg13g2_nand2b_1 _11641_ (.Y(_05196_),
    .B(_05194_),
    .A_N(_05195_));
 sg13g2_nand2b_1 _11642_ (.Y(_05197_),
    .B(_05195_),
    .A_N(_05194_));
 sg13g2_nand3_1 _11643_ (.B(_05196_),
    .C(_05197_),
    .A(net2859),
    .Y(_05198_));
 sg13g2_xnor2_1 _11644_ (.Y(_05199_),
    .A(net3368),
    .B(\u_toplayer.u_layer2.u_neuron.acc[21] ));
 sg13g2_a21oi_1 _11645_ (.A1(net3368),
    .A2(net3058),
    .Y(_05200_),
    .B1(_05189_));
 sg13g2_o21ai_1 _11646_ (.B1(net2886),
    .Y(_05201_),
    .A1(_05199_),
    .A2(_05200_));
 sg13g2_a21oi_1 _11647_ (.A1(_05199_),
    .A2(_05200_),
    .Y(_05202_),
    .B1(_05201_));
 sg13g2_nor2_1 _11648_ (.A(net2752),
    .B(_05202_),
    .Y(_05203_));
 sg13g2_a22oi_1 _11649_ (.Y(_00698_),
    .B1(_05198_),
    .B2(_05203_),
    .A2(net2753),
    .A1(_01112_));
 sg13g2_nor2_1 _11650_ (.A(_01111_),
    .B(_01149_),
    .Y(_05204_));
 sg13g2_xnor2_1 _11651_ (.Y(_05205_),
    .A(\u_toplayer.u_layer2.u_neuron.acc[22] ),
    .B(net3193));
 sg13g2_nand3_1 _11652_ (.B(_05180_),
    .C(_05194_),
    .A(_05179_),
    .Y(_05206_));
 sg13g2_o21ai_1 _11653_ (.B1(net3192),
    .Y(_05207_),
    .A1(\u_toplayer.u_layer2.u_neuron.acc[21] ),
    .A2(net3058));
 sg13g2_nand3_1 _11654_ (.B(_05206_),
    .C(_05207_),
    .A(_05205_),
    .Y(_05208_));
 sg13g2_a21oi_1 _11655_ (.A1(_05206_),
    .A2(_05207_),
    .Y(_05209_),
    .B1(_05205_));
 sg13g2_nor2_1 _11656_ (.A(net2860),
    .B(_05209_),
    .Y(_05210_));
 sg13g2_o21ai_1 _11657_ (.B1(net3368),
    .Y(_05211_),
    .A1(\u_toplayer.u_layer2.u_neuron.acc[21] ),
    .A2(\u_toplayer.u_layer2.u_neuron.acc[20] ));
 sg13g2_o21ai_1 _11658_ (.B1(_05211_),
    .Y(_05212_),
    .A1(_05190_),
    .A2(_05199_));
 sg13g2_and2_1 _11659_ (.A(net3368),
    .B(\u_toplayer.u_layer2.u_neuron.acc[22] ),
    .X(_05213_));
 sg13g2_or2_1 _11660_ (.X(_05214_),
    .B(\u_toplayer.u_layer2.u_neuron.acc[22] ),
    .A(net3368));
 sg13g2_nand2b_1 _11661_ (.Y(_05215_),
    .B(_05214_),
    .A_N(_05213_));
 sg13g2_xnor2_1 _11662_ (.Y(_05216_),
    .A(_05212_),
    .B(_05215_));
 sg13g2_a221oi_1 _11663_ (.B2(net2886),
    .C1(net2752),
    .B1(_05216_),
    .A1(_05208_),
    .Y(_05217_),
    .A2(_05210_));
 sg13g2_a21oi_1 _11664_ (.A1(_01111_),
    .A2(net2752),
    .Y(_00699_),
    .B1(_05217_));
 sg13g2_xor2_1 _11665_ (.B(net3192),
    .A(\u_toplayer.u_layer2.u_neuron.acc[23] ),
    .X(_05218_));
 sg13g2_or3_1 _11666_ (.A(_05204_),
    .B(_05209_),
    .C(_05218_),
    .X(_05219_));
 sg13g2_o21ai_1 _11667_ (.B1(_05218_),
    .Y(_05220_),
    .A1(_05204_),
    .A2(_05209_));
 sg13g2_nand3_1 _11668_ (.B(_05219_),
    .C(_05220_),
    .A(net2859),
    .Y(_05221_));
 sg13g2_a21oi_1 _11669_ (.A1(_05212_),
    .A2(_05214_),
    .Y(_05222_),
    .B1(_05213_));
 sg13g2_xnor2_1 _11670_ (.Y(_05223_),
    .A(net3368),
    .B(\u_toplayer.u_layer2.u_neuron.acc[23] ));
 sg13g2_o21ai_1 _11671_ (.B1(net2886),
    .Y(_05224_),
    .A1(_05222_),
    .A2(_05223_));
 sg13g2_a21oi_1 _11672_ (.A1(_05222_),
    .A2(_05223_),
    .Y(_05225_),
    .B1(_05224_));
 sg13g2_nor2_1 _11673_ (.A(net2752),
    .B(_05225_),
    .Y(_05226_));
 sg13g2_a22oi_1 _11674_ (.Y(_00700_),
    .B1(_05221_),
    .B2(_05226_),
    .A2(net2752),
    .A1(_01110_));
 sg13g2_nand2_2 _11675_ (.Y(_05227_),
    .A(net921),
    .B(net987));
 sg13g2_nor4_1 _11676_ (.A(\u_toplayer.u_layer1.statel1[5] ),
    .B(\u_toplayer.u_layer1.statel1[4] ),
    .C(\u_toplayer.u_layer1.statel1[3] ),
    .D(\u_toplayer.u_layer1.statel1[2] ),
    .Y(_05228_));
 sg13g2_nand3_1 _11677_ (.B(_01028_),
    .C(_05228_),
    .A(_01027_),
    .Y(_05229_));
 sg13g2_inv_1 _11678_ (.Y(_05230_),
    .A(_05229_));
 sg13g2_a21oi_1 _11679_ (.A1(_05227_),
    .A2(_05230_),
    .Y(_05231_),
    .B1(_00029_));
 sg13g2_nor4_2 _11680_ (.A(\u_toplayer.done_layer1 ),
    .B(_01026_),
    .C(_05227_),
    .Y(_05232_),
    .D(_05229_));
 sg13g2_and2_1 _11681_ (.A(_05231_),
    .B(_05232_),
    .X(_05233_));
 sg13g2_mux2_1 _11682_ (.A0(net3057),
    .A1(net597),
    .S(_05233_),
    .X(_00701_));
 sg13g2_nand2_2 _11683_ (.Y(_05234_),
    .A(net3057),
    .B(\u_toplayer.u_layer1.neuron_index[1] ));
 sg13g2_nand3_1 _11684_ (.B(net1146),
    .C(net2818),
    .A(net3057),
    .Y(_05235_));
 sg13g2_a21o_1 _11685_ (.A2(net2818),
    .A1(net3057),
    .B1(net1146),
    .X(_05236_));
 sg13g2_and2_1 _11686_ (.A(_05235_),
    .B(_05236_),
    .X(_00702_));
 sg13g2_and3_1 _11687_ (.X(_05237_),
    .A(net3057),
    .B(\u_toplayer.u_layer1.neuron_index[1] ),
    .C(net3055));
 sg13g2_xnor2_1 _11688_ (.Y(_00703_),
    .A(net3055),
    .B(net1147));
 sg13g2_nand3_1 _11689_ (.B(net2818),
    .C(_05237_),
    .A(net3053),
    .Y(_05238_));
 sg13g2_a21o_1 _11690_ (.A2(net2945),
    .A1(net2818),
    .B1(net3053),
    .X(_05239_));
 sg13g2_and2_1 _11691_ (.A(_05238_),
    .B(_05239_),
    .X(_00704_));
 sg13g2_nand4_1 _11692_ (.B(\u_toplayer.u_layer1.neuron_index[4] ),
    .C(net2818),
    .A(net3053),
    .Y(_05240_),
    .D(net2947));
 sg13g2_xnor2_1 _11693_ (.Y(_00705_),
    .A(net1028),
    .B(_05238_));
 sg13g2_or2_2 _11694_ (.X(_05241_),
    .B(_05240_),
    .A(\u_toplayer.u_layer1.neuron_index[5] ));
 sg13g2_xnor2_1 _11695_ (.Y(_00706_),
    .A(net1010),
    .B(_05240_));
 sg13g2_nor3_1 _11696_ (.A(\u_toplayer.done_layer3 ),
    .B(net126),
    .C(_01025_),
    .Y(_00707_));
 sg13g2_a21o_1 _11697_ (.A2(net907),
    .A1(net126),
    .B1(\u_toplayer.done_layer3 ),
    .X(_00708_));
 sg13g2_nand3_1 _11698_ (.B(_01384_),
    .C(_01387_),
    .A(_00050_),
    .Y(_05242_));
 sg13g2_or2_1 _11699_ (.X(_05243_),
    .B(_05242_),
    .A(\u_toplayer.u_layer1.neuron_index[5] ));
 sg13g2_xnor2_1 _11700_ (.Y(_05244_),
    .A(\u_toplayer.u_layer1.neuron_index[4] ),
    .B(_01386_));
 sg13g2_nand2b_1 _11701_ (.Y(_05245_),
    .B(net2818),
    .A_N(_05244_));
 sg13g2_nor2_1 _11702_ (.A(net2874),
    .B(net2790),
    .Y(_05246_));
 sg13g2_nor2_1 _11703_ (.A(net815),
    .B(net2742),
    .Y(_05247_));
 sg13g2_a21oi_1 _11704_ (.A1(_01178_),
    .A2(net2742),
    .Y(_00709_),
    .B1(_05247_));
 sg13g2_nor2_1 _11705_ (.A(net824),
    .B(net2744),
    .Y(_05248_));
 sg13g2_a21oi_1 _11706_ (.A1(_01179_),
    .A2(net2743),
    .Y(_00710_),
    .B1(_05248_));
 sg13g2_nor2_1 _11707_ (.A(net820),
    .B(net2742),
    .Y(_05249_));
 sg13g2_a21oi_1 _11708_ (.A1(_01180_),
    .A2(net2742),
    .Y(_00711_),
    .B1(_05249_));
 sg13g2_nor2_1 _11709_ (.A(net817),
    .B(net2743),
    .Y(_05250_));
 sg13g2_a21oi_1 _11710_ (.A1(_01181_),
    .A2(net2743),
    .Y(_00712_),
    .B1(_05250_));
 sg13g2_nor2_1 _11711_ (.A(net876),
    .B(net2742),
    .Y(_05251_));
 sg13g2_a21oi_1 _11712_ (.A1(_01182_),
    .A2(net2742),
    .Y(_00713_),
    .B1(_05251_));
 sg13g2_nor2_1 _11713_ (.A(net906),
    .B(net2742),
    .Y(_05252_));
 sg13g2_a21oi_1 _11714_ (.A1(_01183_),
    .A2(net2742),
    .Y(_00714_),
    .B1(_05252_));
 sg13g2_nor2_1 _11715_ (.A(net915),
    .B(net2744),
    .Y(_05253_));
 sg13g2_a21oi_1 _11716_ (.A1(_01184_),
    .A2(net2744),
    .Y(_00715_),
    .B1(_05253_));
 sg13g2_mux2_1 _11717_ (.A0(net879),
    .A1(net3031),
    .S(net2744),
    .X(_00716_));
 sg13g2_xnor2_1 _11718_ (.Y(_05254_),
    .A(\u_toplayer.u_layer1.neuron_index[5] ),
    .B(_05242_));
 sg13g2_nand2_1 _11719_ (.Y(_05255_),
    .A(net2818),
    .B(_05244_));
 sg13g2_nor2_2 _11720_ (.A(_05254_),
    .B(net2777),
    .Y(_05256_));
 sg13g2_and2_1 _11721_ (.A(\u_toplayer.u_layer1.neuron_index[0] ),
    .B(_01384_),
    .X(_05257_));
 sg13g2_nor2b_1 _11722_ (.A(net3054),
    .B_N(net2911),
    .Y(_05258_));
 sg13g2_nand2_2 _11723_ (.Y(_05259_),
    .A(net2741),
    .B(_05258_));
 sg13g2_nand2_1 _11724_ (.Y(_05260_),
    .A(net668),
    .B(_05259_));
 sg13g2_xnor2_1 _11725_ (.Y(_05261_),
    .A(net3054),
    .B(net2980));
 sg13g2_nor2b_2 _11726_ (.A(_05254_),
    .B_N(_05261_),
    .Y(_05262_));
 sg13g2_nand2_1 _11727_ (.Y(_05263_),
    .A(\u_toplayer.u_layer1.sum[0] ),
    .B(net2912));
 sg13g2_nand3_1 _11728_ (.B(net2911),
    .C(net2851),
    .A(net3046),
    .Y(_05264_));
 sg13g2_o21ai_1 _11729_ (.B1(_05260_),
    .Y(_00717_),
    .A1(net2779),
    .A2(_05264_));
 sg13g2_nand2_1 _11730_ (.Y(_05265_),
    .A(net182),
    .B(_05259_));
 sg13g2_nand2_1 _11731_ (.Y(_05266_),
    .A(\u_toplayer.u_layer1.sum[1] ),
    .B(net2913));
 sg13g2_nand3_1 _11732_ (.B(net2913),
    .C(net2851),
    .A(net3044),
    .Y(_05267_));
 sg13g2_o21ai_1 _11733_ (.B1(_05265_),
    .Y(_00718_),
    .A1(net2778),
    .A2(_05267_));
 sg13g2_nand2_1 _11734_ (.Y(_05268_),
    .A(net262),
    .B(_05259_));
 sg13g2_nand2_1 _11735_ (.Y(_05269_),
    .A(net3043),
    .B(net2912));
 sg13g2_nand3_1 _11736_ (.B(net2911),
    .C(net2851),
    .A(\u_toplayer.u_layer1.sum[2] ),
    .Y(_05270_));
 sg13g2_o21ai_1 _11737_ (.B1(_05268_),
    .Y(_00719_),
    .A1(net2779),
    .A2(_05270_));
 sg13g2_nand2_1 _11738_ (.Y(_05271_),
    .A(net220),
    .B(_05259_));
 sg13g2_nand2_1 _11739_ (.Y(_05272_),
    .A(net3040),
    .B(net2912));
 sg13g2_nand3_1 _11740_ (.B(net2911),
    .C(net2851),
    .A(net3040),
    .Y(_05273_));
 sg13g2_o21ai_1 _11741_ (.B1(_05271_),
    .Y(_00720_),
    .A1(net2778),
    .A2(_05273_));
 sg13g2_nand2_1 _11742_ (.Y(_05274_),
    .A(net466),
    .B(_05259_));
 sg13g2_nand2_1 _11743_ (.Y(_05275_),
    .A(net3039),
    .B(net2913));
 sg13g2_nand3_1 _11744_ (.B(net2911),
    .C(net2851),
    .A(net3038),
    .Y(_05276_));
 sg13g2_o21ai_1 _11745_ (.B1(_05274_),
    .Y(_00721_),
    .A1(net2778),
    .A2(_05276_));
 sg13g2_nand2_1 _11746_ (.Y(_05277_),
    .A(net286),
    .B(_05259_));
 sg13g2_nand2_1 _11747_ (.Y(_05278_),
    .A(\u_toplayer.u_layer1.sum[5] ),
    .B(net2912));
 sg13g2_nand3_1 _11748_ (.B(net2911),
    .C(net2851),
    .A(\u_toplayer.u_layer1.sum[5] ),
    .Y(_05279_));
 sg13g2_o21ai_1 _11749_ (.B1(_05277_),
    .Y(_00722_),
    .A1(net2778),
    .A2(_05279_));
 sg13g2_nand2_1 _11750_ (.Y(_05280_),
    .A(net289),
    .B(_05259_));
 sg13g2_nand2_1 _11751_ (.Y(_05281_),
    .A(net3034),
    .B(net2912));
 sg13g2_nand3_1 _11752_ (.B(net2911),
    .C(net2850),
    .A(net3034),
    .Y(_05282_));
 sg13g2_o21ai_1 _11753_ (.B1(_05280_),
    .Y(_00723_),
    .A1(net2776),
    .A2(_05282_));
 sg13g2_nand2_1 _11754_ (.Y(_05283_),
    .A(net341),
    .B(_05259_));
 sg13g2_nand2_1 _11755_ (.Y(_05284_),
    .A(net3033),
    .B(net2912));
 sg13g2_nand3_1 _11756_ (.B(net2911),
    .C(net2850),
    .A(net3031),
    .Y(_05285_));
 sg13g2_o21ai_1 _11757_ (.B1(_05283_),
    .Y(_00724_),
    .A1(net2776),
    .A2(_05285_));
 sg13g2_nor2b_2 _11758_ (.A(\u_toplayer.u_layer1.neuron_index[0] ),
    .B_N(\u_toplayer.u_layer1.neuron_index[1] ),
    .Y(_05286_));
 sg13g2_nor2b_1 _11759_ (.A(net3056),
    .B_N(_05286_),
    .Y(_05287_));
 sg13g2_nor2b_1 _11760_ (.A(net3054),
    .B_N(net2910),
    .Y(_05288_));
 sg13g2_nand2_2 _11761_ (.Y(_05289_),
    .A(net2741),
    .B(_05288_));
 sg13g2_nand2_1 _11762_ (.Y(_05290_),
    .A(net690),
    .B(_05289_));
 sg13g2_nand4_1 _11763_ (.B(net2868),
    .C(net2846),
    .A(net3047),
    .Y(_05291_),
    .D(net2908));
 sg13g2_o21ai_1 _11764_ (.B1(_05290_),
    .Y(_00725_),
    .A1(net2773),
    .A2(_05291_));
 sg13g2_nand2_1 _11765_ (.Y(_05292_),
    .A(net806),
    .B(_05289_));
 sg13g2_nand3_1 _11766_ (.B(net2873),
    .C(net2910),
    .A(net3045),
    .Y(_05293_));
 sg13g2_nand4_1 _11767_ (.B(net2869),
    .C(net2848),
    .A(net3044),
    .Y(_05294_),
    .D(net2908));
 sg13g2_o21ai_1 _11768_ (.B1(_05292_),
    .Y(_00726_),
    .A1(net2775),
    .A2(_05294_));
 sg13g2_nand2_1 _11769_ (.Y(_05295_),
    .A(net467),
    .B(_05289_));
 sg13g2_nand3_1 _11770_ (.B(net2873),
    .C(net2910),
    .A(net3043),
    .Y(_05296_));
 sg13g2_nand4_1 _11771_ (.B(net2868),
    .C(net2845),
    .A(net3042),
    .Y(_05297_),
    .D(net2908));
 sg13g2_o21ai_1 _11772_ (.B1(_05295_),
    .Y(_00727_),
    .A1(net2772),
    .A2(_05297_));
 sg13g2_nand2_1 _11773_ (.Y(_05298_),
    .A(net544),
    .B(_05289_));
 sg13g2_nand3_1 _11774_ (.B(net2872),
    .C(net2909),
    .A(net3040),
    .Y(_05299_));
 sg13g2_nand4_1 _11775_ (.B(net2869),
    .C(net2848),
    .A(net3041),
    .Y(_05300_),
    .D(net2908));
 sg13g2_o21ai_1 _11776_ (.B1(_05298_),
    .Y(_00728_),
    .A1(net2775),
    .A2(_05300_));
 sg13g2_nand2_1 _11777_ (.Y(_05301_),
    .A(net367),
    .B(_05289_));
 sg13g2_nand4_1 _11778_ (.B(net2868),
    .C(net2848),
    .A(net3038),
    .Y(_05302_),
    .D(net2908));
 sg13g2_o21ai_1 _11779_ (.B1(_05301_),
    .Y(_00729_),
    .A1(net2775),
    .A2(_05302_));
 sg13g2_nand2_1 _11780_ (.Y(_05303_),
    .A(net564),
    .B(_05289_));
 sg13g2_nand3_1 _11781_ (.B(net2873),
    .C(net2909),
    .A(net3037),
    .Y(_05304_));
 sg13g2_nand4_1 _11782_ (.B(net2869),
    .C(net2848),
    .A(net3036),
    .Y(_05305_),
    .D(net2908));
 sg13g2_o21ai_1 _11783_ (.B1(_05303_),
    .Y(_00730_),
    .A1(net2775),
    .A2(_05305_));
 sg13g2_nand2_1 _11784_ (.Y(_05306_),
    .A(net562),
    .B(_05289_));
 sg13g2_nand4_1 _11785_ (.B(net2868),
    .C(net2845),
    .A(net3035),
    .Y(_05307_),
    .D(net2908));
 sg13g2_o21ai_1 _11786_ (.B1(_05306_),
    .Y(_00731_),
    .A1(net2776),
    .A2(_05307_));
 sg13g2_nand2_1 _11787_ (.Y(_05308_),
    .A(net692),
    .B(_05289_));
 sg13g2_nand3_1 _11788_ (.B(net2873),
    .C(net2909),
    .A(net3033),
    .Y(_05309_));
 sg13g2_nand4_1 _11789_ (.B(net2868),
    .C(net2845),
    .A(net3031),
    .Y(_05310_),
    .D(net2908));
 sg13g2_o21ai_1 _11790_ (.B1(_05308_),
    .Y(_00732_),
    .A1(net2772),
    .A2(_05310_));
 sg13g2_nor2_2 _11791_ (.A(net3056),
    .B(_05234_),
    .Y(_05311_));
 sg13g2_nor3_2 _11792_ (.A(net3056),
    .B(net3054),
    .C(_05234_),
    .Y(_05312_));
 sg13g2_nand2_2 _11793_ (.Y(_05313_),
    .A(_05256_),
    .B(_05312_));
 sg13g2_nand2_1 _11794_ (.Y(_05314_),
    .A(net378),
    .B(_05313_));
 sg13g2_nand2_1 _11795_ (.Y(_05315_),
    .A(net3046),
    .B(net2906));
 sg13g2_nand3_1 _11796_ (.B(net2846),
    .C(net2907),
    .A(net3047),
    .Y(_05316_));
 sg13g2_o21ai_1 _11797_ (.B1(_05314_),
    .Y(_00733_),
    .A1(net2773),
    .A2(_05316_));
 sg13g2_nand2_1 _11798_ (.Y(_05317_),
    .A(net392),
    .B(_05313_));
 sg13g2_nand2_1 _11799_ (.Y(_05318_),
    .A(net3045),
    .B(_05311_));
 sg13g2_nand3_1 _11800_ (.B(net2850),
    .C(net2907),
    .A(net3044),
    .Y(_05319_));
 sg13g2_o21ai_1 _11801_ (.B1(_05317_),
    .Y(_00734_),
    .A1(net2776),
    .A2(_05319_));
 sg13g2_nand2_1 _11802_ (.Y(_05320_),
    .A(net575),
    .B(_05313_));
 sg13g2_nand2_1 _11803_ (.Y(_05321_),
    .A(net3043),
    .B(net2906));
 sg13g2_nand3_1 _11804_ (.B(net2845),
    .C(net2907),
    .A(net3042),
    .Y(_05322_));
 sg13g2_o21ai_1 _11805_ (.B1(_05320_),
    .Y(_00735_),
    .A1(net2772),
    .A2(_05322_));
 sg13g2_nand2_1 _11806_ (.Y(_05323_),
    .A(net186),
    .B(_05313_));
 sg13g2_nand2_1 _11807_ (.Y(_05324_),
    .A(net3040),
    .B(net2906));
 sg13g2_nand3_1 _11808_ (.B(net2848),
    .C(net2907),
    .A(net3041),
    .Y(_05325_));
 sg13g2_o21ai_1 _11809_ (.B1(_05323_),
    .Y(_00736_),
    .A1(net2775),
    .A2(_05325_));
 sg13g2_nand2_1 _11810_ (.Y(_05326_),
    .A(net296),
    .B(_05313_));
 sg13g2_nand2_1 _11811_ (.Y(_05327_),
    .A(\u_toplayer.u_layer1.sum[4] ),
    .B(net2906));
 sg13g2_nand3_1 _11812_ (.B(net2848),
    .C(net2907),
    .A(net3038),
    .Y(_05328_));
 sg13g2_o21ai_1 _11813_ (.B1(_05326_),
    .Y(_00737_),
    .A1(net2775),
    .A2(_05328_));
 sg13g2_nand2_1 _11814_ (.Y(_05329_),
    .A(net539),
    .B(_05313_));
 sg13g2_nand2_1 _11815_ (.Y(_05330_),
    .A(net3037),
    .B(net2906));
 sg13g2_nand3_1 _11816_ (.B(net2848),
    .C(net2907),
    .A(net3036),
    .Y(_05331_));
 sg13g2_o21ai_1 _11817_ (.B1(_05329_),
    .Y(_00738_),
    .A1(net2775),
    .A2(_05331_));
 sg13g2_nand2_1 _11818_ (.Y(_05332_),
    .A(net291),
    .B(_05313_));
 sg13g2_nand2_1 _11819_ (.Y(_05333_),
    .A(net3034),
    .B(net2906));
 sg13g2_nand3_1 _11820_ (.B(net2845),
    .C(net2907),
    .A(net3035),
    .Y(_05334_));
 sg13g2_o21ai_1 _11821_ (.B1(_05332_),
    .Y(_00739_),
    .A1(net2776),
    .A2(_05334_));
 sg13g2_nand2_1 _11822_ (.Y(_05335_),
    .A(net607),
    .B(_05313_));
 sg13g2_nand2_1 _11823_ (.Y(_05336_),
    .A(net3033),
    .B(_05311_));
 sg13g2_nand3_1 _11824_ (.B(net2845),
    .C(net2907),
    .A(net3031),
    .Y(_05337_));
 sg13g2_o21ai_1 _11825_ (.B1(_05335_),
    .Y(_00740_),
    .A1(net2773),
    .A2(_05337_));
 sg13g2_nor2b_1 _11826_ (.A(\u_toplayer.u_layer1.neuron_index[1] ),
    .B_N(net3055),
    .Y(_05338_));
 sg13g2_nor2b_1 _11827_ (.A(net3057),
    .B_N(_05338_),
    .Y(_05339_));
 sg13g2_nand3b_1 _11828_ (.B(net2741),
    .C(net2903),
    .Y(_05340_),
    .A_N(net3053));
 sg13g2_nand2_1 _11829_ (.Y(_05341_),
    .A(net280),
    .B(_05340_));
 sg13g2_nand2_1 _11830_ (.Y(_05342_),
    .A(\u_toplayer.u_layer1.sum[0] ),
    .B(net2905));
 sg13g2_nand3_1 _11831_ (.B(net2843),
    .C(net2903),
    .A(net3047),
    .Y(_05343_));
 sg13g2_o21ai_1 _11832_ (.B1(_05341_),
    .Y(_00741_),
    .A1(net2769),
    .A2(_05343_));
 sg13g2_nand2_1 _11833_ (.Y(_05344_),
    .A(net499),
    .B(_05340_));
 sg13g2_nand2_1 _11834_ (.Y(_05345_),
    .A(net3045),
    .B(net2904));
 sg13g2_nand3_1 _11835_ (.B(net2843),
    .C(net2903),
    .A(net3044),
    .Y(_05346_));
 sg13g2_o21ai_1 _11836_ (.B1(_05344_),
    .Y(_00742_),
    .A1(net2769),
    .A2(_05346_));
 sg13g2_nand2_1 _11837_ (.Y(_05347_),
    .A(net450),
    .B(_05340_));
 sg13g2_nand2_1 _11838_ (.Y(_05348_),
    .A(net3043),
    .B(net2904));
 sg13g2_nand3_1 _11839_ (.B(net2847),
    .C(net2903),
    .A(net3042),
    .Y(_05349_));
 sg13g2_o21ai_1 _11840_ (.B1(_05347_),
    .Y(_00743_),
    .A1(net2771),
    .A2(_05349_));
 sg13g2_nand2_1 _11841_ (.Y(_05350_),
    .A(net325),
    .B(_05340_));
 sg13g2_nand2_1 _11842_ (.Y(_05351_),
    .A(net3040),
    .B(net2904));
 sg13g2_nand3_1 _11843_ (.B(net2847),
    .C(net2903),
    .A(net3041),
    .Y(_05352_));
 sg13g2_o21ai_1 _11844_ (.B1(_05350_),
    .Y(_00744_),
    .A1(net2771),
    .A2(_05352_));
 sg13g2_nand2_1 _11845_ (.Y(_05353_),
    .A(net342),
    .B(_05340_));
 sg13g2_nand2_1 _11846_ (.Y(_05354_),
    .A(net3039),
    .B(net2904));
 sg13g2_nand3_1 _11847_ (.B(net2849),
    .C(net2905),
    .A(net3038),
    .Y(_05355_));
 sg13g2_o21ai_1 _11848_ (.B1(_05353_),
    .Y(_00745_),
    .A1(net2774),
    .A2(_05355_));
 sg13g2_nand2_1 _11849_ (.Y(_05356_),
    .A(net794),
    .B(_05340_));
 sg13g2_nand2_1 _11850_ (.Y(_05357_),
    .A(net3037),
    .B(net2904));
 sg13g2_nand3_1 _11851_ (.B(net2849),
    .C(net2905),
    .A(net3036),
    .Y(_05358_));
 sg13g2_o21ai_1 _11852_ (.B1(_05356_),
    .Y(_00746_),
    .A1(net2774),
    .A2(_05358_));
 sg13g2_nand2_1 _11853_ (.Y(_05359_),
    .A(net891),
    .B(_05340_));
 sg13g2_nand2_1 _11854_ (.Y(_05360_),
    .A(\u_toplayer.u_layer1.sum[6] ),
    .B(net2904));
 sg13g2_nand3_1 _11855_ (.B(net2843),
    .C(net2903),
    .A(net3035),
    .Y(_05361_));
 sg13g2_o21ai_1 _11856_ (.B1(_05359_),
    .Y(_00747_),
    .A1(net2769),
    .A2(_05361_));
 sg13g2_nand2_1 _11857_ (.Y(_05362_),
    .A(net543),
    .B(_05340_));
 sg13g2_nand2_1 _11858_ (.Y(_05363_),
    .A(net3033),
    .B(net2905));
 sg13g2_nand3_1 _11859_ (.B(net2843),
    .C(net2903),
    .A(net3031),
    .Y(_05364_));
 sg13g2_o21ai_1 _11860_ (.B1(_05362_),
    .Y(_00748_),
    .A1(net2769),
    .A2(_05364_));
 sg13g2_and2_1 _11861_ (.A(net3057),
    .B(_05338_),
    .X(_05365_));
 sg13g2_nor2b_1 _11862_ (.A(net3053),
    .B_N(net2900),
    .Y(_05366_));
 sg13g2_nand2_2 _11863_ (.Y(_05367_),
    .A(net2741),
    .B(_05366_));
 sg13g2_nand2_1 _11864_ (.Y(_05368_),
    .A(net200),
    .B(_05367_));
 sg13g2_nand2_1 _11865_ (.Y(_05369_),
    .A(net3047),
    .B(net2901));
 sg13g2_nand3_1 _11866_ (.B(net2843),
    .C(net2900),
    .A(net3047),
    .Y(_05370_));
 sg13g2_o21ai_1 _11867_ (.B1(_05368_),
    .Y(_00749_),
    .A1(net2769),
    .A2(_05370_));
 sg13g2_nand2_1 _11868_ (.Y(_05371_),
    .A(net363),
    .B(_05367_));
 sg13g2_nand2_1 _11869_ (.Y(_05372_),
    .A(net3045),
    .B(net2901));
 sg13g2_nand3_1 _11870_ (.B(net2843),
    .C(net2900),
    .A(net3044),
    .Y(_05373_));
 sg13g2_o21ai_1 _11871_ (.B1(_05371_),
    .Y(_00750_),
    .A1(net2769),
    .A2(_05373_));
 sg13g2_nand2_1 _11872_ (.Y(_05374_),
    .A(net602),
    .B(_05367_));
 sg13g2_nand2_1 _11873_ (.Y(_05375_),
    .A(\u_toplayer.u_layer1.sum[2] ),
    .B(net2901));
 sg13g2_nand3_1 _11874_ (.B(net2844),
    .C(net2900),
    .A(net3042),
    .Y(_05376_));
 sg13g2_o21ai_1 _11875_ (.B1(_05374_),
    .Y(_00751_),
    .A1(net2771),
    .A2(_05376_));
 sg13g2_nand2_1 _11876_ (.Y(_05377_),
    .A(net719),
    .B(_05367_));
 sg13g2_nand2_1 _11877_ (.Y(_05378_),
    .A(\u_toplayer.u_layer1.sum[3] ),
    .B(net2901));
 sg13g2_nand3_1 _11878_ (.B(net2844),
    .C(net2900),
    .A(net3041),
    .Y(_05379_));
 sg13g2_o21ai_1 _11879_ (.B1(_05377_),
    .Y(_00752_),
    .A1(net2771),
    .A2(_05379_));
 sg13g2_nand2_1 _11880_ (.Y(_05380_),
    .A(net809),
    .B(_05367_));
 sg13g2_nand2_1 _11881_ (.Y(_05381_),
    .A(\u_toplayer.u_layer1.sum[4] ),
    .B(net2902));
 sg13g2_nand3_1 _11882_ (.B(net2849),
    .C(net2902),
    .A(net3038),
    .Y(_05382_));
 sg13g2_o21ai_1 _11883_ (.B1(_05380_),
    .Y(_00753_),
    .A1(net2774),
    .A2(_05382_));
 sg13g2_nand2_1 _11884_ (.Y(_05383_),
    .A(net542),
    .B(_05367_));
 sg13g2_nand2_1 _11885_ (.Y(_05384_),
    .A(net3037),
    .B(net2902));
 sg13g2_nand3_1 _11886_ (.B(net2849),
    .C(net2900),
    .A(net3036),
    .Y(_05385_));
 sg13g2_o21ai_1 _11887_ (.B1(_05383_),
    .Y(_00754_),
    .A1(net2774),
    .A2(_05385_));
 sg13g2_nand2_1 _11888_ (.Y(_05386_),
    .A(net782),
    .B(_05367_));
 sg13g2_nand2_1 _11889_ (.Y(_05387_),
    .A(\u_toplayer.u_layer1.sum[6] ),
    .B(net2901));
 sg13g2_nand3_1 _11890_ (.B(net2843),
    .C(net2900),
    .A(net3035),
    .Y(_05388_));
 sg13g2_o21ai_1 _11891_ (.B1(_05386_),
    .Y(_00755_),
    .A1(net2769),
    .A2(_05388_));
 sg13g2_nand2_1 _11892_ (.Y(_05389_),
    .A(net169),
    .B(_05367_));
 sg13g2_nand2_1 _11893_ (.Y(_05390_),
    .A(net3033),
    .B(net2901));
 sg13g2_nand3_1 _11894_ (.B(net2843),
    .C(net2900),
    .A(net3031),
    .Y(_05391_));
 sg13g2_o21ai_1 _11895_ (.B1(_05389_),
    .Y(_00756_),
    .A1(net2769),
    .A2(_05391_));
 sg13g2_and2_1 _11896_ (.A(net3056),
    .B(_05286_),
    .X(_05392_));
 sg13g2_nor2b_1 _11897_ (.A(net3054),
    .B_N(net2899),
    .Y(_05393_));
 sg13g2_nand2_2 _11898_ (.Y(_05394_),
    .A(net2741),
    .B(_05393_));
 sg13g2_nand2_1 _11899_ (.Y(_05395_),
    .A(net610),
    .B(_05394_));
 sg13g2_nand4_1 _11900_ (.B(net2868),
    .C(net2844),
    .A(net3047),
    .Y(_05396_),
    .D(net2898));
 sg13g2_o21ai_1 _11901_ (.B1(_05395_),
    .Y(_00757_),
    .A1(net2770),
    .A2(_05396_));
 sg13g2_nand2_1 _11902_ (.Y(_05397_),
    .A(net264),
    .B(_05394_));
 sg13g2_nand3_1 _11903_ (.B(net3045),
    .C(_05286_),
    .A(net3056),
    .Y(_05398_));
 sg13g2_nand4_1 _11904_ (.B(net2871),
    .C(net2846),
    .A(net3044),
    .Y(_05399_),
    .D(net2898));
 sg13g2_o21ai_1 _11905_ (.B1(_05397_),
    .Y(_00758_),
    .A1(net2772),
    .A2(_05399_));
 sg13g2_nand2_1 _11906_ (.Y(_05400_),
    .A(net534),
    .B(_05394_));
 sg13g2_nand3_1 _11907_ (.B(net3043),
    .C(_05286_),
    .A(net3056),
    .Y(_05401_));
 sg13g2_nand4_1 _11908_ (.B(net2868),
    .C(net2845),
    .A(net3042),
    .Y(_05402_),
    .D(net2898));
 sg13g2_o21ai_1 _11909_ (.B1(_05400_),
    .Y(_00759_),
    .A1(net2770),
    .A2(_05402_));
 sg13g2_nand2_1 _11910_ (.Y(_05403_),
    .A(net274),
    .B(_05394_));
 sg13g2_nand3_1 _11911_ (.B(net3041),
    .C(_05286_),
    .A(net3055),
    .Y(_05404_));
 sg13g2_nand4_1 _11912_ (.B(net2868),
    .C(net2845),
    .A(net3041),
    .Y(_05405_),
    .D(net2898));
 sg13g2_o21ai_1 _11913_ (.B1(_05403_),
    .Y(_00760_),
    .A1(net2770),
    .A2(_05405_));
 sg13g2_nand2_1 _11914_ (.Y(_05406_),
    .A(net320),
    .B(_05394_));
 sg13g2_nand3_1 _11915_ (.B(net3038),
    .C(_05286_),
    .A(net3055),
    .Y(_05407_));
 sg13g2_nand4_1 _11916_ (.B(net2870),
    .C(net2849),
    .A(net3039),
    .Y(_05408_),
    .D(net2899));
 sg13g2_o21ai_1 _11917_ (.B1(_05406_),
    .Y(_00761_),
    .A1(net2774),
    .A2(_05408_));
 sg13g2_nand2_1 _11918_ (.Y(_05409_),
    .A(net723),
    .B(_05394_));
 sg13g2_nand3_1 _11919_ (.B(net3036),
    .C(_05286_),
    .A(net3055),
    .Y(_05410_));
 sg13g2_nand4_1 _11920_ (.B(net2869),
    .C(net2848),
    .A(net3036),
    .Y(_05411_),
    .D(net2898));
 sg13g2_o21ai_1 _11921_ (.B1(_05409_),
    .Y(_00762_),
    .A1(net2775),
    .A2(_05411_));
 sg13g2_nand2_1 _11922_ (.Y(_05412_),
    .A(net732),
    .B(_05394_));
 sg13g2_nand4_1 _11923_ (.B(net2871),
    .C(net2846),
    .A(net3035),
    .Y(_05413_),
    .D(net2898));
 sg13g2_o21ai_1 _11924_ (.B1(_05412_),
    .Y(_00763_),
    .A1(net2772),
    .A2(_05413_));
 sg13g2_nand2_1 _11925_ (.Y(_05414_),
    .A(net408),
    .B(_05394_));
 sg13g2_nand3_1 _11926_ (.B(net3032),
    .C(_05286_),
    .A(net3056),
    .Y(_05415_));
 sg13g2_nand4_1 _11927_ (.B(net2871),
    .C(net2846),
    .A(net3031),
    .Y(_05416_),
    .D(net2898));
 sg13g2_o21ai_1 _11928_ (.B1(_05414_),
    .Y(_00764_),
    .A1(net2772),
    .A2(_05416_));
 sg13g2_nor2b_1 _11929_ (.A(net3054),
    .B_N(net2945),
    .Y(_05417_));
 sg13g2_nand2_2 _11930_ (.Y(_05418_),
    .A(net2741),
    .B(_05417_));
 sg13g2_nand2_1 _11931_ (.Y(_05419_),
    .A(net178),
    .B(_05418_));
 sg13g2_nand2_1 _11932_ (.Y(_05420_),
    .A(net3046),
    .B(net2946));
 sg13g2_nand3_1 _11933_ (.B(net2945),
    .C(net2844),
    .A(net3047),
    .Y(_05421_));
 sg13g2_o21ai_1 _11934_ (.B1(_05419_),
    .Y(_00765_),
    .A1(net2770),
    .A2(_05421_));
 sg13g2_nand2_1 _11935_ (.Y(_05422_),
    .A(net530),
    .B(_05418_));
 sg13g2_nand2_1 _11936_ (.Y(_05423_),
    .A(\u_toplayer.u_layer1.sum[1] ),
    .B(net2946));
 sg13g2_nand3_1 _11937_ (.B(net2945),
    .C(net2846),
    .A(net3044),
    .Y(_05424_));
 sg13g2_o21ai_1 _11938_ (.B1(_05422_),
    .Y(_00766_),
    .A1(net2772),
    .A2(_05424_));
 sg13g2_nand2_1 _11939_ (.Y(_05425_),
    .A(net415),
    .B(_05418_));
 sg13g2_nand2_1 _11940_ (.Y(_05426_),
    .A(net3042),
    .B(net2946));
 sg13g2_nand3_1 _11941_ (.B(net2945),
    .C(net2844),
    .A(net3042),
    .Y(_05427_));
 sg13g2_o21ai_1 _11942_ (.B1(_05425_),
    .Y(_00767_),
    .A1(net2770),
    .A2(_05427_));
 sg13g2_nand2_1 _11943_ (.Y(_05428_),
    .A(net462),
    .B(_05418_));
 sg13g2_nand2_1 _11944_ (.Y(_05429_),
    .A(net3040),
    .B(net2946));
 sg13g2_nand3_1 _11945_ (.B(net2945),
    .C(net2844),
    .A(net3041),
    .Y(_05430_));
 sg13g2_o21ai_1 _11946_ (.B1(_05428_),
    .Y(_00768_),
    .A1(net2770),
    .A2(_05430_));
 sg13g2_nand2_1 _11947_ (.Y(_05431_),
    .A(net608),
    .B(_05418_));
 sg13g2_nand2_1 _11948_ (.Y(_05432_),
    .A(net3038),
    .B(net2946));
 sg13g2_nand3_1 _11949_ (.B(net2947),
    .C(net2849),
    .A(net3038),
    .Y(_05433_));
 sg13g2_o21ai_1 _11950_ (.B1(_05431_),
    .Y(_00769_),
    .A1(net2774),
    .A2(_05433_));
 sg13g2_nand2_1 _11951_ (.Y(_05434_),
    .A(net482),
    .B(_05418_));
 sg13g2_nand2_1 _11952_ (.Y(_05435_),
    .A(net3036),
    .B(net2946));
 sg13g2_nand3_1 _11953_ (.B(net2947),
    .C(net2849),
    .A(net3037),
    .Y(_05436_));
 sg13g2_o21ai_1 _11954_ (.B1(_05434_),
    .Y(_00770_),
    .A1(net2774),
    .A2(_05436_));
 sg13g2_nand2_1 _11955_ (.Y(_05437_),
    .A(net175),
    .B(_05418_));
 sg13g2_nand2_1 _11956_ (.Y(_05438_),
    .A(net3034),
    .B(net2946));
 sg13g2_nand3_1 _11957_ (.B(net2945),
    .C(net2844),
    .A(net3035),
    .Y(_05439_));
 sg13g2_o21ai_1 _11958_ (.B1(_05437_),
    .Y(_00771_),
    .A1(net2770),
    .A2(_05439_));
 sg13g2_nand2_1 _11959_ (.Y(_05440_),
    .A(net531),
    .B(_05418_));
 sg13g2_nand2_1 _11960_ (.Y(_05441_),
    .A(net3032),
    .B(net2946));
 sg13g2_nand3_1 _11961_ (.B(net2945),
    .C(net2846),
    .A(net3031),
    .Y(_05442_));
 sg13g2_o21ai_1 _11962_ (.B1(_05440_),
    .Y(_00772_),
    .A1(net2772),
    .A2(_05442_));
 sg13g2_and2_2 _11963_ (.A(net3054),
    .B(net2741),
    .X(_05443_));
 sg13g2_nand2_2 _11964_ (.Y(_05444_),
    .A(net2982),
    .B(_05443_));
 sg13g2_nand2_1 _11965_ (.Y(_05445_),
    .A(net639),
    .B(_05444_));
 sg13g2_nand3_1 _11966_ (.B(net2980),
    .C(net2870),
    .A(net3046),
    .Y(_05446_));
 sg13g2_nand4_1 _11967_ (.B(net2982),
    .C(net2872),
    .A(net3046),
    .Y(_05447_),
    .D(net2852));
 sg13g2_o21ai_1 _11968_ (.B1(_05445_),
    .Y(_00773_),
    .A1(net2780),
    .A2(_05447_));
 sg13g2_nand2_1 _11969_ (.Y(_05448_),
    .A(net432),
    .B(_05444_));
 sg13g2_nand3_1 _11970_ (.B(net2981),
    .C(net2870),
    .A(net3044),
    .Y(_05449_));
 sg13g2_nand4_1 _11971_ (.B(net2983),
    .C(net2872),
    .A(net3045),
    .Y(_05450_),
    .D(net2852));
 sg13g2_o21ai_1 _11972_ (.B1(_05448_),
    .Y(_00774_),
    .A1(net2780),
    .A2(_05450_));
 sg13g2_nand2_1 _11973_ (.Y(_05451_),
    .A(net328),
    .B(_05444_));
 sg13g2_nand3_1 _11974_ (.B(net2981),
    .C(net2870),
    .A(net3042),
    .Y(_05452_));
 sg13g2_nand4_1 _11975_ (.B(net2982),
    .C(net2872),
    .A(net3043),
    .Y(_05453_),
    .D(net2852));
 sg13g2_o21ai_1 _11976_ (.B1(_05451_),
    .Y(_00775_),
    .A1(net2779),
    .A2(_05453_));
 sg13g2_nand2_1 _11977_ (.Y(_05454_),
    .A(net730),
    .B(_05444_));
 sg13g2_nand3_1 _11978_ (.B(net2981),
    .C(net2869),
    .A(net3041),
    .Y(_05455_));
 sg13g2_nand4_1 _11979_ (.B(net2982),
    .C(net2872),
    .A(net3040),
    .Y(_05456_),
    .D(net2852));
 sg13g2_o21ai_1 _11980_ (.B1(_05454_),
    .Y(_00776_),
    .A1(net2779),
    .A2(_05456_));
 sg13g2_nand2_1 _11981_ (.Y(_05457_),
    .A(net717),
    .B(_05444_));
 sg13g2_nand3_1 _11982_ (.B(net2980),
    .C(net2870),
    .A(net3039),
    .Y(_05458_));
 sg13g2_nand4_1 _11983_ (.B(net2983),
    .C(net2872),
    .A(net3039),
    .Y(_05459_),
    .D(net2852));
 sg13g2_o21ai_1 _11984_ (.B1(_05457_),
    .Y(_00777_),
    .A1(net2780),
    .A2(_05459_));
 sg13g2_nand2_1 _11985_ (.Y(_05460_),
    .A(net376),
    .B(_05444_));
 sg13g2_nand3_1 _11986_ (.B(net2980),
    .C(net2869),
    .A(net3036),
    .Y(_05461_));
 sg13g2_nand4_1 _11987_ (.B(net2982),
    .C(net2872),
    .A(net3037),
    .Y(_05462_),
    .D(net2852));
 sg13g2_o21ai_1 _11988_ (.B1(_05460_),
    .Y(_00778_),
    .A1(net2779),
    .A2(_05462_));
 sg13g2_nand2_1 _11989_ (.Y(_05463_),
    .A(net640),
    .B(_05444_));
 sg13g2_nand3_1 _11990_ (.B(net2980),
    .C(net2869),
    .A(net3035),
    .Y(_05464_));
 sg13g2_nand4_1 _11991_ (.B(net2982),
    .C(net2872),
    .A(net3034),
    .Y(_05465_),
    .D(net2851));
 sg13g2_o21ai_1 _11992_ (.B1(_05463_),
    .Y(_00779_),
    .A1(net2779),
    .A2(_05465_));
 sg13g2_nand2_1 _11993_ (.Y(_05466_),
    .A(net514),
    .B(_05444_));
 sg13g2_nand3_1 _11994_ (.B(net2980),
    .C(net2869),
    .A(net3032),
    .Y(_05467_));
 sg13g2_nand4_1 _11995_ (.B(net2982),
    .C(net2873),
    .A(net3033),
    .Y(_05468_),
    .D(net2851));
 sg13g2_o21ai_1 _11996_ (.B1(_05466_),
    .Y(_00780_),
    .A1(net2779),
    .A2(_05468_));
 sg13g2_nand2_2 _11997_ (.Y(_05469_),
    .A(net2912),
    .B(_05443_));
 sg13g2_nand2_1 _11998_ (.Y(_05470_),
    .A(net351),
    .B(_05469_));
 sg13g2_nand2b_1 _11999_ (.Y(_05471_),
    .B(net2741),
    .A_N(_05261_));
 sg13g2_nor2_2 _12000_ (.A(_05254_),
    .B(_05261_),
    .Y(_05472_));
 sg13g2_o21ai_1 _12001_ (.B1(_05470_),
    .Y(_00781_),
    .A1(_05263_),
    .A2(net2723));
 sg13g2_nand2_1 _12002_ (.Y(_05473_),
    .A(net451),
    .B(_05469_));
 sg13g2_o21ai_1 _12003_ (.B1(_05473_),
    .Y(_00782_),
    .A1(_05266_),
    .A2(net2724));
 sg13g2_nand2_1 _12004_ (.Y(_05474_),
    .A(net678),
    .B(_05469_));
 sg13g2_o21ai_1 _12005_ (.B1(_05474_),
    .Y(_00783_),
    .A1(_05269_),
    .A2(net2724));
 sg13g2_nand2_1 _12006_ (.Y(_05475_),
    .A(net701),
    .B(_05469_));
 sg13g2_o21ai_1 _12007_ (.B1(_05475_),
    .Y(_00784_),
    .A1(_05272_),
    .A2(net2724));
 sg13g2_nand2_1 _12008_ (.Y(_05476_),
    .A(net297),
    .B(_05469_));
 sg13g2_o21ai_1 _12009_ (.B1(_05476_),
    .Y(_00785_),
    .A1(_05275_),
    .A2(net2724));
 sg13g2_nand2_1 _12010_ (.Y(_05477_),
    .A(net711),
    .B(_05469_));
 sg13g2_o21ai_1 _12011_ (.B1(_05477_),
    .Y(_00786_),
    .A1(_05278_),
    .A2(net2723));
 sg13g2_nand2_1 _12012_ (.Y(_05478_),
    .A(net502),
    .B(_05469_));
 sg13g2_o21ai_1 _12013_ (.B1(_05478_),
    .Y(_00787_),
    .A1(_05281_),
    .A2(net2723));
 sg13g2_nand2_1 _12014_ (.Y(_05479_),
    .A(net571),
    .B(_05469_));
 sg13g2_o21ai_1 _12015_ (.B1(_05479_),
    .Y(_00788_),
    .A1(_05284_),
    .A2(net2724));
 sg13g2_nand2_2 _12016_ (.Y(_05480_),
    .A(net2909),
    .B(_05443_));
 sg13g2_nand2_1 _12017_ (.Y(_05481_),
    .A(net442),
    .B(_05480_));
 sg13g2_nand4_1 _12018_ (.B(net2874),
    .C(net2909),
    .A(net3046),
    .Y(_05482_),
    .D(_05472_));
 sg13g2_o21ai_1 _12019_ (.B1(_05481_),
    .Y(_00789_),
    .A1(net2778),
    .A2(_05482_));
 sg13g2_nand2_1 _12020_ (.Y(_05483_),
    .A(net558),
    .B(_05480_));
 sg13g2_o21ai_1 _12021_ (.B1(_05483_),
    .Y(_00790_),
    .A1(_05293_),
    .A2(net2725));
 sg13g2_nand2_1 _12022_ (.Y(_05484_),
    .A(net519),
    .B(_05480_));
 sg13g2_o21ai_1 _12023_ (.B1(_05484_),
    .Y(_00791_),
    .A1(_05296_),
    .A2(net2725));
 sg13g2_nand2_1 _12024_ (.Y(_05485_),
    .A(net729),
    .B(_05480_));
 sg13g2_o21ai_1 _12025_ (.B1(_05485_),
    .Y(_00792_),
    .A1(_05299_),
    .A2(net2726));
 sg13g2_nand2_1 _12026_ (.Y(_05486_),
    .A(net425),
    .B(_05480_));
 sg13g2_nand4_1 _12027_ (.B(net2874),
    .C(net2909),
    .A(net3039),
    .Y(_05487_),
    .D(_05472_));
 sg13g2_o21ai_1 _12028_ (.B1(_05486_),
    .Y(_00793_),
    .A1(net2778),
    .A2(_05487_));
 sg13g2_nand2_1 _12029_ (.Y(_05488_),
    .A(net242),
    .B(_05480_));
 sg13g2_o21ai_1 _12030_ (.B1(_05488_),
    .Y(_00794_),
    .A1(_05304_),
    .A2(net2725));
 sg13g2_nand2_1 _12031_ (.Y(_05489_),
    .A(net672),
    .B(_05480_));
 sg13g2_nand4_1 _12032_ (.B(net2874),
    .C(net2909),
    .A(net3034),
    .Y(_05490_),
    .D(_05472_));
 sg13g2_o21ai_1 _12033_ (.B1(_05489_),
    .Y(_00795_),
    .A1(net2778),
    .A2(_05490_));
 sg13g2_nand2_1 _12034_ (.Y(_05491_),
    .A(net573),
    .B(_05480_));
 sg13g2_o21ai_1 _12035_ (.B1(_05491_),
    .Y(_00796_),
    .A1(_05309_),
    .A2(net2726));
 sg13g2_nand2_2 _12036_ (.Y(_05492_),
    .A(net2906),
    .B(_05443_));
 sg13g2_nand2_1 _12037_ (.Y(_05493_),
    .A(net354),
    .B(_05492_));
 sg13g2_o21ai_1 _12038_ (.B1(_05493_),
    .Y(_00797_),
    .A1(_05315_),
    .A2(net2725));
 sg13g2_nand2_1 _12039_ (.Y(_05494_),
    .A(net199),
    .B(_05492_));
 sg13g2_o21ai_1 _12040_ (.B1(_05494_),
    .Y(_00798_),
    .A1(_05318_),
    .A2(net2725));
 sg13g2_nand2_1 _12041_ (.Y(_05495_),
    .A(net617),
    .B(_05492_));
 sg13g2_o21ai_1 _12042_ (.B1(_05495_),
    .Y(_00799_),
    .A1(_05321_),
    .A2(net2725));
 sg13g2_nand2_1 _12043_ (.Y(_05496_),
    .A(net460),
    .B(_05492_));
 sg13g2_o21ai_1 _12044_ (.B1(_05496_),
    .Y(_00800_),
    .A1(_05324_),
    .A2(net2726));
 sg13g2_nand2_1 _12045_ (.Y(_05497_),
    .A(net783),
    .B(_05492_));
 sg13g2_o21ai_1 _12046_ (.B1(_05497_),
    .Y(_00801_),
    .A1(_05327_),
    .A2(net2721));
 sg13g2_nand2_1 _12047_ (.Y(_05498_),
    .A(net222),
    .B(_05492_));
 sg13g2_o21ai_1 _12048_ (.B1(_05498_),
    .Y(_00802_),
    .A1(_05330_),
    .A2(net2725));
 sg13g2_nand2_1 _12049_ (.Y(_05499_),
    .A(net345),
    .B(_05492_));
 sg13g2_o21ai_1 _12050_ (.B1(_05499_),
    .Y(_00803_),
    .A1(_05333_),
    .A2(net2721));
 sg13g2_nand2_1 _12051_ (.Y(_05500_),
    .A(net699),
    .B(_05492_));
 sg13g2_o21ai_1 _12052_ (.B1(_05500_),
    .Y(_00804_),
    .A1(_05336_),
    .A2(net2725));
 sg13g2_nand2_2 _12053_ (.Y(_05501_),
    .A(net2904),
    .B(_05443_));
 sg13g2_nand2_1 _12054_ (.Y(_05502_),
    .A(net365),
    .B(_05501_));
 sg13g2_o21ai_1 _12055_ (.B1(_05502_),
    .Y(_00805_),
    .A1(_05342_),
    .A2(net2719));
 sg13g2_nand2_1 _12056_ (.Y(_05503_),
    .A(net418),
    .B(_05501_));
 sg13g2_o21ai_1 _12057_ (.B1(_05503_),
    .Y(_00806_),
    .A1(_05345_),
    .A2(net2722));
 sg13g2_nand2_1 _12058_ (.Y(_05504_),
    .A(net561),
    .B(_05501_));
 sg13g2_o21ai_1 _12059_ (.B1(_05504_),
    .Y(_00807_),
    .A1(_05348_),
    .A2(net2718));
 sg13g2_nand2_1 _12060_ (.Y(_05505_),
    .A(net720),
    .B(_05501_));
 sg13g2_o21ai_1 _12061_ (.B1(_05505_),
    .Y(_00808_),
    .A1(_05351_),
    .A2(net2722));
 sg13g2_nand2_1 _12062_ (.Y(_05506_),
    .A(net582),
    .B(_05501_));
 sg13g2_o21ai_1 _12063_ (.B1(_05506_),
    .Y(_00809_),
    .A1(_05354_),
    .A2(net2718));
 sg13g2_nand2_1 _12064_ (.Y(_05507_),
    .A(net374),
    .B(_05501_));
 sg13g2_o21ai_1 _12065_ (.B1(_05507_),
    .Y(_00810_),
    .A1(_05357_),
    .A2(net2718));
 sg13g2_nand2_1 _12066_ (.Y(_05508_),
    .A(net298),
    .B(_05501_));
 sg13g2_o21ai_1 _12067_ (.B1(_05508_),
    .Y(_00811_),
    .A1(_05360_),
    .A2(net2718));
 sg13g2_nand2_1 _12068_ (.Y(_05509_),
    .A(net311),
    .B(_05501_));
 sg13g2_o21ai_1 _12069_ (.B1(_05509_),
    .Y(_00812_),
    .A1(_05363_),
    .A2(net2718));
 sg13g2_nand2_2 _12070_ (.Y(_05510_),
    .A(net2901),
    .B(_05443_));
 sg13g2_nand2_1 _12071_ (.Y(_05511_),
    .A(net726),
    .B(_05510_));
 sg13g2_o21ai_1 _12072_ (.B1(_05511_),
    .Y(_00813_),
    .A1(_05369_),
    .A2(net2723));
 sg13g2_nand2_1 _12073_ (.Y(_05512_),
    .A(net885),
    .B(_05510_));
 sg13g2_o21ai_1 _12074_ (.B1(_05512_),
    .Y(_00814_),
    .A1(_05372_),
    .A2(net2722));
 sg13g2_nand2_1 _12075_ (.Y(_05513_),
    .A(net623),
    .B(_05510_));
 sg13g2_o21ai_1 _12076_ (.B1(_05513_),
    .Y(_00815_),
    .A1(_05375_),
    .A2(net2722));
 sg13g2_nand2_1 _12077_ (.Y(_05514_),
    .A(net688),
    .B(_05510_));
 sg13g2_o21ai_1 _12078_ (.B1(_05514_),
    .Y(_00816_),
    .A1(_05378_),
    .A2(net2722));
 sg13g2_nand2_1 _12079_ (.Y(_05515_),
    .A(net755),
    .B(_05510_));
 sg13g2_o21ai_1 _12080_ (.B1(_05515_),
    .Y(_00817_),
    .A1(_05381_),
    .A2(net2722));
 sg13g2_nand2_1 _12081_ (.Y(_05516_),
    .A(net379),
    .B(_05510_));
 sg13g2_o21ai_1 _12082_ (.B1(_05516_),
    .Y(_00818_),
    .A1(_05384_),
    .A2(net2722));
 sg13g2_nand2_1 _12083_ (.Y(_05517_),
    .A(net774),
    .B(_05510_));
 sg13g2_o21ai_1 _12084_ (.B1(_05517_),
    .Y(_00819_),
    .A1(_05387_),
    .A2(net2723));
 sg13g2_nand2_1 _12085_ (.Y(_05518_),
    .A(net278),
    .B(_05510_));
 sg13g2_o21ai_1 _12086_ (.B1(_05518_),
    .Y(_00820_),
    .A1(_05390_),
    .A2(net2722));
 sg13g2_nand2_2 _12087_ (.Y(_05519_),
    .A(net2899),
    .B(_05443_));
 sg13g2_nand2_1 _12088_ (.Y(_05520_),
    .A(net540),
    .B(_05519_));
 sg13g2_nand4_1 _12089_ (.B(net2874),
    .C(net2899),
    .A(net3046),
    .Y(_05521_),
    .D(_05472_));
 sg13g2_o21ai_1 _12090_ (.B1(_05520_),
    .Y(_00821_),
    .A1(net2778),
    .A2(_05521_));
 sg13g2_nand2_1 _12091_ (.Y(_05522_),
    .A(net416),
    .B(_05519_));
 sg13g2_o21ai_1 _12092_ (.B1(_05522_),
    .Y(_00822_),
    .A1(_05398_),
    .A2(net2719));
 sg13g2_nand2_1 _12093_ (.Y(_05523_),
    .A(net245),
    .B(_05519_));
 sg13g2_o21ai_1 _12094_ (.B1(_05523_),
    .Y(_00823_),
    .A1(_05401_),
    .A2(net2717));
 sg13g2_nand2_1 _12095_ (.Y(_05524_),
    .A(net423),
    .B(_05519_));
 sg13g2_o21ai_1 _12096_ (.B1(_05524_),
    .Y(_00824_),
    .A1(_05404_),
    .A2(net2717));
 sg13g2_nand2_1 _12097_ (.Y(_05525_),
    .A(net748),
    .B(_05519_));
 sg13g2_o21ai_1 _12098_ (.B1(_05525_),
    .Y(_00825_),
    .A1(_05407_),
    .A2(net2717));
 sg13g2_nand2_1 _12099_ (.Y(_05526_),
    .A(net552),
    .B(_05519_));
 sg13g2_o21ai_1 _12100_ (.B1(_05526_),
    .Y(_00826_),
    .A1(_05410_),
    .A2(net2717));
 sg13g2_nand2_1 _12101_ (.Y(_05527_),
    .A(net633),
    .B(_05519_));
 sg13g2_nand4_1 _12102_ (.B(net2870),
    .C(net2899),
    .A(net3034),
    .Y(_05528_),
    .D(_05472_));
 sg13g2_o21ai_1 _12103_ (.B1(_05527_),
    .Y(_00827_),
    .A1(net2774),
    .A2(_05528_));
 sg13g2_nand2_1 _12104_ (.Y(_05529_),
    .A(net463),
    .B(_05519_));
 sg13g2_o21ai_1 _12105_ (.B1(_05529_),
    .Y(_00828_),
    .A1(_05415_),
    .A2(net2717));
 sg13g2_nand2_2 _12106_ (.Y(_05530_),
    .A(net2947),
    .B(_05443_));
 sg13g2_nand2_1 _12107_ (.Y(_05531_),
    .A(net584),
    .B(_05530_));
 sg13g2_o21ai_1 _12108_ (.B1(_05531_),
    .Y(_00829_),
    .A1(_05420_),
    .A2(net2718));
 sg13g2_nand2_1 _12109_ (.Y(_05532_),
    .A(net179),
    .B(_05530_));
 sg13g2_o21ai_1 _12110_ (.B1(_05532_),
    .Y(_00830_),
    .A1(_05423_),
    .A2(net2719));
 sg13g2_nand2_1 _12111_ (.Y(_05533_),
    .A(net798),
    .B(_05530_));
 sg13g2_o21ai_1 _12112_ (.B1(_05533_),
    .Y(_00831_),
    .A1(_05426_),
    .A2(net2717));
 sg13g2_nand2_1 _12113_ (.Y(_05534_),
    .A(net198),
    .B(_05530_));
 sg13g2_o21ai_1 _12114_ (.B1(_05534_),
    .Y(_00832_),
    .A1(_05429_),
    .A2(net2718));
 sg13g2_nand2_1 _12115_ (.Y(_05535_),
    .A(net259),
    .B(_05530_));
 sg13g2_o21ai_1 _12116_ (.B1(_05535_),
    .Y(_00833_),
    .A1(_05432_),
    .A2(net2718));
 sg13g2_nand2_1 _12117_ (.Y(_05536_),
    .A(net611),
    .B(_05530_));
 sg13g2_o21ai_1 _12118_ (.B1(_05536_),
    .Y(_00834_),
    .A1(_05435_),
    .A2(net2717));
 sg13g2_nand2_1 _12119_ (.Y(_05537_),
    .A(net276),
    .B(_05530_));
 sg13g2_o21ai_1 _12120_ (.B1(_05537_),
    .Y(_00835_),
    .A1(_05438_),
    .A2(net2719));
 sg13g2_nand2_1 _12121_ (.Y(_05538_),
    .A(net373),
    .B(_05530_));
 sg13g2_o21ai_1 _12122_ (.B1(_05538_),
    .Y(_00836_),
    .A1(_05441_),
    .A2(net2717));
 sg13g2_nand2_2 _12123_ (.Y(_05539_),
    .A(net1210),
    .B(_05256_));
 sg13g2_nand2_1 _12124_ (.Y(_05540_),
    .A(net215),
    .B(_05539_));
 sg13g2_o21ai_1 _12125_ (.B1(net216),
    .Y(_00837_),
    .A1(_05446_),
    .A2(net2720));
 sg13g2_nand2_1 _12126_ (.Y(_05541_),
    .A(net238),
    .B(_05539_));
 sg13g2_o21ai_1 _12127_ (.B1(net239),
    .Y(_00838_),
    .A1(_05449_),
    .A2(net2720));
 sg13g2_nand2_1 _12128_ (.Y(_05542_),
    .A(net385),
    .B(_05539_));
 sg13g2_o21ai_1 _12129_ (.B1(net386),
    .Y(_00839_),
    .A1(_05452_),
    .A2(net2720));
 sg13g2_nand2_1 _12130_ (.Y(_05543_),
    .A(net265),
    .B(_05539_));
 sg13g2_o21ai_1 _12131_ (.B1(_05543_),
    .Y(_00840_),
    .A1(_05455_),
    .A2(net2720));
 sg13g2_nand2_1 _12132_ (.Y(_05544_),
    .A(net517),
    .B(_05539_));
 sg13g2_o21ai_1 _12133_ (.B1(_05544_),
    .Y(_00841_),
    .A1(_05458_),
    .A2(net2720));
 sg13g2_nand2_1 _12134_ (.Y(_05545_),
    .A(net254),
    .B(_05539_));
 sg13g2_o21ai_1 _12135_ (.B1(net255),
    .Y(_00842_),
    .A1(_05461_),
    .A2(net2720));
 sg13g2_nand2_1 _12136_ (.Y(_05546_),
    .A(net713),
    .B(_05539_));
 sg13g2_o21ai_1 _12137_ (.B1(net714),
    .Y(_00843_),
    .A1(_05464_),
    .A2(net2720));
 sg13g2_nand2_1 _12138_ (.Y(_05547_),
    .A(net669),
    .B(_05539_));
 sg13g2_o21ai_1 _12139_ (.B1(net670),
    .Y(_00844_),
    .A1(_05467_),
    .A2(net2720));
 sg13g2_nor2_2 _12140_ (.A(net2789),
    .B(_05254_),
    .Y(_05548_));
 sg13g2_nand2_2 _12141_ (.Y(_05549_),
    .A(_05258_),
    .B(_05548_));
 sg13g2_nand2_1 _12142_ (.Y(_05550_),
    .A(net762),
    .B(_05549_));
 sg13g2_o21ai_1 _12143_ (.B1(_05550_),
    .Y(_00845_),
    .A1(net2791),
    .A2(_05264_));
 sg13g2_nand2_1 _12144_ (.Y(_05551_),
    .A(net667),
    .B(_05549_));
 sg13g2_o21ai_1 _12145_ (.B1(_05551_),
    .Y(_00846_),
    .A1(net2788),
    .A2(_05267_));
 sg13g2_nand2_1 _12146_ (.Y(_05552_),
    .A(net738),
    .B(_05549_));
 sg13g2_o21ai_1 _12147_ (.B1(_05552_),
    .Y(_00847_),
    .A1(net2791),
    .A2(_05270_));
 sg13g2_nand2_1 _12148_ (.Y(_05553_),
    .A(net691),
    .B(_05549_));
 sg13g2_o21ai_1 _12149_ (.B1(_05553_),
    .Y(_00848_),
    .A1(net2791),
    .A2(_05273_));
 sg13g2_nand2_1 _12150_ (.Y(_05554_),
    .A(net599),
    .B(_05549_));
 sg13g2_o21ai_1 _12151_ (.B1(_05554_),
    .Y(_00849_),
    .A1(net2790),
    .A2(_05276_));
 sg13g2_nand2_1 _12152_ (.Y(_05555_),
    .A(net799),
    .B(_05549_));
 sg13g2_o21ai_1 _12153_ (.B1(_05555_),
    .Y(_00850_),
    .A1(net2790),
    .A2(_05279_));
 sg13g2_nand2_1 _12154_ (.Y(_05556_),
    .A(net545),
    .B(_05549_));
 sg13g2_o21ai_1 _12155_ (.B1(_05556_),
    .Y(_00851_),
    .A1(net2788),
    .A2(_05282_));
 sg13g2_nand2_1 _12156_ (.Y(_05557_),
    .A(net788),
    .B(_05549_));
 sg13g2_o21ai_1 _12157_ (.B1(_05557_),
    .Y(_00852_),
    .A1(net2788),
    .A2(_05285_));
 sg13g2_nand2_2 _12158_ (.Y(_05558_),
    .A(_05288_),
    .B(_05548_));
 sg13g2_nand2_1 _12159_ (.Y(_05559_),
    .A(net495),
    .B(_05558_));
 sg13g2_o21ai_1 _12160_ (.B1(_05559_),
    .Y(_00853_),
    .A1(net2785),
    .A2(_05291_));
 sg13g2_nand2_1 _12161_ (.Y(_05560_),
    .A(net649),
    .B(_05558_));
 sg13g2_o21ai_1 _12162_ (.B1(_05560_),
    .Y(_00854_),
    .A1(net2788),
    .A2(_05294_));
 sg13g2_nand2_1 _12163_ (.Y(_05561_),
    .A(net548),
    .B(_05558_));
 sg13g2_o21ai_1 _12164_ (.B1(_05561_),
    .Y(_00855_),
    .A1(net2784),
    .A2(_05297_));
 sg13g2_nand2_1 _12165_ (.Y(_05562_),
    .A(net781),
    .B(_05558_));
 sg13g2_o21ai_1 _12166_ (.B1(_05562_),
    .Y(_00856_),
    .A1(net2787),
    .A2(_05300_));
 sg13g2_nand2_1 _12167_ (.Y(_05563_),
    .A(net406),
    .B(_05558_));
 sg13g2_o21ai_1 _12168_ (.B1(_05563_),
    .Y(_00857_),
    .A1(net2787),
    .A2(_05302_));
 sg13g2_nand2_1 _12169_ (.Y(_05564_),
    .A(net727),
    .B(_05558_));
 sg13g2_o21ai_1 _12170_ (.B1(_05564_),
    .Y(_00858_),
    .A1(net2787),
    .A2(_05305_));
 sg13g2_nand2_1 _12171_ (.Y(_05565_),
    .A(net285),
    .B(_05558_));
 sg13g2_o21ai_1 _12172_ (.B1(_05565_),
    .Y(_00859_),
    .A1(net2788),
    .A2(_05307_));
 sg13g2_nand2_1 _12173_ (.Y(_05566_),
    .A(net449),
    .B(_05558_));
 sg13g2_o21ai_1 _12174_ (.B1(_05566_),
    .Y(_00860_),
    .A1(net2785),
    .A2(_05310_));
 sg13g2_nand2_2 _12175_ (.Y(_05567_),
    .A(_05312_),
    .B(_05548_));
 sg13g2_nand2_1 _12176_ (.Y(_05568_),
    .A(net549),
    .B(_05567_));
 sg13g2_o21ai_1 _12177_ (.B1(_05568_),
    .Y(_00861_),
    .A1(net2785),
    .A2(_05316_));
 sg13g2_nand2_1 _12178_ (.Y(_05569_),
    .A(net213),
    .B(_05567_));
 sg13g2_o21ai_1 _12179_ (.B1(_05569_),
    .Y(_00862_),
    .A1(net2788),
    .A2(_05319_));
 sg13g2_nand2_1 _12180_ (.Y(_05570_),
    .A(net498),
    .B(_05567_));
 sg13g2_o21ai_1 _12181_ (.B1(_05570_),
    .Y(_00863_),
    .A1(net2784),
    .A2(_05322_));
 sg13g2_nand2_1 _12182_ (.Y(_05571_),
    .A(net234),
    .B(_05567_));
 sg13g2_o21ai_1 _12183_ (.B1(_05571_),
    .Y(_00864_),
    .A1(net2787),
    .A2(_05325_));
 sg13g2_nand2_1 _12184_ (.Y(_05572_),
    .A(net193),
    .B(_05567_));
 sg13g2_o21ai_1 _12185_ (.B1(_05572_),
    .Y(_00865_),
    .A1(net2787),
    .A2(_05328_));
 sg13g2_nand2_1 _12186_ (.Y(_05573_),
    .A(net197),
    .B(_05567_));
 sg13g2_o21ai_1 _12187_ (.B1(_05573_),
    .Y(_00866_),
    .A1(net2787),
    .A2(_05331_));
 sg13g2_nand2_1 _12188_ (.Y(_05574_),
    .A(net419),
    .B(_05567_));
 sg13g2_o21ai_1 _12189_ (.B1(_05574_),
    .Y(_00867_),
    .A1(net2788),
    .A2(_05334_));
 sg13g2_nand2_1 _12190_ (.Y(_05575_),
    .A(net183),
    .B(_05567_));
 sg13g2_o21ai_1 _12191_ (.B1(_05575_),
    .Y(_00868_),
    .A1(net2784),
    .A2(_05337_));
 sg13g2_nand3b_1 _12192_ (.B(net2903),
    .C(_05548_),
    .Y(_05576_),
    .A_N(net3053));
 sg13g2_nand2_1 _12193_ (.Y(_05577_),
    .A(net427),
    .B(_05576_));
 sg13g2_o21ai_1 _12194_ (.B1(_05577_),
    .Y(_00869_),
    .A1(net2781),
    .A2(_05343_));
 sg13g2_nand2_1 _12195_ (.Y(_05578_),
    .A(net801),
    .B(_05576_));
 sg13g2_o21ai_1 _12196_ (.B1(_05578_),
    .Y(_00870_),
    .A1(net2781),
    .A2(_05346_));
 sg13g2_nand2_1 _12197_ (.Y(_05579_),
    .A(net241),
    .B(_05576_));
 sg13g2_o21ai_1 _12198_ (.B1(_05579_),
    .Y(_00871_),
    .A1(net2783),
    .A2(_05349_));
 sg13g2_nand2_1 _12199_ (.Y(_05580_),
    .A(net329),
    .B(_05576_));
 sg13g2_o21ai_1 _12200_ (.B1(_05580_),
    .Y(_00872_),
    .A1(net2783),
    .A2(_05352_));
 sg13g2_nand2_1 _12201_ (.Y(_05581_),
    .A(net761),
    .B(_05576_));
 sg13g2_o21ai_1 _12202_ (.B1(_05581_),
    .Y(_00873_),
    .A1(net2786),
    .A2(_05355_));
 sg13g2_nand2_1 _12203_ (.Y(_05582_),
    .A(net488),
    .B(_05576_));
 sg13g2_o21ai_1 _12204_ (.B1(_05582_),
    .Y(_00874_),
    .A1(net2786),
    .A2(_05358_));
 sg13g2_nand2_1 _12205_ (.Y(_05583_),
    .A(net557),
    .B(_05576_));
 sg13g2_o21ai_1 _12206_ (.B1(_05583_),
    .Y(_00875_),
    .A1(net2782),
    .A2(_05361_));
 sg13g2_nand2_1 _12207_ (.Y(_05584_),
    .A(net331),
    .B(_05576_));
 sg13g2_o21ai_1 _12208_ (.B1(_05584_),
    .Y(_00876_),
    .A1(net2781),
    .A2(_05364_));
 sg13g2_nand2_2 _12209_ (.Y(_05585_),
    .A(_05366_),
    .B(_05548_));
 sg13g2_nand2_1 _12210_ (.Y(_05586_),
    .A(net184),
    .B(_05585_));
 sg13g2_o21ai_1 _12211_ (.B1(_05586_),
    .Y(_00877_),
    .A1(net2781),
    .A2(_05370_));
 sg13g2_nand2_1 _12212_ (.Y(_05587_),
    .A(net358),
    .B(_05585_));
 sg13g2_o21ai_1 _12213_ (.B1(_05587_),
    .Y(_00878_),
    .A1(net2781),
    .A2(_05373_));
 sg13g2_nand2_1 _12214_ (.Y(_05588_),
    .A(net766),
    .B(_05585_));
 sg13g2_o21ai_1 _12215_ (.B1(_05588_),
    .Y(_00879_),
    .A1(net2783),
    .A2(_05376_));
 sg13g2_nand2_1 _12216_ (.Y(_05589_),
    .A(net473),
    .B(_05585_));
 sg13g2_o21ai_1 _12217_ (.B1(_05589_),
    .Y(_00880_),
    .A1(net2783),
    .A2(_05379_));
 sg13g2_nand2_1 _12218_ (.Y(_05590_),
    .A(net778),
    .B(_05585_));
 sg13g2_o21ai_1 _12219_ (.B1(_05590_),
    .Y(_00881_),
    .A1(net2786),
    .A2(_05382_));
 sg13g2_nand2_1 _12220_ (.Y(_05591_),
    .A(net288),
    .B(_05585_));
 sg13g2_o21ai_1 _12221_ (.B1(_05591_),
    .Y(_00882_),
    .A1(net2786),
    .A2(_05385_));
 sg13g2_nand2_1 _12222_ (.Y(_05592_),
    .A(net677),
    .B(_05585_));
 sg13g2_o21ai_1 _12223_ (.B1(_05592_),
    .Y(_00883_),
    .A1(net2781),
    .A2(_05388_));
 sg13g2_nand2_1 _12224_ (.Y(_05593_),
    .A(net634),
    .B(_05585_));
 sg13g2_o21ai_1 _12225_ (.B1(_05593_),
    .Y(_00884_),
    .A1(net2781),
    .A2(_05391_));
 sg13g2_nand2_2 _12226_ (.Y(_05594_),
    .A(_05393_),
    .B(_05548_));
 sg13g2_nand2_1 _12227_ (.Y(_05595_),
    .A(net513),
    .B(_05594_));
 sg13g2_o21ai_1 _12228_ (.B1(_05595_),
    .Y(_00885_),
    .A1(net2782),
    .A2(_05396_));
 sg13g2_nand2_1 _12229_ (.Y(_05596_),
    .A(net627),
    .B(_05594_));
 sg13g2_o21ai_1 _12230_ (.B1(_05596_),
    .Y(_00886_),
    .A1(net2784),
    .A2(_05399_));
 sg13g2_nand2_1 _12231_ (.Y(_05597_),
    .A(net581),
    .B(_05594_));
 sg13g2_o21ai_1 _12232_ (.B1(_05597_),
    .Y(_00887_),
    .A1(net2782),
    .A2(_05402_));
 sg13g2_nand2_1 _12233_ (.Y(_05598_),
    .A(net270),
    .B(_05594_));
 sg13g2_o21ai_1 _12234_ (.B1(_05598_),
    .Y(_00888_),
    .A1(net2782),
    .A2(_05405_));
 sg13g2_nand2_1 _12235_ (.Y(_05599_),
    .A(net335),
    .B(_05594_));
 sg13g2_o21ai_1 _12236_ (.B1(_05599_),
    .Y(_00889_),
    .A1(net2786),
    .A2(_05408_));
 sg13g2_nand2_1 _12237_ (.Y(_05600_),
    .A(net375),
    .B(_05594_));
 sg13g2_o21ai_1 _12238_ (.B1(_05600_),
    .Y(_00890_),
    .A1(net2787),
    .A2(_05411_));
 sg13g2_nand2_1 _12239_ (.Y(_05601_),
    .A(net333),
    .B(_05594_));
 sg13g2_o21ai_1 _12240_ (.B1(_05601_),
    .Y(_00891_),
    .A1(net2784),
    .A2(_05413_));
 sg13g2_nand2_1 _12241_ (.Y(_05602_),
    .A(net348),
    .B(_05594_));
 sg13g2_o21ai_1 _12242_ (.B1(_05602_),
    .Y(_00892_),
    .A1(net2784),
    .A2(_05416_));
 sg13g2_nand2_2 _12243_ (.Y(_05603_),
    .A(_05417_),
    .B(_05548_));
 sg13g2_nand2_1 _12244_ (.Y(_05604_),
    .A(net313),
    .B(_05603_));
 sg13g2_o21ai_1 _12245_ (.B1(_05604_),
    .Y(_00893_),
    .A1(net2781),
    .A2(_05421_));
 sg13g2_nand2_1 _12246_ (.Y(_05605_),
    .A(net802),
    .B(_05603_));
 sg13g2_o21ai_1 _12247_ (.B1(_05605_),
    .Y(_00894_),
    .A1(net2784),
    .A2(_05424_));
 sg13g2_nand2_1 _12248_ (.Y(_05606_),
    .A(net181),
    .B(_05603_));
 sg13g2_o21ai_1 _12249_ (.B1(_05606_),
    .Y(_00895_),
    .A1(net2782),
    .A2(_05427_));
 sg13g2_nand2_1 _12250_ (.Y(_05607_),
    .A(net283),
    .B(_05603_));
 sg13g2_o21ai_1 _12251_ (.B1(_05607_),
    .Y(_00896_),
    .A1(net2782),
    .A2(_05430_));
 sg13g2_nand2_1 _12252_ (.Y(_05608_),
    .A(net546),
    .B(_05603_));
 sg13g2_o21ai_1 _12253_ (.B1(_05608_),
    .Y(_00897_),
    .A1(net2786),
    .A2(_05433_));
 sg13g2_nand2_1 _12254_ (.Y(_05609_),
    .A(net284),
    .B(_05603_));
 sg13g2_o21ai_1 _12255_ (.B1(_05609_),
    .Y(_00898_),
    .A1(net2787),
    .A2(_05436_));
 sg13g2_nand2_1 _12256_ (.Y(_05610_),
    .A(net804),
    .B(_05603_));
 sg13g2_o21ai_1 _12257_ (.B1(_05610_),
    .Y(_00899_),
    .A1(net2782),
    .A2(_05439_));
 sg13g2_nand2_1 _12258_ (.Y(_05611_),
    .A(net474),
    .B(_05603_));
 sg13g2_o21ai_1 _12259_ (.B1(_05611_),
    .Y(_00900_),
    .A1(net2784),
    .A2(_05442_));
 sg13g2_and2_2 _12260_ (.A(net3054),
    .B(_05548_),
    .X(_05612_));
 sg13g2_nand2_2 _12261_ (.Y(_05613_),
    .A(net2982),
    .B(_05612_));
 sg13g2_nand2_1 _12262_ (.Y(_05614_),
    .A(net795),
    .B(_05613_));
 sg13g2_o21ai_1 _12263_ (.B1(_05614_),
    .Y(_00901_),
    .A1(net2790),
    .A2(_05447_));
 sg13g2_nand2_1 _12264_ (.Y(_05615_),
    .A(net521),
    .B(_05613_));
 sg13g2_o21ai_1 _12265_ (.B1(_05615_),
    .Y(_00902_),
    .A1(net2792),
    .A2(_05450_));
 sg13g2_nand2_1 _12266_ (.Y(_05616_),
    .A(net516),
    .B(_05613_));
 sg13g2_o21ai_1 _12267_ (.B1(_05616_),
    .Y(_00903_),
    .A1(net2792),
    .A2(_05453_));
 sg13g2_nand2_1 _12268_ (.Y(_05617_),
    .A(net355),
    .B(_05613_));
 sg13g2_o21ai_1 _12269_ (.B1(_05617_),
    .Y(_00904_),
    .A1(net2792),
    .A2(_05456_));
 sg13g2_nand2_1 _12270_ (.Y(_05618_),
    .A(net448),
    .B(_05613_));
 sg13g2_o21ai_1 _12271_ (.B1(_05618_),
    .Y(_00905_),
    .A1(net2791),
    .A2(_05459_));
 sg13g2_nand2_1 _12272_ (.Y(_05619_),
    .A(net687),
    .B(_05613_));
 sg13g2_o21ai_1 _12273_ (.B1(_05619_),
    .Y(_00906_),
    .A1(net2791),
    .A2(_05462_));
 sg13g2_nand2_1 _12274_ (.Y(_05620_),
    .A(net505),
    .B(_05613_));
 sg13g2_o21ai_1 _12275_ (.B1(_05620_),
    .Y(_00907_),
    .A1(net2791),
    .A2(_05465_));
 sg13g2_nand2_1 _12276_ (.Y(_05621_),
    .A(net292),
    .B(_05613_));
 sg13g2_o21ai_1 _12277_ (.B1(_05621_),
    .Y(_00908_),
    .A1(net2791),
    .A2(_05468_));
 sg13g2_nand2_2 _12278_ (.Y(_05622_),
    .A(net2912),
    .B(_05612_));
 sg13g2_nand2_1 _12279_ (.Y(_05623_),
    .A(net490),
    .B(_05622_));
 sg13g2_nand2b_1 _12280_ (.Y(_05624_),
    .B(_05472_),
    .A_N(net2786));
 sg13g2_o21ai_1 _12281_ (.B1(_05623_),
    .Y(_00909_),
    .A1(_05263_),
    .A2(net2738));
 sg13g2_nand2_1 _12282_ (.Y(_05625_),
    .A(net779),
    .B(_05622_));
 sg13g2_o21ai_1 _12283_ (.B1(_05625_),
    .Y(_00910_),
    .A1(_05266_),
    .A2(net2738));
 sg13g2_nand2_1 _12284_ (.Y(_05626_),
    .A(net431),
    .B(_05622_));
 sg13g2_o21ai_1 _12285_ (.B1(_05626_),
    .Y(_00911_),
    .A1(_05269_),
    .A2(net2738));
 sg13g2_nand2_1 _12286_ (.Y(_05627_),
    .A(net673),
    .B(_05622_));
 sg13g2_o21ai_1 _12287_ (.B1(_05627_),
    .Y(_00912_),
    .A1(_05272_),
    .A2(net2738));
 sg13g2_nand2_1 _12288_ (.Y(_05628_),
    .A(net219),
    .B(_05622_));
 sg13g2_o21ai_1 _12289_ (.B1(_05628_),
    .Y(_00913_),
    .A1(_05275_),
    .A2(net2738));
 sg13g2_nand2_1 _12290_ (.Y(_05629_),
    .A(net736),
    .B(_05622_));
 sg13g2_o21ai_1 _12291_ (.B1(_05629_),
    .Y(_00914_),
    .A1(_05278_),
    .A2(net2737));
 sg13g2_nand2_1 _12292_ (.Y(_05630_),
    .A(net359),
    .B(_05622_));
 sg13g2_o21ai_1 _12293_ (.B1(_05630_),
    .Y(_00915_),
    .A1(_05281_),
    .A2(net2737));
 sg13g2_nand2_1 _12294_ (.Y(_05631_),
    .A(net694),
    .B(_05622_));
 sg13g2_o21ai_1 _12295_ (.B1(_05631_),
    .Y(_00916_),
    .A1(_05284_),
    .A2(net2738));
 sg13g2_nand2_2 _12296_ (.Y(_05632_),
    .A(net2909),
    .B(_05612_));
 sg13g2_nand2_1 _12297_ (.Y(_05633_),
    .A(net659),
    .B(_05632_));
 sg13g2_o21ai_1 _12298_ (.B1(_05633_),
    .Y(_00917_),
    .A1(net2790),
    .A2(_05482_));
 sg13g2_nand2_1 _12299_ (.Y(_05634_),
    .A(net827),
    .B(_05632_));
 sg13g2_o21ai_1 _12300_ (.B1(_05634_),
    .Y(_00918_),
    .A1(_05293_),
    .A2(net2739));
 sg13g2_nand2_1 _12301_ (.Y(_05635_),
    .A(net759),
    .B(_05632_));
 sg13g2_o21ai_1 _12302_ (.B1(_05635_),
    .Y(_00919_),
    .A1(_05296_),
    .A2(net2739));
 sg13g2_nand2_1 _12303_ (.Y(_05636_),
    .A(net253),
    .B(_05632_));
 sg13g2_o21ai_1 _12304_ (.B1(_05636_),
    .Y(_00920_),
    .A1(_05299_),
    .A2(net2740));
 sg13g2_nand2_1 _12305_ (.Y(_05637_),
    .A(net478),
    .B(_05632_));
 sg13g2_o21ai_1 _12306_ (.B1(_05637_),
    .Y(_00921_),
    .A1(net2790),
    .A2(_05487_));
 sg13g2_nand2_1 _12307_ (.Y(_05638_),
    .A(net763),
    .B(_05632_));
 sg13g2_o21ai_1 _12308_ (.B1(_05638_),
    .Y(_00922_),
    .A1(_05304_),
    .A2(net2739));
 sg13g2_nand2_1 _12309_ (.Y(_05639_),
    .A(net813),
    .B(_05632_));
 sg13g2_o21ai_1 _12310_ (.B1(_05639_),
    .Y(_00923_),
    .A1(net2790),
    .A2(_05490_));
 sg13g2_nand2_1 _12311_ (.Y(_05640_),
    .A(net446),
    .B(_05632_));
 sg13g2_o21ai_1 _12312_ (.B1(_05640_),
    .Y(_00924_),
    .A1(_05309_),
    .A2(net2740));
 sg13g2_nand2_2 _12313_ (.Y(_05641_),
    .A(net2906),
    .B(_05612_));
 sg13g2_nand2_1 _12314_ (.Y(_05642_),
    .A(net675),
    .B(_05641_));
 sg13g2_o21ai_1 _12315_ (.B1(_05642_),
    .Y(_00925_),
    .A1(_05315_),
    .A2(net2736));
 sg13g2_nand2_1 _12316_ (.Y(_05643_),
    .A(net646),
    .B(_05641_));
 sg13g2_o21ai_1 _12317_ (.B1(_05643_),
    .Y(_00926_),
    .A1(_05318_),
    .A2(net2739));
 sg13g2_nand2_1 _12318_ (.Y(_05644_),
    .A(net596),
    .B(_05641_));
 sg13g2_o21ai_1 _12319_ (.B1(_05644_),
    .Y(_00927_),
    .A1(_05321_),
    .A2(net2739));
 sg13g2_nand2_1 _12320_ (.Y(_05645_),
    .A(net209),
    .B(_05641_));
 sg13g2_o21ai_1 _12321_ (.B1(_05645_),
    .Y(_00928_),
    .A1(_05324_),
    .A2(net2739));
 sg13g2_nand2_1 _12322_ (.Y(_05646_),
    .A(net679),
    .B(_05641_));
 sg13g2_o21ai_1 _12323_ (.B1(_05646_),
    .Y(_00929_),
    .A1(_05327_),
    .A2(net2736));
 sg13g2_nand2_1 _12324_ (.Y(_05647_),
    .A(net718),
    .B(_05641_));
 sg13g2_o21ai_1 _12325_ (.B1(_05647_),
    .Y(_00930_),
    .A1(_05330_),
    .A2(net2739));
 sg13g2_nand2_1 _12326_ (.Y(_05648_),
    .A(net457),
    .B(_05641_));
 sg13g2_o21ai_1 _12327_ (.B1(_05648_),
    .Y(_00931_),
    .A1(_05333_),
    .A2(net2736));
 sg13g2_nand2_1 _12328_ (.Y(_05649_),
    .A(net853),
    .B(_05641_));
 sg13g2_o21ai_1 _12329_ (.B1(_05649_),
    .Y(_00932_),
    .A1(_05336_),
    .A2(net2739));
 sg13g2_nand2_2 _12330_ (.Y(_05650_),
    .A(net2904),
    .B(_05612_));
 sg13g2_nand2_1 _12331_ (.Y(_05651_),
    .A(net305),
    .B(_05650_));
 sg13g2_o21ai_1 _12332_ (.B1(_05651_),
    .Y(_00933_),
    .A1(_05342_),
    .A2(net2735));
 sg13g2_nand2_1 _12333_ (.Y(_05652_),
    .A(net698),
    .B(_05650_));
 sg13g2_o21ai_1 _12334_ (.B1(_05652_),
    .Y(_00934_),
    .A1(_05345_),
    .A2(net2734));
 sg13g2_nand2_1 _12335_ (.Y(_05653_),
    .A(net361),
    .B(_05650_));
 sg13g2_o21ai_1 _12336_ (.B1(_05653_),
    .Y(_00935_),
    .A1(_05348_),
    .A2(net2734));
 sg13g2_nand2_1 _12337_ (.Y(_05654_),
    .A(net458),
    .B(_05650_));
 sg13g2_o21ai_1 _12338_ (.B1(_05654_),
    .Y(_00936_),
    .A1(_05351_),
    .A2(net2734));
 sg13g2_nand2_1 _12339_ (.Y(_05655_),
    .A(net330),
    .B(_05650_));
 sg13g2_o21ai_1 _12340_ (.B1(_05655_),
    .Y(_00937_),
    .A1(_05354_),
    .A2(net2734));
 sg13g2_nand2_1 _12341_ (.Y(_05656_),
    .A(net400),
    .B(_05650_));
 sg13g2_o21ai_1 _12342_ (.B1(_05656_),
    .Y(_00938_),
    .A1(_05357_),
    .A2(net2734));
 sg13g2_nand2_1 _12343_ (.Y(_05657_),
    .A(net321),
    .B(_05650_));
 sg13g2_o21ai_1 _12344_ (.B1(_05657_),
    .Y(_00939_),
    .A1(_05360_),
    .A2(net2736));
 sg13g2_nand2_1 _12345_ (.Y(_05658_),
    .A(net326),
    .B(_05650_));
 sg13g2_o21ai_1 _12346_ (.B1(_05658_),
    .Y(_00940_),
    .A1(_05363_),
    .A2(net2735));
 sg13g2_nand2_2 _12347_ (.Y(_05659_),
    .A(net2901),
    .B(_05612_));
 sg13g2_nand2_1 _12348_ (.Y(_05660_),
    .A(net645),
    .B(_05659_));
 sg13g2_o21ai_1 _12349_ (.B1(_05660_),
    .Y(_00941_),
    .A1(_05369_),
    .A2(net2734));
 sg13g2_nand2_1 _12350_ (.Y(_05661_),
    .A(net541),
    .B(_05659_));
 sg13g2_o21ai_1 _12351_ (.B1(_05661_),
    .Y(_00942_),
    .A1(_05372_),
    .A2(net2737));
 sg13g2_nand2_1 _12352_ (.Y(_05662_),
    .A(net421),
    .B(_05659_));
 sg13g2_o21ai_1 _12353_ (.B1(_05662_),
    .Y(_00943_),
    .A1(_05375_),
    .A2(net2737));
 sg13g2_nand2_1 _12354_ (.Y(_05663_),
    .A(net468),
    .B(_05659_));
 sg13g2_o21ai_1 _12355_ (.B1(_05663_),
    .Y(_00944_),
    .A1(_05378_),
    .A2(net2737));
 sg13g2_nand2_1 _12356_ (.Y(_05664_),
    .A(net492),
    .B(_05659_));
 sg13g2_o21ai_1 _12357_ (.B1(_05664_),
    .Y(_00945_),
    .A1(_05381_),
    .A2(net2737));
 sg13g2_nand2_1 _12358_ (.Y(_05665_),
    .A(net615),
    .B(_05659_));
 sg13g2_o21ai_1 _12359_ (.B1(_05665_),
    .Y(_00946_),
    .A1(_05384_),
    .A2(net2737));
 sg13g2_nand2_1 _12360_ (.Y(_05666_),
    .A(net567),
    .B(_05659_));
 sg13g2_o21ai_1 _12361_ (.B1(_05666_),
    .Y(_00947_),
    .A1(_05387_),
    .A2(net2734));
 sg13g2_nand2_1 _12362_ (.Y(_05667_),
    .A(net370),
    .B(_05659_));
 sg13g2_o21ai_1 _12363_ (.B1(_05667_),
    .Y(_00948_),
    .A1(_05390_),
    .A2(net2737));
 sg13g2_nand2_2 _12364_ (.Y(_05668_),
    .A(net2898),
    .B(_05612_));
 sg13g2_nand2_1 _12365_ (.Y(_05669_),
    .A(net745),
    .B(_05668_));
 sg13g2_o21ai_1 _12366_ (.B1(_05669_),
    .Y(_00949_),
    .A1(net2790),
    .A2(_05521_));
 sg13g2_nand2_1 _12367_ (.Y(_05670_),
    .A(net476),
    .B(_05668_));
 sg13g2_o21ai_1 _12368_ (.B1(_05670_),
    .Y(_00950_),
    .A1(_05398_),
    .A2(net2733));
 sg13g2_nand2_1 _12369_ (.Y(_05671_),
    .A(net724),
    .B(_05668_));
 sg13g2_o21ai_1 _12370_ (.B1(_05671_),
    .Y(_00951_),
    .A1(_05401_),
    .A2(net2732));
 sg13g2_nand2_1 _12371_ (.Y(_05672_),
    .A(net401),
    .B(_05668_));
 sg13g2_o21ai_1 _12372_ (.B1(_05672_),
    .Y(_00952_),
    .A1(_05404_),
    .A2(net2732));
 sg13g2_nand2_1 _12373_ (.Y(_05673_),
    .A(net576),
    .B(_05668_));
 sg13g2_o21ai_1 _12374_ (.B1(_05673_),
    .Y(_00953_),
    .A1(_05407_),
    .A2(net2732));
 sg13g2_nand2_1 _12375_ (.Y(_05674_),
    .A(net500),
    .B(_05668_));
 sg13g2_o21ai_1 _12376_ (.B1(_05674_),
    .Y(_00954_),
    .A1(_05410_),
    .A2(net2732));
 sg13g2_nand2_1 _12377_ (.Y(_05675_),
    .A(net308),
    .B(_05668_));
 sg13g2_o21ai_1 _12378_ (.B1(_05675_),
    .Y(_00955_),
    .A1(net2786),
    .A2(_05528_));
 sg13g2_nand2_1 _12379_ (.Y(_05676_),
    .A(net792),
    .B(_05668_));
 sg13g2_o21ai_1 _12380_ (.B1(_05676_),
    .Y(_00956_),
    .A1(_05415_),
    .A2(net2733));
 sg13g2_nand2_1 _12381_ (.Y(_05677_),
    .A(net307),
    .B(_05241_));
 sg13g2_o21ai_1 _12382_ (.B1(_05677_),
    .Y(_00957_),
    .A1(_05420_),
    .A2(net2736));
 sg13g2_nand2_1 _12383_ (.Y(_05678_),
    .A(net413),
    .B(_05241_));
 sg13g2_o21ai_1 _12384_ (.B1(_05678_),
    .Y(_00958_),
    .A1(_05423_),
    .A2(net2733));
 sg13g2_nand2_1 _12385_ (.Y(_05679_),
    .A(net258),
    .B(_05241_));
 sg13g2_o21ai_1 _12386_ (.B1(_05679_),
    .Y(_00959_),
    .A1(_05426_),
    .A2(net2732));
 sg13g2_nand2_1 _12387_ (.Y(_05680_),
    .A(net167),
    .B(_05241_));
 sg13g2_o21ai_1 _12388_ (.B1(_05680_),
    .Y(_00960_),
    .A1(_05429_),
    .A2(net2732));
 sg13g2_nand2_1 _12389_ (.Y(_05681_),
    .A(net272),
    .B(_05241_));
 sg13g2_o21ai_1 _12390_ (.B1(_05681_),
    .Y(_00961_),
    .A1(_05432_),
    .A2(net2734));
 sg13g2_nand2_1 _12391_ (.Y(_05682_),
    .A(net206),
    .B(_05241_));
 sg13g2_o21ai_1 _12392_ (.B1(_05682_),
    .Y(_00962_),
    .A1(_05435_),
    .A2(net2732));
 sg13g2_nand2_1 _12393_ (.Y(_05683_),
    .A(net369),
    .B(_05241_));
 sg13g2_o21ai_1 _12394_ (.B1(_05683_),
    .Y(_00963_),
    .A1(_05438_),
    .A2(net2733));
 sg13g2_nand2_1 _12395_ (.Y(_05684_),
    .A(net733),
    .B(_05241_));
 sg13g2_o21ai_1 _12396_ (.B1(_05684_),
    .Y(_00964_),
    .A1(_05441_),
    .A2(net2732));
 sg13g2_mux2_1 _12397_ (.A0(net3403),
    .A1(net992),
    .S(_03746_),
    .X(_00965_));
 sg13g2_mux2_1 _12398_ (.A0(net3399),
    .A1(net997),
    .S(net2857),
    .X(_00966_));
 sg13g2_mux2_1 _12399_ (.A0(net3395),
    .A1(net1018),
    .S(net2857),
    .X(_00967_));
 sg13g2_mux2_1 _12400_ (.A0(net3392),
    .A1(net1020),
    .S(net2857),
    .X(_00968_));
 sg13g2_nand2_1 _12401_ (.Y(_05685_),
    .A(net845),
    .B(net2857));
 sg13g2_o21ai_1 _12402_ (.B1(_05685_),
    .Y(_00969_),
    .A1(_01046_),
    .A2(net2857));
 sg13g2_mux2_1 _12403_ (.A0(net3385),
    .A1(net1019),
    .S(net2857),
    .X(_00970_));
 sg13g2_mux2_1 _12404_ (.A0(net3381),
    .A1(net1014),
    .S(net2857),
    .X(_00971_));
 sg13g2_nor2_1 _12405_ (.A(net3378),
    .B(_03746_),
    .Y(_05686_));
 sg13g2_a21oi_1 _12406_ (.A1(_01176_),
    .A2(_03746_),
    .Y(_00972_),
    .B1(_05686_));
 sg13g2_nor4_2 _12407_ (.A(\u_toplayer.u_layer1.u_neuron.instCtrl.state[0] ),
    .B(_01030_),
    .C(net968),
    .Y(_05687_),
    .D(_03748_));
 sg13g2_nor4_1 _12408_ (.A(net3027),
    .B(\u_toplayer.u_layer1.u_neuron.acc[10] ),
    .C(\u_toplayer.u_layer1.u_neuron.acc[11] ),
    .D(\u_toplayer.u_layer1.u_neuron.acc[9] ),
    .Y(_05688_));
 sg13g2_nor4_1 _12409_ (.A(\u_toplayer.u_layer1.u_neuron.acc[7] ),
    .B(\u_toplayer.u_layer1.u_neuron.acc[15] ),
    .C(\u_toplayer.u_layer1.u_neuron.acc[14] ),
    .D(\u_toplayer.u_layer1.u_neuron.acc[12] ),
    .Y(_05689_));
 sg13g2_nor4_1 _12410_ (.A(\u_toplayer.u_layer1.u_neuron.acc[8] ),
    .B(\u_toplayer.u_layer1.u_neuron.acc[22] ),
    .C(\u_toplayer.u_layer1.u_neuron.acc[21] ),
    .D(\u_toplayer.u_layer1.u_neuron.acc[20] ),
    .Y(_05690_));
 sg13g2_nor4_1 _12411_ (.A(net3025),
    .B(\u_toplayer.u_layer1.u_neuron.acc[19] ),
    .C(net3026),
    .D(\u_toplayer.u_layer1.u_neuron.acc[17] ),
    .Y(_05691_));
 sg13g2_and3_1 _12412_ (.X(_05692_),
    .A(_05688_),
    .B(_05689_),
    .C(_05691_));
 sg13g2_a21oi_2 _12413_ (.B1(\u_toplayer.u_layer1.u_neuron.acc[23] ),
    .Y(_05693_),
    .A2(_05692_),
    .A1(_05690_));
 sg13g2_nor4_1 _12414_ (.A(\u_toplayer.u_layer1.u_neuron.acc[3] ),
    .B(\u_toplayer.u_layer1.u_neuron.acc[2] ),
    .C(\u_toplayer.u_layer1.u_neuron.acc[1] ),
    .D(\u_toplayer.u_layer1.u_neuron.acc[0] ),
    .Y(_05694_));
 sg13g2_nor3_1 _12415_ (.A(_01152_),
    .B(\u_toplayer.u_layer1.u_neuron.acc[6] ),
    .C(\u_toplayer.u_layer1.u_neuron.acc[5] ),
    .Y(_05695_));
 sg13g2_nand3_1 _12416_ (.B(_05694_),
    .C(_05695_),
    .A(_01155_),
    .Y(_05696_));
 sg13g2_nand4_1 _12417_ (.B(net3029),
    .C(\u_toplayer.u_layer1.u_neuron.acc[11] ),
    .A(net3027),
    .Y(_05697_),
    .D(\u_toplayer.u_layer1.u_neuron.acc[9] ));
 sg13g2_nand4_1 _12418_ (.B(\u_toplayer.u_layer1.u_neuron.acc[15] ),
    .C(\u_toplayer.u_layer1.u_neuron.acc[14] ),
    .A(\u_toplayer.u_layer1.u_neuron.acc[7] ),
    .Y(_05698_),
    .D(net3028));
 sg13g2_nand4_1 _12419_ (.B(\u_toplayer.u_layer1.u_neuron.acc[22] ),
    .C(\u_toplayer.u_layer1.u_neuron.acc[21] ),
    .A(\u_toplayer.u_layer1.u_neuron.acc[8] ),
    .Y(_05699_),
    .D(\u_toplayer.u_layer1.u_neuron.acc[20] ));
 sg13g2_nand4_1 _12420_ (.B(\u_toplayer.u_layer1.u_neuron.acc[19] ),
    .C(net3026),
    .A(net3025),
    .Y(_05700_),
    .D(\u_toplayer.u_layer1.u_neuron.acc[17] ));
 sg13g2_nor4_2 _12421_ (.A(_05697_),
    .B(_05698_),
    .C(_05699_),
    .Y(_05701_),
    .D(_05700_));
 sg13g2_a21oi_1 _12422_ (.A1(_05696_),
    .A2(_05701_),
    .Y(_05702_),
    .B1(_01166_));
 sg13g2_nor2b_2 _12423_ (.A(_05702_),
    .B_N(_05687_),
    .Y(_05703_));
 sg13g2_o21ai_1 _12424_ (.B1(_05703_),
    .Y(_05704_),
    .A1(\u_toplayer.u_layer1.u_neuron.acc[0] ),
    .A2(_05693_));
 sg13g2_o21ai_1 _12425_ (.B1(_05704_),
    .Y(_00973_),
    .A1(_01178_),
    .A2(net2842));
 sg13g2_o21ai_1 _12426_ (.B1(_05703_),
    .Y(_05705_),
    .A1(\u_toplayer.u_layer1.u_neuron.acc[1] ),
    .A2(_05693_));
 sg13g2_o21ai_1 _12427_ (.B1(_05705_),
    .Y(_00974_),
    .A1(_01179_),
    .A2(net2842));
 sg13g2_o21ai_1 _12428_ (.B1(_05703_),
    .Y(_05706_),
    .A1(\u_toplayer.u_layer1.u_neuron.acc[2] ),
    .A2(_05693_));
 sg13g2_o21ai_1 _12429_ (.B1(_05706_),
    .Y(_00975_),
    .A1(_01180_),
    .A2(net2842));
 sg13g2_o21ai_1 _12430_ (.B1(_05703_),
    .Y(_05707_),
    .A1(\u_toplayer.u_layer1.u_neuron.acc[3] ),
    .A2(_05693_));
 sg13g2_o21ai_1 _12431_ (.B1(_05707_),
    .Y(_00976_),
    .A1(_01181_),
    .A2(net2842));
 sg13g2_o21ai_1 _12432_ (.B1(_05703_),
    .Y(_05708_),
    .A1(\u_toplayer.u_layer1.u_neuron.acc[4] ),
    .A2(_05693_));
 sg13g2_o21ai_1 _12433_ (.B1(_05708_),
    .Y(_00977_),
    .A1(_01182_),
    .A2(net2842));
 sg13g2_o21ai_1 _12434_ (.B1(_05703_),
    .Y(_05709_),
    .A1(net3030),
    .A2(_05693_));
 sg13g2_o21ai_1 _12435_ (.B1(_05709_),
    .Y(_00978_),
    .A1(_01183_),
    .A2(net2842));
 sg13g2_o21ai_1 _12436_ (.B1(_05703_),
    .Y(_05710_),
    .A1(\u_toplayer.u_layer1.u_neuron.acc[6] ),
    .A2(_05693_));
 sg13g2_o21ai_1 _12437_ (.B1(_05710_),
    .Y(_00979_),
    .A1(_01184_),
    .A2(net2842));
 sg13g2_nor2_1 _12438_ (.A(net3033),
    .B(net969),
    .Y(_05711_));
 sg13g2_a21oi_1 _12439_ (.A1(_01166_),
    .A2(net2842),
    .Y(_00980_),
    .B1(net970));
 sg13g2_nor2_1 _12440_ (.A(\u_toplayer.done_layer1 ),
    .B(_05231_),
    .Y(_05712_));
 sg13g2_nor2_2 _12441_ (.A(_05232_),
    .B(_05712_),
    .Y(_05713_));
 sg13g2_o21ai_1 _12442_ (.B1(\u_toplayer.u_layer1.statel1[0] ),
    .Y(_05714_),
    .A1(_05232_),
    .A2(_05712_));
 sg13g2_xnor2_1 _12443_ (.Y(_00981_),
    .A(net987),
    .B(_05713_));
 sg13g2_nor2_1 _12444_ (.A(_05227_),
    .B(_05713_),
    .Y(_05715_));
 sg13g2_xnor2_1 _12445_ (.Y(_00982_),
    .A(net921),
    .B(_05714_));
 sg13g2_nor2_1 _12446_ (.A(net994),
    .B(_05715_),
    .Y(_05716_));
 sg13g2_and2_1 _12447_ (.A(net994),
    .B(_05715_),
    .X(_05717_));
 sg13g2_nor3_1 _12448_ (.A(net2818),
    .B(_05716_),
    .C(_05717_),
    .Y(_00983_));
 sg13g2_xor2_1 _12449_ (.B(_05717_),
    .A(net960),
    .X(_00984_));
 sg13g2_nand3_1 _12450_ (.B(net960),
    .C(_05717_),
    .A(net1103),
    .Y(_05718_));
 sg13g2_a21o_1 _12451_ (.A2(_05717_),
    .A1(net960),
    .B1(net1103),
    .X(_05719_));
 sg13g2_and2_1 _12452_ (.A(_05718_),
    .B(_05719_),
    .X(_00985_));
 sg13g2_nand4_1 _12453_ (.B(\u_toplayer.u_layer1.statel1[4] ),
    .C(net960),
    .A(net877),
    .Y(_05720_),
    .D(net994));
 sg13g2_nor3_1 _12454_ (.A(_05227_),
    .B(_05713_),
    .C(_05720_),
    .Y(_05721_));
 sg13g2_xnor2_1 _12455_ (.Y(_00986_),
    .A(net877),
    .B(_05718_));
 sg13g2_and2_1 _12456_ (.A(\u_toplayer.u_layer1.statel1[6] ),
    .B(_05721_),
    .X(_05722_));
 sg13g2_xnor2_1 _12457_ (.Y(_00987_),
    .A(_01027_),
    .B(_05721_));
 sg13g2_xnor2_1 _12458_ (.Y(_00988_),
    .A(_01028_),
    .B(_05722_));
 sg13g2_nand2_1 _12459_ (.Y(_05723_),
    .A(net625),
    .B(_05713_));
 sg13g2_nand4_1 _12460_ (.B(\u_toplayer.u_layer1.statel1[0] ),
    .C(\u_toplayer.u_layer1.statel1[6] ),
    .A(\u_toplayer.u_layer1.statel1[1] ),
    .Y(_05724_),
    .D(\u_toplayer.u_layer1.statel1[7] ));
 sg13g2_o21ai_1 _12461_ (.B1(_00029_),
    .Y(_05725_),
    .A1(_05720_),
    .A2(_05724_));
 sg13g2_nand2b_1 _12462_ (.Y(_05726_),
    .B(_05725_),
    .A_N(_05231_));
 sg13g2_o21ai_1 _12463_ (.B1(_05723_),
    .Y(_00989_),
    .A1(_05713_),
    .A2(_05726_));
 sg13g2_nand2_1 _12464_ (.Y(_05727_),
    .A(\u_toplayer.u_layer1.u_neuron.acc[0] ),
    .B(net825));
 sg13g2_a21oi_1 _12465_ (.A1(_01158_),
    .A2(_01174_),
    .Y(_05728_),
    .B1(net3230));
 sg13g2_nand2_1 _12466_ (.Y(_05729_),
    .A(\u_toplayer.u_layer1.u_neuron.acc[0] ),
    .B(\u_toplayer.u_layer1.u_neuron.b[0] ));
 sg13g2_xor2_1 _12467_ (.B(net992),
    .A(\u_toplayer.u_layer1.u_neuron.acc[0] ),
    .X(_05730_));
 sg13g2_a221oi_1 _12468_ (.B2(net2855),
    .C1(net2832),
    .B1(_05730_),
    .A1(_05727_),
    .Y(_05731_),
    .A2(_05728_));
 sg13g2_a21oi_1 _12469_ (.A1(_01158_),
    .A2(net2832),
    .Y(_00990_),
    .B1(_05731_));
 sg13g2_nand2_1 _12470_ (.Y(_05732_),
    .A(\u_toplayer.u_layer1.u_neuron.acc[1] ),
    .B(\u_toplayer.u_layer1.u_neuron.mult[1] ));
 sg13g2_xnor2_1 _12471_ (.Y(_05733_),
    .A(\u_toplayer.u_layer1.u_neuron.acc[1] ),
    .B(\u_toplayer.u_layer1.u_neuron.mult[1] ));
 sg13g2_a21oi_1 _12472_ (.A1(_05727_),
    .A2(_05733_),
    .Y(_05734_),
    .B1(net3230));
 sg13g2_o21ai_1 _12473_ (.B1(_05734_),
    .Y(_05735_),
    .A1(_05727_),
    .A2(_05733_));
 sg13g2_nand2_1 _12474_ (.Y(_05736_),
    .A(\u_toplayer.u_layer1.u_neuron.acc[1] ),
    .B(\u_toplayer.u_layer1.u_neuron.b[1] ));
 sg13g2_xnor2_1 _12475_ (.Y(_05737_),
    .A(\u_toplayer.u_layer1.u_neuron.acc[1] ),
    .B(\u_toplayer.u_layer1.u_neuron.b[1] ));
 sg13g2_xnor2_1 _12476_ (.Y(_05738_),
    .A(_05729_),
    .B(_05737_));
 sg13g2_o21ai_1 _12477_ (.B1(_05735_),
    .Y(_05739_),
    .A1(net2853),
    .A2(_05738_));
 sg13g2_mux2_1 _12478_ (.A0(_05739_),
    .A1(net1133),
    .S(net2837),
    .X(_00991_));
 sg13g2_nand2_1 _12479_ (.Y(_05740_),
    .A(\u_toplayer.u_layer1.u_neuron.acc[2] ),
    .B(\u_toplayer.u_layer1.u_neuron.mult[2] ));
 sg13g2_inv_1 _12480_ (.Y(_05741_),
    .A(_05740_));
 sg13g2_or2_1 _12481_ (.X(_05742_),
    .B(\u_toplayer.u_layer1.u_neuron.mult[2] ),
    .A(\u_toplayer.u_layer1.u_neuron.acc[2] ));
 sg13g2_nand2_1 _12482_ (.Y(_05743_),
    .A(_05740_),
    .B(_05742_));
 sg13g2_o21ai_1 _12483_ (.B1(_05732_),
    .Y(_05744_),
    .A1(_05727_),
    .A2(_05733_));
 sg13g2_xnor2_1 _12484_ (.Y(_05745_),
    .A(_05743_),
    .B(_05744_));
 sg13g2_nand2_1 _12485_ (.Y(_05746_),
    .A(net3023),
    .B(_05745_));
 sg13g2_and2_1 _12486_ (.A(\u_toplayer.u_layer1.u_neuron.acc[2] ),
    .B(\u_toplayer.u_layer1.u_neuron.b[2] ),
    .X(_05747_));
 sg13g2_xor2_1 _12487_ (.B(\u_toplayer.u_layer1.u_neuron.b[2] ),
    .A(\u_toplayer.u_layer1.u_neuron.acc[2] ),
    .X(_05748_));
 sg13g2_o21ai_1 _12488_ (.B1(_05736_),
    .Y(_05749_),
    .A1(_05729_),
    .A2(_05737_));
 sg13g2_o21ai_1 _12489_ (.B1(net2855),
    .Y(_05750_),
    .A1(_05748_),
    .A2(_05749_));
 sg13g2_a21oi_1 _12490_ (.A1(_05748_),
    .A2(_05749_),
    .Y(_05751_),
    .B1(_05750_));
 sg13g2_nor2_1 _12491_ (.A(net2830),
    .B(_05751_),
    .Y(_05752_));
 sg13g2_a22oi_1 _12492_ (.Y(_00992_),
    .B1(_05746_),
    .B2(_05752_),
    .A2(net2830),
    .A1(_01157_));
 sg13g2_nand2_1 _12493_ (.Y(_05753_),
    .A(\u_toplayer.u_layer1.u_neuron.acc[3] ),
    .B(\u_toplayer.u_layer1.u_neuron.mult[3] ));
 sg13g2_xnor2_1 _12494_ (.Y(_05754_),
    .A(\u_toplayer.u_layer1.u_neuron.acc[3] ),
    .B(\u_toplayer.u_layer1.u_neuron.mult[3] ));
 sg13g2_a21oi_1 _12495_ (.A1(_05742_),
    .A2(_05744_),
    .Y(_05755_),
    .B1(_05741_));
 sg13g2_xor2_1 _12496_ (.B(_05755_),
    .A(_05754_),
    .X(_05756_));
 sg13g2_nand2_1 _12497_ (.Y(_05757_),
    .A(\u_toplayer.u_layer1.u_neuron.acc[3] ),
    .B(\u_toplayer.u_layer1.u_neuron.b[3] ));
 sg13g2_xnor2_1 _12498_ (.Y(_05758_),
    .A(\u_toplayer.u_layer1.u_neuron.acc[3] ),
    .B(\u_toplayer.u_layer1.u_neuron.b[3] ));
 sg13g2_a21oi_1 _12499_ (.A1(_05748_),
    .A2(_05749_),
    .Y(_05759_),
    .B1(_05747_));
 sg13g2_a21oi_1 _12500_ (.A1(_05758_),
    .A2(_05759_),
    .Y(_05760_),
    .B1(net2853));
 sg13g2_o21ai_1 _12501_ (.B1(_05760_),
    .Y(_05761_),
    .A1(_05758_),
    .A2(_05759_));
 sg13g2_a21oi_1 _12502_ (.A1(net3023),
    .A2(_05756_),
    .Y(_05762_),
    .B1(net2830));
 sg13g2_a22oi_1 _12503_ (.Y(_00993_),
    .B1(_05761_),
    .B2(_05762_),
    .A2(net2830),
    .A1(_01156_));
 sg13g2_and2_1 _12504_ (.A(\u_toplayer.u_layer1.u_neuron.acc[4] ),
    .B(\u_toplayer.u_layer1.u_neuron.mult[4] ),
    .X(_05763_));
 sg13g2_xor2_1 _12505_ (.B(\u_toplayer.u_layer1.u_neuron.mult[4] ),
    .A(\u_toplayer.u_layer1.u_neuron.acc[4] ),
    .X(_05764_));
 sg13g2_o21ai_1 _12506_ (.B1(_05753_),
    .Y(_05765_),
    .A1(_05754_),
    .A2(_05755_));
 sg13g2_and2_1 _12507_ (.A(_05764_),
    .B(_05765_),
    .X(_05766_));
 sg13g2_xor2_1 _12508_ (.B(_05765_),
    .A(_05764_),
    .X(_05767_));
 sg13g2_a21oi_1 _12509_ (.A1(net3023),
    .A2(_05767_),
    .Y(_05768_),
    .B1(net2830));
 sg13g2_and2_1 _12510_ (.A(\u_toplayer.u_layer1.u_neuron.acc[4] ),
    .B(\u_toplayer.u_layer1.u_neuron.b[4] ),
    .X(_05769_));
 sg13g2_xor2_1 _12511_ (.B(\u_toplayer.u_layer1.u_neuron.b[4] ),
    .A(\u_toplayer.u_layer1.u_neuron.acc[4] ),
    .X(_05770_));
 sg13g2_o21ai_1 _12512_ (.B1(_05757_),
    .Y(_05771_),
    .A1(_05758_),
    .A2(_05759_));
 sg13g2_o21ai_1 _12513_ (.B1(net2855),
    .Y(_05772_),
    .A1(_05770_),
    .A2(_05771_));
 sg13g2_a21o_1 _12514_ (.A2(_05771_),
    .A1(_05770_),
    .B1(_05772_),
    .X(_05773_));
 sg13g2_a22oi_1 _12515_ (.Y(_00994_),
    .B1(_05768_),
    .B2(_05773_),
    .A2(net2830),
    .A1(_01155_));
 sg13g2_nor2_1 _12516_ (.A(_05763_),
    .B(_05766_),
    .Y(_05774_));
 sg13g2_nor2_1 _12517_ (.A(net3030),
    .B(\u_toplayer.u_layer1.u_neuron.mult[5] ),
    .Y(_05775_));
 sg13g2_xor2_1 _12518_ (.B(\u_toplayer.u_layer1.u_neuron.mult[5] ),
    .A(net3030),
    .X(_05776_));
 sg13g2_xnor2_1 _12519_ (.Y(_05777_),
    .A(_05774_),
    .B(_05776_));
 sg13g2_a21oi_1 _12520_ (.A1(_05770_),
    .A2(_05771_),
    .Y(_05778_),
    .B1(_05769_));
 sg13g2_nor2_1 _12521_ (.A(net3030),
    .B(\u_toplayer.u_layer1.u_neuron.b[5] ),
    .Y(_05779_));
 sg13g2_xnor2_1 _12522_ (.Y(_05780_),
    .A(net3030),
    .B(net1019));
 sg13g2_a21oi_1 _12523_ (.A1(_05778_),
    .A2(_05780_),
    .Y(_05781_),
    .B1(net2853));
 sg13g2_o21ai_1 _12524_ (.B1(_05781_),
    .Y(_05782_),
    .A1(_05778_),
    .A2(_05780_));
 sg13g2_a21oi_1 _12525_ (.A1(net3023),
    .A2(_05777_),
    .Y(_05783_),
    .B1(net2830));
 sg13g2_a22oi_1 _12526_ (.Y(_00995_),
    .B1(_05782_),
    .B2(_05783_),
    .A2(net2830),
    .A1(_01154_));
 sg13g2_and2_1 _12527_ (.A(\u_toplayer.u_layer1.u_neuron.acc[6] ),
    .B(\u_toplayer.u_layer1.u_neuron.b[6] ),
    .X(_05784_));
 sg13g2_xnor2_1 _12528_ (.Y(_05785_),
    .A(\u_toplayer.u_layer1.u_neuron.acc[6] ),
    .B(\u_toplayer.u_layer1.u_neuron.b[6] ));
 sg13g2_a221oi_1 _12529_ (.B2(_05771_),
    .C1(_05769_),
    .B1(_05770_),
    .A1(net3030),
    .Y(_05786_),
    .A2(\u_toplayer.u_layer1.u_neuron.b[5] ));
 sg13g2_o21ai_1 _12530_ (.B1(_05785_),
    .Y(_05787_),
    .A1(_05779_),
    .A2(_05786_));
 sg13g2_nor3_2 _12531_ (.A(_05779_),
    .B(_05785_),
    .C(_05786_),
    .Y(_05788_));
 sg13g2_nor2_1 _12532_ (.A(net2853),
    .B(_05788_),
    .Y(_05789_));
 sg13g2_nand2_1 _12533_ (.Y(_05790_),
    .A(\u_toplayer.u_layer1.u_neuron.acc[6] ),
    .B(\u_toplayer.u_layer1.u_neuron.mult[6] ));
 sg13g2_xnor2_1 _12534_ (.Y(_05791_),
    .A(\u_toplayer.u_layer1.u_neuron.acc[6] ),
    .B(net945));
 sg13g2_a221oi_1 _12535_ (.B2(_05765_),
    .C1(_05763_),
    .B1(_05764_),
    .A1(net3030),
    .Y(_05792_),
    .A2(\u_toplayer.u_layer1.u_neuron.mult[5] ));
 sg13g2_or3_1 _12536_ (.A(_05775_),
    .B(_05791_),
    .C(_05792_),
    .X(_05793_));
 sg13g2_o21ai_1 _12537_ (.B1(_05791_),
    .Y(_05794_),
    .A1(_05775_),
    .A2(_05792_));
 sg13g2_nand3_1 _12538_ (.B(_05793_),
    .C(_05794_),
    .A(net3023),
    .Y(_05795_));
 sg13g2_a21oi_1 _12539_ (.A1(_05787_),
    .A2(_05789_),
    .Y(_05796_),
    .B1(net2831));
 sg13g2_a22oi_1 _12540_ (.Y(_00996_),
    .B1(_05795_),
    .B2(_05796_),
    .A2(net2831),
    .A1(_01153_));
 sg13g2_nand2_1 _12541_ (.Y(_05797_),
    .A(\u_toplayer.u_layer1.u_neuron.acc[7] ),
    .B(net3048));
 sg13g2_xnor2_1 _12542_ (.Y(_05798_),
    .A(\u_toplayer.u_layer1.u_neuron.acc[7] ),
    .B(net3049));
 sg13g2_inv_1 _12543_ (.Y(_05799_),
    .A(_05798_));
 sg13g2_nor3_1 _12544_ (.A(_05784_),
    .B(_05788_),
    .C(_05799_),
    .Y(_05800_));
 sg13g2_o21ai_1 _12545_ (.B1(_05799_),
    .Y(_05801_),
    .A1(_05784_),
    .A2(_05788_));
 sg13g2_nand3b_1 _12546_ (.B(_05801_),
    .C(net2855),
    .Y(_05802_),
    .A_N(_05800_));
 sg13g2_nand2_1 _12547_ (.Y(_05803_),
    .A(\u_toplayer.u_layer1.u_neuron.acc[7] ),
    .B(\u_toplayer.u_layer1.u_neuron.mult[7] ));
 sg13g2_inv_1 _12548_ (.Y(_05804_),
    .A(_05803_));
 sg13g2_xnor2_1 _12549_ (.Y(_05805_),
    .A(\u_toplayer.u_layer1.u_neuron.acc[7] ),
    .B(\u_toplayer.u_layer1.u_neuron.mult[7] ));
 sg13g2_a21oi_1 _12550_ (.A1(_05790_),
    .A2(_05793_),
    .Y(_05806_),
    .B1(_05805_));
 sg13g2_nand3_1 _12551_ (.B(_05793_),
    .C(_05805_),
    .A(_05790_),
    .Y(_05807_));
 sg13g2_nand2b_1 _12552_ (.Y(_05808_),
    .B(_05807_),
    .A_N(_05806_));
 sg13g2_nor2_1 _12553_ (.A(net3230),
    .B(_05808_),
    .Y(_05809_));
 sg13g2_nor2_1 _12554_ (.A(net2831),
    .B(_05809_),
    .Y(_05810_));
 sg13g2_a22oi_1 _12555_ (.Y(_00997_),
    .B1(_05802_),
    .B2(_05810_),
    .A2(net2831),
    .A1(_01152_));
 sg13g2_or2_1 _12556_ (.X(_05811_),
    .B(_05806_),
    .A(_05804_));
 sg13g2_and2_1 _12557_ (.A(\u_toplayer.u_layer1.u_neuron.acc[8] ),
    .B(\u_toplayer.u_layer1.u_neuron.mult[8] ),
    .X(_05812_));
 sg13g2_xor2_1 _12558_ (.B(\u_toplayer.u_layer1.u_neuron.mult[8] ),
    .A(\u_toplayer.u_layer1.u_neuron.acc[8] ),
    .X(_05813_));
 sg13g2_xor2_1 _12559_ (.B(_05813_),
    .A(_05811_),
    .X(_05814_));
 sg13g2_nand2_1 _12560_ (.Y(_05815_),
    .A(\u_toplayer.u_layer1.u_neuron.acc[8] ),
    .B(net3048));
 sg13g2_xnor2_1 _12561_ (.Y(_05816_),
    .A(\u_toplayer.u_layer1.u_neuron.acc[8] ),
    .B(net3048));
 sg13g2_a21o_1 _12562_ (.A2(_05801_),
    .A1(_05797_),
    .B1(_05816_),
    .X(_05817_));
 sg13g2_nand3_1 _12563_ (.B(_05801_),
    .C(_05816_),
    .A(_05797_),
    .Y(_05818_));
 sg13g2_and2_1 _12564_ (.A(net2855),
    .B(_05818_),
    .X(_05819_));
 sg13g2_a221oi_1 _12565_ (.B2(_05819_),
    .C1(net2834),
    .B1(_05817_),
    .A1(net3021),
    .Y(_05820_),
    .A2(_05814_));
 sg13g2_a21oi_1 _12566_ (.A1(_01165_),
    .A2(net2834),
    .Y(_00998_),
    .B1(_05820_));
 sg13g2_nor2_1 _12567_ (.A(\u_toplayer.u_layer1.u_neuron.acc[9] ),
    .B(\u_toplayer.u_layer1.u_neuron.mult[9] ),
    .Y(_05821_));
 sg13g2_nand2_1 _12568_ (.Y(_05822_),
    .A(\u_toplayer.u_layer1.u_neuron.acc[9] ),
    .B(\u_toplayer.u_layer1.u_neuron.mult[9] ));
 sg13g2_nor2b_1 _12569_ (.A(_05821_),
    .B_N(_05822_),
    .Y(_05823_));
 sg13g2_a21oi_1 _12570_ (.A1(_05811_),
    .A2(_05813_),
    .Y(_05824_),
    .B1(_05812_));
 sg13g2_xnor2_1 _12571_ (.Y(_05825_),
    .A(_05823_),
    .B(_05824_));
 sg13g2_xnor2_1 _12572_ (.Y(_05826_),
    .A(\u_toplayer.u_layer1.u_neuron.acc[9] ),
    .B(net3048));
 sg13g2_and2_1 _12573_ (.A(_05815_),
    .B(_05817_),
    .X(_05827_));
 sg13g2_a21oi_1 _12574_ (.A1(_05826_),
    .A2(_05827_),
    .Y(_05828_),
    .B1(net2854));
 sg13g2_o21ai_1 _12575_ (.B1(_05828_),
    .Y(_05829_),
    .A1(_05826_),
    .A2(_05827_));
 sg13g2_a21oi_1 _12576_ (.A1(net3023),
    .A2(_05825_),
    .Y(_05830_),
    .B1(net2832));
 sg13g2_a22oi_1 _12577_ (.Y(_00999_),
    .B1(_05829_),
    .B2(_05830_),
    .A2(net2834),
    .A1(_01164_));
 sg13g2_and2_1 _12578_ (.A(net3029),
    .B(\u_toplayer.u_layer1.u_neuron.mult[10] ),
    .X(_05831_));
 sg13g2_xor2_1 _12579_ (.B(\u_toplayer.u_layer1.u_neuron.mult[10] ),
    .A(net3029),
    .X(_05832_));
 sg13g2_and2_1 _12580_ (.A(_05813_),
    .B(_05823_),
    .X(_05833_));
 sg13g2_o21ai_1 _12581_ (.B1(_05833_),
    .Y(_05834_),
    .A1(_05804_),
    .A2(_05806_));
 sg13g2_nand2b_1 _12582_ (.Y(_05835_),
    .B(_05812_),
    .A_N(_05821_));
 sg13g2_nand3_1 _12583_ (.B(_05834_),
    .C(_05835_),
    .A(_05822_),
    .Y(_05836_));
 sg13g2_xor2_1 _12584_ (.B(_05836_),
    .A(_05832_),
    .X(_05837_));
 sg13g2_nand2_1 _12585_ (.Y(_05838_),
    .A(net3029),
    .B(net3049));
 sg13g2_xor2_1 _12586_ (.B(net3049),
    .A(net3029),
    .X(_05839_));
 sg13g2_xnor2_1 _12587_ (.Y(_05840_),
    .A(net3029),
    .B(net3049));
 sg13g2_o21ai_1 _12588_ (.B1(net3048),
    .Y(_05841_),
    .A1(\u_toplayer.u_layer1.u_neuron.acc[9] ),
    .A2(\u_toplayer.u_layer1.u_neuron.acc[8] ));
 sg13g2_a22oi_1 _12589_ (.Y(_05842_),
    .B1(_05817_),
    .B2(_05841_),
    .A2(_01176_),
    .A1(_01164_));
 sg13g2_nand2_1 _12590_ (.Y(_05843_),
    .A(_05839_),
    .B(_05842_));
 sg13g2_o21ai_1 _12591_ (.B1(net2855),
    .Y(_05844_),
    .A1(_05839_),
    .A2(_05842_));
 sg13g2_nand2b_1 _12592_ (.Y(_05845_),
    .B(_05843_),
    .A_N(_05844_));
 sg13g2_a21oi_1 _12593_ (.A1(net3023),
    .A2(_05837_),
    .Y(_05846_),
    .B1(net2832));
 sg13g2_a22oi_1 _12594_ (.Y(_01000_),
    .B1(_05845_),
    .B2(_05846_),
    .A2(net2833),
    .A1(_01162_));
 sg13g2_nor2_1 _12595_ (.A(\u_toplayer.u_layer1.u_neuron.acc[11] ),
    .B(\u_toplayer.u_layer1.u_neuron.mult[11] ),
    .Y(_05847_));
 sg13g2_xor2_1 _12596_ (.B(\u_toplayer.u_layer1.u_neuron.mult[11] ),
    .A(\u_toplayer.u_layer1.u_neuron.acc[11] ),
    .X(_05848_));
 sg13g2_a21oi_1 _12597_ (.A1(_05832_),
    .A2(_05836_),
    .Y(_05849_),
    .B1(_05831_));
 sg13g2_xnor2_1 _12598_ (.Y(_05850_),
    .A(_05848_),
    .B(_05849_));
 sg13g2_xnor2_1 _12599_ (.Y(_05851_),
    .A(\u_toplayer.u_layer1.u_neuron.acc[11] ),
    .B(net3049));
 sg13g2_a21oi_1 _12600_ (.A1(_05838_),
    .A2(_05843_),
    .Y(_05852_),
    .B1(_05851_));
 sg13g2_nand3_1 _12601_ (.B(_05843_),
    .C(_05851_),
    .A(_05838_),
    .Y(_05853_));
 sg13g2_nor2_1 _12602_ (.A(net2853),
    .B(_05852_),
    .Y(_05854_));
 sg13g2_a221oi_1 _12603_ (.B2(_05854_),
    .C1(net2832),
    .B1(_05853_),
    .A1(net3023),
    .Y(_05855_),
    .A2(_05850_));
 sg13g2_a21oi_1 _12604_ (.A1(_01163_),
    .A2(net2832),
    .Y(_01001_),
    .B1(_05855_));
 sg13g2_a21oi_1 _12605_ (.A1(\u_toplayer.u_layer1.u_neuron.acc[11] ),
    .A2(\u_toplayer.u_layer1.u_neuron.mult[11] ),
    .Y(_05856_),
    .B1(_05831_));
 sg13g2_nor2_1 _12606_ (.A(_05847_),
    .B(_05856_),
    .Y(_05857_));
 sg13g2_inv_1 _12607_ (.Y(_05858_),
    .A(_05857_));
 sg13g2_and2_1 _12608_ (.A(_05832_),
    .B(_05848_),
    .X(_05859_));
 sg13g2_inv_1 _12609_ (.Y(_05860_),
    .A(_05859_));
 sg13g2_and3_1 _12610_ (.X(_05861_),
    .A(_05822_),
    .B(_05835_),
    .C(_05858_));
 sg13g2_a21oi_1 _12611_ (.A1(_05836_),
    .A2(_05859_),
    .Y(_05862_),
    .B1(_05857_));
 sg13g2_nand2_1 _12612_ (.Y(_05863_),
    .A(net3028),
    .B(\u_toplayer.u_layer1.u_neuron.mult[12] ));
 sg13g2_xor2_1 _12613_ (.B(\u_toplayer.u_layer1.u_neuron.mult[12] ),
    .A(net3028),
    .X(_05864_));
 sg13g2_nand2b_1 _12614_ (.Y(_05865_),
    .B(_05864_),
    .A_N(_05862_));
 sg13g2_xnor2_1 _12615_ (.Y(_05866_),
    .A(_05862_),
    .B(_05864_));
 sg13g2_and2_1 _12616_ (.A(net3028),
    .B(net3048),
    .X(_05867_));
 sg13g2_xor2_1 _12617_ (.B(net3048),
    .A(net3028),
    .X(_05868_));
 sg13g2_inv_1 _12618_ (.Y(_05869_),
    .A(_05868_));
 sg13g2_or4_1 _12619_ (.A(_05816_),
    .B(_05826_),
    .C(_05840_),
    .D(_05851_),
    .X(_05870_));
 sg13g2_a21oi_1 _12620_ (.A1(_05797_),
    .A2(_05801_),
    .Y(_05871_),
    .B1(_05870_));
 sg13g2_o21ai_1 _12621_ (.B1(net3048),
    .Y(_05872_),
    .A1(net3029),
    .A2(\u_toplayer.u_layer1.u_neuron.acc[11] ));
 sg13g2_and2_1 _12622_ (.A(_05841_),
    .B(_05872_),
    .X(_05873_));
 sg13g2_nand2b_1 _12623_ (.Y(_05874_),
    .B(_05873_),
    .A_N(_05871_));
 sg13g2_o21ai_1 _12624_ (.B1(net2856),
    .Y(_05875_),
    .A1(_05868_),
    .A2(_05874_));
 sg13g2_a21oi_1 _12625_ (.A1(_05868_),
    .A2(_05874_),
    .Y(_05876_),
    .B1(_05875_));
 sg13g2_a21oi_1 _12626_ (.A1(net3021),
    .A2(_05866_),
    .Y(_05877_),
    .B1(_05876_));
 sg13g2_nand2_1 _12627_ (.Y(_05878_),
    .A(net3028),
    .B(net2833));
 sg13g2_o21ai_1 _12628_ (.B1(_05878_),
    .Y(_01002_),
    .A1(net2833),
    .A2(_05877_));
 sg13g2_nor2_1 _12629_ (.A(\u_toplayer.u_layer1.u_neuron.acc[13] ),
    .B(\u_toplayer.u_layer1.u_neuron.mult[13] ),
    .Y(_05879_));
 sg13g2_xnor2_1 _12630_ (.Y(_05880_),
    .A(net3027),
    .B(\u_toplayer.u_layer1.u_neuron.mult[13] ));
 sg13g2_inv_1 _12631_ (.Y(_05881_),
    .A(_05880_));
 sg13g2_nand2_1 _12632_ (.Y(_05882_),
    .A(_05863_),
    .B(_05865_));
 sg13g2_xnor2_1 _12633_ (.Y(_05883_),
    .A(_05881_),
    .B(_05882_));
 sg13g2_nor2_1 _12634_ (.A(net3230),
    .B(_05883_),
    .Y(_05884_));
 sg13g2_xnor2_1 _12635_ (.Y(_05885_),
    .A(net3027),
    .B(net3052));
 sg13g2_a21oi_1 _12636_ (.A1(_05868_),
    .A2(_05874_),
    .Y(_05886_),
    .B1(_05867_));
 sg13g2_o21ai_1 _12637_ (.B1(net2856),
    .Y(_05887_),
    .A1(_05885_),
    .A2(_05886_));
 sg13g2_a21oi_1 _12638_ (.A1(_05885_),
    .A2(_05886_),
    .Y(_05888_),
    .B1(_05887_));
 sg13g2_nor3_1 _12639_ (.A(net2834),
    .B(_05884_),
    .C(_05888_),
    .Y(_05889_));
 sg13g2_a21oi_1 _12640_ (.A1(_01161_),
    .A2(net2833),
    .Y(_01003_),
    .B1(_05889_));
 sg13g2_nand2_1 _12641_ (.Y(_05890_),
    .A(\u_toplayer.u_layer1.u_neuron.acc[14] ),
    .B(\u_toplayer.u_layer1.u_neuron.mult[14] ));
 sg13g2_xnor2_1 _12642_ (.Y(_05891_),
    .A(\u_toplayer.u_layer1.u_neuron.acc[14] ),
    .B(\u_toplayer.u_layer1.u_neuron.mult[14] ));
 sg13g2_a22oi_1 _12643_ (.Y(_05892_),
    .B1(\u_toplayer.u_layer1.u_neuron.mult[13] ),
    .B2(net3027),
    .A2(\u_toplayer.u_layer1.u_neuron.mult[12] ),
    .A1(net3028));
 sg13g2_a21oi_1 _12644_ (.A1(_05865_),
    .A2(_05892_),
    .Y(_05893_),
    .B1(_05879_));
 sg13g2_nand2b_1 _12645_ (.Y(_05894_),
    .B(_05893_),
    .A_N(_05891_));
 sg13g2_xnor2_1 _12646_ (.Y(_05895_),
    .A(_05891_),
    .B(_05893_));
 sg13g2_nand2_1 _12647_ (.Y(_05896_),
    .A(\u_toplayer.u_layer1.u_neuron.acc[14] ),
    .B(net3052));
 sg13g2_xnor2_1 _12648_ (.Y(_05897_),
    .A(\u_toplayer.u_layer1.u_neuron.acc[14] ),
    .B(net3052));
 sg13g2_o21ai_1 _12649_ (.B1(net3052),
    .Y(_05898_),
    .A1(net3028),
    .A2(net3027));
 sg13g2_o21ai_1 _12650_ (.B1(_05886_),
    .Y(_05899_),
    .A1(_01161_),
    .A2(_01176_));
 sg13g2_o21ai_1 _12651_ (.B1(_05899_),
    .Y(_05900_),
    .A1(net3027),
    .A2(net3052));
 sg13g2_or2_1 _12652_ (.X(_05901_),
    .B(_05900_),
    .A(_05897_));
 sg13g2_a21oi_1 _12653_ (.A1(_05897_),
    .A2(_05900_),
    .Y(_05902_),
    .B1(net2854));
 sg13g2_a221oi_1 _12654_ (.B2(_05902_),
    .C1(net2833),
    .B1(_05901_),
    .A1(net3021),
    .Y(_05903_),
    .A2(_05895_));
 sg13g2_a21oi_1 _12655_ (.A1(_01160_),
    .A2(net2833),
    .Y(_01004_),
    .B1(_05903_));
 sg13g2_nor2_1 _12656_ (.A(\u_toplayer.u_layer1.u_neuron.acc[15] ),
    .B(net3144),
    .Y(_05904_));
 sg13g2_nand2_1 _12657_ (.Y(_05905_),
    .A(\u_toplayer.u_layer1.u_neuron.acc[15] ),
    .B(net3144));
 sg13g2_nand2b_1 _12658_ (.Y(_05906_),
    .B(_05905_),
    .A_N(_05904_));
 sg13g2_and2_1 _12659_ (.A(_05890_),
    .B(_05894_),
    .X(_05907_));
 sg13g2_xor2_1 _12660_ (.B(_05907_),
    .A(_05906_),
    .X(_05908_));
 sg13g2_xnor2_1 _12661_ (.Y(_05909_),
    .A(\u_toplayer.u_layer1.u_neuron.acc[15] ),
    .B(net3052));
 sg13g2_nand3_1 _12662_ (.B(_05901_),
    .C(_05909_),
    .A(_05896_),
    .Y(_05910_));
 sg13g2_a21oi_1 _12663_ (.A1(_05896_),
    .A2(_05901_),
    .Y(_05911_),
    .B1(_05909_));
 sg13g2_nor2_1 _12664_ (.A(net2854),
    .B(_05911_),
    .Y(_05912_));
 sg13g2_a221oi_1 _12665_ (.B2(_05912_),
    .C1(net2833),
    .B1(_05910_),
    .A1(net3021),
    .Y(_05913_),
    .A2(_05908_));
 sg13g2_a21oi_1 _12666_ (.A1(_01159_),
    .A2(net2833),
    .Y(_01005_),
    .B1(_05913_));
 sg13g2_nor2_1 _12667_ (.A(_05891_),
    .B(_05906_),
    .Y(_05914_));
 sg13g2_nand3_1 _12668_ (.B(_05881_),
    .C(_05914_),
    .A(_05864_),
    .Y(_05915_));
 sg13g2_a221oi_1 _12669_ (.B2(_05834_),
    .C1(_05915_),
    .B1(_05861_),
    .A1(_05858_),
    .Y(_05916_),
    .A2(_05860_));
 sg13g2_nor4_1 _12670_ (.A(_05879_),
    .B(_05891_),
    .C(_05892_),
    .D(_05906_),
    .Y(_05917_));
 sg13g2_o21ai_1 _12671_ (.B1(_05905_),
    .Y(_05918_),
    .A1(_05890_),
    .A2(_05904_));
 sg13g2_or2_1 _12672_ (.X(_05919_),
    .B(_05918_),
    .A(_05917_));
 sg13g2_or2_1 _12673_ (.X(_05920_),
    .B(_05919_),
    .A(_05916_));
 sg13g2_and2_1 _12674_ (.A(net3026),
    .B(net3142),
    .X(_05921_));
 sg13g2_xor2_1 _12675_ (.B(net3143),
    .A(net3026),
    .X(_05922_));
 sg13g2_inv_1 _12676_ (.Y(_05923_),
    .A(_05922_));
 sg13g2_o21ai_1 _12677_ (.B1(net3022),
    .Y(_05924_),
    .A1(_05920_),
    .A2(_05922_));
 sg13g2_a21o_1 _12678_ (.A2(_05922_),
    .A1(_05920_),
    .B1(_05924_),
    .X(_05925_));
 sg13g2_nor4_1 _12679_ (.A(_05869_),
    .B(_05885_),
    .C(_05897_),
    .D(_05909_),
    .Y(_05926_));
 sg13g2_o21ai_1 _12680_ (.B1(net3052),
    .Y(_05927_),
    .A1(\u_toplayer.u_layer1.u_neuron.acc[15] ),
    .A2(\u_toplayer.u_layer1.u_neuron.acc[14] ));
 sg13g2_nand3_1 _12681_ (.B(_05898_),
    .C(_05927_),
    .A(_05873_),
    .Y(_05928_));
 sg13g2_a21oi_2 _12682_ (.B1(_05928_),
    .Y(_05929_),
    .A2(_05926_),
    .A1(_05871_));
 sg13g2_nand2_1 _12683_ (.Y(_05930_),
    .A(net3026),
    .B(net3051));
 sg13g2_xnor2_1 _12684_ (.Y(_05931_),
    .A(net3026),
    .B(net3051));
 sg13g2_or2_1 _12685_ (.X(_05932_),
    .B(_05931_),
    .A(_05929_));
 sg13g2_a21oi_1 _12686_ (.A1(_05929_),
    .A2(_05931_),
    .Y(_05933_),
    .B1(net2854));
 sg13g2_a21oi_1 _12687_ (.A1(_05932_),
    .A2(_05933_),
    .Y(_05934_),
    .B1(net2836));
 sg13g2_a22oi_1 _12688_ (.Y(_01006_),
    .B1(_05925_),
    .B2(_05934_),
    .A2(net2835),
    .A1(_01172_));
 sg13g2_xnor2_1 _12689_ (.Y(_05935_),
    .A(\u_toplayer.u_layer1.u_neuron.acc[17] ),
    .B(net3142));
 sg13g2_a21oi_1 _12690_ (.A1(_05920_),
    .A2(_05922_),
    .Y(_05936_),
    .B1(_05921_));
 sg13g2_xor2_1 _12691_ (.B(_05936_),
    .A(_05935_),
    .X(_05937_));
 sg13g2_xnor2_1 _12692_ (.Y(_05938_),
    .A(\u_toplayer.u_layer1.u_neuron.acc[17] ),
    .B(net3051));
 sg13g2_nand3_1 _12693_ (.B(_05932_),
    .C(_05938_),
    .A(_05930_),
    .Y(_05939_));
 sg13g2_a21oi_1 _12694_ (.A1(_05930_),
    .A2(_05932_),
    .Y(_05940_),
    .B1(_05938_));
 sg13g2_nor2_1 _12695_ (.A(net2854),
    .B(_05940_),
    .Y(_05941_));
 sg13g2_a221oi_1 _12696_ (.B2(_05941_),
    .C1(net2836),
    .B1(_05939_),
    .A1(net3022),
    .Y(_05942_),
    .A2(_05937_));
 sg13g2_a21oi_1 _12697_ (.A1(_01173_),
    .A2(net2836),
    .Y(_01007_),
    .B1(_05942_));
 sg13g2_xor2_1 _12698_ (.B(net3143),
    .A(\u_toplayer.u_layer1.u_neuron.acc[18] ),
    .X(_05943_));
 sg13g2_nor2_1 _12699_ (.A(_05923_),
    .B(_05935_),
    .Y(_05944_));
 sg13g2_o21ai_1 _12700_ (.B1(_05944_),
    .Y(_05945_),
    .A1(_05916_),
    .A2(_05919_));
 sg13g2_o21ai_1 _12701_ (.B1(net3143),
    .Y(_05946_),
    .A1(net3026),
    .A2(\u_toplayer.u_layer1.u_neuron.acc[17] ));
 sg13g2_nand2_1 _12702_ (.Y(_05947_),
    .A(_05945_),
    .B(_05946_));
 sg13g2_and2_1 _12703_ (.A(_05943_),
    .B(_05947_),
    .X(_05948_));
 sg13g2_o21ai_1 _12704_ (.B1(net3022),
    .Y(_05949_),
    .A1(_05943_),
    .A2(_05947_));
 sg13g2_xnor2_1 _12705_ (.Y(_05950_),
    .A(net3025),
    .B(net3051));
 sg13g2_or2_1 _12706_ (.X(_05951_),
    .B(_05938_),
    .A(_05932_));
 sg13g2_o21ai_1 _12707_ (.B1(net3051),
    .Y(_05952_),
    .A1(net3026),
    .A2(\u_toplayer.u_layer1.u_neuron.acc[17] ));
 sg13g2_a21o_1 _12708_ (.A2(_05952_),
    .A1(_05951_),
    .B1(_05950_),
    .X(_05953_));
 sg13g2_nand3_1 _12709_ (.B(_05951_),
    .C(_05952_),
    .A(_05950_),
    .Y(_05954_));
 sg13g2_nand3_1 _12710_ (.B(_05953_),
    .C(_05954_),
    .A(net2856),
    .Y(_05955_));
 sg13g2_o21ai_1 _12711_ (.B1(_05955_),
    .Y(_05956_),
    .A1(_05948_),
    .A2(_05949_));
 sg13g2_mux2_1 _12712_ (.A0(_05956_),
    .A1(net3025),
    .S(net2836),
    .X(_01008_));
 sg13g2_xor2_1 _12713_ (.B(net3143),
    .A(\u_toplayer.u_layer1.u_neuron.acc[19] ),
    .X(_05957_));
 sg13g2_a21oi_1 _12714_ (.A1(net3025),
    .A2(net3143),
    .Y(_05958_),
    .B1(_05948_));
 sg13g2_xnor2_1 _12715_ (.Y(_05959_),
    .A(_05957_),
    .B(_05958_));
 sg13g2_nand2_1 _12716_ (.Y(_05960_),
    .A(net3021),
    .B(_05959_));
 sg13g2_xor2_1 _12717_ (.B(net3051),
    .A(\u_toplayer.u_layer1.u_neuron.acc[19] ),
    .X(_05961_));
 sg13g2_o21ai_1 _12718_ (.B1(_05953_),
    .Y(_05962_),
    .A1(_01170_),
    .A2(_01176_));
 sg13g2_o21ai_1 _12719_ (.B1(net2856),
    .Y(_05963_),
    .A1(_05961_),
    .A2(_05962_));
 sg13g2_a21oi_1 _12720_ (.A1(_05961_),
    .A2(_05962_),
    .Y(_05964_),
    .B1(_05963_));
 sg13g2_nor2_1 _12721_ (.A(net2836),
    .B(_05964_),
    .Y(_05965_));
 sg13g2_a22oi_1 _12722_ (.Y(_01009_),
    .B1(_05960_),
    .B2(_05965_),
    .A2(net2836),
    .A1(_01171_));
 sg13g2_nand2_1 _12723_ (.Y(_05966_),
    .A(_05943_),
    .B(_05957_));
 sg13g2_o21ai_1 _12724_ (.B1(net3143),
    .Y(_05967_),
    .A1(net3025),
    .A2(\u_toplayer.u_layer1.u_neuron.acc[19] ));
 sg13g2_and2_1 _12725_ (.A(_05946_),
    .B(_05967_),
    .X(_05968_));
 sg13g2_o21ai_1 _12726_ (.B1(_05968_),
    .Y(_05969_),
    .A1(_05945_),
    .A2(_05966_));
 sg13g2_and2_1 _12727_ (.A(\u_toplayer.u_layer1.u_neuron.acc[20] ),
    .B(net3142),
    .X(_05970_));
 sg13g2_xor2_1 _12728_ (.B(net3142),
    .A(\u_toplayer.u_layer1.u_neuron.acc[20] ),
    .X(_05971_));
 sg13g2_and2_1 _12729_ (.A(_05969_),
    .B(_05971_),
    .X(_05972_));
 sg13g2_o21ai_1 _12730_ (.B1(net3022),
    .Y(_05973_),
    .A1(_05969_),
    .A2(_05971_));
 sg13g2_or2_1 _12731_ (.X(_05974_),
    .B(_05973_),
    .A(_05972_));
 sg13g2_xor2_1 _12732_ (.B(net3050),
    .A(\u_toplayer.u_layer1.u_neuron.acc[20] ),
    .X(_05975_));
 sg13g2_nand2b_1 _12733_ (.Y(_05976_),
    .B(_05961_),
    .A_N(_05950_));
 sg13g2_nor4_2 _12734_ (.A(_05929_),
    .B(_05931_),
    .C(_05938_),
    .Y(_05977_),
    .D(_05976_));
 sg13g2_o21ai_1 _12735_ (.B1(net3050),
    .Y(_05978_),
    .A1(net3025),
    .A2(\u_toplayer.u_layer1.u_neuron.acc[19] ));
 sg13g2_nand2_1 _12736_ (.Y(_05979_),
    .A(_05952_),
    .B(_05978_));
 sg13g2_o21ai_1 _12737_ (.B1(_05975_),
    .Y(_05980_),
    .A1(_05977_),
    .A2(_05979_));
 sg13g2_nor3_1 _12738_ (.A(_05975_),
    .B(_05977_),
    .C(_05979_),
    .Y(_05981_));
 sg13g2_nor2_1 _12739_ (.A(net2853),
    .B(_05981_),
    .Y(_05982_));
 sg13g2_a21oi_1 _12740_ (.A1(_05980_),
    .A2(_05982_),
    .Y(_05983_),
    .B1(net2835));
 sg13g2_a22oi_1 _12741_ (.Y(_01010_),
    .B1(_05974_),
    .B2(_05983_),
    .A2(net2835),
    .A1(_01169_));
 sg13g2_xor2_1 _12742_ (.B(net3142),
    .A(\u_toplayer.u_layer1.u_neuron.acc[21] ),
    .X(_05984_));
 sg13g2_nor3_1 _12743_ (.A(_05970_),
    .B(_05972_),
    .C(_05984_),
    .Y(_05985_));
 sg13g2_o21ai_1 _12744_ (.B1(_05984_),
    .Y(_05986_),
    .A1(_05970_),
    .A2(_05972_));
 sg13g2_nor2_1 _12745_ (.A(net3230),
    .B(_05985_),
    .Y(_05987_));
 sg13g2_xnor2_1 _12746_ (.Y(_05988_),
    .A(\u_toplayer.u_layer1.u_neuron.acc[21] ),
    .B(net3050));
 sg13g2_o21ai_1 _12747_ (.B1(_05980_),
    .Y(_05989_),
    .A1(_01169_),
    .A2(_01176_));
 sg13g2_xnor2_1 _12748_ (.Y(_05990_),
    .A(_05988_),
    .B(_05989_));
 sg13g2_a221oi_1 _12749_ (.B2(net2856),
    .C1(net2835),
    .B1(_05990_),
    .A1(_05986_),
    .Y(_05991_),
    .A2(_05987_));
 sg13g2_a21oi_1 _12750_ (.A1(_01168_),
    .A2(net2835),
    .Y(_01011_),
    .B1(_05991_));
 sg13g2_xnor2_1 _12751_ (.Y(_05992_),
    .A(\u_toplayer.u_layer1.u_neuron.acc[22] ),
    .B(net3142));
 sg13g2_nand3_1 _12752_ (.B(_05971_),
    .C(_05984_),
    .A(_05969_),
    .Y(_05993_));
 sg13g2_o21ai_1 _12753_ (.B1(net3142),
    .Y(_05994_),
    .A1(\u_toplayer.u_layer1.u_neuron.acc[21] ),
    .A2(\u_toplayer.u_layer1.u_neuron.acc[20] ));
 sg13g2_a21oi_1 _12754_ (.A1(_05993_),
    .A2(_05994_),
    .Y(_05995_),
    .B1(_05992_));
 sg13g2_and3_1 _12755_ (.X(_05996_),
    .A(_05992_),
    .B(_05993_),
    .C(_05994_));
 sg13g2_nor3_1 _12756_ (.A(net3230),
    .B(_05995_),
    .C(_05996_),
    .Y(_05997_));
 sg13g2_nand2_1 _12757_ (.Y(_05998_),
    .A(\u_toplayer.u_layer1.u_neuron.acc[22] ),
    .B(net3050));
 sg13g2_xor2_1 _12758_ (.B(net3050),
    .A(\u_toplayer.u_layer1.u_neuron.acc[22] ),
    .X(_05999_));
 sg13g2_o21ai_1 _12759_ (.B1(net3050),
    .Y(_06000_),
    .A1(\u_toplayer.u_layer1.u_neuron.acc[21] ),
    .A2(\u_toplayer.u_layer1.u_neuron.acc[20] ));
 sg13g2_o21ai_1 _12760_ (.B1(_06000_),
    .Y(_06001_),
    .A1(_05980_),
    .A2(_05988_));
 sg13g2_nand2_1 _12761_ (.Y(_06002_),
    .A(_05999_),
    .B(_06001_));
 sg13g2_o21ai_1 _12762_ (.B1(net2855),
    .Y(_06003_),
    .A1(_05999_),
    .A2(_06001_));
 sg13g2_nand2b_1 _12763_ (.Y(_06004_),
    .B(_06002_),
    .A_N(_06003_));
 sg13g2_nor2_1 _12764_ (.A(net2835),
    .B(_05997_),
    .Y(_06005_));
 sg13g2_a22oi_1 _12765_ (.Y(_01012_),
    .B1(_06004_),
    .B2(_06005_),
    .A2(net2835),
    .A1(_01167_));
 sg13g2_a21oi_1 _12766_ (.A1(\u_toplayer.u_layer1.u_neuron.acc[22] ),
    .A2(net3142),
    .Y(_06006_),
    .B1(_05995_));
 sg13g2_xor2_1 _12767_ (.B(net3144),
    .A(\u_toplayer.u_layer1.u_neuron.acc[23] ),
    .X(_06007_));
 sg13g2_xnor2_1 _12768_ (.Y(_06008_),
    .A(_06006_),
    .B(_06007_));
 sg13g2_xnor2_1 _12769_ (.Y(_06009_),
    .A(\u_toplayer.u_layer1.u_neuron.acc[23] ),
    .B(net3050));
 sg13g2_a21oi_1 _12770_ (.A1(_05998_),
    .A2(_06002_),
    .Y(_06010_),
    .B1(_06009_));
 sg13g2_nand3_1 _12771_ (.B(_06002_),
    .C(_06009_),
    .A(_05998_),
    .Y(_06011_));
 sg13g2_nor2_1 _12772_ (.A(net2853),
    .B(_06010_),
    .Y(_06012_));
 sg13g2_a221oi_1 _12773_ (.B2(_06012_),
    .C1(net2835),
    .B1(_06011_),
    .A1(net3022),
    .Y(_06013_),
    .A2(_06008_));
 sg13g2_a21oi_1 _12774_ (.A1(_01166_),
    .A2(net2834),
    .Y(_01013_),
    .B1(_06013_));
 sg13g2_nor3_1 _12775_ (.A(_01022_),
    .B(net124),
    .C(\u_toplayer.done_layer1 ),
    .Y(_01014_));
 sg13g2_a21o_1 _12776_ (.A2(net124),
    .A1(net812),
    .B1(net943),
    .X(_01015_));
 sg13g2_nor3_1 _12777_ (.A(_01023_),
    .B(net130),
    .C(\u_toplayer.done_layer2 ),
    .Y(_01016_));
 sg13g2_a21o_1 _12778_ (.A2(net130),
    .A1(net925),
    .B1(\u_toplayer.done_layer2 ),
    .X(_01017_));
 sg13g2_buf_1 _12779_ (.A(net120),
    .X(_00347_));
 sg13g2_buf_1 _12780_ (.A(net121),
    .X(_00346_));
 sg13g2_inv_1 _12782__3 (.Y(net22),
    .A(clknet_4_8_0_clk));
 sg13g2_inv_1 _12783__4 (.Y(net23),
    .A(clknet_4_8_0_clk));
 sg13g2_inv_1 _12784__5 (.Y(net24),
    .A(clknet_4_8_0_clk));
 sg13g2_inv_1 _12785__6 (.Y(net25),
    .A(clknet_4_8_0_clk));
 sg13g2_inv_1 _12786__7 (.Y(net26),
    .A(clknet_4_14_0_clk));
 sg13g2_inv_1 _12787__8 (.Y(net27),
    .A(clknet_4_11_0_clk));
 sg13g2_inv_1 _12788__9 (.Y(net28),
    .A(clknet_4_10_0_clk));
 sg13g2_inv_1 _12789__10 (.Y(net29),
    .A(clknet_4_10_0_clk));
 sg13g2_inv_1 _12790__11 (.Y(net30),
    .A(clknet_4_14_0_clk));
 sg13g2_inv_1 _12791__12 (.Y(net31),
    .A(clknet_4_15_0_clk));
 sg13g2_inv_1 _12792__13 (.Y(net32),
    .A(clknet_4_14_0_clk));
 sg13g2_inv_1 _12793__14 (.Y(net33),
    .A(clknet_4_13_0_clk));
 sg13g2_inv_1 _12794__15 (.Y(net34),
    .A(clknet_4_13_0_clk));
 sg13g2_inv_1 _12795__16 (.Y(net35),
    .A(clknet_4_9_0_clk));
 sg13g2_inv_1 _12796__17 (.Y(net36),
    .A(clknet_4_10_0_clk));
 sg13g2_inv_1 _12797__18 (.Y(net37),
    .A(clknet_4_11_0_clk));
 sg13g2_inv_1 _12798__19 (.Y(net38),
    .A(clknet_4_10_0_clk));
 sg13g2_inv_1 _12799__20 (.Y(net39),
    .A(clknet_4_15_0_clk));
 sg13g2_inv_1 _12800__21 (.Y(net40),
    .A(clknet_4_14_0_clk));
 sg13g2_inv_1 _12801__22 (.Y(net41),
    .A(clknet_4_13_0_clk));
 sg13g2_inv_1 _12802__23 (.Y(net42),
    .A(clknet_4_4_0_clk));
 sg13g2_inv_1 _12803__24 (.Y(net43),
    .A(clknet_4_0_0_clk));
 sg13g2_inv_1 _12804__25 (.Y(net44),
    .A(clknet_4_0_0_clk));
 sg13g2_inv_1 _12805__26 (.Y(net45),
    .A(clknet_4_0_0_clk));
 sg13g2_inv_1 _12806__27 (.Y(net46),
    .A(clknet_4_4_0_clk));
 sg13g2_inv_1 _12807__28 (.Y(net47),
    .A(clknet_4_5_0_clk));
 sg13g2_inv_1 _12808__29 (.Y(net48),
    .A(clknet_4_5_0_clk));
 sg13g2_inv_1 _12809__30 (.Y(net49),
    .A(clknet_4_6_0_clk));
 sg13g2_inv_1 _12810__31 (.Y(net50),
    .A(clknet_4_5_0_clk));
 sg13g2_inv_1 _12811__32 (.Y(net51),
    .A(clknet_4_4_0_clk));
 sg13g2_inv_1 _12812__33 (.Y(net52),
    .A(clknet_4_0_0_clk));
 sg13g2_inv_1 _12813__34 (.Y(net53),
    .A(clknet_4_0_0_clk));
 sg13g2_inv_1 _12814__35 (.Y(net54),
    .A(clknet_4_4_0_clk));
 sg13g2_inv_1 _12815__36 (.Y(net55),
    .A(clknet_4_5_0_clk));
 sg13g2_inv_1 _12816__37 (.Y(net56),
    .A(clknet_4_5_0_clk));
 sg13g2_inv_1 _12817__38 (.Y(net57),
    .A(clknet_4_4_0_clk));
 sg13g2_inv_1 _12818__39 (.Y(net58),
    .A(clknet_4_1_0_clk));
 sg13g2_inv_1 _12819__40 (.Y(net59),
    .A(clknet_4_1_0_clk));
 sg13g2_inv_1 _12820__41 (.Y(net60),
    .A(clknet_4_1_0_clk));
 sg13g2_inv_1 _12821__42 (.Y(net61),
    .A(clknet_4_0_0_clk));
 sg13g2_inv_1 _12822__43 (.Y(net62),
    .A(clknet_4_4_0_clk));
 sg13g2_inv_1 _12823__44 (.Y(net63),
    .A(clknet_4_6_0_clk));
 sg13g2_inv_1 _12824__45 (.Y(net64),
    .A(clknet_4_7_0_clk));
 sg13g2_inv_1 _12825__46 (.Y(net65),
    .A(clknet_4_12_0_clk));
 sg13g2_inv_1 _12826__47 (.Y(net66),
    .A(clknet_4_7_0_clk));
 sg13g2_inv_1 _12827__48 (.Y(net67),
    .A(clknet_4_1_0_clk));
 sg13g2_inv_1 _12828__49 (.Y(net68),
    .A(clknet_4_3_0_clk));
 sg13g2_inv_1 _12829__50 (.Y(net69),
    .A(clknet_4_1_0_clk));
 sg13g2_inv_1 _12830__51 (.Y(net70),
    .A(clknet_4_1_0_clk));
 sg13g2_inv_1 _12831__52 (.Y(net71),
    .A(clknet_4_6_0_clk));
 sg13g2_inv_1 _12832__53 (.Y(net72),
    .A(clknet_4_12_0_clk));
 sg13g2_inv_1 _12833__54 (.Y(net73),
    .A(clknet_4_12_0_clk));
 sg13g2_inv_1 _12834__55 (.Y(net74),
    .A(clknet_4_6_0_clk));
 sg13g2_inv_1 _12835__56 (.Y(net75),
    .A(clknet_4_9_0_clk));
 sg13g2_inv_1 _12836__57 (.Y(net76),
    .A(clknet_4_9_0_clk));
 sg13g2_inv_1 _12837__58 (.Y(net77),
    .A(clknet_4_3_0_clk));
 sg13g2_inv_1 _12838__59 (.Y(net78),
    .A(clknet_4_12_0_clk));
 sg13g2_inv_1 _12839__60 (.Y(net79),
    .A(clknet_4_5_0_clk));
 sg13g2_inv_1 _12840__61 (.Y(net80),
    .A(clknet_4_7_0_clk));
 sg13g2_inv_1 _12841__62 (.Y(net81),
    .A(clknet_4_7_0_clk));
 sg13g2_inv_1 _12842__63 (.Y(net82),
    .A(clknet_4_6_0_clk));
 sg13g2_inv_1 _12843__64 (.Y(net83),
    .A(clknet_4_9_0_clk));
 sg13g2_inv_1 _12844__65 (.Y(net84),
    .A(clknet_4_3_0_clk));
 sg13g2_inv_1 _12845__66 (.Y(net85),
    .A(clknet_4_3_0_clk));
 sg13g2_inv_1 _12846__67 (.Y(net86),
    .A(clknet_4_12_0_clk));
 sg13g2_inv_1 _12847__68 (.Y(net87),
    .A(clknet_4_6_0_clk));
 sg13g2_inv_1 _12848__69 (.Y(net88),
    .A(clknet_4_7_0_clk));
 sg13g2_inv_1 _12849__70 (.Y(net89),
    .A(clknet_4_7_0_clk));
 sg13g2_inv_1 _12850__71 (.Y(net90),
    .A(clknet_4_13_0_clk));
 sg13g2_inv_1 _12851__72 (.Y(net91),
    .A(clknet_4_11_0_clk));
 sg13g2_inv_1 _12852__73 (.Y(net92),
    .A(clknet_4_10_0_clk));
 sg13g2_inv_1 _12853__74 (.Y(net93),
    .A(clknet_4_11_0_clk));
 sg13g2_inv_1 _12854__75 (.Y(net94),
    .A(clknet_4_14_0_clk));
 sg13g2_inv_1 _12855__76 (.Y(net95),
    .A(clknet_4_15_0_clk));
 sg13g2_inv_1 _12856__77 (.Y(net96),
    .A(clknet_4_15_0_clk));
 sg13g2_inv_1 _12857__78 (.Y(net97),
    .A(clknet_4_13_0_clk));
 sg13g2_inv_1 _12858__79 (.Y(net98),
    .A(clknet_4_12_0_clk));
 sg13g2_inv_1 _12859__80 (.Y(net99),
    .A(clknet_4_11_0_clk));
 sg13g2_inv_1 _12860__81 (.Y(net100),
    .A(clknet_4_10_0_clk));
 sg13g2_inv_1 _12861__82 (.Y(net101),
    .A(clknet_4_11_0_clk));
 sg13g2_inv_1 _12862__83 (.Y(net102),
    .A(clknet_4_14_0_clk));
 sg13g2_inv_1 _12863__84 (.Y(net103),
    .A(clknet_4_15_0_clk));
 sg13g2_inv_1 _12864__85 (.Y(net104),
    .A(clknet_4_15_0_clk));
 sg13g2_inv_1 _12865__86 (.Y(net105),
    .A(clknet_4_13_0_clk));
 sg13g2_inv_1 _12866__87 (.Y(net106),
    .A(clknet_4_9_0_clk));
 sg13g2_inv_1 _12867__88 (.Y(net107),
    .A(clknet_4_2_0_clk));
 sg13g2_inv_1 _12868__89 (.Y(net108),
    .A(clknet_4_2_0_clk));
 sg13g2_inv_1 _12869__90 (.Y(net109),
    .A(clknet_4_8_0_clk));
 sg13g2_inv_1 _12870__91 (.Y(net110),
    .A(clknet_4_2_0_clk));
 sg13g2_inv_1 _12871__92 (.Y(net111),
    .A(clknet_4_2_0_clk));
 sg13g2_inv_1 _12872__93 (.Y(net112),
    .A(clknet_4_8_0_clk));
 sg13g2_inv_1 _12873__94 (.Y(net113),
    .A(clknet_4_2_0_clk));
 sg13g2_inv_1 _12874__95 (.Y(net114),
    .A(clknet_4_3_0_clk));
 sg13g2_inv_1 _12875__96 (.Y(net115),
    .A(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_regs_0_clk (.A(clk),
    .X(clk_regs));
 sg13g2_buf_1 _12876_ (.A(net128),
    .X(_00674_));
 sg13g2_buf_1 _12877_ (.A(net132),
    .X(_00675_));
 sg13g2_dfrbp_1 _12878_ (.CLK(clknet_leaf_82_clk_regs),
    .RESET_B(net3494),
    .D(net1175),
    .Q_N(_06876_),
    .Q(\u_toplayer.u_layer2.u_neuron.instCtrl.state[0] ));
 sg13g2_dfrbp_1 _12879_ (.CLK(clknet_leaf_82_clk_regs),
    .RESET_B(net3494),
    .D(net1073),
    .Q_N(_06877_),
    .Q(\u_toplayer.u_layer2.u_neuron.instCtrl.state[1] ));
 sg13g2_dfrbp_1 _12880_ (.CLK(clknet_leaf_82_clk_regs),
    .RESET_B(net3493),
    .D(net1135),
    .Q_N(_00040_),
    .Q(\u_toplayer.u_layer2.u_neuron.instCtrl.state[2] ));
 sg13g2_dfrbp_1 _12881_ (.CLK(clknet_leaf_82_clk_regs),
    .RESET_B(net3506),
    .D(net1001),
    .Q_N(_00041_),
    .Q(\u_toplayer.u_layer2.u_neuron.instCtrl.state[3] ));
 sg13g2_dfrbp_1 _12882_ (.CLK(clknet_leaf_82_clk_regs),
    .RESET_B(net3496),
    .D(net934),
    .Q_N(_00042_),
    .Q(\u_toplayer.u_layer2.u_neuron.instCtrl.state[4] ));
 sg13g2_dfrbp_1 _12883_ (.CLK(clknet_leaf_88_clk_regs),
    .RESET_B(net3506),
    .D(net873),
    .Q_N(_00032_),
    .Q(\u_toplayer.u_layer2.u_neuron.instCtrl.state[5] ));
 sg13g2_dfrbp_1 _12884_ (.CLK(clknet_leaf_47_clk_regs),
    .RESET_B(net3556),
    .D(net119),
    .Q_N(_00043_),
    .Q(\u_toplayer.u_layer1.u_neuron.instCtrl.state[0] ));
 sg13g2_dfrbp_1 _12885_ (.CLK(clknet_leaf_47_clk_regs),
    .RESET_B(net3556),
    .D(_00001_),
    .Q_N(_06878_),
    .Q(\u_toplayer.u_layer1.u_neuron.instCtrl.state[1] ));
 sg13g2_dfrbp_1 _12886_ (.CLK(clknet_leaf_47_clk_regs),
    .RESET_B(net3556),
    .D(net1108),
    .Q_N(_00045_),
    .Q(\u_toplayer.u_layer1.u_neuron.instCtrl.state[2] ));
 sg13g2_dfrbp_1 _12887_ (.CLK(clknet_leaf_47_clk_regs),
    .RESET_B(net3556),
    .D(net919),
    .Q_N(_00046_),
    .Q(\u_toplayer.u_layer1.u_neuron.instCtrl.state[3] ));
 sg13g2_dfrbp_1 _12888_ (.CLK(clknet_leaf_47_clk_regs),
    .RESET_B(net3552),
    .D(net512),
    .Q_N(_00047_),
    .Q(\u_toplayer.u_layer1.u_neuron.instCtrl.state[4] ));
 sg13g2_dfrbp_1 _12889_ (.CLK(clknet_leaf_47_clk_regs),
    .RESET_B(net3552),
    .D(net570),
    .Q_N(_00048_),
    .Q(\u_toplayer.u_layer1.u_neuron.instCtrl.state[5] ));
 sg13g2_dfrbp_1 _12890_ (.CLK(clknet_leaf_38_clk_regs),
    .RESET_B(net3552),
    .D(net555),
    .Q_N(_00049_),
    .Q(\u_toplayer.u_layer1.u_neuron.instCtrl.state[6] ));
 sg13g2_dfrbp_1 _12891_ (.CLK(clknet_leaf_47_clk_regs),
    .RESET_B(net3556),
    .D(net772),
    .Q_N(_00044_),
    .Q(\u_toplayer.u_layer1.u_neuron.instCtrl.state[7] ));
 sg13g2_dfrbp_1 _12892_ (.CLK(clknet_leaf_38_clk_regs),
    .RESET_B(net3556),
    .D(net1041),
    .Q_N(_00030_),
    .Q(\u_toplayer.u_layer1.u_neuron.instCtrl.state[8] ));
 sg13g2_dfrbp_1 _12893_ (.CLK(clknet_leaf_29_clk_regs),
    .RESET_B(net3475),
    .D(net902),
    .Q_N(_06875_),
    .Q(\u_toplayer.u_outlayer.u_neuron.mult[0] ));
 sg13g2_dfrbp_1 _12894_ (.CLK(clknet_leaf_29_clk_regs),
    .RESET_B(net3475),
    .D(_00150_),
    .Q_N(_06874_),
    .Q(\u_toplayer.u_outlayer.u_neuron.mult[1] ));
 sg13g2_dfrbp_1 _12895_ (.CLK(clknet_leaf_29_clk_regs),
    .RESET_B(net3477),
    .D(_00151_),
    .Q_N(_06873_),
    .Q(\u_toplayer.u_outlayer.u_neuron.mult[2] ));
 sg13g2_dfrbp_1 _12896_ (.CLK(clknet_leaf_26_clk_regs),
    .RESET_B(net3474),
    .D(_00152_),
    .Q_N(_06872_),
    .Q(\u_toplayer.u_outlayer.u_neuron.mult[3] ));
 sg13g2_dfrbp_1 _12897_ (.CLK(clknet_leaf_26_clk_regs),
    .RESET_B(net3474),
    .D(net875),
    .Q_N(_06871_),
    .Q(\u_toplayer.u_outlayer.u_neuron.mult[4] ));
 sg13g2_dfrbp_1 _12898_ (.CLK(clknet_leaf_26_clk_regs),
    .RESET_B(net3474),
    .D(_00154_),
    .Q_N(_06870_),
    .Q(\u_toplayer.u_outlayer.u_neuron.mult[5] ));
 sg13g2_dfrbp_1 _12899_ (.CLK(clknet_leaf_27_clk_regs),
    .RESET_B(net3476),
    .D(_00155_),
    .Q_N(_06869_),
    .Q(\u_toplayer.u_outlayer.u_neuron.mult[6] ));
 sg13g2_dfrbp_1 _12900_ (.CLK(clknet_leaf_27_clk_regs),
    .RESET_B(net3476),
    .D(_00156_),
    .Q_N(_06868_),
    .Q(\u_toplayer.u_outlayer.u_neuron.mult[7] ));
 sg13g2_dfrbp_1 _12901_ (.CLK(clknet_leaf_27_clk_regs),
    .RESET_B(net3476),
    .D(_00157_),
    .Q_N(_06867_),
    .Q(\u_toplayer.u_outlayer.u_neuron.mult[8] ));
 sg13g2_dfrbp_1 _12902_ (.CLK(clknet_leaf_27_clk_regs),
    .RESET_B(net3476),
    .D(_00158_),
    .Q_N(_06866_),
    .Q(\u_toplayer.u_outlayer.u_neuron.mult[9] ));
 sg13g2_dfrbp_1 _12903_ (.CLK(clknet_leaf_27_clk_regs),
    .RESET_B(net3476),
    .D(_00159_),
    .Q_N(_06865_),
    .Q(\u_toplayer.u_outlayer.u_neuron.mult[10] ));
 sg13g2_dfrbp_1 _12904_ (.CLK(clknet_leaf_27_clk_regs),
    .RESET_B(net3470),
    .D(_00160_),
    .Q_N(_06864_),
    .Q(\u_toplayer.u_outlayer.u_neuron.mult[11] ));
 sg13g2_dfrbp_1 _12905_ (.CLK(clknet_leaf_29_clk_regs),
    .RESET_B(net3477),
    .D(_00161_),
    .Q_N(_06863_),
    .Q(\u_toplayer.u_outlayer.u_neuron.mult[12] ));
 sg13g2_dfrbp_1 _12906_ (.CLK(clknet_leaf_29_clk_regs),
    .RESET_B(net3485),
    .D(_00162_),
    .Q_N(_06862_),
    .Q(\u_toplayer.u_outlayer.u_neuron.mult[13] ));
 sg13g2_dfrbp_1 _12907_ (.CLK(clknet_leaf_29_clk_regs),
    .RESET_B(net3485),
    .D(_00163_),
    .Q_N(_06861_),
    .Q(\u_toplayer.u_outlayer.u_neuron.mult[14] ));
 sg13g2_dfrbp_1 _12908_ (.CLK(clknet_leaf_29_clk_regs),
    .RESET_B(net3485),
    .D(_00164_),
    .Q_N(_06860_),
    .Q(\u_toplayer.u_outlayer.u_neuron.mult[15] ));
 sg13g2_dfrbp_1 _12909_ (.CLK(clknet_leaf_21_clk_regs),
    .RESET_B(net3466),
    .D(net1126),
    .Q_N(_06859_),
    .Q(\u_toplayer.u_outlayer.u_neuron.din[0] ));
 sg13g2_dfrbp_1 _12910_ (.CLK(clknet_leaf_21_clk_regs),
    .RESET_B(net3467),
    .D(net1094),
    .Q_N(_06858_),
    .Q(\u_toplayer.u_outlayer.u_neuron.din[1] ));
 sg13g2_dfrbp_1 _12911_ (.CLK(clknet_leaf_28_clk_regs),
    .RESET_B(net3467),
    .D(_00167_),
    .Q_N(_06857_),
    .Q(\u_toplayer.u_outlayer.u_neuron.din[2] ));
 sg13g2_dfrbp_1 _12912_ (.CLK(clknet_leaf_21_clk_regs),
    .RESET_B(net3466),
    .D(net1139),
    .Q_N(_06856_),
    .Q(\u_toplayer.u_outlayer.u_neuron.din[3] ));
 sg13g2_dfrbp_1 _12913_ (.CLK(clknet_leaf_31_clk_regs),
    .RESET_B(net3481),
    .D(_00169_),
    .Q_N(_06855_),
    .Q(\u_toplayer.u_outlayer.u_neuron.din[4] ));
 sg13g2_dfrbp_1 _12914_ (.CLK(clknet_leaf_31_clk_regs),
    .RESET_B(net3480),
    .D(net1057),
    .Q_N(_06854_),
    .Q(\u_toplayer.u_outlayer.u_neuron.din[5] ));
 sg13g2_dfrbp_1 _12915_ (.CLK(clknet_leaf_31_clk_regs),
    .RESET_B(net3480),
    .D(net1097),
    .Q_N(_06853_),
    .Q(\u_toplayer.u_outlayer.u_neuron.din[6] ));
 sg13g2_dfrbp_1 _12916_ (.CLK(clknet_leaf_28_clk_regs),
    .RESET_B(net3485),
    .D(net1091),
    .Q_N(_06852_),
    .Q(\u_toplayer.u_outlayer.u_neuron.din[7] ));
 sg13g2_dfrbp_1 _12917_ (.CLK(clknet_leaf_25_clk_regs),
    .RESET_B(net3475),
    .D(net905),
    .Q_N(_06851_),
    .Q(uo_out[0]));
 sg13g2_dfrbp_1 _12918_ (.CLK(clknet_leaf_26_clk_regs),
    .RESET_B(net3475),
    .D(_00174_),
    .Q_N(_06850_),
    .Q(uo_out[1]));
 sg13g2_dfrbp_1 _12919_ (.CLK(clknet_leaf_25_clk_regs),
    .RESET_B(net3474),
    .D(net808),
    .Q_N(_06849_),
    .Q(uo_out[2]));
 sg13g2_dfrbp_1 _12920_ (.CLK(clknet_leaf_25_clk_regs),
    .RESET_B(net3474),
    .D(net850),
    .Q_N(_06848_),
    .Q(uo_out[3]));
 sg13g2_dfrbp_1 _12921_ (.CLK(clknet_leaf_25_clk_regs),
    .RESET_B(net3474),
    .D(net900),
    .Q_N(_06847_),
    .Q(uo_out[4]));
 sg13g2_dfrbp_1 _12922_ (.CLK(clknet_leaf_25_clk_regs),
    .RESET_B(net3472),
    .D(net909),
    .Q_N(_06846_),
    .Q(uo_out[5]));
 sg13g2_dfrbp_1 _12923_ (.CLK(clknet_leaf_25_clk_regs),
    .RESET_B(net3472),
    .D(net867),
    .Q_N(_06845_),
    .Q(uo_out[6]));
 sg13g2_dfrbp_1 _12924_ (.CLK(clknet_leaf_24_clk_regs),
    .RESET_B(net3472),
    .D(net985),
    .Q_N(_06844_),
    .Q(uo_out[7]));
 sg13g2_dfrbp_1 _12925_ (.CLK(clknet_leaf_34_clk_regs),
    .RESET_B(net3484),
    .D(net928),
    .Q_N(_06843_),
    .Q(\u_toplayer.u_layer3.u_neuron.mult[0] ));
 sg13g2_dfrbp_1 _12926_ (.CLK(clknet_leaf_34_clk_regs),
    .RESET_B(net3484),
    .D(_00182_),
    .Q_N(_06842_),
    .Q(\u_toplayer.u_layer3.u_neuron.mult[1] ));
 sg13g2_dfrbp_1 _12927_ (.CLK(clknet_leaf_34_clk_regs),
    .RESET_B(net3484),
    .D(_00183_),
    .Q_N(_06841_),
    .Q(\u_toplayer.u_layer3.u_neuron.mult[2] ));
 sg13g2_dfrbp_1 _12928_ (.CLK(clknet_leaf_34_clk_regs),
    .RESET_B(net3484),
    .D(_00184_),
    .Q_N(_06840_),
    .Q(\u_toplayer.u_layer3.u_neuron.mult[3] ));
 sg13g2_dfrbp_1 _12929_ (.CLK(clknet_leaf_34_clk_regs),
    .RESET_B(net3483),
    .D(_00185_),
    .Q_N(_06839_),
    .Q(\u_toplayer.u_layer3.u_neuron.mult[4] ));
 sg13g2_dfrbp_1 _12930_ (.CLK(clknet_leaf_36_clk_regs),
    .RESET_B(net3549),
    .D(_00186_),
    .Q_N(_06838_),
    .Q(\u_toplayer.u_layer3.u_neuron.mult[5] ));
 sg13g2_dfrbp_1 _12931_ (.CLK(clknet_leaf_35_clk_regs),
    .RESET_B(net3483),
    .D(_00187_),
    .Q_N(_06837_),
    .Q(\u_toplayer.u_layer3.u_neuron.mult[6] ));
 sg13g2_dfrbp_1 _12932_ (.CLK(clknet_leaf_36_clk_regs),
    .RESET_B(net3549),
    .D(_00188_),
    .Q_N(_06836_),
    .Q(\u_toplayer.u_layer3.u_neuron.mult[7] ));
 sg13g2_dfrbp_1 _12933_ (.CLK(clknet_leaf_37_clk_regs),
    .RESET_B(net3549),
    .D(_00189_),
    .Q_N(_06835_),
    .Q(\u_toplayer.u_layer3.u_neuron.mult[8] ));
 sg13g2_dfrbp_1 _12934_ (.CLK(clknet_leaf_37_clk_regs),
    .RESET_B(net3549),
    .D(_00190_),
    .Q_N(_06834_),
    .Q(\u_toplayer.u_layer3.u_neuron.mult[9] ));
 sg13g2_dfrbp_1 _12935_ (.CLK(clknet_leaf_38_clk_regs),
    .RESET_B(net3549),
    .D(_00191_),
    .Q_N(_06833_),
    .Q(\u_toplayer.u_layer3.u_neuron.mult[10] ));
 sg13g2_dfrbp_1 _12936_ (.CLK(clknet_leaf_38_clk_regs),
    .RESET_B(net3549),
    .D(_00192_),
    .Q_N(_06832_),
    .Q(\u_toplayer.u_layer3.u_neuron.mult[11] ));
 sg13g2_dfrbp_1 _12937_ (.CLK(clknet_leaf_38_clk_regs),
    .RESET_B(net3552),
    .D(_00193_),
    .Q_N(_06831_),
    .Q(\u_toplayer.u_layer3.u_neuron.mult[12] ));
 sg13g2_dfrbp_1 _12938_ (.CLK(clknet_leaf_37_clk_regs),
    .RESET_B(net3549),
    .D(_00194_),
    .Q_N(_06830_),
    .Q(\u_toplayer.u_layer3.u_neuron.mult[13] ));
 sg13g2_dfrbp_1 _12939_ (.CLK(clknet_leaf_36_clk_regs),
    .RESET_B(net3550),
    .D(_00195_),
    .Q_N(_06829_),
    .Q(\u_toplayer.u_layer3.u_neuron.mult[14] ));
 sg13g2_dfrbp_1 _12940_ (.CLK(clknet_leaf_37_clk_regs),
    .RESET_B(net3552),
    .D(_00196_),
    .Q_N(_06828_),
    .Q(\u_toplayer.u_layer3.u_neuron.mult[15] ));
 sg13g2_dfrbp_1 _12941_ (.CLK(clknet_leaf_26_clk_regs),
    .RESET_B(net3475),
    .D(_00197_),
    .Q_N(_06827_),
    .Q(\u_toplayer.u_outlayer.u_neuron.acc[0] ));
 sg13g2_dfrbp_1 _12942_ (.CLK(clknet_leaf_26_clk_regs),
    .RESET_B(net3475),
    .D(_00198_),
    .Q_N(_06826_),
    .Q(\u_toplayer.u_outlayer.u_neuron.acc[1] ));
 sg13g2_dfrbp_1 _12943_ (.CLK(clknet_leaf_26_clk_regs),
    .RESET_B(net3475),
    .D(_00199_),
    .Q_N(_06825_),
    .Q(\u_toplayer.u_outlayer.u_neuron.acc[2] ));
 sg13g2_dfrbp_1 _12944_ (.CLK(clknet_leaf_26_clk_regs),
    .RESET_B(net3474),
    .D(_00200_),
    .Q_N(_06824_),
    .Q(\u_toplayer.u_outlayer.u_neuron.acc[3] ));
 sg13g2_dfrbp_1 _12945_ (.CLK(clknet_leaf_25_clk_regs),
    .RESET_B(net3474),
    .D(_00201_),
    .Q_N(_06823_),
    .Q(\u_toplayer.u_outlayer.u_neuron.acc[4] ));
 sg13g2_dfrbp_1 _12946_ (.CLK(clknet_leaf_24_clk_regs),
    .RESET_B(net3471),
    .D(_00202_),
    .Q_N(_06822_),
    .Q(\u_toplayer.u_outlayer.u_neuron.acc[5] ));
 sg13g2_dfrbp_1 _12947_ (.CLK(clknet_leaf_25_clk_regs),
    .RESET_B(net3472),
    .D(_00203_),
    .Q_N(_06821_),
    .Q(\u_toplayer.u_outlayer.u_neuron.acc[6] ));
 sg13g2_dfrbp_1 _12948_ (.CLK(clknet_leaf_23_clk_regs),
    .RESET_B(net3470),
    .D(net1162),
    .Q_N(_06820_),
    .Q(\u_toplayer.u_outlayer.u_neuron.acc[7] ));
 sg13g2_dfrbp_1 _12949_ (.CLK(clknet_leaf_22_clk_regs),
    .RESET_B(net3470),
    .D(_00205_),
    .Q_N(_06819_),
    .Q(\u_toplayer.u_outlayer.u_neuron.acc[8] ));
 sg13g2_dfrbp_1 _12950_ (.CLK(clknet_leaf_22_clk_regs),
    .RESET_B(net3470),
    .D(_00206_),
    .Q_N(_06818_),
    .Q(\u_toplayer.u_outlayer.u_neuron.acc[9] ));
 sg13g2_dfrbp_1 _12951_ (.CLK(clknet_leaf_21_clk_regs),
    .RESET_B(net3473),
    .D(_00207_),
    .Q_N(_06817_),
    .Q(\u_toplayer.u_outlayer.u_neuron.acc[10] ));
 sg13g2_dfrbp_1 _12952_ (.CLK(clknet_leaf_27_clk_regs),
    .RESET_B(net3470),
    .D(_00208_),
    .Q_N(_06816_),
    .Q(\u_toplayer.u_outlayer.u_neuron.acc[11] ));
 sg13g2_dfrbp_1 _12953_ (.CLK(clknet_leaf_22_clk_regs),
    .RESET_B(net3470),
    .D(_00209_),
    .Q_N(_06815_),
    .Q(\u_toplayer.u_outlayer.u_neuron.acc[12] ));
 sg13g2_dfrbp_1 _12954_ (.CLK(clknet_leaf_22_clk_regs),
    .RESET_B(net3470),
    .D(_00210_),
    .Q_N(_06814_),
    .Q(\u_toplayer.u_outlayer.u_neuron.acc[13] ));
 sg13g2_dfrbp_1 _12955_ (.CLK(clknet_leaf_22_clk_regs),
    .RESET_B(net3470),
    .D(_00211_),
    .Q_N(_06813_),
    .Q(\u_toplayer.u_outlayer.u_neuron.acc[14] ));
 sg13g2_dfrbp_1 _12956_ (.CLK(clknet_leaf_23_clk_regs),
    .RESET_B(net3471),
    .D(_00212_),
    .Q_N(_06812_),
    .Q(\u_toplayer.u_outlayer.u_neuron.acc[15] ));
 sg13g2_dfrbp_1 _12957_ (.CLK(clknet_leaf_24_clk_regs),
    .RESET_B(net3471),
    .D(_00213_),
    .Q_N(_06811_),
    .Q(\u_toplayer.u_outlayer.u_neuron.acc[16] ));
 sg13g2_dfrbp_1 _12958_ (.CLK(clknet_leaf_24_clk_regs),
    .RESET_B(net3471),
    .D(_00214_),
    .Q_N(_06810_),
    .Q(\u_toplayer.u_outlayer.u_neuron.acc[17] ));
 sg13g2_dfrbp_1 _12959_ (.CLK(clknet_leaf_24_clk_regs),
    .RESET_B(net3471),
    .D(_00215_),
    .Q_N(_06809_),
    .Q(\u_toplayer.u_outlayer.u_neuron.acc[18] ));
 sg13g2_dfrbp_1 _12960_ (.CLK(clknet_leaf_24_clk_regs),
    .RESET_B(net3471),
    .D(_00216_),
    .Q_N(_06808_),
    .Q(\u_toplayer.u_outlayer.u_neuron.acc[19] ));
 sg13g2_dfrbp_1 _12961_ (.CLK(clknet_leaf_23_clk_regs),
    .RESET_B(net3471),
    .D(_00217_),
    .Q_N(_06807_),
    .Q(\u_toplayer.u_outlayer.u_neuron.acc[20] ));
 sg13g2_dfrbp_1 _12962_ (.CLK(clknet_leaf_23_clk_regs),
    .RESET_B(net3471),
    .D(_00218_),
    .Q_N(_06806_),
    .Q(\u_toplayer.u_outlayer.u_neuron.acc[21] ));
 sg13g2_dfrbp_1 _12963_ (.CLK(clknet_leaf_23_clk_regs),
    .RESET_B(net3472),
    .D(_00219_),
    .Q_N(_06805_),
    .Q(\u_toplayer.u_outlayer.u_neuron.acc[22] ));
 sg13g2_dfrbp_1 _12964_ (.CLK(clknet_leaf_24_clk_regs),
    .RESET_B(net3472),
    .D(_00220_),
    .Q_N(_06804_),
    .Q(\u_toplayer.u_outlayer.u_neuron.acc[23] ));
 sg13g2_dfrbp_1 _12965_ (.CLK(net20),
    .RESET_B(net3422),
    .D(net832),
    .Q_N(_00052_),
    .Q(\u_toplayer.u_layer3.neuron_index[0] ));
 sg13g2_dfrbp_1 _12966_ (.CLK(net21),
    .RESET_B(net3423),
    .D(_00222_),
    .Q_N(_06803_),
    .Q(\u_toplayer.u_layer3.neuron_index[1] ));
 sg13g2_dfrbp_1 _12967_ (.CLK(net22),
    .RESET_B(net3424),
    .D(net1099),
    .Q_N(_06802_),
    .Q(\u_toplayer.u_layer3.neuron_index[2] ));
 sg13g2_dfrbp_1 _12968_ (.CLK(net23),
    .RESET_B(net3424),
    .D(net1191),
    .Q_N(_06801_),
    .Q(\u_toplayer.u_layer3.neuron_index[3] ));
 sg13g2_dfrbp_1 _12969_ (.CLK(net24),
    .RESET_B(net3425),
    .D(net1035),
    .Q_N(_06800_),
    .Q(\u_toplayer.u_layer3.neuron_index[4] ));
 sg13g2_dfrbp_1 _12970_ (.CLK(net25),
    .RESET_B(net3425),
    .D(net1025),
    .Q_N(_06799_),
    .Q(\u_toplayer.u_layer3.neuron_index[5] ));
 sg13g2_dfrbp_1 _12971_ (.CLK(clknet_leaf_49_clk_regs),
    .RESET_B(net3550),
    .D(net930),
    .Q_N(_06798_),
    .Q(\u_toplayer.u_layer2.u_neuron.mult[0] ));
 sg13g2_dfrbp_1 _12972_ (.CLK(clknet_leaf_35_clk_regs),
    .RESET_B(net3550),
    .D(_00228_),
    .Q_N(_06797_),
    .Q(\u_toplayer.u_layer2.u_neuron.mult[1] ));
 sg13g2_dfrbp_1 _12973_ (.CLK(clknet_leaf_35_clk_regs),
    .RESET_B(net3550),
    .D(_00229_),
    .Q_N(_06796_),
    .Q(\u_toplayer.u_layer2.u_neuron.mult[2] ));
 sg13g2_dfrbp_1 _12974_ (.CLK(clknet_leaf_34_clk_regs),
    .RESET_B(net3550),
    .D(_00230_),
    .Q_N(_06795_),
    .Q(\u_toplayer.u_layer2.u_neuron.mult[3] ));
 sg13g2_dfrbp_1 _12975_ (.CLK(clknet_leaf_17_clk_regs),
    .RESET_B(net3550),
    .D(_00231_),
    .Q_N(_06794_),
    .Q(\u_toplayer.u_layer2.u_neuron.mult[4] ));
 sg13g2_dfrbp_1 _12976_ (.CLK(clknet_leaf_91_clk_regs),
    .RESET_B(net3550),
    .D(_00232_),
    .Q_N(_06793_),
    .Q(\u_toplayer.u_layer2.u_neuron.mult[5] ));
 sg13g2_dfrbp_1 _12977_ (.CLK(clknet_leaf_17_clk_regs),
    .RESET_B(net3508),
    .D(_00233_),
    .Q_N(_06792_),
    .Q(\u_toplayer.u_layer2.u_neuron.mult[6] ));
 sg13g2_dfrbp_1 _12978_ (.CLK(clknet_leaf_17_clk_regs),
    .RESET_B(net3508),
    .D(_00234_),
    .Q_N(_06791_),
    .Q(\u_toplayer.u_layer2.u_neuron.mult[7] ));
 sg13g2_dfrbp_1 _12979_ (.CLK(clknet_leaf_17_clk_regs),
    .RESET_B(net3454),
    .D(_00235_),
    .Q_N(_06790_),
    .Q(\u_toplayer.u_layer2.u_neuron.mult[8] ));
 sg13g2_dfrbp_1 _12980_ (.CLK(clknet_leaf_17_clk_regs),
    .RESET_B(net3454),
    .D(_00236_),
    .Q_N(_06789_),
    .Q(\u_toplayer.u_layer2.u_neuron.mult[9] ));
 sg13g2_dfrbp_1 _12981_ (.CLK(clknet_leaf_16_clk_regs),
    .RESET_B(net3453),
    .D(_00237_),
    .Q_N(_06788_),
    .Q(\u_toplayer.u_layer2.u_neuron.mult[10] ));
 sg13g2_dfrbp_1 _12982_ (.CLK(clknet_leaf_15_clk_regs),
    .RESET_B(net3453),
    .D(_00238_),
    .Q_N(_06787_),
    .Q(\u_toplayer.u_layer2.u_neuron.mult[11] ));
 sg13g2_dfrbp_1 _12983_ (.CLK(clknet_leaf_16_clk_regs),
    .RESET_B(net3454),
    .D(_00239_),
    .Q_N(_06786_),
    .Q(\u_toplayer.u_layer2.u_neuron.mult[12] ));
 sg13g2_dfrbp_1 _12984_ (.CLK(clknet_leaf_16_clk_regs),
    .RESET_B(net3454),
    .D(_00240_),
    .Q_N(_06785_),
    .Q(\u_toplayer.u_layer2.u_neuron.mult[13] ));
 sg13g2_dfrbp_1 _12985_ (.CLK(clknet_leaf_92_clk_regs),
    .RESET_B(net3452),
    .D(_00241_),
    .Q_N(_06784_),
    .Q(\u_toplayer.u_layer2.u_neuron.mult[14] ));
 sg13g2_dfrbp_1 _12986_ (.CLK(clknet_leaf_16_clk_regs),
    .RESET_B(net3454),
    .D(_00242_),
    .Q_N(_06783_),
    .Q(\u_toplayer.u_layer2.u_neuron.mult[15] ));
 sg13g2_dfrbp_1 _12987_ (.CLK(net26),
    .RESET_B(net3466),
    .D(_00243_),
    .Q_N(_06782_),
    .Q(\u_toplayer.outreg[0] ));
 sg13g2_dfrbp_1 _12988_ (.CLK(net27),
    .RESET_B(net3464),
    .D(_00244_),
    .Q_N(_06781_),
    .Q(\u_toplayer.outreg[1] ));
 sg13g2_dfrbp_1 _12989_ (.CLK(net28),
    .RESET_B(net3479),
    .D(_00245_),
    .Q_N(_06780_),
    .Q(\u_toplayer.outreg[2] ));
 sg13g2_dfrbp_1 _12990_ (.CLK(net29),
    .RESET_B(net3463),
    .D(_00246_),
    .Q_N(_06779_),
    .Q(\u_toplayer.outreg[3] ));
 sg13g2_dfrbp_1 _12991_ (.CLK(net30),
    .RESET_B(net3478),
    .D(_00247_),
    .Q_N(_06778_),
    .Q(\u_toplayer.outreg[4] ));
 sg13g2_dfrbp_1 _12992_ (.CLK(net31),
    .RESET_B(net3480),
    .D(_00248_),
    .Q_N(_06777_),
    .Q(\u_toplayer.outreg[5] ));
 sg13g2_dfrbp_1 _12993_ (.CLK(net32),
    .RESET_B(net3480),
    .D(_00249_),
    .Q_N(_06776_),
    .Q(\u_toplayer.outreg[6] ));
 sg13g2_dfrbp_1 _12994_ (.CLK(net33),
    .RESET_B(net3466),
    .D(_00250_),
    .Q_N(_06775_),
    .Q(\u_toplayer.outreg[7] ));
 sg13g2_dfrbp_1 _12995_ (.CLK(net34),
    .RESET_B(net3466),
    .D(_00251_),
    .Q_N(_06774_),
    .Q(\u_toplayer.outreg[8] ));
 sg13g2_dfrbp_1 _12996_ (.CLK(net35),
    .RESET_B(net3463),
    .D(_00252_),
    .Q_N(_06773_),
    .Q(\u_toplayer.outreg[9] ));
 sg13g2_dfrbp_1 _12997_ (.CLK(net36),
    .RESET_B(net3479),
    .D(_00253_),
    .Q_N(_06772_),
    .Q(\u_toplayer.outreg[10] ));
 sg13g2_dfrbp_1 _12998_ (.CLK(net37),
    .RESET_B(net3463),
    .D(_00254_),
    .Q_N(_06771_),
    .Q(\u_toplayer.outreg[11] ));
 sg13g2_dfrbp_1 _12999_ (.CLK(net38),
    .RESET_B(net3478),
    .D(_00255_),
    .Q_N(_06770_),
    .Q(\u_toplayer.outreg[12] ));
 sg13g2_dfrbp_1 _13000_ (.CLK(net39),
    .RESET_B(net3480),
    .D(_00256_),
    .Q_N(_06769_),
    .Q(\u_toplayer.outreg[13] ));
 sg13g2_dfrbp_1 _13001_ (.CLK(net40),
    .RESET_B(net3480),
    .D(net156),
    .Q_N(_06768_),
    .Q(\u_toplayer.outreg[14] ));
 sg13g2_dfrbp_1 _13002_ (.CLK(net41),
    .RESET_B(net3466),
    .D(_00258_),
    .Q_N(_06767_),
    .Q(\u_toplayer.outreg[15] ));
 sg13g2_dfrbp_1 _13003_ (.CLK(net42),
    .RESET_B(net3459),
    .D(_00259_),
    .Q_N(_06766_),
    .Q(\u_toplayer.outreg[16] ));
 sg13g2_dfrbp_1 _13004_ (.CLK(net43),
    .RESET_B(net3457),
    .D(_00260_),
    .Q_N(_06765_),
    .Q(\u_toplayer.outreg[17] ));
 sg13g2_dfrbp_1 _13005_ (.CLK(net44),
    .RESET_B(net3458),
    .D(_00261_),
    .Q_N(_06764_),
    .Q(\u_toplayer.outreg[18] ));
 sg13g2_dfrbp_1 _13006_ (.CLK(net45),
    .RESET_B(net3458),
    .D(_00262_),
    .Q_N(_06763_),
    .Q(\u_toplayer.outreg[19] ));
 sg13g2_dfrbp_1 _13007_ (.CLK(net46),
    .RESET_B(net3457),
    .D(_00263_),
    .Q_N(_06762_),
    .Q(\u_toplayer.outreg[20] ));
 sg13g2_dfrbp_1 _13008_ (.CLK(net47),
    .RESET_B(net3459),
    .D(_00264_),
    .Q_N(_06761_),
    .Q(\u_toplayer.outreg[21] ));
 sg13g2_dfrbp_1 _13009_ (.CLK(net48),
    .RESET_B(net3459),
    .D(_00265_),
    .Q_N(_06760_),
    .Q(\u_toplayer.outreg[22] ));
 sg13g2_dfrbp_1 _13010_ (.CLK(net49),
    .RESET_B(net3460),
    .D(_00266_),
    .Q_N(_06759_),
    .Q(\u_toplayer.outreg[23] ));
 sg13g2_dfrbp_1 _13011_ (.CLK(net50),
    .RESET_B(net3459),
    .D(_00267_),
    .Q_N(_06758_),
    .Q(\u_toplayer.outreg[24] ));
 sg13g2_dfrbp_1 _13012_ (.CLK(net51),
    .RESET_B(net3457),
    .D(_00268_),
    .Q_N(_06757_),
    .Q(\u_toplayer.outreg[25] ));
 sg13g2_dfrbp_1 _13013_ (.CLK(net52),
    .RESET_B(net3458),
    .D(_00269_),
    .Q_N(_06756_),
    .Q(\u_toplayer.outreg[26] ));
 sg13g2_dfrbp_1 _13014_ (.CLK(net53),
    .RESET_B(net3458),
    .D(_00270_),
    .Q_N(_06755_),
    .Q(\u_toplayer.outreg[27] ));
 sg13g2_dfrbp_1 _13015_ (.CLK(net54),
    .RESET_B(net3457),
    .D(_00271_),
    .Q_N(_06754_),
    .Q(\u_toplayer.outreg[28] ));
 sg13g2_dfrbp_1 _13016_ (.CLK(net55),
    .RESET_B(net3459),
    .D(_00272_),
    .Q_N(_06753_),
    .Q(\u_toplayer.outreg[29] ));
 sg13g2_dfrbp_1 _13017_ (.CLK(net56),
    .RESET_B(net3459),
    .D(_00273_),
    .Q_N(_06752_),
    .Q(\u_toplayer.outreg[30] ));
 sg13g2_dfrbp_1 _13018_ (.CLK(net57),
    .RESET_B(net3460),
    .D(net154),
    .Q_N(_06751_),
    .Q(\u_toplayer.outreg[31] ));
 sg13g2_dfrbp_1 _13019_ (.CLK(net58),
    .RESET_B(net3457),
    .D(_00275_),
    .Q_N(_06750_),
    .Q(\u_toplayer.outreg[32] ));
 sg13g2_dfrbp_1 _13020_ (.CLK(net59),
    .RESET_B(net3457),
    .D(_00276_),
    .Q_N(_06749_),
    .Q(\u_toplayer.outreg[33] ));
 sg13g2_dfrbp_1 _13021_ (.CLK(net60),
    .RESET_B(net3461),
    .D(_00277_),
    .Q_N(_06748_),
    .Q(\u_toplayer.outreg[34] ));
 sg13g2_dfrbp_1 _13022_ (.CLK(net61),
    .RESET_B(net3458),
    .D(_00278_),
    .Q_N(_06747_),
    .Q(\u_toplayer.outreg[35] ));
 sg13g2_dfrbp_1 _13023_ (.CLK(net62),
    .RESET_B(net3458),
    .D(_00279_),
    .Q_N(_06746_),
    .Q(\u_toplayer.outreg[36] ));
 sg13g2_dfrbp_1 _13024_ (.CLK(net63),
    .RESET_B(net3459),
    .D(_00280_),
    .Q_N(_06745_),
    .Q(\u_toplayer.outreg[37] ));
 sg13g2_dfrbp_1 _13025_ (.CLK(net64),
    .RESET_B(net3465),
    .D(_00281_),
    .Q_N(_06744_),
    .Q(\u_toplayer.outreg[38] ));
 sg13g2_dfrbp_1 _13026_ (.CLK(net65),
    .RESET_B(net3460),
    .D(net136),
    .Q_N(_06743_),
    .Q(\u_toplayer.outreg[39] ));
 sg13g2_dfrbp_1 _13027_ (.CLK(net66),
    .RESET_B(net3462),
    .D(_00283_),
    .Q_N(_06742_),
    .Q(\u_toplayer.outreg[40] ));
 sg13g2_dfrbp_1 _13028_ (.CLK(net67),
    .RESET_B(net3457),
    .D(_00284_),
    .Q_N(_06741_),
    .Q(\u_toplayer.outreg[41] ));
 sg13g2_dfrbp_1 _13029_ (.CLK(net68),
    .RESET_B(net3461),
    .D(_00285_),
    .Q_N(_06740_),
    .Q(\u_toplayer.outreg[42] ));
 sg13g2_dfrbp_1 _13030_ (.CLK(net69),
    .RESET_B(net3461),
    .D(_00286_),
    .Q_N(_06739_),
    .Q(\u_toplayer.outreg[43] ));
 sg13g2_dfrbp_1 _13031_ (.CLK(net70),
    .RESET_B(net3457),
    .D(_00287_),
    .Q_N(_06738_),
    .Q(\u_toplayer.outreg[44] ));
 sg13g2_dfrbp_1 _13032_ (.CLK(net71),
    .RESET_B(net3465),
    .D(_00288_),
    .Q_N(_06737_),
    .Q(\u_toplayer.outreg[45] ));
 sg13g2_dfrbp_1 _13033_ (.CLK(net72),
    .RESET_B(net3465),
    .D(net218),
    .Q_N(_06736_),
    .Q(\u_toplayer.outreg[46] ));
 sg13g2_dfrbp_1 _13034_ (.CLK(net73),
    .RESET_B(net3465),
    .D(_00290_),
    .Q_N(_06735_),
    .Q(\u_toplayer.outreg[47] ));
 sg13g2_dfrbp_1 _13035_ (.CLK(net74),
    .RESET_B(net3459),
    .D(_00291_),
    .Q_N(_06734_),
    .Q(\u_toplayer.outreg[48] ));
 sg13g2_dfrbp_1 _13036_ (.CLK(net75),
    .RESET_B(net3461),
    .D(_00292_),
    .Q_N(_06733_),
    .Q(\u_toplayer.outreg[49] ));
 sg13g2_dfrbp_1 _13037_ (.CLK(net76),
    .RESET_B(net3461),
    .D(_00293_),
    .Q_N(_06732_),
    .Q(\u_toplayer.outreg[50] ));
 sg13g2_dfrbp_1 _13038_ (.CLK(net77),
    .RESET_B(net3461),
    .D(_00294_),
    .Q_N(_06731_),
    .Q(\u_toplayer.outreg[51] ));
 sg13g2_dfrbp_1 _13039_ (.CLK(net78),
    .RESET_B(net3462),
    .D(_00295_),
    .Q_N(_06730_),
    .Q(\u_toplayer.outreg[52] ));
 sg13g2_dfrbp_1 _13040_ (.CLK(net79),
    .RESET_B(net3460),
    .D(_00296_),
    .Q_N(_06729_),
    .Q(\u_toplayer.outreg[53] ));
 sg13g2_dfrbp_1 _13041_ (.CLK(net80),
    .RESET_B(net3465),
    .D(_00297_),
    .Q_N(_06728_),
    .Q(\u_toplayer.outreg[54] ));
 sg13g2_dfrbp_1 _13042_ (.CLK(net81),
    .RESET_B(net3468),
    .D(_00298_),
    .Q_N(_06727_),
    .Q(\u_toplayer.outreg[55] ));
 sg13g2_dfrbp_1 _13043_ (.CLK(net82),
    .RESET_B(net3460),
    .D(_00299_),
    .Q_N(_06726_),
    .Q(\u_toplayer.outreg[56] ));
 sg13g2_dfrbp_1 _13044_ (.CLK(net83),
    .RESET_B(net3462),
    .D(_00300_),
    .Q_N(_06725_),
    .Q(\u_toplayer.outreg[57] ));
 sg13g2_dfrbp_1 _13045_ (.CLK(net84),
    .RESET_B(net3461),
    .D(_00301_),
    .Q_N(_06724_),
    .Q(\u_toplayer.outreg[58] ));
 sg13g2_dfrbp_1 _13046_ (.CLK(net85),
    .RESET_B(net3461),
    .D(_00302_),
    .Q_N(_06723_),
    .Q(\u_toplayer.outreg[59] ));
 sg13g2_dfrbp_1 _13047_ (.CLK(net86),
    .RESET_B(net3462),
    .D(_00303_),
    .Q_N(_06722_),
    .Q(\u_toplayer.outreg[60] ));
 sg13g2_dfrbp_1 _13048_ (.CLK(net87),
    .RESET_B(net3460),
    .D(_00304_),
    .Q_N(_06721_),
    .Q(\u_toplayer.outreg[61] ));
 sg13g2_dfrbp_1 _13049_ (.CLK(net88),
    .RESET_B(net3465),
    .D(_00305_),
    .Q_N(_06720_),
    .Q(\u_toplayer.outreg[62] ));
 sg13g2_dfrbp_1 _13050_ (.CLK(net89),
    .RESET_B(net3468),
    .D(_00306_),
    .Q_N(_06719_),
    .Q(\u_toplayer.outreg[63] ));
 sg13g2_dfrbp_1 _13051_ (.CLK(net90),
    .RESET_B(net3465),
    .D(_00307_),
    .Q_N(_06718_),
    .Q(\u_toplayer.outreg[64] ));
 sg13g2_dfrbp_1 _13052_ (.CLK(net91),
    .RESET_B(net3463),
    .D(_00308_),
    .Q_N(_06717_),
    .Q(\u_toplayer.outreg[65] ));
 sg13g2_dfrbp_1 _13053_ (.CLK(net92),
    .RESET_B(net3478),
    .D(_00309_),
    .Q_N(_06716_),
    .Q(\u_toplayer.outreg[66] ));
 sg13g2_dfrbp_1 _13054_ (.CLK(net93),
    .RESET_B(net3463),
    .D(_00310_),
    .Q_N(_06715_),
    .Q(\u_toplayer.outreg[67] ));
 sg13g2_dfrbp_1 _13055_ (.CLK(net94),
    .RESET_B(net3478),
    .D(_00311_),
    .Q_N(_06714_),
    .Q(\u_toplayer.outreg[68] ));
 sg13g2_dfrbp_1 _13056_ (.CLK(net95),
    .RESET_B(net3481),
    .D(_00312_),
    .Q_N(_06713_),
    .Q(\u_toplayer.outreg[69] ));
 sg13g2_dfrbp_1 _13057_ (.CLK(net96),
    .RESET_B(net3481),
    .D(_00313_),
    .Q_N(_06712_),
    .Q(\u_toplayer.outreg[70] ));
 sg13g2_dfrbp_1 _13058_ (.CLK(net97),
    .RESET_B(net3467),
    .D(_00314_),
    .Q_N(_06711_),
    .Q(\u_toplayer.outreg[71] ));
 sg13g2_dfrbp_1 _13059_ (.CLK(net98),
    .RESET_B(net3465),
    .D(_00315_),
    .Q_N(_06710_),
    .Q(\u_toplayer.outreg[72] ));
 sg13g2_dfrbp_1 _13060_ (.CLK(net99),
    .RESET_B(net3463),
    .D(_00316_),
    .Q_N(_06709_),
    .Q(\u_toplayer.outreg[73] ));
 sg13g2_dfrbp_1 _13061_ (.CLK(net100),
    .RESET_B(net3463),
    .D(_00317_),
    .Q_N(_06708_),
    .Q(\u_toplayer.outreg[74] ));
 sg13g2_dfrbp_1 _13062_ (.CLK(net101),
    .RESET_B(net3463),
    .D(_00318_),
    .Q_N(_06707_),
    .Q(\u_toplayer.outreg[75] ));
 sg13g2_dfrbp_1 _13063_ (.CLK(net102),
    .RESET_B(net3478),
    .D(_00319_),
    .Q_N(_06706_),
    .Q(\u_toplayer.outreg[76] ));
 sg13g2_dfrbp_1 _13064_ (.CLK(net103),
    .RESET_B(net3466),
    .D(_00320_),
    .Q_N(_06705_),
    .Q(\u_toplayer.outreg[77] ));
 sg13g2_dfrbp_1 _13065_ (.CLK(net104),
    .RESET_B(net3466),
    .D(net389),
    .Q_N(_06704_),
    .Q(\u_toplayer.outreg[78] ));
 sg13g2_dfrbp_1 _13066_ (.CLK(net105),
    .RESET_B(net3467),
    .D(_00322_),
    .Q_N(_06703_),
    .Q(\u_toplayer.outreg[79] ));
 sg13g2_dfrbp_1 _13067_ (.CLK(net106),
    .RESET_B(net3422),
    .D(net893),
    .Q_N(_06879_),
    .Q(\u_toplayer.done_layer3 ));
 sg13g2_dfrbp_1 _13068_ (.CLK(clknet_leaf_21_clk_regs),
    .RESET_B(net3473),
    .D(_00025_),
    .Q_N(_06880_),
    .Q(\u_toplayer.u_outlayer.u_neuron.instCtrl.state[0] ));
 sg13g2_dfrbp_1 _13069_ (.CLK(clknet_leaf_21_clk_regs),
    .RESET_B(net3468),
    .D(_00026_),
    .Q_N(_00036_),
    .Q(\u_toplayer.u_outlayer.u_neuron.instCtrl.state[1] ));
 sg13g2_dfrbp_1 _13070_ (.CLK(clknet_leaf_21_clk_regs),
    .RESET_B(net3476),
    .D(_00027_),
    .Q_N(_00035_),
    .Q(\u_toplayer.u_outlayer.u_neuron.instCtrl.state[2] ));
 sg13g2_dfrbp_1 _13071_ (.CLK(clknet_leaf_21_clk_regs),
    .RESET_B(net3476),
    .D(net959),
    .Q_N(_06702_),
    .Q(\u_toplayer.u_outlayer.u_neuron.instCtrl.state[3] ));
 sg13g2_dfrbp_1 _13072_ (.CLK(clknet_leaf_48_clk_regs),
    .RESET_B(net3561),
    .D(_00324_),
    .Q_N(_06701_),
    .Q(\u_toplayer.u_layer3.u_neuron.din[0] ));
 sg13g2_dfrbp_1 _13073_ (.CLK(clknet_leaf_46_clk_regs),
    .RESET_B(net3561),
    .D(_00325_),
    .Q_N(_06700_),
    .Q(\u_toplayer.u_layer3.u_neuron.din[1] ));
 sg13g2_dfrbp_1 _13074_ (.CLK(clknet_leaf_46_clk_regs),
    .RESET_B(net3561),
    .D(_00326_),
    .Q_N(_06699_),
    .Q(\u_toplayer.u_layer3.u_neuron.din[2] ));
 sg13g2_dfrbp_1 _13075_ (.CLK(clknet_leaf_46_clk_regs),
    .RESET_B(net3561),
    .D(_00327_),
    .Q_N(_06698_),
    .Q(\u_toplayer.u_layer3.u_neuron.din[3] ));
 sg13g2_dfrbp_1 _13076_ (.CLK(clknet_leaf_46_clk_regs),
    .RESET_B(net3561),
    .D(_00328_),
    .Q_N(_06697_),
    .Q(\u_toplayer.u_layer3.u_neuron.din[4] ));
 sg13g2_dfrbp_1 _13077_ (.CLK(clknet_leaf_90_clk_regs),
    .RESET_B(net3515),
    .D(_00329_),
    .Q_N(_06696_),
    .Q(\u_toplayer.u_layer3.u_neuron.din[5] ));
 sg13g2_dfrbp_1 _13078_ (.CLK(clknet_leaf_87_clk_regs),
    .RESET_B(net3511),
    .D(_00330_),
    .Q_N(_06695_),
    .Q(\u_toplayer.u_layer3.u_neuron.din[6] ));
 sg13g2_dfrbp_1 _13079_ (.CLK(clknet_leaf_88_clk_regs),
    .RESET_B(net3510),
    .D(_00331_),
    .Q_N(_06694_),
    .Q(\u_toplayer.u_layer3.u_neuron.din[7] ));
 sg13g2_dfrbp_1 _13080_ (.CLK(clknet_leaf_18_clk_regs),
    .RESET_B(net3482),
    .D(_00332_),
    .Q_N(_06693_),
    .Q(\u_toplayer.u_layer3.sum[0] ));
 sg13g2_dfrbp_1 _13081_ (.CLK(clknet_leaf_18_clk_regs),
    .RESET_B(net3479),
    .D(net1027),
    .Q_N(_06692_),
    .Q(\u_toplayer.u_layer3.sum[1] ));
 sg13g2_dfrbp_1 _13082_ (.CLK(clknet_leaf_18_clk_regs),
    .RESET_B(net3478),
    .D(net1054),
    .Q_N(_06691_),
    .Q(\u_toplayer.u_layer3.sum[2] ));
 sg13g2_dfrbp_1 _13083_ (.CLK(clknet_leaf_18_clk_regs),
    .RESET_B(net3478),
    .D(net1077),
    .Q_N(_06690_),
    .Q(\u_toplayer.u_layer3.sum[3] ));
 sg13g2_dfrbp_1 _13084_ (.CLK(clknet_leaf_18_clk_regs),
    .RESET_B(net3478),
    .D(net1031),
    .Q_N(_06689_),
    .Q(\u_toplayer.u_layer3.sum[4] ));
 sg13g2_dfrbp_1 _13085_ (.CLK(clknet_leaf_19_clk_regs),
    .RESET_B(net3482),
    .D(net1102),
    .Q_N(_06688_),
    .Q(\u_toplayer.u_layer3.sum[5] ));
 sg13g2_dfrbp_1 _13086_ (.CLK(clknet_leaf_19_clk_regs),
    .RESET_B(net3480),
    .D(net1045),
    .Q_N(_06687_),
    .Q(\u_toplayer.u_layer3.sum[6] ));
 sg13g2_dfrbp_1 _13087_ (.CLK(clknet_leaf_31_clk_regs),
    .RESET_B(net3480),
    .D(net1033),
    .Q_N(_06686_),
    .Q(\u_toplayer.u_layer3.sum[7] ));
 sg13g2_dfrbp_1 _13088_ (.CLK(net107),
    .RESET_B(net3423),
    .D(net841),
    .Q_N(_06685_),
    .Q(\u_toplayer.u_layer3.stateout[0] ));
 sg13g2_dfrbp_1 _13089_ (.CLK(net108),
    .RESET_B(net3423),
    .D(_00341_),
    .Q_N(_06684_),
    .Q(\u_toplayer.u_layer3.stateout[1] ));
 sg13g2_dfrbp_1 _13090_ (.CLK(net109),
    .RESET_B(net3422),
    .D(net941),
    .Q_N(_06683_),
    .Q(\u_toplayer.u_layer3.stateout[2] ));
 sg13g2_dfrbp_1 _13091_ (.CLK(net110),
    .RESET_B(net3426),
    .D(net864),
    .Q_N(_06682_),
    .Q(\u_toplayer.u_layer3.stateout[3] ));
 sg13g2_dfrbp_1 _13092_ (.CLK(net111),
    .RESET_B(net3417),
    .D(_00344_),
    .Q_N(_06681_),
    .Q(\u_toplayer.u_layer3.stateout[4] ));
 sg13g2_dfrbp_1 _13093_ (.CLK(net112),
    .RESET_B(net3422),
    .D(net896),
    .Q_N(_06680_),
    .Q(\u_toplayer.u_layer3.stateout[5] ));
 sg13g2_dfrbp_1 _13094_ (.CLK(net113),
    .RESET_B(net3417),
    .D(_00346_),
    .Q_N(_06679_),
    .Q(\u_toplayer.u_layer3.stateout[6] ));
 sg13g2_dfrbp_1 _13095_ (.CLK(net114),
    .RESET_B(net3417),
    .D(_00347_),
    .Q_N(_06678_),
    .Q(\u_toplayer.u_layer3.stateout[7] ));
 sg13g2_dfrbp_1 _13096_ (.CLK(net115),
    .RESET_B(net3423),
    .D(net117),
    .Q_N(_00033_),
    .Q(\u_toplayer.u_layer3.stateout[8] ));
 sg13g2_dfrbp_1 _13097_ (.CLK(clknet_leaf_18_clk_regs),
    .RESET_B(net3482),
    .D(net1048),
    .Q_N(_06677_),
    .Q(\u_toplayer.u_layer3.u_neuron.acc[0] ));
 sg13g2_dfrbp_1 _13098_ (.CLK(clknet_leaf_18_clk_regs),
    .RESET_B(net3482),
    .D(net1087),
    .Q_N(_06676_),
    .Q(\u_toplayer.u_layer3.u_neuron.acc[1] ));
 sg13g2_dfrbp_1 _13099_ (.CLK(clknet_leaf_18_clk_regs),
    .RESET_B(net3484),
    .D(_00351_),
    .Q_N(_06675_),
    .Q(\u_toplayer.u_layer3.u_neuron.acc[2] ));
 sg13g2_dfrbp_1 _13100_ (.CLK(clknet_leaf_32_clk_regs),
    .RESET_B(net3484),
    .D(_00352_),
    .Q_N(_06674_),
    .Q(\u_toplayer.u_layer3.u_neuron.acc[3] ));
 sg13g2_dfrbp_1 _13101_ (.CLK(clknet_leaf_32_clk_regs),
    .RESET_B(net3481),
    .D(_00353_),
    .Q_N(_06673_),
    .Q(\u_toplayer.u_layer3.u_neuron.acc[4] ));
 sg13g2_dfrbp_1 _13102_ (.CLK(clknet_leaf_34_clk_regs),
    .RESET_B(net3483),
    .D(_00354_),
    .Q_N(_06672_),
    .Q(\u_toplayer.u_layer3.u_neuron.acc[5] ));
 sg13g2_dfrbp_1 _13103_ (.CLK(clknet_leaf_33_clk_regs),
    .RESET_B(net3483),
    .D(_00355_),
    .Q_N(_06671_),
    .Q(\u_toplayer.u_layer3.u_neuron.acc[6] ));
 sg13g2_dfrbp_1 _13104_ (.CLK(clknet_leaf_33_clk_regs),
    .RESET_B(net3484),
    .D(_00356_),
    .Q_N(_06670_),
    .Q(\u_toplayer.u_layer3.u_neuron.acc[7] ));
 sg13g2_dfrbp_1 _13105_ (.CLK(clknet_leaf_36_clk_regs),
    .RESET_B(net3483),
    .D(_00357_),
    .Q_N(_06669_),
    .Q(\u_toplayer.u_layer3.u_neuron.acc[8] ));
 sg13g2_dfrbp_1 _13106_ (.CLK(clknet_leaf_37_clk_regs),
    .RESET_B(net3549),
    .D(_00358_),
    .Q_N(_06668_),
    .Q(\u_toplayer.u_layer3.u_neuron.acc[9] ));
 sg13g2_dfrbp_1 _13107_ (.CLK(clknet_leaf_41_clk_regs),
    .RESET_B(net3485),
    .D(_00359_),
    .Q_N(_06667_),
    .Q(\u_toplayer.u_layer3.u_neuron.acc[10] ));
 sg13g2_dfrbp_1 _13108_ (.CLK(clknet_leaf_36_clk_regs),
    .RESET_B(net3553),
    .D(_00360_),
    .Q_N(_06666_),
    .Q(\u_toplayer.u_layer3.u_neuron.acc[11] ));
 sg13g2_dfrbp_1 _13109_ (.CLK(clknet_leaf_33_clk_regs),
    .RESET_B(net3486),
    .D(_00361_),
    .Q_N(_06665_),
    .Q(\u_toplayer.u_layer3.u_neuron.acc[12] ));
 sg13g2_dfrbp_1 _13110_ (.CLK(clknet_leaf_36_clk_regs),
    .RESET_B(net3483),
    .D(_00362_),
    .Q_N(_06664_),
    .Q(\u_toplayer.u_layer3.u_neuron.acc[13] ));
 sg13g2_dfrbp_1 _13111_ (.CLK(clknet_leaf_33_clk_regs),
    .RESET_B(net3483),
    .D(_00363_),
    .Q_N(_06663_),
    .Q(\u_toplayer.u_layer3.u_neuron.acc[14] ));
 sg13g2_dfrbp_1 _13112_ (.CLK(clknet_leaf_33_clk_regs),
    .RESET_B(net3483),
    .D(_00364_),
    .Q_N(_06662_),
    .Q(\u_toplayer.u_layer3.u_neuron.acc[15] ));
 sg13g2_dfrbp_1 _13113_ (.CLK(clknet_leaf_30_clk_regs),
    .RESET_B(net3485),
    .D(_00365_),
    .Q_N(_06661_),
    .Q(\u_toplayer.u_layer3.u_neuron.acc[16] ));
 sg13g2_dfrbp_1 _13114_ (.CLK(clknet_leaf_30_clk_regs),
    .RESET_B(net3486),
    .D(_00366_),
    .Q_N(_06660_),
    .Q(\u_toplayer.u_layer3.u_neuron.acc[17] ));
 sg13g2_dfrbp_1 _13115_ (.CLK(clknet_leaf_30_clk_regs),
    .RESET_B(net3486),
    .D(_00367_),
    .Q_N(_06659_),
    .Q(\u_toplayer.u_layer3.u_neuron.acc[18] ));
 sg13g2_dfrbp_1 _13116_ (.CLK(clknet_leaf_30_clk_regs),
    .RESET_B(net3485),
    .D(_00368_),
    .Q_N(_06658_),
    .Q(\u_toplayer.u_layer3.u_neuron.acc[19] ));
 sg13g2_dfrbp_1 _13117_ (.CLK(clknet_leaf_31_clk_regs),
    .RESET_B(net3485),
    .D(_00369_),
    .Q_N(_06657_),
    .Q(\u_toplayer.u_layer3.u_neuron.acc[20] ));
 sg13g2_dfrbp_1 _13118_ (.CLK(clknet_leaf_31_clk_regs),
    .RESET_B(net3481),
    .D(_00370_),
    .Q_N(_06656_),
    .Q(\u_toplayer.u_layer3.u_neuron.acc[21] ));
 sg13g2_dfrbp_1 _13119_ (.CLK(clknet_leaf_31_clk_regs),
    .RESET_B(net3481),
    .D(_00371_),
    .Q_N(_06655_),
    .Q(\u_toplayer.u_layer3.u_neuron.acc[22] ));
 sg13g2_dfrbp_1 _13120_ (.CLK(clknet_leaf_31_clk_regs),
    .RESET_B(net3481),
    .D(_00372_),
    .Q_N(_06654_),
    .Q(\u_toplayer.u_layer3.u_neuron.acc[23] ));
 sg13g2_dfrbp_1 _13121_ (.CLK(clknet_leaf_77_clk_regs),
    .RESET_B(net3497),
    .D(net735),
    .Q_N(_00051_),
    .Q(\u_toplayer.u_layer2.neuron_index[0] ));
 sg13g2_dfrbp_1 _13122_ (.CLK(clknet_leaf_77_clk_regs),
    .RESET_B(net3498),
    .D(_00374_),
    .Q_N(_06653_),
    .Q(\u_toplayer.u_layer2.neuron_index[1] ));
 sg13g2_dfrbp_1 _13123_ (.CLK(clknet_leaf_76_clk_regs),
    .RESET_B(net3498),
    .D(_00375_),
    .Q_N(_06652_),
    .Q(\u_toplayer.u_layer2.neuron_index[2] ));
 sg13g2_dfrbp_1 _13124_ (.CLK(clknet_leaf_77_clk_regs),
    .RESET_B(net3497),
    .D(_00376_),
    .Q_N(_06651_),
    .Q(\u_toplayer.u_layer2.neuron_index[3] ));
 sg13g2_dfrbp_1 _13125_ (.CLK(clknet_leaf_77_clk_regs),
    .RESET_B(net3497),
    .D(_00377_),
    .Q_N(_06650_),
    .Q(\u_toplayer.u_layer2.neuron_index[4] ));
 sg13g2_dfrbp_1 _13126_ (.CLK(clknet_leaf_77_clk_regs),
    .RESET_B(net3500),
    .D(net983),
    .Q_N(_06649_),
    .Q(\u_toplayer.u_layer2.neuron_index[5] ));
 sg13g2_dfrbp_1 _13127_ (.CLK(clknet_leaf_39_clk_regs),
    .RESET_B(net3557),
    .D(_00379_),
    .Q_N(_06648_),
    .Q(\u_toplayer.u_layer1.u_neuron.mult[0] ));
 sg13g2_dfrbp_1 _13128_ (.CLK(clknet_leaf_36_clk_regs),
    .RESET_B(net3553),
    .D(_00380_),
    .Q_N(_06647_),
    .Q(\u_toplayer.u_layer1.u_neuron.mult[1] ));
 sg13g2_dfrbp_1 _13129_ (.CLK(clknet_leaf_41_clk_regs),
    .RESET_B(net3553),
    .D(_00381_),
    .Q_N(_06646_),
    .Q(\u_toplayer.u_layer1.u_neuron.mult[2] ));
 sg13g2_dfrbp_1 _13130_ (.CLK(clknet_leaf_40_clk_regs),
    .RESET_B(net3553),
    .D(_00382_),
    .Q_N(_06645_),
    .Q(\u_toplayer.u_layer1.u_neuron.mult[3] ));
 sg13g2_dfrbp_1 _13131_ (.CLK(clknet_leaf_41_clk_regs),
    .RESET_B(net3553),
    .D(_00383_),
    .Q_N(_06644_),
    .Q(\u_toplayer.u_layer1.u_neuron.mult[4] ));
 sg13g2_dfrbp_1 _13132_ (.CLK(clknet_leaf_41_clk_regs),
    .RESET_B(net3554),
    .D(_00384_),
    .Q_N(_06643_),
    .Q(\u_toplayer.u_layer1.u_neuron.mult[5] ));
 sg13g2_dfrbp_1 _13133_ (.CLK(clknet_leaf_40_clk_regs),
    .RESET_B(net3554),
    .D(_00385_),
    .Q_N(_06642_),
    .Q(\u_toplayer.u_layer1.u_neuron.mult[6] ));
 sg13g2_dfrbp_1 _13134_ (.CLK(clknet_leaf_40_clk_regs),
    .RESET_B(net3553),
    .D(_00386_),
    .Q_N(_06641_),
    .Q(\u_toplayer.u_layer1.u_neuron.mult[7] ));
 sg13g2_dfrbp_1 _13135_ (.CLK(clknet_leaf_42_clk_regs),
    .RESET_B(net3553),
    .D(_00387_),
    .Q_N(_06640_),
    .Q(\u_toplayer.u_layer1.u_neuron.mult[8] ));
 sg13g2_dfrbp_1 _13136_ (.CLK(clknet_leaf_42_clk_regs),
    .RESET_B(net3555),
    .D(_00388_),
    .Q_N(_06639_),
    .Q(\u_toplayer.u_layer1.u_neuron.mult[9] ));
 sg13g2_dfrbp_1 _13137_ (.CLK(clknet_leaf_42_clk_regs),
    .RESET_B(net3555),
    .D(_00389_),
    .Q_N(_06638_),
    .Q(\u_toplayer.u_layer1.u_neuron.mult[10] ));
 sg13g2_dfrbp_1 _13138_ (.CLK(clknet_leaf_42_clk_regs),
    .RESET_B(net3555),
    .D(_00390_),
    .Q_N(_06637_),
    .Q(\u_toplayer.u_layer1.u_neuron.mult[11] ));
 sg13g2_dfrbp_1 _13139_ (.CLK(clknet_leaf_43_clk_regs),
    .RESET_B(net3559),
    .D(_00391_),
    .Q_N(_06636_),
    .Q(\u_toplayer.u_layer1.u_neuron.mult[12] ));
 sg13g2_dfrbp_1 _13140_ (.CLK(clknet_leaf_43_clk_regs),
    .RESET_B(net3559),
    .D(_00392_),
    .Q_N(_06635_),
    .Q(\u_toplayer.u_layer1.u_neuron.mult[13] ));
 sg13g2_dfrbp_1 _13141_ (.CLK(clknet_leaf_42_clk_regs),
    .RESET_B(net3559),
    .D(_00393_),
    .Q_N(_06634_),
    .Q(\u_toplayer.u_layer1.u_neuron.mult[14] ));
 sg13g2_dfrbp_1 _13142_ (.CLK(clknet_leaf_42_clk_regs),
    .RESET_B(net3559),
    .D(_00394_),
    .Q_N(_06633_),
    .Q(\u_toplayer.u_layer1.u_neuron.mult[15] ));
 sg13g2_dfrbp_1 _13143_ (.CLK(clknet_leaf_74_clk_regs),
    .RESET_B(net3521),
    .D(_00395_),
    .Q_N(_06632_),
    .Q(\u_toplayer.reg_layer2[0] ));
 sg13g2_dfrbp_1 _13144_ (.CLK(clknet_leaf_85_clk_regs),
    .RESET_B(net3523),
    .D(_00396_),
    .Q_N(_06631_),
    .Q(\u_toplayer.reg_layer2[1] ));
 sg13g2_dfrbp_1 _13145_ (.CLK(clknet_leaf_74_clk_regs),
    .RESET_B(net3522),
    .D(_00397_),
    .Q_N(_06630_),
    .Q(\u_toplayer.reg_layer2[2] ));
 sg13g2_dfrbp_1 _13146_ (.CLK(clknet_leaf_65_clk_regs),
    .RESET_B(net3521),
    .D(_00398_),
    .Q_N(_06629_),
    .Q(\u_toplayer.reg_layer2[3] ));
 sg13g2_dfrbp_1 _13147_ (.CLK(clknet_leaf_86_clk_regs),
    .RESET_B(net3523),
    .D(_00399_),
    .Q_N(_06628_),
    .Q(\u_toplayer.reg_layer2[4] ));
 sg13g2_dfrbp_1 _13148_ (.CLK(clknet_leaf_74_clk_regs),
    .RESET_B(net3521),
    .D(_00400_),
    .Q_N(_06627_),
    .Q(\u_toplayer.reg_layer2[5] ));
 sg13g2_dfrbp_1 _13149_ (.CLK(clknet_leaf_75_clk_regs),
    .RESET_B(net3521),
    .D(_00401_),
    .Q_N(_06626_),
    .Q(\u_toplayer.reg_layer2[6] ));
 sg13g2_dfrbp_1 _13150_ (.CLK(clknet_leaf_74_clk_regs),
    .RESET_B(net3517),
    .D(_00402_),
    .Q_N(_06625_),
    .Q(\u_toplayer.reg_layer2[7] ));
 sg13g2_dfrbp_1 _13151_ (.CLK(clknet_leaf_75_clk_regs),
    .RESET_B(net3521),
    .D(_00403_),
    .Q_N(_06624_),
    .Q(\u_toplayer.reg_layer2[8] ));
 sg13g2_dfrbp_1 _13152_ (.CLK(clknet_leaf_85_clk_regs),
    .RESET_B(net3502),
    .D(_00404_),
    .Q_N(_06623_),
    .Q(\u_toplayer.reg_layer2[9] ));
 sg13g2_dfrbp_1 _13153_ (.CLK(clknet_leaf_74_clk_regs),
    .RESET_B(net3521),
    .D(_00405_),
    .Q_N(_06622_),
    .Q(\u_toplayer.reg_layer2[10] ));
 sg13g2_dfrbp_1 _13154_ (.CLK(clknet_leaf_85_clk_regs),
    .RESET_B(net3523),
    .D(_00406_),
    .Q_N(_06621_),
    .Q(\u_toplayer.reg_layer2[11] ));
 sg13g2_dfrbp_1 _13155_ (.CLK(clknet_leaf_86_clk_regs),
    .RESET_B(net3523),
    .D(net847),
    .Q_N(_06620_),
    .Q(\u_toplayer.reg_layer2[12] ));
 sg13g2_dfrbp_1 _13156_ (.CLK(clknet_leaf_85_clk_regs),
    .RESET_B(net3503),
    .D(_00408_),
    .Q_N(_06619_),
    .Q(\u_toplayer.reg_layer2[13] ));
 sg13g2_dfrbp_1 _13157_ (.CLK(clknet_leaf_75_clk_regs),
    .RESET_B(net3502),
    .D(_00409_),
    .Q_N(_06618_),
    .Q(\u_toplayer.reg_layer2[14] ));
 sg13g2_dfrbp_1 _13158_ (.CLK(clknet_leaf_76_clk_regs),
    .RESET_B(net3498),
    .D(_00410_),
    .Q_N(_06617_),
    .Q(\u_toplayer.reg_layer2[15] ));
 sg13g2_dfrbp_1 _13159_ (.CLK(clknet_leaf_78_clk_regs),
    .RESET_B(net3497),
    .D(_00411_),
    .Q_N(_06616_),
    .Q(\u_toplayer.reg_layer2[16] ));
 sg13g2_dfrbp_1 _13160_ (.CLK(clknet_leaf_83_clk_regs),
    .RESET_B(net3501),
    .D(_00412_),
    .Q_N(_06615_),
    .Q(\u_toplayer.reg_layer2[17] ));
 sg13g2_dfrbp_1 _13161_ (.CLK(clknet_leaf_84_clk_regs),
    .RESET_B(net3501),
    .D(_00413_),
    .Q_N(_06614_),
    .Q(\u_toplayer.reg_layer2[18] ));
 sg13g2_dfrbp_1 _13162_ (.CLK(clknet_leaf_83_clk_regs),
    .RESET_B(net3495),
    .D(_00414_),
    .Q_N(_06613_),
    .Q(\u_toplayer.reg_layer2[19] ));
 sg13g2_dfrbp_1 _13163_ (.CLK(clknet_leaf_88_clk_regs),
    .RESET_B(net3501),
    .D(_00415_),
    .Q_N(_06612_),
    .Q(\u_toplayer.reg_layer2[20] ));
 sg13g2_dfrbp_1 _13164_ (.CLK(clknet_leaf_84_clk_regs),
    .RESET_B(net3495),
    .D(_00416_),
    .Q_N(_06611_),
    .Q(\u_toplayer.reg_layer2[21] ));
 sg13g2_dfrbp_1 _13165_ (.CLK(clknet_leaf_81_clk_regs),
    .RESET_B(net3495),
    .D(_00417_),
    .Q_N(_06610_),
    .Q(\u_toplayer.reg_layer2[22] ));
 sg13g2_dfrbp_1 _13166_ (.CLK(clknet_leaf_78_clk_regs),
    .RESET_B(net3497),
    .D(_00418_),
    .Q_N(_06609_),
    .Q(\u_toplayer.reg_layer2[23] ));
 sg13g2_dfrbp_1 _13167_ (.CLK(clknet_leaf_78_clk_regs),
    .RESET_B(net3497),
    .D(_00419_),
    .Q_N(_06608_),
    .Q(\u_toplayer.reg_layer2[24] ));
 sg13g2_dfrbp_1 _13168_ (.CLK(clknet_leaf_83_clk_regs),
    .RESET_B(net3501),
    .D(net481),
    .Q_N(_06607_),
    .Q(\u_toplayer.reg_layer2[25] ));
 sg13g2_dfrbp_1 _13169_ (.CLK(clknet_leaf_84_clk_regs),
    .RESET_B(net3501),
    .D(_00421_),
    .Q_N(_06606_),
    .Q(\u_toplayer.reg_layer2[26] ));
 sg13g2_dfrbp_1 _13170_ (.CLK(clknet_leaf_83_clk_regs),
    .RESET_B(net3496),
    .D(_00422_),
    .Q_N(_06605_),
    .Q(\u_toplayer.reg_layer2[27] ));
 sg13g2_dfrbp_1 _13171_ (.CLK(clknet_leaf_83_clk_regs),
    .RESET_B(net3501),
    .D(_00423_),
    .Q_N(_06604_),
    .Q(\u_toplayer.reg_layer2[28] ));
 sg13g2_dfrbp_1 _13172_ (.CLK(clknet_leaf_82_clk_regs),
    .RESET_B(net3495),
    .D(_00424_),
    .Q_N(_06603_),
    .Q(\u_toplayer.reg_layer2[29] ));
 sg13g2_dfrbp_1 _13173_ (.CLK(clknet_leaf_80_clk_regs),
    .RESET_B(net3491),
    .D(_00425_),
    .Q_N(_06602_),
    .Q(\u_toplayer.reg_layer2[30] ));
 sg13g2_dfrbp_1 _13174_ (.CLK(clknet_leaf_81_clk_regs),
    .RESET_B(net3491),
    .D(_00426_),
    .Q_N(_06601_),
    .Q(\u_toplayer.reg_layer2[31] ));
 sg13g2_dfrbp_1 _13175_ (.CLK(clknet_leaf_70_clk_regs),
    .RESET_B(net3524),
    .D(_00427_),
    .Q_N(_06600_),
    .Q(\u_toplayer.reg_layer2[32] ));
 sg13g2_dfrbp_1 _13176_ (.CLK(clknet_leaf_66_clk_regs),
    .RESET_B(net3527),
    .D(_00428_),
    .Q_N(_06599_),
    .Q(\u_toplayer.reg_layer2[33] ));
 sg13g2_dfrbp_1 _13177_ (.CLK(clknet_leaf_69_clk_regs),
    .RESET_B(net3531),
    .D(net838),
    .Q_N(_06598_),
    .Q(\u_toplayer.reg_layer2[34] ));
 sg13g2_dfrbp_1 _13178_ (.CLK(clknet_leaf_68_clk_regs),
    .RESET_B(net3527),
    .D(net686),
    .Q_N(_06597_),
    .Q(\u_toplayer.reg_layer2[35] ));
 sg13g2_dfrbp_1 _13179_ (.CLK(clknet_leaf_70_clk_regs),
    .RESET_B(net3526),
    .D(_00431_),
    .Q_N(_06596_),
    .Q(\u_toplayer.reg_layer2[36] ));
 sg13g2_dfrbp_1 _13180_ (.CLK(clknet_leaf_73_clk_regs),
    .RESET_B(net3525),
    .D(net527),
    .Q_N(_06595_),
    .Q(\u_toplayer.reg_layer2[37] ));
 sg13g2_dfrbp_1 _13181_ (.CLK(clknet_leaf_71_clk_regs),
    .RESET_B(net3518),
    .D(net173),
    .Q_N(_06594_),
    .Q(\u_toplayer.reg_layer2[38] ));
 sg13g2_dfrbp_1 _13182_ (.CLK(clknet_leaf_71_clk_regs),
    .RESET_B(net3518),
    .D(net743),
    .Q_N(_06593_),
    .Q(\u_toplayer.reg_layer2[39] ));
 sg13g2_dfrbp_1 _13183_ (.CLK(clknet_leaf_70_clk_regs),
    .RESET_B(net3524),
    .D(_00435_),
    .Q_N(_06592_),
    .Q(\u_toplayer.reg_layer2[40] ));
 sg13g2_dfrbp_1 _13184_ (.CLK(clknet_leaf_67_clk_regs),
    .RESET_B(net3527),
    .D(_00436_),
    .Q_N(_06591_),
    .Q(\u_toplayer.reg_layer2[41] ));
 sg13g2_dfrbp_1 _13185_ (.CLK(clknet_leaf_69_clk_regs),
    .RESET_B(net3531),
    .D(net843),
    .Q_N(_06590_),
    .Q(\u_toplayer.reg_layer2[42] ));
 sg13g2_dfrbp_1 _13186_ (.CLK(clknet_leaf_68_clk_regs),
    .RESET_B(net3530),
    .D(net456),
    .Q_N(_06589_),
    .Q(\u_toplayer.reg_layer2[43] ));
 sg13g2_dfrbp_1 _13187_ (.CLK(clknet_leaf_70_clk_regs),
    .RESET_B(net3526),
    .D(_00439_),
    .Q_N(_06588_),
    .Q(\u_toplayer.reg_layer2[44] ));
 sg13g2_dfrbp_1 _13188_ (.CLK(clknet_leaf_69_clk_regs),
    .RESET_B(net3525),
    .D(net454),
    .Q_N(_06587_),
    .Q(\u_toplayer.reg_layer2[45] ));
 sg13g2_dfrbp_1 _13189_ (.CLK(clknet_leaf_70_clk_regs),
    .RESET_B(net3524),
    .D(net790),
    .Q_N(_06586_),
    .Q(\u_toplayer.reg_layer2[46] ));
 sg13g2_dfrbp_1 _13190_ (.CLK(clknet_leaf_71_clk_regs),
    .RESET_B(net3524),
    .D(net189),
    .Q_N(_06585_),
    .Q(\u_toplayer.reg_layer2[47] ));
 sg13g2_dfrbp_1 _13191_ (.CLK(clknet_leaf_71_clk_regs),
    .RESET_B(net3518),
    .D(net525),
    .Q_N(_06584_),
    .Q(\u_toplayer.reg_layer2[48] ));
 sg13g2_dfrbp_1 _13192_ (.CLK(clknet_leaf_66_clk_regs),
    .RESET_B(net3522),
    .D(net652),
    .Q_N(_06583_),
    .Q(\u_toplayer.reg_layer2[49] ));
 sg13g2_dfrbp_1 _13193_ (.CLK(clknet_leaf_73_clk_regs),
    .RESET_B(net3516),
    .D(net232),
    .Q_N(_06582_),
    .Q(\u_toplayer.reg_layer2[50] ));
 sg13g2_dfrbp_1 _13194_ (.CLK(clknet_leaf_67_clk_regs),
    .RESET_B(net3522),
    .D(_00446_),
    .Q_N(_06581_),
    .Q(\u_toplayer.reg_layer2[51] ));
 sg13g2_dfrbp_1 _13195_ (.CLK(clknet_leaf_73_clk_regs),
    .RESET_B(net3519),
    .D(net629),
    .Q_N(_06580_),
    .Q(\u_toplayer.reg_layer2[52] ));
 sg13g2_dfrbp_1 _13196_ (.CLK(clknet_leaf_72_clk_regs),
    .RESET_B(net3517),
    .D(net566),
    .Q_N(_06579_),
    .Q(\u_toplayer.reg_layer2[53] ));
 sg13g2_dfrbp_1 _13197_ (.CLK(clknet_leaf_77_clk_regs),
    .RESET_B(net3498),
    .D(_00449_),
    .Q_N(_06578_),
    .Q(\u_toplayer.reg_layer2[54] ));
 sg13g2_dfrbp_1 _13198_ (.CLK(clknet_leaf_72_clk_regs),
    .RESET_B(net3516),
    .D(_00450_),
    .Q_N(_06577_),
    .Q(\u_toplayer.reg_layer2[55] ));
 sg13g2_dfrbp_1 _13199_ (.CLK(clknet_leaf_71_clk_regs),
    .RESET_B(net3518),
    .D(_00451_),
    .Q_N(_06576_),
    .Q(\u_toplayer.reg_layer2[56] ));
 sg13g2_dfrbp_1 _13200_ (.CLK(clknet_leaf_74_clk_regs),
    .RESET_B(net3521),
    .D(_00452_),
    .Q_N(_06575_),
    .Q(\u_toplayer.reg_layer2[57] ));
 sg13g2_dfrbp_1 _13201_ (.CLK(clknet_leaf_72_clk_regs),
    .RESET_B(net3516),
    .D(_00453_),
    .Q_N(_06574_),
    .Q(\u_toplayer.reg_layer2[58] ));
 sg13g2_dfrbp_1 _13202_ (.CLK(clknet_leaf_66_clk_regs),
    .RESET_B(net3522),
    .D(_00454_),
    .Q_N(_06573_),
    .Q(\u_toplayer.reg_layer2[59] ));
 sg13g2_dfrbp_1 _13203_ (.CLK(clknet_leaf_73_clk_regs),
    .RESET_B(net3518),
    .D(_00455_),
    .Q_N(_06572_),
    .Q(\u_toplayer.reg_layer2[60] ));
 sg13g2_dfrbp_1 _13204_ (.CLK(clknet_leaf_76_clk_regs),
    .RESET_B(net3499),
    .D(_00456_),
    .Q_N(_06571_),
    .Q(\u_toplayer.reg_layer2[61] ));
 sg13g2_dfrbp_1 _13205_ (.CLK(clknet_leaf_76_clk_regs),
    .RESET_B(net3498),
    .D(_00457_),
    .Q_N(_06570_),
    .Q(\u_toplayer.reg_layer2[62] ));
 sg13g2_dfrbp_1 _13206_ (.CLK(clknet_leaf_72_clk_regs),
    .RESET_B(net3516),
    .D(_00458_),
    .Q_N(_06569_),
    .Q(\u_toplayer.reg_layer2[63] ));
 sg13g2_dfrbp_1 _13207_ (.CLK(clknet_leaf_56_clk_regs),
    .RESET_B(net3538),
    .D(_00459_),
    .Q_N(_06568_),
    .Q(\u_toplayer.reg_layer2[64] ));
 sg13g2_dfrbp_1 _13208_ (.CLK(clknet_leaf_52_clk_regs),
    .RESET_B(net3537),
    .D(_00460_),
    .Q_N(_06567_),
    .Q(\u_toplayer.reg_layer2[65] ));
 sg13g2_dfrbp_1 _13209_ (.CLK(clknet_leaf_57_clk_regs),
    .RESET_B(net3538),
    .D(_00461_),
    .Q_N(_06566_),
    .Q(\u_toplayer.reg_layer2[66] ));
 sg13g2_dfrbp_1 _13210_ (.CLK(clknet_leaf_57_clk_regs),
    .RESET_B(net3540),
    .D(_00462_),
    .Q_N(_06565_),
    .Q(\u_toplayer.reg_layer2[67] ));
 sg13g2_dfrbp_1 _13211_ (.CLK(clknet_leaf_55_clk_regs),
    .RESET_B(net3534),
    .D(_00463_),
    .Q_N(_06564_),
    .Q(\u_toplayer.reg_layer2[68] ));
 sg13g2_dfrbp_1 _13212_ (.CLK(clknet_leaf_57_clk_regs),
    .RESET_B(net3537),
    .D(_00464_),
    .Q_N(_06563_),
    .Q(\u_toplayer.reg_layer2[69] ));
 sg13g2_dfrbp_1 _13213_ (.CLK(clknet_leaf_55_clk_regs),
    .RESET_B(net3535),
    .D(_00465_),
    .Q_N(_06562_),
    .Q(\u_toplayer.reg_layer2[70] ));
 sg13g2_dfrbp_1 _13214_ (.CLK(clknet_leaf_55_clk_regs),
    .RESET_B(net3532),
    .D(_00466_),
    .Q_N(_06561_),
    .Q(\u_toplayer.reg_layer2[71] ));
 sg13g2_dfrbp_1 _13215_ (.CLK(clknet_leaf_56_clk_regs),
    .RESET_B(net3538),
    .D(net439),
    .Q_N(_06560_),
    .Q(\u_toplayer.reg_layer2[72] ));
 sg13g2_dfrbp_1 _13216_ (.CLK(clknet_leaf_57_clk_regs),
    .RESET_B(net3539),
    .D(net754),
    .Q_N(_06559_),
    .Q(\u_toplayer.reg_layer2[73] ));
 sg13g2_dfrbp_1 _13217_ (.CLK(clknet_leaf_58_clk_regs),
    .RESET_B(net3539),
    .D(net497),
    .Q_N(_06558_),
    .Q(\u_toplayer.reg_layer2[74] ));
 sg13g2_dfrbp_1 _13218_ (.CLK(clknet_leaf_58_clk_regs),
    .RESET_B(net3539),
    .D(_00470_),
    .Q_N(_06557_),
    .Q(\u_toplayer.reg_layer2[75] ));
 sg13g2_dfrbp_1 _13219_ (.CLK(clknet_leaf_64_clk_regs),
    .RESET_B(net3534),
    .D(_00471_),
    .Q_N(_06556_),
    .Q(\u_toplayer.reg_layer2[76] ));
 sg13g2_dfrbp_1 _13220_ (.CLK(clknet_leaf_59_clk_regs),
    .RESET_B(net3538),
    .D(net666),
    .Q_N(_06555_),
    .Q(\u_toplayer.reg_layer2[77] ));
 sg13g2_dfrbp_1 _13221_ (.CLK(clknet_leaf_55_clk_regs),
    .RESET_B(net3534),
    .D(net340),
    .Q_N(_06554_),
    .Q(\u_toplayer.reg_layer2[78] ));
 sg13g2_dfrbp_1 _13222_ (.CLK(clknet_leaf_65_clk_regs),
    .RESET_B(net3534),
    .D(net705),
    .Q_N(_06553_),
    .Q(\u_toplayer.reg_layer2[79] ));
 sg13g2_dfrbp_1 _13223_ (.CLK(clknet_leaf_54_clk_regs),
    .RESET_B(net3532),
    .D(_00475_),
    .Q_N(_06552_),
    .Q(\u_toplayer.reg_layer2[80] ));
 sg13g2_dfrbp_1 _13224_ (.CLK(clknet_leaf_50_clk_regs),
    .RESET_B(net3513),
    .D(_00476_),
    .Q_N(_06551_),
    .Q(\u_toplayer.reg_layer2[81] ));
 sg13g2_dfrbp_1 _13225_ (.CLK(clknet_leaf_53_clk_regs),
    .RESET_B(net3537),
    .D(_00477_),
    .Q_N(_06550_),
    .Q(\u_toplayer.reg_layer2[82] ));
 sg13g2_dfrbp_1 _13226_ (.CLK(clknet_leaf_52_clk_regs),
    .RESET_B(net3540),
    .D(_00478_),
    .Q_N(_06549_),
    .Q(\u_toplayer.reg_layer2[83] ));
 sg13g2_dfrbp_1 _13227_ (.CLK(clknet_leaf_54_clk_regs),
    .RESET_B(net3533),
    .D(_00479_),
    .Q_N(_06548_),
    .Q(\u_toplayer.reg_layer2[84] ));
 sg13g2_dfrbp_1 _13228_ (.CLK(clknet_leaf_53_clk_regs),
    .RESET_B(net3513),
    .D(_00480_),
    .Q_N(_06547_),
    .Q(\u_toplayer.reg_layer2[85] ));
 sg13g2_dfrbp_1 _13229_ (.CLK(clknet_leaf_87_clk_regs),
    .RESET_B(net3510),
    .D(_00481_),
    .Q_N(_06546_),
    .Q(\u_toplayer.reg_layer2[86] ));
 sg13g2_dfrbp_1 _13230_ (.CLK(clknet_leaf_54_clk_regs),
    .RESET_B(net3533),
    .D(_00482_),
    .Q_N(_06545_),
    .Q(\u_toplayer.reg_layer2[87] ));
 sg13g2_dfrbp_1 _13231_ (.CLK(clknet_leaf_54_clk_regs),
    .RESET_B(net3532),
    .D(_00483_),
    .Q_N(_06544_),
    .Q(\u_toplayer.reg_layer2[88] ));
 sg13g2_dfrbp_1 _13232_ (.CLK(clknet_leaf_51_clk_regs),
    .RESET_B(net3513),
    .D(_00484_),
    .Q_N(_06543_),
    .Q(\u_toplayer.reg_layer2[89] ));
 sg13g2_dfrbp_1 _13233_ (.CLK(clknet_leaf_53_clk_regs),
    .RESET_B(net3537),
    .D(_00485_),
    .Q_N(_06542_),
    .Q(\u_toplayer.reg_layer2[90] ));
 sg13g2_dfrbp_1 _13234_ (.CLK(clknet_leaf_52_clk_regs),
    .RESET_B(net3540),
    .D(_00486_),
    .Q_N(_06541_),
    .Q(\u_toplayer.reg_layer2[91] ));
 sg13g2_dfrbp_1 _13235_ (.CLK(clknet_leaf_54_clk_regs),
    .RESET_B(net3533),
    .D(_00487_),
    .Q_N(_06540_),
    .Q(\u_toplayer.reg_layer2[92] ));
 sg13g2_dfrbp_1 _13236_ (.CLK(clknet_leaf_53_clk_regs),
    .RESET_B(net3513),
    .D(_00488_),
    .Q_N(_06539_),
    .Q(\u_toplayer.reg_layer2[93] ));
 sg13g2_dfrbp_1 _13237_ (.CLK(clknet_leaf_87_clk_regs),
    .RESET_B(net3510),
    .D(_00489_),
    .Q_N(_06538_),
    .Q(\u_toplayer.reg_layer2[94] ));
 sg13g2_dfrbp_1 _13238_ (.CLK(clknet_leaf_86_clk_regs),
    .RESET_B(net3532),
    .D(_00490_),
    .Q_N(_06537_),
    .Q(\u_toplayer.reg_layer2[95] ));
 sg13g2_dfrbp_1 _13239_ (.CLK(clknet_leaf_59_clk_regs),
    .RESET_B(net3546),
    .D(net382),
    .Q_N(_06536_),
    .Q(\u_toplayer.reg_layer2[96] ));
 sg13g2_dfrbp_1 _13240_ (.CLK(clknet_leaf_56_clk_regs),
    .RESET_B(net3541),
    .D(net398),
    .Q_N(_06535_),
    .Q(\u_toplayer.reg_layer2[97] ));
 sg13g2_dfrbp_1 _13241_ (.CLK(clknet_leaf_60_clk_regs),
    .RESET_B(net3545),
    .D(_00493_),
    .Q_N(_06534_),
    .Q(\u_toplayer.reg_layer2[98] ));
 sg13g2_dfrbp_1 _13242_ (.CLK(clknet_leaf_60_clk_regs),
    .RESET_B(net3545),
    .D(_00494_),
    .Q_N(_06533_),
    .Q(\u_toplayer.reg_layer2[99] ));
 sg13g2_dfrbp_1 _13243_ (.CLK(clknet_leaf_62_clk_regs),
    .RESET_B(net3542),
    .D(_00495_),
    .Q_N(_06532_),
    .Q(\u_toplayer.reg_layer2[100] ));
 sg13g2_dfrbp_1 _13244_ (.CLK(clknet_leaf_60_clk_regs),
    .RESET_B(net3545),
    .D(_00496_),
    .Q_N(_06531_),
    .Q(\u_toplayer.reg_layer2[101] ));
 sg13g2_dfrbp_1 _13245_ (.CLK(clknet_leaf_62_clk_regs),
    .RESET_B(net3543),
    .D(_00497_),
    .Q_N(_06530_),
    .Q(\u_toplayer.reg_layer2[102] ));
 sg13g2_dfrbp_1 _13246_ (.CLK(clknet_leaf_62_clk_regs),
    .RESET_B(net3542),
    .D(_00498_),
    .Q_N(_06529_),
    .Q(\u_toplayer.reg_layer2[103] ));
 sg13g2_dfrbp_1 _13247_ (.CLK(clknet_leaf_58_clk_regs),
    .RESET_B(net3546),
    .D(net208),
    .Q_N(_06528_),
    .Q(\u_toplayer.reg_layer2[104] ));
 sg13g2_dfrbp_1 _13248_ (.CLK(clknet_leaf_59_clk_regs),
    .RESET_B(net3546),
    .D(_00500_),
    .Q_N(_06527_),
    .Q(\u_toplayer.reg_layer2[105] ));
 sg13g2_dfrbp_1 _13249_ (.CLK(clknet_leaf_59_clk_regs),
    .RESET_B(net3547),
    .D(_00501_),
    .Q_N(_06526_),
    .Q(\u_toplayer.reg_layer2[106] ));
 sg13g2_dfrbp_1 _13250_ (.CLK(clknet_leaf_60_clk_regs),
    .RESET_B(net3545),
    .D(net227),
    .Q_N(_06525_),
    .Q(\u_toplayer.reg_layer2[107] ));
 sg13g2_dfrbp_1 _13251_ (.CLK(clknet_leaf_62_clk_regs),
    .RESET_B(net3542),
    .D(net229),
    .Q_N(_06524_),
    .Q(\u_toplayer.reg_layer2[108] ));
 sg13g2_dfrbp_1 _13252_ (.CLK(clknet_leaf_60_clk_regs),
    .RESET_B(net3545),
    .D(_00504_),
    .Q_N(_06523_),
    .Q(\u_toplayer.reg_layer2[109] ));
 sg13g2_dfrbp_1 _13253_ (.CLK(clknet_leaf_62_clk_regs),
    .RESET_B(net3543),
    .D(_00505_),
    .Q_N(_06522_),
    .Q(\u_toplayer.reg_layer2[110] ));
 sg13g2_dfrbp_1 _13254_ (.CLK(clknet_leaf_61_clk_regs),
    .RESET_B(net3544),
    .D(_00506_),
    .Q_N(_06521_),
    .Q(\u_toplayer.reg_layer2[111] ));
 sg13g2_dfrbp_1 _13255_ (.CLK(clknet_leaf_64_clk_regs),
    .RESET_B(net3541),
    .D(_00507_),
    .Q_N(_06520_),
    .Q(\u_toplayer.reg_layer2[112] ));
 sg13g2_dfrbp_1 _13256_ (.CLK(clknet_leaf_64_clk_regs),
    .RESET_B(net3528),
    .D(_00508_),
    .Q_N(_06519_),
    .Q(\u_toplayer.reg_layer2[113] ));
 sg13g2_dfrbp_1 _13257_ (.CLK(clknet_leaf_61_clk_regs),
    .RESET_B(net3542),
    .D(_00509_),
    .Q_N(_06518_),
    .Q(\u_toplayer.reg_layer2[114] ));
 sg13g2_dfrbp_1 _13258_ (.CLK(clknet_leaf_61_clk_regs),
    .RESET_B(net3544),
    .D(_00510_),
    .Q_N(_06517_),
    .Q(\u_toplayer.reg_layer2[115] ));
 sg13g2_dfrbp_1 _13259_ (.CLK(clknet_leaf_63_clk_regs),
    .RESET_B(net3529),
    .D(_00511_),
    .Q_N(_06516_),
    .Q(\u_toplayer.reg_layer2[116] ));
 sg13g2_dfrbp_1 _13260_ (.CLK(clknet_leaf_63_clk_regs),
    .RESET_B(net3527),
    .D(_00512_),
    .Q_N(_06515_),
    .Q(\u_toplayer.reg_layer2[117] ));
 sg13g2_dfrbp_1 _13261_ (.CLK(clknet_leaf_64_clk_regs),
    .RESET_B(net3542),
    .D(_00513_),
    .Q_N(_06514_),
    .Q(\u_toplayer.reg_layer2[118] ));
 sg13g2_dfrbp_1 _13262_ (.CLK(clknet_leaf_63_clk_regs),
    .RESET_B(net3529),
    .D(_00514_),
    .Q_N(_06513_),
    .Q(\u_toplayer.reg_layer2[119] ));
 sg13g2_dfrbp_1 _13263_ (.CLK(clknet_leaf_66_clk_regs),
    .RESET_B(net3522),
    .D(_00515_),
    .Q_N(_06512_),
    .Q(\u_toplayer.reg_layer2[120] ));
 sg13g2_dfrbp_1 _13264_ (.CLK(clknet_leaf_65_clk_regs),
    .RESET_B(net3528),
    .D(_00516_),
    .Q_N(_06511_),
    .Q(\u_toplayer.reg_layer2[121] ));
 sg13g2_dfrbp_1 _13265_ (.CLK(clknet_leaf_61_clk_regs),
    .RESET_B(net3543),
    .D(_00517_),
    .Q_N(_06510_),
    .Q(\u_toplayer.reg_layer2[122] ));
 sg13g2_dfrbp_1 _13266_ (.CLK(clknet_leaf_61_clk_regs),
    .RESET_B(net3541),
    .D(_00518_),
    .Q_N(_06509_),
    .Q(\u_toplayer.reg_layer2[123] ));
 sg13g2_dfrbp_1 _13267_ (.CLK(clknet_leaf_68_clk_regs),
    .RESET_B(net3530),
    .D(_00519_),
    .Q_N(_06508_),
    .Q(\u_toplayer.reg_layer2[124] ));
 sg13g2_dfrbp_1 _13268_ (.CLK(clknet_leaf_67_clk_regs),
    .RESET_B(net3528),
    .D(_00520_),
    .Q_N(_06507_),
    .Q(\u_toplayer.reg_layer2[125] ));
 sg13g2_dfrbp_1 _13269_ (.CLK(clknet_leaf_61_clk_regs),
    .RESET_B(net3542),
    .D(_00521_),
    .Q_N(_06506_),
    .Q(\u_toplayer.reg_layer2[126] ));
 sg13g2_dfrbp_1 _13270_ (.CLK(clknet_leaf_68_clk_regs),
    .RESET_B(net3529),
    .D(_00522_),
    .Q_N(_06505_),
    .Q(\u_toplayer.reg_layer2[127] ));
 sg13g2_dfrbp_1 _13271_ (.CLK(clknet_leaf_75_clk_regs),
    .RESET_B(net3502),
    .D(_00523_),
    .Q_N(_06504_),
    .Q(\u_toplayer.reg_layer2[128] ));
 sg13g2_dfrbp_1 _13272_ (.CLK(clknet_leaf_88_clk_regs),
    .RESET_B(net3511),
    .D(_00524_),
    .Q_N(_06503_),
    .Q(\u_toplayer.reg_layer2[129] ));
 sg13g2_dfrbp_1 _13273_ (.CLK(clknet_leaf_85_clk_regs),
    .RESET_B(net3503),
    .D(_00525_),
    .Q_N(_06502_),
    .Q(\u_toplayer.reg_layer2[130] ));
 sg13g2_dfrbp_1 _13274_ (.CLK(clknet_leaf_85_clk_regs),
    .RESET_B(net3502),
    .D(_00526_),
    .Q_N(_06501_),
    .Q(\u_toplayer.reg_layer2[131] ));
 sg13g2_dfrbp_1 _13275_ (.CLK(clknet_leaf_86_clk_regs),
    .RESET_B(net3510),
    .D(_00527_),
    .Q_N(_06500_),
    .Q(\u_toplayer.reg_layer2[132] ));
 sg13g2_dfrbp_1 _13276_ (.CLK(clknet_leaf_84_clk_regs),
    .RESET_B(net3502),
    .D(_00528_),
    .Q_N(_06499_),
    .Q(\u_toplayer.reg_layer2[133] ));
 sg13g2_dfrbp_1 _13277_ (.CLK(clknet_leaf_75_clk_regs),
    .RESET_B(net3502),
    .D(_00529_),
    .Q_N(_06498_),
    .Q(\u_toplayer.reg_layer2[134] ));
 sg13g2_dfrbp_1 _13278_ (.CLK(clknet_leaf_75_clk_regs),
    .RESET_B(net3499),
    .D(_00530_),
    .Q_N(_06497_),
    .Q(\u_toplayer.reg_layer2[135] ));
 sg13g2_dfrbp_1 _13279_ (.CLK(clknet_leaf_76_clk_regs),
    .RESET_B(net3499),
    .D(_00531_),
    .Q_N(_06496_),
    .Q(\u_toplayer.reg_layer2[136] ));
 sg13g2_dfrbp_1 _13280_ (.CLK(clknet_leaf_85_clk_regs),
    .RESET_B(net3502),
    .D(_00532_),
    .Q_N(_06495_),
    .Q(\u_toplayer.reg_layer2[137] ));
 sg13g2_dfrbp_1 _13281_ (.CLK(clknet_leaf_75_clk_regs),
    .RESET_B(net3503),
    .D(_00533_),
    .Q_N(_06494_),
    .Q(\u_toplayer.reg_layer2[138] ));
 sg13g2_dfrbp_1 _13282_ (.CLK(clknet_leaf_85_clk_regs),
    .RESET_B(net3503),
    .D(_00534_),
    .Q_N(_06493_),
    .Q(\u_toplayer.reg_layer2[139] ));
 sg13g2_dfrbp_1 _13283_ (.CLK(clknet_leaf_86_clk_regs),
    .RESET_B(net3510),
    .D(net648),
    .Q_N(_06492_),
    .Q(\u_toplayer.reg_layer2[140] ));
 sg13g2_dfrbp_1 _13284_ (.CLK(clknet_leaf_84_clk_regs),
    .RESET_B(net3503),
    .D(_00536_),
    .Q_N(_06491_),
    .Q(\u_toplayer.reg_layer2[141] ));
 sg13g2_dfrbp_1 _13285_ (.CLK(clknet_leaf_75_clk_regs),
    .RESET_B(net3502),
    .D(_00537_),
    .Q_N(_06490_),
    .Q(\u_toplayer.reg_layer2[142] ));
 sg13g2_dfrbp_1 _13286_ (.CLK(clknet_leaf_76_clk_regs),
    .RESET_B(net3499),
    .D(_00538_),
    .Q_N(_06489_),
    .Q(\u_toplayer.reg_layer2[143] ));
 sg13g2_dfrbp_1 _13287_ (.CLK(clknet_leaf_78_clk_regs),
    .RESET_B(net3497),
    .D(_00539_),
    .Q_N(_06488_),
    .Q(\u_toplayer.reg_layer2[144] ));
 sg13g2_dfrbp_1 _13288_ (.CLK(clknet_leaf_88_clk_regs),
    .RESET_B(net3511),
    .D(_00540_),
    .Q_N(_06487_),
    .Q(\u_toplayer.reg_layer2[145] ));
 sg13g2_dfrbp_1 _13289_ (.CLK(clknet_leaf_84_clk_regs),
    .RESET_B(net3501),
    .D(_00541_),
    .Q_N(_06486_),
    .Q(\u_toplayer.reg_layer2[146] ));
 sg13g2_dfrbp_1 _13290_ (.CLK(clknet_leaf_83_clk_regs),
    .RESET_B(net3495),
    .D(_00542_),
    .Q_N(_06485_),
    .Q(\u_toplayer.reg_layer2[147] ));
 sg13g2_dfrbp_1 _13291_ (.CLK(clknet_leaf_88_clk_regs),
    .RESET_B(net3511),
    .D(_00543_),
    .Q_N(_06484_),
    .Q(\u_toplayer.reg_layer2[148] ));
 sg13g2_dfrbp_1 _13292_ (.CLK(clknet_leaf_81_clk_regs),
    .RESET_B(net3495),
    .D(_00544_),
    .Q_N(_06483_),
    .Q(\u_toplayer.reg_layer2[149] ));
 sg13g2_dfrbp_1 _13293_ (.CLK(clknet_leaf_81_clk_regs),
    .RESET_B(net3491),
    .D(_00545_),
    .Q_N(_06482_),
    .Q(\u_toplayer.reg_layer2[150] ));
 sg13g2_dfrbp_1 _13294_ (.CLK(clknet_leaf_81_clk_regs),
    .RESET_B(net3491),
    .D(_00546_),
    .Q_N(_06481_),
    .Q(\u_toplayer.reg_layer2[151] ));
 sg13g2_dfrbp_1 _13295_ (.CLK(clknet_leaf_78_clk_regs),
    .RESET_B(net3497),
    .D(_00547_),
    .Q_N(_06480_),
    .Q(\u_toplayer.reg_layer2[152] ));
 sg13g2_dfrbp_1 _13296_ (.CLK(clknet_leaf_84_clk_regs),
    .RESET_B(net3501),
    .D(_00548_),
    .Q_N(_06479_),
    .Q(\u_toplayer.reg_layer2[153] ));
 sg13g2_dfrbp_1 _13297_ (.CLK(clknet_leaf_83_clk_regs),
    .RESET_B(net3504),
    .D(_00549_),
    .Q_N(_06478_),
    .Q(\u_toplayer.reg_layer2[154] ));
 sg13g2_dfrbp_1 _13298_ (.CLK(clknet_leaf_83_clk_regs),
    .RESET_B(net3495),
    .D(_00550_),
    .Q_N(_06477_),
    .Q(\u_toplayer.reg_layer2[155] ));
 sg13g2_dfrbp_1 _13299_ (.CLK(clknet_leaf_84_clk_regs),
    .RESET_B(net3504),
    .D(_00551_),
    .Q_N(_06476_),
    .Q(\u_toplayer.reg_layer2[156] ));
 sg13g2_dfrbp_1 _13300_ (.CLK(clknet_leaf_81_clk_regs),
    .RESET_B(net3495),
    .D(_00552_),
    .Q_N(_06475_),
    .Q(\u_toplayer.reg_layer2[157] ));
 sg13g2_dfrbp_1 _13301_ (.CLK(clknet_leaf_80_clk_regs),
    .RESET_B(net3491),
    .D(_00553_),
    .Q_N(_06474_),
    .Q(\u_toplayer.reg_layer2[158] ));
 sg13g2_dfrbp_1 _13302_ (.CLK(clknet_leaf_81_clk_regs),
    .RESET_B(net3490),
    .D(_00554_),
    .Q_N(_06473_),
    .Q(\u_toplayer.reg_layer2[159] ));
 sg13g2_dfrbp_1 _13303_ (.CLK(clknet_leaf_70_clk_regs),
    .RESET_B(net3524),
    .D(_00555_),
    .Q_N(_06472_),
    .Q(\u_toplayer.reg_layer2[160] ));
 sg13g2_dfrbp_1 _13304_ (.CLK(clknet_leaf_67_clk_regs),
    .RESET_B(net3527),
    .D(_00556_),
    .Q_N(_06471_),
    .Q(\u_toplayer.reg_layer2[161] ));
 sg13g2_dfrbp_1 _13305_ (.CLK(clknet_leaf_69_clk_regs),
    .RESET_B(net3526),
    .D(net436),
    .Q_N(_06470_),
    .Q(\u_toplayer.reg_layer2[162] ));
 sg13g2_dfrbp_1 _13306_ (.CLK(clknet_leaf_68_clk_regs),
    .RESET_B(net3530),
    .D(net601),
    .Q_N(_06469_),
    .Q(\u_toplayer.reg_layer2[163] ));
 sg13g2_dfrbp_1 _13307_ (.CLK(clknet_leaf_67_clk_regs),
    .RESET_B(net3526),
    .D(_00559_),
    .Q_N(_06468_),
    .Q(\u_toplayer.reg_layer2[164] ));
 sg13g2_dfrbp_1 _13308_ (.CLK(clknet_leaf_67_clk_regs),
    .RESET_B(net3525),
    .D(net315),
    .Q_N(_06467_),
    .Q(\u_toplayer.reg_layer2[165] ));
 sg13g2_dfrbp_1 _13309_ (.CLK(clknet_leaf_71_clk_regs),
    .RESET_B(net3518),
    .D(net337),
    .Q_N(_06466_),
    .Q(\u_toplayer.reg_layer2[166] ));
 sg13g2_dfrbp_1 _13310_ (.CLK(clknet_leaf_73_clk_regs),
    .RESET_B(net3525),
    .D(net529),
    .Q_N(_06465_),
    .Q(\u_toplayer.reg_layer2[167] ));
 sg13g2_dfrbp_1 _13311_ (.CLK(clknet_leaf_70_clk_regs),
    .RESET_B(net3524),
    .D(_00563_),
    .Q_N(_06464_),
    .Q(\u_toplayer.reg_layer2[168] ));
 sg13g2_dfrbp_1 _13312_ (.CLK(clknet_leaf_67_clk_regs),
    .RESET_B(net3527),
    .D(_00564_),
    .Q_N(_06463_),
    .Q(\u_toplayer.reg_layer2[169] ));
 sg13g2_dfrbp_1 _13313_ (.CLK(clknet_leaf_69_clk_regs),
    .RESET_B(net3526),
    .D(net829),
    .Q_N(_06462_),
    .Q(\u_toplayer.reg_layer2[170] ));
 sg13g2_dfrbp_1 _13314_ (.CLK(clknet_leaf_68_clk_regs),
    .RESET_B(net3530),
    .D(net777),
    .Q_N(_06461_),
    .Q(\u_toplayer.reg_layer2[171] ));
 sg13g2_dfrbp_1 _13315_ (.CLK(clknet_leaf_69_clk_regs),
    .RESET_B(net3526),
    .D(_00567_),
    .Q_N(_06460_),
    .Q(\u_toplayer.reg_layer2[172] ));
 sg13g2_dfrbp_1 _13316_ (.CLK(clknet_leaf_69_clk_regs),
    .RESET_B(net3524),
    .D(net508),
    .Q_N(_06459_),
    .Q(\u_toplayer.reg_layer2[173] ));
 sg13g2_dfrbp_1 _13317_ (.CLK(clknet_leaf_70_clk_regs),
    .RESET_B(net3524),
    .D(net485),
    .Q_N(_06458_),
    .Q(\u_toplayer.reg_layer2[174] ));
 sg13g2_dfrbp_1 _13318_ (.CLK(clknet_leaf_69_clk_regs),
    .RESET_B(net3525),
    .D(net622),
    .Q_N(_06457_),
    .Q(\u_toplayer.reg_layer2[175] ));
 sg13g2_dfrbp_1 _13319_ (.CLK(clknet_leaf_71_clk_regs),
    .RESET_B(net3518),
    .D(net631),
    .Q_N(_06456_),
    .Q(\u_toplayer.reg_layer2[176] ));
 sg13g2_dfrbp_1 _13320_ (.CLK(clknet_leaf_67_clk_regs),
    .RESET_B(net3519),
    .D(net797),
    .Q_N(_06455_),
    .Q(\u_toplayer.reg_layer2[177] ));
 sg13g2_dfrbp_1 _13321_ (.CLK(clknet_leaf_73_clk_regs),
    .RESET_B(net3516),
    .D(net248),
    .Q_N(_06454_),
    .Q(\u_toplayer.reg_layer2[178] ));
 sg13g2_dfrbp_1 _13322_ (.CLK(clknet_leaf_66_clk_regs),
    .RESET_B(net3522),
    .D(_00574_),
    .Q_N(_06453_),
    .Q(\u_toplayer.reg_layer2[179] ));
 sg13g2_dfrbp_1 _13323_ (.CLK(clknet_leaf_73_clk_regs),
    .RESET_B(net3519),
    .D(net586),
    .Q_N(_06452_),
    .Q(\u_toplayer.reg_layer2[180] ));
 sg13g2_dfrbp_1 _13324_ (.CLK(clknet_leaf_72_clk_regs),
    .RESET_B(net3517),
    .D(net765),
    .Q_N(_06451_),
    .Q(\u_toplayer.reg_layer2[181] ));
 sg13g2_dfrbp_1 _13325_ (.CLK(clknet_leaf_76_clk_regs),
    .RESET_B(net3498),
    .D(_00577_),
    .Q_N(_06450_),
    .Q(\u_toplayer.reg_layer2[182] ));
 sg13g2_dfrbp_1 _13326_ (.CLK(clknet_leaf_73_clk_regs),
    .RESET_B(net3516),
    .D(_00578_),
    .Q_N(_06449_),
    .Q(\u_toplayer.reg_layer2[183] ));
 sg13g2_dfrbp_1 _13327_ (.CLK(clknet_leaf_71_clk_regs),
    .RESET_B(net3518),
    .D(_00579_),
    .Q_N(_06448_),
    .Q(\u_toplayer.reg_layer2[184] ));
 sg13g2_dfrbp_1 _13328_ (.CLK(clknet_leaf_74_clk_regs),
    .RESET_B(net3517),
    .D(_00580_),
    .Q_N(_06447_),
    .Q(\u_toplayer.reg_layer2[185] ));
 sg13g2_dfrbp_1 _13329_ (.CLK(clknet_leaf_72_clk_regs),
    .RESET_B(net3516),
    .D(_00581_),
    .Q_N(_06446_),
    .Q(\u_toplayer.reg_layer2[186] ));
 sg13g2_dfrbp_1 _13330_ (.CLK(clknet_leaf_66_clk_regs),
    .RESET_B(net3522),
    .D(_00582_),
    .Q_N(_06445_),
    .Q(\u_toplayer.reg_layer2[187] ));
 sg13g2_dfrbp_1 _13331_ (.CLK(clknet_leaf_74_clk_regs),
    .RESET_B(net3519),
    .D(_00583_),
    .Q_N(_06444_),
    .Q(\u_toplayer.reg_layer2[188] ));
 sg13g2_dfrbp_1 _13332_ (.CLK(clknet_leaf_72_clk_regs),
    .RESET_B(net3498),
    .D(_00584_),
    .Q_N(_06443_),
    .Q(\u_toplayer.reg_layer2[189] ));
 sg13g2_dfrbp_1 _13333_ (.CLK(clknet_leaf_76_clk_regs),
    .RESET_B(net3498),
    .D(_00585_),
    .Q_N(_06442_),
    .Q(\u_toplayer.reg_layer2[190] ));
 sg13g2_dfrbp_1 _13334_ (.CLK(clknet_leaf_72_clk_regs),
    .RESET_B(net3516),
    .D(_00586_),
    .Q_N(_06441_),
    .Q(\u_toplayer.reg_layer2[191] ));
 sg13g2_dfrbp_1 _13335_ (.CLK(clknet_leaf_55_clk_regs),
    .RESET_B(net3534),
    .D(_00587_),
    .Q_N(_06440_),
    .Q(\u_toplayer.reg_layer2[192] ));
 sg13g2_dfrbp_1 _13336_ (.CLK(clknet_leaf_57_clk_regs),
    .RESET_B(net3537),
    .D(_00588_),
    .Q_N(_06439_),
    .Q(\u_toplayer.reg_layer2[193] ));
 sg13g2_dfrbp_1 _13337_ (.CLK(clknet_leaf_57_clk_regs),
    .RESET_B(net3538),
    .D(_00589_),
    .Q_N(_06438_),
    .Q(\u_toplayer.reg_layer2[194] ));
 sg13g2_dfrbp_1 _13338_ (.CLK(clknet_leaf_57_clk_regs),
    .RESET_B(net3539),
    .D(_00590_),
    .Q_N(_06437_),
    .Q(\u_toplayer.reg_layer2[195] ));
 sg13g2_dfrbp_1 _13339_ (.CLK(clknet_leaf_65_clk_regs),
    .RESET_B(net3534),
    .D(_00591_),
    .Q_N(_06436_),
    .Q(\u_toplayer.reg_layer2[196] ));
 sg13g2_dfrbp_1 _13340_ (.CLK(clknet_leaf_55_clk_regs),
    .RESET_B(net3535),
    .D(_00592_),
    .Q_N(_06435_),
    .Q(\u_toplayer.reg_layer2[197] ));
 sg13g2_dfrbp_1 _13341_ (.CLK(clknet_leaf_55_clk_regs),
    .RESET_B(net3535),
    .D(_00593_),
    .Q_N(_06434_),
    .Q(\u_toplayer.reg_layer2[198] ));
 sg13g2_dfrbp_1 _13342_ (.CLK(clknet_leaf_65_clk_regs),
    .RESET_B(net3521),
    .D(_00594_),
    .Q_N(_06433_),
    .Q(\u_toplayer.reg_layer2[199] ));
 sg13g2_dfrbp_1 _13343_ (.CLK(clknet_leaf_56_clk_regs),
    .RESET_B(net3538),
    .D(net237),
    .Q_N(_06432_),
    .Q(\u_toplayer.reg_layer2[200] ));
 sg13g2_dfrbp_1 _13344_ (.CLK(clknet_leaf_57_clk_regs),
    .RESET_B(net3539),
    .D(net445),
    .Q_N(_06431_),
    .Q(\u_toplayer.reg_layer2[201] ));
 sg13g2_dfrbp_1 _13345_ (.CLK(clknet_leaf_58_clk_regs),
    .RESET_B(net3538),
    .D(net205),
    .Q_N(_06430_),
    .Q(\u_toplayer.reg_layer2[202] ));
 sg13g2_dfrbp_1 _13346_ (.CLK(clknet_leaf_58_clk_regs),
    .RESET_B(net3539),
    .D(_00598_),
    .Q_N(_06429_),
    .Q(\u_toplayer.reg_layer2[203] ));
 sg13g2_dfrbp_1 _13347_ (.CLK(clknet_leaf_65_clk_regs),
    .RESET_B(net3534),
    .D(_00599_),
    .Q_N(_06428_),
    .Q(\u_toplayer.reg_layer2[204] ));
 sg13g2_dfrbp_1 _13348_ (.CLK(clknet_leaf_56_clk_regs),
    .RESET_B(net3538),
    .D(net394),
    .Q_N(_06427_),
    .Q(\u_toplayer.reg_layer2[205] ));
 sg13g2_dfrbp_1 _13349_ (.CLK(clknet_leaf_55_clk_regs),
    .RESET_B(net3535),
    .D(net319),
    .Q_N(_06426_),
    .Q(\u_toplayer.reg_layer2[206] ));
 sg13g2_dfrbp_1 _13350_ (.CLK(clknet_leaf_65_clk_regs),
    .RESET_B(net3534),
    .D(net708),
    .Q_N(_06425_),
    .Q(\u_toplayer.reg_layer2[207] ));
 sg13g2_dfrbp_1 _13351_ (.CLK(clknet_leaf_54_clk_regs),
    .RESET_B(net3533),
    .D(_00603_),
    .Q_N(_06424_),
    .Q(\u_toplayer.reg_layer2[208] ));
 sg13g2_dfrbp_1 _13352_ (.CLK(clknet_leaf_50_clk_regs),
    .RESET_B(net3513),
    .D(_00604_),
    .Q_N(_06423_),
    .Q(\u_toplayer.reg_layer2[209] ));
 sg13g2_dfrbp_1 _13353_ (.CLK(clknet_leaf_52_clk_regs),
    .RESET_B(net3537),
    .D(_00605_),
    .Q_N(_06422_),
    .Q(\u_toplayer.reg_layer2[210] ));
 sg13g2_dfrbp_1 _13354_ (.CLK(clknet_leaf_51_clk_regs),
    .RESET_B(net3513),
    .D(_00606_),
    .Q_N(_06421_),
    .Q(\u_toplayer.reg_layer2[211] ));
 sg13g2_dfrbp_1 _13355_ (.CLK(clknet_leaf_54_clk_regs),
    .RESET_B(net3532),
    .D(_00607_),
    .Q_N(_06420_),
    .Q(\u_toplayer.reg_layer2[212] ));
 sg13g2_dfrbp_1 _13356_ (.CLK(clknet_leaf_53_clk_regs),
    .RESET_B(net3513),
    .D(_00608_),
    .Q_N(_06419_),
    .Q(\u_toplayer.reg_layer2[213] ));
 sg13g2_dfrbp_1 _13357_ (.CLK(clknet_leaf_87_clk_regs),
    .RESET_B(net3510),
    .D(_00609_),
    .Q_N(_06418_),
    .Q(\u_toplayer.reg_layer2[214] ));
 sg13g2_dfrbp_1 _13358_ (.CLK(clknet_leaf_86_clk_regs),
    .RESET_B(net3532),
    .D(_00610_),
    .Q_N(_06417_),
    .Q(\u_toplayer.reg_layer2[215] ));
 sg13g2_dfrbp_1 _13359_ (.CLK(clknet_leaf_53_clk_regs),
    .RESET_B(net3537),
    .D(_00611_),
    .Q_N(_06416_),
    .Q(\u_toplayer.reg_layer2[216] ));
 sg13g2_dfrbp_1 _13360_ (.CLK(clknet_leaf_51_clk_regs),
    .RESET_B(net3513),
    .D(_00612_),
    .Q_N(_06415_),
    .Q(\u_toplayer.reg_layer2[217] ));
 sg13g2_dfrbp_1 _13361_ (.CLK(clknet_leaf_53_clk_regs),
    .RESET_B(net3537),
    .D(_00613_),
    .Q_N(_06414_),
    .Q(\u_toplayer.reg_layer2[218] ));
 sg13g2_dfrbp_1 _13362_ (.CLK(clknet_leaf_51_clk_regs),
    .RESET_B(net3514),
    .D(_00614_),
    .Q_N(_06413_),
    .Q(\u_toplayer.reg_layer2[219] ));
 sg13g2_dfrbp_1 _13363_ (.CLK(clknet_leaf_86_clk_regs),
    .RESET_B(net3532),
    .D(_00615_),
    .Q_N(_06412_),
    .Q(\u_toplayer.reg_layer2[220] ));
 sg13g2_dfrbp_1 _13364_ (.CLK(clknet_leaf_53_clk_regs),
    .RESET_B(net3510),
    .D(_00616_),
    .Q_N(_06411_),
    .Q(\u_toplayer.reg_layer2[221] ));
 sg13g2_dfrbp_1 _13365_ (.CLK(clknet_leaf_87_clk_regs),
    .RESET_B(net3510),
    .D(_00617_),
    .Q_N(_06410_),
    .Q(\u_toplayer.reg_layer2[222] ));
 sg13g2_dfrbp_1 _13366_ (.CLK(clknet_leaf_86_clk_regs),
    .RESET_B(net3532),
    .D(_00618_),
    .Q_N(_06409_),
    .Q(\u_toplayer.reg_layer2[223] ));
 sg13g2_dfrbp_1 _13367_ (.CLK(clknet_leaf_58_clk_regs),
    .RESET_B(net3546),
    .D(net510),
    .Q_N(_06408_),
    .Q(\u_toplayer.reg_layer2[224] ));
 sg13g2_dfrbp_1 _13368_ (.CLK(clknet_leaf_56_clk_regs),
    .RESET_B(net3541),
    .D(net551),
    .Q_N(_06407_),
    .Q(\u_toplayer.reg_layer2[225] ));
 sg13g2_dfrbp_1 _13369_ (.CLK(clknet_leaf_59_clk_regs),
    .RESET_B(net3545),
    .D(_00621_),
    .Q_N(_06406_),
    .Q(\u_toplayer.reg_layer2[226] ));
 sg13g2_dfrbp_1 _13370_ (.CLK(clknet_leaf_59_clk_regs),
    .RESET_B(net3546),
    .D(_00622_),
    .Q_N(_06405_),
    .Q(\u_toplayer.reg_layer2[227] ));
 sg13g2_dfrbp_1 _13371_ (.CLK(clknet_leaf_63_clk_regs),
    .RESET_B(net3529),
    .D(_00623_),
    .Q_N(_06404_),
    .Q(\u_toplayer.reg_layer2[228] ));
 sg13g2_dfrbp_1 _13372_ (.CLK(clknet_leaf_60_clk_regs),
    .RESET_B(net3545),
    .D(_00624_),
    .Q_N(_06403_),
    .Q(\u_toplayer.reg_layer2[229] ));
 sg13g2_dfrbp_1 _13373_ (.CLK(clknet_leaf_61_clk_regs),
    .RESET_B(net3543),
    .D(_00625_),
    .Q_N(_06402_),
    .Q(\u_toplayer.reg_layer2[230] ));
 sg13g2_dfrbp_1 _13374_ (.CLK(clknet_leaf_62_clk_regs),
    .RESET_B(net3543),
    .D(_00626_),
    .Q_N(_06401_),
    .Q(\u_toplayer.reg_layer2[231] ));
 sg13g2_dfrbp_1 _13375_ (.CLK(clknet_leaf_58_clk_regs),
    .RESET_B(net3546),
    .D(net658),
    .Q_N(_06400_),
    .Q(\u_toplayer.reg_layer2[232] ));
 sg13g2_dfrbp_1 _13376_ (.CLK(clknet_leaf_58_clk_regs),
    .RESET_B(net3546),
    .D(_00628_),
    .Q_N(_06399_),
    .Q(\u_toplayer.reg_layer2[233] ));
 sg13g2_dfrbp_1 _13377_ (.CLK(clknet_leaf_59_clk_regs),
    .RESET_B(net3547),
    .D(_00629_),
    .Q_N(_06398_),
    .Q(\u_toplayer.reg_layer2[234] ));
 sg13g2_dfrbp_1 _13378_ (.CLK(clknet_leaf_59_clk_regs),
    .RESET_B(net3546),
    .D(net441),
    .Q_N(_06397_),
    .Q(\u_toplayer.reg_layer2[235] ));
 sg13g2_dfrbp_1 _13379_ (.CLK(clknet_leaf_63_clk_regs),
    .RESET_B(net3529),
    .D(net303),
    .Q_N(_06396_),
    .Q(\u_toplayer.reg_layer2[236] ));
 sg13g2_dfrbp_1 _13380_ (.CLK(clknet_leaf_60_clk_regs),
    .RESET_B(net3545),
    .D(_00632_),
    .Q_N(_06395_),
    .Q(\u_toplayer.reg_layer2[237] ));
 sg13g2_dfrbp_1 _13381_ (.CLK(clknet_leaf_60_clk_regs),
    .RESET_B(net3543),
    .D(_00633_),
    .Q_N(_06394_),
    .Q(\u_toplayer.reg_layer2[238] ));
 sg13g2_dfrbp_1 _13382_ (.CLK(clknet_leaf_62_clk_regs),
    .RESET_B(net3543),
    .D(_00634_),
    .Q_N(_06393_),
    .Q(\u_toplayer.reg_layer2[239] ));
 sg13g2_dfrbp_1 _13383_ (.CLK(clknet_leaf_56_clk_regs),
    .RESET_B(net3541),
    .D(_00635_),
    .Q_N(_06392_),
    .Q(\u_toplayer.reg_layer2[240] ));
 sg13g2_dfrbp_1 _13384_ (.CLK(clknet_leaf_64_clk_regs),
    .RESET_B(net3528),
    .D(_00636_),
    .Q_N(_06391_),
    .Q(\u_toplayer.reg_layer2[241] ));
 sg13g2_dfrbp_1 _13385_ (.CLK(clknet_leaf_64_clk_regs),
    .RESET_B(net3541),
    .D(_00637_),
    .Q_N(_06390_),
    .Q(\u_toplayer.reg_layer2[242] ));
 sg13g2_dfrbp_1 _13386_ (.CLK(clknet_leaf_64_clk_regs),
    .RESET_B(net3541),
    .D(_00638_),
    .Q_N(_06389_),
    .Q(\u_toplayer.reg_layer2[243] ));
 sg13g2_dfrbp_1 _13387_ (.CLK(clknet_leaf_63_clk_regs),
    .RESET_B(net3529),
    .D(_00639_),
    .Q_N(_06388_),
    .Q(\u_toplayer.reg_layer2[244] ));
 sg13g2_dfrbp_1 _13388_ (.CLK(clknet_leaf_63_clk_regs),
    .RESET_B(net3527),
    .D(_00640_),
    .Q_N(_06387_),
    .Q(\u_toplayer.reg_layer2[245] ));
 sg13g2_dfrbp_1 _13389_ (.CLK(clknet_leaf_64_clk_regs),
    .RESET_B(net3542),
    .D(_00641_),
    .Q_N(_06386_),
    .Q(\u_toplayer.reg_layer2[246] ));
 sg13g2_dfrbp_1 _13390_ (.CLK(clknet_leaf_63_clk_regs),
    .RESET_B(net3529),
    .D(_00642_),
    .Q_N(_06385_),
    .Q(\u_toplayer.reg_layer2[247] ));
 sg13g2_dfrbp_1 _13391_ (.CLK(clknet_leaf_66_clk_regs),
    .RESET_B(net3522),
    .D(_00643_),
    .Q_N(_06384_),
    .Q(\u_toplayer.reg_layer2[248] ));
 sg13g2_dfrbp_1 _13392_ (.CLK(clknet_leaf_65_clk_regs),
    .RESET_B(net3528),
    .D(_00644_),
    .Q_N(_06383_),
    .Q(\u_toplayer.reg_layer2[249] ));
 sg13g2_dfrbp_1 _13393_ (.CLK(clknet_leaf_61_clk_regs),
    .RESET_B(net3544),
    .D(_00645_),
    .Q_N(_06382_),
    .Q(\u_toplayer.reg_layer2[250] ));
 sg13g2_dfrbp_1 _13394_ (.CLK(clknet_leaf_56_clk_regs),
    .RESET_B(net3541),
    .D(_00646_),
    .Q_N(_06381_),
    .Q(\u_toplayer.reg_layer2[251] ));
 sg13g2_dfrbp_1 _13395_ (.CLK(clknet_leaf_68_clk_regs),
    .RESET_B(net3529),
    .D(_00647_),
    .Q_N(_06380_),
    .Q(\u_toplayer.reg_layer2[252] ));
 sg13g2_dfrbp_1 _13396_ (.CLK(clknet_leaf_66_clk_regs),
    .RESET_B(net3527),
    .D(_00648_),
    .Q_N(_06379_),
    .Q(\u_toplayer.reg_layer2[253] ));
 sg13g2_dfrbp_1 _13397_ (.CLK(clknet_leaf_62_clk_regs),
    .RESET_B(net3542),
    .D(_00649_),
    .Q_N(_06378_),
    .Q(\u_toplayer.reg_layer2[254] ));
 sg13g2_dfrbp_1 _13398_ (.CLK(clknet_leaf_68_clk_regs),
    .RESET_B(net3530),
    .D(_00650_),
    .Q_N(_06377_),
    .Q(\u_toplayer.reg_layer2[255] ));
 sg13g2_dfrbp_1 _13399_ (.CLK(clknet_leaf_79_clk_regs),
    .RESET_B(net3491),
    .D(net981),
    .Q_N(_06881_),
    .Q(\u_toplayer.done_layer2 ));
 sg13g2_dfrbp_1 _13400_ (.CLK(clknet_leaf_52_clk_regs),
    .RESET_B(net3551),
    .D(_00019_),
    .Q_N(_06882_),
    .Q(\u_toplayer.u_layer3.u_neuron.instCtrl.state[0] ));
 sg13g2_dfrbp_1 _13401_ (.CLK(clknet_leaf_52_clk_regs),
    .RESET_B(net3551),
    .D(net882),
    .Q_N(_06883_),
    .Q(\u_toplayer.u_layer3.u_neuron.instCtrl.state[1] ));
 sg13g2_dfrbp_1 _13402_ (.CLK(clknet_leaf_52_clk_regs),
    .RESET_B(net3514),
    .D(_00021_),
    .Q_N(_00037_),
    .Q(\u_toplayer.u_layer3.u_neuron.instCtrl.state[2] ));
 sg13g2_dfrbp_1 _13403_ (.CLK(clknet_leaf_52_clk_regs),
    .RESET_B(net3514),
    .D(net1006),
    .Q_N(_00038_),
    .Q(\u_toplayer.u_layer3.u_neuron.instCtrl.state[3] ));
 sg13g2_dfrbp_1 _13404_ (.CLK(clknet_leaf_51_clk_regs),
    .RESET_B(net3551),
    .D(net967),
    .Q_N(_00039_),
    .Q(\u_toplayer.u_layer3.u_neuron.instCtrl.state[4] ));
 sg13g2_dfrbp_1 _13405_ (.CLK(clknet_leaf_48_clk_regs),
    .RESET_B(net3551),
    .D(net683),
    .Q_N(_00034_),
    .Q(\u_toplayer.u_layer3.u_neuron.instCtrl.state[5] ));
 sg13g2_dfrbp_1 _13406_ (.CLK(clknet_leaf_92_clk_regs),
    .RESET_B(net3451),
    .D(_00652_),
    .Q_N(_06376_),
    .Q(\u_toplayer.u_layer2.u_neuron.din[0] ));
 sg13g2_dfrbp_1 _13407_ (.CLK(clknet_leaf_16_clk_regs),
    .RESET_B(net3453),
    .D(_00653_),
    .Q_N(_06375_),
    .Q(\u_toplayer.u_layer2.u_neuron.din[1] ));
 sg13g2_dfrbp_1 _13408_ (.CLK(clknet_leaf_15_clk_regs),
    .RESET_B(net3453),
    .D(net1142),
    .Q_N(_06374_),
    .Q(\u_toplayer.u_layer2.u_neuron.din[2] ));
 sg13g2_dfrbp_1 _13409_ (.CLK(clknet_leaf_15_clk_regs),
    .RESET_B(net3448),
    .D(_00655_),
    .Q_N(_06373_),
    .Q(\u_toplayer.u_layer2.u_neuron.din[3] ));
 sg13g2_dfrbp_1 _13410_ (.CLK(clknet_leaf_14_clk_regs),
    .RESET_B(net3449),
    .D(_00656_),
    .Q_N(_06372_),
    .Q(\u_toplayer.u_layer2.u_neuron.din[4] ));
 sg13g2_dfrbp_1 _13411_ (.CLK(clknet_leaf_15_clk_regs),
    .RESET_B(net3448),
    .D(_00657_),
    .Q_N(_06371_),
    .Q(\u_toplayer.u_layer2.u_neuron.din[5] ));
 sg13g2_dfrbp_1 _13412_ (.CLK(clknet_leaf_15_clk_regs),
    .RESET_B(net3449),
    .D(_00658_),
    .Q_N(_06370_),
    .Q(\u_toplayer.u_layer2.u_neuron.din[6] ));
 sg13g2_dfrbp_1 _13413_ (.CLK(clknet_leaf_15_clk_regs),
    .RESET_B(net3448),
    .D(_00659_),
    .Q_N(_06369_),
    .Q(\u_toplayer.u_layer2.u_neuron.din[7] ));
 sg13g2_dfrbp_1 _13414_ (.CLK(clknet_leaf_51_clk_regs),
    .RESET_B(net3512),
    .D(_00660_),
    .Q_N(_06368_),
    .Q(\u_toplayer.u_layer2.sum[0] ));
 sg13g2_dfrbp_1 _13415_ (.CLK(clknet_leaf_51_clk_regs),
    .RESET_B(net3512),
    .D(_00661_),
    .Q_N(_06367_),
    .Q(\u_toplayer.u_layer2.sum[1] ));
 sg13g2_dfrbp_1 _13416_ (.CLK(clknet_leaf_51_clk_regs),
    .RESET_B(net3512),
    .D(_00662_),
    .Q_N(_06366_),
    .Q(\u_toplayer.u_layer2.sum[2] ));
 sg13g2_dfrbp_1 _13417_ (.CLK(clknet_leaf_50_clk_regs),
    .RESET_B(net3512),
    .D(_00663_),
    .Q_N(_06365_),
    .Q(\u_toplayer.u_layer2.sum[3] ));
 sg13g2_dfrbp_1 _13418_ (.CLK(clknet_leaf_50_clk_regs),
    .RESET_B(net3512),
    .D(_00664_),
    .Q_N(_06364_),
    .Q(\u_toplayer.u_layer2.sum[4] ));
 sg13g2_dfrbp_1 _13419_ (.CLK(clknet_leaf_50_clk_regs),
    .RESET_B(net3512),
    .D(_00665_),
    .Q_N(_06363_),
    .Q(\u_toplayer.u_layer2.sum[5] ));
 sg13g2_dfrbp_1 _13420_ (.CLK(clknet_leaf_50_clk_regs),
    .RESET_B(net3512),
    .D(_00666_),
    .Q_N(_06362_),
    .Q(\u_toplayer.u_layer2.sum[6] ));
 sg13g2_dfrbp_1 _13421_ (.CLK(clknet_leaf_87_clk_regs),
    .RESET_B(net3511),
    .D(_00667_),
    .Q_N(_06361_),
    .Q(\u_toplayer.u_layer2.sum[7] ));
 sg13g2_dfrbp_1 _13422_ (.CLK(clknet_leaf_79_clk_regs),
    .RESET_B(net3490),
    .D(_00668_),
    .Q_N(_06360_),
    .Q(\u_toplayer.u_layer2.statel2[0] ));
 sg13g2_dfrbp_1 _13423_ (.CLK(clknet_leaf_79_clk_regs),
    .RESET_B(net3490),
    .D(_00669_),
    .Q_N(_06359_),
    .Q(\u_toplayer.u_layer2.statel2[1] ));
 sg13g2_dfrbp_1 _13424_ (.CLK(clknet_leaf_79_clk_regs),
    .RESET_B(net3490),
    .D(_00670_),
    .Q_N(_06358_),
    .Q(\u_toplayer.u_layer2.statel2[2] ));
 sg13g2_dfrbp_1 _13425_ (.CLK(clknet_leaf_79_clk_regs),
    .RESET_B(net3488),
    .D(_00671_),
    .Q_N(_06357_),
    .Q(\u_toplayer.u_layer2.statel2[3] ));
 sg13g2_dfrbp_1 _13426_ (.CLK(clknet_leaf_79_clk_regs),
    .RESET_B(net3488),
    .D(_00672_),
    .Q_N(_06356_),
    .Q(\u_toplayer.u_layer2.statel2[4] ));
 sg13g2_dfrbp_1 _13427_ (.CLK(clknet_leaf_79_clk_regs),
    .RESET_B(net3490),
    .D(net938),
    .Q_N(_06355_),
    .Q(\u_toplayer.u_layer2.statel2[5] ));
 sg13g2_dfrbp_1 _13428_ (.CLK(clknet_leaf_78_clk_regs),
    .RESET_B(net3490),
    .D(_00674_),
    .Q_N(_06354_),
    .Q(\u_toplayer.u_layer2.statel2[6] ));
 sg13g2_dfrbp_1 _13429_ (.CLK(clknet_leaf_78_clk_regs),
    .RESET_B(net3490),
    .D(_00675_),
    .Q_N(_06353_),
    .Q(\u_toplayer.u_layer2.statel2[7] ));
 sg13g2_dfrbp_1 _13430_ (.CLK(clknet_leaf_78_clk_regs),
    .RESET_B(net3490),
    .D(net123),
    .Q_N(_00031_),
    .Q(\u_toplayer.u_layer2.statel2[8] ));
 sg13g2_dfrbp_1 _13431_ (.CLK(clknet_leaf_49_clk_regs),
    .RESET_B(net3551),
    .D(net1038),
    .Q_N(_06352_),
    .Q(\u_toplayer.u_layer2.u_neuron.acc[0] ));
 sg13g2_dfrbp_1 _13432_ (.CLK(clknet_leaf_48_clk_regs),
    .RESET_B(net3551),
    .D(_00678_),
    .Q_N(_06351_),
    .Q(\u_toplayer.u_layer2.u_neuron.acc[1] ));
 sg13g2_dfrbp_1 _13433_ (.CLK(clknet_leaf_49_clk_regs),
    .RESET_B(net3551),
    .D(_00679_),
    .Q_N(_06350_),
    .Q(\u_toplayer.u_layer2.u_neuron.acc[2] ));
 sg13g2_dfrbp_1 _13434_ (.CLK(clknet_leaf_49_clk_regs),
    .RESET_B(net3551),
    .D(_00680_),
    .Q_N(_06349_),
    .Q(\u_toplayer.u_layer2.u_neuron.acc[3] ));
 sg13g2_dfrbp_1 _13435_ (.CLK(clknet_leaf_49_clk_regs),
    .RESET_B(net3514),
    .D(_00681_),
    .Q_N(_06348_),
    .Q(\u_toplayer.u_layer2.u_neuron.acc[4] ));
 sg13g2_dfrbp_1 _13436_ (.CLK(clknet_leaf_50_clk_regs),
    .RESET_B(net3514),
    .D(_00682_),
    .Q_N(_06347_),
    .Q(\u_toplayer.u_layer2.u_neuron.acc[5] ));
 sg13g2_dfrbp_1 _13437_ (.CLK(clknet_leaf_49_clk_regs),
    .RESET_B(net3508),
    .D(_00683_),
    .Q_N(_06346_),
    .Q(\u_toplayer.u_layer2.u_neuron.acc[6] ));
 sg13g2_dfrbp_1 _13438_ (.CLK(clknet_leaf_50_clk_regs),
    .RESET_B(net3508),
    .D(_00684_),
    .Q_N(_06345_),
    .Q(\u_toplayer.u_layer2.u_neuron.acc[7] ));
 sg13g2_dfrbp_1 _13439_ (.CLK(clknet_leaf_90_clk_regs),
    .RESET_B(net3509),
    .D(_00685_),
    .Q_N(_06344_),
    .Q(\u_toplayer.u_layer2.u_neuron.acc[8] ));
 sg13g2_dfrbp_1 _13440_ (.CLK(clknet_leaf_90_clk_regs),
    .RESET_B(net3508),
    .D(_00686_),
    .Q_N(_06343_),
    .Q(\u_toplayer.u_layer2.u_neuron.acc[9] ));
 sg13g2_dfrbp_1 _13441_ (.CLK(clknet_leaf_91_clk_regs),
    .RESET_B(net3508),
    .D(_00687_),
    .Q_N(_06342_),
    .Q(\u_toplayer.u_layer2.u_neuron.acc[10] ));
 sg13g2_dfrbp_1 _13442_ (.CLK(clknet_leaf_91_clk_regs),
    .RESET_B(net3454),
    .D(_00688_),
    .Q_N(_06341_),
    .Q(\u_toplayer.u_layer2.u_neuron.acc[11] ));
 sg13g2_dfrbp_1 _13443_ (.CLK(clknet_leaf_91_clk_regs),
    .RESET_B(net3508),
    .D(_00689_),
    .Q_N(_06340_),
    .Q(\u_toplayer.u_layer2.u_neuron.acc[12] ));
 sg13g2_dfrbp_1 _13444_ (.CLK(clknet_leaf_92_clk_regs),
    .RESET_B(net3507),
    .D(_00690_),
    .Q_N(_06339_),
    .Q(\u_toplayer.u_layer2.u_neuron.acc[13] ));
 sg13g2_dfrbp_1 _13445_ (.CLK(clknet_leaf_92_clk_regs),
    .RESET_B(net3507),
    .D(_00691_),
    .Q_N(_06338_),
    .Q(\u_toplayer.u_layer2.u_neuron.acc[14] ));
 sg13g2_dfrbp_1 _13446_ (.CLK(clknet_leaf_92_clk_regs),
    .RESET_B(net3506),
    .D(_00692_),
    .Q_N(_06337_),
    .Q(\u_toplayer.u_layer2.u_neuron.acc[15] ));
 sg13g2_dfrbp_1 _13447_ (.CLK(clknet_4_12_0_clk_regs),
    .RESET_B(net3507),
    .D(_00693_),
    .Q_N(_06336_),
    .Q(\u_toplayer.u_layer2.u_neuron.acc[16] ));
 sg13g2_dfrbp_1 _13448_ (.CLK(clknet_leaf_93_clk_regs),
    .RESET_B(net3507),
    .D(net1105),
    .Q_N(_06335_),
    .Q(\u_toplayer.u_layer2.u_neuron.acc[17] ));
 sg13g2_dfrbp_1 _13449_ (.CLK(clknet_leaf_88_clk_regs),
    .RESET_B(net3507),
    .D(net1169),
    .Q_N(_06334_),
    .Q(\u_toplayer.u_layer2.u_neuron.acc[18] ));
 sg13g2_dfrbp_1 _13450_ (.CLK(clknet_leaf_88_clk_regs),
    .RESET_B(net3507),
    .D(_00696_),
    .Q_N(_06333_),
    .Q(\u_toplayer.u_layer2.u_neuron.acc[19] ));
 sg13g2_dfrbp_1 _13451_ (.CLK(clknet_leaf_87_clk_regs),
    .RESET_B(net3511),
    .D(_00697_),
    .Q_N(_06332_),
    .Q(\u_toplayer.u_layer2.u_neuron.acc[20] ));
 sg13g2_dfrbp_1 _13452_ (.CLK(clknet_leaf_87_clk_regs),
    .RESET_B(net3511),
    .D(_00698_),
    .Q_N(_06331_),
    .Q(\u_toplayer.u_layer2.u_neuron.acc[21] ));
 sg13g2_dfrbp_1 _13453_ (.CLK(clknet_leaf_90_clk_regs),
    .RESET_B(net3509),
    .D(_00699_),
    .Q_N(_06330_),
    .Q(\u_toplayer.u_layer2.u_neuron.acc[22] ));
 sg13g2_dfrbp_1 _13454_ (.CLK(clknet_leaf_90_clk_regs),
    .RESET_B(net3512),
    .D(_00700_),
    .Q_N(_06329_),
    .Q(\u_toplayer.u_layer2.u_neuron.acc[23] ));
 sg13g2_dfrbp_1 _13455_ (.CLK(clknet_leaf_109_clk_regs),
    .RESET_B(net3409),
    .D(net598),
    .Q_N(_00050_),
    .Q(\u_toplayer.u_layer1.neuron_index[0] ));
 sg13g2_dfrbp_1 _13456_ (.CLK(clknet_leaf_109_clk_regs),
    .RESET_B(net3409),
    .D(_00702_),
    .Q_N(_06328_),
    .Q(\u_toplayer.u_layer1.neuron_index[1] ));
 sg13g2_dfrbp_1 _13457_ (.CLK(clknet_leaf_109_clk_regs),
    .RESET_B(net3409),
    .D(_00703_),
    .Q_N(_06327_),
    .Q(\u_toplayer.u_layer1.neuron_index[2] ));
 sg13g2_dfrbp_1 _13458_ (.CLK(clknet_leaf_108_clk_regs),
    .RESET_B(net3409),
    .D(_00704_),
    .Q_N(_06326_),
    .Q(\u_toplayer.u_layer1.neuron_index[3] ));
 sg13g2_dfrbp_1 _13459_ (.CLK(clknet_leaf_108_clk_regs),
    .RESET_B(net3409),
    .D(net1029),
    .Q_N(_06325_),
    .Q(\u_toplayer.u_layer1.neuron_index[4] ));
 sg13g2_dfrbp_1 _13460_ (.CLK(clknet_leaf_108_clk_regs),
    .RESET_B(net3434),
    .D(net1011),
    .Q_N(_06324_),
    .Q(\u_toplayer.u_layer1.neuron_index[5] ));
 sg13g2_dfrbp_1 _13461_ (.CLK(clknet_leaf_20_clk_regs),
    .RESET_B(net3417),
    .D(net127),
    .Q_N(_06323_),
    .Q(\u_toplayer.delay_counter_layer3[0] ));
 sg13g2_dfrbp_1 _13462_ (.CLK(clknet_leaf_20_clk_regs),
    .RESET_B(net3417),
    .D(_00708_),
    .Q_N(_06884_),
    .Q(\u_toplayer.delay_counter_layer3[1] ));
 sg13g2_dfrbp_1 _13463_ (.CLK(clknet_leaf_110_clk_regs),
    .RESET_B(net3408),
    .D(_00012_),
    .Q_N(_06322_),
    .Q(\u_toplayer.done_layer1 ));
 sg13g2_dfrbp_1 _13464_ (.CLK(clknet_leaf_14_clk_regs),
    .RESET_B(net3446),
    .D(_00709_),
    .Q_N(_06321_),
    .Q(\u_toplayer.reg_layer1[0] ));
 sg13g2_dfrbp_1 _13465_ (.CLK(clknet_leaf_14_clk_regs),
    .RESET_B(net3449),
    .D(_00710_),
    .Q_N(_06320_),
    .Q(\u_toplayer.reg_layer1[1] ));
 sg13g2_dfrbp_1 _13466_ (.CLK(clknet_leaf_95_clk_regs),
    .RESET_B(net3451),
    .D(_00711_),
    .Q_N(_06319_),
    .Q(\u_toplayer.reg_layer1[2] ));
 sg13g2_dfrbp_1 _13467_ (.CLK(clknet_leaf_16_clk_regs),
    .RESET_B(net3453),
    .D(_00712_),
    .Q_N(_06318_),
    .Q(\u_toplayer.reg_layer1[3] ));
 sg13g2_dfrbp_1 _13468_ (.CLK(clknet_leaf_95_clk_regs),
    .RESET_B(net3451),
    .D(_00713_),
    .Q_N(_06317_),
    .Q(\u_toplayer.reg_layer1[4] ));
 sg13g2_dfrbp_1 _13469_ (.CLK(clknet_leaf_95_clk_regs),
    .RESET_B(net3446),
    .D(_00714_),
    .Q_N(_06316_),
    .Q(\u_toplayer.reg_layer1[5] ));
 sg13g2_dfrbp_1 _13470_ (.CLK(clknet_leaf_14_clk_regs),
    .RESET_B(net3449),
    .D(_00715_),
    .Q_N(_06315_),
    .Q(\u_toplayer.reg_layer1[6] ));
 sg13g2_dfrbp_1 _13471_ (.CLK(clknet_leaf_15_clk_regs),
    .RESET_B(net3448),
    .D(_00716_),
    .Q_N(_06314_),
    .Q(\u_toplayer.reg_layer1[7] ));
 sg13g2_dfrbp_1 _13472_ (.CLK(clknet_leaf_13_clk_regs),
    .RESET_B(net3447),
    .D(_00717_),
    .Q_N(_06313_),
    .Q(\u_toplayer.reg_layer1[8] ));
 sg13g2_dfrbp_1 _13473_ (.CLK(clknet_leaf_15_clk_regs),
    .RESET_B(net3448),
    .D(_00718_),
    .Q_N(_06312_),
    .Q(\u_toplayer.reg_layer1[9] ));
 sg13g2_dfrbp_1 _13474_ (.CLK(clknet_leaf_14_clk_regs),
    .RESET_B(net3447),
    .D(net263),
    .Q_N(_06311_),
    .Q(\u_toplayer.reg_layer1[10] ));
 sg13g2_dfrbp_1 _13475_ (.CLK(clknet_leaf_14_clk_regs),
    .RESET_B(net3449),
    .D(_00720_),
    .Q_N(_06310_),
    .Q(\u_toplayer.reg_layer1[11] ));
 sg13g2_dfrbp_1 _13476_ (.CLK(clknet_leaf_13_clk_regs),
    .RESET_B(net3446),
    .D(_00721_),
    .Q_N(_06309_),
    .Q(\u_toplayer.reg_layer1[12] ));
 sg13g2_dfrbp_1 _13477_ (.CLK(clknet_leaf_13_clk_regs),
    .RESET_B(net3446),
    .D(net287),
    .Q_N(_06308_),
    .Q(\u_toplayer.reg_layer1[13] ));
 sg13g2_dfrbp_1 _13478_ (.CLK(clknet_leaf_10_clk_regs),
    .RESET_B(net3448),
    .D(_00723_),
    .Q_N(_06307_),
    .Q(\u_toplayer.reg_layer1[14] ));
 sg13g2_dfrbp_1 _13479_ (.CLK(clknet_leaf_10_clk_regs),
    .RESET_B(net3448),
    .D(_00724_),
    .Q_N(_06306_),
    .Q(\u_toplayer.reg_layer1[15] ));
 sg13g2_dfrbp_1 _13480_ (.CLK(clknet_leaf_8_clk_regs),
    .RESET_B(net3416),
    .D(_00725_),
    .Q_N(_06305_),
    .Q(\u_toplayer.reg_layer1[16] ));
 sg13g2_dfrbp_1 _13481_ (.CLK(clknet_leaf_9_clk_regs),
    .RESET_B(net3424),
    .D(_00726_),
    .Q_N(_06304_),
    .Q(\u_toplayer.reg_layer1[17] ));
 sg13g2_dfrbp_1 _13482_ (.CLK(clknet_leaf_5_clk_regs),
    .RESET_B(net3418),
    .D(_00727_),
    .Q_N(_06303_),
    .Q(\u_toplayer.reg_layer1[18] ));
 sg13g2_dfrbp_1 _13483_ (.CLK(clknet_leaf_11_clk_regs),
    .RESET_B(net3424),
    .D(_00728_),
    .Q_N(_06302_),
    .Q(\u_toplayer.reg_layer1[19] ));
 sg13g2_dfrbp_1 _13484_ (.CLK(clknet_leaf_11_clk_regs),
    .RESET_B(net3418),
    .D(_00729_),
    .Q_N(_06301_),
    .Q(\u_toplayer.reg_layer1[20] ));
 sg13g2_dfrbp_1 _13485_ (.CLK(clknet_leaf_11_clk_regs),
    .RESET_B(net3420),
    .D(_00730_),
    .Q_N(_06300_),
    .Q(\u_toplayer.reg_layer1[21] ));
 sg13g2_dfrbp_1 _13486_ (.CLK(clknet_leaf_9_clk_regs),
    .RESET_B(net3422),
    .D(_00731_),
    .Q_N(_06299_),
    .Q(\u_toplayer.reg_layer1[22] ));
 sg13g2_dfrbp_1 _13487_ (.CLK(clknet_leaf_9_clk_regs),
    .RESET_B(net3422),
    .D(_00732_),
    .Q_N(_06298_),
    .Q(\u_toplayer.reg_layer1[23] ));
 sg13g2_dfrbp_1 _13488_ (.CLK(clknet_leaf_8_clk_regs),
    .RESET_B(net3416),
    .D(_00733_),
    .Q_N(_06297_),
    .Q(\u_toplayer.reg_layer1[24] ));
 sg13g2_dfrbp_1 _13489_ (.CLK(clknet_leaf_10_clk_regs),
    .RESET_B(net3424),
    .D(_00734_),
    .Q_N(_06296_),
    .Q(\u_toplayer.reg_layer1[25] ));
 sg13g2_dfrbp_1 _13490_ (.CLK(clknet_leaf_5_clk_regs),
    .RESET_B(net3418),
    .D(_00735_),
    .Q_N(_06295_),
    .Q(\u_toplayer.reg_layer1[26] ));
 sg13g2_dfrbp_1 _13491_ (.CLK(clknet_leaf_11_clk_regs),
    .RESET_B(net3424),
    .D(_00736_),
    .Q_N(_06294_),
    .Q(\u_toplayer.reg_layer1[27] ));
 sg13g2_dfrbp_1 _13492_ (.CLK(clknet_leaf_5_clk_regs),
    .RESET_B(net3418),
    .D(_00737_),
    .Q_N(_06293_),
    .Q(\u_toplayer.reg_layer1[28] ));
 sg13g2_dfrbp_1 _13493_ (.CLK(clknet_leaf_12_clk_regs),
    .RESET_B(net3419),
    .D(_00738_),
    .Q_N(_06292_),
    .Q(\u_toplayer.reg_layer1[29] ));
 sg13g2_dfrbp_1 _13494_ (.CLK(clknet_leaf_9_clk_regs),
    .RESET_B(net3422),
    .D(_00739_),
    .Q_N(_06291_),
    .Q(\u_toplayer.reg_layer1[30] ));
 sg13g2_dfrbp_1 _13495_ (.CLK(clknet_leaf_9_clk_regs),
    .RESET_B(net3422),
    .D(_00740_),
    .Q_N(_06290_),
    .Q(\u_toplayer.reg_layer1[31] ));
 sg13g2_dfrbp_1 _13496_ (.CLK(clknet_leaf_0_clk_regs),
    .RESET_B(net3407),
    .D(_00741_),
    .Q_N(_06289_),
    .Q(\u_toplayer.reg_layer1[32] ));
 sg13g2_dfrbp_1 _13497_ (.CLK(clknet_leaf_1_clk_regs),
    .RESET_B(net3405),
    .D(_00742_),
    .Q_N(_06288_),
    .Q(\u_toplayer.reg_layer1[33] ));
 sg13g2_dfrbp_1 _13498_ (.CLK(clknet_leaf_2_clk_regs),
    .RESET_B(net3411),
    .D(_00743_),
    .Q_N(_06287_),
    .Q(\u_toplayer.reg_layer1[34] ));
 sg13g2_dfrbp_1 _13499_ (.CLK(clknet_leaf_2_clk_regs),
    .RESET_B(net3411),
    .D(_00744_),
    .Q_N(_06286_),
    .Q(\u_toplayer.reg_layer1[35] ));
 sg13g2_dfrbp_1 _13500_ (.CLK(clknet_leaf_108_clk_regs),
    .RESET_B(net3413),
    .D(_00745_),
    .Q_N(_06285_),
    .Q(\u_toplayer.reg_layer1[36] ));
 sg13g2_dfrbp_1 _13501_ (.CLK(clknet_leaf_3_clk_regs),
    .RESET_B(net3411),
    .D(_00746_),
    .Q_N(_06284_),
    .Q(\u_toplayer.reg_layer1[37] ));
 sg13g2_dfrbp_1 _13502_ (.CLK(clknet_leaf_1_clk_regs),
    .RESET_B(net3406),
    .D(_00747_),
    .Q_N(_06283_),
    .Q(\u_toplayer.reg_layer1[38] ));
 sg13g2_dfrbp_1 _13503_ (.CLK(clknet_leaf_1_clk_regs),
    .RESET_B(net3405),
    .D(_00748_),
    .Q_N(_06282_),
    .Q(\u_toplayer.reg_layer1[39] ));
 sg13g2_dfrbp_1 _13504_ (.CLK(clknet_leaf_0_clk_regs),
    .RESET_B(net3407),
    .D(_00749_),
    .Q_N(_06281_),
    .Q(\u_toplayer.reg_layer1[40] ));
 sg13g2_dfrbp_1 _13505_ (.CLK(clknet_leaf_2_clk_regs),
    .RESET_B(net3407),
    .D(_00750_),
    .Q_N(_06280_),
    .Q(\u_toplayer.reg_layer1[41] ));
 sg13g2_dfrbp_1 _13506_ (.CLK(clknet_leaf_0_clk_regs),
    .RESET_B(net3410),
    .D(_00751_),
    .Q_N(_06279_),
    .Q(\u_toplayer.reg_layer1[42] ));
 sg13g2_dfrbp_1 _13507_ (.CLK(clknet_leaf_3_clk_regs),
    .RESET_B(net3410),
    .D(_00752_),
    .Q_N(_06278_),
    .Q(\u_toplayer.reg_layer1[43] ));
 sg13g2_dfrbp_1 _13508_ (.CLK(clknet_leaf_3_clk_regs),
    .RESET_B(net3410),
    .D(_00753_),
    .Q_N(_06277_),
    .Q(\u_toplayer.reg_layer1[44] ));
 sg13g2_dfrbp_1 _13509_ (.CLK(clknet_leaf_3_clk_regs),
    .RESET_B(net3413),
    .D(_00754_),
    .Q_N(_06276_),
    .Q(\u_toplayer.reg_layer1[45] ));
 sg13g2_dfrbp_1 _13510_ (.CLK(clknet_leaf_1_clk_regs),
    .RESET_B(net3405),
    .D(_00755_),
    .Q_N(_06275_),
    .Q(\u_toplayer.reg_layer1[46] ));
 sg13g2_dfrbp_1 _13511_ (.CLK(clknet_leaf_0_clk_regs),
    .RESET_B(net3405),
    .D(_00756_),
    .Q_N(_06274_),
    .Q(\u_toplayer.reg_layer1[47] ));
 sg13g2_dfrbp_1 _13512_ (.CLK(clknet_leaf_6_clk_regs),
    .RESET_B(net3406),
    .D(_00757_),
    .Q_N(_06273_),
    .Q(\u_toplayer.reg_layer1[48] ));
 sg13g2_dfrbp_1 _13513_ (.CLK(clknet_leaf_8_clk_regs),
    .RESET_B(net3415),
    .D(_00758_),
    .Q_N(_06272_),
    .Q(\u_toplayer.reg_layer1[49] ));
 sg13g2_dfrbp_1 _13514_ (.CLK(clknet_leaf_6_clk_regs),
    .RESET_B(net3412),
    .D(_00759_),
    .Q_N(_06271_),
    .Q(\u_toplayer.reg_layer1[50] ));
 sg13g2_dfrbp_1 _13515_ (.CLK(clknet_leaf_6_clk_regs),
    .RESET_B(net3412),
    .D(_00760_),
    .Q_N(_06270_),
    .Q(\u_toplayer.reg_layer1[51] ));
 sg13g2_dfrbp_1 _13516_ (.CLK(clknet_leaf_4_clk_regs),
    .RESET_B(net3413),
    .D(_00761_),
    .Q_N(_06269_),
    .Q(\u_toplayer.reg_layer1[52] ));
 sg13g2_dfrbp_1 _13517_ (.CLK(clknet_leaf_4_clk_regs),
    .RESET_B(net3419),
    .D(_00762_),
    .Q_N(_06268_),
    .Q(\u_toplayer.reg_layer1[53] ));
 sg13g2_dfrbp_1 _13518_ (.CLK(clknet_leaf_7_clk_regs),
    .RESET_B(net3415),
    .D(_00763_),
    .Q_N(_06267_),
    .Q(\u_toplayer.reg_layer1[54] ));
 sg13g2_dfrbp_1 _13519_ (.CLK(clknet_leaf_7_clk_regs),
    .RESET_B(net3415),
    .D(_00764_),
    .Q_N(_06266_),
    .Q(\u_toplayer.reg_layer1[55] ));
 sg13g2_dfrbp_1 _13520_ (.CLK(clknet_leaf_6_clk_regs),
    .RESET_B(net3406),
    .D(_00765_),
    .Q_N(_06265_),
    .Q(\u_toplayer.reg_layer1[56] ));
 sg13g2_dfrbp_1 _13521_ (.CLK(clknet_leaf_8_clk_regs),
    .RESET_B(net3416),
    .D(_00766_),
    .Q_N(_06264_),
    .Q(\u_toplayer.reg_layer1[57] ));
 sg13g2_dfrbp_1 _13522_ (.CLK(clknet_leaf_2_clk_regs),
    .RESET_B(net3412),
    .D(_00767_),
    .Q_N(_06263_),
    .Q(\u_toplayer.reg_layer1[58] ));
 sg13g2_dfrbp_1 _13523_ (.CLK(clknet_leaf_2_clk_regs),
    .RESET_B(net3411),
    .D(_00768_),
    .Q_N(_06262_),
    .Q(\u_toplayer.reg_layer1[59] ));
 sg13g2_dfrbp_1 _13524_ (.CLK(clknet_leaf_4_clk_regs),
    .RESET_B(net3413),
    .D(_00769_),
    .Q_N(_06261_),
    .Q(\u_toplayer.reg_layer1[60] ));
 sg13g2_dfrbp_1 _13525_ (.CLK(clknet_leaf_3_clk_regs),
    .RESET_B(net3414),
    .D(_00770_),
    .Q_N(_06260_),
    .Q(\u_toplayer.reg_layer1[61] ));
 sg13g2_dfrbp_1 _13526_ (.CLK(clknet_leaf_7_clk_regs),
    .RESET_B(net3406),
    .D(_00771_),
    .Q_N(_06259_),
    .Q(\u_toplayer.reg_layer1[62] ));
 sg13g2_dfrbp_1 _13527_ (.CLK(clknet_leaf_7_clk_regs),
    .RESET_B(net3415),
    .D(_00772_),
    .Q_N(_06258_),
    .Q(\u_toplayer.reg_layer1[63] ));
 sg13g2_dfrbp_1 _13528_ (.CLK(clknet_leaf_97_clk_regs),
    .RESET_B(net3440),
    .D(_00773_),
    .Q_N(_06257_),
    .Q(\u_toplayer.reg_layer1[64] ));
 sg13g2_dfrbp_1 _13529_ (.CLK(clknet_leaf_99_clk_regs),
    .RESET_B(net3493),
    .D(_00774_),
    .Q_N(_06256_),
    .Q(\u_toplayer.reg_layer1[65] ));
 sg13g2_dfrbp_1 _13530_ (.CLK(clknet_leaf_99_clk_regs),
    .RESET_B(net3493),
    .D(_00775_),
    .Q_N(_06255_),
    .Q(\u_toplayer.reg_layer1[66] ));
 sg13g2_dfrbp_1 _13531_ (.CLK(clknet_leaf_82_clk_regs),
    .RESET_B(net3493),
    .D(_00776_),
    .Q_N(_06254_),
    .Q(\u_toplayer.reg_layer1[67] ));
 sg13g2_dfrbp_1 _13532_ (.CLK(clknet_leaf_99_clk_regs),
    .RESET_B(net3441),
    .D(_00777_),
    .Q_N(_06253_),
    .Q(\u_toplayer.reg_layer1[68] ));
 sg13g2_dfrbp_1 _13533_ (.CLK(clknet_leaf_97_clk_regs),
    .RESET_B(net3440),
    .D(net377),
    .Q_N(_06252_),
    .Q(\u_toplayer.reg_layer1[69] ));
 sg13g2_dfrbp_1 _13534_ (.CLK(clknet_leaf_97_clk_regs),
    .RESET_B(net3442),
    .D(_00779_),
    .Q_N(_06251_),
    .Q(\u_toplayer.reg_layer1[70] ));
 sg13g2_dfrbp_1 _13535_ (.CLK(clknet_leaf_82_clk_regs),
    .RESET_B(net3494),
    .D(net515),
    .Q_N(_06250_),
    .Q(\u_toplayer.reg_layer1[71] ));
 sg13g2_dfrbp_1 _13536_ (.CLK(clknet_leaf_97_clk_regs),
    .RESET_B(net3440),
    .D(net352),
    .Q_N(_06249_),
    .Q(\u_toplayer.reg_layer1[72] ));
 sg13g2_dfrbp_1 _13537_ (.CLK(clknet_leaf_100_clk_regs),
    .RESET_B(net3488),
    .D(net452),
    .Q_N(_06248_),
    .Q(\u_toplayer.reg_layer1[73] ));
 sg13g2_dfrbp_1 _13538_ (.CLK(clknet_leaf_80_clk_regs),
    .RESET_B(net3489),
    .D(_00783_),
    .Q_N(_06247_),
    .Q(\u_toplayer.reg_layer1[74] ));
 sg13g2_dfrbp_1 _13539_ (.CLK(clknet_leaf_80_clk_regs),
    .RESET_B(net3489),
    .D(_00784_),
    .Q_N(_06246_),
    .Q(\u_toplayer.reg_layer1[75] ));
 sg13g2_dfrbp_1 _13540_ (.CLK(clknet_leaf_100_clk_regs),
    .RESET_B(net3438),
    .D(_00785_),
    .Q_N(_06245_),
    .Q(\u_toplayer.reg_layer1[76] ));
 sg13g2_dfrbp_1 _13541_ (.CLK(clknet_leaf_99_clk_regs),
    .RESET_B(net3441),
    .D(net712),
    .Q_N(_06244_),
    .Q(\u_toplayer.reg_layer1[77] ));
 sg13g2_dfrbp_1 _13542_ (.CLK(clknet_leaf_100_clk_regs),
    .RESET_B(net3438),
    .D(_00787_),
    .Q_N(_06243_),
    .Q(\u_toplayer.reg_layer1[78] ));
 sg13g2_dfrbp_1 _13543_ (.CLK(clknet_leaf_81_clk_regs),
    .RESET_B(net3493),
    .D(net572),
    .Q_N(_06242_),
    .Q(\u_toplayer.reg_layer1[79] ));
 sg13g2_dfrbp_1 _13544_ (.CLK(clknet_leaf_95_clk_regs),
    .RESET_B(net3450),
    .D(_00789_),
    .Q_N(_06241_),
    .Q(\u_toplayer.reg_layer1[80] ));
 sg13g2_dfrbp_1 _13545_ (.CLK(clknet_leaf_93_clk_regs),
    .RESET_B(net3452),
    .D(_00790_),
    .Q_N(_06240_),
    .Q(\u_toplayer.reg_layer1[81] ));
 sg13g2_dfrbp_1 _13546_ (.CLK(clknet_leaf_94_clk_regs),
    .RESET_B(net3452),
    .D(_00791_),
    .Q_N(_06239_),
    .Q(\u_toplayer.reg_layer1[82] ));
 sg13g2_dfrbp_1 _13547_ (.CLK(clknet_leaf_98_clk_regs),
    .RESET_B(net3506),
    .D(_00792_),
    .Q_N(_06238_),
    .Q(\u_toplayer.reg_layer1[83] ));
 sg13g2_dfrbp_1 _13548_ (.CLK(clknet_leaf_96_clk_regs),
    .RESET_B(net3433),
    .D(_00793_),
    .Q_N(_06237_),
    .Q(\u_toplayer.reg_layer1[84] ));
 sg13g2_dfrbp_1 _13549_ (.CLK(clknet_leaf_94_clk_regs),
    .RESET_B(net3450),
    .D(_00794_),
    .Q_N(_06236_),
    .Q(\u_toplayer.reg_layer1[85] ));
 sg13g2_dfrbp_1 _13550_ (.CLK(clknet_leaf_96_clk_regs),
    .RESET_B(net3446),
    .D(_00795_),
    .Q_N(_06235_),
    .Q(\u_toplayer.reg_layer1[86] ));
 sg13g2_dfrbp_1 _13551_ (.CLK(clknet_leaf_93_clk_regs),
    .RESET_B(net3452),
    .D(net574),
    .Q_N(_06234_),
    .Q(\u_toplayer.reg_layer1[87] ));
 sg13g2_dfrbp_1 _13552_ (.CLK(clknet_leaf_95_clk_regs),
    .RESET_B(net3450),
    .D(_00797_),
    .Q_N(_06233_),
    .Q(\u_toplayer.reg_layer1[88] ));
 sg13g2_dfrbp_1 _13553_ (.CLK(clknet_leaf_93_clk_regs),
    .RESET_B(net3441),
    .D(_00798_),
    .Q_N(_06232_),
    .Q(\u_toplayer.reg_layer1[89] ));
 sg13g2_dfrbp_1 _13554_ (.CLK(clknet_leaf_93_clk_regs),
    .RESET_B(net3452),
    .D(_00799_),
    .Q_N(_06231_),
    .Q(\u_toplayer.reg_layer1[90] ));
 sg13g2_dfrbp_1 _13555_ (.CLK(clknet_leaf_98_clk_regs),
    .RESET_B(net3494),
    .D(_00800_),
    .Q_N(_06230_),
    .Q(\u_toplayer.reg_layer1[91] ));
 sg13g2_dfrbp_1 _13556_ (.CLK(clknet_leaf_96_clk_regs),
    .RESET_B(net3442),
    .D(net784),
    .Q_N(_06229_),
    .Q(\u_toplayer.reg_layer1[92] ));
 sg13g2_dfrbp_1 _13557_ (.CLK(clknet_leaf_94_clk_regs),
    .RESET_B(net3450),
    .D(_00802_),
    .Q_N(_06228_),
    .Q(\u_toplayer.reg_layer1[93] ));
 sg13g2_dfrbp_1 _13558_ (.CLK(clknet_leaf_96_clk_regs),
    .RESET_B(net3450),
    .D(_00803_),
    .Q_N(_06227_),
    .Q(\u_toplayer.reg_layer1[94] ));
 sg13g2_dfrbp_1 _13559_ (.CLK(clknet_leaf_93_clk_regs),
    .RESET_B(net3506),
    .D(net700),
    .Q_N(_06226_),
    .Q(\u_toplayer.reg_layer1[95] ));
 sg13g2_dfrbp_1 _13560_ (.CLK(clknet_leaf_106_clk_regs),
    .RESET_B(net3432),
    .D(net366),
    .Q_N(_06225_),
    .Q(\u_toplayer.reg_layer1[96] ));
 sg13g2_dfrbp_1 _13561_ (.CLK(clknet_leaf_102_clk_regs),
    .RESET_B(net3436),
    .D(_00806_),
    .Q_N(_06224_),
    .Q(\u_toplayer.reg_layer1[97] ));
 sg13g2_dfrbp_1 _13562_ (.CLK(clknet_leaf_103_clk_regs),
    .RESET_B(net3435),
    .D(_00807_),
    .Q_N(_06223_),
    .Q(\u_toplayer.reg_layer1[98] ));
 sg13g2_dfrbp_1 _13563_ (.CLK(clknet_leaf_103_clk_regs),
    .RESET_B(net3435),
    .D(_00808_),
    .Q_N(_06222_),
    .Q(\u_toplayer.reg_layer1[99] ));
 sg13g2_dfrbp_1 _13564_ (.CLK(clknet_leaf_104_clk_regs),
    .RESET_B(net3429),
    .D(_00809_),
    .Q_N(_06221_),
    .Q(\u_toplayer.reg_layer1[100] ));
 sg13g2_dfrbp_1 _13565_ (.CLK(clknet_leaf_104_clk_regs),
    .RESET_B(net3429),
    .D(_00810_),
    .Q_N(_06220_),
    .Q(\u_toplayer.reg_layer1[101] ));
 sg13g2_dfrbp_1 _13566_ (.CLK(clknet_leaf_106_clk_regs),
    .RESET_B(net3432),
    .D(net299),
    .Q_N(_06219_),
    .Q(\u_toplayer.reg_layer1[102] ));
 sg13g2_dfrbp_1 _13567_ (.CLK(clknet_leaf_106_clk_regs),
    .RESET_B(net3430),
    .D(net312),
    .Q_N(_06218_),
    .Q(\u_toplayer.reg_layer1[103] ));
 sg13g2_dfrbp_1 _13568_ (.CLK(clknet_leaf_102_clk_regs),
    .RESET_B(net3436),
    .D(_00813_),
    .Q_N(_06217_),
    .Q(\u_toplayer.reg_layer1[104] ));
 sg13g2_dfrbp_1 _13569_ (.CLK(clknet_leaf_101_clk_regs),
    .RESET_B(net3437),
    .D(_00814_),
    .Q_N(_06216_),
    .Q(\u_toplayer.reg_layer1[105] ));
 sg13g2_dfrbp_1 _13570_ (.CLK(clknet_leaf_101_clk_regs),
    .RESET_B(net3437),
    .D(net624),
    .Q_N(_06215_),
    .Q(\u_toplayer.reg_layer1[106] ));
 sg13g2_dfrbp_1 _13571_ (.CLK(clknet_leaf_101_clk_regs),
    .RESET_B(net3437),
    .D(net689),
    .Q_N(_06214_),
    .Q(\u_toplayer.reg_layer1[107] ));
 sg13g2_dfrbp_1 _13572_ (.CLK(clknet_leaf_102_clk_regs),
    .RESET_B(net3435),
    .D(net756),
    .Q_N(_06213_),
    .Q(\u_toplayer.reg_layer1[108] ));
 sg13g2_dfrbp_1 _13573_ (.CLK(clknet_leaf_101_clk_regs),
    .RESET_B(net3437),
    .D(_00818_),
    .Q_N(_06212_),
    .Q(\u_toplayer.reg_layer1[109] ));
 sg13g2_dfrbp_1 _13574_ (.CLK(clknet_leaf_103_clk_regs),
    .RESET_B(net3440),
    .D(net775),
    .Q_N(_06211_),
    .Q(\u_toplayer.reg_layer1[110] ));
 sg13g2_dfrbp_1 _13575_ (.CLK(clknet_leaf_102_clk_regs),
    .RESET_B(net3435),
    .D(net279),
    .Q_N(_06210_),
    .Q(\u_toplayer.reg_layer1[111] ));
 sg13g2_dfrbp_1 _13576_ (.CLK(clknet_leaf_107_clk_regs),
    .RESET_B(net3433),
    .D(_00821_),
    .Q_N(_06209_),
    .Q(\u_toplayer.reg_layer1[112] ));
 sg13g2_dfrbp_1 _13577_ (.CLK(clknet_leaf_105_clk_regs),
    .RESET_B(net3432),
    .D(net417),
    .Q_N(_06208_),
    .Q(\u_toplayer.reg_layer1[113] ));
 sg13g2_dfrbp_1 _13578_ (.CLK(clknet_leaf_104_clk_regs),
    .RESET_B(net3428),
    .D(net246),
    .Q_N(_06207_),
    .Q(\u_toplayer.reg_layer1[114] ));
 sg13g2_dfrbp_1 _13579_ (.CLK(clknet_leaf_104_clk_regs),
    .RESET_B(net3429),
    .D(net424),
    .Q_N(_06206_),
    .Q(\u_toplayer.reg_layer1[115] ));
 sg13g2_dfrbp_1 _13580_ (.CLK(clknet_leaf_105_clk_regs),
    .RESET_B(net3430),
    .D(net749),
    .Q_N(_06205_),
    .Q(\u_toplayer.reg_layer1[116] ));
 sg13g2_dfrbp_1 _13581_ (.CLK(clknet_leaf_110_clk_regs),
    .RESET_B(net3428),
    .D(net553),
    .Q_N(_06204_),
    .Q(\u_toplayer.reg_layer1[117] ));
 sg13g2_dfrbp_1 _13582_ (.CLK(clknet_leaf_108_clk_regs),
    .RESET_B(net3434),
    .D(_00827_),
    .Q_N(_06203_),
    .Q(\u_toplayer.reg_layer1[118] ));
 sg13g2_dfrbp_1 _13583_ (.CLK(clknet_leaf_109_clk_regs),
    .RESET_B(net3431),
    .D(net464),
    .Q_N(_06202_),
    .Q(\u_toplayer.reg_layer1[119] ));
 sg13g2_dfrbp_1 _13584_ (.CLK(clknet_leaf_107_clk_regs),
    .RESET_B(net3432),
    .D(_00829_),
    .Q_N(_06201_),
    .Q(\u_toplayer.reg_layer1[120] ));
 sg13g2_dfrbp_1 _13585_ (.CLK(clknet_leaf_105_clk_regs),
    .RESET_B(net3430),
    .D(net180),
    .Q_N(_06200_),
    .Q(\u_toplayer.reg_layer1[121] ));
 sg13g2_dfrbp_1 _13586_ (.CLK(clknet_leaf_104_clk_regs),
    .RESET_B(net3428),
    .D(_00831_),
    .Q_N(_06199_),
    .Q(\u_toplayer.reg_layer1[122] ));
 sg13g2_dfrbp_1 _13587_ (.CLK(clknet_leaf_104_clk_regs),
    .RESET_B(net3429),
    .D(_00832_),
    .Q_N(_06198_),
    .Q(\u_toplayer.reg_layer1[123] ));
 sg13g2_dfrbp_1 _13588_ (.CLK(clknet_leaf_105_clk_regs),
    .RESET_B(net3429),
    .D(_00833_),
    .Q_N(_06197_),
    .Q(\u_toplayer.reg_layer1[124] ));
 sg13g2_dfrbp_1 _13589_ (.CLK(clknet_leaf_110_clk_regs),
    .RESET_B(net3428),
    .D(_00834_),
    .Q_N(_06196_),
    .Q(\u_toplayer.reg_layer1[125] ));
 sg13g2_dfrbp_1 _13590_ (.CLK(clknet_leaf_107_clk_regs),
    .RESET_B(net3434),
    .D(_00835_),
    .Q_N(_06195_),
    .Q(\u_toplayer.reg_layer1[126] ));
 sg13g2_dfrbp_1 _13591_ (.CLK(clknet_leaf_109_clk_regs),
    .RESET_B(net3431),
    .D(_00836_),
    .Q_N(_06194_),
    .Q(\u_toplayer.reg_layer1[127] ));
 sg13g2_dfrbp_1 _13592_ (.CLK(clknet_leaf_12_clk_regs),
    .RESET_B(net3444),
    .D(_00837_),
    .Q_N(_06193_),
    .Q(\u_toplayer.reg_layer1[128] ));
 sg13g2_dfrbp_1 _13593_ (.CLK(clknet_leaf_10_clk_regs),
    .RESET_B(net3445),
    .D(_00838_),
    .Q_N(_06192_),
    .Q(\u_toplayer.reg_layer1[129] ));
 sg13g2_dfrbp_1 _13594_ (.CLK(clknet_leaf_12_clk_regs),
    .RESET_B(net3444),
    .D(_00839_),
    .Q_N(_06191_),
    .Q(\u_toplayer.reg_layer1[130] ));
 sg13g2_dfrbp_1 _13595_ (.CLK(clknet_leaf_13_clk_regs),
    .RESET_B(net3445),
    .D(_00840_),
    .Q_N(_06190_),
    .Q(\u_toplayer.reg_layer1[131] ));
 sg13g2_dfrbp_1 _13596_ (.CLK(clknet_leaf_107_clk_regs),
    .RESET_B(net3434),
    .D(net518),
    .Q_N(_06189_),
    .Q(\u_toplayer.reg_layer1[132] ));
 sg13g2_dfrbp_1 _13597_ (.CLK(clknet_leaf_12_clk_regs),
    .RESET_B(net3444),
    .D(_00842_),
    .Q_N(_06188_),
    .Q(\u_toplayer.reg_layer1[133] ));
 sg13g2_dfrbp_1 _13598_ (.CLK(clknet_leaf_12_clk_regs),
    .RESET_B(net3445),
    .D(net715),
    .Q_N(_06187_),
    .Q(\u_toplayer.reg_layer1[134] ));
 sg13g2_dfrbp_1 _13599_ (.CLK(clknet_leaf_12_clk_regs),
    .RESET_B(net3420),
    .D(_00844_),
    .Q_N(_06186_),
    .Q(\u_toplayer.reg_layer1[135] ));
 sg13g2_dfrbp_1 _13600_ (.CLK(clknet_leaf_13_clk_regs),
    .RESET_B(net3444),
    .D(_00845_),
    .Q_N(_06185_),
    .Q(\u_toplayer.reg_layer1[136] ));
 sg13g2_dfrbp_1 _13601_ (.CLK(clknet_leaf_14_clk_regs),
    .RESET_B(net3444),
    .D(_00846_),
    .Q_N(_06184_),
    .Q(\u_toplayer.reg_layer1[137] ));
 sg13g2_dfrbp_1 _13602_ (.CLK(clknet_leaf_13_clk_regs),
    .RESET_B(net3446),
    .D(net739),
    .Q_N(_06183_),
    .Q(\u_toplayer.reg_layer1[138] ));
 sg13g2_dfrbp_1 _13603_ (.CLK(clknet_leaf_13_clk_regs),
    .RESET_B(net3444),
    .D(_00848_),
    .Q_N(_06182_),
    .Q(\u_toplayer.reg_layer1[139] ));
 sg13g2_dfrbp_1 _13604_ (.CLK(clknet_leaf_13_clk_regs),
    .RESET_B(net3444),
    .D(_00849_),
    .Q_N(_06181_),
    .Q(\u_toplayer.reg_layer1[140] ));
 sg13g2_dfrbp_1 _13605_ (.CLK(clknet_leaf_12_clk_regs),
    .RESET_B(net3444),
    .D(net800),
    .Q_N(_06180_),
    .Q(\u_toplayer.reg_layer1[141] ));
 sg13g2_dfrbp_1 _13606_ (.CLK(clknet_leaf_10_clk_regs),
    .RESET_B(net3448),
    .D(_00851_),
    .Q_N(_06179_),
    .Q(\u_toplayer.reg_layer1[142] ));
 sg13g2_dfrbp_1 _13607_ (.CLK(clknet_leaf_10_clk_regs),
    .RESET_B(net3445),
    .D(_00852_),
    .Q_N(_06178_),
    .Q(\u_toplayer.reg_layer1[143] ));
 sg13g2_dfrbp_1 _13608_ (.CLK(clknet_leaf_9_clk_regs),
    .RESET_B(net3416),
    .D(_00853_),
    .Q_N(_06177_),
    .Q(\u_toplayer.reg_layer1[144] ));
 sg13g2_dfrbp_1 _13609_ (.CLK(clknet_leaf_10_clk_regs),
    .RESET_B(net3424),
    .D(_00854_),
    .Q_N(_06176_),
    .Q(\u_toplayer.reg_layer1[145] ));
 sg13g2_dfrbp_1 _13610_ (.CLK(clknet_leaf_5_clk_regs),
    .RESET_B(net3418),
    .D(_00855_),
    .Q_N(_06175_),
    .Q(\u_toplayer.reg_layer1[146] ));
 sg13g2_dfrbp_1 _13611_ (.CLK(clknet_leaf_11_clk_regs),
    .RESET_B(net3420),
    .D(_00856_),
    .Q_N(_06174_),
    .Q(\u_toplayer.reg_layer1[147] ));
 sg13g2_dfrbp_1 _13612_ (.CLK(clknet_leaf_11_clk_regs),
    .RESET_B(net3419),
    .D(_00857_),
    .Q_N(_06173_),
    .Q(\u_toplayer.reg_layer1[148] ));
 sg13g2_dfrbp_1 _13613_ (.CLK(clknet_leaf_4_clk_regs),
    .RESET_B(net3419),
    .D(_00858_),
    .Q_N(_06172_),
    .Q(\u_toplayer.reg_layer1[149] ));
 sg13g2_dfrbp_1 _13614_ (.CLK(clknet_leaf_11_clk_regs),
    .RESET_B(net3418),
    .D(_00859_),
    .Q_N(_06171_),
    .Q(\u_toplayer.reg_layer1[150] ));
 sg13g2_dfrbp_1 _13615_ (.CLK(clknet_leaf_9_clk_regs),
    .RESET_B(net3421),
    .D(_00860_),
    .Q_N(_06170_),
    .Q(\u_toplayer.reg_layer1[151] ));
 sg13g2_dfrbp_1 _13616_ (.CLK(clknet_leaf_8_clk_regs),
    .RESET_B(net3416),
    .D(_00861_),
    .Q_N(_06169_),
    .Q(\u_toplayer.reg_layer1[152] ));
 sg13g2_dfrbp_1 _13617_ (.CLK(clknet_leaf_10_clk_regs),
    .RESET_B(net3424),
    .D(_00862_),
    .Q_N(_06168_),
    .Q(\u_toplayer.reg_layer1[153] ));
 sg13g2_dfrbp_1 _13618_ (.CLK(clknet_leaf_5_clk_regs),
    .RESET_B(net3418),
    .D(_00863_),
    .Q_N(_06167_),
    .Q(\u_toplayer.reg_layer1[154] ));
 sg13g2_dfrbp_1 _13619_ (.CLK(clknet_leaf_12_clk_regs),
    .RESET_B(net3420),
    .D(net235),
    .Q_N(_06166_),
    .Q(\u_toplayer.reg_layer1[155] ));
 sg13g2_dfrbp_1 _13620_ (.CLK(clknet_leaf_5_clk_regs),
    .RESET_B(net3419),
    .D(_00865_),
    .Q_N(_06165_),
    .Q(\u_toplayer.reg_layer1[156] ));
 sg13g2_dfrbp_1 _13621_ (.CLK(clknet_leaf_4_clk_regs),
    .RESET_B(net3419),
    .D(_00866_),
    .Q_N(_06164_),
    .Q(\u_toplayer.reg_layer1[157] ));
 sg13g2_dfrbp_1 _13622_ (.CLK(clknet_leaf_11_clk_regs),
    .RESET_B(net3418),
    .D(_00867_),
    .Q_N(_06163_),
    .Q(\u_toplayer.reg_layer1[158] ));
 sg13g2_dfrbp_1 _13623_ (.CLK(clknet_leaf_5_clk_regs),
    .RESET_B(net3421),
    .D(_00868_),
    .Q_N(_06162_),
    .Q(\u_toplayer.reg_layer1[159] ));
 sg13g2_dfrbp_1 _13624_ (.CLK(clknet_leaf_0_clk_regs),
    .RESET_B(net3407),
    .D(_00869_),
    .Q_N(_06161_),
    .Q(\u_toplayer.reg_layer1[160] ));
 sg13g2_dfrbp_1 _13625_ (.CLK(clknet_leaf_1_clk_regs),
    .RESET_B(net3405),
    .D(_00870_),
    .Q_N(_06160_),
    .Q(\u_toplayer.reg_layer1[161] ));
 sg13g2_dfrbp_1 _13626_ (.CLK(clknet_leaf_2_clk_regs),
    .RESET_B(net3411),
    .D(_00871_),
    .Q_N(_06159_),
    .Q(\u_toplayer.reg_layer1[162] ));
 sg13g2_dfrbp_1 _13627_ (.CLK(clknet_leaf_2_clk_regs),
    .RESET_B(net3411),
    .D(_00872_),
    .Q_N(_06158_),
    .Q(\u_toplayer.reg_layer1[163] ));
 sg13g2_dfrbp_1 _13628_ (.CLK(clknet_leaf_108_clk_regs),
    .RESET_B(net3413),
    .D(_00873_),
    .Q_N(_06157_),
    .Q(\u_toplayer.reg_layer1[164] ));
 sg13g2_dfrbp_1 _13629_ (.CLK(clknet_leaf_3_clk_regs),
    .RESET_B(net3413),
    .D(_00874_),
    .Q_N(_06156_),
    .Q(\u_toplayer.reg_layer1[165] ));
 sg13g2_dfrbp_1 _13630_ (.CLK(clknet_leaf_1_clk_regs),
    .RESET_B(net3406),
    .D(_00875_),
    .Q_N(_06155_),
    .Q(\u_toplayer.reg_layer1[166] ));
 sg13g2_dfrbp_1 _13631_ (.CLK(clknet_leaf_0_clk_regs),
    .RESET_B(net3405),
    .D(_00876_),
    .Q_N(_06154_),
    .Q(\u_toplayer.reg_layer1[167] ));
 sg13g2_dfrbp_1 _13632_ (.CLK(clknet_leaf_0_clk_regs),
    .RESET_B(net3407),
    .D(_00877_),
    .Q_N(_06153_),
    .Q(\u_toplayer.reg_layer1[168] ));
 sg13g2_dfrbp_1 _13633_ (.CLK(clknet_leaf_1_clk_regs),
    .RESET_B(net3407),
    .D(_00878_),
    .Q_N(_06152_),
    .Q(\u_toplayer.reg_layer1[169] ));
 sg13g2_dfrbp_1 _13634_ (.CLK(clknet_leaf_111_clk_regs),
    .RESET_B(net3410),
    .D(_00879_),
    .Q_N(_06151_),
    .Q(\u_toplayer.reg_layer1[170] ));
 sg13g2_dfrbp_1 _13635_ (.CLK(clknet_leaf_3_clk_regs),
    .RESET_B(net3411),
    .D(_00880_),
    .Q_N(_06150_),
    .Q(\u_toplayer.reg_layer1[171] ));
 sg13g2_dfrbp_1 _13636_ (.CLK(clknet_leaf_108_clk_regs),
    .RESET_B(net3409),
    .D(_00881_),
    .Q_N(_06149_),
    .Q(\u_toplayer.reg_layer1[172] ));
 sg13g2_dfrbp_1 _13637_ (.CLK(clknet_leaf_3_clk_regs),
    .RESET_B(net3413),
    .D(_00882_),
    .Q_N(_06148_),
    .Q(\u_toplayer.reg_layer1[173] ));
 sg13g2_dfrbp_1 _13638_ (.CLK(clknet_leaf_1_clk_regs),
    .RESET_B(net3405),
    .D(_00883_),
    .Q_N(_06147_),
    .Q(\u_toplayer.reg_layer1[174] ));
 sg13g2_dfrbp_1 _13639_ (.CLK(clknet_leaf_0_clk_regs),
    .RESET_B(net3405),
    .D(_00884_),
    .Q_N(_06146_),
    .Q(\u_toplayer.reg_layer1[175] ));
 sg13g2_dfrbp_1 _13640_ (.CLK(clknet_leaf_7_clk_regs),
    .RESET_B(net3407),
    .D(_00885_),
    .Q_N(_06145_),
    .Q(\u_toplayer.reg_layer1[176] ));
 sg13g2_dfrbp_1 _13641_ (.CLK(clknet_leaf_8_clk_regs),
    .RESET_B(net3415),
    .D(_00886_),
    .Q_N(_06144_),
    .Q(\u_toplayer.reg_layer1[177] ));
 sg13g2_dfrbp_1 _13642_ (.CLK(clknet_leaf_6_clk_regs),
    .RESET_B(net3412),
    .D(_00887_),
    .Q_N(_06143_),
    .Q(\u_toplayer.reg_layer1[178] ));
 sg13g2_dfrbp_1 _13643_ (.CLK(clknet_leaf_6_clk_regs),
    .RESET_B(net3411),
    .D(_00888_),
    .Q_N(_06142_),
    .Q(\u_toplayer.reg_layer1[179] ));
 sg13g2_dfrbp_1 _13644_ (.CLK(clknet_leaf_4_clk_regs),
    .RESET_B(net3413),
    .D(_00889_),
    .Q_N(_06141_),
    .Q(\u_toplayer.reg_layer1[180] ));
 sg13g2_dfrbp_1 _13645_ (.CLK(clknet_leaf_5_clk_regs),
    .RESET_B(net3419),
    .D(_00890_),
    .Q_N(_06140_),
    .Q(\u_toplayer.reg_layer1[181] ));
 sg13g2_dfrbp_1 _13646_ (.CLK(clknet_leaf_7_clk_regs),
    .RESET_B(net3415),
    .D(_00891_),
    .Q_N(_06139_),
    .Q(\u_toplayer.reg_layer1[182] ));
 sg13g2_dfrbp_1 _13647_ (.CLK(clknet_leaf_7_clk_regs),
    .RESET_B(net3415),
    .D(_00892_),
    .Q_N(_06138_),
    .Q(\u_toplayer.reg_layer1[183] ));
 sg13g2_dfrbp_1 _13648_ (.CLK(clknet_leaf_6_clk_regs),
    .RESET_B(net3406),
    .D(_00893_),
    .Q_N(_06137_),
    .Q(\u_toplayer.reg_layer1[184] ));
 sg13g2_dfrbp_1 _13649_ (.CLK(clknet_leaf_8_clk_regs),
    .RESET_B(net3415),
    .D(_00894_),
    .Q_N(_06136_),
    .Q(\u_toplayer.reg_layer1[185] ));
 sg13g2_dfrbp_1 _13650_ (.CLK(clknet_leaf_6_clk_regs),
    .RESET_B(net3412),
    .D(_00895_),
    .Q_N(_06135_),
    .Q(\u_toplayer.reg_layer1[186] ));
 sg13g2_dfrbp_1 _13651_ (.CLK(clknet_leaf_2_clk_regs),
    .RESET_B(net3412),
    .D(_00896_),
    .Q_N(_06134_),
    .Q(\u_toplayer.reg_layer1[187] ));
 sg13g2_dfrbp_1 _13652_ (.CLK(clknet_leaf_4_clk_regs),
    .RESET_B(net3414),
    .D(_00897_),
    .Q_N(_06133_),
    .Q(\u_toplayer.reg_layer1[188] ));
 sg13g2_dfrbp_1 _13653_ (.CLK(clknet_leaf_4_clk_regs),
    .RESET_B(net3419),
    .D(_00898_),
    .Q_N(_06132_),
    .Q(\u_toplayer.reg_layer1[189] ));
 sg13g2_dfrbp_1 _13654_ (.CLK(clknet_leaf_7_clk_regs),
    .RESET_B(net3406),
    .D(_00899_),
    .Q_N(_06131_),
    .Q(\u_toplayer.reg_layer1[190] ));
 sg13g2_dfrbp_1 _13655_ (.CLK(clknet_leaf_8_clk_regs),
    .RESET_B(net3417),
    .D(_00900_),
    .Q_N(_06130_),
    .Q(\u_toplayer.reg_layer1[191] ));
 sg13g2_dfrbp_1 _13656_ (.CLK(clknet_leaf_96_clk_regs),
    .RESET_B(net3440),
    .D(_00901_),
    .Q_N(_06129_),
    .Q(\u_toplayer.reg_layer1[192] ));
 sg13g2_dfrbp_1 _13657_ (.CLK(clknet_leaf_99_clk_regs),
    .RESET_B(net3493),
    .D(_00902_),
    .Q_N(_06128_),
    .Q(\u_toplayer.reg_layer1[193] ));
 sg13g2_dfrbp_1 _13658_ (.CLK(clknet_leaf_98_clk_regs),
    .RESET_B(net3441),
    .D(_00903_),
    .Q_N(_06127_),
    .Q(\u_toplayer.reg_layer1[194] ));
 sg13g2_dfrbp_1 _13659_ (.CLK(clknet_leaf_99_clk_regs),
    .RESET_B(net3493),
    .D(_00904_),
    .Q_N(_06126_),
    .Q(\u_toplayer.reg_layer1[195] ));
 sg13g2_dfrbp_1 _13660_ (.CLK(clknet_leaf_99_clk_regs),
    .RESET_B(net3441),
    .D(_00905_),
    .Q_N(_06125_),
    .Q(\u_toplayer.reg_layer1[196] ));
 sg13g2_dfrbp_1 _13661_ (.CLK(clknet_leaf_97_clk_regs),
    .RESET_B(net3440),
    .D(_00906_),
    .Q_N(_06124_),
    .Q(\u_toplayer.reg_layer1[197] ));
 sg13g2_dfrbp_1 _13662_ (.CLK(clknet_leaf_97_clk_regs),
    .RESET_B(net3441),
    .D(_00907_),
    .Q_N(_06123_),
    .Q(\u_toplayer.reg_layer1[198] ));
 sg13g2_dfrbp_1 _13663_ (.CLK(clknet_leaf_98_clk_regs),
    .RESET_B(net3494),
    .D(net293),
    .Q_N(_06122_),
    .Q(\u_toplayer.reg_layer1[199] ));
 sg13g2_dfrbp_1 _13664_ (.CLK(clknet_leaf_97_clk_regs),
    .RESET_B(net3440),
    .D(net491),
    .Q_N(_06121_),
    .Q(\u_toplayer.reg_layer1[200] ));
 sg13g2_dfrbp_1 _13665_ (.CLK(clknet_leaf_100_clk_regs),
    .RESET_B(net3489),
    .D(net780),
    .Q_N(_06120_),
    .Q(\u_toplayer.reg_layer1[201] ));
 sg13g2_dfrbp_1 _13666_ (.CLK(clknet_leaf_80_clk_regs),
    .RESET_B(net3489),
    .D(_00911_),
    .Q_N(_06119_),
    .Q(\u_toplayer.reg_layer1[202] ));
 sg13g2_dfrbp_1 _13667_ (.CLK(clknet_leaf_80_clk_regs),
    .RESET_B(net3489),
    .D(_00912_),
    .Q_N(_06118_),
    .Q(\u_toplayer.reg_layer1[203] ));
 sg13g2_dfrbp_1 _13668_ (.CLK(clknet_leaf_100_clk_regs),
    .RESET_B(net3438),
    .D(_00913_),
    .Q_N(_06117_),
    .Q(\u_toplayer.reg_layer1[204] ));
 sg13g2_dfrbp_1 _13669_ (.CLK(clknet_leaf_99_clk_regs),
    .RESET_B(net3441),
    .D(net737),
    .Q_N(_06116_),
    .Q(\u_toplayer.reg_layer1[205] ));
 sg13g2_dfrbp_1 _13670_ (.CLK(clknet_leaf_100_clk_regs),
    .RESET_B(net3438),
    .D(_00915_),
    .Q_N(_06115_),
    .Q(\u_toplayer.reg_layer1[206] ));
 sg13g2_dfrbp_1 _13671_ (.CLK(clknet_leaf_80_clk_regs),
    .RESET_B(net3493),
    .D(net695),
    .Q_N(_06114_),
    .Q(\u_toplayer.reg_layer1[207] ));
 sg13g2_dfrbp_1 _13672_ (.CLK(clknet_leaf_95_clk_regs),
    .RESET_B(net3446),
    .D(_00917_),
    .Q_N(_06113_),
    .Q(\u_toplayer.reg_layer1[208] ));
 sg13g2_dfrbp_1 _13673_ (.CLK(clknet_leaf_94_clk_regs),
    .RESET_B(net3452),
    .D(_00918_),
    .Q_N(_06112_),
    .Q(\u_toplayer.reg_layer1[209] ));
 sg13g2_dfrbp_1 _13674_ (.CLK(clknet_leaf_92_clk_regs),
    .RESET_B(net3455),
    .D(_00919_),
    .Q_N(_06111_),
    .Q(\u_toplayer.reg_layer1[210] ));
 sg13g2_dfrbp_1 _13675_ (.CLK(clknet_leaf_98_clk_regs),
    .RESET_B(net3506),
    .D(_00920_),
    .Q_N(_06110_),
    .Q(\u_toplayer.reg_layer1[211] ));
 sg13g2_dfrbp_1 _13676_ (.CLK(clknet_leaf_96_clk_regs),
    .RESET_B(net3433),
    .D(_00921_),
    .Q_N(_06109_),
    .Q(\u_toplayer.reg_layer1[212] ));
 sg13g2_dfrbp_1 _13677_ (.CLK(clknet_leaf_94_clk_regs),
    .RESET_B(net3451),
    .D(_00922_),
    .Q_N(_06108_),
    .Q(\u_toplayer.reg_layer1[213] ));
 sg13g2_dfrbp_1 _13678_ (.CLK(clknet_leaf_95_clk_regs),
    .RESET_B(net3446),
    .D(_00923_),
    .Q_N(_06107_),
    .Q(\u_toplayer.reg_layer1[214] ));
 sg13g2_dfrbp_1 _13679_ (.CLK(clknet_leaf_98_clk_regs),
    .RESET_B(net3506),
    .D(net447),
    .Q_N(_06106_),
    .Q(\u_toplayer.reg_layer1[215] ));
 sg13g2_dfrbp_1 _13680_ (.CLK(clknet_leaf_93_clk_regs),
    .RESET_B(net3450),
    .D(_00925_),
    .Q_N(_06105_),
    .Q(\u_toplayer.reg_layer1[216] ));
 sg13g2_dfrbp_1 _13681_ (.CLK(clknet_leaf_98_clk_regs),
    .RESET_B(net3441),
    .D(_00926_),
    .Q_N(_06104_),
    .Q(\u_toplayer.reg_layer1[217] ));
 sg13g2_dfrbp_1 _13682_ (.CLK(clknet_leaf_92_clk_regs),
    .RESET_B(net3452),
    .D(_00927_),
    .Q_N(_06103_),
    .Q(\u_toplayer.reg_layer1[218] ));
 sg13g2_dfrbp_1 _13683_ (.CLK(clknet_leaf_98_clk_regs),
    .RESET_B(net3494),
    .D(_00928_),
    .Q_N(_06102_),
    .Q(\u_toplayer.reg_layer1[219] ));
 sg13g2_dfrbp_1 _13684_ (.CLK(clknet_leaf_96_clk_regs),
    .RESET_B(net3442),
    .D(net680),
    .Q_N(_06101_),
    .Q(\u_toplayer.reg_layer1[220] ));
 sg13g2_dfrbp_1 _13685_ (.CLK(clknet_leaf_97_clk_regs),
    .RESET_B(net3450),
    .D(_00930_),
    .Q_N(_06100_),
    .Q(\u_toplayer.reg_layer1[221] ));
 sg13g2_dfrbp_1 _13686_ (.CLK(clknet_leaf_96_clk_regs),
    .RESET_B(net3450),
    .D(_00931_),
    .Q_N(_06099_),
    .Q(\u_toplayer.reg_layer1[222] ));
 sg13g2_dfrbp_1 _13687_ (.CLK(clknet_leaf_93_clk_regs),
    .RESET_B(net3506),
    .D(net854),
    .Q_N(_06098_),
    .Q(\u_toplayer.reg_layer1[223] ));
 sg13g2_dfrbp_1 _13688_ (.CLK(clknet_leaf_106_clk_regs),
    .RESET_B(net3430),
    .D(net306),
    .Q_N(_06097_),
    .Q(\u_toplayer.reg_layer1[224] ));
 sg13g2_dfrbp_1 _13689_ (.CLK(clknet_leaf_103_clk_regs),
    .RESET_B(net3436),
    .D(_00934_),
    .Q_N(_06096_),
    .Q(\u_toplayer.reg_layer1[225] ));
 sg13g2_dfrbp_1 _13690_ (.CLK(clknet_leaf_103_clk_regs),
    .RESET_B(net3436),
    .D(_00935_),
    .Q_N(_06095_),
    .Q(\u_toplayer.reg_layer1[226] ));
 sg13g2_dfrbp_1 _13691_ (.CLK(clknet_leaf_102_clk_regs),
    .RESET_B(net3435),
    .D(_00936_),
    .Q_N(_06094_),
    .Q(\u_toplayer.reg_layer1[227] ));
 sg13g2_dfrbp_1 _13692_ (.CLK(clknet_leaf_104_clk_regs),
    .RESET_B(net3429),
    .D(_00937_),
    .Q_N(_06093_),
    .Q(\u_toplayer.reg_layer1[228] ));
 sg13g2_dfrbp_1 _13693_ (.CLK(clknet_leaf_103_clk_regs),
    .RESET_B(net3435),
    .D(_00938_),
    .Q_N(_06092_),
    .Q(\u_toplayer.reg_layer1[229] ));
 sg13g2_dfrbp_1 _13694_ (.CLK(clknet_leaf_106_clk_regs),
    .RESET_B(net3432),
    .D(net322),
    .Q_N(_06091_),
    .Q(\u_toplayer.reg_layer1[230] ));
 sg13g2_dfrbp_1 _13695_ (.CLK(clknet_leaf_106_clk_regs),
    .RESET_B(net3430),
    .D(net327),
    .Q_N(_06090_),
    .Q(\u_toplayer.reg_layer1[231] ));
 sg13g2_dfrbp_1 _13696_ (.CLK(clknet_leaf_103_clk_regs),
    .RESET_B(net3436),
    .D(_00941_),
    .Q_N(_06089_),
    .Q(\u_toplayer.reg_layer1[232] ));
 sg13g2_dfrbp_1 _13697_ (.CLK(clknet_leaf_100_clk_regs),
    .RESET_B(net3437),
    .D(_00942_),
    .Q_N(_06088_),
    .Q(\u_toplayer.reg_layer1[233] ));
 sg13g2_dfrbp_1 _13698_ (.CLK(clknet_leaf_101_clk_regs),
    .RESET_B(net3437),
    .D(net422),
    .Q_N(_06087_),
    .Q(\u_toplayer.reg_layer1[234] ));
 sg13g2_dfrbp_1 _13699_ (.CLK(clknet_leaf_102_clk_regs),
    .RESET_B(net3437),
    .D(net469),
    .Q_N(_06086_),
    .Q(\u_toplayer.reg_layer1[235] ));
 sg13g2_dfrbp_1 _13700_ (.CLK(clknet_leaf_102_clk_regs),
    .RESET_B(net3435),
    .D(net493),
    .Q_N(_06085_),
    .Q(\u_toplayer.reg_layer1[236] ));
 sg13g2_dfrbp_1 _13701_ (.CLK(clknet_leaf_101_clk_regs),
    .RESET_B(net3437),
    .D(_00946_),
    .Q_N(_06084_),
    .Q(\u_toplayer.reg_layer1[237] ));
 sg13g2_dfrbp_1 _13702_ (.CLK(clknet_leaf_106_clk_regs),
    .RESET_B(net3440),
    .D(net568),
    .Q_N(_06083_),
    .Q(\u_toplayer.reg_layer1[238] ));
 sg13g2_dfrbp_1 _13703_ (.CLK(clknet_leaf_102_clk_regs),
    .RESET_B(net3435),
    .D(net371),
    .Q_N(_06082_),
    .Q(\u_toplayer.reg_layer1[239] ));
 sg13g2_dfrbp_1 _13704_ (.CLK(clknet_leaf_107_clk_regs),
    .RESET_B(net3433),
    .D(_00949_),
    .Q_N(_06081_),
    .Q(\u_toplayer.reg_layer1[240] ));
 sg13g2_dfrbp_1 _13705_ (.CLK(clknet_leaf_107_clk_regs),
    .RESET_B(net3432),
    .D(net477),
    .Q_N(_06080_),
    .Q(\u_toplayer.reg_layer1[241] ));
 sg13g2_dfrbp_1 _13706_ (.CLK(clknet_leaf_105_clk_regs),
    .RESET_B(net3428),
    .D(net725),
    .Q_N(_06079_),
    .Q(\u_toplayer.reg_layer1[242] ));
 sg13g2_dfrbp_1 _13707_ (.CLK(clknet_leaf_105_clk_regs),
    .RESET_B(net3429),
    .D(net402),
    .Q_N(_06078_),
    .Q(\u_toplayer.reg_layer1[243] ));
 sg13g2_dfrbp_1 _13708_ (.CLK(clknet_leaf_105_clk_regs),
    .RESET_B(net3430),
    .D(net577),
    .Q_N(_06077_),
    .Q(\u_toplayer.reg_layer1[244] ));
 sg13g2_dfrbp_1 _13709_ (.CLK(clknet_leaf_109_clk_regs),
    .RESET_B(net3428),
    .D(net501),
    .Q_N(_06076_),
    .Q(\u_toplayer.reg_layer1[245] ));
 sg13g2_dfrbp_1 _13710_ (.CLK(clknet_leaf_107_clk_regs),
    .RESET_B(net3434),
    .D(_00955_),
    .Q_N(_06075_),
    .Q(\u_toplayer.reg_layer1[246] ));
 sg13g2_dfrbp_1 _13711_ (.CLK(clknet_leaf_109_clk_regs),
    .RESET_B(net3434),
    .D(net793),
    .Q_N(_06074_),
    .Q(\u_toplayer.reg_layer1[247] ));
 sg13g2_dfrbp_1 _13712_ (.CLK(clknet_leaf_106_clk_regs),
    .RESET_B(net3432),
    .D(_00957_),
    .Q_N(_06073_),
    .Q(\u_toplayer.reg_layer1[248] ));
 sg13g2_dfrbp_1 _13713_ (.CLK(clknet_leaf_107_clk_regs),
    .RESET_B(net3432),
    .D(net414),
    .Q_N(_06072_),
    .Q(\u_toplayer.reg_layer1[249] ));
 sg13g2_dfrbp_1 _13714_ (.CLK(clknet_leaf_110_clk_regs),
    .RESET_B(net3431),
    .D(_00959_),
    .Q_N(_06071_),
    .Q(\u_toplayer.reg_layer1[250] ));
 sg13g2_dfrbp_1 _13715_ (.CLK(clknet_leaf_104_clk_regs),
    .RESET_B(net3429),
    .D(_00960_),
    .Q_N(_06070_),
    .Q(\u_toplayer.reg_layer1[251] ));
 sg13g2_dfrbp_1 _13716_ (.CLK(clknet_leaf_105_clk_regs),
    .RESET_B(net3430),
    .D(_00961_),
    .Q_N(_06069_),
    .Q(\u_toplayer.reg_layer1[252] ));
 sg13g2_dfrbp_1 _13717_ (.CLK(clknet_leaf_110_clk_regs),
    .RESET_B(net3428),
    .D(_00962_),
    .Q_N(_06068_),
    .Q(\u_toplayer.reg_layer1[253] ));
 sg13g2_dfrbp_1 _13718_ (.CLK(clknet_leaf_108_clk_regs),
    .RESET_B(net3434),
    .D(_00963_),
    .Q_N(_06067_),
    .Q(\u_toplayer.reg_layer1[254] ));
 sg13g2_dfrbp_1 _13719_ (.CLK(clknet_leaf_109_clk_regs),
    .RESET_B(net3428),
    .D(_00964_),
    .Q_N(_06066_),
    .Q(\u_toplayer.reg_layer1[255] ));
 sg13g2_dfrbp_1 _13720_ (.CLK(clknet_leaf_38_clk_regs),
    .RESET_B(net3557),
    .D(_00965_),
    .Q_N(_06065_),
    .Q(\u_toplayer.u_layer1.u_neuron.b[0] ));
 sg13g2_dfrbp_1 _13721_ (.CLK(clknet_leaf_38_clk_regs),
    .RESET_B(net3557),
    .D(_00966_),
    .Q_N(_06064_),
    .Q(\u_toplayer.u_layer1.u_neuron.b[1] ));
 sg13g2_dfrbp_1 _13722_ (.CLK(clknet_leaf_41_clk_regs),
    .RESET_B(net3555),
    .D(_00967_),
    .Q_N(_06063_),
    .Q(\u_toplayer.u_layer1.u_neuron.b[2] ));
 sg13g2_dfrbp_1 _13723_ (.CLK(clknet_leaf_42_clk_regs),
    .RESET_B(net3557),
    .D(_00968_),
    .Q_N(_06062_),
    .Q(\u_toplayer.u_layer1.u_neuron.b[3] ));
 sg13g2_dfrbp_1 _13724_ (.CLK(clknet_leaf_40_clk_regs),
    .RESET_B(net3555),
    .D(_00969_),
    .Q_N(_06061_),
    .Q(\u_toplayer.u_layer1.u_neuron.b[4] ));
 sg13g2_dfrbp_1 _13725_ (.CLK(clknet_leaf_41_clk_regs),
    .RESET_B(net3554),
    .D(_00970_),
    .Q_N(_06060_),
    .Q(\u_toplayer.u_layer1.u_neuron.b[5] ));
 sg13g2_dfrbp_1 _13726_ (.CLK(clknet_leaf_42_clk_regs),
    .RESET_B(net3557),
    .D(_00971_),
    .Q_N(_06059_),
    .Q(\u_toplayer.u_layer1.u_neuron.b[6] ));
 sg13g2_dfrbp_1 _13727_ (.CLK(clknet_leaf_44_clk_regs),
    .RESET_B(net3556),
    .D(_00972_),
    .Q_N(_06058_),
    .Q(\u_toplayer.u_layer1.u_neuron.b[7] ));
 sg13g2_dfrbp_1 _13728_ (.CLK(clknet_leaf_95_clk_regs),
    .RESET_B(net3451),
    .D(_00973_),
    .Q_N(_06057_),
    .Q(\u_toplayer.u_layer1.sum[0] ));
 sg13g2_dfrbp_1 _13729_ (.CLK(clknet_leaf_16_clk_regs),
    .RESET_B(net3453),
    .D(_00974_),
    .Q_N(_06056_),
    .Q(\u_toplayer.u_layer1.sum[1] ));
 sg13g2_dfrbp_1 _13730_ (.CLK(clknet_leaf_94_clk_regs),
    .RESET_B(net3451),
    .D(_00975_),
    .Q_N(_06055_),
    .Q(\u_toplayer.u_layer1.sum[2] ));
 sg13g2_dfrbp_1 _13731_ (.CLK(clknet_leaf_14_clk_regs),
    .RESET_B(net3453),
    .D(_00976_),
    .Q_N(_06054_),
    .Q(\u_toplayer.u_layer1.sum[3] ));
 sg13g2_dfrbp_1 _13732_ (.CLK(clknet_leaf_94_clk_regs),
    .RESET_B(net3452),
    .D(_00977_),
    .Q_N(_06053_),
    .Q(\u_toplayer.u_layer1.sum[4] ));
 sg13g2_dfrbp_1 _13733_ (.CLK(clknet_leaf_94_clk_regs),
    .RESET_B(net3451),
    .D(_00978_),
    .Q_N(_06052_),
    .Q(\u_toplayer.u_layer1.sum[5] ));
 sg13g2_dfrbp_1 _13734_ (.CLK(clknet_leaf_16_clk_regs),
    .RESET_B(net3453),
    .D(_00979_),
    .Q_N(_06051_),
    .Q(\u_toplayer.u_layer1.sum[6] ));
 sg13g2_dfrbp_1 _13735_ (.CLK(clknet_leaf_36_clk_regs),
    .RESET_B(net3553),
    .D(net971),
    .Q_N(_06050_),
    .Q(\u_toplayer.u_layer1.sum[7] ));
 sg13g2_dfrbp_1 _13736_ (.CLK(clknet_leaf_110_clk_regs),
    .RESET_B(net3408),
    .D(_00981_),
    .Q_N(_06049_),
    .Q(\u_toplayer.u_layer1.statel1[0] ));
 sg13g2_dfrbp_1 _13737_ (.CLK(clknet_leaf_110_clk_regs),
    .RESET_B(net3408),
    .D(net922),
    .Q_N(_06048_),
    .Q(\u_toplayer.u_layer1.statel1[1] ));
 sg13g2_dfrbp_1 _13738_ (.CLK(clknet_leaf_111_clk_regs),
    .RESET_B(net3408),
    .D(_00983_),
    .Q_N(_06047_),
    .Q(\u_toplayer.u_layer1.statel1[2] ));
 sg13g2_dfrbp_1 _13739_ (.CLK(clknet_leaf_111_clk_regs),
    .RESET_B(net3410),
    .D(net961),
    .Q_N(_06046_),
    .Q(\u_toplayer.u_layer1.statel1[3] ));
 sg13g2_dfrbp_1 _13740_ (.CLK(clknet_leaf_111_clk_regs),
    .RESET_B(net3410),
    .D(_00985_),
    .Q_N(_06045_),
    .Q(\u_toplayer.u_layer1.statel1[4] ));
 sg13g2_dfrbp_1 _13741_ (.CLK(clknet_leaf_111_clk_regs),
    .RESET_B(net3408),
    .D(net878),
    .Q_N(_06044_),
    .Q(\u_toplayer.u_layer1.statel1[5] ));
 sg13g2_dfrbp_1 _13742_ (.CLK(clknet_leaf_111_clk_regs),
    .RESET_B(net3408),
    .D(net1016),
    .Q_N(_06043_),
    .Q(\u_toplayer.u_layer1.statel1[6] ));
 sg13g2_dfrbp_1 _13743_ (.CLK(clknet_leaf_110_clk_regs),
    .RESET_B(net3408),
    .D(net973),
    .Q_N(_06042_),
    .Q(\u_toplayer.u_layer1.statel1[7] ));
 sg13g2_dfrbp_1 _13744_ (.CLK(clknet_leaf_111_clk_regs),
    .RESET_B(net3408),
    .D(net626),
    .Q_N(_00029_),
    .Q(\u_toplayer.u_layer1.statel1[8] ));
 sg13g2_dfrbp_1 _13745_ (.CLK(clknet_leaf_39_clk_regs),
    .RESET_B(net3557),
    .D(_00990_),
    .Q_N(_06041_),
    .Q(\u_toplayer.u_layer1.u_neuron.acc[0] ));
 sg13g2_dfrbp_1 _13746_ (.CLK(clknet_leaf_38_clk_regs),
    .RESET_B(net3557),
    .D(_00991_),
    .Q_N(_06040_),
    .Q(\u_toplayer.u_layer1.u_neuron.acc[1] ));
 sg13g2_dfrbp_1 _13747_ (.CLK(clknet_leaf_37_clk_regs),
    .RESET_B(net3554),
    .D(_00992_),
    .Q_N(_06039_),
    .Q(\u_toplayer.u_layer1.u_neuron.acc[2] ));
 sg13g2_dfrbp_1 _13748_ (.CLK(clknet_leaf_37_clk_regs),
    .RESET_B(net3554),
    .D(_00993_),
    .Q_N(_06038_),
    .Q(\u_toplayer.u_layer1.u_neuron.acc[3] ));
 sg13g2_dfrbp_1 _13749_ (.CLK(clknet_leaf_37_clk_regs),
    .RESET_B(net3554),
    .D(_00994_),
    .Q_N(_06037_),
    .Q(\u_toplayer.u_layer1.u_neuron.acc[4] ));
 sg13g2_dfrbp_1 _13750_ (.CLK(clknet_leaf_39_clk_regs),
    .RESET_B(net3554),
    .D(_00995_),
    .Q_N(_06036_),
    .Q(\u_toplayer.u_layer1.u_neuron.acc[5] ));
 sg13g2_dfrbp_1 _13751_ (.CLK(clknet_leaf_39_clk_regs),
    .RESET_B(net3555),
    .D(_00996_),
    .Q_N(_06035_),
    .Q(\u_toplayer.u_layer1.u_neuron.acc[6] ));
 sg13g2_dfrbp_1 _13752_ (.CLK(clknet_leaf_39_clk_regs),
    .RESET_B(net3557),
    .D(_00997_),
    .Q_N(_06034_),
    .Q(\u_toplayer.u_layer1.u_neuron.acc[7] ));
 sg13g2_dfrbp_1 _13753_ (.CLK(clknet_leaf_44_clk_regs),
    .RESET_B(net3558),
    .D(_00998_),
    .Q_N(_06033_),
    .Q(\u_toplayer.u_layer1.u_neuron.acc[8] ));
 sg13g2_dfrbp_1 _13754_ (.CLK(clknet_leaf_39_clk_regs),
    .RESET_B(net3558),
    .D(_00999_),
    .Q_N(_06032_),
    .Q(\u_toplayer.u_layer1.u_neuron.acc[9] ));
 sg13g2_dfrbp_1 _13755_ (.CLK(clknet_leaf_43_clk_regs),
    .RESET_B(net3559),
    .D(_01000_),
    .Q_N(_06031_),
    .Q(\u_toplayer.u_layer1.u_neuron.acc[10] ));
 sg13g2_dfrbp_1 _13756_ (.CLK(clknet_leaf_43_clk_regs),
    .RESET_B(net3559),
    .D(_01001_),
    .Q_N(_06030_),
    .Q(\u_toplayer.u_layer1.u_neuron.acc[11] ));
 sg13g2_dfrbp_1 _13757_ (.CLK(clknet_leaf_43_clk_regs),
    .RESET_B(net3560),
    .D(_01002_),
    .Q_N(_06029_),
    .Q(\u_toplayer.u_layer1.u_neuron.acc[12] ));
 sg13g2_dfrbp_1 _13758_ (.CLK(clknet_leaf_43_clk_regs),
    .RESET_B(net3556),
    .D(_01003_),
    .Q_N(_06028_),
    .Q(\u_toplayer.u_layer1.u_neuron.acc[13] ));
 sg13g2_dfrbp_1 _13759_ (.CLK(clknet_leaf_43_clk_regs),
    .RESET_B(net3559),
    .D(_01004_),
    .Q_N(_06027_),
    .Q(\u_toplayer.u_layer1.u_neuron.acc[14] ));
 sg13g2_dfrbp_1 _13760_ (.CLK(clknet_leaf_44_clk_regs),
    .RESET_B(net3559),
    .D(_01005_),
    .Q_N(_06026_),
    .Q(\u_toplayer.u_layer1.u_neuron.acc[15] ));
 sg13g2_dfrbp_1 _13761_ (.CLK(clknet_leaf_44_clk_regs),
    .RESET_B(net3562),
    .D(_01006_),
    .Q_N(_06025_),
    .Q(\u_toplayer.u_layer1.u_neuron.acc[16] ));
 sg13g2_dfrbp_1 _13762_ (.CLK(clknet_leaf_44_clk_regs),
    .RESET_B(net3562),
    .D(_01007_),
    .Q_N(_06024_),
    .Q(\u_toplayer.u_layer1.u_neuron.acc[17] ));
 sg13g2_dfrbp_1 _13763_ (.CLK(clknet_leaf_44_clk_regs),
    .RESET_B(net3561),
    .D(_01008_),
    .Q_N(_06023_),
    .Q(\u_toplayer.u_layer1.u_neuron.acc[18] ));
 sg13g2_dfrbp_1 _13764_ (.CLK(clknet_leaf_44_clk_regs),
    .RESET_B(net3562),
    .D(_01009_),
    .Q_N(_06022_),
    .Q(\u_toplayer.u_layer1.u_neuron.acc[19] ));
 sg13g2_dfrbp_1 _13765_ (.CLK(clknet_leaf_45_clk_regs),
    .RESET_B(net3561),
    .D(_01010_),
    .Q_N(_06021_),
    .Q(\u_toplayer.u_layer1.u_neuron.acc[20] ));
 sg13g2_dfrbp_1 _13766_ (.CLK(clknet_leaf_45_clk_regs),
    .RESET_B(net3561),
    .D(_01011_),
    .Q_N(_06020_),
    .Q(\u_toplayer.u_layer1.u_neuron.acc[21] ));
 sg13g2_dfrbp_1 _13767_ (.CLK(clknet_leaf_45_clk_regs),
    .RESET_B(net3562),
    .D(_01012_),
    .Q_N(_06019_),
    .Q(\u_toplayer.u_layer1.u_neuron.acc[22] ));
 sg13g2_dfrbp_1 _13768_ (.CLK(clknet_leaf_39_clk_regs),
    .RESET_B(net3558),
    .D(_01013_),
    .Q_N(_06018_),
    .Q(\u_toplayer.u_layer1.u_neuron.acc[23] ));
 sg13g2_dfrbp_1 _13769_ (.CLK(clknet_leaf_101_clk_regs),
    .RESET_B(net3488),
    .D(net125),
    .Q_N(_06017_),
    .Q(\u_toplayer.delay_counter_layer1[0] ));
 sg13g2_dfrbp_1 _13770_ (.CLK(clknet_leaf_101_clk_regs),
    .RESET_B(net3488),
    .D(_01015_),
    .Q_N(_06885_),
    .Q(\u_toplayer.delay_counter_layer1[1] ));
 sg13g2_dfrbp_1 _13771_ (.CLK(clknet_leaf_20_clk_regs),
    .RESET_B(net3417),
    .D(_00011_),
    .Q_N(_06886_),
    .Q(\u_toplayer.delayed_done_layer3 ));
 sg13g2_dfrbp_1 _13772_ (.CLK(clknet_leaf_91_clk_regs),
    .RESET_B(net3508),
    .D(_00009_),
    .Q_N(_06887_),
    .Q(\u_toplayer.delayed_done_layer2 ));
 sg13g2_dfrbp_1 _13773_ (.CLK(clknet_leaf_79_clk_regs),
    .RESET_B(net3488),
    .D(_00010_),
    .Q_N(_06016_),
    .Q(\u_toplayer.delayed_done_layer1 ));
 sg13g2_dfrbp_1 _13774_ (.CLK(clknet_leaf_80_clk_regs),
    .RESET_B(net3488),
    .D(net131),
    .Q_N(_06015_),
    .Q(\u_toplayer.delay_counter_layer2[0] ));
 sg13g2_dfrbp_1 _13775_ (.CLK(clknet_leaf_100_clk_regs),
    .RESET_B(net3488),
    .D(net926),
    .Q_N(_06014_),
    .Q(\u_toplayer.delay_counter_layer2[1] ));
 sg13g2_tielo tt_um_neural_navigators_5 (.L_LO(net5));
 sg13g2_tielo tt_um_neural_navigators_6 (.L_LO(net6));
 sg13g2_tielo tt_um_neural_navigators_7 (.L_LO(net7));
 sg13g2_tielo tt_um_neural_navigators_8 (.L_LO(net8));
 sg13g2_tielo tt_um_neural_navigators_9 (.L_LO(net9));
 sg13g2_tielo tt_um_neural_navigators_10 (.L_LO(net10));
 sg13g2_tielo tt_um_neural_navigators_11 (.L_LO(net11));
 sg13g2_tielo tt_um_neural_navigators_12 (.L_LO(net12));
 sg13g2_tielo tt_um_neural_navigators_13 (.L_LO(net13));
 sg13g2_tielo tt_um_neural_navigators_14 (.L_LO(net14));
 sg13g2_tielo tt_um_neural_navigators_15 (.L_LO(net15));
 sg13g2_tielo tt_um_neural_navigators_16 (.L_LO(net16));
 sg13g2_tielo tt_um_neural_navigators_17 (.L_LO(net17));
 sg13g2_tielo tt_um_neural_navigators_18 (.L_LO(net18));
 sg13g2_tielo tt_um_neural_navigators_19 (.L_LO(net19));
 sg13g2_inv_1 _07055__1 (.Y(net20),
    .A(clknet_4_9_0_clk));
 sg13g2_buf_2 fanout2692 (.A(net2693),
    .X(net2692));
 sg13g2_buf_4 fanout2693 (.X(net2693),
    .A(net2701));
 sg13g2_buf_4 fanout2694 (.X(net2694),
    .A(net2696));
 sg13g2_buf_2 fanout2695 (.A(net2696),
    .X(net2695));
 sg13g2_buf_2 fanout2696 (.A(net2700),
    .X(net2696));
 sg13g2_buf_4 fanout2697 (.X(net2697),
    .A(net2699));
 sg13g2_buf_2 fanout2698 (.A(net2699),
    .X(net2698));
 sg13g2_buf_2 fanout2699 (.A(net2700),
    .X(net2699));
 sg13g2_buf_2 fanout2700 (.A(net2701),
    .X(net2700));
 sg13g2_buf_2 fanout2701 (.A(_04539_),
    .X(net2701));
 sg13g2_buf_2 fanout2702 (.A(net2704),
    .X(net2702));
 sg13g2_buf_1 fanout2703 (.A(net2704),
    .X(net2703));
 sg13g2_buf_2 fanout2704 (.A(_04392_),
    .X(net2704));
 sg13g2_buf_2 fanout2705 (.A(_04392_),
    .X(net2705));
 sg13g2_buf_2 fanout2706 (.A(net2711),
    .X(net2706));
 sg13g2_buf_4 fanout2707 (.X(net2707),
    .A(net2711));
 sg13g2_buf_4 fanout2708 (.X(net2708),
    .A(net2710));
 sg13g2_buf_2 fanout2709 (.A(net2710),
    .X(net2709));
 sg13g2_buf_4 fanout2710 (.X(net2710),
    .A(net2711));
 sg13g2_buf_2 fanout2711 (.A(_04392_),
    .X(net2711));
 sg13g2_buf_4 fanout2712 (.X(net2712),
    .A(_04464_));
 sg13g2_buf_4 fanout2713 (.X(net2713),
    .A(_04464_));
 sg13g2_buf_4 fanout2714 (.X(net2714),
    .A(net2715));
 sg13g2_buf_4 fanout2715 (.X(net2715),
    .A(_04175_));
 sg13g2_buf_4 fanout2716 (.X(net2716),
    .A(_04174_));
 sg13g2_buf_2 fanout2717 (.A(net2719),
    .X(net2717));
 sg13g2_buf_4 fanout2718 (.X(net2718),
    .A(net2719));
 sg13g2_buf_2 fanout2719 (.A(net2721),
    .X(net2719));
 sg13g2_buf_2 fanout2720 (.A(net2721),
    .X(net2720));
 sg13g2_buf_2 fanout2721 (.A(_05471_),
    .X(net2721));
 sg13g2_buf_2 fanout2722 (.A(net2724),
    .X(net2722));
 sg13g2_buf_2 fanout2723 (.A(net2724),
    .X(net2723));
 sg13g2_buf_2 fanout2724 (.A(net2726),
    .X(net2724));
 sg13g2_buf_2 fanout2725 (.A(net2726),
    .X(net2725));
 sg13g2_buf_2 fanout2726 (.A(_05471_),
    .X(net2726));
 sg13g2_buf_2 fanout2727 (.A(_02653_),
    .X(net2727));
 sg13g2_buf_2 fanout2728 (.A(_01945_),
    .X(net2728));
 sg13g2_buf_2 fanout2729 (.A(_01945_),
    .X(net2729));
 sg13g2_buf_2 fanout2730 (.A(_01943_),
    .X(net2730));
 sg13g2_buf_2 fanout2731 (.A(_01943_),
    .X(net2731));
 sg13g2_buf_2 fanout2732 (.A(net2735),
    .X(net2732));
 sg13g2_buf_1 fanout2733 (.A(net2735),
    .X(net2733));
 sg13g2_buf_4 fanout2734 (.X(net2734),
    .A(net2735));
 sg13g2_buf_2 fanout2735 (.A(net2736),
    .X(net2735));
 sg13g2_buf_2 fanout2736 (.A(_05624_),
    .X(net2736));
 sg13g2_buf_2 fanout2737 (.A(net2738),
    .X(net2737));
 sg13g2_buf_2 fanout2738 (.A(net2740),
    .X(net2738));
 sg13g2_buf_4 fanout2739 (.X(net2739),
    .A(net2740));
 sg13g2_buf_2 fanout2740 (.A(_05624_),
    .X(net2740));
 sg13g2_buf_4 fanout2741 (.X(net2741),
    .A(_05256_));
 sg13g2_buf_2 fanout2742 (.A(net2743),
    .X(net2742));
 sg13g2_buf_1 fanout2743 (.A(net2744),
    .X(net2743));
 sg13g2_buf_2 fanout2744 (.A(_05246_),
    .X(net2744));
 sg13g2_buf_2 fanout2745 (.A(net2746),
    .X(net2745));
 sg13g2_buf_1 fanout2746 (.A(net2747),
    .X(net2746));
 sg13g2_buf_2 fanout2747 (.A(_03756_),
    .X(net2747));
 sg13g2_buf_2 fanout2748 (.A(_02650_),
    .X(net2748));
 sg13g2_buf_2 fanout2749 (.A(_02650_),
    .X(net2749));
 sg13g2_buf_2 fanout2750 (.A(net2751),
    .X(net2750));
 sg13g2_buf_2 fanout2751 (.A(net2756),
    .X(net2751));
 sg13g2_buf_2 fanout2752 (.A(net2753),
    .X(net2752));
 sg13g2_buf_2 fanout2753 (.A(net2756),
    .X(net2753));
 sg13g2_buf_2 fanout2754 (.A(net2756),
    .X(net2754));
 sg13g2_buf_2 fanout2755 (.A(net2756),
    .X(net2755));
 sg13g2_buf_2 fanout2756 (.A(_02649_),
    .X(net2756));
 sg13g2_buf_2 fanout2757 (.A(net2759),
    .X(net2757));
 sg13g2_buf_2 fanout2758 (.A(net2759),
    .X(net2758));
 sg13g2_buf_4 fanout2759 (.X(net2759),
    .A(_01942_));
 sg13g2_buf_2 fanout2760 (.A(net2761),
    .X(net2760));
 sg13g2_buf_2 fanout2761 (.A(net2764),
    .X(net2761));
 sg13g2_buf_2 fanout2762 (.A(net2764),
    .X(net2762));
 sg13g2_buf_1 fanout2763 (.A(net2764),
    .X(net2763));
 sg13g2_buf_2 fanout2764 (.A(_01941_),
    .X(net2764));
 sg13g2_buf_2 fanout2765 (.A(_01256_),
    .X(net2765));
 sg13g2_buf_4 fanout2766 (.X(net2766),
    .A(_01254_));
 sg13g2_buf_2 fanout2767 (.A(_01252_),
    .X(net2767));
 sg13g2_buf_4 fanout2768 (.X(net2768),
    .A(_01250_));
 sg13g2_buf_2 fanout2769 (.A(net2770),
    .X(net2769));
 sg13g2_buf_4 fanout2770 (.X(net2770),
    .A(net2773));
 sg13g2_buf_1 fanout2771 (.A(net2773),
    .X(net2771));
 sg13g2_buf_4 fanout2772 (.X(net2772),
    .A(net2773));
 sg13g2_buf_2 fanout2773 (.A(net2777),
    .X(net2773));
 sg13g2_buf_2 fanout2774 (.A(net2777),
    .X(net2774));
 sg13g2_buf_2 fanout2775 (.A(net2776),
    .X(net2775));
 sg13g2_buf_2 fanout2776 (.A(net2777),
    .X(net2776));
 sg13g2_buf_2 fanout2777 (.A(net2780),
    .X(net2777));
 sg13g2_buf_4 fanout2778 (.X(net2778),
    .A(net2779));
 sg13g2_buf_4 fanout2779 (.X(net2779),
    .A(net2780));
 sg13g2_buf_2 fanout2780 (.A(_05255_),
    .X(net2780));
 sg13g2_buf_2 fanout2781 (.A(net2782),
    .X(net2781));
 sg13g2_buf_2 fanout2782 (.A(net2785),
    .X(net2782));
 sg13g2_buf_1 fanout2783 (.A(net2785),
    .X(net2783));
 sg13g2_buf_4 fanout2784 (.X(net2784),
    .A(net2785));
 sg13g2_buf_2 fanout2785 (.A(net2789),
    .X(net2785));
 sg13g2_buf_4 fanout2786 (.X(net2786),
    .A(net2789));
 sg13g2_buf_2 fanout2787 (.A(net2788),
    .X(net2787));
 sg13g2_buf_4 fanout2788 (.X(net2788),
    .A(net2789));
 sg13g2_buf_2 fanout2789 (.A(net2792),
    .X(net2789));
 sg13g2_buf_4 fanout2790 (.X(net2790),
    .A(net2791));
 sg13g2_buf_4 fanout2791 (.X(net2791),
    .A(net2792));
 sg13g2_buf_2 fanout2792 (.A(_05245_),
    .X(net2792));
 sg13g2_buf_4 fanout2793 (.X(net2793),
    .A(net2795));
 sg13g2_buf_2 fanout2794 (.A(net2795),
    .X(net2794));
 sg13g2_buf_4 fanout2795 (.X(net2795),
    .A(net2796));
 sg13g2_buf_2 fanout2796 (.A(_04182_),
    .X(net2796));
 sg13g2_buf_4 fanout2797 (.X(net2797),
    .A(net2801));
 sg13g2_buf_2 fanout2798 (.A(net2800),
    .X(net2798));
 sg13g2_buf_1 fanout2799 (.A(net2800),
    .X(net2799));
 sg13g2_buf_2 fanout2800 (.A(net2801),
    .X(net2800));
 sg13g2_buf_2 fanout2801 (.A(net2802),
    .X(net2801));
 sg13g2_buf_4 fanout2802 (.X(net2802),
    .A(_04182_));
 sg13g2_buf_2 fanout2803 (.A(net2806),
    .X(net2803));
 sg13g2_buf_2 fanout2804 (.A(net2806),
    .X(net2804));
 sg13g2_buf_4 fanout2805 (.X(net2805),
    .A(net2806));
 sg13g2_buf_2 fanout2806 (.A(net2807),
    .X(net2806));
 sg13g2_buf_2 fanout2807 (.A(net2813),
    .X(net2807));
 sg13g2_buf_4 fanout2808 (.X(net2808),
    .A(net2812));
 sg13g2_buf_1 fanout2809 (.A(net2812),
    .X(net2809));
 sg13g2_buf_4 fanout2810 (.X(net2810),
    .A(net2811));
 sg13g2_buf_2 fanout2811 (.A(net2812),
    .X(net2811));
 sg13g2_buf_4 fanout2812 (.X(net2812),
    .A(net2813));
 sg13g2_buf_4 fanout2813 (.X(net2813),
    .A(_04168_));
 sg13g2_buf_2 fanout2814 (.A(net2815),
    .X(net2814));
 sg13g2_buf_2 fanout2815 (.A(_03754_),
    .X(net2815));
 sg13g2_buf_2 fanout2816 (.A(_03375_),
    .X(net2816));
 sg13g2_buf_4 fanout2817 (.X(net2817),
    .A(_01938_));
 sg13g2_buf_2 fanout2818 (.A(_05233_),
    .X(net2818));
 sg13g2_buf_2 fanout2819 (.A(_04907_),
    .X(net2819));
 sg13g2_buf_2 fanout2820 (.A(net2823),
    .X(net2820));
 sg13g2_buf_1 fanout2821 (.A(net2823),
    .X(net2821));
 sg13g2_buf_2 fanout2822 (.A(net2823),
    .X(net2822));
 sg13g2_buf_2 fanout2823 (.A(net2824),
    .X(net2823));
 sg13g2_buf_2 fanout2824 (.A(_04179_),
    .X(net2824));
 sg13g2_buf_4 fanout2825 (.X(net2825),
    .A(net2828));
 sg13g2_buf_2 fanout2826 (.A(net2827),
    .X(net2826));
 sg13g2_buf_2 fanout2827 (.A(net2828),
    .X(net2827));
 sg13g2_buf_2 fanout2828 (.A(net2829),
    .X(net2828));
 sg13g2_buf_2 fanout2829 (.A(_04179_),
    .X(net2829));
 sg13g2_buf_2 fanout2830 (.A(net2831),
    .X(net2830));
 sg13g2_buf_2 fanout2831 (.A(net2832),
    .X(net2831));
 sg13g2_buf_2 fanout2832 (.A(net2837),
    .X(net2832));
 sg13g2_buf_2 fanout2833 (.A(net2834),
    .X(net2833));
 sg13g2_buf_2 fanout2834 (.A(net2837),
    .X(net2834));
 sg13g2_buf_2 fanout2835 (.A(net2837),
    .X(net2835));
 sg13g2_buf_2 fanout2836 (.A(net2837),
    .X(net2836));
 sg13g2_buf_2 fanout2837 (.A(_03750_),
    .X(net2837));
 sg13g2_buf_4 fanout2838 (.X(net2838),
    .A(_01219_));
 sg13g2_buf_4 fanout2839 (.X(net2839),
    .A(net2841));
 sg13g2_buf_4 fanout2840 (.X(net2840),
    .A(net2841));
 sg13g2_buf_2 fanout2841 (.A(_01215_),
    .X(net2841));
 sg13g2_buf_4 fanout2842 (.X(net2842),
    .A(_05687_));
 sg13g2_buf_2 fanout2843 (.A(net2844),
    .X(net2843));
 sg13g2_buf_2 fanout2844 (.A(net2847),
    .X(net2844));
 sg13g2_buf_2 fanout2845 (.A(net2846),
    .X(net2845));
 sg13g2_buf_2 fanout2846 (.A(net2847),
    .X(net2846));
 sg13g2_buf_1 fanout2847 (.A(net2850),
    .X(net2847));
 sg13g2_buf_2 fanout2848 (.A(net2849),
    .X(net2848));
 sg13g2_buf_2 fanout2849 (.A(net2850),
    .X(net2849));
 sg13g2_buf_2 fanout2850 (.A(_05262_),
    .X(net2850));
 sg13g2_buf_4 fanout2851 (.X(net2851),
    .A(_05262_));
 sg13g2_buf_2 fanout2852 (.A(_05262_),
    .X(net2852));
 sg13g2_buf_4 fanout2853 (.X(net2853),
    .A(_03752_));
 sg13g2_buf_2 fanout2854 (.A(_03752_),
    .X(net2854));
 sg13g2_buf_4 fanout2855 (.X(net2855),
    .A(_03751_));
 sg13g2_buf_2 fanout2856 (.A(_03751_),
    .X(net2856));
 sg13g2_buf_4 fanout2857 (.X(net2857),
    .A(_03746_));
 sg13g2_buf_4 fanout2858 (.X(net2858),
    .A(_02644_));
 sg13g2_buf_2 fanout2859 (.A(_02644_),
    .X(net2859));
 sg13g2_buf_2 fanout2860 (.A(net2861),
    .X(net2860));
 sg13g2_buf_4 fanout2861 (.X(net2861),
    .A(_02643_));
 sg13g2_buf_4 fanout2862 (.X(net2862),
    .A(_01936_));
 sg13g2_buf_1 fanout2863 (.A(_01936_),
    .X(net2863));
 sg13g2_buf_2 fanout2864 (.A(net2865),
    .X(net2864));
 sg13g2_buf_4 fanout2865 (.X(net2865),
    .A(_01935_));
 sg13g2_buf_4 fanout2866 (.X(net2866),
    .A(_01217_));
 sg13g2_buf_4 fanout2867 (.X(net2867),
    .A(_01216_));
 sg13g2_buf_2 fanout2868 (.A(net2871),
    .X(net2868));
 sg13g2_buf_2 fanout2869 (.A(net2870),
    .X(net2869));
 sg13g2_buf_2 fanout2870 (.A(net2871),
    .X(net2870));
 sg13g2_buf_2 fanout2871 (.A(_05243_),
    .X(net2871));
 sg13g2_buf_2 fanout2872 (.A(net2873),
    .X(net2872));
 sg13g2_buf_2 fanout2873 (.A(net2874),
    .X(net2873));
 sg13g2_buf_2 fanout2874 (.A(_05243_),
    .X(net2874));
 sg13g2_buf_2 fanout2875 (.A(net2877),
    .X(net2875));
 sg13g2_buf_2 fanout2876 (.A(net2877),
    .X(net2876));
 sg13g2_buf_2 fanout2877 (.A(_04204_),
    .X(net2877));
 sg13g2_buf_2 fanout2878 (.A(net2880),
    .X(net2878));
 sg13g2_buf_2 fanout2879 (.A(net2880),
    .X(net2879));
 sg13g2_buf_2 fanout2880 (.A(_04163_),
    .X(net2880));
 sg13g2_buf_2 fanout2881 (.A(net2883),
    .X(net2881));
 sg13g2_buf_1 fanout2882 (.A(net2883),
    .X(net2882));
 sg13g2_buf_2 fanout2883 (.A(_04163_),
    .X(net2883));
 sg13g2_buf_2 fanout2884 (.A(_02639_),
    .X(net2884));
 sg13g2_buf_1 fanout2885 (.A(_02639_),
    .X(net2885));
 sg13g2_buf_2 fanout2886 (.A(net2887),
    .X(net2886));
 sg13g2_buf_2 fanout2887 (.A(_02638_),
    .X(net2887));
 sg13g2_buf_2 fanout2888 (.A(net2890),
    .X(net2888));
 sg13g2_buf_2 fanout2889 (.A(net2890),
    .X(net2889));
 sg13g2_buf_2 fanout2890 (.A(_02343_),
    .X(net2890));
 sg13g2_buf_2 fanout2891 (.A(_02343_),
    .X(net2891));
 sg13g2_buf_2 fanout2892 (.A(net2893),
    .X(net2892));
 sg13g2_buf_2 fanout2893 (.A(_02342_),
    .X(net2893));
 sg13g2_buf_4 fanout2894 (.X(net2894),
    .A(_01931_));
 sg13g2_buf_2 fanout2895 (.A(_01931_),
    .X(net2895));
 sg13g2_buf_4 fanout2896 (.X(net2896),
    .A(_01930_));
 sg13g2_buf_2 fanout2897 (.A(_01930_),
    .X(net2897));
 sg13g2_buf_4 fanout2898 (.X(net2898),
    .A(_05392_));
 sg13g2_buf_2 fanout2899 (.A(_05392_),
    .X(net2899));
 sg13g2_buf_2 fanout2900 (.A(net2902),
    .X(net2900));
 sg13g2_buf_2 fanout2901 (.A(net2902),
    .X(net2901));
 sg13g2_buf_2 fanout2902 (.A(_05365_),
    .X(net2902));
 sg13g2_buf_2 fanout2903 (.A(net2905),
    .X(net2903));
 sg13g2_buf_4 fanout2904 (.X(net2904),
    .A(net2905));
 sg13g2_buf_2 fanout2905 (.A(_05339_),
    .X(net2905));
 sg13g2_buf_4 fanout2906 (.X(net2906),
    .A(_05311_));
 sg13g2_buf_4 fanout2907 (.X(net2907),
    .A(_05311_));
 sg13g2_buf_2 fanout2908 (.A(net2910),
    .X(net2908));
 sg13g2_buf_4 fanout2909 (.X(net2909),
    .A(net2910));
 sg13g2_buf_2 fanout2910 (.A(_05287_),
    .X(net2910));
 sg13g2_buf_4 fanout2911 (.X(net2911),
    .A(net2913));
 sg13g2_buf_4 fanout2912 (.X(net2912),
    .A(net2913));
 sg13g2_buf_4 fanout2913 (.X(net2913),
    .A(_05257_));
 sg13g2_buf_2 fanout2914 (.A(net2915),
    .X(net2914));
 sg13g2_buf_2 fanout2915 (.A(_04615_),
    .X(net2915));
 sg13g2_buf_2 fanout2916 (.A(net2918),
    .X(net2916));
 sg13g2_buf_4 fanout2917 (.X(net2917),
    .A(net2918));
 sg13g2_buf_4 fanout2918 (.X(net2918),
    .A(_04285_));
 sg13g2_buf_2 fanout2919 (.A(net2921),
    .X(net2919));
 sg13g2_buf_4 fanout2920 (.X(net2920),
    .A(net2921));
 sg13g2_buf_2 fanout2921 (.A(_04258_),
    .X(net2921));
 sg13g2_buf_2 fanout2922 (.A(_04231_),
    .X(net2922));
 sg13g2_buf_2 fanout2923 (.A(_04231_),
    .X(net2923));
 sg13g2_buf_2 fanout2924 (.A(_04170_),
    .X(net2924));
 sg13g2_buf_2 fanout2925 (.A(_04170_),
    .X(net2925));
 sg13g2_buf_4 fanout2926 (.X(net2926),
    .A(net2928));
 sg13g2_buf_4 fanout2927 (.X(net2927),
    .A(net2928));
 sg13g2_buf_2 fanout2928 (.A(_03738_),
    .X(net2928));
 sg13g2_buf_2 fanout2929 (.A(net2930),
    .X(net2929));
 sg13g2_buf_2 fanout2930 (.A(_03734_),
    .X(net2930));
 sg13g2_buf_4 fanout2931 (.X(net2931),
    .A(_03734_));
 sg13g2_buf_4 fanout2932 (.X(net2932),
    .A(_02346_));
 sg13g2_buf_4 fanout2933 (.X(net2933),
    .A(_02345_));
 sg13g2_buf_2 fanout2934 (.A(_02345_),
    .X(net2934));
 sg13g2_buf_2 fanout2935 (.A(net2937),
    .X(net2935));
 sg13g2_buf_1 fanout2936 (.A(net2937),
    .X(net2936));
 sg13g2_buf_2 fanout2937 (.A(_01939_),
    .X(net2937));
 sg13g2_buf_2 fanout2938 (.A(_01898_),
    .X(net2938));
 sg13g2_buf_2 fanout2939 (.A(_01803_),
    .X(net2939));
 sg13g2_buf_2 fanout2940 (.A(net2941),
    .X(net2940));
 sg13g2_buf_2 fanout2941 (.A(_01392_),
    .X(net2941));
 sg13g2_buf_2 fanout2942 (.A(net2944),
    .X(net2942));
 sg13g2_buf_2 fanout2943 (.A(net2944),
    .X(net2943));
 sg13g2_buf_4 fanout2944 (.X(net2944),
    .A(_01391_));
 sg13g2_buf_4 fanout2945 (.X(net2945),
    .A(_05237_));
 sg13g2_buf_4 fanout2946 (.X(net2946),
    .A(net2947));
 sg13g2_buf_2 fanout2947 (.A(_05237_),
    .X(net2947));
 sg13g2_buf_2 fanout2948 (.A(net2949),
    .X(net2948));
 sg13g2_buf_2 fanout2949 (.A(_04164_),
    .X(net2949));
 sg13g2_buf_4 fanout2950 (.X(net2950),
    .A(_04164_));
 sg13g2_buf_4 fanout2951 (.X(net2951),
    .A(_02877_));
 sg13g2_buf_2 fanout2952 (.A(_02780_),
    .X(net2952));
 sg13g2_buf_1 fanout2953 (.A(_02780_),
    .X(net2953));
 sg13g2_buf_4 fanout2954 (.X(net2954),
    .A(net2955));
 sg13g2_buf_4 fanout2955 (.X(net2955),
    .A(net2956));
 sg13g2_buf_2 fanout2956 (.A(_02642_),
    .X(net2956));
 sg13g2_buf_4 fanout2957 (.X(net2957),
    .A(net2958));
 sg13g2_buf_2 fanout2958 (.A(net2959),
    .X(net2958));
 sg13g2_buf_4 fanout2959 (.X(net2959),
    .A(_02642_));
 sg13g2_buf_4 fanout2960 (.X(net2960),
    .A(net2961));
 sg13g2_buf_2 fanout2961 (.A(net2962),
    .X(net2961));
 sg13g2_buf_2 fanout2962 (.A(net2964),
    .X(net2962));
 sg13g2_buf_4 fanout2963 (.X(net2963),
    .A(net2964));
 sg13g2_buf_2 fanout2964 (.A(_02642_),
    .X(net2964));
 sg13g2_buf_4 fanout2965 (.X(net2965),
    .A(net2966));
 sg13g2_buf_4 fanout2966 (.X(net2966),
    .A(net2967));
 sg13g2_buf_4 fanout2967 (.X(net2967),
    .A(net2970));
 sg13g2_buf_4 fanout2968 (.X(net2968),
    .A(net2969));
 sg13g2_buf_4 fanout2969 (.X(net2969),
    .A(net2970));
 sg13g2_buf_2 fanout2970 (.A(_01934_),
    .X(net2970));
 sg13g2_buf_4 fanout2971 (.X(net2971),
    .A(net2972));
 sg13g2_buf_4 fanout2972 (.X(net2972),
    .A(net2974));
 sg13g2_buf_4 fanout2973 (.X(net2973),
    .A(net2974));
 sg13g2_buf_2 fanout2974 (.A(_01934_),
    .X(net2974));
 sg13g2_buf_2 fanout2975 (.A(_01572_),
    .X(net2975));
 sg13g2_buf_4 fanout2976 (.X(net2976),
    .A(net2978));
 sg13g2_buf_4 fanout2977 (.X(net2977),
    .A(net2978));
 sg13g2_buf_4 fanout2978 (.X(net2978),
    .A(_01390_));
 sg13g2_buf_4 fanout2979 (.X(net2979),
    .A(_01389_));
 sg13g2_buf_4 fanout2980 (.X(net2980),
    .A(net2981));
 sg13g2_buf_2 fanout2981 (.A(net2983),
    .X(net2981));
 sg13g2_buf_2 fanout2982 (.A(net2983),
    .X(net2982));
 sg13g2_buf_2 fanout2983 (.A(_01385_),
    .X(net2983));
 sg13g2_buf_2 fanout2984 (.A(net2986),
    .X(net2984));
 sg13g2_buf_2 fanout2985 (.A(net2986),
    .X(net2985));
 sg13g2_buf_2 fanout2986 (.A(net2995),
    .X(net2986));
 sg13g2_buf_4 fanout2987 (.X(net2987),
    .A(net2989));
 sg13g2_buf_2 fanout2988 (.A(net2989),
    .X(net2988));
 sg13g2_buf_2 fanout2989 (.A(net2995),
    .X(net2989));
 sg13g2_buf_2 fanout2990 (.A(net2994),
    .X(net2990));
 sg13g2_buf_2 fanout2991 (.A(net2994),
    .X(net2991));
 sg13g2_buf_2 fanout2992 (.A(net2994),
    .X(net2992));
 sg13g2_buf_1 fanout2993 (.A(net2994),
    .X(net2993));
 sg13g2_buf_2 fanout2994 (.A(net2995),
    .X(net2994));
 sg13g2_buf_2 fanout2995 (.A(_01352_),
    .X(net2995));
 sg13g2_buf_2 fanout2996 (.A(net2997),
    .X(net2996));
 sg13g2_buf_2 fanout2997 (.A(_01349_),
    .X(net2997));
 sg13g2_buf_2 fanout2998 (.A(net2999),
    .X(net2998));
 sg13g2_buf_2 fanout2999 (.A(net3000),
    .X(net2999));
 sg13g2_buf_4 fanout3000 (.X(net3000),
    .A(net3003));
 sg13g2_buf_2 fanout3001 (.A(net3002),
    .X(net3001));
 sg13g2_buf_2 fanout3002 (.A(net3003),
    .X(net3002));
 sg13g2_buf_2 fanout3003 (.A(net3007),
    .X(net3003));
 sg13g2_buf_2 fanout3004 (.A(net3005),
    .X(net3004));
 sg13g2_buf_2 fanout3005 (.A(net3006),
    .X(net3005));
 sg13g2_buf_2 fanout3006 (.A(net3007),
    .X(net3006));
 sg13g2_buf_2 fanout3007 (.A(_01335_),
    .X(net3007));
 sg13g2_buf_2 fanout3008 (.A(net3010),
    .X(net3008));
 sg13g2_buf_1 fanout3009 (.A(net3010),
    .X(net3009));
 sg13g2_buf_2 fanout3010 (.A(_01333_),
    .X(net3010));
 sg13g2_buf_4 fanout3011 (.X(net3011),
    .A(net3013));
 sg13g2_buf_4 fanout3012 (.X(net3012),
    .A(net3013));
 sg13g2_buf_2 fanout3013 (.A(_01324_),
    .X(net3013));
 sg13g2_buf_2 fanout3014 (.A(net3016),
    .X(net3014));
 sg13g2_buf_2 fanout3015 (.A(net3016),
    .X(net3015));
 sg13g2_buf_2 fanout3016 (.A(_01321_),
    .X(net3016));
 sg13g2_buf_2 fanout3017 (.A(net3018),
    .X(net3017));
 sg13g2_buf_2 fanout3018 (.A(_01036_),
    .X(net3018));
 sg13g2_buf_4 fanout3019 (.X(net3019),
    .A(_01035_));
 sg13g2_buf_2 fanout3020 (.A(_01035_),
    .X(net3020));
 sg13g2_buf_4 fanout3021 (.X(net3021),
    .A(_01029_));
 sg13g2_buf_2 fanout3022 (.A(_01029_),
    .X(net3022));
 sg13g2_buf_2 fanout3023 (.A(_01029_),
    .X(net3023));
 sg13g2_buf_2 fanout3024 (.A(net1193),
    .X(net3024));
 sg13g2_buf_2 fanout3025 (.A(net1204),
    .X(net3025));
 sg13g2_buf_2 fanout3026 (.A(\u_toplayer.u_layer1.u_neuron.acc[16] ),
    .X(net3026));
 sg13g2_buf_2 fanout3027 (.A(net1198),
    .X(net3027));
 sg13g2_buf_2 fanout3028 (.A(net1165),
    .X(net3028));
 sg13g2_buf_4 fanout3029 (.X(net3029),
    .A(net1145));
 sg13g2_buf_2 fanout3030 (.A(net1192),
    .X(net3030));
 sg13g2_buf_4 fanout3031 (.X(net3031),
    .A(net3032));
 sg13g2_buf_2 fanout3032 (.A(net3033),
    .X(net3032));
 sg13g2_buf_8 fanout3033 (.A(\u_toplayer.u_layer1.sum[7] ),
    .X(net3033));
 sg13g2_buf_4 fanout3034 (.X(net3034),
    .A(net3035));
 sg13g2_buf_4 fanout3035 (.X(net3035),
    .A(\u_toplayer.u_layer1.sum[6] ));
 sg13g2_buf_4 fanout3036 (.X(net3036),
    .A(net3037));
 sg13g2_buf_4 fanout3037 (.X(net3037),
    .A(\u_toplayer.u_layer1.sum[5] ));
 sg13g2_buf_4 fanout3038 (.X(net3038),
    .A(net3039));
 sg13g2_buf_4 fanout3039 (.X(net3039),
    .A(\u_toplayer.u_layer1.sum[4] ));
 sg13g2_buf_4 fanout3040 (.X(net3040),
    .A(\u_toplayer.u_layer1.sum[3] ));
 sg13g2_buf_4 fanout3041 (.X(net3041),
    .A(\u_toplayer.u_layer1.sum[3] ));
 sg13g2_buf_4 fanout3042 (.X(net3042),
    .A(net3043));
 sg13g2_buf_4 fanout3043 (.X(net3043),
    .A(\u_toplayer.u_layer1.sum[2] ));
 sg13g2_buf_4 fanout3044 (.X(net3044),
    .A(net3045));
 sg13g2_buf_4 fanout3045 (.X(net3045),
    .A(\u_toplayer.u_layer1.sum[1] ));
 sg13g2_buf_4 fanout3046 (.X(net3046),
    .A(net3047));
 sg13g2_buf_4 fanout3047 (.X(net3047),
    .A(\u_toplayer.u_layer1.sum[0] ));
 sg13g2_buf_2 fanout3048 (.A(net3049),
    .X(net3048));
 sg13g2_buf_2 fanout3049 (.A(\u_toplayer.u_layer1.u_neuron.b[7] ),
    .X(net3049));
 sg13g2_buf_4 fanout3050 (.X(net3050),
    .A(net1188));
 sg13g2_buf_2 fanout3051 (.A(net3052),
    .X(net3051));
 sg13g2_buf_2 fanout3052 (.A(\u_toplayer.u_layer1.u_neuron.b[7] ),
    .X(net3052));
 sg13g2_buf_2 fanout3053 (.A(net1043),
    .X(net3053));
 sg13g2_buf_4 fanout3054 (.X(net3054),
    .A(\u_toplayer.u_layer1.neuron_index[3] ));
 sg13g2_buf_2 fanout3055 (.A(net3056),
    .X(net3055));
 sg13g2_buf_4 fanout3056 (.X(net3056),
    .A(\u_toplayer.u_layer1.neuron_index[2] ));
 sg13g2_buf_2 fanout3057 (.A(\u_toplayer.u_layer1.neuron_index[0] ),
    .X(net3057));
 sg13g2_buf_2 fanout3058 (.A(net1203),
    .X(net3058));
 sg13g2_buf_2 fanout3059 (.A(net1194),
    .X(net3059));
 sg13g2_buf_2 fanout3060 (.A(net1189),
    .X(net3060));
 sg13g2_buf_2 fanout3061 (.A(net1195),
    .X(net3061));
 sg13g2_buf_2 fanout3062 (.A(net1182),
    .X(net3062));
 sg13g2_buf_2 fanout3063 (.A(net821),
    .X(net3063));
 sg13g2_buf_2 fanout3064 (.A(net785),
    .X(net3064));
 sg13g2_buf_4 fanout3065 (.X(net3065),
    .A(net3066));
 sg13g2_buf_4 fanout3066 (.X(net3066),
    .A(\u_toplayer.u_layer2.sum[7] ));
 sg13g2_buf_4 fanout3067 (.X(net3067),
    .A(net3068));
 sg13g2_buf_4 fanout3068 (.X(net3068),
    .A(\u_toplayer.u_layer2.sum[6] ));
 sg13g2_buf_4 fanout3069 (.X(net3069),
    .A(net3070));
 sg13g2_buf_4 fanout3070 (.X(net3070),
    .A(\u_toplayer.u_layer2.sum[5] ));
 sg13g2_buf_4 fanout3071 (.X(net3071),
    .A(net3073));
 sg13g2_buf_4 fanout3072 (.X(net3072),
    .A(net3073));
 sg13g2_buf_4 fanout3073 (.X(net3073),
    .A(\u_toplayer.u_layer2.sum[4] ));
 sg13g2_buf_4 fanout3074 (.X(net3074),
    .A(net3075));
 sg13g2_buf_4 fanout3075 (.X(net3075),
    .A(\u_toplayer.u_layer2.sum[3] ));
 sg13g2_buf_4 fanout3076 (.X(net3076),
    .A(net3077));
 sg13g2_buf_4 fanout3077 (.X(net3077),
    .A(\u_toplayer.u_layer2.sum[2] ));
 sg13g2_buf_4 fanout3078 (.X(net3078),
    .A(\u_toplayer.u_layer2.sum[1] ));
 sg13g2_buf_4 fanout3079 (.X(net3079),
    .A(net1205));
 sg13g2_buf_4 fanout3080 (.X(net3080),
    .A(net3081));
 sg13g2_buf_4 fanout3081 (.X(net3081),
    .A(\u_toplayer.u_layer2.sum[0] ));
 sg13g2_buf_4 fanout3082 (.X(net3082),
    .A(net3083));
 sg13g2_buf_4 fanout3083 (.X(net3083),
    .A(\u_toplayer.u_layer2.u_neuron.din[7] ));
 sg13g2_buf_2 fanout3084 (.A(net1207),
    .X(net3084));
 sg13g2_buf_4 fanout3085 (.X(net3085),
    .A(net1197));
 sg13g2_buf_4 fanout3086 (.X(net3086),
    .A(net1160));
 sg13g2_buf_2 fanout3087 (.A(\u_toplayer.u_layer2.u_neuron.din[4] ),
    .X(net3087));
 sg13g2_buf_2 fanout3088 (.A(net1187),
    .X(net3088));
 sg13g2_buf_2 fanout3089 (.A(\u_toplayer.u_layer2.u_neuron.din[3] ),
    .X(net3089));
 sg13g2_buf_4 fanout3090 (.X(net3090),
    .A(net1141));
 sg13g2_buf_2 fanout3091 (.A(\u_toplayer.u_layer2.u_neuron.din[2] ),
    .X(net3091));
 sg13g2_buf_4 fanout3092 (.X(net3092),
    .A(net1152));
 sg13g2_buf_2 fanout3093 (.A(\u_toplayer.u_layer2.u_neuron.din[1] ),
    .X(net3093));
 sg13g2_buf_4 fanout3094 (.X(net3094),
    .A(net1186));
 sg13g2_buf_2 fanout3095 (.A(\u_toplayer.u_layer2.u_neuron.din[0] ),
    .X(net3095));
 sg13g2_buf_2 fanout3096 (.A(net3098),
    .X(net3096));
 sg13g2_buf_2 fanout3097 (.A(net3098),
    .X(net3097));
 sg13g2_buf_4 fanout3098 (.X(net3098),
    .A(\u_toplayer.u_layer3.u_neuron.instCtrl.state[4] ));
 sg13g2_buf_2 fanout3099 (.A(net3101),
    .X(net3099));
 sg13g2_buf_2 fanout3100 (.A(net3101),
    .X(net3100));
 sg13g2_buf_2 fanout3101 (.A(\u_toplayer.u_layer3.u_neuron.instCtrl.state[3] ),
    .X(net3101));
 sg13g2_buf_4 fanout3102 (.X(net3102),
    .A(net3105));
 sg13g2_buf_2 fanout3103 (.A(net3105),
    .X(net3103));
 sg13g2_buf_1 fanout3104 (.A(net3105),
    .X(net3104));
 sg13g2_buf_2 fanout3105 (.A(\u_toplayer.u_layer3.u_neuron.instCtrl.state[2] ),
    .X(net3105));
 sg13g2_buf_2 fanout3106 (.A(net3107),
    .X(net3106));
 sg13g2_buf_4 fanout3107 (.X(net3107),
    .A(net3110));
 sg13g2_buf_4 fanout3108 (.X(net3108),
    .A(net3109));
 sg13g2_buf_4 fanout3109 (.X(net3109),
    .A(net3110));
 sg13g2_buf_2 fanout3110 (.A(net3116),
    .X(net3110));
 sg13g2_buf_2 fanout3111 (.A(net3112),
    .X(net3111));
 sg13g2_buf_4 fanout3112 (.X(net3112),
    .A(net3116));
 sg13g2_buf_2 fanout3113 (.A(net3114),
    .X(net3113));
 sg13g2_buf_2 fanout3114 (.A(net3115),
    .X(net3114));
 sg13g2_buf_4 fanout3115 (.X(net3115),
    .A(net3116));
 sg13g2_buf_2 fanout3116 (.A(\u_toplayer.u_layer3.u_neuron.instCtrl.state[1] ),
    .X(net3116));
 sg13g2_buf_2 fanout3117 (.A(net3120),
    .X(net3117));
 sg13g2_buf_2 fanout3118 (.A(net3119),
    .X(net3118));
 sg13g2_buf_2 fanout3119 (.A(net3120),
    .X(net3119));
 sg13g2_buf_2 fanout3120 (.A(net3128),
    .X(net3120));
 sg13g2_buf_2 fanout3121 (.A(net3122),
    .X(net3121));
 sg13g2_buf_2 fanout3122 (.A(net3128),
    .X(net3122));
 sg13g2_buf_2 fanout3123 (.A(net3128),
    .X(net3123));
 sg13g2_buf_1 fanout3124 (.A(net3127),
    .X(net3124));
 sg13g2_buf_2 fanout3125 (.A(net3126),
    .X(net3125));
 sg13g2_buf_1 fanout3126 (.A(net3127),
    .X(net3126));
 sg13g2_buf_4 fanout3127 (.X(net3127),
    .A(net3128));
 sg13g2_buf_2 fanout3128 (.A(\u_toplayer.u_layer3.u_neuron.instCtrl.state[0] ),
    .X(net3128));
 sg13g2_buf_2 fanout3129 (.A(net3131),
    .X(net3129));
 sg13g2_buf_2 fanout3130 (.A(net3131),
    .X(net3130));
 sg13g2_buf_1 fanout3131 (.A(net3135),
    .X(net3131));
 sg13g2_buf_2 fanout3132 (.A(net3134),
    .X(net3132));
 sg13g2_buf_1 fanout3133 (.A(net3134),
    .X(net3133));
 sg13g2_buf_4 fanout3134 (.X(net3134),
    .A(net3135));
 sg13g2_buf_1 fanout3135 (.A(\u_toplayer.u_layer3.u_neuron.instCtrl.state[0] ),
    .X(net3135));
 sg13g2_buf_2 fanout3136 (.A(net3137),
    .X(net3136));
 sg13g2_buf_2 fanout3137 (.A(net3141),
    .X(net3137));
 sg13g2_buf_2 fanout3138 (.A(net3140),
    .X(net3138));
 sg13g2_buf_1 fanout3139 (.A(net3140),
    .X(net3139));
 sg13g2_buf_2 fanout3140 (.A(net3141),
    .X(net3140));
 sg13g2_buf_1 fanout3141 (.A(\u_toplayer.u_layer3.u_neuron.instCtrl.state[0] ),
    .X(net3141));
 sg13g2_buf_2 fanout3142 (.A(net3144),
    .X(net3142));
 sg13g2_buf_2 fanout3143 (.A(net3144),
    .X(net3143));
 sg13g2_buf_2 fanout3144 (.A(net1209),
    .X(net3144));
 sg13g2_buf_4 fanout3145 (.X(net3145),
    .A(net3146));
 sg13g2_buf_2 fanout3146 (.A(\u_toplayer.u_layer2.neuron_index[3] ),
    .X(net3146));
 sg13g2_buf_2 fanout3147 (.A(net3148),
    .X(net3147));
 sg13g2_buf_2 fanout3148 (.A(\u_toplayer.u_layer2.neuron_index[3] ),
    .X(net3148));
 sg13g2_buf_4 fanout3149 (.X(net3149),
    .A(net3150));
 sg13g2_buf_2 fanout3150 (.A(\u_toplayer.u_layer2.neuron_index[2] ),
    .X(net3150));
 sg13g2_buf_2 fanout3151 (.A(net3152),
    .X(net3151));
 sg13g2_buf_2 fanout3152 (.A(net3153),
    .X(net3152));
 sg13g2_buf_2 fanout3153 (.A(\u_toplayer.u_layer2.neuron_index[2] ),
    .X(net3153));
 sg13g2_buf_2 fanout3154 (.A(\u_toplayer.u_layer3.u_neuron.acc[20] ),
    .X(net3154));
 sg13g2_buf_2 fanout3155 (.A(net1179),
    .X(net3155));
 sg13g2_buf_2 fanout3156 (.A(\u_toplayer.u_layer3.u_neuron.acc[16] ),
    .X(net3156));
 sg13g2_buf_2 fanout3157 (.A(net1167),
    .X(net3157));
 sg13g2_buf_4 fanout3158 (.X(net3158),
    .A(\u_toplayer.u_layer3.u_neuron.acc[8] ));
 sg13g2_buf_2 fanout3159 (.A(net1183),
    .X(net3159));
 sg13g2_buf_2 fanout3160 (.A(net3161),
    .X(net3160));
 sg13g2_buf_2 fanout3161 (.A(net3162),
    .X(net3161));
 sg13g2_buf_2 fanout3162 (.A(net1177),
    .X(net3162));
 sg13g2_buf_2 fanout3163 (.A(\u_toplayer.u_layer3.u_neuron.din[6] ),
    .X(net3163));
 sg13g2_buf_1 fanout3164 (.A(\u_toplayer.u_layer3.u_neuron.din[6] ),
    .X(net3164));
 sg13g2_buf_2 fanout3165 (.A(net3166),
    .X(net3165));
 sg13g2_buf_1 fanout3166 (.A(net3167),
    .X(net3166));
 sg13g2_buf_1 fanout3167 (.A(\u_toplayer.u_layer3.u_neuron.din[5] ),
    .X(net3167));
 sg13g2_buf_2 fanout3168 (.A(net3170),
    .X(net3168));
 sg13g2_buf_2 fanout3169 (.A(net3170),
    .X(net3169));
 sg13g2_buf_2 fanout3170 (.A(net1080),
    .X(net3170));
 sg13g2_buf_2 fanout3171 (.A(net3172),
    .X(net3171));
 sg13g2_buf_2 fanout3172 (.A(net3173),
    .X(net3172));
 sg13g2_buf_2 fanout3173 (.A(net1092),
    .X(net3173));
 sg13g2_buf_2 fanout3174 (.A(net3175),
    .X(net3174));
 sg13g2_buf_2 fanout3175 (.A(net1166),
    .X(net3175));
 sg13g2_buf_2 fanout3176 (.A(net3177),
    .X(net3176));
 sg13g2_buf_2 fanout3177 (.A(net1131),
    .X(net3177));
 sg13g2_buf_2 fanout3178 (.A(\u_toplayer.u_layer3.u_neuron.din[0] ),
    .X(net3178));
 sg13g2_buf_4 fanout3179 (.X(net3179),
    .A(\u_toplayer.u_outlayer.u_neuron.instCtrl.state[3] ));
 sg13g2_buf_2 fanout3180 (.A(\u_toplayer.u_outlayer.u_neuron.instCtrl.state[3] ),
    .X(net3180));
 sg13g2_buf_2 fanout3181 (.A(net3183),
    .X(net3181));
 sg13g2_buf_2 fanout3182 (.A(net3183),
    .X(net3182));
 sg13g2_buf_2 fanout3183 (.A(\u_toplayer.u_outlayer.u_neuron.instCtrl.state[2] ),
    .X(net3183));
 sg13g2_buf_2 fanout3184 (.A(net3186),
    .X(net3184));
 sg13g2_buf_2 fanout3185 (.A(net3186),
    .X(net3185));
 sg13g2_buf_4 fanout3186 (.X(net3186),
    .A(\u_toplayer.u_outlayer.u_neuron.instCtrl.state[1] ));
 sg13g2_buf_4 fanout3187 (.X(net3187),
    .A(net3188));
 sg13g2_buf_4 fanout3188 (.X(net3188),
    .A(net3191));
 sg13g2_buf_4 fanout3189 (.X(net3189),
    .A(net3190));
 sg13g2_buf_4 fanout3190 (.X(net3190),
    .A(net3191));
 sg13g2_buf_2 fanout3191 (.A(\u_toplayer.u_outlayer.u_neuron.instCtrl.state[0] ),
    .X(net3191));
 sg13g2_buf_2 fanout3192 (.A(net3193),
    .X(net3192));
 sg13g2_buf_4 fanout3193 (.X(net3193),
    .A(net3194));
 sg13g2_buf_2 fanout3194 (.A(net1059),
    .X(net3194));
 sg13g2_buf_2 fanout3195 (.A(net1208),
    .X(net3195));
 sg13g2_buf_2 fanout3196 (.A(net1196),
    .X(net3196));
 sg13g2_buf_2 fanout3197 (.A(\u_toplayer.u_outlayer.u_neuron.acc[16] ),
    .X(net3197));
 sg13g2_buf_2 fanout3198 (.A(net1201),
    .X(net3198));
 sg13g2_buf_2 fanout3199 (.A(net1184),
    .X(net3199));
 sg13g2_buf_2 fanout3200 (.A(net1202),
    .X(net3200));
 sg13g2_buf_2 fanout3201 (.A(net822),
    .X(net3201));
 sg13g2_buf_2 fanout3202 (.A(net3203),
    .X(net3202));
 sg13g2_buf_2 fanout3203 (.A(net3204),
    .X(net3203));
 sg13g2_buf_2 fanout3204 (.A(net1128),
    .X(net3204));
 sg13g2_buf_2 fanout3205 (.A(net3207),
    .X(net3205));
 sg13g2_buf_1 fanout3206 (.A(net3207),
    .X(net3206));
 sg13g2_buf_1 fanout3207 (.A(net3208),
    .X(net3207));
 sg13g2_buf_2 fanout3208 (.A(net1090),
    .X(net3208));
 sg13g2_buf_2 fanout3209 (.A(net3210),
    .X(net3209));
 sg13g2_buf_1 fanout3210 (.A(net3211),
    .X(net3210));
 sg13g2_buf_2 fanout3211 (.A(net1096),
    .X(net3211));
 sg13g2_buf_2 fanout3212 (.A(net3213),
    .X(net3212));
 sg13g2_buf_1 fanout3213 (.A(net3214),
    .X(net3213));
 sg13g2_buf_2 fanout3214 (.A(net1056),
    .X(net3214));
 sg13g2_buf_2 fanout3215 (.A(net3216),
    .X(net3215));
 sg13g2_buf_4 fanout3216 (.X(net3216),
    .A(net1148));
 sg13g2_buf_4 fanout3217 (.X(net3217),
    .A(net1138));
 sg13g2_buf_2 fanout3218 (.A(\u_toplayer.u_outlayer.u_neuron.din[3] ),
    .X(net3218));
 sg13g2_buf_2 fanout3219 (.A(net1123),
    .X(net3219));
 sg13g2_buf_2 fanout3220 (.A(\u_toplayer.u_outlayer.u_neuron.din[2] ),
    .X(net3220));
 sg13g2_buf_2 fanout3221 (.A(net3222),
    .X(net3221));
 sg13g2_buf_1 fanout3222 (.A(net3223),
    .X(net3222));
 sg13g2_buf_2 fanout3223 (.A(net1093),
    .X(net3223));
 sg13g2_buf_2 fanout3224 (.A(net3225),
    .X(net3224));
 sg13g2_buf_2 fanout3225 (.A(net1125),
    .X(net3225));
 sg13g2_buf_2 fanout3226 (.A(net3228),
    .X(net3226));
 sg13g2_buf_2 fanout3227 (.A(net3228),
    .X(net3227));
 sg13g2_buf_2 fanout3228 (.A(\u_toplayer.u_outlayer.u_neuron.mult[15] ),
    .X(net3228));
 sg13g2_buf_2 fanout3229 (.A(net968),
    .X(net3229));
 sg13g2_buf_4 fanout3230 (.X(net3230),
    .A(net1039));
 sg13g2_buf_2 fanout3231 (.A(net3233),
    .X(net3231));
 sg13g2_buf_1 fanout3232 (.A(net3233),
    .X(net3232));
 sg13g2_buf_1 fanout3233 (.A(net3234),
    .X(net3233));
 sg13g2_buf_2 fanout3234 (.A(\u_toplayer.u_layer2.u_neuron.instCtrl.state[4] ),
    .X(net3234));
 sg13g2_buf_2 fanout3235 (.A(net3236),
    .X(net3235));
 sg13g2_buf_2 fanout3236 (.A(net3237),
    .X(net3236));
 sg13g2_buf_1 fanout3237 (.A(net3238),
    .X(net3237));
 sg13g2_buf_2 fanout3238 (.A(\u_toplayer.u_layer2.u_neuron.instCtrl.state[3] ),
    .X(net3238));
 sg13g2_buf_2 fanout3239 (.A(net3240),
    .X(net3239));
 sg13g2_buf_2 fanout3240 (.A(net3241),
    .X(net3240));
 sg13g2_buf_2 fanout3241 (.A(net3242),
    .X(net3241));
 sg13g2_buf_2 fanout3242 (.A(net1134),
    .X(net3242));
 sg13g2_buf_2 fanout3243 (.A(net3245),
    .X(net3243));
 sg13g2_buf_1 fanout3244 (.A(net3245),
    .X(net3244));
 sg13g2_buf_2 fanout3245 (.A(net3248),
    .X(net3245));
 sg13g2_buf_2 fanout3246 (.A(net3247),
    .X(net3246));
 sg13g2_buf_2 fanout3247 (.A(net3248),
    .X(net3247));
 sg13g2_buf_2 fanout3248 (.A(\u_toplayer.u_layer2.u_neuron.instCtrl.state[1] ),
    .X(net3248));
 sg13g2_buf_2 fanout3249 (.A(net3250),
    .X(net3249));
 sg13g2_buf_2 fanout3250 (.A(net3251),
    .X(net3250));
 sg13g2_buf_2 fanout3251 (.A(net3252),
    .X(net3251));
 sg13g2_buf_2 fanout3252 (.A(\u_toplayer.u_layer2.u_neuron.instCtrl.state[1] ),
    .X(net3252));
 sg13g2_buf_2 fanout3253 (.A(net3255),
    .X(net3253));
 sg13g2_buf_2 fanout3254 (.A(net3255),
    .X(net3254));
 sg13g2_buf_2 fanout3255 (.A(\u_toplayer.u_layer2.u_neuron.instCtrl.state[1] ),
    .X(net3255));
 sg13g2_buf_2 fanout3256 (.A(net3257),
    .X(net3256));
 sg13g2_buf_2 fanout3257 (.A(net3258),
    .X(net3257));
 sg13g2_buf_2 fanout3258 (.A(net3259),
    .X(net3258));
 sg13g2_buf_2 fanout3259 (.A(net3264),
    .X(net3259));
 sg13g2_buf_2 fanout3260 (.A(net3264),
    .X(net3260));
 sg13g2_buf_1 fanout3261 (.A(net3262),
    .X(net3261));
 sg13g2_buf_2 fanout3262 (.A(net3264),
    .X(net3262));
 sg13g2_buf_2 fanout3263 (.A(net3264),
    .X(net3263));
 sg13g2_buf_2 fanout3264 (.A(\u_toplayer.u_layer2.u_neuron.instCtrl.state[0] ),
    .X(net3264));
 sg13g2_buf_2 fanout3265 (.A(net3268),
    .X(net3265));
 sg13g2_buf_2 fanout3266 (.A(net3268),
    .X(net3266));
 sg13g2_buf_2 fanout3267 (.A(net3268),
    .X(net3267));
 sg13g2_buf_2 fanout3268 (.A(net3272),
    .X(net3268));
 sg13g2_buf_2 fanout3269 (.A(net3272),
    .X(net3269));
 sg13g2_buf_2 fanout3270 (.A(net3272),
    .X(net3270));
 sg13g2_buf_1 fanout3271 (.A(net3272),
    .X(net3271));
 sg13g2_buf_2 fanout3272 (.A(\u_toplayer.u_layer2.u_neuron.instCtrl.state[0] ),
    .X(net3272));
 sg13g2_buf_2 fanout3273 (.A(net3274),
    .X(net3273));
 sg13g2_buf_2 fanout3274 (.A(net3277),
    .X(net3274));
 sg13g2_buf_2 fanout3275 (.A(net3277),
    .X(net3275));
 sg13g2_buf_2 fanout3276 (.A(net3277),
    .X(net3276));
 sg13g2_buf_2 fanout3277 (.A(\u_toplayer.u_layer2.u_neuron.instCtrl.state[0] ),
    .X(net3277));
 sg13g2_buf_2 fanout3278 (.A(_03930_),
    .X(net3278));
 sg13g2_buf_2 fanout3279 (.A(net3280),
    .X(net3279));
 sg13g2_buf_4 fanout3280 (.X(net3280),
    .A(_01049_));
 sg13g2_buf_2 fanout3281 (.A(net3283),
    .X(net3281));
 sg13g2_buf_2 fanout3282 (.A(net3283),
    .X(net3282));
 sg13g2_buf_4 fanout3283 (.X(net3283),
    .A(_01049_));
 sg13g2_buf_2 fanout3284 (.A(net3286),
    .X(net3284));
 sg13g2_buf_2 fanout3285 (.A(net3286),
    .X(net3285));
 sg13g2_buf_4 fanout3286 (.X(net3286),
    .A(uio_in[7]));
 sg13g2_buf_2 fanout3287 (.A(net3288),
    .X(net3287));
 sg13g2_buf_4 fanout3288 (.X(net3288),
    .A(net3292));
 sg13g2_buf_2 fanout3289 (.A(net3290),
    .X(net3289));
 sg13g2_buf_4 fanout3290 (.X(net3290),
    .A(net3291));
 sg13g2_buf_4 fanout3291 (.X(net3291),
    .A(net3292));
 sg13g2_buf_2 fanout3292 (.A(uio_in[6]),
    .X(net3292));
 sg13g2_buf_2 fanout3293 (.A(net3295),
    .X(net3293));
 sg13g2_buf_2 fanout3294 (.A(net3295),
    .X(net3294));
 sg13g2_buf_2 fanout3295 (.A(net3298),
    .X(net3295));
 sg13g2_buf_4 fanout3296 (.X(net3296),
    .A(net3297));
 sg13g2_buf_4 fanout3297 (.X(net3297),
    .A(net3298));
 sg13g2_buf_2 fanout3298 (.A(uio_in[5]),
    .X(net3298));
 sg13g2_buf_2 fanout3299 (.A(net3300),
    .X(net3299));
 sg13g2_buf_2 fanout3300 (.A(net3306),
    .X(net3300));
 sg13g2_buf_4 fanout3301 (.X(net3301),
    .A(net3306));
 sg13g2_buf_2 fanout3302 (.A(net3304),
    .X(net3302));
 sg13g2_buf_1 fanout3303 (.A(net3304),
    .X(net3303));
 sg13g2_buf_4 fanout3304 (.X(net3304),
    .A(net3306));
 sg13g2_buf_2 fanout3305 (.A(net3306),
    .X(net3305));
 sg13g2_buf_4 fanout3306 (.X(net3306),
    .A(uio_in[4]));
 sg13g2_buf_2 fanout3307 (.A(net3313),
    .X(net3307));
 sg13g2_buf_2 fanout3308 (.A(net3310),
    .X(net3308));
 sg13g2_buf_2 fanout3309 (.A(net3310),
    .X(net3309));
 sg13g2_buf_2 fanout3310 (.A(net3313),
    .X(net3310));
 sg13g2_buf_2 fanout3311 (.A(net3313),
    .X(net3311));
 sg13g2_buf_2 fanout3312 (.A(net3313),
    .X(net3312));
 sg13g2_buf_4 fanout3313 (.X(net3313),
    .A(net3320));
 sg13g2_buf_2 fanout3314 (.A(net3316),
    .X(net3314));
 sg13g2_buf_2 fanout3315 (.A(net3320),
    .X(net3315));
 sg13g2_buf_1 fanout3316 (.A(net3320),
    .X(net3316));
 sg13g2_buf_2 fanout3317 (.A(net3318),
    .X(net3317));
 sg13g2_buf_2 fanout3318 (.A(net3319),
    .X(net3318));
 sg13g2_buf_1 fanout3319 (.A(net3320),
    .X(net3319));
 sg13g2_buf_4 fanout3320 (.X(net3320),
    .A(uio_in[3]));
 sg13g2_buf_2 fanout3321 (.A(net3322),
    .X(net3321));
 sg13g2_buf_2 fanout3322 (.A(net3323),
    .X(net3322));
 sg13g2_buf_2 fanout3323 (.A(net3324),
    .X(net3323));
 sg13g2_buf_2 fanout3324 (.A(uio_in[2]),
    .X(net3324));
 sg13g2_buf_2 fanout3325 (.A(net3326),
    .X(net3325));
 sg13g2_buf_2 fanout3326 (.A(net3327),
    .X(net3326));
 sg13g2_buf_2 fanout3327 (.A(uio_in[2]),
    .X(net3327));
 sg13g2_buf_2 fanout3328 (.A(net3331),
    .X(net3328));
 sg13g2_buf_2 fanout3329 (.A(net3330),
    .X(net3329));
 sg13g2_buf_2 fanout3330 (.A(net3331),
    .X(net3330));
 sg13g2_buf_2 fanout3331 (.A(net3333),
    .X(net3331));
 sg13g2_buf_2 fanout3332 (.A(net3333),
    .X(net3332));
 sg13g2_buf_2 fanout3333 (.A(uio_in[2]),
    .X(net3333));
 sg13g2_buf_2 fanout3334 (.A(net3337),
    .X(net3334));
 sg13g2_buf_2 fanout3335 (.A(net3336),
    .X(net3335));
 sg13g2_buf_4 fanout3336 (.X(net3336),
    .A(net3337));
 sg13g2_buf_2 fanout3337 (.A(uio_in[1]),
    .X(net3337));
 sg13g2_buf_2 fanout3338 (.A(net3342),
    .X(net3338));
 sg13g2_buf_2 fanout3339 (.A(net3342),
    .X(net3339));
 sg13g2_buf_2 fanout3340 (.A(net3342),
    .X(net3340));
 sg13g2_buf_1 fanout3341 (.A(net3342),
    .X(net3341));
 sg13g2_buf_2 fanout3342 (.A(uio_in[1]),
    .X(net3342));
 sg13g2_buf_2 fanout3343 (.A(net3344),
    .X(net3343));
 sg13g2_buf_2 fanout3344 (.A(uio_in[1]),
    .X(net3344));
 sg13g2_buf_2 fanout3345 (.A(net3346),
    .X(net3345));
 sg13g2_buf_4 fanout3346 (.X(net3346),
    .A(net3347));
 sg13g2_buf_4 fanout3347 (.X(net3347),
    .A(net3));
 sg13g2_buf_2 fanout3348 (.A(net3350),
    .X(net3348));
 sg13g2_buf_2 fanout3349 (.A(net3350),
    .X(net3349));
 sg13g2_buf_1 fanout3350 (.A(net3356),
    .X(net3350));
 sg13g2_buf_2 fanout3351 (.A(net3356),
    .X(net3351));
 sg13g2_buf_2 fanout3352 (.A(net3356),
    .X(net3352));
 sg13g2_buf_2 fanout3353 (.A(net3355),
    .X(net3353));
 sg13g2_buf_1 fanout3354 (.A(net3355),
    .X(net3354));
 sg13g2_buf_4 fanout3355 (.X(net3355),
    .A(net3356));
 sg13g2_buf_2 fanout3356 (.A(net3),
    .X(net3356));
 sg13g2_buf_2 fanout3357 (.A(net3363),
    .X(net3357));
 sg13g2_buf_2 fanout3358 (.A(net3359),
    .X(net3358));
 sg13g2_buf_2 fanout3359 (.A(net3362),
    .X(net3359));
 sg13g2_buf_2 fanout3360 (.A(net3361),
    .X(net3360));
 sg13g2_buf_2 fanout3361 (.A(net3362),
    .X(net3361));
 sg13g2_buf_2 fanout3362 (.A(net3363),
    .X(net3362));
 sg13g2_buf_2 fanout3363 (.A(net2),
    .X(net3363));
 sg13g2_buf_4 fanout3364 (.X(net3364),
    .A(net3365));
 sg13g2_buf_1 fanout3365 (.A(net3366),
    .X(net3365));
 sg13g2_buf_2 fanout3366 (.A(net3369),
    .X(net3366));
 sg13g2_buf_2 fanout3367 (.A(net3369),
    .X(net3367));
 sg13g2_buf_2 fanout3368 (.A(net3369),
    .X(net3368));
 sg13g2_buf_2 fanout3369 (.A(net3379),
    .X(net3369));
 sg13g2_buf_2 fanout3370 (.A(net3375),
    .X(net3370));
 sg13g2_buf_2 fanout3371 (.A(net3375),
    .X(net3371));
 sg13g2_buf_2 fanout3372 (.A(net3374),
    .X(net3372));
 sg13g2_buf_1 fanout3373 (.A(net3374),
    .X(net3373));
 sg13g2_buf_2 fanout3374 (.A(net3375),
    .X(net3374));
 sg13g2_buf_2 fanout3375 (.A(net3376),
    .X(net3375));
 sg13g2_buf_2 fanout3376 (.A(net3379),
    .X(net3376));
 sg13g2_buf_2 fanout3377 (.A(net3378),
    .X(net3377));
 sg13g2_buf_4 fanout3378 (.X(net3378),
    .A(net3379));
 sg13g2_buf_2 fanout3379 (.A(net2),
    .X(net3379));
 sg13g2_buf_2 fanout3380 (.A(net3381),
    .X(net3380));
 sg13g2_buf_2 fanout3381 (.A(net3382),
    .X(net3381));
 sg13g2_buf_2 fanout3382 (.A(net3383),
    .X(net3382));
 sg13g2_buf_4 fanout3383 (.X(net3383),
    .A(net1));
 sg13g2_buf_2 fanout3384 (.A(net3385),
    .X(net3384));
 sg13g2_buf_4 fanout3385 (.X(net3385),
    .A(net3386));
 sg13g2_buf_4 fanout3386 (.X(net3386),
    .A(net3387));
 sg13g2_buf_2 fanout3387 (.A(ui_in[5]),
    .X(net3387));
 sg13g2_buf_2 fanout3388 (.A(net3389),
    .X(net3388));
 sg13g2_buf_2 fanout3389 (.A(net3390),
    .X(net3389));
 sg13g2_buf_8 fanout3390 (.A(ui_in[4]),
    .X(net3390));
 sg13g2_buf_2 fanout3391 (.A(net3392),
    .X(net3391));
 sg13g2_buf_2 fanout3392 (.A(net3393),
    .X(net3392));
 sg13g2_buf_8 fanout3393 (.A(ui_in[3]),
    .X(net3393));
 sg13g2_buf_2 fanout3394 (.A(net3395),
    .X(net3394));
 sg13g2_buf_2 fanout3395 (.A(net3396),
    .X(net3395));
 sg13g2_buf_4 fanout3396 (.X(net3396),
    .A(ui_in[2]));
 sg13g2_buf_2 fanout3397 (.A(net3398),
    .X(net3397));
 sg13g2_buf_4 fanout3398 (.X(net3398),
    .A(net3399));
 sg13g2_buf_4 fanout3399 (.X(net3399),
    .A(net3400));
 sg13g2_buf_4 fanout3400 (.X(net3400),
    .A(ui_in[1]));
 sg13g2_buf_2 fanout3401 (.A(net3402),
    .X(net3401));
 sg13g2_buf_2 fanout3402 (.A(net3403),
    .X(net3402));
 sg13g2_buf_4 fanout3403 (.X(net3403),
    .A(net3404));
 sg13g2_buf_4 fanout3404 (.X(net3404),
    .A(ui_in[0]));
 sg13g2_buf_4 fanout3405 (.X(net3405),
    .A(net3406));
 sg13g2_buf_4 fanout3406 (.X(net3406),
    .A(net3407));
 sg13g2_buf_4 fanout3407 (.X(net3407),
    .A(net3427));
 sg13g2_buf_4 fanout3408 (.X(net3408),
    .A(net3410));
 sg13g2_buf_4 fanout3409 (.X(net3409),
    .A(net3410));
 sg13g2_buf_4 fanout3410 (.X(net3410),
    .A(net3427));
 sg13g2_buf_4 fanout3411 (.X(net3411),
    .A(net3414));
 sg13g2_buf_4 fanout3412 (.X(net3412),
    .A(net3414));
 sg13g2_buf_4 fanout3413 (.X(net3413),
    .A(net3414));
 sg13g2_buf_2 fanout3414 (.A(net3427),
    .X(net3414));
 sg13g2_buf_4 fanout3415 (.X(net3415),
    .A(net3416));
 sg13g2_buf_4 fanout3416 (.X(net3416),
    .A(net3417));
 sg13g2_buf_4 fanout3417 (.X(net3417),
    .A(net3426));
 sg13g2_buf_4 fanout3418 (.X(net3418),
    .A(net3421));
 sg13g2_buf_4 fanout3419 (.X(net3419),
    .A(net3421));
 sg13g2_buf_2 fanout3420 (.A(net3421),
    .X(net3420));
 sg13g2_buf_2 fanout3421 (.A(net3426),
    .X(net3421));
 sg13g2_buf_4 fanout3422 (.X(net3422),
    .A(net3425));
 sg13g2_buf_2 fanout3423 (.A(net3425),
    .X(net3423));
 sg13g2_buf_4 fanout3424 (.X(net3424),
    .A(net3425));
 sg13g2_buf_2 fanout3425 (.A(net3426),
    .X(net3425));
 sg13g2_buf_2 fanout3426 (.A(net3427),
    .X(net3426));
 sg13g2_buf_2 fanout3427 (.A(net3487),
    .X(net3427));
 sg13g2_buf_4 fanout3428 (.X(net3428),
    .A(net3431));
 sg13g2_buf_4 fanout3429 (.X(net3429),
    .A(net3431));
 sg13g2_buf_4 fanout3430 (.X(net3430),
    .A(net3431));
 sg13g2_buf_2 fanout3431 (.A(net3443),
    .X(net3431));
 sg13g2_buf_4 fanout3432 (.X(net3432),
    .A(net3443));
 sg13g2_buf_2 fanout3433 (.A(net3434),
    .X(net3433));
 sg13g2_buf_4 fanout3434 (.X(net3434),
    .A(net3443));
 sg13g2_buf_4 fanout3435 (.X(net3435),
    .A(net3439));
 sg13g2_buf_2 fanout3436 (.A(net3439),
    .X(net3436));
 sg13g2_buf_4 fanout3437 (.X(net3437),
    .A(net3439));
 sg13g2_buf_2 fanout3438 (.A(net3439),
    .X(net3438));
 sg13g2_buf_2 fanout3439 (.A(net3443),
    .X(net3439));
 sg13g2_buf_4 fanout3440 (.X(net3440),
    .A(net3442));
 sg13g2_buf_4 fanout3441 (.X(net3441),
    .A(net3442));
 sg13g2_buf_2 fanout3442 (.A(net3443),
    .X(net3442));
 sg13g2_buf_2 fanout3443 (.A(net3487),
    .X(net3443));
 sg13g2_buf_4 fanout3444 (.X(net3444),
    .A(net3447));
 sg13g2_buf_2 fanout3445 (.A(net3447),
    .X(net3445));
 sg13g2_buf_4 fanout3446 (.X(net3446),
    .A(net3447));
 sg13g2_buf_2 fanout3447 (.A(net3456),
    .X(net3447));
 sg13g2_buf_4 fanout3448 (.X(net3448),
    .A(net3456));
 sg13g2_buf_2 fanout3449 (.A(net3456),
    .X(net3449));
 sg13g2_buf_4 fanout3450 (.X(net3450),
    .A(net3451));
 sg13g2_buf_4 fanout3451 (.X(net3451),
    .A(net3455));
 sg13g2_buf_4 fanout3452 (.X(net3452),
    .A(net3455));
 sg13g2_buf_4 fanout3453 (.X(net3453),
    .A(net3455));
 sg13g2_buf_4 fanout3454 (.X(net3454),
    .A(net3455));
 sg13g2_buf_2 fanout3455 (.A(net3456),
    .X(net3455));
 sg13g2_buf_2 fanout3456 (.A(net3487),
    .X(net3456));
 sg13g2_buf_4 fanout3457 (.X(net3457),
    .A(net3458));
 sg13g2_buf_4 fanout3458 (.X(net3458),
    .A(net3469));
 sg13g2_buf_4 fanout3459 (.X(net3459),
    .A(net3460));
 sg13g2_buf_4 fanout3460 (.X(net3460),
    .A(net3469));
 sg13g2_buf_4 fanout3461 (.X(net3461),
    .A(net3464));
 sg13g2_buf_2 fanout3462 (.A(net3464),
    .X(net3462));
 sg13g2_buf_4 fanout3463 (.X(net3463),
    .A(net3464));
 sg13g2_buf_2 fanout3464 (.A(net3469),
    .X(net3464));
 sg13g2_buf_4 fanout3465 (.X(net3465),
    .A(net3468));
 sg13g2_buf_4 fanout3466 (.X(net3466),
    .A(net3468));
 sg13g2_buf_2 fanout3467 (.A(net3468),
    .X(net3467));
 sg13g2_buf_2 fanout3468 (.A(net3469),
    .X(net3468));
 sg13g2_buf_2 fanout3469 (.A(net3487),
    .X(net3469));
 sg13g2_buf_4 fanout3470 (.X(net3470),
    .A(net3473));
 sg13g2_buf_4 fanout3471 (.X(net3471),
    .A(net3473));
 sg13g2_buf_4 fanout3472 (.X(net3472),
    .A(net3473));
 sg13g2_buf_2 fanout3473 (.A(net3477),
    .X(net3473));
 sg13g2_buf_4 fanout3474 (.X(net3474),
    .A(net3475));
 sg13g2_buf_4 fanout3475 (.X(net3475),
    .A(net3476));
 sg13g2_buf_4 fanout3476 (.X(net3476),
    .A(net3477));
 sg13g2_buf_2 fanout3477 (.A(net3487),
    .X(net3477));
 sg13g2_buf_4 fanout3478 (.X(net3478),
    .A(net3479));
 sg13g2_buf_2 fanout3479 (.A(net3482),
    .X(net3479));
 sg13g2_buf_4 fanout3480 (.X(net3480),
    .A(net3481));
 sg13g2_buf_4 fanout3481 (.X(net3481),
    .A(net3482));
 sg13g2_buf_4 fanout3482 (.X(net3482),
    .A(net3486));
 sg13g2_buf_4 fanout3483 (.X(net3483),
    .A(net3484));
 sg13g2_buf_4 fanout3484 (.X(net3484),
    .A(net3486));
 sg13g2_buf_8 fanout3485 (.A(net3486),
    .X(net3485));
 sg13g2_buf_4 fanout3486 (.X(net3486),
    .A(net3487));
 sg13g2_buf_8 fanout3487 (.A(rst_n),
    .X(net3487));
 sg13g2_buf_4 fanout3488 (.X(net3488),
    .A(net3492));
 sg13g2_buf_2 fanout3489 (.A(net3492),
    .X(net3489));
 sg13g2_buf_4 fanout3490 (.X(net3490),
    .A(net3492));
 sg13g2_buf_4 fanout3491 (.X(net3491),
    .A(net3492));
 sg13g2_buf_2 fanout3492 (.A(net3505),
    .X(net3492));
 sg13g2_buf_4 fanout3493 (.X(net3493),
    .A(net3496));
 sg13g2_buf_4 fanout3494 (.X(net3494),
    .A(net3496));
 sg13g2_buf_4 fanout3495 (.X(net3495),
    .A(net3496));
 sg13g2_buf_2 fanout3496 (.A(net3505),
    .X(net3496));
 sg13g2_buf_4 fanout3497 (.X(net3497),
    .A(net3500));
 sg13g2_buf_4 fanout3498 (.X(net3498),
    .A(net3500));
 sg13g2_buf_2 fanout3499 (.A(net3500),
    .X(net3499));
 sg13g2_buf_2 fanout3500 (.A(net3505),
    .X(net3500));
 sg13g2_buf_4 fanout3501 (.X(net3501),
    .A(net3504));
 sg13g2_buf_4 fanout3502 (.X(net3502),
    .A(net3504));
 sg13g2_buf_2 fanout3503 (.A(net3504),
    .X(net3503));
 sg13g2_buf_2 fanout3504 (.A(net3505),
    .X(net3504));
 sg13g2_buf_2 fanout3505 (.A(net3564),
    .X(net3505));
 sg13g2_buf_4 fanout3506 (.X(net3506),
    .A(net3507));
 sg13g2_buf_4 fanout3507 (.X(net3507),
    .A(net3509));
 sg13g2_buf_4 fanout3508 (.X(net3508),
    .A(net3509));
 sg13g2_buf_2 fanout3509 (.A(net3515),
    .X(net3509));
 sg13g2_buf_4 fanout3510 (.X(net3510),
    .A(net3511));
 sg13g2_buf_4 fanout3511 (.X(net3511),
    .A(net3515));
 sg13g2_buf_4 fanout3512 (.X(net3512),
    .A(net3514));
 sg13g2_buf_4 fanout3513 (.X(net3513),
    .A(net3514));
 sg13g2_buf_4 fanout3514 (.X(net3514),
    .A(net3515));
 sg13g2_buf_2 fanout3515 (.A(net3564),
    .X(net3515));
 sg13g2_buf_4 fanout3516 (.X(net3516),
    .A(net3520));
 sg13g2_buf_2 fanout3517 (.A(net3520),
    .X(net3517));
 sg13g2_buf_4 fanout3518 (.X(net3518),
    .A(net3520));
 sg13g2_buf_2 fanout3519 (.A(net3520),
    .X(net3519));
 sg13g2_buf_2 fanout3520 (.A(net3548),
    .X(net3520));
 sg13g2_buf_4 fanout3521 (.X(net3521),
    .A(net3523));
 sg13g2_buf_4 fanout3522 (.X(net3522),
    .A(net3523));
 sg13g2_buf_4 fanout3523 (.X(net3523),
    .A(net3548));
 sg13g2_buf_4 fanout3524 (.X(net3524),
    .A(net3526));
 sg13g2_buf_2 fanout3525 (.A(net3526),
    .X(net3525));
 sg13g2_buf_4 fanout3526 (.X(net3526),
    .A(net3531));
 sg13g2_buf_4 fanout3527 (.X(net3527),
    .A(net3531));
 sg13g2_buf_4 fanout3528 (.X(net3528),
    .A(net3531));
 sg13g2_buf_4 fanout3529 (.X(net3529),
    .A(net3530));
 sg13g2_buf_4 fanout3530 (.X(net3530),
    .A(net3531));
 sg13g2_buf_2 fanout3531 (.A(net3548),
    .X(net3531));
 sg13g2_buf_4 fanout3532 (.X(net3532),
    .A(net3536));
 sg13g2_buf_2 fanout3533 (.A(net3536),
    .X(net3533));
 sg13g2_buf_4 fanout3534 (.X(net3534),
    .A(net3536));
 sg13g2_buf_2 fanout3535 (.A(net3536),
    .X(net3535));
 sg13g2_buf_1 fanout3536 (.A(net3548),
    .X(net3536));
 sg13g2_buf_4 fanout3537 (.X(net3537),
    .A(net3540));
 sg13g2_buf_4 fanout3538 (.X(net3538),
    .A(net3540));
 sg13g2_buf_4 fanout3539 (.X(net3539),
    .A(net3540));
 sg13g2_buf_2 fanout3540 (.A(net3548),
    .X(net3540));
 sg13g2_buf_4 fanout3541 (.X(net3541),
    .A(net3544));
 sg13g2_buf_4 fanout3542 (.X(net3542),
    .A(net3543));
 sg13g2_buf_4 fanout3543 (.X(net3543),
    .A(net3544));
 sg13g2_buf_2 fanout3544 (.A(net3547),
    .X(net3544));
 sg13g2_buf_4 fanout3545 (.X(net3545),
    .A(net3547));
 sg13g2_buf_4 fanout3546 (.X(net3546),
    .A(net3547));
 sg13g2_buf_2 fanout3547 (.A(net3548),
    .X(net3547));
 sg13g2_buf_4 fanout3548 (.X(net3548),
    .A(net3564));
 sg13g2_buf_4 fanout3549 (.X(net3549),
    .A(net3550));
 sg13g2_buf_4 fanout3550 (.X(net3550),
    .A(net3552));
 sg13g2_buf_4 fanout3551 (.X(net3551),
    .A(net3552));
 sg13g2_buf_4 fanout3552 (.X(net3552),
    .A(net3563));
 sg13g2_buf_4 fanout3553 (.X(net3553),
    .A(net3554));
 sg13g2_buf_4 fanout3554 (.X(net3554),
    .A(net3555));
 sg13g2_buf_4 fanout3555 (.X(net3555),
    .A(net3563));
 sg13g2_buf_4 fanout3556 (.X(net3556),
    .A(net3558));
 sg13g2_buf_4 fanout3557 (.X(net3557),
    .A(net3560));
 sg13g2_buf_2 fanout3558 (.A(net3560),
    .X(net3558));
 sg13g2_buf_4 fanout3559 (.X(net3559),
    .A(net3560));
 sg13g2_buf_2 fanout3560 (.A(net3563),
    .X(net3560));
 sg13g2_buf_4 fanout3561 (.X(net3561),
    .A(net3563));
 sg13g2_buf_2 fanout3562 (.A(net3563),
    .X(net3562));
 sg13g2_buf_4 fanout3563 (.X(net3563),
    .A(net3564));
 sg13g2_buf_2 fanout3564 (.A(rst_n),
    .X(net3564));
 sg13g2_buf_2 input1 (.A(ui_in[6]),
    .X(net1));
 sg13g2_buf_4 input2 (.X(net2),
    .A(ui_in[7]));
 sg13g2_buf_2 input3 (.A(uio_in[0]),
    .X(net3));
 sg13g2_tielo tt_um_neural_navigators_4 (.L_LO(net4));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_buf_2 clkbuf_leaf_0_clk_regs (.A(clknet_4_1_0_clk_regs),
    .X(clknet_leaf_0_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_1_clk_regs (.A(clknet_4_1_0_clk_regs),
    .X(clknet_leaf_1_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_2_clk_regs (.A(clknet_4_1_0_clk_regs),
    .X(clknet_leaf_2_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_3_clk_regs (.A(clknet_4_0_0_clk_regs),
    .X(clknet_leaf_3_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_4_clk_regs (.A(clknet_4_0_0_clk_regs),
    .X(clknet_leaf_4_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_5_clk_regs (.A(clknet_4_1_0_clk_regs),
    .X(clknet_leaf_5_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_6_clk_regs (.A(clknet_4_1_0_clk_regs),
    .X(clknet_leaf_6_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_7_clk_regs (.A(clknet_4_1_0_clk_regs),
    .X(clknet_leaf_7_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_8_clk_regs (.A(clknet_4_1_0_clk_regs),
    .X(clknet_leaf_8_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_9_clk_regs (.A(clknet_4_4_0_clk_regs),
    .X(clknet_leaf_9_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_10_clk_regs (.A(clknet_4_4_0_clk_regs),
    .X(clknet_leaf_10_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_11_clk_regs (.A(clknet_4_4_0_clk_regs),
    .X(clknet_leaf_11_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_12_clk_regs (.A(clknet_4_4_0_clk_regs),
    .X(clknet_leaf_12_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_13_clk_regs (.A(clknet_4_6_0_clk_regs),
    .X(clknet_leaf_13_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_14_clk_regs (.A(clknet_4_6_0_clk_regs),
    .X(clknet_leaf_14_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_15_clk_regs (.A(clknet_4_6_0_clk_regs),
    .X(clknet_leaf_15_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_16_clk_regs (.A(clknet_4_6_0_clk_regs),
    .X(clknet_leaf_16_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_17_clk_regs (.A(clknet_4_6_0_clk_regs),
    .X(clknet_leaf_17_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_18_clk_regs (.A(clknet_4_7_0_clk_regs),
    .X(clknet_leaf_18_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_19_clk_regs (.A(clknet_4_7_0_clk_regs),
    .X(clknet_leaf_19_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_20_clk_regs (.A(clknet_4_4_0_clk_regs),
    .X(clknet_leaf_20_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_21_clk_regs (.A(clknet_4_4_0_clk_regs),
    .X(clknet_leaf_21_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_22_clk_regs (.A(clknet_4_5_0_clk_regs),
    .X(clknet_leaf_22_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_23_clk_regs (.A(clknet_4_5_0_clk_regs),
    .X(clknet_leaf_23_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_24_clk_regs (.A(clknet_4_5_0_clk_regs),
    .X(clknet_leaf_24_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_25_clk_regs (.A(clknet_4_5_0_clk_regs),
    .X(clknet_leaf_25_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_26_clk_regs (.A(clknet_4_5_0_clk_regs),
    .X(clknet_leaf_26_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_27_clk_regs (.A(clknet_4_4_0_clk_regs),
    .X(clknet_leaf_27_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_28_clk_regs (.A(clknet_4_5_0_clk_regs),
    .X(clknet_leaf_28_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_29_clk_regs (.A(clknet_4_5_0_clk_regs),
    .X(clknet_leaf_29_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_30_clk_regs (.A(clknet_4_7_0_clk_regs),
    .X(clknet_leaf_30_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_31_clk_regs (.A(clknet_4_7_0_clk_regs),
    .X(clknet_leaf_31_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_32_clk_regs (.A(clknet_4_7_0_clk_regs),
    .X(clknet_leaf_32_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_33_clk_regs (.A(clknet_4_7_0_clk_regs),
    .X(clknet_leaf_33_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_34_clk_regs (.A(clknet_4_7_0_clk_regs),
    .X(clknet_leaf_34_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_35_clk_regs (.A(clknet_4_13_0_clk_regs),
    .X(clknet_leaf_35_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_36_clk_regs (.A(clknet_4_14_0_clk_regs),
    .X(clknet_leaf_36_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_37_clk_regs (.A(clknet_4_14_0_clk_regs),
    .X(clknet_leaf_37_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_38_clk_regs (.A(clknet_4_14_0_clk_regs),
    .X(clknet_leaf_38_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_39_clk_regs (.A(clknet_4_15_0_clk_regs),
    .X(clknet_leaf_39_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_40_clk_regs (.A(clknet_4_15_0_clk_regs),
    .X(clknet_leaf_40_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_41_clk_regs (.A(clknet_4_15_0_clk_regs),
    .X(clknet_leaf_41_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_42_clk_regs (.A(clknet_4_15_0_clk_regs),
    .X(clknet_leaf_42_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_43_clk_regs (.A(clknet_4_15_0_clk_regs),
    .X(clknet_leaf_43_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_44_clk_regs (.A(clknet_4_15_0_clk_regs),
    .X(clknet_leaf_44_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_45_clk_regs (.A(clknet_4_15_0_clk_regs),
    .X(clknet_leaf_45_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_46_clk_regs (.A(clknet_4_14_0_clk_regs),
    .X(clknet_leaf_46_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_47_clk_regs (.A(clknet_4_14_0_clk_regs),
    .X(clknet_leaf_47_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_48_clk_regs (.A(clknet_4_14_0_clk_regs),
    .X(clknet_leaf_48_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_49_clk_regs (.A(clknet_4_13_0_clk_regs),
    .X(clknet_leaf_49_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_50_clk_regs (.A(clknet_4_13_0_clk_regs),
    .X(clknet_leaf_50_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_51_clk_regs (.A(clknet_4_13_0_clk_regs),
    .X(clknet_leaf_51_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_52_clk_regs (.A(clknet_4_14_0_clk_regs),
    .X(clknet_leaf_52_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_53_clk_regs (.A(clknet_4_13_0_clk_regs),
    .X(clknet_leaf_53_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_54_clk_regs (.A(clknet_4_12_0_clk_regs),
    .X(clknet_leaf_54_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_55_clk_regs (.A(clknet_4_11_0_clk_regs),
    .X(clknet_leaf_55_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_56_clk_regs (.A(clknet_4_11_0_clk_regs),
    .X(clknet_leaf_56_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_57_clk_regs (.A(clknet_4_13_0_clk_regs),
    .X(clknet_leaf_57_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_58_clk_regs (.A(clknet_4_11_0_clk_regs),
    .X(clknet_leaf_58_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_59_clk_regs (.A(clknet_4_11_0_clk_regs),
    .X(clknet_leaf_59_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_60_clk_regs (.A(clknet_4_11_0_clk_regs),
    .X(clknet_leaf_60_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_61_clk_regs (.A(clknet_4_11_0_clk_regs),
    .X(clknet_leaf_61_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_62_clk_regs (.A(clknet_4_11_0_clk_regs),
    .X(clknet_leaf_62_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_63_clk_regs (.A(clknet_4_10_0_clk_regs),
    .X(clknet_leaf_63_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_64_clk_regs (.A(clknet_4_10_0_clk_regs),
    .X(clknet_leaf_64_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_65_clk_regs (.A(clknet_4_9_0_clk_regs),
    .X(clknet_leaf_65_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_66_clk_regs (.A(clknet_4_9_0_clk_regs),
    .X(clknet_leaf_66_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_67_clk_regs (.A(clknet_4_10_0_clk_regs),
    .X(clknet_leaf_67_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_68_clk_regs (.A(clknet_4_10_0_clk_regs),
    .X(clknet_leaf_68_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_69_clk_regs (.A(clknet_4_10_0_clk_regs),
    .X(clknet_leaf_69_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_70_clk_regs (.A(clknet_4_10_0_clk_regs),
    .X(clknet_leaf_70_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_71_clk_regs (.A(clknet_4_10_0_clk_regs),
    .X(clknet_leaf_71_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_72_clk_regs (.A(clknet_4_9_0_clk_regs),
    .X(clknet_leaf_72_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_73_clk_regs (.A(clknet_4_9_0_clk_regs),
    .X(clknet_leaf_73_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_74_clk_regs (.A(clknet_4_9_0_clk_regs),
    .X(clknet_leaf_74_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_75_clk_regs (.A(clknet_4_9_0_clk_regs),
    .X(clknet_leaf_75_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_76_clk_regs (.A(clknet_4_9_0_clk_regs),
    .X(clknet_leaf_76_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_77_clk_regs (.A(clknet_4_8_0_clk_regs),
    .X(clknet_leaf_77_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_78_clk_regs (.A(clknet_4_8_0_clk_regs),
    .X(clknet_leaf_78_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_79_clk_regs (.A(clknet_4_8_0_clk_regs),
    .X(clknet_leaf_79_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_80_clk_regs (.A(clknet_4_8_0_clk_regs),
    .X(clknet_leaf_80_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_81_clk_regs (.A(clknet_4_8_0_clk_regs),
    .X(clknet_leaf_81_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_82_clk_regs (.A(clknet_4_8_0_clk_regs),
    .X(clknet_leaf_82_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_83_clk_regs (.A(clknet_4_12_0_clk_regs),
    .X(clknet_leaf_83_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_84_clk_regs (.A(clknet_4_12_0_clk_regs),
    .X(clknet_leaf_84_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_85_clk_regs (.A(clknet_4_8_0_clk_regs),
    .X(clknet_leaf_85_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_86_clk_regs (.A(clknet_4_12_0_clk_regs),
    .X(clknet_leaf_86_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_87_clk_regs (.A(clknet_4_12_0_clk_regs),
    .X(clknet_leaf_87_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_88_clk_regs (.A(clknet_4_12_0_clk_regs),
    .X(clknet_leaf_88_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_90_clk_regs (.A(clknet_4_13_0_clk_regs),
    .X(clknet_leaf_90_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_91_clk_regs (.A(clknet_4_6_0_clk_regs),
    .X(clknet_leaf_91_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_92_clk_regs (.A(clknet_4_3_0_clk_regs),
    .X(clknet_leaf_92_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_93_clk_regs (.A(clknet_4_3_0_clk_regs),
    .X(clknet_leaf_93_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_94_clk_regs (.A(clknet_4_3_0_clk_regs),
    .X(clknet_leaf_94_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_95_clk_regs (.A(clknet_4_3_0_clk_regs),
    .X(clknet_leaf_95_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_96_clk_regs (.A(clknet_4_3_0_clk_regs),
    .X(clknet_leaf_96_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_97_clk_regs (.A(clknet_4_3_0_clk_regs),
    .X(clknet_leaf_97_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_98_clk_regs (.A(clknet_4_3_0_clk_regs),
    .X(clknet_leaf_98_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_99_clk_regs (.A(clknet_4_2_0_clk_regs),
    .X(clknet_leaf_99_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_100_clk_regs (.A(clknet_4_2_0_clk_regs),
    .X(clknet_leaf_100_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_101_clk_regs (.A(clknet_4_2_0_clk_regs),
    .X(clknet_leaf_101_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_102_clk_regs (.A(clknet_4_2_0_clk_regs),
    .X(clknet_leaf_102_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_103_clk_regs (.A(clknet_4_2_0_clk_regs),
    .X(clknet_leaf_103_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_104_clk_regs (.A(clknet_4_2_0_clk_regs),
    .X(clknet_leaf_104_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_105_clk_regs (.A(clknet_4_0_0_clk_regs),
    .X(clknet_leaf_105_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_106_clk_regs (.A(clknet_4_2_0_clk_regs),
    .X(clknet_leaf_106_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_107_clk_regs (.A(clknet_4_6_0_clk_regs),
    .X(clknet_leaf_107_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_108_clk_regs (.A(clknet_4_0_0_clk_regs),
    .X(clknet_leaf_108_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_109_clk_regs (.A(clknet_4_0_0_clk_regs),
    .X(clknet_leaf_109_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_110_clk_regs (.A(clknet_4_0_0_clk_regs),
    .X(clknet_leaf_110_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_111_clk_regs (.A(clknet_4_0_0_clk_regs),
    .X(clknet_leaf_111_clk_regs));
 sg13g2_buf_2 clkbuf_0_clk_regs (.A(clk_regs),
    .X(clknet_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_0_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_0_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_1_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_1_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_2_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_2_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_3_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_3_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_4_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_4_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_5_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_5_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_6_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_6_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_7_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_7_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_8_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_8_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_9_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_9_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_10_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_10_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_11_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_11_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_12_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_12_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_13_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_13_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_14_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_14_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_15_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_15_0_clk_regs));
 sg13g2_buf_1 clkload0 (.A(clknet_4_0_0_clk_regs));
 sg13g2_buf_1 clkload1 (.A(clknet_4_1_0_clk_regs));
 sg13g2_buf_1 clkload2 (.A(clknet_4_2_0_clk_regs));
 sg13g2_buf_1 clkload3 (.A(clknet_4_3_0_clk_regs));
 sg13g2_buf_1 clkload4 (.A(clknet_4_4_0_clk_regs));
 sg13g2_buf_1 clkload5 (.A(clknet_4_5_0_clk_regs));
 sg13g2_buf_1 clkload6 (.A(clknet_4_6_0_clk_regs));
 sg13g2_buf_1 clkload7 (.A(clknet_4_7_0_clk_regs));
 sg13g2_buf_1 clkload8 (.A(clknet_4_8_0_clk_regs));
 sg13g2_buf_1 clkload9 (.A(clknet_4_9_0_clk_regs));
 sg13g2_buf_1 clkload10 (.A(clknet_4_10_0_clk_regs));
 sg13g2_buf_1 clkload11 (.A(clknet_4_11_0_clk_regs));
 sg13g2_buf_1 clkload12 (.A(clknet_4_13_0_clk_regs));
 sg13g2_buf_1 clkload13 (.A(clknet_4_14_0_clk_regs));
 sg13g2_buf_1 clkload14 (.A(clknet_4_15_0_clk_regs));
 sg13g2_inv_1 clkload15 (.A(clknet_leaf_111_clk_regs));
 sg13g2_inv_1 clkload16 (.A(clknet_leaf_103_clk_regs));
 sg13g2_inv_1 clkload17 (.A(clknet_leaf_92_clk_regs));
 sg13g2_inv_1 clkload18 (.A(clknet_leaf_9_clk_regs));
 sg13g2_inv_4 clkload19 (.A(clknet_leaf_20_clk_regs));
 sg13g2_inv_1 clkload20 (.A(clknet_leaf_27_clk_regs));
 sg13g2_inv_4 clkload21 (.A(clknet_leaf_22_clk_regs));
 sg13g2_inv_4 clkload22 (.A(clknet_leaf_23_clk_regs));
 sg13g2_inv_1 clkload23 (.A(clknet_leaf_24_clk_regs));
 sg13g2_inv_8 clkload24 (.A(clknet_leaf_28_clk_regs));
 sg13g2_inv_1 clkload25 (.A(clknet_leaf_29_clk_regs));
 sg13g2_inv_4 clkload26 (.A(clknet_leaf_17_clk_regs));
 sg13g2_inv_4 clkload27 (.A(clknet_leaf_91_clk_regs));
 sg13g2_inv_8 clkload28 (.A(clknet_leaf_19_clk_regs));
 sg13g2_inv_4 clkload29 (.A(clknet_leaf_30_clk_regs));
 sg13g2_inv_8 clkload30 (.A(clknet_leaf_32_clk_regs));
 sg13g2_inv_4 clkload31 (.A(clknet_leaf_33_clk_regs));
 sg13g2_inv_1 clkload32 (.A(clknet_leaf_34_clk_regs));
 sg13g2_inv_2 clkload33 (.A(clknet_leaf_77_clk_regs));
 sg13g2_inv_1 clkload34 (.A(clknet_leaf_54_clk_regs));
 sg13g2_inv_4 clkload35 (.A(clknet_leaf_35_clk_regs));
 sg13g2_inv_2 clkload36 (.A(clknet_leaf_49_clk_regs));
 sg13g2_inv_4 clkload37 (.A(clknet_leaf_90_clk_regs));
 sg13g2_inv_4 clkload38 (.A(clknet_leaf_46_clk_regs));
 sg13g2_inv_1 clkload39 (.A(clknet_leaf_47_clk_regs));
 sg13g2_inv_4 clkload40 (.A(clknet_leaf_48_clk_regs));
 sg13g2_inv_1 clkload41 (.A(clknet_leaf_39_clk_regs));
 sg13g2_inv_4 clkload42 (.A(clknet_leaf_40_clk_regs));
 sg13g2_inv_2 clkload43 (.A(clknet_leaf_41_clk_regs));
 sg13g2_inv_1 clkload44 (.A(clknet_leaf_43_clk_regs));
 sg13g2_inv_1 clkload45 (.A(clknet_leaf_44_clk_regs));
 sg13g2_inv_4 clkload46 (.A(clknet_leaf_45_clk_regs));
 sg13g2_dlygate4sd3_1 hold1 (.A(_00033_),
    .X(net116));
 sg13g2_dlygate4sd3_1 hold2 (.A(_00348_),
    .X(net117));
 sg13g2_dlygate4sd3_1 hold3 (.A(_00043_),
    .X(net118));
 sg13g2_dlygate4sd3_1 hold4 (.A(_00000_),
    .X(net119));
 sg13g2_dlygate4sd3_1 hold5 (.A(\u_toplayer.u_layer3.stateout[7] ),
    .X(net120));
 sg13g2_dlygate4sd3_1 hold6 (.A(\u_toplayer.u_layer3.stateout[6] ),
    .X(net121));
 sg13g2_dlygate4sd3_1 hold7 (.A(_00031_),
    .X(net122));
 sg13g2_dlygate4sd3_1 hold8 (.A(_00676_),
    .X(net123));
 sg13g2_dlygate4sd3_1 hold9 (.A(\u_toplayer.delay_counter_layer1[0] ),
    .X(net124));
 sg13g2_dlygate4sd3_1 hold10 (.A(_01014_),
    .X(net125));
 sg13g2_dlygate4sd3_1 hold11 (.A(\u_toplayer.delay_counter_layer3[0] ),
    .X(net126));
 sg13g2_dlygate4sd3_1 hold12 (.A(_00707_),
    .X(net127));
 sg13g2_dlygate4sd3_1 hold13 (.A(\u_toplayer.u_layer2.statel2[6] ),
    .X(net128));
 sg13g2_dlygate4sd3_1 hold14 (.A(\u_toplayer.outreg[38] ),
    .X(net129));
 sg13g2_dlygate4sd3_1 hold15 (.A(\u_toplayer.delay_counter_layer2[0] ),
    .X(net130));
 sg13g2_dlygate4sd3_1 hold16 (.A(_01016_),
    .X(net131));
 sg13g2_dlygate4sd3_1 hold17 (.A(\u_toplayer.u_layer2.statel2[7] ),
    .X(net132));
 sg13g2_dlygate4sd3_1 hold18 (.A(\u_toplayer.outreg[32] ),
    .X(net133));
 sg13g2_dlygate4sd3_1 hold19 (.A(\u_toplayer.outreg[37] ),
    .X(net134));
 sg13g2_dlygate4sd3_1 hold20 (.A(\u_toplayer.outreg[39] ),
    .X(net135));
 sg13g2_dlygate4sd3_1 hold21 (.A(_00282_),
    .X(net136));
 sg13g2_dlygate4sd3_1 hold22 (.A(\u_toplayer.outreg[34] ),
    .X(net137));
 sg13g2_dlygate4sd3_1 hold23 (.A(\u_toplayer.outreg[36] ),
    .X(net138));
 sg13g2_dlygate4sd3_1 hold24 (.A(\u_toplayer.outreg[43] ),
    .X(net139));
 sg13g2_dlygate4sd3_1 hold25 (.A(\u_toplayer.outreg[20] ),
    .X(net140));
 sg13g2_dlygate4sd3_1 hold26 (.A(\u_toplayer.outreg[11] ),
    .X(net141));
 sg13g2_dlygate4sd3_1 hold27 (.A(\u_toplayer.outreg[74] ),
    .X(net142));
 sg13g2_dlygate4sd3_1 hold28 (.A(\u_toplayer.outreg[21] ),
    .X(net143));
 sg13g2_dlygate4sd3_1 hold29 (.A(\u_toplayer.outreg[47] ),
    .X(net144));
 sg13g2_dlygate4sd3_1 hold30 (.A(\u_toplayer.outreg[24] ),
    .X(net145));
 sg13g2_dlygate4sd3_1 hold31 (.A(\u_toplayer.outreg[33] ),
    .X(net146));
 sg13g2_dlygate4sd3_1 hold32 (.A(\u_toplayer.outreg[44] ),
    .X(net147));
 sg13g2_dlygate4sd3_1 hold33 (.A(\u_toplayer.outreg[79] ),
    .X(net148));
 sg13g2_dlygate4sd3_1 hold34 (.A(\u_toplayer.outreg[13] ),
    .X(net149));
 sg13g2_dlygate4sd3_1 hold35 (.A(\u_toplayer.outreg[8] ),
    .X(net150));
 sg13g2_dlygate4sd3_1 hold36 (.A(\u_toplayer.outreg[12] ),
    .X(net151));
 sg13g2_dlygate4sd3_1 hold37 (.A(\u_toplayer.outreg[40] ),
    .X(net152));
 sg13g2_dlygate4sd3_1 hold38 (.A(\u_toplayer.outreg[31] ),
    .X(net153));
 sg13g2_dlygate4sd3_1 hold39 (.A(_00274_),
    .X(net154));
 sg13g2_dlygate4sd3_1 hold40 (.A(\u_toplayer.outreg[14] ),
    .X(net155));
 sg13g2_dlygate4sd3_1 hold41 (.A(_00257_),
    .X(net156));
 sg13g2_dlygate4sd3_1 hold42 (.A(\u_toplayer.outreg[17] ),
    .X(net157));
 sg13g2_dlygate4sd3_1 hold43 (.A(\u_toplayer.outreg[72] ),
    .X(net158));
 sg13g2_dlygate4sd3_1 hold44 (.A(\u_toplayer.outreg[45] ),
    .X(net159));
 sg13g2_dlygate4sd3_1 hold45 (.A(\u_toplayer.outreg[29] ),
    .X(net160));
 sg13g2_dlygate4sd3_1 hold46 (.A(\u_toplayer.outreg[35] ),
    .X(net161));
 sg13g2_dlygate4sd3_1 hold47 (.A(\u_toplayer.outreg[42] ),
    .X(net162));
 sg13g2_dlygate4sd3_1 hold48 (.A(\u_toplayer.reg_layer2[218] ),
    .X(net163));
 sg13g2_dlygate4sd3_1 hold49 (.A(\u_toplayer.outreg[0] ),
    .X(net164));
 sg13g2_dlygate4sd3_1 hold50 (.A(\u_toplayer.outreg[4] ),
    .X(net165));
 sg13g2_dlygate4sd3_1 hold51 (.A(\u_toplayer.reg_layer2[92] ),
    .X(net166));
 sg13g2_dlygate4sd3_1 hold52 (.A(\u_toplayer.reg_layer1[251] ),
    .X(net167));
 sg13g2_dlygate4sd3_1 hold53 (.A(\u_toplayer.outreg[19] ),
    .X(net168));
 sg13g2_dlygate4sd3_1 hold54 (.A(\u_toplayer.reg_layer1[47] ),
    .X(net169));
 sg13g2_dlygate4sd3_1 hold55 (.A(\u_toplayer.outreg[25] ),
    .X(net170));
 sg13g2_dlygate4sd3_1 hold56 (.A(\u_toplayer.outreg[18] ),
    .X(net171));
 sg13g2_dlygate4sd3_1 hold57 (.A(\u_toplayer.reg_layer2[38] ),
    .X(net172));
 sg13g2_dlygate4sd3_1 hold58 (.A(_00433_),
    .X(net173));
 sg13g2_dlygate4sd3_1 hold59 (.A(\u_toplayer.reg_layer2[168] ),
    .X(net174));
 sg13g2_dlygate4sd3_1 hold60 (.A(\u_toplayer.reg_layer1[62] ),
    .X(net175));
 sg13g2_dlygate4sd3_1 hold61 (.A(\u_toplayer.reg_layer2[154] ),
    .X(net176));
 sg13g2_dlygate4sd3_1 hold62 (.A(\u_toplayer.outreg[6] ),
    .X(net177));
 sg13g2_dlygate4sd3_1 hold63 (.A(\u_toplayer.reg_layer1[56] ),
    .X(net178));
 sg13g2_dlygate4sd3_1 hold64 (.A(\u_toplayer.reg_layer1[121] ),
    .X(net179));
 sg13g2_dlygate4sd3_1 hold65 (.A(_00830_),
    .X(net180));
 sg13g2_dlygate4sd3_1 hold66 (.A(\u_toplayer.reg_layer1[186] ),
    .X(net181));
 sg13g2_dlygate4sd3_1 hold67 (.A(\u_toplayer.reg_layer1[9] ),
    .X(net182));
 sg13g2_dlygate4sd3_1 hold68 (.A(\u_toplayer.reg_layer1[159] ),
    .X(net183));
 sg13g2_dlygate4sd3_1 hold69 (.A(\u_toplayer.reg_layer1[168] ),
    .X(net184));
 sg13g2_dlygate4sd3_1 hold70 (.A(\u_toplayer.reg_layer2[90] ),
    .X(net185));
 sg13g2_dlygate4sd3_1 hold71 (.A(\u_toplayer.reg_layer1[27] ),
    .X(net186));
 sg13g2_dlygate4sd3_1 hold72 (.A(\u_toplayer.outreg[27] ),
    .X(net187));
 sg13g2_dlygate4sd3_1 hold73 (.A(\u_toplayer.reg_layer2[47] ),
    .X(net188));
 sg13g2_dlygate4sd3_1 hold74 (.A(_00442_),
    .X(net189));
 sg13g2_dlygate4sd3_1 hold75 (.A(\u_toplayer.outreg[23] ),
    .X(net190));
 sg13g2_dlygate4sd3_1 hold76 (.A(\u_toplayer.reg_layer2[185] ),
    .X(net191));
 sg13g2_dlygate4sd3_1 hold77 (.A(\u_toplayer.outreg[22] ),
    .X(net192));
 sg13g2_dlygate4sd3_1 hold78 (.A(\u_toplayer.reg_layer1[156] ),
    .X(net193));
 sg13g2_dlygate4sd3_1 hold79 (.A(\u_toplayer.reg_layer2[59] ),
    .X(net194));
 sg13g2_dlygate4sd3_1 hold80 (.A(\u_toplayer.outreg[41] ),
    .X(net195));
 sg13g2_dlygate4sd3_1 hold81 (.A(\u_toplayer.outreg[77] ),
    .X(net196));
 sg13g2_dlygate4sd3_1 hold82 (.A(\u_toplayer.reg_layer1[157] ),
    .X(net197));
 sg13g2_dlygate4sd3_1 hold83 (.A(\u_toplayer.reg_layer1[123] ),
    .X(net198));
 sg13g2_dlygate4sd3_1 hold84 (.A(\u_toplayer.reg_layer1[89] ),
    .X(net199));
 sg13g2_dlygate4sd3_1 hold85 (.A(\u_toplayer.reg_layer1[40] ),
    .X(net200));
 sg13g2_dlygate4sd3_1 hold86 (.A(\u_toplayer.reg_layer2[89] ),
    .X(net201));
 sg13g2_dlygate4sd3_1 hold87 (.A(\u_toplayer.reg_layer2[91] ),
    .X(net202));
 sg13g2_dlygate4sd3_1 hold88 (.A(\u_toplayer.reg_layer2[184] ),
    .X(net203));
 sg13g2_dlygate4sd3_1 hold89 (.A(\u_toplayer.reg_layer2[202] ),
    .X(net204));
 sg13g2_dlygate4sd3_1 hold90 (.A(_00597_),
    .X(net205));
 sg13g2_dlygate4sd3_1 hold91 (.A(\u_toplayer.reg_layer1[253] ),
    .X(net206));
 sg13g2_dlygate4sd3_1 hold92 (.A(\u_toplayer.reg_layer2[104] ),
    .X(net207));
 sg13g2_dlygate4sd3_1 hold93 (.A(_00499_),
    .X(net208));
 sg13g2_dlygate4sd3_1 hold94 (.A(\u_toplayer.reg_layer1[219] ),
    .X(net209));
 sg13g2_dlygate4sd3_1 hold95 (.A(\u_toplayer.reg_layer2[26] ),
    .X(net210));
 sg13g2_dlygate4sd3_1 hold96 (.A(\u_toplayer.outreg[9] ),
    .X(net211));
 sg13g2_dlygate4sd3_1 hold97 (.A(\u_toplayer.outreg[73] ),
    .X(net212));
 sg13g2_dlygate4sd3_1 hold98 (.A(\u_toplayer.reg_layer1[153] ),
    .X(net213));
 sg13g2_dlygate4sd3_1 hold99 (.A(\u_toplayer.reg_layer2[95] ),
    .X(net214));
 sg13g2_dlygate4sd3_1 hold100 (.A(\u_toplayer.reg_layer1[128] ),
    .X(net215));
 sg13g2_dlygate4sd3_1 hold101 (.A(_05540_),
    .X(net216));
 sg13g2_dlygate4sd3_1 hold102 (.A(\u_toplayer.outreg[46] ),
    .X(net217));
 sg13g2_dlygate4sd3_1 hold103 (.A(_00289_),
    .X(net218));
 sg13g2_dlygate4sd3_1 hold104 (.A(\u_toplayer.reg_layer1[204] ),
    .X(net219));
 sg13g2_dlygate4sd3_1 hold105 (.A(\u_toplayer.reg_layer1[11] ),
    .X(net220));
 sg13g2_dlygate4sd3_1 hold106 (.A(\u_toplayer.reg_layer2[155] ),
    .X(net221));
 sg13g2_dlygate4sd3_1 hold107 (.A(\u_toplayer.reg_layer1[93] ),
    .X(net222));
 sg13g2_dlygate4sd3_1 hold108 (.A(\u_toplayer.reg_layer2[221] ),
    .X(net223));
 sg13g2_dlygate4sd3_1 hold109 (.A(\u_toplayer.outreg[76] ),
    .X(net224));
 sg13g2_dlygate4sd3_1 hold110 (.A(\u_toplayer.reg_layer2[127] ),
    .X(net225));
 sg13g2_dlygate4sd3_1 hold111 (.A(\u_toplayer.reg_layer2[107] ),
    .X(net226));
 sg13g2_dlygate4sd3_1 hold112 (.A(_00502_),
    .X(net227));
 sg13g2_dlygate4sd3_1 hold113 (.A(\u_toplayer.reg_layer2[108] ),
    .X(net228));
 sg13g2_dlygate4sd3_1 hold114 (.A(_00503_),
    .X(net229));
 sg13g2_dlygate4sd3_1 hold115 (.A(\u_toplayer.reg_layer2[126] ),
    .X(net230));
 sg13g2_dlygate4sd3_1 hold116 (.A(\u_toplayer.reg_layer2[50] ),
    .X(net231));
 sg13g2_dlygate4sd3_1 hold117 (.A(_00445_),
    .X(net232));
 sg13g2_dlygate4sd3_1 hold118 (.A(\u_toplayer.reg_layer2[85] ),
    .X(net233));
 sg13g2_dlygate4sd3_1 hold119 (.A(\u_toplayer.reg_layer1[155] ),
    .X(net234));
 sg13g2_dlygate4sd3_1 hold120 (.A(_00864_),
    .X(net235));
 sg13g2_dlygate4sd3_1 hold121 (.A(\u_toplayer.reg_layer2[200] ),
    .X(net236));
 sg13g2_dlygate4sd3_1 hold122 (.A(_00595_),
    .X(net237));
 sg13g2_dlygate4sd3_1 hold123 (.A(\u_toplayer.reg_layer1[129] ),
    .X(net238));
 sg13g2_dlygate4sd3_1 hold124 (.A(_05541_),
    .X(net239));
 sg13g2_dlygate4sd3_1 hold125 (.A(\u_toplayer.outreg[10] ),
    .X(net240));
 sg13g2_dlygate4sd3_1 hold126 (.A(\u_toplayer.reg_layer1[162] ),
    .X(net241));
 sg13g2_dlygate4sd3_1 hold127 (.A(\u_toplayer.reg_layer1[85] ),
    .X(net242));
 sg13g2_dlygate4sd3_1 hold128 (.A(\u_toplayer.reg_layer2[15] ),
    .X(net243));
 sg13g2_dlygate4sd3_1 hold129 (.A(\u_toplayer.reg_layer2[13] ),
    .X(net244));
 sg13g2_dlygate4sd3_1 hold130 (.A(\u_toplayer.reg_layer1[114] ),
    .X(net245));
 sg13g2_dlygate4sd3_1 hold131 (.A(_00823_),
    .X(net246));
 sg13g2_dlygate4sd3_1 hold132 (.A(\u_toplayer.reg_layer2[178] ),
    .X(net247));
 sg13g2_dlygate4sd3_1 hold133 (.A(_00573_),
    .X(net248));
 sg13g2_dlygate4sd3_1 hold134 (.A(\u_toplayer.outreg[15] ),
    .X(net249));
 sg13g2_dlygate4sd3_1 hold135 (.A(\u_toplayer.reg_layer2[93] ),
    .X(net250));
 sg13g2_dlygate4sd3_1 hold136 (.A(\u_toplayer.reg_layer2[119] ),
    .X(net251));
 sg13g2_dlygate4sd3_1 hold137 (.A(\u_toplayer.outreg[30] ),
    .X(net252));
 sg13g2_dlygate4sd3_1 hold138 (.A(\u_toplayer.reg_layer1[211] ),
    .X(net253));
 sg13g2_dlygate4sd3_1 hold139 (.A(\u_toplayer.reg_layer1[133] ),
    .X(net254));
 sg13g2_dlygate4sd3_1 hold140 (.A(_05545_),
    .X(net255));
 sg13g2_dlygate4sd3_1 hold141 (.A(\u_toplayer.reg_layer2[125] ),
    .X(net256));
 sg13g2_dlygate4sd3_1 hold142 (.A(\u_toplayer.reg_layer2[189] ),
    .X(net257));
 sg13g2_dlygate4sd3_1 hold143 (.A(\u_toplayer.reg_layer1[250] ),
    .X(net258));
 sg13g2_dlygate4sd3_1 hold144 (.A(\u_toplayer.reg_layer1[124] ),
    .X(net259));
 sg13g2_dlygate4sd3_1 hold145 (.A(\u_toplayer.reg_layer2[94] ),
    .X(net260));
 sg13g2_dlygate4sd3_1 hold146 (.A(\u_toplayer.outreg[2] ),
    .X(net261));
 sg13g2_dlygate4sd3_1 hold147 (.A(\u_toplayer.reg_layer1[10] ),
    .X(net262));
 sg13g2_dlygate4sd3_1 hold148 (.A(_00719_),
    .X(net263));
 sg13g2_dlygate4sd3_1 hold149 (.A(\u_toplayer.reg_layer1[49] ),
    .X(net264));
 sg13g2_dlygate4sd3_1 hold150 (.A(\u_toplayer.reg_layer1[131] ),
    .X(net265));
 sg13g2_dlygate4sd3_1 hold151 (.A(\u_toplayer.reg_layer2[250] ),
    .X(net266));
 sg13g2_dlygate4sd3_1 hold152 (.A(\u_toplayer.reg_layer2[118] ),
    .X(net267));
 sg13g2_dlygate4sd3_1 hold153 (.A(\u_toplayer.reg_layer2[217] ),
    .X(net268));
 sg13g2_dlygate4sd3_1 hold154 (.A(\u_toplayer.reg_layer2[61] ),
    .X(net269));
 sg13g2_dlygate4sd3_1 hold155 (.A(\u_toplayer.reg_layer1[179] ),
    .X(net270));
 sg13g2_dlygate4sd3_1 hold156 (.A(\u_toplayer.reg_layer2[116] ),
    .X(net271));
 sg13g2_dlygate4sd3_1 hold157 (.A(\u_toplayer.reg_layer1[252] ),
    .X(net272));
 sg13g2_dlygate4sd3_1 hold158 (.A(\u_toplayer.reg_layer2[123] ),
    .X(net273));
 sg13g2_dlygate4sd3_1 hold159 (.A(\u_toplayer.reg_layer1[51] ),
    .X(net274));
 sg13g2_dlygate4sd3_1 hold160 (.A(\u_toplayer.reg_layer2[82] ),
    .X(net275));
 sg13g2_dlygate4sd3_1 hold161 (.A(\u_toplayer.reg_layer1[126] ),
    .X(net276));
 sg13g2_dlygate4sd3_1 hold162 (.A(\u_toplayer.reg_layer2[187] ),
    .X(net277));
 sg13g2_dlygate4sd3_1 hold163 (.A(\u_toplayer.reg_layer1[111] ),
    .X(net278));
 sg13g2_dlygate4sd3_1 hold164 (.A(_00820_),
    .X(net279));
 sg13g2_dlygate4sd3_1 hold165 (.A(\u_toplayer.reg_layer1[32] ),
    .X(net280));
 sg13g2_dlygate4sd3_1 hold166 (.A(\u_toplayer.outreg[5] ),
    .X(net281));
 sg13g2_dlygate4sd3_1 hold167 (.A(\u_toplayer.reg_layer2[44] ),
    .X(net282));
 sg13g2_dlygate4sd3_1 hold168 (.A(\u_toplayer.reg_layer1[187] ),
    .X(net283));
 sg13g2_dlygate4sd3_1 hold169 (.A(\u_toplayer.reg_layer1[189] ),
    .X(net284));
 sg13g2_dlygate4sd3_1 hold170 (.A(\u_toplayer.reg_layer1[150] ),
    .X(net285));
 sg13g2_dlygate4sd3_1 hold171 (.A(\u_toplayer.reg_layer1[13] ),
    .X(net286));
 sg13g2_dlygate4sd3_1 hold172 (.A(_00722_),
    .X(net287));
 sg13g2_dlygate4sd3_1 hold173 (.A(\u_toplayer.reg_layer1[173] ),
    .X(net288));
 sg13g2_dlygate4sd3_1 hold174 (.A(\u_toplayer.reg_layer1[14] ),
    .X(net289));
 sg13g2_dlygate4sd3_1 hold175 (.A(\u_toplayer.reg_layer2[247] ),
    .X(net290));
 sg13g2_dlygate4sd3_1 hold176 (.A(\u_toplayer.reg_layer1[30] ),
    .X(net291));
 sg13g2_dlygate4sd3_1 hold177 (.A(\u_toplayer.reg_layer1[199] ),
    .X(net292));
 sg13g2_dlygate4sd3_1 hold178 (.A(_00908_),
    .X(net293));
 sg13g2_dlygate4sd3_1 hold179 (.A(\u_toplayer.reg_layer2[115] ),
    .X(net294));
 sg13g2_dlygate4sd3_1 hold180 (.A(\u_toplayer.reg_layer2[111] ),
    .X(net295));
 sg13g2_dlygate4sd3_1 hold181 (.A(\u_toplayer.reg_layer1[28] ),
    .X(net296));
 sg13g2_dlygate4sd3_1 hold182 (.A(\u_toplayer.reg_layer1[76] ),
    .X(net297));
 sg13g2_dlygate4sd3_1 hold183 (.A(\u_toplayer.reg_layer1[102] ),
    .X(net298));
 sg13g2_dlygate4sd3_1 hold184 (.A(_00811_),
    .X(net299));
 sg13g2_dlygate4sd3_1 hold185 (.A(\u_toplayer.reg_layer2[238] ),
    .X(net300));
 sg13g2_dlygate4sd3_1 hold186 (.A(\u_toplayer.reg_layer2[210] ),
    .X(net301));
 sg13g2_dlygate4sd3_1 hold187 (.A(\u_toplayer.reg_layer2[236] ),
    .X(net302));
 sg13g2_dlygate4sd3_1 hold188 (.A(_00631_),
    .X(net303));
 sg13g2_dlygate4sd3_1 hold189 (.A(\u_toplayer.reg_layer2[117] ),
    .X(net304));
 sg13g2_dlygate4sd3_1 hold190 (.A(\u_toplayer.reg_layer1[224] ),
    .X(net305));
 sg13g2_dlygate4sd3_1 hold191 (.A(_00933_),
    .X(net306));
 sg13g2_dlygate4sd3_1 hold192 (.A(\u_toplayer.reg_layer1[248] ),
    .X(net307));
 sg13g2_dlygate4sd3_1 hold193 (.A(\u_toplayer.reg_layer1[246] ),
    .X(net308));
 sg13g2_dlygate4sd3_1 hold194 (.A(\u_toplayer.reg_layer2[241] ),
    .X(net309));
 sg13g2_dlygate4sd3_1 hold195 (.A(\u_toplayer.reg_layer2[164] ),
    .X(net310));
 sg13g2_dlygate4sd3_1 hold196 (.A(\u_toplayer.reg_layer1[103] ),
    .X(net311));
 sg13g2_dlygate4sd3_1 hold197 (.A(_00812_),
    .X(net312));
 sg13g2_dlygate4sd3_1 hold198 (.A(\u_toplayer.reg_layer1[184] ),
    .X(net313));
 sg13g2_dlygate4sd3_1 hold199 (.A(\u_toplayer.reg_layer2[165] ),
    .X(net314));
 sg13g2_dlygate4sd3_1 hold200 (.A(_00560_),
    .X(net315));
 sg13g2_dlygate4sd3_1 hold201 (.A(\u_toplayer.reg_layer2[198] ),
    .X(net316));
 sg13g2_dlygate4sd3_1 hold202 (.A(\u_toplayer.reg_layer2[80] ),
    .X(net317));
 sg13g2_dlygate4sd3_1 hold203 (.A(\u_toplayer.reg_layer2[206] ),
    .X(net318));
 sg13g2_dlygate4sd3_1 hold204 (.A(_00601_),
    .X(net319));
 sg13g2_dlygate4sd3_1 hold205 (.A(\u_toplayer.reg_layer1[52] ),
    .X(net320));
 sg13g2_dlygate4sd3_1 hold206 (.A(\u_toplayer.reg_layer1[230] ),
    .X(net321));
 sg13g2_dlygate4sd3_1 hold207 (.A(_00939_),
    .X(net322));
 sg13g2_dlygate4sd3_1 hold208 (.A(\u_toplayer.reg_layer2[239] ),
    .X(net323));
 sg13g2_dlygate4sd3_1 hold209 (.A(\u_toplayer.reg_layer2[252] ),
    .X(net324));
 sg13g2_dlygate4sd3_1 hold210 (.A(\u_toplayer.reg_layer1[35] ),
    .X(net325));
 sg13g2_dlygate4sd3_1 hold211 (.A(\u_toplayer.reg_layer1[231] ),
    .X(net326));
 sg13g2_dlygate4sd3_1 hold212 (.A(_00940_),
    .X(net327));
 sg13g2_dlygate4sd3_1 hold213 (.A(\u_toplayer.reg_layer1[66] ),
    .X(net328));
 sg13g2_dlygate4sd3_1 hold214 (.A(\u_toplayer.reg_layer1[163] ),
    .X(net329));
 sg13g2_dlygate4sd3_1 hold215 (.A(\u_toplayer.reg_layer1[228] ),
    .X(net330));
 sg13g2_dlygate4sd3_1 hold216 (.A(\u_toplayer.reg_layer1[167] ),
    .X(net331));
 sg13g2_dlygate4sd3_1 hold217 (.A(\u_toplayer.reg_layer2[226] ),
    .X(net332));
 sg13g2_dlygate4sd3_1 hold218 (.A(\u_toplayer.reg_layer1[182] ),
    .X(net333));
 sg13g2_dlygate4sd3_1 hold219 (.A(\u_toplayer.reg_layer2[128] ),
    .X(net334));
 sg13g2_dlygate4sd3_1 hold220 (.A(\u_toplayer.reg_layer1[180] ),
    .X(net335));
 sg13g2_dlygate4sd3_1 hold221 (.A(\u_toplayer.reg_layer2[166] ),
    .X(net336));
 sg13g2_dlygate4sd3_1 hold222 (.A(_00561_),
    .X(net337));
 sg13g2_dlygate4sd3_1 hold223 (.A(\u_toplayer.reg_layer2[87] ),
    .X(net338));
 sg13g2_dlygate4sd3_1 hold224 (.A(\u_toplayer.reg_layer2[78] ),
    .X(net339));
 sg13g2_dlygate4sd3_1 hold225 (.A(_00473_),
    .X(net340));
 sg13g2_dlygate4sd3_1 hold226 (.A(\u_toplayer.reg_layer1[15] ),
    .X(net341));
 sg13g2_dlygate4sd3_1 hold227 (.A(\u_toplayer.reg_layer1[36] ),
    .X(net342));
 sg13g2_dlygate4sd3_1 hold228 (.A(\u_toplayer.reg_layer2[84] ),
    .X(net343));
 sg13g2_dlygate4sd3_1 hold229 (.A(\u_toplayer.reg_layer2[245] ),
    .X(net344));
 sg13g2_dlygate4sd3_1 hold230 (.A(\u_toplayer.reg_layer1[94] ),
    .X(net345));
 sg13g2_dlygate4sd3_1 hold231 (.A(\u_toplayer.outreg[75] ),
    .X(net346));
 sg13g2_dlygate4sd3_1 hold232 (.A(\u_toplayer.reg_layer2[100] ),
    .X(net347));
 sg13g2_dlygate4sd3_1 hold233 (.A(\u_toplayer.reg_layer1[183] ),
    .X(net348));
 sg13g2_dlygate4sd3_1 hold234 (.A(\u_toplayer.reg_layer2[17] ),
    .X(net349));
 sg13g2_dlygate4sd3_1 hold235 (.A(\u_toplayer.reg_layer2[212] ),
    .X(net350));
 sg13g2_dlygate4sd3_1 hold236 (.A(\u_toplayer.reg_layer1[72] ),
    .X(net351));
 sg13g2_dlygate4sd3_1 hold237 (.A(_00781_),
    .X(net352));
 sg13g2_dlygate4sd3_1 hold238 (.A(\u_toplayer.reg_layer2[190] ),
    .X(net353));
 sg13g2_dlygate4sd3_1 hold239 (.A(\u_toplayer.reg_layer1[88] ),
    .X(net354));
 sg13g2_dlygate4sd3_1 hold240 (.A(\u_toplayer.reg_layer1[195] ),
    .X(net355));
 sg13g2_dlygate4sd3_1 hold241 (.A(\u_toplayer.reg_layer2[150] ),
    .X(net356));
 sg13g2_dlygate4sd3_1 hold242 (.A(\u_toplayer.reg_layer2[230] ),
    .X(net357));
 sg13g2_dlygate4sd3_1 hold243 (.A(\u_toplayer.reg_layer1[169] ),
    .X(net358));
 sg13g2_dlygate4sd3_1 hold244 (.A(\u_toplayer.reg_layer1[206] ),
    .X(net359));
 sg13g2_dlygate4sd3_1 hold245 (.A(\u_toplayer.reg_layer2[153] ),
    .X(net360));
 sg13g2_dlygate4sd3_1 hold246 (.A(\u_toplayer.reg_layer1[226] ),
    .X(net361));
 sg13g2_dlygate4sd3_1 hold247 (.A(\u_toplayer.reg_layer2[186] ),
    .X(net362));
 sg13g2_dlygate4sd3_1 hold248 (.A(\u_toplayer.reg_layer1[41] ),
    .X(net363));
 sg13g2_dlygate4sd3_1 hold249 (.A(\u_toplayer.reg_layer2[28] ),
    .X(net364));
 sg13g2_dlygate4sd3_1 hold250 (.A(\u_toplayer.reg_layer1[96] ),
    .X(net365));
 sg13g2_dlygate4sd3_1 hold251 (.A(_00805_),
    .X(net366));
 sg13g2_dlygate4sd3_1 hold252 (.A(\u_toplayer.reg_layer1[20] ),
    .X(net367));
 sg13g2_dlygate4sd3_1 hold253 (.A(\u_toplayer.reg_layer2[138] ),
    .X(net368));
 sg13g2_dlygate4sd3_1 hold254 (.A(\u_toplayer.reg_layer1[254] ),
    .X(net369));
 sg13g2_dlygate4sd3_1 hold255 (.A(\u_toplayer.reg_layer1[239] ),
    .X(net370));
 sg13g2_dlygate4sd3_1 hold256 (.A(_00948_),
    .X(net371));
 sg13g2_dlygate4sd3_1 hold257 (.A(\u_toplayer.reg_layer2[146] ),
    .X(net372));
 sg13g2_dlygate4sd3_1 hold258 (.A(\u_toplayer.reg_layer1[127] ),
    .X(net373));
 sg13g2_dlygate4sd3_1 hold259 (.A(\u_toplayer.reg_layer1[101] ),
    .X(net374));
 sg13g2_dlygate4sd3_1 hold260 (.A(\u_toplayer.reg_layer1[181] ),
    .X(net375));
 sg13g2_dlygate4sd3_1 hold261 (.A(\u_toplayer.reg_layer1[69] ),
    .X(net376));
 sg13g2_dlygate4sd3_1 hold262 (.A(_00778_),
    .X(net377));
 sg13g2_dlygate4sd3_1 hold263 (.A(\u_toplayer.reg_layer1[24] ),
    .X(net378));
 sg13g2_dlygate4sd3_1 hold264 (.A(\u_toplayer.reg_layer1[109] ),
    .X(net379));
 sg13g2_dlygate4sd3_1 hold265 (.A(\u_toplayer.outreg[26] ),
    .X(net380));
 sg13g2_dlygate4sd3_1 hold266 (.A(\u_toplayer.reg_layer2[96] ),
    .X(net381));
 sg13g2_dlygate4sd3_1 hold267 (.A(_00491_),
    .X(net382));
 sg13g2_dlygate4sd3_1 hold268 (.A(\u_toplayer.reg_layer2[9] ),
    .X(net383));
 sg13g2_dlygate4sd3_1 hold269 (.A(\u_toplayer.reg_layer2[220] ),
    .X(net384));
 sg13g2_dlygate4sd3_1 hold270 (.A(\u_toplayer.reg_layer1[130] ),
    .X(net385));
 sg13g2_dlygate4sd3_1 hold271 (.A(_05542_),
    .X(net386));
 sg13g2_dlygate4sd3_1 hold272 (.A(\u_toplayer.reg_layer2[99] ),
    .X(net387));
 sg13g2_dlygate4sd3_1 hold273 (.A(\u_toplayer.outreg[78] ),
    .X(net388));
 sg13g2_dlygate4sd3_1 hold274 (.A(_00321_),
    .X(net389));
 sg13g2_dlygate4sd3_1 hold275 (.A(\u_toplayer.reg_layer2[114] ),
    .X(net390));
 sg13g2_dlygate4sd3_1 hold276 (.A(\u_toplayer.reg_layer2[216] ),
    .X(net391));
 sg13g2_dlygate4sd3_1 hold277 (.A(\u_toplayer.reg_layer1[25] ),
    .X(net392));
 sg13g2_dlygate4sd3_1 hold278 (.A(\u_toplayer.reg_layer2[205] ),
    .X(net393));
 sg13g2_dlygate4sd3_1 hold279 (.A(_00600_),
    .X(net394));
 sg13g2_dlygate4sd3_1 hold280 (.A(\u_toplayer.outreg[1] ),
    .X(net395));
 sg13g2_dlygate4sd3_1 hold281 (.A(\u_toplayer.reg_layer2[103] ),
    .X(net396));
 sg13g2_dlygate4sd3_1 hold282 (.A(\u_toplayer.reg_layer2[97] ),
    .X(net397));
 sg13g2_dlygate4sd3_1 hold283 (.A(_00492_),
    .X(net398));
 sg13g2_dlygate4sd3_1 hold284 (.A(\u_toplayer.reg_layer2[66] ),
    .X(net399));
 sg13g2_dlygate4sd3_1 hold285 (.A(\u_toplayer.reg_layer1[229] ),
    .X(net400));
 sg13g2_dlygate4sd3_1 hold286 (.A(\u_toplayer.reg_layer1[243] ),
    .X(net401));
 sg13g2_dlygate4sd3_1 hold287 (.A(_00952_),
    .X(net402));
 sg13g2_dlygate4sd3_1 hold288 (.A(\u_toplayer.reg_layer2[253] ),
    .X(net403));
 sg13g2_dlygate4sd3_1 hold289 (.A(\u_toplayer.reg_layer2[63] ),
    .X(net404));
 sg13g2_dlygate4sd3_1 hold290 (.A(\u_toplayer.reg_layer2[188] ),
    .X(net405));
 sg13g2_dlygate4sd3_1 hold291 (.A(\u_toplayer.reg_layer1[148] ),
    .X(net406));
 sg13g2_dlygate4sd3_1 hold292 (.A(\u_toplayer.reg_layer2[135] ),
    .X(net407));
 sg13g2_dlygate4sd3_1 hold293 (.A(\u_toplayer.reg_layer1[55] ),
    .X(net408));
 sg13g2_dlygate4sd3_1 hold294 (.A(\u_toplayer.reg_layer2[20] ),
    .X(net409));
 sg13g2_dlygate4sd3_1 hold295 (.A(\u_toplayer.reg_layer2[183] ),
    .X(net410));
 sg13g2_dlygate4sd3_1 hold296 (.A(\u_toplayer.reg_layer2[223] ),
    .X(net411));
 sg13g2_dlygate4sd3_1 hold297 (.A(\u_toplayer.reg_layer2[18] ),
    .X(net412));
 sg13g2_dlygate4sd3_1 hold298 (.A(\u_toplayer.reg_layer1[249] ),
    .X(net413));
 sg13g2_dlygate4sd3_1 hold299 (.A(_00958_),
    .X(net414));
 sg13g2_dlygate4sd3_1 hold300 (.A(\u_toplayer.reg_layer1[58] ),
    .X(net415));
 sg13g2_dlygate4sd3_1 hold301 (.A(\u_toplayer.reg_layer1[113] ),
    .X(net416));
 sg13g2_dlygate4sd3_1 hold302 (.A(_00822_),
    .X(net417));
 sg13g2_dlygate4sd3_1 hold303 (.A(\u_toplayer.reg_layer1[97] ),
    .X(net418));
 sg13g2_dlygate4sd3_1 hold304 (.A(\u_toplayer.reg_layer1[158] ),
    .X(net419));
 sg13g2_dlygate4sd3_1 hold305 (.A(\u_toplayer.reg_layer2[21] ),
    .X(net420));
 sg13g2_dlygate4sd3_1 hold306 (.A(\u_toplayer.reg_layer1[234] ),
    .X(net421));
 sg13g2_dlygate4sd3_1 hold307 (.A(_00943_),
    .X(net422));
 sg13g2_dlygate4sd3_1 hold308 (.A(\u_toplayer.reg_layer1[115] ),
    .X(net423));
 sg13g2_dlygate4sd3_1 hold309 (.A(_00824_),
    .X(net424));
 sg13g2_dlygate4sd3_1 hold310 (.A(\u_toplayer.reg_layer1[84] ),
    .X(net425));
 sg13g2_dlygate4sd3_1 hold311 (.A(\u_toplayer.outreg[16] ),
    .X(net426));
 sg13g2_dlygate4sd3_1 hold312 (.A(\u_toplayer.reg_layer1[160] ),
    .X(net427));
 sg13g2_dlygate4sd3_1 hold313 (.A(\u_toplayer.reg_layer2[106] ),
    .X(net428));
 sg13g2_dlygate4sd3_1 hold314 (.A(\u_toplayer.reg_layer2[70] ),
    .X(net429));
 sg13g2_dlygate4sd3_1 hold315 (.A(\u_toplayer.reg_layer2[251] ),
    .X(net430));
 sg13g2_dlygate4sd3_1 hold316 (.A(\u_toplayer.reg_layer1[202] ),
    .X(net431));
 sg13g2_dlygate4sd3_1 hold317 (.A(\u_toplayer.reg_layer1[65] ),
    .X(net432));
 sg13g2_dlygate4sd3_1 hold318 (.A(\u_toplayer.reg_layer2[62] ),
    .X(net433));
 sg13g2_dlygate4sd3_1 hold319 (.A(\u_toplayer.reg_layer2[193] ),
    .X(net434));
 sg13g2_dlygate4sd3_1 hold320 (.A(\u_toplayer.reg_layer2[162] ),
    .X(net435));
 sg13g2_dlygate4sd3_1 hold321 (.A(_00557_),
    .X(net436));
 sg13g2_dlygate4sd3_1 hold322 (.A(\u_toplayer.reg_layer2[68] ),
    .X(net437));
 sg13g2_dlygate4sd3_1 hold323 (.A(\u_toplayer.reg_layer2[72] ),
    .X(net438));
 sg13g2_dlygate4sd3_1 hold324 (.A(_00467_),
    .X(net439));
 sg13g2_dlygate4sd3_1 hold325 (.A(\u_toplayer.reg_layer2[235] ),
    .X(net440));
 sg13g2_dlygate4sd3_1 hold326 (.A(_00630_),
    .X(net441));
 sg13g2_dlygate4sd3_1 hold327 (.A(\u_toplayer.reg_layer1[80] ),
    .X(net442));
 sg13g2_dlygate4sd3_1 hold328 (.A(\u_toplayer.reg_layer2[69] ),
    .X(net443));
 sg13g2_dlygate4sd3_1 hold329 (.A(\u_toplayer.reg_layer2[201] ),
    .X(net444));
 sg13g2_dlygate4sd3_1 hold330 (.A(_00596_),
    .X(net445));
 sg13g2_dlygate4sd3_1 hold331 (.A(\u_toplayer.reg_layer1[215] ),
    .X(net446));
 sg13g2_dlygate4sd3_1 hold332 (.A(_00924_),
    .X(net447));
 sg13g2_dlygate4sd3_1 hold333 (.A(\u_toplayer.reg_layer1[196] ),
    .X(net448));
 sg13g2_dlygate4sd3_1 hold334 (.A(\u_toplayer.reg_layer1[151] ),
    .X(net449));
 sg13g2_dlygate4sd3_1 hold335 (.A(\u_toplayer.reg_layer1[34] ),
    .X(net450));
 sg13g2_dlygate4sd3_1 hold336 (.A(\u_toplayer.reg_layer1[73] ),
    .X(net451));
 sg13g2_dlygate4sd3_1 hold337 (.A(_00782_),
    .X(net452));
 sg13g2_dlygate4sd3_1 hold338 (.A(\u_toplayer.reg_layer2[45] ),
    .X(net453));
 sg13g2_dlygate4sd3_1 hold339 (.A(_00440_),
    .X(net454));
 sg13g2_dlygate4sd3_1 hold340 (.A(\u_toplayer.reg_layer2[43] ),
    .X(net455));
 sg13g2_dlygate4sd3_1 hold341 (.A(_00438_),
    .X(net456));
 sg13g2_dlygate4sd3_1 hold342 (.A(\u_toplayer.reg_layer1[222] ),
    .X(net457));
 sg13g2_dlygate4sd3_1 hold343 (.A(\u_toplayer.reg_layer1[227] ),
    .X(net458));
 sg13g2_dlygate4sd3_1 hold344 (.A(\u_toplayer.reg_layer2[246] ),
    .X(net459));
 sg13g2_dlygate4sd3_1 hold345 (.A(\u_toplayer.reg_layer1[91] ),
    .X(net460));
 sg13g2_dlygate4sd3_1 hold346 (.A(\u_toplayer.reg_layer2[40] ),
    .X(net461));
 sg13g2_dlygate4sd3_1 hold347 (.A(\u_toplayer.reg_layer1[59] ),
    .X(net462));
 sg13g2_dlygate4sd3_1 hold348 (.A(\u_toplayer.reg_layer1[119] ),
    .X(net463));
 sg13g2_dlygate4sd3_1 hold349 (.A(_00828_),
    .X(net464));
 sg13g2_dlygate4sd3_1 hold350 (.A(\u_toplayer.reg_layer2[76] ),
    .X(net465));
 sg13g2_dlygate4sd3_1 hold351 (.A(\u_toplayer.reg_layer1[12] ),
    .X(net466));
 sg13g2_dlygate4sd3_1 hold352 (.A(\u_toplayer.reg_layer1[18] ),
    .X(net467));
 sg13g2_dlygate4sd3_1 hold353 (.A(\u_toplayer.reg_layer1[235] ),
    .X(net468));
 sg13g2_dlygate4sd3_1 hold354 (.A(_00944_),
    .X(net469));
 sg13g2_dlygate4sd3_1 hold355 (.A(\u_toplayer.reg_layer2[254] ),
    .X(net470));
 sg13g2_dlygate4sd3_1 hold356 (.A(\u_toplayer.reg_layer2[110] ),
    .X(net471));
 sg13g2_dlygate4sd3_1 hold357 (.A(\u_toplayer.reg_layer2[145] ),
    .X(net472));
 sg13g2_dlygate4sd3_1 hold358 (.A(\u_toplayer.reg_layer1[171] ),
    .X(net473));
 sg13g2_dlygate4sd3_1 hold359 (.A(\u_toplayer.reg_layer1[191] ),
    .X(net474));
 sg13g2_dlygate4sd3_1 hold360 (.A(\u_toplayer.reg_layer2[249] ),
    .X(net475));
 sg13g2_dlygate4sd3_1 hold361 (.A(\u_toplayer.reg_layer1[241] ),
    .X(net476));
 sg13g2_dlygate4sd3_1 hold362 (.A(_00950_),
    .X(net477));
 sg13g2_dlygate4sd3_1 hold363 (.A(\u_toplayer.reg_layer1[212] ),
    .X(net478));
 sg13g2_dlygate4sd3_1 hold364 (.A(\u_toplayer.reg_layer2[233] ),
    .X(net479));
 sg13g2_dlygate4sd3_1 hold365 (.A(\u_toplayer.reg_layer2[25] ),
    .X(net480));
 sg13g2_dlygate4sd3_1 hold366 (.A(_00420_),
    .X(net481));
 sg13g2_dlygate4sd3_1 hold367 (.A(\u_toplayer.reg_layer1[61] ),
    .X(net482));
 sg13g2_dlygate4sd3_1 hold368 (.A(\u_toplayer.reg_layer2[105] ),
    .X(net483));
 sg13g2_dlygate4sd3_1 hold369 (.A(\u_toplayer.reg_layer2[174] ),
    .X(net484));
 sg13g2_dlygate4sd3_1 hold370 (.A(_00569_),
    .X(net485));
 sg13g2_dlygate4sd3_1 hold371 (.A(\u_toplayer.reg_layer2[10] ),
    .X(net486));
 sg13g2_dlygate4sd3_1 hold372 (.A(\u_toplayer.reg_layer2[213] ),
    .X(net487));
 sg13g2_dlygate4sd3_1 hold373 (.A(\u_toplayer.reg_layer1[165] ),
    .X(net488));
 sg13g2_dlygate4sd3_1 hold374 (.A(\u_toplayer.reg_layer2[24] ),
    .X(net489));
 sg13g2_dlygate4sd3_1 hold375 (.A(\u_toplayer.reg_layer1[200] ),
    .X(net490));
 sg13g2_dlygate4sd3_1 hold376 (.A(_00909_),
    .X(net491));
 sg13g2_dlygate4sd3_1 hold377 (.A(\u_toplayer.reg_layer1[236] ),
    .X(net492));
 sg13g2_dlygate4sd3_1 hold378 (.A(_00945_),
    .X(net493));
 sg13g2_dlygate4sd3_1 hold379 (.A(\u_toplayer.reg_layer2[11] ),
    .X(net494));
 sg13g2_dlygate4sd3_1 hold380 (.A(\u_toplayer.reg_layer1[144] ),
    .X(net495));
 sg13g2_dlygate4sd3_1 hold381 (.A(\u_toplayer.reg_layer2[74] ),
    .X(net496));
 sg13g2_dlygate4sd3_1 hold382 (.A(_00469_),
    .X(net497));
 sg13g2_dlygate4sd3_1 hold383 (.A(\u_toplayer.reg_layer1[154] ),
    .X(net498));
 sg13g2_dlygate4sd3_1 hold384 (.A(\u_toplayer.reg_layer1[33] ),
    .X(net499));
 sg13g2_dlygate4sd3_1 hold385 (.A(\u_toplayer.reg_layer1[245] ),
    .X(net500));
 sg13g2_dlygate4sd3_1 hold386 (.A(_00954_),
    .X(net501));
 sg13g2_dlygate4sd3_1 hold387 (.A(\u_toplayer.reg_layer1[78] ),
    .X(net502));
 sg13g2_dlygate4sd3_1 hold388 (.A(\u_toplayer.reg_layer2[197] ),
    .X(net503));
 sg13g2_dlygate4sd3_1 hold389 (.A(\u_toplayer.outreg[7] ),
    .X(net504));
 sg13g2_dlygate4sd3_1 hold390 (.A(\u_toplayer.reg_layer1[198] ),
    .X(net505));
 sg13g2_dlygate4sd3_1 hold391 (.A(\u_toplayer.reg_layer2[113] ),
    .X(net506));
 sg13g2_dlygate4sd3_1 hold392 (.A(\u_toplayer.reg_layer2[173] ),
    .X(net507));
 sg13g2_dlygate4sd3_1 hold393 (.A(_00568_),
    .X(net508));
 sg13g2_dlygate4sd3_1 hold394 (.A(\u_toplayer.reg_layer2[224] ),
    .X(net509));
 sg13g2_dlygate4sd3_1 hold395 (.A(_00619_),
    .X(net510));
 sg13g2_dlygate4sd3_1 hold396 (.A(\u_toplayer.u_layer1.u_neuron.instCtrl.state[4] ),
    .X(net511));
 sg13g2_dlygate4sd3_1 hold397 (.A(_00004_),
    .X(net512));
 sg13g2_dlygate4sd3_1 hold398 (.A(\u_toplayer.reg_layer1[176] ),
    .X(net513));
 sg13g2_dlygate4sd3_1 hold399 (.A(\u_toplayer.reg_layer1[71] ),
    .X(net514));
 sg13g2_dlygate4sd3_1 hold400 (.A(_00780_),
    .X(net515));
 sg13g2_dlygate4sd3_1 hold401 (.A(\u_toplayer.reg_layer1[194] ),
    .X(net516));
 sg13g2_dlygate4sd3_1 hold402 (.A(\u_toplayer.reg_layer1[132] ),
    .X(net517));
 sg13g2_dlygate4sd3_1 hold403 (.A(_00841_),
    .X(net518));
 sg13g2_dlygate4sd3_1 hold404 (.A(\u_toplayer.reg_layer1[82] ),
    .X(net519));
 sg13g2_dlygate4sd3_1 hold405 (.A(\u_toplayer.reg_layer2[231] ),
    .X(net520));
 sg13g2_dlygate4sd3_1 hold406 (.A(\u_toplayer.reg_layer1[193] ),
    .X(net521));
 sg13g2_dlygate4sd3_1 hold407 (.A(\u_toplayer.reg_layer2[229] ),
    .X(net522));
 sg13g2_dlygate4sd3_1 hold408 (.A(\u_toplayer.reg_layer2[137] ),
    .X(net523));
 sg13g2_dlygate4sd3_1 hold409 (.A(\u_toplayer.reg_layer2[48] ),
    .X(net524));
 sg13g2_dlygate4sd3_1 hold410 (.A(_00443_),
    .X(net525));
 sg13g2_dlygate4sd3_1 hold411 (.A(\u_toplayer.reg_layer2[37] ),
    .X(net526));
 sg13g2_dlygate4sd3_1 hold412 (.A(_00432_),
    .X(net527));
 sg13g2_dlygate4sd3_1 hold413 (.A(\u_toplayer.reg_layer2[167] ),
    .X(net528));
 sg13g2_dlygate4sd3_1 hold414 (.A(_00562_),
    .X(net529));
 sg13g2_dlygate4sd3_1 hold415 (.A(\u_toplayer.reg_layer1[57] ),
    .X(net530));
 sg13g2_dlygate4sd3_1 hold416 (.A(\u_toplayer.reg_layer1[63] ),
    .X(net531));
 sg13g2_dlygate4sd3_1 hold417 (.A(\u_toplayer.reg_layer2[136] ),
    .X(net532));
 sg13g2_dlygate4sd3_1 hold418 (.A(\u_toplayer.reg_layer2[142] ),
    .X(net533));
 sg13g2_dlygate4sd3_1 hold419 (.A(\u_toplayer.reg_layer1[50] ),
    .X(net534));
 sg13g2_dlygate4sd3_1 hold420 (.A(\u_toplayer.reg_layer2[191] ),
    .X(net535));
 sg13g2_dlygate4sd3_1 hold421 (.A(\u_toplayer.reg_layer2[244] ),
    .X(net536));
 sg13g2_dlygate4sd3_1 hold422 (.A(\u_toplayer.reg_layer2[29] ),
    .X(net537));
 sg13g2_dlygate4sd3_1 hold423 (.A(\u_toplayer.reg_layer2[65] ),
    .X(net538));
 sg13g2_dlygate4sd3_1 hold424 (.A(\u_toplayer.reg_layer1[29] ),
    .X(net539));
 sg13g2_dlygate4sd3_1 hold425 (.A(\u_toplayer.reg_layer1[112] ),
    .X(net540));
 sg13g2_dlygate4sd3_1 hold426 (.A(\u_toplayer.reg_layer1[233] ),
    .X(net541));
 sg13g2_dlygate4sd3_1 hold427 (.A(\u_toplayer.reg_layer1[45] ),
    .X(net542));
 sg13g2_dlygate4sd3_1 hold428 (.A(\u_toplayer.reg_layer1[39] ),
    .X(net543));
 sg13g2_dlygate4sd3_1 hold429 (.A(\u_toplayer.reg_layer1[19] ),
    .X(net544));
 sg13g2_dlygate4sd3_1 hold430 (.A(\u_toplayer.reg_layer1[142] ),
    .X(net545));
 sg13g2_dlygate4sd3_1 hold431 (.A(\u_toplayer.reg_layer1[188] ),
    .X(net546));
 sg13g2_dlygate4sd3_1 hold432 (.A(\u_toplayer.reg_layer2[196] ),
    .X(net547));
 sg13g2_dlygate4sd3_1 hold433 (.A(\u_toplayer.reg_layer1[146] ),
    .X(net548));
 sg13g2_dlygate4sd3_1 hold434 (.A(\u_toplayer.reg_layer1[152] ),
    .X(net549));
 sg13g2_dlygate4sd3_1 hold435 (.A(\u_toplayer.reg_layer2[225] ),
    .X(net550));
 sg13g2_dlygate4sd3_1 hold436 (.A(_00620_),
    .X(net551));
 sg13g2_dlygate4sd3_1 hold437 (.A(\u_toplayer.reg_layer1[117] ),
    .X(net552));
 sg13g2_dlygate4sd3_1 hold438 (.A(_00826_),
    .X(net553));
 sg13g2_dlygate4sd3_1 hold439 (.A(\u_toplayer.u_layer1.u_neuron.instCtrl.state[6] ),
    .X(net554));
 sg13g2_dlygate4sd3_1 hold440 (.A(_00006_),
    .X(net555));
 sg13g2_dlygate4sd3_1 hold441 (.A(\u_toplayer.reg_layer2[75] ),
    .X(net556));
 sg13g2_dlygate4sd3_1 hold442 (.A(\u_toplayer.reg_layer1[166] ),
    .X(net557));
 sg13g2_dlygate4sd3_1 hold443 (.A(\u_toplayer.reg_layer1[81] ),
    .X(net558));
 sg13g2_dlygate4sd3_1 hold444 (.A(\u_toplayer.reg_layer2[60] ),
    .X(net559));
 sg13g2_dlygate4sd3_1 hold445 (.A(\u_toplayer.reg_layer2[141] ),
    .X(net560));
 sg13g2_dlygate4sd3_1 hold446 (.A(\u_toplayer.reg_layer1[98] ),
    .X(net561));
 sg13g2_dlygate4sd3_1 hold447 (.A(\u_toplayer.reg_layer1[22] ),
    .X(net562));
 sg13g2_dlygate4sd3_1 hold448 (.A(\u_toplayer.reg_layer2[199] ),
    .X(net563));
 sg13g2_dlygate4sd3_1 hold449 (.A(\u_toplayer.reg_layer1[21] ),
    .X(net564));
 sg13g2_dlygate4sd3_1 hold450 (.A(\u_toplayer.reg_layer2[53] ),
    .X(net565));
 sg13g2_dlygate4sd3_1 hold451 (.A(_00448_),
    .X(net566));
 sg13g2_dlygate4sd3_1 hold452 (.A(\u_toplayer.reg_layer1[238] ),
    .X(net567));
 sg13g2_dlygate4sd3_1 hold453 (.A(_00947_),
    .X(net568));
 sg13g2_dlygate4sd3_1 hold454 (.A(\u_toplayer.u_layer1.u_neuron.instCtrl.state[5] ),
    .X(net569));
 sg13g2_dlygate4sd3_1 hold455 (.A(_00005_),
    .X(net570));
 sg13g2_dlygate4sd3_1 hold456 (.A(\u_toplayer.reg_layer1[79] ),
    .X(net571));
 sg13g2_dlygate4sd3_1 hold457 (.A(_00788_),
    .X(net572));
 sg13g2_dlygate4sd3_1 hold458 (.A(\u_toplayer.reg_layer1[87] ),
    .X(net573));
 sg13g2_dlygate4sd3_1 hold459 (.A(_00796_),
    .X(net574));
 sg13g2_dlygate4sd3_1 hold460 (.A(\u_toplayer.reg_layer1[26] ),
    .X(net575));
 sg13g2_dlygate4sd3_1 hold461 (.A(\u_toplayer.reg_layer1[244] ),
    .X(net576));
 sg13g2_dlygate4sd3_1 hold462 (.A(_00953_),
    .X(net577));
 sg13g2_dlygate4sd3_1 hold463 (.A(\u_toplayer.reg_layer2[14] ),
    .X(net578));
 sg13g2_dlygate4sd3_1 hold464 (.A(\u_toplayer.reg_layer2[121] ),
    .X(net579));
 sg13g2_dlygate4sd3_1 hold465 (.A(\u_toplayer.reg_layer2[64] ),
    .X(net580));
 sg13g2_dlygate4sd3_1 hold466 (.A(\u_toplayer.reg_layer1[178] ),
    .X(net581));
 sg13g2_dlygate4sd3_1 hold467 (.A(\u_toplayer.reg_layer1[100] ),
    .X(net582));
 sg13g2_dlygate4sd3_1 hold468 (.A(\u_toplayer.reg_layer2[243] ),
    .X(net583));
 sg13g2_dlygate4sd3_1 hold469 (.A(\u_toplayer.reg_layer1[120] ),
    .X(net584));
 sg13g2_dlygate4sd3_1 hold470 (.A(\u_toplayer.reg_layer2[180] ),
    .X(net585));
 sg13g2_dlygate4sd3_1 hold471 (.A(_00575_),
    .X(net586));
 sg13g2_dlygate4sd3_1 hold472 (.A(\u_toplayer.reg_layer2[27] ),
    .X(net587));
 sg13g2_dlygate4sd3_1 hold473 (.A(\u_toplayer.reg_layer2[101] ),
    .X(net588));
 sg13g2_dlygate4sd3_1 hold474 (.A(\u_toplayer.reg_layer2[242] ),
    .X(net589));
 sg13g2_dlygate4sd3_1 hold475 (.A(\u_toplayer.reg_layer2[57] ),
    .X(net590));
 sg13g2_dlygate4sd3_1 hold476 (.A(\u_toplayer.outreg[3] ),
    .X(net591));
 sg13g2_dlygate4sd3_1 hold477 (.A(\u_toplayer.reg_layer2[22] ),
    .X(net592));
 sg13g2_dlygate4sd3_1 hold478 (.A(\u_toplayer.reg_layer2[159] ),
    .X(net593));
 sg13g2_dlygate4sd3_1 hold479 (.A(\u_toplayer.outreg[28] ),
    .X(net594));
 sg13g2_dlygate4sd3_1 hold480 (.A(\u_toplayer.reg_layer2[179] ),
    .X(net595));
 sg13g2_dlygate4sd3_1 hold481 (.A(\u_toplayer.reg_layer1[218] ),
    .X(net596));
 sg13g2_dlygate4sd3_1 hold482 (.A(_00050_),
    .X(net597));
 sg13g2_dlygate4sd3_1 hold483 (.A(_00701_),
    .X(net598));
 sg13g2_dlygate4sd3_1 hold484 (.A(\u_toplayer.reg_layer1[140] ),
    .X(net599));
 sg13g2_dlygate4sd3_1 hold485 (.A(\u_toplayer.reg_layer2[163] ),
    .X(net600));
 sg13g2_dlygate4sd3_1 hold486 (.A(_00558_),
    .X(net601));
 sg13g2_dlygate4sd3_1 hold487 (.A(\u_toplayer.reg_layer1[42] ),
    .X(net602));
 sg13g2_dlygate4sd3_1 hold488 (.A(\u_toplayer.reg_layer2[32] ),
    .X(net603));
 sg13g2_dlygate4sd3_1 hold489 (.A(\u_toplayer.reg_layer2[156] ),
    .X(net604));
 sg13g2_dlygate4sd3_1 hold490 (.A(\u_toplayer.reg_layer2[19] ),
    .X(net605));
 sg13g2_dlygate4sd3_1 hold491 (.A(\u_toplayer.reg_layer2[83] ),
    .X(net606));
 sg13g2_dlygate4sd3_1 hold492 (.A(\u_toplayer.reg_layer1[31] ),
    .X(net607));
 sg13g2_dlygate4sd3_1 hold493 (.A(\u_toplayer.reg_layer1[60] ),
    .X(net608));
 sg13g2_dlygate4sd3_1 hold494 (.A(\u_toplayer.reg_layer2[36] ),
    .X(net609));
 sg13g2_dlygate4sd3_1 hold495 (.A(\u_toplayer.reg_layer1[48] ),
    .X(net610));
 sg13g2_dlygate4sd3_1 hold496 (.A(\u_toplayer.reg_layer1[125] ),
    .X(net611));
 sg13g2_dlygate4sd3_1 hold497 (.A(\u_toplayer.reg_layer2[56] ),
    .X(net612));
 sg13g2_dlygate4sd3_1 hold498 (.A(\u_toplayer.reg_layer2[55] ),
    .X(net613));
 sg13g2_dlygate4sd3_1 hold499 (.A(\u_toplayer.reg_layer2[147] ),
    .X(net614));
 sg13g2_dlygate4sd3_1 hold500 (.A(\u_toplayer.reg_layer1[237] ),
    .X(net615));
 sg13g2_dlygate4sd3_1 hold501 (.A(\u_toplayer.reg_layer2[33] ),
    .X(net616));
 sg13g2_dlygate4sd3_1 hold502 (.A(\u_toplayer.reg_layer1[90] ),
    .X(net617));
 sg13g2_dlygate4sd3_1 hold503 (.A(\u_toplayer.reg_layer2[237] ),
    .X(net618));
 sg13g2_dlygate4sd3_1 hold504 (.A(\u_toplayer.reg_layer2[112] ),
    .X(net619));
 sg13g2_dlygate4sd3_1 hold505 (.A(\u_toplayer.reg_layer2[131] ),
    .X(net620));
 sg13g2_dlygate4sd3_1 hold506 (.A(\u_toplayer.reg_layer2[175] ),
    .X(net621));
 sg13g2_dlygate4sd3_1 hold507 (.A(_00570_),
    .X(net622));
 sg13g2_dlygate4sd3_1 hold508 (.A(\u_toplayer.reg_layer1[106] ),
    .X(net623));
 sg13g2_dlygate4sd3_1 hold509 (.A(_00815_),
    .X(net624));
 sg13g2_dlygate4sd3_1 hold510 (.A(\u_toplayer.u_layer1.statel1[8] ),
    .X(net625));
 sg13g2_dlygate4sd3_1 hold511 (.A(_00989_),
    .X(net626));
 sg13g2_dlygate4sd3_1 hold512 (.A(\u_toplayer.reg_layer1[177] ),
    .X(net627));
 sg13g2_dlygate4sd3_1 hold513 (.A(\u_toplayer.reg_layer2[52] ),
    .X(net628));
 sg13g2_dlygate4sd3_1 hold514 (.A(_00447_),
    .X(net629));
 sg13g2_dlygate4sd3_1 hold515 (.A(\u_toplayer.reg_layer2[176] ),
    .X(net630));
 sg13g2_dlygate4sd3_1 hold516 (.A(_00571_),
    .X(net631));
 sg13g2_dlygate4sd3_1 hold517 (.A(\u_toplayer.reg_layer2[102] ),
    .X(net632));
 sg13g2_dlygate4sd3_1 hold518 (.A(\u_toplayer.reg_layer1[118] ),
    .X(net633));
 sg13g2_dlygate4sd3_1 hold519 (.A(\u_toplayer.reg_layer1[175] ),
    .X(net634));
 sg13g2_dlygate4sd3_1 hold520 (.A(\u_toplayer.reg_layer2[98] ),
    .X(net635));
 sg13g2_dlygate4sd3_1 hold521 (.A(\u_toplayer.reg_layer2[161] ),
    .X(net636));
 sg13g2_dlygate4sd3_1 hold522 (.A(\u_toplayer.reg_layer2[139] ),
    .X(net637));
 sg13g2_dlygate4sd3_1 hold523 (.A(\u_toplayer.reg_layer2[58] ),
    .X(net638));
 sg13g2_dlygate4sd3_1 hold524 (.A(\u_toplayer.reg_layer1[64] ),
    .X(net639));
 sg13g2_dlygate4sd3_1 hold525 (.A(\u_toplayer.reg_layer1[70] ),
    .X(net640));
 sg13g2_dlygate4sd3_1 hold526 (.A(\u_toplayer.reg_layer2[151] ),
    .X(net641));
 sg13g2_dlygate4sd3_1 hold527 (.A(\u_toplayer.reg_layer2[182] ),
    .X(net642));
 sg13g2_dlygate4sd3_1 hold528 (.A(\u_toplayer.reg_layer2[148] ),
    .X(net643));
 sg13g2_dlygate4sd3_1 hold529 (.A(\u_toplayer.reg_layer2[109] ),
    .X(net644));
 sg13g2_dlygate4sd3_1 hold530 (.A(\u_toplayer.reg_layer1[232] ),
    .X(net645));
 sg13g2_dlygate4sd3_1 hold531 (.A(\u_toplayer.reg_layer1[217] ),
    .X(net646));
 sg13g2_dlygate4sd3_1 hold532 (.A(\u_toplayer.reg_layer2[140] ),
    .X(net647));
 sg13g2_dlygate4sd3_1 hold533 (.A(_00535_),
    .X(net648));
 sg13g2_dlygate4sd3_1 hold534 (.A(\u_toplayer.reg_layer1[145] ),
    .X(net649));
 sg13g2_dlygate4sd3_1 hold535 (.A(\u_toplayer.reg_layer2[209] ),
    .X(net650));
 sg13g2_dlygate4sd3_1 hold536 (.A(\u_toplayer.reg_layer2[49] ),
    .X(net651));
 sg13g2_dlygate4sd3_1 hold537 (.A(_00444_),
    .X(net652));
 sg13g2_dlygate4sd3_1 hold538 (.A(\u_toplayer.reg_layer2[169] ),
    .X(net653));
 sg13g2_dlygate4sd3_1 hold539 (.A(\u_toplayer.reg_layer2[23] ),
    .X(net654));
 sg13g2_dlygate4sd3_1 hold540 (.A(\u_toplayer.reg_layer2[88] ),
    .X(net655));
 sg13g2_dlygate4sd3_1 hold541 (.A(\u_toplayer.reg_layer2[228] ),
    .X(net656));
 sg13g2_dlygate4sd3_1 hold542 (.A(\u_toplayer.reg_layer2[232] ),
    .X(net657));
 sg13g2_dlygate4sd3_1 hold543 (.A(_00627_),
    .X(net658));
 sg13g2_dlygate4sd3_1 hold544 (.A(\u_toplayer.reg_layer1[208] ),
    .X(net659));
 sg13g2_dlygate4sd3_1 hold545 (.A(\u_toplayer.reg_layer2[255] ),
    .X(net660));
 sg13g2_dlygate4sd3_1 hold546 (.A(\u_toplayer.reg_layer2[130] ),
    .X(net661));
 sg13g2_dlygate4sd3_1 hold547 (.A(\u_toplayer.reg_layer2[219] ),
    .X(net662));
 sg13g2_dlygate4sd3_1 hold548 (.A(\u_toplayer.reg_layer2[132] ),
    .X(net663));
 sg13g2_dlygate4sd3_1 hold549 (.A(\u_toplayer.reg_layer2[122] ),
    .X(net664));
 sg13g2_dlygate4sd3_1 hold550 (.A(\u_toplayer.reg_layer2[77] ),
    .X(net665));
 sg13g2_dlygate4sd3_1 hold551 (.A(_00472_),
    .X(net666));
 sg13g2_dlygate4sd3_1 hold552 (.A(\u_toplayer.reg_layer1[137] ),
    .X(net667));
 sg13g2_dlygate4sd3_1 hold553 (.A(\u_toplayer.reg_layer1[8] ),
    .X(net668));
 sg13g2_dlygate4sd3_1 hold554 (.A(\u_toplayer.reg_layer1[135] ),
    .X(net669));
 sg13g2_dlygate4sd3_1 hold555 (.A(_05547_),
    .X(net670));
 sg13g2_dlygate4sd3_1 hold556 (.A(\u_toplayer.reg_layer2[234] ),
    .X(net671));
 sg13g2_dlygate4sd3_1 hold557 (.A(\u_toplayer.reg_layer1[86] ),
    .X(net672));
 sg13g2_dlygate4sd3_1 hold558 (.A(\u_toplayer.reg_layer1[203] ),
    .X(net673));
 sg13g2_dlygate4sd3_1 hold559 (.A(\u_toplayer.reg_layer2[194] ),
    .X(net674));
 sg13g2_dlygate4sd3_1 hold560 (.A(\u_toplayer.reg_layer1[216] ),
    .X(net675));
 sg13g2_dlygate4sd3_1 hold561 (.A(\u_toplayer.reg_layer2[51] ),
    .X(net676));
 sg13g2_dlygate4sd3_1 hold562 (.A(\u_toplayer.reg_layer1[174] ),
    .X(net677));
 sg13g2_dlygate4sd3_1 hold563 (.A(\u_toplayer.reg_layer1[74] ),
    .X(net678));
 sg13g2_dlygate4sd3_1 hold564 (.A(\u_toplayer.reg_layer1[220] ),
    .X(net679));
 sg13g2_dlygate4sd3_1 hold565 (.A(_00929_),
    .X(net680));
 sg13g2_dlygate4sd3_1 hold566 (.A(_00039_),
    .X(net681));
 sg13g2_dlygate4sd3_1 hold567 (.A(_01343_),
    .X(net682));
 sg13g2_dlygate4sd3_1 hold568 (.A(_00024_),
    .X(net683));
 sg13g2_dlygate4sd3_1 hold569 (.A(\u_toplayer.reg_layer2[149] ),
    .X(net684));
 sg13g2_dlygate4sd3_1 hold570 (.A(\u_toplayer.reg_layer2[35] ),
    .X(net685));
 sg13g2_dlygate4sd3_1 hold571 (.A(_00430_),
    .X(net686));
 sg13g2_dlygate4sd3_1 hold572 (.A(\u_toplayer.reg_layer1[197] ),
    .X(net687));
 sg13g2_dlygate4sd3_1 hold573 (.A(\u_toplayer.reg_layer1[107] ),
    .X(net688));
 sg13g2_dlygate4sd3_1 hold574 (.A(_00816_),
    .X(net689));
 sg13g2_dlygate4sd3_1 hold575 (.A(\u_toplayer.reg_layer1[16] ),
    .X(net690));
 sg13g2_dlygate4sd3_1 hold576 (.A(\u_toplayer.reg_layer1[139] ),
    .X(net691));
 sg13g2_dlygate4sd3_1 hold577 (.A(\u_toplayer.reg_layer1[23] ),
    .X(net692));
 sg13g2_dlygate4sd3_1 hold578 (.A(\u_toplayer.reg_layer2[227] ),
    .X(net693));
 sg13g2_dlygate4sd3_1 hold579 (.A(\u_toplayer.reg_layer1[207] ),
    .X(net694));
 sg13g2_dlygate4sd3_1 hold580 (.A(_00916_),
    .X(net695));
 sg13g2_dlygate4sd3_1 hold581 (.A(\u_toplayer.reg_layer2[172] ),
    .X(net696));
 sg13g2_dlygate4sd3_1 hold582 (.A(\u_toplayer.reg_layer2[192] ),
    .X(net697));
 sg13g2_dlygate4sd3_1 hold583 (.A(\u_toplayer.reg_layer1[225] ),
    .X(net698));
 sg13g2_dlygate4sd3_1 hold584 (.A(\u_toplayer.reg_layer1[95] ),
    .X(net699));
 sg13g2_dlygate4sd3_1 hold585 (.A(_00804_),
    .X(net700));
 sg13g2_dlygate4sd3_1 hold586 (.A(\u_toplayer.reg_layer1[75] ),
    .X(net701));
 sg13g2_dlygate4sd3_1 hold587 (.A(\u_toplayer.reg_layer2[41] ),
    .X(net702));
 sg13g2_dlygate4sd3_1 hold588 (.A(\u_toplayer.reg_layer2[143] ),
    .X(net703));
 sg13g2_dlygate4sd3_1 hold589 (.A(\u_toplayer.reg_layer2[79] ),
    .X(net704));
 sg13g2_dlygate4sd3_1 hold590 (.A(_00474_),
    .X(net705));
 sg13g2_dlygate4sd3_1 hold591 (.A(\u_toplayer.reg_layer2[133] ),
    .X(net706));
 sg13g2_dlygate4sd3_1 hold592 (.A(\u_toplayer.reg_layer2[207] ),
    .X(net707));
 sg13g2_dlygate4sd3_1 hold593 (.A(_00602_),
    .X(net708));
 sg13g2_dlygate4sd3_1 hold594 (.A(\u_toplayer.reg_layer2[67] ),
    .X(net709));
 sg13g2_dlygate4sd3_1 hold595 (.A(\u_toplayer.reg_layer2[195] ),
    .X(net710));
 sg13g2_dlygate4sd3_1 hold596 (.A(\u_toplayer.reg_layer1[77] ),
    .X(net711));
 sg13g2_dlygate4sd3_1 hold597 (.A(_00786_),
    .X(net712));
 sg13g2_dlygate4sd3_1 hold598 (.A(\u_toplayer.reg_layer1[134] ),
    .X(net713));
 sg13g2_dlygate4sd3_1 hold599 (.A(_05546_),
    .X(net714));
 sg13g2_dlygate4sd3_1 hold600 (.A(_00843_),
    .X(net715));
 sg13g2_dlygate4sd3_1 hold601 (.A(\u_toplayer.reg_layer2[203] ),
    .X(net716));
 sg13g2_dlygate4sd3_1 hold602 (.A(\u_toplayer.reg_layer1[68] ),
    .X(net717));
 sg13g2_dlygate4sd3_1 hold603 (.A(\u_toplayer.reg_layer1[221] ),
    .X(net718));
 sg13g2_dlygate4sd3_1 hold604 (.A(\u_toplayer.reg_layer1[43] ),
    .X(net719));
 sg13g2_dlygate4sd3_1 hold605 (.A(\u_toplayer.reg_layer1[99] ),
    .X(net720));
 sg13g2_dlygate4sd3_1 hold606 (.A(\u_toplayer.u_layer3.u_neuron.acc[16] ),
    .X(net721));
 sg13g2_dlygate4sd3_1 hold607 (.A(\u_toplayer.reg_layer2[208] ),
    .X(net722));
 sg13g2_dlygate4sd3_1 hold608 (.A(\u_toplayer.reg_layer1[53] ),
    .X(net723));
 sg13g2_dlygate4sd3_1 hold609 (.A(\u_toplayer.reg_layer1[242] ),
    .X(net724));
 sg13g2_dlygate4sd3_1 hold610 (.A(_00951_),
    .X(net725));
 sg13g2_dlygate4sd3_1 hold611 (.A(\u_toplayer.reg_layer1[104] ),
    .X(net726));
 sg13g2_dlygate4sd3_1 hold612 (.A(\u_toplayer.reg_layer1[149] ),
    .X(net727));
 sg13g2_dlygate4sd3_1 hold613 (.A(\u_toplayer.reg_layer2[240] ),
    .X(net728));
 sg13g2_dlygate4sd3_1 hold614 (.A(\u_toplayer.reg_layer1[83] ),
    .X(net729));
 sg13g2_dlygate4sd3_1 hold615 (.A(\u_toplayer.reg_layer1[67] ),
    .X(net730));
 sg13g2_dlygate4sd3_1 hold616 (.A(\u_toplayer.reg_layer2[8] ),
    .X(net731));
 sg13g2_dlygate4sd3_1 hold617 (.A(\u_toplayer.reg_layer1[54] ),
    .X(net732));
 sg13g2_dlygate4sd3_1 hold618 (.A(\u_toplayer.reg_layer1[255] ),
    .X(net733));
 sg13g2_dlygate4sd3_1 hold619 (.A(_00051_),
    .X(net734));
 sg13g2_dlygate4sd3_1 hold620 (.A(_00373_),
    .X(net735));
 sg13g2_dlygate4sd3_1 hold621 (.A(\u_toplayer.reg_layer1[205] ),
    .X(net736));
 sg13g2_dlygate4sd3_1 hold622 (.A(_00914_),
    .X(net737));
 sg13g2_dlygate4sd3_1 hold623 (.A(\u_toplayer.reg_layer1[138] ),
    .X(net738));
 sg13g2_dlygate4sd3_1 hold624 (.A(_00847_),
    .X(net739));
 sg13g2_dlygate4sd3_1 hold625 (.A(\u_toplayer.reg_layer2[211] ),
    .X(net740));
 sg13g2_dlygate4sd3_1 hold626 (.A(\u_toplayer.reg_layer2[30] ),
    .X(net741));
 sg13g2_dlygate4sd3_1 hold627 (.A(\u_toplayer.reg_layer2[39] ),
    .X(net742));
 sg13g2_dlygate4sd3_1 hold628 (.A(_00434_),
    .X(net743));
 sg13g2_dlygate4sd3_1 hold629 (.A(\u_toplayer.outreg[66] ),
    .X(net744));
 sg13g2_dlygate4sd3_1 hold630 (.A(\u_toplayer.reg_layer1[240] ),
    .X(net745));
 sg13g2_dlygate4sd3_1 hold631 (.A(\u_toplayer.reg_layer2[16] ),
    .X(net746));
 sg13g2_dlygate4sd3_1 hold632 (.A(\u_toplayer.reg_layer2[86] ),
    .X(net747));
 sg13g2_dlygate4sd3_1 hold633 (.A(\u_toplayer.reg_layer1[116] ),
    .X(net748));
 sg13g2_dlygate4sd3_1 hold634 (.A(_00825_),
    .X(net749));
 sg13g2_dlygate4sd3_1 hold635 (.A(\u_toplayer.reg_layer2[81] ),
    .X(net750));
 sg13g2_dlygate4sd3_1 hold636 (.A(\u_toplayer.reg_layer2[158] ),
    .X(net751));
 sg13g2_dlygate4sd3_1 hold637 (.A(\u_toplayer.outreg[65] ),
    .X(net752));
 sg13g2_dlygate4sd3_1 hold638 (.A(\u_toplayer.reg_layer2[73] ),
    .X(net753));
 sg13g2_dlygate4sd3_1 hold639 (.A(_00468_),
    .X(net754));
 sg13g2_dlygate4sd3_1 hold640 (.A(\u_toplayer.reg_layer1[108] ),
    .X(net755));
 sg13g2_dlygate4sd3_1 hold641 (.A(_00817_),
    .X(net756));
 sg13g2_dlygate4sd3_1 hold642 (.A(\u_toplayer.reg_layer2[204] ),
    .X(net757));
 sg13g2_dlygate4sd3_1 hold643 (.A(\u_toplayer.reg_layer2[31] ),
    .X(net758));
 sg13g2_dlygate4sd3_1 hold644 (.A(\u_toplayer.reg_layer1[210] ),
    .X(net759));
 sg13g2_dlygate4sd3_1 hold645 (.A(\u_toplayer.reg_layer2[71] ),
    .X(net760));
 sg13g2_dlygate4sd3_1 hold646 (.A(\u_toplayer.reg_layer1[164] ),
    .X(net761));
 sg13g2_dlygate4sd3_1 hold647 (.A(\u_toplayer.reg_layer1[136] ),
    .X(net762));
 sg13g2_dlygate4sd3_1 hold648 (.A(\u_toplayer.reg_layer1[213] ),
    .X(net763));
 sg13g2_dlygate4sd3_1 hold649 (.A(\u_toplayer.reg_layer2[181] ),
    .X(net764));
 sg13g2_dlygate4sd3_1 hold650 (.A(_00576_),
    .X(net765));
 sg13g2_dlygate4sd3_1 hold651 (.A(\u_toplayer.reg_layer1[170] ),
    .X(net766));
 sg13g2_dlygate4sd3_1 hold652 (.A(\u_toplayer.reg_layer2[160] ),
    .X(net767));
 sg13g2_dlygate4sd3_1 hold653 (.A(\u_toplayer.reg_layer2[215] ),
    .X(net768));
 sg13g2_dlygate4sd3_1 hold654 (.A(\u_toplayer.u_layer1.u_neuron.mult[2] ),
    .X(net769));
 sg13g2_dlygate4sd3_1 hold655 (.A(\u_toplayer.u_layer1.u_neuron.instCtrl.state[7] ),
    .X(net770));
 sg13g2_dlygate4sd3_1 hold656 (.A(_01380_),
    .X(net771));
 sg13g2_dlygate4sd3_1 hold657 (.A(_00007_),
    .X(net772));
 sg13g2_dlygate4sd3_1 hold658 (.A(\u_toplayer.reg_layer2[157] ),
    .X(net773));
 sg13g2_dlygate4sd3_1 hold659 (.A(\u_toplayer.reg_layer1[110] ),
    .X(net774));
 sg13g2_dlygate4sd3_1 hold660 (.A(_00819_),
    .X(net775));
 sg13g2_dlygate4sd3_1 hold661 (.A(\u_toplayer.reg_layer2[171] ),
    .X(net776));
 sg13g2_dlygate4sd3_1 hold662 (.A(_00566_),
    .X(net777));
 sg13g2_dlygate4sd3_1 hold663 (.A(\u_toplayer.reg_layer1[172] ),
    .X(net778));
 sg13g2_dlygate4sd3_1 hold664 (.A(\u_toplayer.reg_layer1[201] ),
    .X(net779));
 sg13g2_dlygate4sd3_1 hold665 (.A(_00910_),
    .X(net780));
 sg13g2_dlygate4sd3_1 hold666 (.A(\u_toplayer.reg_layer1[147] ),
    .X(net781));
 sg13g2_dlygate4sd3_1 hold667 (.A(\u_toplayer.reg_layer1[46] ),
    .X(net782));
 sg13g2_dlygate4sd3_1 hold668 (.A(\u_toplayer.reg_layer1[92] ),
    .X(net783));
 sg13g2_dlygate4sd3_1 hold669 (.A(_00801_),
    .X(net784));
 sg13g2_dlygate4sd3_1 hold670 (.A(\u_toplayer.u_layer2.u_neuron.acc[1] ),
    .X(net785));
 sg13g2_dlygate4sd3_1 hold671 (.A(\u_toplayer.outreg[67] ),
    .X(net786));
 sg13g2_dlygate4sd3_1 hold672 (.A(\u_toplayer.outreg[64] ),
    .X(net787));
 sg13g2_dlygate4sd3_1 hold673 (.A(\u_toplayer.reg_layer1[143] ),
    .X(net788));
 sg13g2_dlygate4sd3_1 hold674 (.A(\u_toplayer.reg_layer2[46] ),
    .X(net789));
 sg13g2_dlygate4sd3_1 hold675 (.A(_00441_),
    .X(net790));
 sg13g2_dlygate4sd3_1 hold676 (.A(\u_toplayer.outreg[71] ),
    .X(net791));
 sg13g2_dlygate4sd3_1 hold677 (.A(\u_toplayer.reg_layer1[247] ),
    .X(net792));
 sg13g2_dlygate4sd3_1 hold678 (.A(_00956_),
    .X(net793));
 sg13g2_dlygate4sd3_1 hold679 (.A(\u_toplayer.reg_layer1[37] ),
    .X(net794));
 sg13g2_dlygate4sd3_1 hold680 (.A(\u_toplayer.reg_layer1[192] ),
    .X(net795));
 sg13g2_dlygate4sd3_1 hold681 (.A(\u_toplayer.reg_layer2[177] ),
    .X(net796));
 sg13g2_dlygate4sd3_1 hold682 (.A(_00572_),
    .X(net797));
 sg13g2_dlygate4sd3_1 hold683 (.A(\u_toplayer.reg_layer1[122] ),
    .X(net798));
 sg13g2_dlygate4sd3_1 hold684 (.A(\u_toplayer.reg_layer1[141] ),
    .X(net799));
 sg13g2_dlygate4sd3_1 hold685 (.A(_00850_),
    .X(net800));
 sg13g2_dlygate4sd3_1 hold686 (.A(\u_toplayer.reg_layer1[161] ),
    .X(net801));
 sg13g2_dlygate4sd3_1 hold687 (.A(\u_toplayer.reg_layer1[185] ),
    .X(net802));
 sg13g2_dlygate4sd3_1 hold688 (.A(\u_toplayer.reg_layer2[54] ),
    .X(net803));
 sg13g2_dlygate4sd3_1 hold689 (.A(\u_toplayer.reg_layer1[190] ),
    .X(net804));
 sg13g2_dlygate4sd3_1 hold690 (.A(\u_toplayer.reg_layer2[222] ),
    .X(net805));
 sg13g2_dlygate4sd3_1 hold691 (.A(\u_toplayer.reg_layer1[17] ),
    .X(net806));
 sg13g2_dlygate4sd3_1 hold692 (.A(uo_out[2]),
    .X(net807));
 sg13g2_dlygate4sd3_1 hold693 (.A(_00175_),
    .X(net808));
 sg13g2_dlygate4sd3_1 hold694 (.A(\u_toplayer.reg_layer1[44] ),
    .X(net809));
 sg13g2_dlygate4sd3_1 hold695 (.A(\u_toplayer.reg_layer2[120] ),
    .X(net810));
 sg13g2_dlygate4sd3_1 hold696 (.A(\u_toplayer.outreg[69] ),
    .X(net811));
 sg13g2_dlygate4sd3_1 hold697 (.A(\u_toplayer.delay_counter_layer1[1] ),
    .X(net812));
 sg13g2_dlygate4sd3_1 hold698 (.A(\u_toplayer.reg_layer1[214] ),
    .X(net813));
 sg13g2_dlygate4sd3_1 hold699 (.A(\u_toplayer.reg_layer2[134] ),
    .X(net814));
 sg13g2_dlygate4sd3_1 hold700 (.A(\u_toplayer.reg_layer1[0] ),
    .X(net815));
 sg13g2_dlygate4sd3_1 hold701 (.A(\u_toplayer.outreg[50] ),
    .X(net816));
 sg13g2_dlygate4sd3_1 hold702 (.A(\u_toplayer.reg_layer1[3] ),
    .X(net817));
 sg13g2_dlygate4sd3_1 hold703 (.A(\u_toplayer.outreg[68] ),
    .X(net818));
 sg13g2_dlygate4sd3_1 hold704 (.A(\u_toplayer.reg_layer2[124] ),
    .X(net819));
 sg13g2_dlygate4sd3_1 hold705 (.A(\u_toplayer.reg_layer1[2] ),
    .X(net820));
 sg13g2_dlygate4sd3_1 hold706 (.A(\u_toplayer.u_layer2.u_neuron.acc[5] ),
    .X(net821));
 sg13g2_dlygate4sd3_1 hold707 (.A(\u_toplayer.u_outlayer.u_neuron.acc[1] ),
    .X(net822));
 sg13g2_dlygate4sd3_1 hold708 (.A(\u_toplayer.u_outlayer.u_neuron.acc[16] ),
    .X(net823));
 sg13g2_dlygate4sd3_1 hold709 (.A(\u_toplayer.reg_layer1[1] ),
    .X(net824));
 sg13g2_dlygate4sd3_1 hold710 (.A(\u_toplayer.u_layer1.u_neuron.mult[0] ),
    .X(net825));
 sg13g2_dlygate4sd3_1 hold711 (.A(\u_toplayer.outreg[52] ),
    .X(net826));
 sg13g2_dlygate4sd3_1 hold712 (.A(\u_toplayer.reg_layer1[209] ),
    .X(net827));
 sg13g2_dlygate4sd3_1 hold713 (.A(\u_toplayer.reg_layer2[170] ),
    .X(net828));
 sg13g2_dlygate4sd3_1 hold714 (.A(_00565_),
    .X(net829));
 sg13g2_dlygate4sd3_1 hold715 (.A(\u_toplayer.u_layer2.u_neuron.mult[2] ),
    .X(net830));
 sg13g2_dlygate4sd3_1 hold716 (.A(_00052_),
    .X(net831));
 sg13g2_dlygate4sd3_1 hold717 (.A(_00221_),
    .X(net832));
 sg13g2_dlygate4sd3_1 hold718 (.A(\u_toplayer.u_outlayer.u_neuron.mult[11] ),
    .X(net833));
 sg13g2_dlygate4sd3_1 hold719 (.A(\u_toplayer.reg_layer2[214] ),
    .X(net834));
 sg13g2_dlygate4sd3_1 hold720 (.A(\u_toplayer.reg_layer2[248] ),
    .X(net835));
 sg13g2_dlygate4sd3_1 hold721 (.A(\u_toplayer.u_outlayer.u_neuron.mult[3] ),
    .X(net836));
 sg13g2_dlygate4sd3_1 hold722 (.A(\u_toplayer.reg_layer2[34] ),
    .X(net837));
 sg13g2_dlygate4sd3_1 hold723 (.A(_00429_),
    .X(net838));
 sg13g2_dlygate4sd3_1 hold724 (.A(\u_toplayer.outreg[49] ),
    .X(net839));
 sg13g2_dlygate4sd3_1 hold725 (.A(\u_toplayer.u_layer3.stateout[0] ),
    .X(net840));
 sg13g2_dlygate4sd3_1 hold726 (.A(_00340_),
    .X(net841));
 sg13g2_dlygate4sd3_1 hold727 (.A(\u_toplayer.reg_layer2[42] ),
    .X(net842));
 sg13g2_dlygate4sd3_1 hold728 (.A(_00437_),
    .X(net843));
 sg13g2_dlygate4sd3_1 hold729 (.A(\u_toplayer.outreg[55] ),
    .X(net844));
 sg13g2_dlygate4sd3_1 hold730 (.A(\u_toplayer.u_layer1.u_neuron.b[4] ),
    .X(net845));
 sg13g2_dlygate4sd3_1 hold731 (.A(\u_toplayer.reg_layer2[12] ),
    .X(net846));
 sg13g2_dlygate4sd3_1 hold732 (.A(_00407_),
    .X(net847));
 sg13g2_dlygate4sd3_1 hold733 (.A(\u_toplayer.outreg[70] ),
    .X(net848));
 sg13g2_dlygate4sd3_1 hold734 (.A(uo_out[3]),
    .X(net849));
 sg13g2_dlygate4sd3_1 hold735 (.A(_00176_),
    .X(net850));
 sg13g2_dlygate4sd3_1 hold736 (.A(\u_toplayer.outreg[62] ),
    .X(net851));
 sg13g2_dlygate4sd3_1 hold737 (.A(\u_toplayer.outreg[57] ),
    .X(net852));
 sg13g2_dlygate4sd3_1 hold738 (.A(\u_toplayer.reg_layer1[223] ),
    .X(net853));
 sg13g2_dlygate4sd3_1 hold739 (.A(_00932_),
    .X(net854));
 sg13g2_dlygate4sd3_1 hold740 (.A(\u_toplayer.outreg[61] ),
    .X(net855));
 sg13g2_dlygate4sd3_1 hold741 (.A(\u_toplayer.u_layer1.u_neuron.mult[10] ),
    .X(net856));
 sg13g2_dlygate4sd3_1 hold742 (.A(\u_toplayer.u_layer3.u_neuron.mult[6] ),
    .X(net857));
 sg13g2_dlygate4sd3_1 hold743 (.A(\u_toplayer.reg_layer2[144] ),
    .X(net858));
 sg13g2_dlygate4sd3_1 hold744 (.A(\u_toplayer.outreg[54] ),
    .X(net859));
 sg13g2_dlygate4sd3_1 hold745 (.A(\u_toplayer.u_layer2.statel2[0] ),
    .X(net860));
 sg13g2_dlygate4sd3_1 hold746 (.A(\u_toplayer.outreg[53] ),
    .X(net861));
 sg13g2_dlygate4sd3_1 hold747 (.A(\u_toplayer.outreg[56] ),
    .X(net862));
 sg13g2_dlygate4sd3_1 hold748 (.A(\u_toplayer.u_layer3.stateout[3] ),
    .X(net863));
 sg13g2_dlygate4sd3_1 hold749 (.A(_00343_),
    .X(net864));
 sg13g2_dlygate4sd3_1 hold750 (.A(\u_toplayer.outreg[51] ),
    .X(net865));
 sg13g2_dlygate4sd3_1 hold751 (.A(uo_out[6]),
    .X(net866));
 sg13g2_dlygate4sd3_1 hold752 (.A(_00179_),
    .X(net867));
 sg13g2_dlygate4sd3_1 hold753 (.A(\u_toplayer.outreg[48] ),
    .X(net868));
 sg13g2_dlygate4sd3_1 hold754 (.A(\u_toplayer.outreg[58] ),
    .X(net869));
 sg13g2_dlygate4sd3_1 hold755 (.A(\u_toplayer.reg_layer2[129] ),
    .X(net870));
 sg13g2_dlygate4sd3_1 hold756 (.A(_00042_),
    .X(net871));
 sg13g2_dlygate4sd3_1 hold757 (.A(_01359_),
    .X(net872));
 sg13g2_dlygate4sd3_1 hold758 (.A(_00018_),
    .X(net873));
 sg13g2_dlygate4sd3_1 hold759 (.A(\u_toplayer.u_outlayer.u_neuron.mult[4] ),
    .X(net874));
 sg13g2_dlygate4sd3_1 hold760 (.A(_00153_),
    .X(net875));
 sg13g2_dlygate4sd3_1 hold761 (.A(\u_toplayer.reg_layer1[4] ),
    .X(net876));
 sg13g2_dlygate4sd3_1 hold762 (.A(\u_toplayer.u_layer1.statel1[5] ),
    .X(net877));
 sg13g2_dlygate4sd3_1 hold763 (.A(_00986_),
    .X(net878));
 sg13g2_dlygate4sd3_1 hold764 (.A(\u_toplayer.reg_layer1[7] ),
    .X(net879));
 sg13g2_dlygate4sd3_1 hold765 (.A(\u_toplayer.reg_layer2[152] ),
    .X(net880));
 sg13g2_dlygate4sd3_1 hold766 (.A(\u_toplayer.u_layer3.u_neuron.instCtrl.state[5] ),
    .X(net881));
 sg13g2_dlygate4sd3_1 hold767 (.A(_00020_),
    .X(net882));
 sg13g2_dlygate4sd3_1 hold768 (.A(uo_out[1]),
    .X(net883));
 sg13g2_dlygate4sd3_1 hold769 (.A(\u_toplayer.outreg[63] ),
    .X(net884));
 sg13g2_dlygate4sd3_1 hold770 (.A(\u_toplayer.reg_layer1[105] ),
    .X(net885));
 sg13g2_dlygate4sd3_1 hold771 (.A(\u_toplayer.u_layer1.u_neuron.acc[16] ),
    .X(net886));
 sg13g2_dlygate4sd3_1 hold772 (.A(\u_toplayer.outreg[60] ),
    .X(net887));
 sg13g2_dlygate4sd3_1 hold773 (.A(\u_toplayer.u_layer2.u_neuron.mult[3] ),
    .X(net888));
 sg13g2_dlygate4sd3_1 hold774 (.A(\u_toplayer.u_layer3.u_neuron.mult[2] ),
    .X(net889));
 sg13g2_dlygate4sd3_1 hold775 (.A(\u_toplayer.u_layer1.u_neuron.mult[8] ),
    .X(net890));
 sg13g2_dlygate4sd3_1 hold776 (.A(\u_toplayer.reg_layer1[38] ),
    .X(net891));
 sg13g2_dlygate4sd3_1 hold777 (.A(\u_toplayer.done_layer3 ),
    .X(net892));
 sg13g2_dlygate4sd3_1 hold778 (.A(_00323_),
    .X(net893));
 sg13g2_dlygate4sd3_1 hold779 (.A(\u_toplayer.outreg[59] ),
    .X(net894));
 sg13g2_dlygate4sd3_1 hold780 (.A(\u_toplayer.u_layer3.stateout[5] ),
    .X(net895));
 sg13g2_dlygate4sd3_1 hold781 (.A(_00345_),
    .X(net896));
 sg13g2_dlygate4sd3_1 hold782 (.A(\u_toplayer.u_layer2.u_neuron.mult[4] ),
    .X(net897));
 sg13g2_dlygate4sd3_1 hold783 (.A(\u_toplayer.u_layer3.u_neuron.acc[20] ),
    .X(net898));
 sg13g2_dlygate4sd3_1 hold784 (.A(uo_out[4]),
    .X(net899));
 sg13g2_dlygate4sd3_1 hold785 (.A(_00177_),
    .X(net900));
 sg13g2_dlygate4sd3_1 hold786 (.A(\u_toplayer.u_outlayer.u_neuron.mult[0] ),
    .X(net901));
 sg13g2_dlygate4sd3_1 hold787 (.A(_00149_),
    .X(net902));
 sg13g2_dlygate4sd3_1 hold788 (.A(uo_out[0]),
    .X(net903));
 sg13g2_dlygate4sd3_1 hold789 (.A(_01899_),
    .X(net904));
 sg13g2_dlygate4sd3_1 hold790 (.A(_00173_),
    .X(net905));
 sg13g2_dlygate4sd3_1 hold791 (.A(\u_toplayer.reg_layer1[5] ),
    .X(net906));
 sg13g2_dlygate4sd3_1 hold792 (.A(\u_toplayer.delay_counter_layer3[1] ),
    .X(net907));
 sg13g2_dlygate4sd3_1 hold793 (.A(uo_out[5]),
    .X(net908));
 sg13g2_dlygate4sd3_1 hold794 (.A(_00178_),
    .X(net909));
 sg13g2_dlygate4sd3_1 hold795 (.A(\u_toplayer.u_layer1.u_neuron.mult[9] ),
    .X(net910));
 sg13g2_dlygate4sd3_1 hold796 (.A(\u_toplayer.reg_layer2[0] ),
    .X(net911));
 sg13g2_dlygate4sd3_1 hold797 (.A(\u_toplayer.reg_layer2[2] ),
    .X(net912));
 sg13g2_dlygate4sd3_1 hold798 (.A(\u_toplayer.reg_layer2[1] ),
    .X(net913));
 sg13g2_dlygate4sd3_1 hold799 (.A(\u_toplayer.reg_layer2[4] ),
    .X(net914));
 sg13g2_dlygate4sd3_1 hold800 (.A(\u_toplayer.reg_layer1[6] ),
    .X(net915));
 sg13g2_dlygate4sd3_1 hold801 (.A(\u_toplayer.u_layer2.u_neuron.mult[8] ),
    .X(net916));
 sg13g2_dlygate4sd3_1 hold802 (.A(\u_toplayer.u_layer3.u_neuron.mult[3] ),
    .X(net917));
 sg13g2_dlygate4sd3_1 hold803 (.A(\u_toplayer.u_layer1.u_neuron.instCtrl.state[3] ),
    .X(net918));
 sg13g2_dlygate4sd3_1 hold804 (.A(_00003_),
    .X(net919));
 sg13g2_dlygate4sd3_1 hold805 (.A(\u_toplayer.u_outlayer.u_neuron.mult[2] ),
    .X(net920));
 sg13g2_dlygate4sd3_1 hold806 (.A(\u_toplayer.u_layer1.statel1[1] ),
    .X(net921));
 sg13g2_dlygate4sd3_1 hold807 (.A(_00982_),
    .X(net922));
 sg13g2_dlygate4sd3_1 hold808 (.A(\u_toplayer.u_layer1.u_neuron.mult[5] ),
    .X(net923));
 sg13g2_dlygate4sd3_1 hold809 (.A(\u_toplayer.u_layer3.u_neuron.acc[8] ),
    .X(net924));
 sg13g2_dlygate4sd3_1 hold810 (.A(\u_toplayer.delay_counter_layer2[1] ),
    .X(net925));
 sg13g2_dlygate4sd3_1 hold811 (.A(_01017_),
    .X(net926));
 sg13g2_dlygate4sd3_1 hold812 (.A(\u_toplayer.u_layer3.u_neuron.mult[0] ),
    .X(net927));
 sg13g2_dlygate4sd3_1 hold813 (.A(_00181_),
    .X(net928));
 sg13g2_dlygate4sd3_1 hold814 (.A(\u_toplayer.u_layer2.u_neuron.mult[0] ),
    .X(net929));
 sg13g2_dlygate4sd3_1 hold815 (.A(_00227_),
    .X(net930));
 sg13g2_dlygate4sd3_1 hold816 (.A(_00041_),
    .X(net931));
 sg13g2_dlygate4sd3_1 hold817 (.A(_01357_),
    .X(net932));
 sg13g2_dlygate4sd3_1 hold818 (.A(_01358_),
    .X(net933));
 sg13g2_dlygate4sd3_1 hold819 (.A(_00017_),
    .X(net934));
 sg13g2_dlygate4sd3_1 hold820 (.A(\u_toplayer.reg_layer2[5] ),
    .X(net935));
 sg13g2_dlygate4sd3_1 hold821 (.A(\u_toplayer.reg_layer2[3] ),
    .X(net936));
 sg13g2_dlygate4sd3_1 hold822 (.A(\u_toplayer.u_layer2.statel2[5] ),
    .X(net937));
 sg13g2_dlygate4sd3_1 hold823 (.A(_00673_),
    .X(net938));
 sg13g2_dlygate4sd3_1 hold824 (.A(\u_toplayer.u_layer3.stateout[2] ),
    .X(net939));
 sg13g2_dlygate4sd3_1 hold825 (.A(_01201_),
    .X(net940));
 sg13g2_dlygate4sd3_1 hold826 (.A(_00342_),
    .X(net941));
 sg13g2_dlygate4sd3_1 hold827 (.A(\u_toplayer.u_layer3.u_neuron.mult[7] ),
    .X(net942));
 sg13g2_dlygate4sd3_1 hold828 (.A(\u_toplayer.done_layer1 ),
    .X(net943));
 sg13g2_dlygate4sd3_1 hold829 (.A(\u_toplayer.u_layer2.u_neuron.mult[7] ),
    .X(net944));
 sg13g2_dlygate4sd3_1 hold830 (.A(\u_toplayer.u_layer1.u_neuron.mult[6] ),
    .X(net945));
 sg13g2_dlygate4sd3_1 hold831 (.A(\u_toplayer.reg_layer2[6] ),
    .X(net946));
 sg13g2_dlygate4sd3_1 hold832 (.A(\u_toplayer.u_layer3.u_neuron.mult[4] ),
    .X(net947));
 sg13g2_dlygate4sd3_1 hold833 (.A(\u_toplayer.u_layer2.u_neuron.mult[5] ),
    .X(net948));
 sg13g2_dlygate4sd3_1 hold834 (.A(\u_toplayer.u_layer2.u_neuron.mult[12] ),
    .X(net949));
 sg13g2_dlygate4sd3_1 hold835 (.A(\u_toplayer.u_layer2.u_neuron.mult[9] ),
    .X(net950));
 sg13g2_dlygate4sd3_1 hold836 (.A(\u_toplayer.u_layer1.u_neuron.mult[11] ),
    .X(net951));
 sg13g2_dlygate4sd3_1 hold837 (.A(\u_toplayer.u_outlayer.u_neuron.mult[6] ),
    .X(net952));
 sg13g2_dlygate4sd3_1 hold838 (.A(\u_toplayer.u_layer1.u_neuron.mult[3] ),
    .X(net953));
 sg13g2_dlygate4sd3_1 hold839 (.A(\u_toplayer.u_layer2.statel2[1] ),
    .X(net954));
 sg13g2_dlygate4sd3_1 hold840 (.A(\u_toplayer.u_outlayer.u_neuron.mult[5] ),
    .X(net955));
 sg13g2_dlygate4sd3_1 hold841 (.A(\u_toplayer.reg_layer2[7] ),
    .X(net956));
 sg13g2_dlygate4sd3_1 hold842 (.A(\u_toplayer.u_layer3.u_neuron.mult[9] ),
    .X(net957));
 sg13g2_dlygate4sd3_1 hold843 (.A(_00035_),
    .X(net958));
 sg13g2_dlygate4sd3_1 hold844 (.A(_00028_),
    .X(net959));
 sg13g2_dlygate4sd3_1 hold845 (.A(\u_toplayer.u_layer1.statel1[3] ),
    .X(net960));
 sg13g2_dlygate4sd3_1 hold846 (.A(_00984_),
    .X(net961));
 sg13g2_dlygate4sd3_1 hold847 (.A(\u_toplayer.u_layer1.u_neuron.mult[7] ),
    .X(net962));
 sg13g2_dlygate4sd3_1 hold848 (.A(\u_toplayer.u_layer3.u_neuron.mult[8] ),
    .X(net963));
 sg13g2_dlygate4sd3_1 hold849 (.A(_00038_),
    .X(net964));
 sg13g2_dlygate4sd3_1 hold850 (.A(_01341_),
    .X(net965));
 sg13g2_dlygate4sd3_1 hold851 (.A(_01342_),
    .X(net966));
 sg13g2_dlygate4sd3_1 hold852 (.A(_00023_),
    .X(net967));
 sg13g2_dlygate4sd3_1 hold853 (.A(_00030_),
    .X(net968));
 sg13g2_dlygate4sd3_1 hold854 (.A(_05687_),
    .X(net969));
 sg13g2_dlygate4sd3_1 hold855 (.A(_05711_),
    .X(net970));
 sg13g2_dlygate4sd3_1 hold856 (.A(_00980_),
    .X(net971));
 sg13g2_dlygate4sd3_1 hold857 (.A(\u_toplayer.u_layer1.statel1[7] ),
    .X(net972));
 sg13g2_dlygate4sd3_1 hold858 (.A(_00988_),
    .X(net973));
 sg13g2_dlygate4sd3_1 hold859 (.A(\u_toplayer.u_layer3.u_neuron.mult[13] ),
    .X(net974));
 sg13g2_dlygate4sd3_1 hold860 (.A(\u_toplayer.u_layer2.u_neuron.mult[6] ),
    .X(net975));
 sg13g2_dlygate4sd3_1 hold861 (.A(\u_toplayer.u_layer1.u_neuron.mult[4] ),
    .X(net976));
 sg13g2_dlygate4sd3_1 hold862 (.A(\u_toplayer.u_layer2.u_neuron.mult[10] ),
    .X(net977));
 sg13g2_dlygate4sd3_1 hold863 (.A(\u_toplayer.u_layer3.stateout[1] ),
    .X(net978));
 sg13g2_dlygate4sd3_1 hold864 (.A(\u_toplayer.u_layer2.statel2[3] ),
    .X(net979));
 sg13g2_dlygate4sd3_1 hold865 (.A(\u_toplayer.done_layer2 ),
    .X(net980));
 sg13g2_dlygate4sd3_1 hold866 (.A(_00651_),
    .X(net981));
 sg13g2_dlygate4sd3_1 hold867 (.A(\u_toplayer.u_layer2.neuron_index[5] ),
    .X(net982));
 sg13g2_dlygate4sd3_1 hold868 (.A(_00378_),
    .X(net983));
 sg13g2_dlygate4sd3_1 hold869 (.A(uo_out[7]),
    .X(net984));
 sg13g2_dlygate4sd3_1 hold870 (.A(_00180_),
    .X(net985));
 sg13g2_dlygate4sd3_1 hold871 (.A(\u_toplayer.u_layer1.u_neuron.mult[1] ),
    .X(net986));
 sg13g2_dlygate4sd3_1 hold872 (.A(\u_toplayer.u_layer1.statel1[0] ),
    .X(net987));
 sg13g2_dlygate4sd3_1 hold873 (.A(\u_toplayer.u_outlayer.u_neuron.mult[7] ),
    .X(net988));
 sg13g2_dlygate4sd3_1 hold874 (.A(\u_toplayer.u_layer1.u_neuron.mult[12] ),
    .X(net989));
 sg13g2_dlygate4sd3_1 hold875 (.A(\u_toplayer.u_layer3.u_neuron.mult[10] ),
    .X(net990));
 sg13g2_dlygate4sd3_1 hold876 (.A(\u_toplayer.u_outlayer.u_neuron.mult[1] ),
    .X(net991));
 sg13g2_dlygate4sd3_1 hold877 (.A(\u_toplayer.u_layer1.u_neuron.b[0] ),
    .X(net992));
 sg13g2_dlygate4sd3_1 hold878 (.A(\u_toplayer.u_layer3.neuron_index[1] ),
    .X(net993));
 sg13g2_dlygate4sd3_1 hold879 (.A(\u_toplayer.u_layer1.statel1[2] ),
    .X(net994));
 sg13g2_dlygate4sd3_1 hold880 (.A(\u_toplayer.u_layer3.u_neuron.mult[1] ),
    .X(net995));
 sg13g2_dlygate4sd3_1 hold881 (.A(\u_toplayer.u_layer3.u_neuron.mult[5] ),
    .X(net996));
 sg13g2_dlygate4sd3_1 hold882 (.A(\u_toplayer.u_layer1.u_neuron.b[1] ),
    .X(net997));
 sg13g2_dlygate4sd3_1 hold883 (.A(\u_toplayer.u_layer3.u_neuron.mult[12] ),
    .X(net998));
 sg13g2_dlygate4sd3_1 hold884 (.A(_00040_),
    .X(net999));
 sg13g2_dlygate4sd3_1 hold885 (.A(_01356_),
    .X(net1000));
 sg13g2_dlygate4sd3_1 hold886 (.A(_00016_),
    .X(net1001));
 sg13g2_dlygate4sd3_1 hold887 (.A(\u_toplayer.u_layer2.u_neuron.mult[14] ),
    .X(net1002));
 sg13g2_dlygate4sd3_1 hold888 (.A(\u_toplayer.u_layer2.u_neuron.mult[1] ),
    .X(net1003));
 sg13g2_dlygate4sd3_1 hold889 (.A(\u_toplayer.u_layer2.u_neuron.mult[13] ),
    .X(net1004));
 sg13g2_dlygate4sd3_1 hold890 (.A(_00037_),
    .X(net1005));
 sg13g2_dlygate4sd3_1 hold891 (.A(_00022_),
    .X(net1006));
 sg13g2_dlygate4sd3_1 hold892 (.A(\u_toplayer.u_layer1.u_neuron.mult[13] ),
    .X(net1007));
 sg13g2_dlygate4sd3_1 hold893 (.A(\u_toplayer.u_outlayer.u_neuron.mult[8] ),
    .X(net1008));
 sg13g2_dlygate4sd3_1 hold894 (.A(\u_toplayer.u_layer2.statel2[2] ),
    .X(net1009));
 sg13g2_dlygate4sd3_1 hold895 (.A(\u_toplayer.u_layer1.neuron_index[5] ),
    .X(net1010));
 sg13g2_dlygate4sd3_1 hold896 (.A(_00706_),
    .X(net1011));
 sg13g2_dlygate4sd3_1 hold897 (.A(\u_toplayer.u_layer3.u_neuron.mult[11] ),
    .X(net1012));
 sg13g2_dlygate4sd3_1 hold898 (.A(\u_toplayer.u_layer2.u_neuron.mult[11] ),
    .X(net1013));
 sg13g2_dlygate4sd3_1 hold899 (.A(\u_toplayer.u_layer1.u_neuron.b[6] ),
    .X(net1014));
 sg13g2_dlygate4sd3_1 hold900 (.A(\u_toplayer.u_layer1.statel1[6] ),
    .X(net1015));
 sg13g2_dlygate4sd3_1 hold901 (.A(_00987_),
    .X(net1016));
 sg13g2_dlygate4sd3_1 hold902 (.A(\u_toplayer.u_outlayer.u_neuron.mult[9] ),
    .X(net1017));
 sg13g2_dlygate4sd3_1 hold903 (.A(\u_toplayer.u_layer1.u_neuron.b[2] ),
    .X(net1018));
 sg13g2_dlygate4sd3_1 hold904 (.A(\u_toplayer.u_layer1.u_neuron.b[5] ),
    .X(net1019));
 sg13g2_dlygate4sd3_1 hold905 (.A(\u_toplayer.u_layer1.u_neuron.b[3] ),
    .X(net1020));
 sg13g2_dlygate4sd3_1 hold906 (.A(\u_toplayer.u_layer3.u_neuron.mult[14] ),
    .X(net1021));
 sg13g2_dlygate4sd3_1 hold907 (.A(\u_toplayer.u_layer3.u_neuron.din[0] ),
    .X(net1022));
 sg13g2_dlygate4sd3_1 hold908 (.A(\u_toplayer.u_layer3.u_neuron.din[5] ),
    .X(net1023));
 sg13g2_dlygate4sd3_1 hold909 (.A(\u_toplayer.u_layer3.neuron_index[5] ),
    .X(net1024));
 sg13g2_dlygate4sd3_1 hold910 (.A(_00226_),
    .X(net1025));
 sg13g2_dlygate4sd3_1 hold911 (.A(\u_toplayer.u_layer3.sum[1] ),
    .X(net1026));
 sg13g2_dlygate4sd3_1 hold912 (.A(_00333_),
    .X(net1027));
 sg13g2_dlygate4sd3_1 hold913 (.A(\u_toplayer.u_layer1.neuron_index[4] ),
    .X(net1028));
 sg13g2_dlygate4sd3_1 hold914 (.A(_00705_),
    .X(net1029));
 sg13g2_dlygate4sd3_1 hold915 (.A(\u_toplayer.u_layer3.sum[4] ),
    .X(net1030));
 sg13g2_dlygate4sd3_1 hold916 (.A(_00336_),
    .X(net1031));
 sg13g2_dlygate4sd3_1 hold917 (.A(\u_toplayer.u_layer3.u_neuron.acc[23] ),
    .X(net1032));
 sg13g2_dlygate4sd3_1 hold918 (.A(_00339_),
    .X(net1033));
 sg13g2_dlygate4sd3_1 hold919 (.A(\u_toplayer.u_layer3.neuron_index[4] ),
    .X(net1034));
 sg13g2_dlygate4sd3_1 hold920 (.A(_00225_),
    .X(net1035));
 sg13g2_dlygate4sd3_1 hold921 (.A(\u_toplayer.u_layer3.stateout[4] ),
    .X(net1036));
 sg13g2_dlygate4sd3_1 hold922 (.A(\u_toplayer.u_layer2.u_neuron.acc[0] ),
    .X(net1037));
 sg13g2_dlygate4sd3_1 hold923 (.A(_00677_),
    .X(net1038));
 sg13g2_dlygate4sd3_1 hold924 (.A(\u_toplayer.u_layer1.u_neuron.instCtrl.state[8] ),
    .X(net1039));
 sg13g2_dlygate4sd3_1 hold925 (.A(_01370_),
    .X(net1040));
 sg13g2_dlygate4sd3_1 hold926 (.A(_00008_),
    .X(net1041));
 sg13g2_dlygate4sd3_1 hold927 (.A(\u_toplayer.u_outlayer.u_neuron.acc[23] ),
    .X(net1042));
 sg13g2_dlygate4sd3_1 hold928 (.A(\u_toplayer.u_layer1.neuron_index[3] ),
    .X(net1043));
 sg13g2_dlygate4sd3_1 hold929 (.A(\u_toplayer.u_layer3.sum[6] ),
    .X(net1044));
 sg13g2_dlygate4sd3_1 hold930 (.A(_00338_),
    .X(net1045));
 sg13g2_dlygate4sd3_1 hold931 (.A(\u_toplayer.u_layer3.u_neuron.acc[17] ),
    .X(net1046));
 sg13g2_dlygate4sd3_1 hold932 (.A(\u_toplayer.u_layer3.u_neuron.acc[0] ),
    .X(net1047));
 sg13g2_dlygate4sd3_1 hold933 (.A(_00349_),
    .X(net1048));
 sg13g2_dlygate4sd3_1 hold934 (.A(\u_toplayer.u_layer1.u_neuron.acc[15] ),
    .X(net1049));
 sg13g2_dlygate4sd3_1 hold935 (.A(\u_toplayer.u_layer2.u_neuron.acc[22] ),
    .X(net1050));
 sg13g2_dlygate4sd3_1 hold936 (.A(\u_toplayer.u_outlayer.u_neuron.acc[21] ),
    .X(net1051));
 sg13g2_dlygate4sd3_1 hold937 (.A(\u_toplayer.u_layer3.u_neuron.acc[19] ),
    .X(net1052));
 sg13g2_dlygate4sd3_1 hold938 (.A(\u_toplayer.u_layer3.sum[2] ),
    .X(net1053));
 sg13g2_dlygate4sd3_1 hold939 (.A(_00334_),
    .X(net1054));
 sg13g2_dlygate4sd3_1 hold940 (.A(\u_toplayer.u_layer2.u_neuron.acc[6] ),
    .X(net1055));
 sg13g2_dlygate4sd3_1 hold941 (.A(\u_toplayer.u_outlayer.u_neuron.din[5] ),
    .X(net1056));
 sg13g2_dlygate4sd3_1 hold942 (.A(_00170_),
    .X(net1057));
 sg13g2_dlygate4sd3_1 hold943 (.A(\u_toplayer.u_outlayer.u_neuron.acc[15] ),
    .X(net1058));
 sg13g2_dlygate4sd3_1 hold944 (.A(\u_toplayer.u_layer2.u_neuron.mult[15] ),
    .X(net1059));
 sg13g2_dlygate4sd3_1 hold945 (.A(\u_toplayer.u_outlayer.u_neuron.mult[12] ),
    .X(net1060));
 sg13g2_dlygate4sd3_1 hold946 (.A(\u_toplayer.u_layer3.u_neuron.acc[2] ),
    .X(net1061));
 sg13g2_dlygate4sd3_1 hold947 (.A(\u_toplayer.u_layer1.u_neuron.acc[21] ),
    .X(net1062));
 sg13g2_dlygate4sd3_1 hold948 (.A(\u_toplayer.u_layer1.u_neuron.acc[17] ),
    .X(net1063));
 sg13g2_dlygate4sd3_1 hold949 (.A(\u_toplayer.u_layer1.u_neuron.acc[23] ),
    .X(net1064));
 sg13g2_dlygate4sd3_1 hold950 (.A(\u_toplayer.u_layer1.u_neuron.instCtrl.state[1] ),
    .X(net1065));
 sg13g2_dlygate4sd3_1 hold951 (.A(_01366_),
    .X(net1066));
 sg13g2_dlygate4sd3_1 hold952 (.A(\u_toplayer.u_outlayer.u_neuron.acc[19] ),
    .X(net1067));
 sg13g2_dlygate4sd3_1 hold953 (.A(\u_toplayer.u_layer3.u_neuron.acc[23] ),
    .X(net1068));
 sg13g2_dlygate4sd3_1 hold954 (.A(\u_toplayer.u_layer1.u_neuron.acc[0] ),
    .X(net1069));
 sg13g2_dlygate4sd3_1 hold955 (.A(\u_toplayer.u_layer2.u_neuron.acc[9] ),
    .X(net1070));
 sg13g2_dlygate4sd3_1 hold956 (.A(\u_toplayer.u_layer2.u_neuron.instCtrl.state[5] ),
    .X(net1071));
 sg13g2_dlygate4sd3_1 hold957 (.A(_01351_),
    .X(net1072));
 sg13g2_dlygate4sd3_1 hold958 (.A(_00014_),
    .X(net1073));
 sg13g2_dlygate4sd3_1 hold959 (.A(\u_toplayer.u_layer1.u_neuron.acc[22] ),
    .X(net1074));
 sg13g2_dlygate4sd3_1 hold960 (.A(\u_toplayer.u_layer2.neuron_index[4] ),
    .X(net1075));
 sg13g2_dlygate4sd3_1 hold961 (.A(\u_toplayer.u_layer3.sum[3] ),
    .X(net1076));
 sg13g2_dlygate4sd3_1 hold962 (.A(_00335_),
    .X(net1077));
 sg13g2_dlygate4sd3_1 hold963 (.A(\u_toplayer.u_outlayer.u_neuron.mult[10] ),
    .X(net1078));
 sg13g2_dlygate4sd3_1 hold964 (.A(\u_toplayer.u_outlayer.u_neuron.acc[17] ),
    .X(net1079));
 sg13g2_dlygate4sd3_1 hold965 (.A(\u_toplayer.u_layer3.u_neuron.din[4] ),
    .X(net1080));
 sg13g2_dlygate4sd3_1 hold966 (.A(\u_toplayer.u_layer2.u_neuron.acc[19] ),
    .X(net1081));
 sg13g2_dlygate4sd3_1 hold967 (.A(\u_toplayer.u_layer1.u_neuron.mult[14] ),
    .X(net1082));
 sg13g2_dlygate4sd3_1 hold968 (.A(\u_toplayer.u_outlayer.u_neuron.acc[11] ),
    .X(net1083));
 sg13g2_dlygate4sd3_1 hold969 (.A(\u_toplayer.u_layer1.u_neuron.acc[2] ),
    .X(net1084));
 sg13g2_dlygate4sd3_1 hold970 (.A(\u_toplayer.u_layer3.sum[0] ),
    .X(net1085));
 sg13g2_dlygate4sd3_1 hold971 (.A(\u_toplayer.u_layer3.u_neuron.acc[1] ),
    .X(net1086));
 sg13g2_dlygate4sd3_1 hold972 (.A(_00350_),
    .X(net1087));
 sg13g2_dlygate4sd3_1 hold973 (.A(\u_toplayer.u_layer3.u_neuron.acc[15] ),
    .X(net1088));
 sg13g2_dlygate4sd3_1 hold974 (.A(\u_toplayer.u_outlayer.u_neuron.acc[0] ),
    .X(net1089));
 sg13g2_dlygate4sd3_1 hold975 (.A(\u_toplayer.u_outlayer.u_neuron.din[7] ),
    .X(net1090));
 sg13g2_dlygate4sd3_1 hold976 (.A(_00172_),
    .X(net1091));
 sg13g2_dlygate4sd3_1 hold977 (.A(\u_toplayer.u_layer3.u_neuron.din[3] ),
    .X(net1092));
 sg13g2_dlygate4sd3_1 hold978 (.A(\u_toplayer.u_outlayer.u_neuron.din[1] ),
    .X(net1093));
 sg13g2_dlygate4sd3_1 hold979 (.A(_00166_),
    .X(net1094));
 sg13g2_dlygate4sd3_1 hold980 (.A(\u_toplayer.u_layer3.u_neuron.acc[13] ),
    .X(net1095));
 sg13g2_dlygate4sd3_1 hold981 (.A(\u_toplayer.u_outlayer.u_neuron.din[6] ),
    .X(net1096));
 sg13g2_dlygate4sd3_1 hold982 (.A(_00171_),
    .X(net1097));
 sg13g2_dlygate4sd3_1 hold983 (.A(\u_toplayer.u_layer3.neuron_index[2] ),
    .X(net1098));
 sg13g2_dlygate4sd3_1 hold984 (.A(_00223_),
    .X(net1099));
 sg13g2_dlygate4sd3_1 hold985 (.A(\u_toplayer.u_outlayer.u_neuron.acc[3] ),
    .X(net1100));
 sg13g2_dlygate4sd3_1 hold986 (.A(\u_toplayer.u_layer3.sum[5] ),
    .X(net1101));
 sg13g2_dlygate4sd3_1 hold987 (.A(_00337_),
    .X(net1102));
 sg13g2_dlygate4sd3_1 hold988 (.A(\u_toplayer.u_layer1.statel1[4] ),
    .X(net1103));
 sg13g2_dlygate4sd3_1 hold989 (.A(\u_toplayer.u_layer2.u_neuron.acc[17] ),
    .X(net1104));
 sg13g2_dlygate4sd3_1 hold990 (.A(_00694_),
    .X(net1105));
 sg13g2_dlygate4sd3_1 hold991 (.A(\u_toplayer.u_layer1.u_neuron.instCtrl.state[2] ),
    .X(net1106));
 sg13g2_dlygate4sd3_1 hold992 (.A(_01371_),
    .X(net1107));
 sg13g2_dlygate4sd3_1 hold993 (.A(_00002_),
    .X(net1108));
 sg13g2_dlygate4sd3_1 hold994 (.A(\u_toplayer.u_layer3.u_neuron.acc[22] ),
    .X(net1109));
 sg13g2_dlygate4sd3_1 hold995 (.A(\u_toplayer.u_outlayer.u_neuron.acc[22] ),
    .X(net1110));
 sg13g2_dlygate4sd3_1 hold996 (.A(\u_toplayer.u_layer3.u_neuron.acc[3] ),
    .X(net1111));
 sg13g2_dlygate4sd3_1 hold997 (.A(\u_toplayer.u_layer1.u_neuron.acc[11] ),
    .X(net1112));
 sg13g2_dlygate4sd3_1 hold998 (.A(\u_toplayer.u_layer3.u_neuron.din[6] ),
    .X(net1113));
 sg13g2_dlygate4sd3_1 hold999 (.A(\u_toplayer.u_layer2.u_neuron.acc[11] ),
    .X(net1114));
 sg13g2_dlygate4sd3_1 hold1000 (.A(\u_toplayer.u_outlayer.u_neuron.mult[15] ),
    .X(net1115));
 sg13g2_dlygate4sd3_1 hold1001 (.A(\u_toplayer.u_outlayer.u_neuron.acc[2] ),
    .X(net1116));
 sg13g2_dlygate4sd3_1 hold1002 (.A(\u_toplayer.u_layer1.u_neuron.acc[14] ),
    .X(net1117));
 sg13g2_dlygate4sd3_1 hold1003 (.A(\u_toplayer.u_outlayer.u_neuron.acc[6] ),
    .X(net1118));
 sg13g2_dlygate4sd3_1 hold1004 (.A(\u_toplayer.u_layer2.u_neuron.acc[23] ),
    .X(net1119));
 sg13g2_dlygate4sd3_1 hold1005 (.A(\u_toplayer.u_layer1.u_neuron.acc[19] ),
    .X(net1120));
 sg13g2_dlygate4sd3_1 hold1006 (.A(\u_toplayer.u_layer3.u_neuron.acc[21] ),
    .X(net1121));
 sg13g2_dlygate4sd3_1 hold1007 (.A(\u_toplayer.u_layer3.u_neuron.acc[4] ),
    .X(net1122));
 sg13g2_dlygate4sd3_1 hold1008 (.A(\u_toplayer.u_outlayer.u_neuron.din[2] ),
    .X(net1123));
 sg13g2_dlygate4sd3_1 hold1009 (.A(\u_toplayer.u_layer2.u_neuron.acc[21] ),
    .X(net1124));
 sg13g2_dlygate4sd3_1 hold1010 (.A(\u_toplayer.u_outlayer.u_neuron.din[0] ),
    .X(net1125));
 sg13g2_dlygate4sd3_1 hold1011 (.A(_00165_),
    .X(net1126));
 sg13g2_dlygate4sd3_1 hold1012 (.A(\u_toplayer.u_outlayer.u_neuron.acc[10] ),
    .X(net1127));
 sg13g2_dlygate4sd3_1 hold1013 (.A(\u_toplayer.u_layer3.u_neuron.mult[15] ),
    .X(net1128));
 sg13g2_dlygate4sd3_1 hold1014 (.A(\u_toplayer.u_layer2.statel2[4] ),
    .X(net1129));
 sg13g2_dlygate4sd3_1 hold1015 (.A(\u_toplayer.u_layer3.u_neuron.acc[6] ),
    .X(net1130));
 sg13g2_dlygate4sd3_1 hold1016 (.A(\u_toplayer.u_layer3.u_neuron.din[1] ),
    .X(net1131));
 sg13g2_dlygate4sd3_1 hold1017 (.A(\u_toplayer.u_layer2.u_neuron.acc[8] ),
    .X(net1132));
 sg13g2_dlygate4sd3_1 hold1018 (.A(\u_toplayer.u_layer1.u_neuron.acc[1] ),
    .X(net1133));
 sg13g2_dlygate4sd3_1 hold1019 (.A(\u_toplayer.u_layer2.u_neuron.instCtrl.state[2] ),
    .X(net1134));
 sg13g2_dlygate4sd3_1 hold1020 (.A(_00015_),
    .X(net1135));
 sg13g2_dlygate4sd3_1 hold1021 (.A(\u_toplayer.u_layer2.u_neuron.acc[7] ),
    .X(net1136));
 sg13g2_dlygate4sd3_1 hold1022 (.A(\u_toplayer.u_layer2.u_neuron.acc[4] ),
    .X(net1137));
 sg13g2_dlygate4sd3_1 hold1023 (.A(\u_toplayer.u_outlayer.u_neuron.din[3] ),
    .X(net1138));
 sg13g2_dlygate4sd3_1 hold1024 (.A(_00168_),
    .X(net1139));
 sg13g2_dlygate4sd3_1 hold1025 (.A(\u_toplayer.u_outlayer.u_neuron.acc[8] ),
    .X(net1140));
 sg13g2_dlygate4sd3_1 hold1026 (.A(\u_toplayer.u_layer2.u_neuron.din[2] ),
    .X(net1141));
 sg13g2_dlygate4sd3_1 hold1027 (.A(_00654_),
    .X(net1142));
 sg13g2_dlygate4sd3_1 hold1028 (.A(\u_toplayer.u_layer1.u_neuron.acc[6] ),
    .X(net1143));
 sg13g2_dlygate4sd3_1 hold1029 (.A(\u_toplayer.u_layer3.u_neuron.acc[11] ),
    .X(net1144));
 sg13g2_dlygate4sd3_1 hold1030 (.A(\u_toplayer.u_layer1.u_neuron.acc[10] ),
    .X(net1145));
 sg13g2_dlygate4sd3_1 hold1031 (.A(\u_toplayer.u_layer1.neuron_index[1] ),
    .X(net1146));
 sg13g2_dlygate4sd3_1 hold1032 (.A(_05235_),
    .X(net1147));
 sg13g2_dlygate4sd3_1 hold1033 (.A(\u_toplayer.u_outlayer.u_neuron.din[4] ),
    .X(net1148));
 sg13g2_dlygate4sd3_1 hold1034 (.A(\u_toplayer.u_layer2.neuron_index[1] ),
    .X(net1149));
 sg13g2_dlygate4sd3_1 hold1035 (.A(_03737_),
    .X(net1150));
 sg13g2_dlygate4sd3_1 hold1036 (.A(\u_toplayer.u_layer3.u_neuron.acc[9] ),
    .X(net1151));
 sg13g2_dlygate4sd3_1 hold1037 (.A(\u_toplayer.u_layer2.u_neuron.din[1] ),
    .X(net1152));
 sg13g2_dlygate4sd3_1 hold1038 (.A(\u_toplayer.u_layer1.u_neuron.acc[3] ),
    .X(net1153));
 sg13g2_dlygate4sd3_1 hold1039 (.A(\u_toplayer.u_layer1.u_neuron.acc[8] ),
    .X(net1154));
 sg13g2_dlygate4sd3_1 hold1040 (.A(\u_toplayer.u_outlayer.u_neuron.acc[14] ),
    .X(net1155));
 sg13g2_dlygate4sd3_1 hold1041 (.A(_00032_),
    .X(net1156));
 sg13g2_dlygate4sd3_1 hold1042 (.A(\u_toplayer.u_layer2.u_neuron.acc[3] ),
    .X(net1157));
 sg13g2_dlygate4sd3_1 hold1043 (.A(\u_toplayer.u_outlayer.u_neuron.acc[12] ),
    .X(net1158));
 sg13g2_dlygate4sd3_1 hold1044 (.A(\u_toplayer.u_layer2.u_neuron.acc[13] ),
    .X(net1159));
 sg13g2_dlygate4sd3_1 hold1045 (.A(\u_toplayer.u_layer2.u_neuron.din[4] ),
    .X(net1160));
 sg13g2_dlygate4sd3_1 hold1046 (.A(\u_toplayer.u_outlayer.u_neuron.acc[7] ),
    .X(net1161));
 sg13g2_dlygate4sd3_1 hold1047 (.A(_00204_),
    .X(net1162));
 sg13g2_dlygate4sd3_1 hold1048 (.A(\u_toplayer.u_layer3.u_neuron.acc[12] ),
    .X(net1163));
 sg13g2_dlygate4sd3_1 hold1049 (.A(\u_toplayer.u_layer2.u_neuron.acc[23] ),
    .X(net1164));
 sg13g2_dlygate4sd3_1 hold1050 (.A(\u_toplayer.u_layer1.u_neuron.acc[12] ),
    .X(net1165));
 sg13g2_dlygate4sd3_1 hold1051 (.A(\u_toplayer.u_layer3.u_neuron.din[2] ),
    .X(net1166));
 sg13g2_dlygate4sd3_1 hold1052 (.A(\u_toplayer.u_layer3.u_neuron.acc[14] ),
    .X(net1167));
 sg13g2_dlygate4sd3_1 hold1053 (.A(\u_toplayer.u_layer2.u_neuron.acc[18] ),
    .X(net1168));
 sg13g2_dlygate4sd3_1 hold1054 (.A(_00695_),
    .X(net1169));
 sg13g2_dlygate4sd3_1 hold1055 (.A(\u_toplayer.u_outlayer.u_neuron.acc[4] ),
    .X(net1170));
 sg13g2_dlygate4sd3_1 hold1056 (.A(\u_toplayer.u_layer3.u_neuron.acc[10] ),
    .X(net1171));
 sg13g2_dlygate4sd3_1 hold1057 (.A(\u_toplayer.u_layer1.u_neuron.acc[4] ),
    .X(net1172));
 sg13g2_dlygate4sd3_1 hold1058 (.A(\u_toplayer.u_layer2.u_neuron.acc[15] ),
    .X(net1173));
 sg13g2_dlygate4sd3_1 hold1059 (.A(\u_toplayer.delayed_done_layer1 ),
    .X(net1174));
 sg13g2_dlygate4sd3_1 hold1060 (.A(_00013_),
    .X(net1175));
 sg13g2_dlygate4sd3_1 hold1061 (.A(\u_toplayer.u_layer2.u_neuron.acc[2] ),
    .X(net1176));
 sg13g2_dlygate4sd3_1 hold1062 (.A(\u_toplayer.u_layer3.u_neuron.din[7] ),
    .X(net1177));
 sg13g2_dlygate4sd3_1 hold1063 (.A(\u_toplayer.u_layer3.u_neuron.instCtrl.state[4] ),
    .X(net1178));
 sg13g2_dlygate4sd3_1 hold1064 (.A(\u_toplayer.u_layer3.u_neuron.acc[18] ),
    .X(net1179));
 sg13g2_dlygate4sd3_1 hold1065 (.A(\u_toplayer.u_layer1.u_neuron.acc[9] ),
    .X(net1180));
 sg13g2_dlygate4sd3_1 hold1066 (.A(\u_toplayer.u_layer1.u_neuron.acc[7] ),
    .X(net1181));
 sg13g2_dlygate4sd3_1 hold1067 (.A(\u_toplayer.u_layer2.u_neuron.acc[10] ),
    .X(net1182));
 sg13g2_dlygate4sd3_1 hold1068 (.A(\u_toplayer.u_layer3.u_neuron.acc[5] ),
    .X(net1183));
 sg13g2_dlygate4sd3_1 hold1069 (.A(\u_toplayer.u_outlayer.u_neuron.acc[9] ),
    .X(net1184));
 sg13g2_dlygate4sd3_1 hold1070 (.A(\u_toplayer.u_layer1.u_neuron.acc[20] ),
    .X(net1185));
 sg13g2_dlygate4sd3_1 hold1071 (.A(\u_toplayer.u_layer2.u_neuron.din[0] ),
    .X(net1186));
 sg13g2_dlygate4sd3_1 hold1072 (.A(\u_toplayer.u_layer2.u_neuron.din[3] ),
    .X(net1187));
 sg13g2_dlygate4sd3_1 hold1073 (.A(\u_toplayer.u_layer1.u_neuron.b[7] ),
    .X(net1188));
 sg13g2_dlygate4sd3_1 hold1074 (.A(\u_toplayer.u_layer2.u_neuron.acc[14] ),
    .X(net1189));
 sg13g2_dlygate4sd3_1 hold1075 (.A(\u_toplayer.u_layer3.neuron_index[3] ),
    .X(net1190));
 sg13g2_dlygate4sd3_1 hold1076 (.A(_00224_),
    .X(net1191));
 sg13g2_dlygate4sd3_1 hold1077 (.A(\u_toplayer.u_layer1.u_neuron.acc[5] ),
    .X(net1192));
 sg13g2_dlygate4sd3_1 hold1078 (.A(\u_toplayer.delayed_done_layer3 ),
    .X(net1193));
 sg13g2_dlygate4sd3_1 hold1079 (.A(\u_toplayer.u_layer2.u_neuron.acc[16] ),
    .X(net1194));
 sg13g2_dlygate4sd3_1 hold1080 (.A(\u_toplayer.u_layer2.u_neuron.acc[12] ),
    .X(net1195));
 sg13g2_dlygate4sd3_1 hold1081 (.A(\u_toplayer.u_outlayer.u_neuron.acc[18] ),
    .X(net1196));
 sg13g2_dlygate4sd3_1 hold1082 (.A(\u_toplayer.u_layer2.u_neuron.din[5] ),
    .X(net1197));
 sg13g2_dlygate4sd3_1 hold1083 (.A(\u_toplayer.u_layer1.u_neuron.acc[13] ),
    .X(net1198));
 sg13g2_dlygate4sd3_1 hold1084 (.A(\u_toplayer.u_outlayer.u_neuron.mult[13] ),
    .X(net1199));
 sg13g2_dlygate4sd3_1 hold1085 (.A(\u_toplayer.u_outlayer.u_neuron.mult[14] ),
    .X(net1200));
 sg13g2_dlygate4sd3_1 hold1086 (.A(\u_toplayer.u_outlayer.u_neuron.acc[13] ),
    .X(net1201));
 sg13g2_dlygate4sd3_1 hold1087 (.A(\u_toplayer.u_outlayer.u_neuron.acc[5] ),
    .X(net1202));
 sg13g2_dlygate4sd3_1 hold1088 (.A(\u_toplayer.u_layer2.u_neuron.acc[20] ),
    .X(net1203));
 sg13g2_dlygate4sd3_1 hold1089 (.A(\u_toplayer.u_layer1.u_neuron.acc[18] ),
    .X(net1204));
 sg13g2_dlygate4sd3_1 hold1090 (.A(\u_toplayer.u_layer2.sum[1] ),
    .X(net1205));
 sg13g2_dlygate4sd3_1 hold1091 (.A(\u_toplayer.u_layer3.u_neuron.acc[7] ),
    .X(net1206));
 sg13g2_dlygate4sd3_1 hold1092 (.A(\u_toplayer.u_layer2.u_neuron.din[6] ),
    .X(net1207));
 sg13g2_dlygate4sd3_1 hold1093 (.A(\u_toplayer.u_outlayer.u_neuron.acc[20] ),
    .X(net1208));
 sg13g2_dlygate4sd3_1 hold1094 (.A(\u_toplayer.u_layer1.u_neuron.mult[15] ),
    .X(net1209));
 sg13g2_dlygate4sd3_1 hold1095 (.A(\u_toplayer.u_layer1.neuron_index[4] ),
    .X(net1210));
 sg13g2_dlygate4sd3_1 hold1096 (.A(\u_toplayer.u_layer3.neuron_index[1] ),
    .X(net1211));
 sg13g2_dlygate4sd3_1 hold1097 (.A(\u_toplayer.u_outlayer.u_neuron.mult[0] ),
    .X(net1212));
 sg13g2_antennanp ANTENNA_1 (.A(_03375_));
 sg13g2_antennanp ANTENNA_2 (.A(_03375_));
 sg13g2_antennanp ANTENNA_3 (.A(clk));
 sg13g2_antennanp ANTENNA_4 (.A(clk));
 sg13g2_antennanp ANTENNA_5 (.A(clk));
 sg13g2_antennanp ANTENNA_6 (.A(clk));
 sg13g2_antennanp ANTENNA_7 (.A(uio_in[6]));
 sg13g2_antennanp ANTENNA_8 (.A(uio_in[7]));
 sg13g2_antennanp ANTENNA_9 (.A(uio_in[7]));
 sg13g2_antennanp ANTENNA_10 (.A(net3487));
 sg13g2_antennanp ANTENNA_11 (.A(net3487));
 sg13g2_antennanp ANTENNA_12 (.A(net3487));
 sg13g2_antennanp ANTENNA_13 (.A(net3487));
 sg13g2_antennanp ANTENNA_14 (.A(net3487));
 sg13g2_antennanp ANTENNA_15 (.A(net3487));
 sg13g2_antennanp ANTENNA_16 (.A(net3487));
 sg13g2_antennanp ANTENNA_17 (.A(net3487));
 sg13g2_antennanp ANTENNA_18 (.A(net3487));
 sg13g2_antennanp ANTENNA_19 (.A(net3487));
 sg13g2_antennanp ANTENNA_20 (.A(net3487));
 sg13g2_antennanp ANTENNA_21 (.A(net3487));
 sg13g2_antennanp ANTENNA_22 (.A(net3487));
 sg13g2_antennanp ANTENNA_23 (.A(clk));
 sg13g2_antennanp ANTENNA_24 (.A(clk));
 sg13g2_antennanp ANTENNA_25 (.A(clk));
 sg13g2_antennanp ANTENNA_26 (.A(clk));
 sg13g2_antennanp ANTENNA_27 (.A(uio_in[6]));
 sg13g2_antennanp ANTENNA_28 (.A(uio_in[7]));
 sg13g2_antennanp ANTENNA_29 (.A(uio_in[7]));
 sg13g2_antennanp ANTENNA_30 (.A(clk));
 sg13g2_antennanp ANTENNA_31 (.A(clk));
 sg13g2_antennanp ANTENNA_32 (.A(clk));
 sg13g2_antennanp ANTENNA_33 (.A(clk));
 sg13g2_antennanp ANTENNA_34 (.A(uio_in[6]));
 sg13g2_antennanp ANTENNA_35 (.A(uio_in[7]));
 sg13g2_antennanp ANTENNA_36 (.A(uio_in[7]));
 sg13g2_antennanp ANTENNA_37 (.A(net3487));
 sg13g2_antennanp ANTENNA_38 (.A(net3487));
 sg13g2_antennanp ANTENNA_39 (.A(net3487));
 sg13g2_antennanp ANTENNA_40 (.A(net3487));
 sg13g2_antennanp ANTENNA_41 (.A(net3487));
 sg13g2_antennanp ANTENNA_42 (.A(net3487));
 sg13g2_antennanp ANTENNA_43 (.A(net3487));
 sg13g2_antennanp ANTENNA_44 (.A(net3487));
 sg13g2_antennanp ANTENNA_45 (.A(net3487));
 sg13g2_antennanp ANTENNA_46 (.A(net3487));
 sg13g2_antennanp ANTENNA_47 (.A(net3487));
 sg13g2_antennanp ANTENNA_48 (.A(net3487));
 sg13g2_antennanp ANTENNA_49 (.A(net3487));
 sg13g2_antennanp ANTENNA_50 (.A(net3487));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_fill_2 FILLER_0_378 ();
 sg13g2_fill_1 FILLER_0_380 ();
 sg13g2_fill_2 FILLER_0_386 ();
 sg13g2_fill_1 FILLER_0_388 ();
 sg13g2_fill_2 FILLER_0_435 ();
 sg13g2_fill_1 FILLER_0_437 ();
 sg13g2_fill_2 FILLER_0_506 ();
 sg13g2_fill_1 FILLER_0_508 ();
 sg13g2_fill_2 FILLER_0_579 ();
 sg13g2_decap_8 FILLER_0_624 ();
 sg13g2_decap_8 FILLER_0_631 ();
 sg13g2_decap_8 FILLER_0_638 ();
 sg13g2_decap_8 FILLER_0_645 ();
 sg13g2_decap_8 FILLER_0_652 ();
 sg13g2_decap_8 FILLER_0_659 ();
 sg13g2_decap_8 FILLER_0_666 ();
 sg13g2_decap_8 FILLER_0_673 ();
 sg13g2_decap_8 FILLER_0_680 ();
 sg13g2_decap_8 FILLER_0_687 ();
 sg13g2_decap_8 FILLER_0_694 ();
 sg13g2_decap_8 FILLER_0_701 ();
 sg13g2_decap_8 FILLER_0_708 ();
 sg13g2_decap_8 FILLER_0_715 ();
 sg13g2_fill_2 FILLER_0_722 ();
 sg13g2_decap_4 FILLER_0_750 ();
 sg13g2_decap_8 FILLER_0_806 ();
 sg13g2_decap_8 FILLER_0_813 ();
 sg13g2_decap_8 FILLER_0_820 ();
 sg13g2_decap_8 FILLER_0_827 ();
 sg13g2_decap_8 FILLER_0_834 ();
 sg13g2_decap_8 FILLER_0_841 ();
 sg13g2_decap_8 FILLER_0_848 ();
 sg13g2_decap_8 FILLER_0_855 ();
 sg13g2_decap_8 FILLER_0_862 ();
 sg13g2_decap_8 FILLER_0_869 ();
 sg13g2_decap_8 FILLER_0_876 ();
 sg13g2_decap_8 FILLER_0_883 ();
 sg13g2_decap_8 FILLER_0_890 ();
 sg13g2_decap_8 FILLER_0_897 ();
 sg13g2_decap_8 FILLER_0_904 ();
 sg13g2_decap_8 FILLER_0_911 ();
 sg13g2_decap_8 FILLER_0_918 ();
 sg13g2_decap_8 FILLER_0_925 ();
 sg13g2_decap_8 FILLER_0_932 ();
 sg13g2_decap_8 FILLER_0_939 ();
 sg13g2_decap_8 FILLER_0_946 ();
 sg13g2_decap_8 FILLER_0_953 ();
 sg13g2_decap_8 FILLER_0_960 ();
 sg13g2_decap_8 FILLER_0_967 ();
 sg13g2_decap_8 FILLER_0_974 ();
 sg13g2_decap_8 FILLER_0_981 ();
 sg13g2_decap_8 FILLER_0_988 ();
 sg13g2_decap_8 FILLER_0_995 ();
 sg13g2_decap_8 FILLER_0_1002 ();
 sg13g2_decap_8 FILLER_0_1009 ();
 sg13g2_decap_8 FILLER_0_1016 ();
 sg13g2_decap_8 FILLER_0_1023 ();
 sg13g2_decap_8 FILLER_0_1030 ();
 sg13g2_decap_8 FILLER_0_1037 ();
 sg13g2_decap_8 FILLER_0_1044 ();
 sg13g2_decap_8 FILLER_0_1051 ();
 sg13g2_decap_8 FILLER_0_1058 ();
 sg13g2_decap_8 FILLER_0_1065 ();
 sg13g2_decap_8 FILLER_0_1072 ();
 sg13g2_decap_8 FILLER_0_1079 ();
 sg13g2_decap_8 FILLER_0_1086 ();
 sg13g2_decap_8 FILLER_0_1093 ();
 sg13g2_decap_8 FILLER_0_1100 ();
 sg13g2_decap_8 FILLER_0_1107 ();
 sg13g2_decap_8 FILLER_0_1114 ();
 sg13g2_decap_8 FILLER_0_1121 ();
 sg13g2_decap_8 FILLER_0_1128 ();
 sg13g2_decap_8 FILLER_0_1135 ();
 sg13g2_decap_8 FILLER_0_1142 ();
 sg13g2_decap_8 FILLER_0_1149 ();
 sg13g2_decap_8 FILLER_0_1156 ();
 sg13g2_decap_8 FILLER_0_1163 ();
 sg13g2_decap_8 FILLER_0_1170 ();
 sg13g2_decap_8 FILLER_0_1177 ();
 sg13g2_decap_8 FILLER_0_1184 ();
 sg13g2_decap_8 FILLER_0_1191 ();
 sg13g2_decap_8 FILLER_0_1198 ();
 sg13g2_decap_8 FILLER_0_1205 ();
 sg13g2_decap_8 FILLER_0_1212 ();
 sg13g2_decap_8 FILLER_0_1219 ();
 sg13g2_decap_8 FILLER_0_1226 ();
 sg13g2_decap_8 FILLER_0_1233 ();
 sg13g2_decap_8 FILLER_0_1240 ();
 sg13g2_decap_8 FILLER_0_1247 ();
 sg13g2_decap_8 FILLER_0_1254 ();
 sg13g2_decap_8 FILLER_0_1261 ();
 sg13g2_decap_8 FILLER_0_1268 ();
 sg13g2_decap_8 FILLER_0_1275 ();
 sg13g2_decap_8 FILLER_0_1282 ();
 sg13g2_decap_8 FILLER_0_1289 ();
 sg13g2_decap_8 FILLER_0_1296 ();
 sg13g2_decap_8 FILLER_0_1303 ();
 sg13g2_decap_8 FILLER_0_1310 ();
 sg13g2_decap_8 FILLER_0_1317 ();
 sg13g2_decap_8 FILLER_0_1324 ();
 sg13g2_decap_8 FILLER_0_1331 ();
 sg13g2_decap_8 FILLER_0_1338 ();
 sg13g2_decap_8 FILLER_0_1345 ();
 sg13g2_decap_8 FILLER_0_1352 ();
 sg13g2_decap_8 FILLER_0_1359 ();
 sg13g2_decap_8 FILLER_0_1366 ();
 sg13g2_decap_8 FILLER_0_1373 ();
 sg13g2_decap_8 FILLER_0_1380 ();
 sg13g2_decap_8 FILLER_0_1387 ();
 sg13g2_decap_8 FILLER_0_1394 ();
 sg13g2_decap_8 FILLER_0_1401 ();
 sg13g2_decap_8 FILLER_0_1408 ();
 sg13g2_decap_8 FILLER_0_1415 ();
 sg13g2_decap_8 FILLER_0_1422 ();
 sg13g2_decap_8 FILLER_0_1429 ();
 sg13g2_decap_8 FILLER_0_1436 ();
 sg13g2_decap_8 FILLER_0_1443 ();
 sg13g2_decap_8 FILLER_0_1450 ();
 sg13g2_decap_8 FILLER_0_1457 ();
 sg13g2_decap_8 FILLER_0_1464 ();
 sg13g2_decap_8 FILLER_0_1471 ();
 sg13g2_decap_8 FILLER_0_1478 ();
 sg13g2_decap_8 FILLER_0_1485 ();
 sg13g2_decap_8 FILLER_0_1492 ();
 sg13g2_decap_8 FILLER_0_1499 ();
 sg13g2_decap_8 FILLER_0_1506 ();
 sg13g2_decap_8 FILLER_0_1513 ();
 sg13g2_decap_8 FILLER_0_1520 ();
 sg13g2_decap_8 FILLER_0_1527 ();
 sg13g2_decap_8 FILLER_0_1534 ();
 sg13g2_decap_8 FILLER_0_1541 ();
 sg13g2_decap_8 FILLER_0_1548 ();
 sg13g2_decap_8 FILLER_0_1555 ();
 sg13g2_decap_8 FILLER_0_1562 ();
 sg13g2_decap_8 FILLER_0_1569 ();
 sg13g2_decap_8 FILLER_0_1576 ();
 sg13g2_decap_8 FILLER_0_1583 ();
 sg13g2_decap_8 FILLER_0_1590 ();
 sg13g2_decap_8 FILLER_0_1597 ();
 sg13g2_decap_8 FILLER_0_1604 ();
 sg13g2_decap_8 FILLER_0_1611 ();
 sg13g2_decap_8 FILLER_0_1618 ();
 sg13g2_decap_8 FILLER_0_1625 ();
 sg13g2_decap_8 FILLER_0_1632 ();
 sg13g2_decap_8 FILLER_0_1639 ();
 sg13g2_decap_8 FILLER_0_1646 ();
 sg13g2_decap_8 FILLER_0_1653 ();
 sg13g2_decap_8 FILLER_0_1660 ();
 sg13g2_decap_8 FILLER_0_1667 ();
 sg13g2_decap_8 FILLER_0_1674 ();
 sg13g2_decap_8 FILLER_0_1681 ();
 sg13g2_decap_8 FILLER_0_1688 ();
 sg13g2_decap_8 FILLER_0_1695 ();
 sg13g2_decap_8 FILLER_0_1702 ();
 sg13g2_decap_8 FILLER_0_1709 ();
 sg13g2_decap_8 FILLER_0_1716 ();
 sg13g2_decap_8 FILLER_0_1723 ();
 sg13g2_decap_8 FILLER_0_1730 ();
 sg13g2_decap_8 FILLER_0_1737 ();
 sg13g2_decap_8 FILLER_0_1744 ();
 sg13g2_decap_8 FILLER_0_1751 ();
 sg13g2_decap_8 FILLER_0_1758 ();
 sg13g2_fill_2 FILLER_0_1765 ();
 sg13g2_fill_1 FILLER_0_1767 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_fill_2 FILLER_1_308 ();
 sg13g2_fill_1 FILLER_1_349 ();
 sg13g2_fill_2 FILLER_1_408 ();
 sg13g2_fill_1 FILLER_1_476 ();
 sg13g2_fill_1 FILLER_1_486 ();
 sg13g2_fill_1 FILLER_1_553 ();
 sg13g2_fill_1 FILLER_1_563 ();
 sg13g2_fill_1 FILLER_1_578 ();
 sg13g2_decap_8 FILLER_1_634 ();
 sg13g2_decap_8 FILLER_1_641 ();
 sg13g2_decap_8 FILLER_1_648 ();
 sg13g2_decap_8 FILLER_1_655 ();
 sg13g2_decap_8 FILLER_1_662 ();
 sg13g2_decap_8 FILLER_1_669 ();
 sg13g2_decap_8 FILLER_1_676 ();
 sg13g2_decap_8 FILLER_1_683 ();
 sg13g2_decap_8 FILLER_1_690 ();
 sg13g2_decap_8 FILLER_1_697 ();
 sg13g2_decap_8 FILLER_1_704 ();
 sg13g2_fill_2 FILLER_1_711 ();
 sg13g2_fill_1 FILLER_1_713 ();
 sg13g2_fill_2 FILLER_1_776 ();
 sg13g2_fill_1 FILLER_1_778 ();
 sg13g2_decap_8 FILLER_1_811 ();
 sg13g2_decap_8 FILLER_1_818 ();
 sg13g2_decap_8 FILLER_1_825 ();
 sg13g2_decap_8 FILLER_1_832 ();
 sg13g2_decap_8 FILLER_1_839 ();
 sg13g2_decap_8 FILLER_1_846 ();
 sg13g2_decap_8 FILLER_1_853 ();
 sg13g2_decap_8 FILLER_1_860 ();
 sg13g2_decap_8 FILLER_1_867 ();
 sg13g2_decap_8 FILLER_1_874 ();
 sg13g2_decap_8 FILLER_1_881 ();
 sg13g2_decap_8 FILLER_1_888 ();
 sg13g2_decap_8 FILLER_1_895 ();
 sg13g2_decap_8 FILLER_1_902 ();
 sg13g2_decap_8 FILLER_1_909 ();
 sg13g2_decap_8 FILLER_1_916 ();
 sg13g2_decap_8 FILLER_1_923 ();
 sg13g2_decap_8 FILLER_1_930 ();
 sg13g2_decap_8 FILLER_1_937 ();
 sg13g2_decap_8 FILLER_1_944 ();
 sg13g2_decap_8 FILLER_1_951 ();
 sg13g2_decap_8 FILLER_1_958 ();
 sg13g2_decap_8 FILLER_1_965 ();
 sg13g2_decap_8 FILLER_1_972 ();
 sg13g2_decap_8 FILLER_1_979 ();
 sg13g2_decap_8 FILLER_1_986 ();
 sg13g2_decap_8 FILLER_1_993 ();
 sg13g2_decap_8 FILLER_1_1000 ();
 sg13g2_decap_8 FILLER_1_1007 ();
 sg13g2_decap_8 FILLER_1_1014 ();
 sg13g2_decap_8 FILLER_1_1021 ();
 sg13g2_decap_8 FILLER_1_1028 ();
 sg13g2_decap_8 FILLER_1_1035 ();
 sg13g2_decap_8 FILLER_1_1042 ();
 sg13g2_decap_8 FILLER_1_1049 ();
 sg13g2_decap_8 FILLER_1_1056 ();
 sg13g2_decap_8 FILLER_1_1063 ();
 sg13g2_decap_8 FILLER_1_1070 ();
 sg13g2_decap_8 FILLER_1_1077 ();
 sg13g2_decap_8 FILLER_1_1084 ();
 sg13g2_decap_8 FILLER_1_1091 ();
 sg13g2_decap_8 FILLER_1_1098 ();
 sg13g2_decap_8 FILLER_1_1105 ();
 sg13g2_decap_8 FILLER_1_1112 ();
 sg13g2_decap_8 FILLER_1_1119 ();
 sg13g2_decap_8 FILLER_1_1126 ();
 sg13g2_decap_8 FILLER_1_1133 ();
 sg13g2_decap_8 FILLER_1_1140 ();
 sg13g2_decap_8 FILLER_1_1147 ();
 sg13g2_decap_8 FILLER_1_1154 ();
 sg13g2_decap_8 FILLER_1_1161 ();
 sg13g2_decap_8 FILLER_1_1168 ();
 sg13g2_decap_8 FILLER_1_1175 ();
 sg13g2_decap_8 FILLER_1_1182 ();
 sg13g2_decap_8 FILLER_1_1189 ();
 sg13g2_decap_8 FILLER_1_1196 ();
 sg13g2_decap_8 FILLER_1_1203 ();
 sg13g2_decap_8 FILLER_1_1210 ();
 sg13g2_decap_8 FILLER_1_1217 ();
 sg13g2_decap_8 FILLER_1_1224 ();
 sg13g2_decap_8 FILLER_1_1231 ();
 sg13g2_decap_8 FILLER_1_1238 ();
 sg13g2_decap_8 FILLER_1_1245 ();
 sg13g2_decap_8 FILLER_1_1252 ();
 sg13g2_decap_8 FILLER_1_1259 ();
 sg13g2_decap_8 FILLER_1_1266 ();
 sg13g2_decap_8 FILLER_1_1273 ();
 sg13g2_decap_8 FILLER_1_1280 ();
 sg13g2_decap_8 FILLER_1_1287 ();
 sg13g2_decap_8 FILLER_1_1294 ();
 sg13g2_decap_8 FILLER_1_1301 ();
 sg13g2_decap_8 FILLER_1_1308 ();
 sg13g2_decap_8 FILLER_1_1315 ();
 sg13g2_decap_8 FILLER_1_1322 ();
 sg13g2_decap_8 FILLER_1_1329 ();
 sg13g2_decap_8 FILLER_1_1336 ();
 sg13g2_decap_8 FILLER_1_1343 ();
 sg13g2_decap_8 FILLER_1_1350 ();
 sg13g2_decap_8 FILLER_1_1357 ();
 sg13g2_decap_8 FILLER_1_1364 ();
 sg13g2_decap_8 FILLER_1_1371 ();
 sg13g2_decap_8 FILLER_1_1378 ();
 sg13g2_decap_8 FILLER_1_1385 ();
 sg13g2_decap_8 FILLER_1_1392 ();
 sg13g2_decap_8 FILLER_1_1399 ();
 sg13g2_decap_8 FILLER_1_1406 ();
 sg13g2_decap_8 FILLER_1_1413 ();
 sg13g2_decap_8 FILLER_1_1420 ();
 sg13g2_decap_8 FILLER_1_1427 ();
 sg13g2_decap_8 FILLER_1_1434 ();
 sg13g2_decap_8 FILLER_1_1441 ();
 sg13g2_decap_8 FILLER_1_1448 ();
 sg13g2_decap_8 FILLER_1_1455 ();
 sg13g2_decap_8 FILLER_1_1462 ();
 sg13g2_decap_8 FILLER_1_1469 ();
 sg13g2_decap_8 FILLER_1_1476 ();
 sg13g2_decap_8 FILLER_1_1483 ();
 sg13g2_decap_8 FILLER_1_1490 ();
 sg13g2_decap_8 FILLER_1_1497 ();
 sg13g2_decap_8 FILLER_1_1504 ();
 sg13g2_decap_8 FILLER_1_1511 ();
 sg13g2_decap_8 FILLER_1_1518 ();
 sg13g2_decap_8 FILLER_1_1525 ();
 sg13g2_decap_8 FILLER_1_1532 ();
 sg13g2_decap_8 FILLER_1_1539 ();
 sg13g2_decap_8 FILLER_1_1546 ();
 sg13g2_decap_8 FILLER_1_1553 ();
 sg13g2_decap_8 FILLER_1_1560 ();
 sg13g2_decap_8 FILLER_1_1567 ();
 sg13g2_decap_8 FILLER_1_1574 ();
 sg13g2_decap_8 FILLER_1_1581 ();
 sg13g2_decap_8 FILLER_1_1588 ();
 sg13g2_decap_8 FILLER_1_1595 ();
 sg13g2_decap_8 FILLER_1_1602 ();
 sg13g2_decap_8 FILLER_1_1609 ();
 sg13g2_decap_8 FILLER_1_1616 ();
 sg13g2_decap_8 FILLER_1_1623 ();
 sg13g2_decap_8 FILLER_1_1630 ();
 sg13g2_decap_8 FILLER_1_1637 ();
 sg13g2_decap_8 FILLER_1_1644 ();
 sg13g2_decap_8 FILLER_1_1651 ();
 sg13g2_decap_8 FILLER_1_1658 ();
 sg13g2_decap_8 FILLER_1_1665 ();
 sg13g2_decap_8 FILLER_1_1672 ();
 sg13g2_decap_8 FILLER_1_1679 ();
 sg13g2_decap_8 FILLER_1_1686 ();
 sg13g2_decap_8 FILLER_1_1693 ();
 sg13g2_decap_8 FILLER_1_1700 ();
 sg13g2_decap_8 FILLER_1_1707 ();
 sg13g2_decap_8 FILLER_1_1714 ();
 sg13g2_decap_8 FILLER_1_1721 ();
 sg13g2_decap_8 FILLER_1_1728 ();
 sg13g2_decap_8 FILLER_1_1735 ();
 sg13g2_decap_8 FILLER_1_1742 ();
 sg13g2_decap_8 FILLER_1_1749 ();
 sg13g2_decap_8 FILLER_1_1756 ();
 sg13g2_decap_4 FILLER_1_1763 ();
 sg13g2_fill_1 FILLER_1_1767 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_4 FILLER_2_210 ();
 sg13g2_fill_1 FILLER_2_214 ();
 sg13g2_decap_8 FILLER_2_233 ();
 sg13g2_fill_2 FILLER_2_240 ();
 sg13g2_fill_1 FILLER_2_242 ();
 sg13g2_decap_8 FILLER_2_253 ();
 sg13g2_decap_8 FILLER_2_260 ();
 sg13g2_decap_8 FILLER_2_267 ();
 sg13g2_decap_8 FILLER_2_274 ();
 sg13g2_decap_8 FILLER_2_281 ();
 sg13g2_decap_8 FILLER_2_288 ();
 sg13g2_decap_4 FILLER_2_295 ();
 sg13g2_fill_1 FILLER_2_299 ();
 sg13g2_fill_2 FILLER_2_358 ();
 sg13g2_fill_1 FILLER_2_360 ();
 sg13g2_fill_2 FILLER_2_370 ();
 sg13g2_fill_1 FILLER_2_372 ();
 sg13g2_fill_1 FILLER_2_442 ();
 sg13g2_fill_2 FILLER_2_448 ();
 sg13g2_fill_1 FILLER_2_450 ();
 sg13g2_fill_2 FILLER_2_483 ();
 sg13g2_fill_1 FILLER_2_507 ();
 sg13g2_fill_2 FILLER_2_522 ();
 sg13g2_fill_1 FILLER_2_524 ();
 sg13g2_decap_8 FILLER_2_639 ();
 sg13g2_decap_8 FILLER_2_646 ();
 sg13g2_decap_8 FILLER_2_653 ();
 sg13g2_decap_8 FILLER_2_660 ();
 sg13g2_decap_8 FILLER_2_667 ();
 sg13g2_decap_8 FILLER_2_674 ();
 sg13g2_decap_8 FILLER_2_681 ();
 sg13g2_decap_8 FILLER_2_688 ();
 sg13g2_fill_2 FILLER_2_695 ();
 sg13g2_fill_2 FILLER_2_723 ();
 sg13g2_fill_1 FILLER_2_725 ();
 sg13g2_fill_1 FILLER_2_735 ();
 sg13g2_decap_8 FILLER_2_812 ();
 sg13g2_decap_8 FILLER_2_819 ();
 sg13g2_decap_8 FILLER_2_826 ();
 sg13g2_decap_8 FILLER_2_833 ();
 sg13g2_decap_8 FILLER_2_840 ();
 sg13g2_decap_8 FILLER_2_847 ();
 sg13g2_decap_8 FILLER_2_854 ();
 sg13g2_decap_8 FILLER_2_861 ();
 sg13g2_fill_2 FILLER_2_868 ();
 sg13g2_decap_8 FILLER_2_878 ();
 sg13g2_decap_8 FILLER_2_885 ();
 sg13g2_decap_8 FILLER_2_892 ();
 sg13g2_decap_8 FILLER_2_899 ();
 sg13g2_decap_8 FILLER_2_906 ();
 sg13g2_decap_8 FILLER_2_913 ();
 sg13g2_decap_8 FILLER_2_934 ();
 sg13g2_decap_4 FILLER_2_941 ();
 sg13g2_decap_8 FILLER_2_948 ();
 sg13g2_decap_8 FILLER_2_955 ();
 sg13g2_decap_8 FILLER_2_962 ();
 sg13g2_decap_8 FILLER_2_969 ();
 sg13g2_decap_8 FILLER_2_976 ();
 sg13g2_decap_8 FILLER_2_983 ();
 sg13g2_decap_8 FILLER_2_990 ();
 sg13g2_fill_1 FILLER_2_997 ();
 sg13g2_decap_4 FILLER_2_1037 ();
 sg13g2_decap_8 FILLER_2_1045 ();
 sg13g2_decap_8 FILLER_2_1052 ();
 sg13g2_decap_8 FILLER_2_1059 ();
 sg13g2_decap_8 FILLER_2_1066 ();
 sg13g2_decap_8 FILLER_2_1073 ();
 sg13g2_decap_8 FILLER_2_1080 ();
 sg13g2_fill_2 FILLER_2_1087 ();
 sg13g2_decap_8 FILLER_2_1093 ();
 sg13g2_decap_8 FILLER_2_1100 ();
 sg13g2_decap_8 FILLER_2_1107 ();
 sg13g2_decap_8 FILLER_2_1114 ();
 sg13g2_decap_8 FILLER_2_1121 ();
 sg13g2_decap_8 FILLER_2_1128 ();
 sg13g2_decap_8 FILLER_2_1135 ();
 sg13g2_decap_8 FILLER_2_1142 ();
 sg13g2_decap_8 FILLER_2_1149 ();
 sg13g2_decap_8 FILLER_2_1156 ();
 sg13g2_decap_8 FILLER_2_1163 ();
 sg13g2_decap_8 FILLER_2_1170 ();
 sg13g2_decap_8 FILLER_2_1177 ();
 sg13g2_decap_8 FILLER_2_1184 ();
 sg13g2_decap_8 FILLER_2_1191 ();
 sg13g2_decap_8 FILLER_2_1198 ();
 sg13g2_decap_8 FILLER_2_1205 ();
 sg13g2_decap_8 FILLER_2_1212 ();
 sg13g2_decap_8 FILLER_2_1219 ();
 sg13g2_decap_8 FILLER_2_1226 ();
 sg13g2_decap_8 FILLER_2_1233 ();
 sg13g2_decap_8 FILLER_2_1240 ();
 sg13g2_decap_8 FILLER_2_1247 ();
 sg13g2_decap_8 FILLER_2_1254 ();
 sg13g2_decap_8 FILLER_2_1261 ();
 sg13g2_decap_8 FILLER_2_1268 ();
 sg13g2_decap_8 FILLER_2_1275 ();
 sg13g2_decap_8 FILLER_2_1282 ();
 sg13g2_decap_8 FILLER_2_1289 ();
 sg13g2_decap_8 FILLER_2_1296 ();
 sg13g2_decap_8 FILLER_2_1303 ();
 sg13g2_decap_8 FILLER_2_1310 ();
 sg13g2_decap_8 FILLER_2_1317 ();
 sg13g2_decap_8 FILLER_2_1324 ();
 sg13g2_decap_8 FILLER_2_1331 ();
 sg13g2_decap_8 FILLER_2_1338 ();
 sg13g2_decap_8 FILLER_2_1345 ();
 sg13g2_decap_8 FILLER_2_1352 ();
 sg13g2_decap_8 FILLER_2_1359 ();
 sg13g2_decap_8 FILLER_2_1366 ();
 sg13g2_decap_8 FILLER_2_1373 ();
 sg13g2_decap_8 FILLER_2_1380 ();
 sg13g2_decap_8 FILLER_2_1387 ();
 sg13g2_decap_8 FILLER_2_1394 ();
 sg13g2_decap_8 FILLER_2_1401 ();
 sg13g2_decap_8 FILLER_2_1408 ();
 sg13g2_decap_8 FILLER_2_1415 ();
 sg13g2_decap_8 FILLER_2_1422 ();
 sg13g2_decap_8 FILLER_2_1429 ();
 sg13g2_decap_8 FILLER_2_1436 ();
 sg13g2_decap_8 FILLER_2_1443 ();
 sg13g2_decap_8 FILLER_2_1450 ();
 sg13g2_decap_8 FILLER_2_1457 ();
 sg13g2_decap_8 FILLER_2_1464 ();
 sg13g2_decap_8 FILLER_2_1471 ();
 sg13g2_decap_8 FILLER_2_1478 ();
 sg13g2_decap_8 FILLER_2_1485 ();
 sg13g2_decap_8 FILLER_2_1492 ();
 sg13g2_decap_8 FILLER_2_1499 ();
 sg13g2_decap_8 FILLER_2_1506 ();
 sg13g2_decap_8 FILLER_2_1513 ();
 sg13g2_decap_8 FILLER_2_1520 ();
 sg13g2_decap_8 FILLER_2_1527 ();
 sg13g2_decap_8 FILLER_2_1534 ();
 sg13g2_decap_8 FILLER_2_1541 ();
 sg13g2_decap_8 FILLER_2_1548 ();
 sg13g2_decap_8 FILLER_2_1555 ();
 sg13g2_decap_8 FILLER_2_1562 ();
 sg13g2_decap_8 FILLER_2_1569 ();
 sg13g2_decap_8 FILLER_2_1576 ();
 sg13g2_decap_8 FILLER_2_1583 ();
 sg13g2_decap_8 FILLER_2_1590 ();
 sg13g2_decap_8 FILLER_2_1597 ();
 sg13g2_decap_8 FILLER_2_1604 ();
 sg13g2_decap_8 FILLER_2_1611 ();
 sg13g2_decap_8 FILLER_2_1618 ();
 sg13g2_decap_8 FILLER_2_1625 ();
 sg13g2_decap_8 FILLER_2_1632 ();
 sg13g2_decap_8 FILLER_2_1639 ();
 sg13g2_decap_8 FILLER_2_1646 ();
 sg13g2_decap_8 FILLER_2_1653 ();
 sg13g2_decap_8 FILLER_2_1660 ();
 sg13g2_decap_8 FILLER_2_1667 ();
 sg13g2_decap_8 FILLER_2_1674 ();
 sg13g2_decap_8 FILLER_2_1681 ();
 sg13g2_decap_8 FILLER_2_1688 ();
 sg13g2_decap_8 FILLER_2_1695 ();
 sg13g2_decap_8 FILLER_2_1702 ();
 sg13g2_decap_8 FILLER_2_1709 ();
 sg13g2_decap_8 FILLER_2_1716 ();
 sg13g2_decap_8 FILLER_2_1723 ();
 sg13g2_decap_8 FILLER_2_1730 ();
 sg13g2_decap_8 FILLER_2_1737 ();
 sg13g2_decap_8 FILLER_2_1744 ();
 sg13g2_decap_8 FILLER_2_1751 ();
 sg13g2_decap_8 FILLER_2_1758 ();
 sg13g2_fill_2 FILLER_2_1765 ();
 sg13g2_fill_1 FILLER_2_1767 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_fill_2 FILLER_3_203 ();
 sg13g2_fill_2 FILLER_3_242 ();
 sg13g2_decap_8 FILLER_3_283 ();
 sg13g2_decap_4 FILLER_3_290 ();
 sg13g2_fill_1 FILLER_3_294 ();
 sg13g2_fill_1 FILLER_3_325 ();
 sg13g2_fill_2 FILLER_3_335 ();
 sg13g2_fill_1 FILLER_3_372 ();
 sg13g2_fill_1 FILLER_3_521 ();
 sg13g2_fill_1 FILLER_3_527 ();
 sg13g2_fill_1 FILLER_3_532 ();
 sg13g2_fill_2 FILLER_3_561 ();
 sg13g2_fill_1 FILLER_3_582 ();
 sg13g2_decap_8 FILLER_3_637 ();
 sg13g2_decap_4 FILLER_3_644 ();
 sg13g2_fill_1 FILLER_3_648 ();
 sg13g2_decap_4 FILLER_3_675 ();
 sg13g2_decap_4 FILLER_3_705 ();
 sg13g2_fill_2 FILLER_3_740 ();
 sg13g2_decap_4 FILLER_3_769 ();
 sg13g2_fill_2 FILLER_3_773 ();
 sg13g2_decap_8 FILLER_3_791 ();
 sg13g2_decap_8 FILLER_3_798 ();
 sg13g2_decap_8 FILLER_3_805 ();
 sg13g2_fill_1 FILLER_3_812 ();
 sg13g2_decap_8 FILLER_3_839 ();
 sg13g2_decap_8 FILLER_3_846 ();
 sg13g2_decap_8 FILLER_3_853 ();
 sg13g2_decap_4 FILLER_3_860 ();
 sg13g2_fill_1 FILLER_3_864 ();
 sg13g2_decap_4 FILLER_3_874 ();
 sg13g2_fill_2 FILLER_3_878 ();
 sg13g2_fill_2 FILLER_3_967 ();
 sg13g2_decap_8 FILLER_3_1055 ();
 sg13g2_decap_8 FILLER_3_1077 ();
 sg13g2_fill_1 FILLER_3_1084 ();
 sg13g2_fill_2 FILLER_3_1089 ();
 sg13g2_fill_1 FILLER_3_1091 ();
 sg13g2_fill_2 FILLER_3_1102 ();
 sg13g2_fill_1 FILLER_3_1104 ();
 sg13g2_decap_4 FILLER_3_1114 ();
 sg13g2_fill_1 FILLER_3_1118 ();
 sg13g2_decap_8 FILLER_3_1132 ();
 sg13g2_decap_8 FILLER_3_1139 ();
 sg13g2_fill_2 FILLER_3_1146 ();
 sg13g2_fill_1 FILLER_3_1148 ();
 sg13g2_decap_4 FILLER_3_1153 ();
 sg13g2_fill_2 FILLER_3_1157 ();
 sg13g2_fill_2 FILLER_3_1176 ();
 sg13g2_decap_8 FILLER_3_1188 ();
 sg13g2_decap_8 FILLER_3_1195 ();
 sg13g2_decap_8 FILLER_3_1202 ();
 sg13g2_decap_8 FILLER_3_1209 ();
 sg13g2_decap_8 FILLER_3_1216 ();
 sg13g2_decap_8 FILLER_3_1223 ();
 sg13g2_decap_8 FILLER_3_1230 ();
 sg13g2_decap_8 FILLER_3_1237 ();
 sg13g2_decap_8 FILLER_3_1244 ();
 sg13g2_decap_8 FILLER_3_1251 ();
 sg13g2_decap_8 FILLER_3_1258 ();
 sg13g2_decap_8 FILLER_3_1265 ();
 sg13g2_decap_8 FILLER_3_1272 ();
 sg13g2_decap_8 FILLER_3_1279 ();
 sg13g2_decap_8 FILLER_3_1286 ();
 sg13g2_decap_8 FILLER_3_1293 ();
 sg13g2_decap_8 FILLER_3_1300 ();
 sg13g2_decap_8 FILLER_3_1307 ();
 sg13g2_decap_8 FILLER_3_1314 ();
 sg13g2_decap_8 FILLER_3_1321 ();
 sg13g2_decap_8 FILLER_3_1328 ();
 sg13g2_decap_8 FILLER_3_1335 ();
 sg13g2_decap_8 FILLER_3_1342 ();
 sg13g2_decap_8 FILLER_3_1349 ();
 sg13g2_decap_8 FILLER_3_1356 ();
 sg13g2_decap_8 FILLER_3_1363 ();
 sg13g2_decap_8 FILLER_3_1370 ();
 sg13g2_decap_8 FILLER_3_1377 ();
 sg13g2_decap_8 FILLER_3_1384 ();
 sg13g2_decap_8 FILLER_3_1391 ();
 sg13g2_decap_8 FILLER_3_1398 ();
 sg13g2_decap_8 FILLER_3_1405 ();
 sg13g2_decap_8 FILLER_3_1412 ();
 sg13g2_decap_8 FILLER_3_1419 ();
 sg13g2_decap_8 FILLER_3_1426 ();
 sg13g2_decap_8 FILLER_3_1433 ();
 sg13g2_decap_8 FILLER_3_1440 ();
 sg13g2_decap_8 FILLER_3_1447 ();
 sg13g2_decap_8 FILLER_3_1454 ();
 sg13g2_decap_8 FILLER_3_1461 ();
 sg13g2_decap_8 FILLER_3_1468 ();
 sg13g2_decap_8 FILLER_3_1475 ();
 sg13g2_decap_8 FILLER_3_1482 ();
 sg13g2_decap_8 FILLER_3_1489 ();
 sg13g2_decap_8 FILLER_3_1496 ();
 sg13g2_decap_8 FILLER_3_1503 ();
 sg13g2_decap_8 FILLER_3_1510 ();
 sg13g2_decap_8 FILLER_3_1517 ();
 sg13g2_decap_8 FILLER_3_1524 ();
 sg13g2_decap_8 FILLER_3_1531 ();
 sg13g2_decap_8 FILLER_3_1538 ();
 sg13g2_decap_8 FILLER_3_1545 ();
 sg13g2_decap_8 FILLER_3_1552 ();
 sg13g2_decap_8 FILLER_3_1559 ();
 sg13g2_decap_8 FILLER_3_1566 ();
 sg13g2_decap_8 FILLER_3_1573 ();
 sg13g2_decap_8 FILLER_3_1580 ();
 sg13g2_decap_8 FILLER_3_1587 ();
 sg13g2_decap_8 FILLER_3_1594 ();
 sg13g2_decap_8 FILLER_3_1601 ();
 sg13g2_decap_8 FILLER_3_1608 ();
 sg13g2_decap_8 FILLER_3_1615 ();
 sg13g2_decap_8 FILLER_3_1622 ();
 sg13g2_decap_8 FILLER_3_1629 ();
 sg13g2_decap_8 FILLER_3_1636 ();
 sg13g2_decap_8 FILLER_3_1643 ();
 sg13g2_decap_8 FILLER_3_1650 ();
 sg13g2_decap_8 FILLER_3_1657 ();
 sg13g2_decap_8 FILLER_3_1664 ();
 sg13g2_decap_8 FILLER_3_1671 ();
 sg13g2_decap_8 FILLER_3_1678 ();
 sg13g2_decap_8 FILLER_3_1685 ();
 sg13g2_decap_8 FILLER_3_1692 ();
 sg13g2_decap_8 FILLER_3_1699 ();
 sg13g2_decap_8 FILLER_3_1706 ();
 sg13g2_decap_8 FILLER_3_1713 ();
 sg13g2_decap_8 FILLER_3_1720 ();
 sg13g2_decap_8 FILLER_3_1727 ();
 sg13g2_decap_8 FILLER_3_1734 ();
 sg13g2_decap_8 FILLER_3_1741 ();
 sg13g2_decap_8 FILLER_3_1748 ();
 sg13g2_decap_8 FILLER_3_1755 ();
 sg13g2_decap_4 FILLER_3_1762 ();
 sg13g2_fill_2 FILLER_3_1766 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_4 FILLER_4_182 ();
 sg13g2_fill_2 FILLER_4_186 ();
 sg13g2_fill_2 FILLER_4_223 ();
 sg13g2_fill_1 FILLER_4_234 ();
 sg13g2_fill_1 FILLER_4_244 ();
 sg13g2_fill_2 FILLER_4_300 ();
 sg13g2_fill_1 FILLER_4_302 ();
 sg13g2_fill_2 FILLER_4_336 ();
 sg13g2_fill_1 FILLER_4_338 ();
 sg13g2_fill_1 FILLER_4_380 ();
 sg13g2_fill_2 FILLER_4_452 ();
 sg13g2_fill_1 FILLER_4_454 ();
 sg13g2_fill_2 FILLER_4_465 ();
 sg13g2_fill_1 FILLER_4_467 ();
 sg13g2_fill_2 FILLER_4_477 ();
 sg13g2_fill_2 FILLER_4_484 ();
 sg13g2_fill_1 FILLER_4_486 ();
 sg13g2_fill_2 FILLER_4_510 ();
 sg13g2_fill_1 FILLER_4_548 ();
 sg13g2_fill_1 FILLER_4_575 ();
 sg13g2_fill_1 FILLER_4_598 ();
 sg13g2_fill_1 FILLER_4_643 ();
 sg13g2_fill_2 FILLER_4_723 ();
 sg13g2_fill_1 FILLER_4_756 ();
 sg13g2_fill_2 FILLER_4_805 ();
 sg13g2_decap_4 FILLER_4_820 ();
 sg13g2_fill_1 FILLER_4_824 ();
 sg13g2_decap_4 FILLER_4_851 ();
 sg13g2_fill_2 FILLER_4_890 ();
 sg13g2_fill_2 FILLER_4_949 ();
 sg13g2_decap_8 FILLER_4_972 ();
 sg13g2_fill_2 FILLER_4_979 ();
 sg13g2_fill_1 FILLER_4_981 ();
 sg13g2_fill_2 FILLER_4_992 ();
 sg13g2_fill_1 FILLER_4_1003 ();
 sg13g2_fill_2 FILLER_4_1022 ();
 sg13g2_fill_1 FILLER_4_1024 ();
 sg13g2_fill_2 FILLER_4_1061 ();
 sg13g2_fill_1 FILLER_4_1063 ();
 sg13g2_fill_2 FILLER_4_1120 ();
 sg13g2_fill_1 FILLER_4_1136 ();
 sg13g2_fill_2 FILLER_4_1178 ();
 sg13g2_fill_1 FILLER_4_1199 ();
 sg13g2_decap_8 FILLER_4_1209 ();
 sg13g2_decap_8 FILLER_4_1216 ();
 sg13g2_decap_8 FILLER_4_1223 ();
 sg13g2_fill_2 FILLER_4_1230 ();
 sg13g2_fill_2 FILLER_4_1236 ();
 sg13g2_fill_2 FILLER_4_1242 ();
 sg13g2_fill_1 FILLER_4_1244 ();
 sg13g2_decap_8 FILLER_4_1249 ();
 sg13g2_decap_8 FILLER_4_1256 ();
 sg13g2_decap_8 FILLER_4_1263 ();
 sg13g2_decap_8 FILLER_4_1270 ();
 sg13g2_decap_8 FILLER_4_1277 ();
 sg13g2_decap_8 FILLER_4_1284 ();
 sg13g2_decap_8 FILLER_4_1291 ();
 sg13g2_decap_8 FILLER_4_1298 ();
 sg13g2_decap_8 FILLER_4_1305 ();
 sg13g2_decap_8 FILLER_4_1312 ();
 sg13g2_decap_8 FILLER_4_1319 ();
 sg13g2_decap_8 FILLER_4_1326 ();
 sg13g2_decap_8 FILLER_4_1333 ();
 sg13g2_decap_8 FILLER_4_1340 ();
 sg13g2_decap_8 FILLER_4_1347 ();
 sg13g2_decap_8 FILLER_4_1354 ();
 sg13g2_decap_8 FILLER_4_1361 ();
 sg13g2_decap_8 FILLER_4_1368 ();
 sg13g2_decap_8 FILLER_4_1375 ();
 sg13g2_decap_8 FILLER_4_1382 ();
 sg13g2_decap_8 FILLER_4_1389 ();
 sg13g2_decap_8 FILLER_4_1396 ();
 sg13g2_decap_8 FILLER_4_1403 ();
 sg13g2_decap_8 FILLER_4_1410 ();
 sg13g2_decap_8 FILLER_4_1417 ();
 sg13g2_decap_8 FILLER_4_1424 ();
 sg13g2_decap_8 FILLER_4_1431 ();
 sg13g2_decap_8 FILLER_4_1438 ();
 sg13g2_decap_8 FILLER_4_1445 ();
 sg13g2_decap_8 FILLER_4_1452 ();
 sg13g2_decap_8 FILLER_4_1459 ();
 sg13g2_decap_8 FILLER_4_1466 ();
 sg13g2_decap_8 FILLER_4_1473 ();
 sg13g2_decap_8 FILLER_4_1480 ();
 sg13g2_decap_8 FILLER_4_1487 ();
 sg13g2_decap_8 FILLER_4_1494 ();
 sg13g2_decap_8 FILLER_4_1501 ();
 sg13g2_decap_8 FILLER_4_1508 ();
 sg13g2_decap_8 FILLER_4_1515 ();
 sg13g2_decap_8 FILLER_4_1522 ();
 sg13g2_decap_8 FILLER_4_1529 ();
 sg13g2_decap_8 FILLER_4_1536 ();
 sg13g2_decap_8 FILLER_4_1543 ();
 sg13g2_decap_8 FILLER_4_1550 ();
 sg13g2_decap_8 FILLER_4_1557 ();
 sg13g2_decap_8 FILLER_4_1564 ();
 sg13g2_decap_8 FILLER_4_1571 ();
 sg13g2_decap_8 FILLER_4_1578 ();
 sg13g2_decap_8 FILLER_4_1585 ();
 sg13g2_decap_8 FILLER_4_1592 ();
 sg13g2_decap_8 FILLER_4_1599 ();
 sg13g2_decap_8 FILLER_4_1606 ();
 sg13g2_decap_8 FILLER_4_1613 ();
 sg13g2_decap_8 FILLER_4_1620 ();
 sg13g2_decap_8 FILLER_4_1627 ();
 sg13g2_decap_8 FILLER_4_1634 ();
 sg13g2_decap_8 FILLER_4_1641 ();
 sg13g2_decap_8 FILLER_4_1648 ();
 sg13g2_decap_8 FILLER_4_1655 ();
 sg13g2_decap_8 FILLER_4_1662 ();
 sg13g2_decap_8 FILLER_4_1669 ();
 sg13g2_decap_8 FILLER_4_1676 ();
 sg13g2_decap_8 FILLER_4_1683 ();
 sg13g2_decap_8 FILLER_4_1690 ();
 sg13g2_decap_8 FILLER_4_1697 ();
 sg13g2_decap_8 FILLER_4_1704 ();
 sg13g2_decap_8 FILLER_4_1711 ();
 sg13g2_decap_8 FILLER_4_1718 ();
 sg13g2_decap_8 FILLER_4_1725 ();
 sg13g2_decap_8 FILLER_4_1732 ();
 sg13g2_decap_8 FILLER_4_1739 ();
 sg13g2_decap_8 FILLER_4_1746 ();
 sg13g2_decap_8 FILLER_4_1753 ();
 sg13g2_decap_8 FILLER_4_1760 ();
 sg13g2_fill_1 FILLER_4_1767 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_4 FILLER_5_175 ();
 sg13g2_fill_1 FILLER_5_179 ();
 sg13g2_fill_2 FILLER_5_219 ();
 sg13g2_fill_1 FILLER_5_221 ();
 sg13g2_fill_1 FILLER_5_230 ();
 sg13g2_fill_2 FILLER_5_327 ();
 sg13g2_fill_1 FILLER_5_338 ();
 sg13g2_fill_2 FILLER_5_447 ();
 sg13g2_fill_1 FILLER_5_458 ();
 sg13g2_fill_1 FILLER_5_560 ();
 sg13g2_decap_4 FILLER_5_641 ();
 sg13g2_fill_2 FILLER_5_661 ();
 sg13g2_decap_8 FILLER_5_672 ();
 sg13g2_fill_2 FILLER_5_679 ();
 sg13g2_fill_1 FILLER_5_681 ();
 sg13g2_fill_1 FILLER_5_698 ();
 sg13g2_fill_1 FILLER_5_720 ();
 sg13g2_fill_2 FILLER_5_756 ();
 sg13g2_fill_2 FILLER_5_771 ();
 sg13g2_fill_2 FILLER_5_791 ();
 sg13g2_decap_8 FILLER_5_802 ();
 sg13g2_fill_2 FILLER_5_809 ();
 sg13g2_decap_8 FILLER_5_846 ();
 sg13g2_fill_1 FILLER_5_853 ();
 sg13g2_decap_4 FILLER_5_860 ();
 sg13g2_decap_8 FILLER_5_874 ();
 sg13g2_fill_2 FILLER_5_899 ();
 sg13g2_decap_4 FILLER_5_910 ();
 sg13g2_fill_1 FILLER_5_923 ();
 sg13g2_fill_1 FILLER_5_934 ();
 sg13g2_fill_2 FILLER_5_941 ();
 sg13g2_fill_2 FILLER_5_990 ();
 sg13g2_fill_2 FILLER_5_996 ();
 sg13g2_fill_2 FILLER_5_1009 ();
 sg13g2_fill_2 FILLER_5_1060 ();
 sg13g2_fill_1 FILLER_5_1062 ();
 sg13g2_fill_1 FILLER_5_1171 ();
 sg13g2_decap_8 FILLER_5_1215 ();
 sg13g2_decap_4 FILLER_5_1222 ();
 sg13g2_fill_1 FILLER_5_1226 ();
 sg13g2_fill_2 FILLER_5_1245 ();
 sg13g2_fill_1 FILLER_5_1247 ();
 sg13g2_fill_1 FILLER_5_1253 ();
 sg13g2_decap_8 FILLER_5_1268 ();
 sg13g2_decap_8 FILLER_5_1275 ();
 sg13g2_decap_8 FILLER_5_1282 ();
 sg13g2_decap_8 FILLER_5_1289 ();
 sg13g2_decap_8 FILLER_5_1296 ();
 sg13g2_decap_8 FILLER_5_1303 ();
 sg13g2_decap_8 FILLER_5_1310 ();
 sg13g2_decap_8 FILLER_5_1317 ();
 sg13g2_decap_8 FILLER_5_1324 ();
 sg13g2_decap_8 FILLER_5_1331 ();
 sg13g2_decap_8 FILLER_5_1338 ();
 sg13g2_decap_8 FILLER_5_1345 ();
 sg13g2_decap_8 FILLER_5_1352 ();
 sg13g2_decap_8 FILLER_5_1359 ();
 sg13g2_decap_8 FILLER_5_1366 ();
 sg13g2_decap_8 FILLER_5_1373 ();
 sg13g2_decap_8 FILLER_5_1380 ();
 sg13g2_decap_8 FILLER_5_1387 ();
 sg13g2_decap_8 FILLER_5_1394 ();
 sg13g2_decap_8 FILLER_5_1401 ();
 sg13g2_decap_8 FILLER_5_1408 ();
 sg13g2_decap_8 FILLER_5_1415 ();
 sg13g2_decap_8 FILLER_5_1422 ();
 sg13g2_decap_8 FILLER_5_1429 ();
 sg13g2_decap_8 FILLER_5_1436 ();
 sg13g2_decap_8 FILLER_5_1443 ();
 sg13g2_decap_8 FILLER_5_1450 ();
 sg13g2_decap_8 FILLER_5_1457 ();
 sg13g2_decap_8 FILLER_5_1464 ();
 sg13g2_decap_8 FILLER_5_1471 ();
 sg13g2_decap_8 FILLER_5_1478 ();
 sg13g2_decap_8 FILLER_5_1485 ();
 sg13g2_decap_8 FILLER_5_1492 ();
 sg13g2_decap_8 FILLER_5_1499 ();
 sg13g2_decap_8 FILLER_5_1506 ();
 sg13g2_decap_8 FILLER_5_1513 ();
 sg13g2_decap_8 FILLER_5_1520 ();
 sg13g2_decap_8 FILLER_5_1527 ();
 sg13g2_decap_8 FILLER_5_1534 ();
 sg13g2_decap_8 FILLER_5_1541 ();
 sg13g2_decap_8 FILLER_5_1548 ();
 sg13g2_decap_8 FILLER_5_1555 ();
 sg13g2_decap_8 FILLER_5_1562 ();
 sg13g2_decap_8 FILLER_5_1569 ();
 sg13g2_decap_8 FILLER_5_1576 ();
 sg13g2_decap_8 FILLER_5_1583 ();
 sg13g2_decap_8 FILLER_5_1590 ();
 sg13g2_decap_8 FILLER_5_1597 ();
 sg13g2_decap_8 FILLER_5_1604 ();
 sg13g2_decap_8 FILLER_5_1611 ();
 sg13g2_decap_8 FILLER_5_1618 ();
 sg13g2_decap_8 FILLER_5_1625 ();
 sg13g2_decap_8 FILLER_5_1632 ();
 sg13g2_decap_8 FILLER_5_1639 ();
 sg13g2_decap_8 FILLER_5_1646 ();
 sg13g2_decap_8 FILLER_5_1653 ();
 sg13g2_decap_8 FILLER_5_1660 ();
 sg13g2_decap_8 FILLER_5_1667 ();
 sg13g2_decap_8 FILLER_5_1674 ();
 sg13g2_decap_8 FILLER_5_1681 ();
 sg13g2_decap_8 FILLER_5_1688 ();
 sg13g2_decap_8 FILLER_5_1695 ();
 sg13g2_decap_8 FILLER_5_1702 ();
 sg13g2_decap_8 FILLER_5_1709 ();
 sg13g2_decap_8 FILLER_5_1716 ();
 sg13g2_decap_8 FILLER_5_1723 ();
 sg13g2_decap_8 FILLER_5_1730 ();
 sg13g2_decap_8 FILLER_5_1737 ();
 sg13g2_decap_8 FILLER_5_1744 ();
 sg13g2_decap_8 FILLER_5_1751 ();
 sg13g2_decap_8 FILLER_5_1758 ();
 sg13g2_fill_2 FILLER_5_1765 ();
 sg13g2_fill_1 FILLER_5_1767 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_fill_1 FILLER_6_182 ();
 sg13g2_fill_1 FILLER_6_218 ();
 sg13g2_fill_2 FILLER_6_255 ();
 sg13g2_fill_2 FILLER_6_272 ();
 sg13g2_fill_1 FILLER_6_274 ();
 sg13g2_fill_1 FILLER_6_280 ();
 sg13g2_fill_2 FILLER_6_295 ();
 sg13g2_fill_1 FILLER_6_297 ();
 sg13g2_fill_1 FILLER_6_328 ();
 sg13g2_fill_2 FILLER_6_397 ();
 sg13g2_fill_2 FILLER_6_409 ();
 sg13g2_fill_1 FILLER_6_490 ();
 sg13g2_fill_2 FILLER_6_505 ();
 sg13g2_fill_1 FILLER_6_516 ();
 sg13g2_fill_1 FILLER_6_638 ();
 sg13g2_decap_4 FILLER_6_724 ();
 sg13g2_fill_1 FILLER_6_789 ();
 sg13g2_decap_4 FILLER_6_816 ();
 sg13g2_fill_2 FILLER_6_820 ();
 sg13g2_fill_2 FILLER_6_861 ();
 sg13g2_fill_2 FILLER_6_878 ();
 sg13g2_decap_4 FILLER_6_892 ();
 sg13g2_decap_4 FILLER_6_913 ();
 sg13g2_fill_2 FILLER_6_917 ();
 sg13g2_fill_1 FILLER_6_942 ();
 sg13g2_fill_2 FILLER_6_1008 ();
 sg13g2_fill_1 FILLER_6_1022 ();
 sg13g2_fill_2 FILLER_6_1065 ();
 sg13g2_fill_1 FILLER_6_1067 ();
 sg13g2_fill_2 FILLER_6_1082 ();
 sg13g2_fill_2 FILLER_6_1181 ();
 sg13g2_fill_1 FILLER_6_1183 ();
 sg13g2_decap_8 FILLER_6_1271 ();
 sg13g2_decap_8 FILLER_6_1278 ();
 sg13g2_decap_8 FILLER_6_1285 ();
 sg13g2_decap_8 FILLER_6_1292 ();
 sg13g2_decap_8 FILLER_6_1299 ();
 sg13g2_decap_8 FILLER_6_1306 ();
 sg13g2_decap_8 FILLER_6_1313 ();
 sg13g2_decap_8 FILLER_6_1320 ();
 sg13g2_decap_8 FILLER_6_1327 ();
 sg13g2_decap_8 FILLER_6_1334 ();
 sg13g2_decap_8 FILLER_6_1341 ();
 sg13g2_decap_8 FILLER_6_1348 ();
 sg13g2_decap_8 FILLER_6_1355 ();
 sg13g2_decap_8 FILLER_6_1362 ();
 sg13g2_decap_8 FILLER_6_1369 ();
 sg13g2_decap_8 FILLER_6_1376 ();
 sg13g2_decap_8 FILLER_6_1383 ();
 sg13g2_decap_8 FILLER_6_1390 ();
 sg13g2_decap_8 FILLER_6_1397 ();
 sg13g2_decap_8 FILLER_6_1404 ();
 sg13g2_decap_8 FILLER_6_1411 ();
 sg13g2_decap_8 FILLER_6_1418 ();
 sg13g2_decap_8 FILLER_6_1425 ();
 sg13g2_decap_8 FILLER_6_1432 ();
 sg13g2_decap_8 FILLER_6_1439 ();
 sg13g2_decap_8 FILLER_6_1446 ();
 sg13g2_decap_8 FILLER_6_1453 ();
 sg13g2_decap_8 FILLER_6_1460 ();
 sg13g2_decap_8 FILLER_6_1467 ();
 sg13g2_decap_8 FILLER_6_1474 ();
 sg13g2_decap_8 FILLER_6_1481 ();
 sg13g2_decap_8 FILLER_6_1488 ();
 sg13g2_decap_8 FILLER_6_1495 ();
 sg13g2_decap_8 FILLER_6_1502 ();
 sg13g2_decap_8 FILLER_6_1509 ();
 sg13g2_decap_8 FILLER_6_1516 ();
 sg13g2_decap_8 FILLER_6_1523 ();
 sg13g2_decap_8 FILLER_6_1530 ();
 sg13g2_decap_8 FILLER_6_1537 ();
 sg13g2_decap_8 FILLER_6_1544 ();
 sg13g2_decap_8 FILLER_6_1551 ();
 sg13g2_decap_8 FILLER_6_1558 ();
 sg13g2_decap_8 FILLER_6_1565 ();
 sg13g2_decap_8 FILLER_6_1572 ();
 sg13g2_decap_8 FILLER_6_1579 ();
 sg13g2_decap_8 FILLER_6_1586 ();
 sg13g2_decap_8 FILLER_6_1593 ();
 sg13g2_decap_8 FILLER_6_1600 ();
 sg13g2_decap_8 FILLER_6_1607 ();
 sg13g2_decap_8 FILLER_6_1614 ();
 sg13g2_decap_8 FILLER_6_1621 ();
 sg13g2_decap_8 FILLER_6_1628 ();
 sg13g2_decap_8 FILLER_6_1635 ();
 sg13g2_decap_8 FILLER_6_1642 ();
 sg13g2_decap_8 FILLER_6_1649 ();
 sg13g2_decap_8 FILLER_6_1656 ();
 sg13g2_decap_8 FILLER_6_1663 ();
 sg13g2_decap_8 FILLER_6_1670 ();
 sg13g2_decap_8 FILLER_6_1677 ();
 sg13g2_decap_8 FILLER_6_1684 ();
 sg13g2_decap_8 FILLER_6_1691 ();
 sg13g2_decap_8 FILLER_6_1698 ();
 sg13g2_decap_8 FILLER_6_1705 ();
 sg13g2_decap_8 FILLER_6_1712 ();
 sg13g2_decap_8 FILLER_6_1719 ();
 sg13g2_decap_8 FILLER_6_1726 ();
 sg13g2_decap_8 FILLER_6_1733 ();
 sg13g2_decap_8 FILLER_6_1740 ();
 sg13g2_decap_8 FILLER_6_1747 ();
 sg13g2_decap_8 FILLER_6_1754 ();
 sg13g2_decap_8 FILLER_6_1761 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_fill_2 FILLER_7_175 ();
 sg13g2_fill_2 FILLER_7_211 ();
 sg13g2_fill_1 FILLER_7_225 ();
 sg13g2_fill_2 FILLER_7_300 ();
 sg13g2_fill_1 FILLER_7_302 ();
 sg13g2_fill_2 FILLER_7_375 ();
 sg13g2_fill_2 FILLER_7_412 ();
 sg13g2_fill_1 FILLER_7_414 ();
 sg13g2_fill_2 FILLER_7_431 ();
 sg13g2_fill_2 FILLER_7_478 ();
 sg13g2_fill_1 FILLER_7_577 ();
 sg13g2_fill_1 FILLER_7_614 ();
 sg13g2_fill_1 FILLER_7_695 ();
 sg13g2_fill_2 FILLER_7_712 ();
 sg13g2_fill_1 FILLER_7_732 ();
 sg13g2_fill_2 FILLER_7_769 ();
 sg13g2_fill_2 FILLER_7_802 ();
 sg13g2_decap_4 FILLER_7_809 ();
 sg13g2_fill_1 FILLER_7_813 ();
 sg13g2_fill_2 FILLER_7_828 ();
 sg13g2_fill_2 FILLER_7_847 ();
 sg13g2_decap_8 FILLER_7_857 ();
 sg13g2_fill_2 FILLER_7_876 ();
 sg13g2_decap_8 FILLER_7_888 ();
 sg13g2_decap_4 FILLER_7_895 ();
 sg13g2_fill_2 FILLER_7_940 ();
 sg13g2_fill_2 FILLER_7_946 ();
 sg13g2_decap_8 FILLER_7_965 ();
 sg13g2_fill_2 FILLER_7_972 ();
 sg13g2_decap_8 FILLER_7_984 ();
 sg13g2_fill_1 FILLER_7_991 ();
 sg13g2_fill_2 FILLER_7_1024 ();
 sg13g2_fill_1 FILLER_7_1026 ();
 sg13g2_fill_2 FILLER_7_1064 ();
 sg13g2_fill_1 FILLER_7_1066 ();
 sg13g2_fill_2 FILLER_7_1108 ();
 sg13g2_fill_2 FILLER_7_1168 ();
 sg13g2_fill_2 FILLER_7_1193 ();
 sg13g2_fill_2 FILLER_7_1242 ();
 sg13g2_decap_8 FILLER_7_1281 ();
 sg13g2_decap_8 FILLER_7_1288 ();
 sg13g2_decap_8 FILLER_7_1295 ();
 sg13g2_decap_8 FILLER_7_1302 ();
 sg13g2_decap_8 FILLER_7_1309 ();
 sg13g2_decap_8 FILLER_7_1316 ();
 sg13g2_decap_8 FILLER_7_1323 ();
 sg13g2_decap_8 FILLER_7_1330 ();
 sg13g2_decap_8 FILLER_7_1337 ();
 sg13g2_decap_8 FILLER_7_1344 ();
 sg13g2_decap_8 FILLER_7_1351 ();
 sg13g2_decap_8 FILLER_7_1358 ();
 sg13g2_decap_8 FILLER_7_1365 ();
 sg13g2_decap_8 FILLER_7_1372 ();
 sg13g2_decap_8 FILLER_7_1379 ();
 sg13g2_decap_8 FILLER_7_1386 ();
 sg13g2_decap_8 FILLER_7_1393 ();
 sg13g2_decap_8 FILLER_7_1400 ();
 sg13g2_decap_8 FILLER_7_1407 ();
 sg13g2_decap_8 FILLER_7_1414 ();
 sg13g2_decap_8 FILLER_7_1421 ();
 sg13g2_decap_8 FILLER_7_1428 ();
 sg13g2_decap_8 FILLER_7_1435 ();
 sg13g2_decap_8 FILLER_7_1442 ();
 sg13g2_decap_8 FILLER_7_1449 ();
 sg13g2_decap_8 FILLER_7_1456 ();
 sg13g2_decap_8 FILLER_7_1463 ();
 sg13g2_decap_8 FILLER_7_1470 ();
 sg13g2_decap_8 FILLER_7_1477 ();
 sg13g2_decap_8 FILLER_7_1484 ();
 sg13g2_decap_8 FILLER_7_1491 ();
 sg13g2_decap_8 FILLER_7_1498 ();
 sg13g2_decap_8 FILLER_7_1505 ();
 sg13g2_decap_8 FILLER_7_1512 ();
 sg13g2_decap_8 FILLER_7_1519 ();
 sg13g2_decap_8 FILLER_7_1526 ();
 sg13g2_decap_8 FILLER_7_1533 ();
 sg13g2_decap_8 FILLER_7_1540 ();
 sg13g2_decap_8 FILLER_7_1547 ();
 sg13g2_decap_8 FILLER_7_1554 ();
 sg13g2_decap_8 FILLER_7_1561 ();
 sg13g2_decap_8 FILLER_7_1568 ();
 sg13g2_decap_8 FILLER_7_1575 ();
 sg13g2_decap_8 FILLER_7_1582 ();
 sg13g2_decap_8 FILLER_7_1589 ();
 sg13g2_decap_8 FILLER_7_1596 ();
 sg13g2_decap_8 FILLER_7_1603 ();
 sg13g2_decap_8 FILLER_7_1610 ();
 sg13g2_decap_8 FILLER_7_1617 ();
 sg13g2_decap_8 FILLER_7_1624 ();
 sg13g2_decap_8 FILLER_7_1631 ();
 sg13g2_decap_8 FILLER_7_1638 ();
 sg13g2_decap_8 FILLER_7_1645 ();
 sg13g2_decap_8 FILLER_7_1652 ();
 sg13g2_decap_8 FILLER_7_1659 ();
 sg13g2_decap_8 FILLER_7_1666 ();
 sg13g2_decap_8 FILLER_7_1673 ();
 sg13g2_decap_8 FILLER_7_1680 ();
 sg13g2_decap_8 FILLER_7_1687 ();
 sg13g2_decap_8 FILLER_7_1694 ();
 sg13g2_decap_8 FILLER_7_1701 ();
 sg13g2_decap_8 FILLER_7_1708 ();
 sg13g2_decap_8 FILLER_7_1715 ();
 sg13g2_decap_8 FILLER_7_1722 ();
 sg13g2_decap_8 FILLER_7_1729 ();
 sg13g2_decap_8 FILLER_7_1736 ();
 sg13g2_decap_8 FILLER_7_1743 ();
 sg13g2_decap_8 FILLER_7_1750 ();
 sg13g2_decap_8 FILLER_7_1757 ();
 sg13g2_decap_4 FILLER_7_1764 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_fill_2 FILLER_8_168 ();
 sg13g2_fill_1 FILLER_8_196 ();
 sg13g2_fill_2 FILLER_8_214 ();
 sg13g2_fill_1 FILLER_8_216 ();
 sg13g2_fill_2 FILLER_8_243 ();
 sg13g2_fill_1 FILLER_8_287 ();
 sg13g2_fill_2 FILLER_8_324 ();
 sg13g2_fill_1 FILLER_8_348 ();
 sg13g2_fill_2 FILLER_8_380 ();
 sg13g2_fill_2 FILLER_8_395 ();
 sg13g2_fill_2 FILLER_8_423 ();
 sg13g2_fill_1 FILLER_8_425 ();
 sg13g2_fill_1 FILLER_8_434 ();
 sg13g2_fill_1 FILLER_8_445 ();
 sg13g2_fill_1 FILLER_8_472 ();
 sg13g2_fill_2 FILLER_8_488 ();
 sg13g2_fill_1 FILLER_8_547 ();
 sg13g2_decap_4 FILLER_8_569 ();
 sg13g2_fill_2 FILLER_8_573 ();
 sg13g2_fill_2 FILLER_8_586 ();
 sg13g2_fill_2 FILLER_8_592 ();
 sg13g2_fill_2 FILLER_8_630 ();
 sg13g2_fill_1 FILLER_8_650 ();
 sg13g2_fill_1 FILLER_8_660 ();
 sg13g2_fill_2 FILLER_8_702 ();
 sg13g2_fill_2 FILLER_8_730 ();
 sg13g2_fill_1 FILLER_8_766 ();
 sg13g2_fill_2 FILLER_8_790 ();
 sg13g2_fill_1 FILLER_8_792 ();
 sg13g2_fill_2 FILLER_8_804 ();
 sg13g2_fill_2 FILLER_8_863 ();
 sg13g2_fill_2 FILLER_8_878 ();
 sg13g2_fill_1 FILLER_8_880 ();
 sg13g2_fill_1 FILLER_8_886 ();
 sg13g2_fill_2 FILLER_8_913 ();
 sg13g2_fill_1 FILLER_8_915 ();
 sg13g2_fill_2 FILLER_8_927 ();
 sg13g2_fill_1 FILLER_8_935 ();
 sg13g2_decap_8 FILLER_8_979 ();
 sg13g2_decap_8 FILLER_8_986 ();
 sg13g2_fill_1 FILLER_8_993 ();
 sg13g2_fill_2 FILLER_8_1000 ();
 sg13g2_fill_1 FILLER_8_1028 ();
 sg13g2_fill_1 FILLER_8_1057 ();
 sg13g2_fill_2 FILLER_8_1086 ();
 sg13g2_fill_2 FILLER_8_1135 ();
 sg13g2_fill_2 FILLER_8_1156 ();
 sg13g2_fill_1 FILLER_8_1158 ();
 sg13g2_fill_2 FILLER_8_1248 ();
 sg13g2_decap_8 FILLER_8_1285 ();
 sg13g2_decap_8 FILLER_8_1292 ();
 sg13g2_decap_8 FILLER_8_1299 ();
 sg13g2_decap_8 FILLER_8_1306 ();
 sg13g2_decap_8 FILLER_8_1313 ();
 sg13g2_decap_8 FILLER_8_1320 ();
 sg13g2_decap_8 FILLER_8_1327 ();
 sg13g2_decap_8 FILLER_8_1334 ();
 sg13g2_decap_8 FILLER_8_1341 ();
 sg13g2_decap_8 FILLER_8_1348 ();
 sg13g2_decap_8 FILLER_8_1355 ();
 sg13g2_decap_8 FILLER_8_1362 ();
 sg13g2_decap_8 FILLER_8_1369 ();
 sg13g2_decap_8 FILLER_8_1376 ();
 sg13g2_decap_8 FILLER_8_1383 ();
 sg13g2_decap_8 FILLER_8_1390 ();
 sg13g2_decap_8 FILLER_8_1397 ();
 sg13g2_decap_8 FILLER_8_1404 ();
 sg13g2_decap_8 FILLER_8_1411 ();
 sg13g2_decap_8 FILLER_8_1418 ();
 sg13g2_decap_8 FILLER_8_1425 ();
 sg13g2_decap_8 FILLER_8_1432 ();
 sg13g2_decap_8 FILLER_8_1439 ();
 sg13g2_decap_8 FILLER_8_1446 ();
 sg13g2_decap_8 FILLER_8_1453 ();
 sg13g2_decap_8 FILLER_8_1460 ();
 sg13g2_decap_8 FILLER_8_1467 ();
 sg13g2_decap_8 FILLER_8_1474 ();
 sg13g2_decap_8 FILLER_8_1481 ();
 sg13g2_decap_8 FILLER_8_1488 ();
 sg13g2_decap_8 FILLER_8_1495 ();
 sg13g2_decap_8 FILLER_8_1502 ();
 sg13g2_decap_8 FILLER_8_1509 ();
 sg13g2_decap_8 FILLER_8_1516 ();
 sg13g2_decap_8 FILLER_8_1523 ();
 sg13g2_decap_8 FILLER_8_1530 ();
 sg13g2_decap_8 FILLER_8_1537 ();
 sg13g2_decap_8 FILLER_8_1544 ();
 sg13g2_decap_8 FILLER_8_1551 ();
 sg13g2_decap_8 FILLER_8_1558 ();
 sg13g2_decap_8 FILLER_8_1565 ();
 sg13g2_decap_8 FILLER_8_1572 ();
 sg13g2_decap_8 FILLER_8_1579 ();
 sg13g2_decap_8 FILLER_8_1586 ();
 sg13g2_decap_8 FILLER_8_1593 ();
 sg13g2_decap_8 FILLER_8_1600 ();
 sg13g2_decap_8 FILLER_8_1607 ();
 sg13g2_decap_8 FILLER_8_1614 ();
 sg13g2_decap_8 FILLER_8_1621 ();
 sg13g2_decap_8 FILLER_8_1628 ();
 sg13g2_decap_8 FILLER_8_1635 ();
 sg13g2_decap_8 FILLER_8_1642 ();
 sg13g2_decap_8 FILLER_8_1649 ();
 sg13g2_decap_8 FILLER_8_1656 ();
 sg13g2_decap_8 FILLER_8_1663 ();
 sg13g2_decap_8 FILLER_8_1670 ();
 sg13g2_decap_8 FILLER_8_1677 ();
 sg13g2_decap_8 FILLER_8_1684 ();
 sg13g2_decap_8 FILLER_8_1691 ();
 sg13g2_decap_8 FILLER_8_1698 ();
 sg13g2_decap_8 FILLER_8_1705 ();
 sg13g2_decap_8 FILLER_8_1712 ();
 sg13g2_decap_8 FILLER_8_1719 ();
 sg13g2_decap_8 FILLER_8_1726 ();
 sg13g2_decap_8 FILLER_8_1733 ();
 sg13g2_decap_8 FILLER_8_1740 ();
 sg13g2_decap_8 FILLER_8_1747 ();
 sg13g2_decap_8 FILLER_8_1754 ();
 sg13g2_decap_8 FILLER_8_1761 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_4 FILLER_9_168 ();
 sg13g2_fill_2 FILLER_9_172 ();
 sg13g2_decap_8 FILLER_9_178 ();
 sg13g2_fill_2 FILLER_9_185 ();
 sg13g2_fill_1 FILLER_9_229 ();
 sg13g2_decap_4 FILLER_9_275 ();
 sg13g2_fill_1 FILLER_9_310 ();
 sg13g2_fill_2 FILLER_9_332 ();
 sg13g2_fill_1 FILLER_9_368 ();
 sg13g2_fill_2 FILLER_9_383 ();
 sg13g2_fill_2 FILLER_9_399 ();
 sg13g2_fill_1 FILLER_9_401 ();
 sg13g2_fill_1 FILLER_9_411 ();
 sg13g2_fill_1 FILLER_9_468 ();
 sg13g2_fill_1 FILLER_9_478 ();
 sg13g2_fill_1 FILLER_9_535 ();
 sg13g2_fill_1 FILLER_9_542 ();
 sg13g2_fill_2 FILLER_9_564 ();
 sg13g2_fill_2 FILLER_9_583 ();
 sg13g2_fill_1 FILLER_9_590 ();
 sg13g2_fill_1 FILLER_9_656 ();
 sg13g2_fill_2 FILLER_9_684 ();
 sg13g2_fill_2 FILLER_9_731 ();
 sg13g2_fill_1 FILLER_9_759 ();
 sg13g2_fill_1 FILLER_9_795 ();
 sg13g2_fill_2 FILLER_9_816 ();
 sg13g2_fill_1 FILLER_9_818 ();
 sg13g2_fill_2 FILLER_9_830 ();
 sg13g2_fill_1 FILLER_9_832 ();
 sg13g2_fill_2 FILLER_9_837 ();
 sg13g2_fill_1 FILLER_9_839 ();
 sg13g2_fill_2 FILLER_9_846 ();
 sg13g2_decap_8 FILLER_9_856 ();
 sg13g2_fill_2 FILLER_9_863 ();
 sg13g2_decap_8 FILLER_9_906 ();
 sg13g2_decap_4 FILLER_9_913 ();
 sg13g2_fill_2 FILLER_9_917 ();
 sg13g2_fill_2 FILLER_9_929 ();
 sg13g2_fill_2 FILLER_9_937 ();
 sg13g2_fill_1 FILLER_9_939 ();
 sg13g2_fill_1 FILLER_9_959 ();
 sg13g2_fill_2 FILLER_9_1017 ();
 sg13g2_fill_2 FILLER_9_1217 ();
 sg13g2_fill_2 FILLER_9_1238 ();
 sg13g2_fill_1 FILLER_9_1254 ();
 sg13g2_fill_1 FILLER_9_1269 ();
 sg13g2_decap_8 FILLER_9_1291 ();
 sg13g2_decap_8 FILLER_9_1298 ();
 sg13g2_decap_8 FILLER_9_1305 ();
 sg13g2_decap_8 FILLER_9_1312 ();
 sg13g2_decap_8 FILLER_9_1319 ();
 sg13g2_decap_8 FILLER_9_1326 ();
 sg13g2_decap_8 FILLER_9_1333 ();
 sg13g2_decap_8 FILLER_9_1340 ();
 sg13g2_decap_8 FILLER_9_1347 ();
 sg13g2_decap_8 FILLER_9_1354 ();
 sg13g2_decap_8 FILLER_9_1361 ();
 sg13g2_decap_8 FILLER_9_1368 ();
 sg13g2_decap_8 FILLER_9_1375 ();
 sg13g2_decap_8 FILLER_9_1382 ();
 sg13g2_decap_8 FILLER_9_1389 ();
 sg13g2_decap_8 FILLER_9_1396 ();
 sg13g2_decap_8 FILLER_9_1403 ();
 sg13g2_decap_8 FILLER_9_1410 ();
 sg13g2_decap_8 FILLER_9_1417 ();
 sg13g2_decap_8 FILLER_9_1424 ();
 sg13g2_decap_8 FILLER_9_1431 ();
 sg13g2_decap_8 FILLER_9_1438 ();
 sg13g2_decap_8 FILLER_9_1445 ();
 sg13g2_decap_8 FILLER_9_1452 ();
 sg13g2_decap_8 FILLER_9_1459 ();
 sg13g2_decap_8 FILLER_9_1466 ();
 sg13g2_decap_8 FILLER_9_1473 ();
 sg13g2_decap_8 FILLER_9_1480 ();
 sg13g2_decap_8 FILLER_9_1487 ();
 sg13g2_decap_8 FILLER_9_1494 ();
 sg13g2_decap_8 FILLER_9_1501 ();
 sg13g2_decap_8 FILLER_9_1508 ();
 sg13g2_decap_8 FILLER_9_1515 ();
 sg13g2_decap_8 FILLER_9_1522 ();
 sg13g2_decap_8 FILLER_9_1529 ();
 sg13g2_decap_8 FILLER_9_1536 ();
 sg13g2_decap_8 FILLER_9_1543 ();
 sg13g2_decap_8 FILLER_9_1550 ();
 sg13g2_decap_8 FILLER_9_1557 ();
 sg13g2_decap_8 FILLER_9_1564 ();
 sg13g2_decap_8 FILLER_9_1571 ();
 sg13g2_decap_8 FILLER_9_1578 ();
 sg13g2_decap_8 FILLER_9_1585 ();
 sg13g2_decap_8 FILLER_9_1592 ();
 sg13g2_decap_8 FILLER_9_1599 ();
 sg13g2_decap_8 FILLER_9_1606 ();
 sg13g2_decap_8 FILLER_9_1613 ();
 sg13g2_decap_8 FILLER_9_1620 ();
 sg13g2_decap_8 FILLER_9_1627 ();
 sg13g2_decap_8 FILLER_9_1634 ();
 sg13g2_decap_8 FILLER_9_1641 ();
 sg13g2_decap_8 FILLER_9_1648 ();
 sg13g2_decap_8 FILLER_9_1655 ();
 sg13g2_decap_8 FILLER_9_1662 ();
 sg13g2_decap_8 FILLER_9_1669 ();
 sg13g2_decap_8 FILLER_9_1676 ();
 sg13g2_decap_8 FILLER_9_1683 ();
 sg13g2_decap_8 FILLER_9_1690 ();
 sg13g2_decap_8 FILLER_9_1697 ();
 sg13g2_decap_8 FILLER_9_1704 ();
 sg13g2_decap_8 FILLER_9_1711 ();
 sg13g2_decap_8 FILLER_9_1718 ();
 sg13g2_decap_8 FILLER_9_1725 ();
 sg13g2_decap_8 FILLER_9_1732 ();
 sg13g2_decap_8 FILLER_9_1739 ();
 sg13g2_decap_8 FILLER_9_1746 ();
 sg13g2_decap_8 FILLER_9_1753 ();
 sg13g2_decap_8 FILLER_9_1760 ();
 sg13g2_fill_1 FILLER_9_1767 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_4 FILLER_10_154 ();
 sg13g2_fill_1 FILLER_10_158 ();
 sg13g2_decap_8 FILLER_10_185 ();
 sg13g2_decap_8 FILLER_10_192 ();
 sg13g2_decap_8 FILLER_10_199 ();
 sg13g2_decap_4 FILLER_10_206 ();
 sg13g2_fill_1 FILLER_10_210 ();
 sg13g2_fill_2 FILLER_10_220 ();
 sg13g2_fill_2 FILLER_10_257 ();
 sg13g2_fill_1 FILLER_10_259 ();
 sg13g2_fill_1 FILLER_10_275 ();
 sg13g2_fill_1 FILLER_10_317 ();
 sg13g2_fill_2 FILLER_10_362 ();
 sg13g2_fill_2 FILLER_10_414 ();
 sg13g2_fill_1 FILLER_10_416 ();
 sg13g2_fill_2 FILLER_10_431 ();
 sg13g2_fill_1 FILLER_10_433 ();
 sg13g2_fill_1 FILLER_10_439 ();
 sg13g2_fill_2 FILLER_10_485 ();
 sg13g2_fill_2 FILLER_10_496 ();
 sg13g2_fill_1 FILLER_10_507 ();
 sg13g2_fill_1 FILLER_10_628 ();
 sg13g2_fill_2 FILLER_10_689 ();
 sg13g2_decap_8 FILLER_10_733 ();
 sg13g2_fill_1 FILLER_10_770 ();
 sg13g2_decap_4 FILLER_10_817 ();
 sg13g2_fill_1 FILLER_10_821 ();
 sg13g2_fill_2 FILLER_10_827 ();
 sg13g2_fill_2 FILLER_10_834 ();
 sg13g2_fill_1 FILLER_10_853 ();
 sg13g2_fill_2 FILLER_10_880 ();
 sg13g2_fill_2 FILLER_10_903 ();
 sg13g2_decap_4 FILLER_10_929 ();
 sg13g2_fill_2 FILLER_10_968 ();
 sg13g2_fill_1 FILLER_10_970 ();
 sg13g2_fill_2 FILLER_10_994 ();
 sg13g2_fill_1 FILLER_10_1010 ();
 sg13g2_fill_2 FILLER_10_1075 ();
 sg13g2_fill_1 FILLER_10_1085 ();
 sg13g2_fill_2 FILLER_10_1106 ();
 sg13g2_fill_1 FILLER_10_1108 ();
 sg13g2_fill_2 FILLER_10_1141 ();
 sg13g2_fill_1 FILLER_10_1143 ();
 sg13g2_fill_1 FILLER_10_1186 ();
 sg13g2_fill_1 FILLER_10_1255 ();
 sg13g2_decap_8 FILLER_10_1286 ();
 sg13g2_decap_8 FILLER_10_1293 ();
 sg13g2_decap_8 FILLER_10_1300 ();
 sg13g2_decap_8 FILLER_10_1307 ();
 sg13g2_decap_8 FILLER_10_1314 ();
 sg13g2_decap_8 FILLER_10_1321 ();
 sg13g2_decap_8 FILLER_10_1328 ();
 sg13g2_decap_8 FILLER_10_1335 ();
 sg13g2_decap_8 FILLER_10_1342 ();
 sg13g2_decap_8 FILLER_10_1349 ();
 sg13g2_decap_8 FILLER_10_1356 ();
 sg13g2_decap_8 FILLER_10_1363 ();
 sg13g2_decap_8 FILLER_10_1370 ();
 sg13g2_decap_8 FILLER_10_1377 ();
 sg13g2_decap_8 FILLER_10_1384 ();
 sg13g2_decap_8 FILLER_10_1391 ();
 sg13g2_decap_8 FILLER_10_1398 ();
 sg13g2_decap_8 FILLER_10_1405 ();
 sg13g2_decap_8 FILLER_10_1412 ();
 sg13g2_decap_8 FILLER_10_1419 ();
 sg13g2_decap_8 FILLER_10_1426 ();
 sg13g2_decap_8 FILLER_10_1433 ();
 sg13g2_decap_8 FILLER_10_1440 ();
 sg13g2_decap_8 FILLER_10_1447 ();
 sg13g2_decap_8 FILLER_10_1454 ();
 sg13g2_decap_8 FILLER_10_1461 ();
 sg13g2_decap_8 FILLER_10_1468 ();
 sg13g2_decap_8 FILLER_10_1475 ();
 sg13g2_decap_8 FILLER_10_1482 ();
 sg13g2_decap_8 FILLER_10_1489 ();
 sg13g2_decap_8 FILLER_10_1496 ();
 sg13g2_decap_8 FILLER_10_1503 ();
 sg13g2_decap_8 FILLER_10_1510 ();
 sg13g2_decap_8 FILLER_10_1517 ();
 sg13g2_decap_8 FILLER_10_1524 ();
 sg13g2_decap_8 FILLER_10_1531 ();
 sg13g2_decap_8 FILLER_10_1538 ();
 sg13g2_decap_8 FILLER_10_1545 ();
 sg13g2_decap_8 FILLER_10_1552 ();
 sg13g2_decap_8 FILLER_10_1559 ();
 sg13g2_decap_8 FILLER_10_1566 ();
 sg13g2_decap_8 FILLER_10_1573 ();
 sg13g2_decap_8 FILLER_10_1580 ();
 sg13g2_decap_8 FILLER_10_1587 ();
 sg13g2_decap_8 FILLER_10_1594 ();
 sg13g2_decap_8 FILLER_10_1601 ();
 sg13g2_decap_8 FILLER_10_1608 ();
 sg13g2_decap_8 FILLER_10_1615 ();
 sg13g2_decap_8 FILLER_10_1622 ();
 sg13g2_decap_8 FILLER_10_1629 ();
 sg13g2_decap_8 FILLER_10_1636 ();
 sg13g2_decap_8 FILLER_10_1643 ();
 sg13g2_decap_8 FILLER_10_1650 ();
 sg13g2_decap_8 FILLER_10_1657 ();
 sg13g2_decap_8 FILLER_10_1664 ();
 sg13g2_decap_8 FILLER_10_1671 ();
 sg13g2_decap_8 FILLER_10_1678 ();
 sg13g2_decap_8 FILLER_10_1685 ();
 sg13g2_decap_8 FILLER_10_1692 ();
 sg13g2_decap_8 FILLER_10_1699 ();
 sg13g2_decap_8 FILLER_10_1706 ();
 sg13g2_decap_8 FILLER_10_1713 ();
 sg13g2_decap_8 FILLER_10_1720 ();
 sg13g2_decap_8 FILLER_10_1727 ();
 sg13g2_decap_8 FILLER_10_1734 ();
 sg13g2_decap_8 FILLER_10_1741 ();
 sg13g2_decap_8 FILLER_10_1748 ();
 sg13g2_decap_8 FILLER_10_1755 ();
 sg13g2_decap_4 FILLER_10_1762 ();
 sg13g2_fill_2 FILLER_10_1766 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_fill_2 FILLER_11_77 ();
 sg13g2_fill_1 FILLER_11_79 ();
 sg13g2_fill_1 FILLER_11_88 ();
 sg13g2_decap_8 FILLER_11_94 ();
 sg13g2_decap_8 FILLER_11_101 ();
 sg13g2_decap_8 FILLER_11_108 ();
 sg13g2_decap_8 FILLER_11_115 ();
 sg13g2_decap_8 FILLER_11_122 ();
 sg13g2_decap_4 FILLER_11_129 ();
 sg13g2_fill_2 FILLER_11_133 ();
 sg13g2_fill_1 FILLER_11_143 ();
 sg13g2_fill_2 FILLER_11_152 ();
 sg13g2_fill_1 FILLER_11_163 ();
 sg13g2_fill_2 FILLER_11_174 ();
 sg13g2_fill_1 FILLER_11_228 ();
 sg13g2_fill_2 FILLER_11_239 ();
 sg13g2_fill_2 FILLER_11_267 ();
 sg13g2_fill_1 FILLER_11_269 ();
 sg13g2_fill_2 FILLER_11_309 ();
 sg13g2_fill_1 FILLER_11_402 ();
 sg13g2_fill_1 FILLER_11_429 ();
 sg13g2_fill_1 FILLER_11_469 ();
 sg13g2_fill_1 FILLER_11_506 ();
 sg13g2_fill_1 FILLER_11_565 ();
 sg13g2_fill_1 FILLER_11_571 ();
 sg13g2_decap_8 FILLER_11_606 ();
 sg13g2_fill_2 FILLER_11_613 ();
 sg13g2_fill_1 FILLER_11_615 ();
 sg13g2_fill_2 FILLER_11_621 ();
 sg13g2_fill_1 FILLER_11_660 ();
 sg13g2_fill_1 FILLER_11_678 ();
 sg13g2_fill_2 FILLER_11_710 ();
 sg13g2_decap_4 FILLER_11_747 ();
 sg13g2_fill_1 FILLER_11_751 ();
 sg13g2_fill_1 FILLER_11_770 ();
 sg13g2_fill_2 FILLER_11_785 ();
 sg13g2_fill_2 FILLER_11_808 ();
 sg13g2_fill_1 FILLER_11_823 ();
 sg13g2_decap_4 FILLER_11_854 ();
 sg13g2_fill_2 FILLER_11_858 ();
 sg13g2_fill_2 FILLER_11_949 ();
 sg13g2_fill_1 FILLER_11_951 ();
 sg13g2_fill_1 FILLER_11_956 ();
 sg13g2_fill_1 FILLER_11_987 ();
 sg13g2_fill_1 FILLER_11_1000 ();
 sg13g2_fill_1 FILLER_11_1017 ();
 sg13g2_fill_2 FILLER_11_1023 ();
 sg13g2_fill_1 FILLER_11_1025 ();
 sg13g2_fill_2 FILLER_11_1064 ();
 sg13g2_decap_4 FILLER_11_1071 ();
 sg13g2_fill_1 FILLER_11_1075 ();
 sg13g2_fill_1 FILLER_11_1143 ();
 sg13g2_fill_2 FILLER_11_1184 ();
 sg13g2_fill_2 FILLER_11_1239 ();
 sg13g2_fill_1 FILLER_11_1241 ();
 sg13g2_fill_2 FILLER_11_1252 ();
 sg13g2_fill_1 FILLER_11_1254 ();
 sg13g2_fill_1 FILLER_11_1264 ();
 sg13g2_decap_8 FILLER_11_1300 ();
 sg13g2_decap_8 FILLER_11_1307 ();
 sg13g2_decap_8 FILLER_11_1314 ();
 sg13g2_decap_8 FILLER_11_1321 ();
 sg13g2_decap_8 FILLER_11_1328 ();
 sg13g2_decap_8 FILLER_11_1335 ();
 sg13g2_decap_8 FILLER_11_1342 ();
 sg13g2_decap_8 FILLER_11_1349 ();
 sg13g2_decap_8 FILLER_11_1356 ();
 sg13g2_decap_8 FILLER_11_1363 ();
 sg13g2_decap_8 FILLER_11_1370 ();
 sg13g2_decap_8 FILLER_11_1377 ();
 sg13g2_decap_8 FILLER_11_1384 ();
 sg13g2_decap_8 FILLER_11_1391 ();
 sg13g2_decap_8 FILLER_11_1398 ();
 sg13g2_decap_8 FILLER_11_1405 ();
 sg13g2_decap_8 FILLER_11_1412 ();
 sg13g2_decap_8 FILLER_11_1419 ();
 sg13g2_decap_8 FILLER_11_1426 ();
 sg13g2_decap_8 FILLER_11_1433 ();
 sg13g2_decap_8 FILLER_11_1440 ();
 sg13g2_decap_8 FILLER_11_1447 ();
 sg13g2_decap_8 FILLER_11_1454 ();
 sg13g2_decap_8 FILLER_11_1461 ();
 sg13g2_decap_8 FILLER_11_1468 ();
 sg13g2_decap_8 FILLER_11_1475 ();
 sg13g2_decap_8 FILLER_11_1482 ();
 sg13g2_decap_8 FILLER_11_1489 ();
 sg13g2_decap_8 FILLER_11_1496 ();
 sg13g2_decap_8 FILLER_11_1503 ();
 sg13g2_decap_8 FILLER_11_1510 ();
 sg13g2_decap_8 FILLER_11_1517 ();
 sg13g2_decap_8 FILLER_11_1524 ();
 sg13g2_decap_8 FILLER_11_1531 ();
 sg13g2_decap_8 FILLER_11_1538 ();
 sg13g2_decap_8 FILLER_11_1545 ();
 sg13g2_decap_8 FILLER_11_1552 ();
 sg13g2_decap_8 FILLER_11_1559 ();
 sg13g2_decap_8 FILLER_11_1566 ();
 sg13g2_decap_8 FILLER_11_1573 ();
 sg13g2_decap_8 FILLER_11_1580 ();
 sg13g2_decap_8 FILLER_11_1587 ();
 sg13g2_decap_8 FILLER_11_1594 ();
 sg13g2_decap_8 FILLER_11_1601 ();
 sg13g2_decap_8 FILLER_11_1608 ();
 sg13g2_decap_8 FILLER_11_1615 ();
 sg13g2_decap_8 FILLER_11_1622 ();
 sg13g2_decap_8 FILLER_11_1629 ();
 sg13g2_decap_8 FILLER_11_1636 ();
 sg13g2_decap_8 FILLER_11_1643 ();
 sg13g2_decap_8 FILLER_11_1650 ();
 sg13g2_decap_8 FILLER_11_1657 ();
 sg13g2_decap_8 FILLER_11_1664 ();
 sg13g2_decap_8 FILLER_11_1671 ();
 sg13g2_decap_8 FILLER_11_1678 ();
 sg13g2_decap_8 FILLER_11_1685 ();
 sg13g2_decap_8 FILLER_11_1692 ();
 sg13g2_decap_8 FILLER_11_1699 ();
 sg13g2_decap_8 FILLER_11_1706 ();
 sg13g2_decap_8 FILLER_11_1713 ();
 sg13g2_decap_8 FILLER_11_1720 ();
 sg13g2_decap_8 FILLER_11_1727 ();
 sg13g2_decap_8 FILLER_11_1734 ();
 sg13g2_decap_8 FILLER_11_1741 ();
 sg13g2_decap_8 FILLER_11_1748 ();
 sg13g2_decap_8 FILLER_11_1755 ();
 sg13g2_decap_4 FILLER_11_1762 ();
 sg13g2_fill_2 FILLER_11_1766 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_4 FILLER_12_56 ();
 sg13g2_fill_2 FILLER_12_60 ();
 sg13g2_fill_1 FILLER_12_71 ();
 sg13g2_fill_2 FILLER_12_82 ();
 sg13g2_fill_2 FILLER_12_136 ();
 sg13g2_fill_2 FILLER_12_173 ();
 sg13g2_fill_1 FILLER_12_211 ();
 sg13g2_fill_2 FILLER_12_236 ();
 sg13g2_fill_1 FILLER_12_238 ();
 sg13g2_fill_2 FILLER_12_279 ();
 sg13g2_fill_1 FILLER_12_281 ();
 sg13g2_fill_2 FILLER_12_290 ();
 sg13g2_fill_1 FILLER_12_292 ();
 sg13g2_fill_2 FILLER_12_307 ();
 sg13g2_fill_1 FILLER_12_309 ();
 sg13g2_fill_1 FILLER_12_379 ();
 sg13g2_fill_2 FILLER_12_420 ();
 sg13g2_fill_1 FILLER_12_422 ();
 sg13g2_fill_2 FILLER_12_440 ();
 sg13g2_fill_1 FILLER_12_442 ();
 sg13g2_fill_1 FILLER_12_530 ();
 sg13g2_fill_2 FILLER_12_581 ();
 sg13g2_fill_2 FILLER_12_623 ();
 sg13g2_fill_1 FILLER_12_625 ();
 sg13g2_fill_1 FILLER_12_652 ();
 sg13g2_fill_1 FILLER_12_689 ();
 sg13g2_fill_1 FILLER_12_705 ();
 sg13g2_fill_2 FILLER_12_718 ();
 sg13g2_decap_8 FILLER_12_729 ();
 sg13g2_fill_1 FILLER_12_762 ();
 sg13g2_fill_2 FILLER_12_833 ();
 sg13g2_fill_1 FILLER_12_835 ();
 sg13g2_fill_1 FILLER_12_840 ();
 sg13g2_fill_2 FILLER_12_891 ();
 sg13g2_fill_1 FILLER_12_893 ();
 sg13g2_fill_1 FILLER_12_899 ();
 sg13g2_fill_1 FILLER_12_919 ();
 sg13g2_fill_1 FILLER_12_946 ();
 sg13g2_fill_2 FILLER_12_961 ();
 sg13g2_fill_1 FILLER_12_963 ();
 sg13g2_decap_8 FILLER_12_974 ();
 sg13g2_decap_4 FILLER_12_981 ();
 sg13g2_decap_4 FILLER_12_994 ();
 sg13g2_fill_2 FILLER_12_1026 ();
 sg13g2_fill_1 FILLER_12_1028 ();
 sg13g2_decap_4 FILLER_12_1065 ();
 sg13g2_fill_2 FILLER_12_1069 ();
 sg13g2_fill_2 FILLER_12_1084 ();
 sg13g2_fill_2 FILLER_12_1091 ();
 sg13g2_fill_1 FILLER_12_1093 ();
 sg13g2_fill_2 FILLER_12_1099 ();
 sg13g2_fill_1 FILLER_12_1101 ();
 sg13g2_fill_2 FILLER_12_1111 ();
 sg13g2_decap_8 FILLER_12_1309 ();
 sg13g2_decap_8 FILLER_12_1316 ();
 sg13g2_decap_8 FILLER_12_1323 ();
 sg13g2_decap_8 FILLER_12_1330 ();
 sg13g2_decap_8 FILLER_12_1337 ();
 sg13g2_decap_8 FILLER_12_1344 ();
 sg13g2_decap_8 FILLER_12_1351 ();
 sg13g2_decap_8 FILLER_12_1358 ();
 sg13g2_decap_8 FILLER_12_1365 ();
 sg13g2_decap_8 FILLER_12_1372 ();
 sg13g2_decap_8 FILLER_12_1379 ();
 sg13g2_decap_8 FILLER_12_1386 ();
 sg13g2_decap_8 FILLER_12_1393 ();
 sg13g2_decap_8 FILLER_12_1400 ();
 sg13g2_decap_8 FILLER_12_1407 ();
 sg13g2_decap_8 FILLER_12_1414 ();
 sg13g2_decap_8 FILLER_12_1421 ();
 sg13g2_decap_8 FILLER_12_1428 ();
 sg13g2_decap_8 FILLER_12_1435 ();
 sg13g2_decap_8 FILLER_12_1442 ();
 sg13g2_decap_8 FILLER_12_1449 ();
 sg13g2_decap_8 FILLER_12_1456 ();
 sg13g2_decap_8 FILLER_12_1463 ();
 sg13g2_decap_8 FILLER_12_1470 ();
 sg13g2_decap_8 FILLER_12_1477 ();
 sg13g2_decap_8 FILLER_12_1484 ();
 sg13g2_decap_8 FILLER_12_1491 ();
 sg13g2_decap_8 FILLER_12_1498 ();
 sg13g2_decap_8 FILLER_12_1505 ();
 sg13g2_decap_8 FILLER_12_1512 ();
 sg13g2_decap_8 FILLER_12_1519 ();
 sg13g2_decap_8 FILLER_12_1526 ();
 sg13g2_decap_8 FILLER_12_1533 ();
 sg13g2_decap_8 FILLER_12_1540 ();
 sg13g2_decap_8 FILLER_12_1547 ();
 sg13g2_decap_8 FILLER_12_1554 ();
 sg13g2_decap_8 FILLER_12_1561 ();
 sg13g2_decap_8 FILLER_12_1568 ();
 sg13g2_decap_8 FILLER_12_1575 ();
 sg13g2_decap_8 FILLER_12_1582 ();
 sg13g2_decap_8 FILLER_12_1589 ();
 sg13g2_decap_8 FILLER_12_1596 ();
 sg13g2_decap_8 FILLER_12_1603 ();
 sg13g2_decap_8 FILLER_12_1610 ();
 sg13g2_decap_8 FILLER_12_1617 ();
 sg13g2_decap_8 FILLER_12_1624 ();
 sg13g2_decap_8 FILLER_12_1631 ();
 sg13g2_decap_8 FILLER_12_1638 ();
 sg13g2_decap_8 FILLER_12_1645 ();
 sg13g2_decap_8 FILLER_12_1652 ();
 sg13g2_decap_8 FILLER_12_1659 ();
 sg13g2_decap_8 FILLER_12_1666 ();
 sg13g2_decap_8 FILLER_12_1673 ();
 sg13g2_decap_8 FILLER_12_1680 ();
 sg13g2_decap_8 FILLER_12_1687 ();
 sg13g2_decap_8 FILLER_12_1694 ();
 sg13g2_decap_8 FILLER_12_1701 ();
 sg13g2_decap_8 FILLER_12_1708 ();
 sg13g2_decap_8 FILLER_12_1715 ();
 sg13g2_decap_8 FILLER_12_1722 ();
 sg13g2_decap_8 FILLER_12_1729 ();
 sg13g2_decap_8 FILLER_12_1736 ();
 sg13g2_decap_8 FILLER_12_1743 ();
 sg13g2_decap_8 FILLER_12_1750 ();
 sg13g2_decap_8 FILLER_12_1757 ();
 sg13g2_decap_4 FILLER_12_1764 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_4 FILLER_13_49 ();
 sg13g2_fill_2 FILLER_13_89 ();
 sg13g2_decap_4 FILLER_13_123 ();
 sg13g2_fill_1 FILLER_13_127 ();
 sg13g2_decap_8 FILLER_13_142 ();
 sg13g2_decap_4 FILLER_13_149 ();
 sg13g2_fill_1 FILLER_13_153 ();
 sg13g2_fill_1 FILLER_13_163 ();
 sg13g2_fill_2 FILLER_13_236 ();
 sg13g2_fill_1 FILLER_13_238 ();
 sg13g2_fill_2 FILLER_13_252 ();
 sg13g2_fill_2 FILLER_13_277 ();
 sg13g2_fill_1 FILLER_13_279 ();
 sg13g2_fill_2 FILLER_13_339 ();
 sg13g2_fill_1 FILLER_13_341 ();
 sg13g2_fill_1 FILLER_13_348 ();
 sg13g2_fill_2 FILLER_13_475 ();
 sg13g2_fill_1 FILLER_13_595 ();
 sg13g2_fill_1 FILLER_13_601 ();
 sg13g2_fill_2 FILLER_13_630 ();
 sg13g2_fill_1 FILLER_13_632 ();
 sg13g2_fill_1 FILLER_13_652 ();
 sg13g2_fill_1 FILLER_13_670 ();
 sg13g2_fill_1 FILLER_13_699 ();
 sg13g2_decap_8 FILLER_13_731 ();
 sg13g2_decap_8 FILLER_13_738 ();
 sg13g2_fill_2 FILLER_13_780 ();
 sg13g2_fill_1 FILLER_13_782 ();
 sg13g2_decap_4 FILLER_13_803 ();
 sg13g2_fill_2 FILLER_13_807 ();
 sg13g2_fill_2 FILLER_13_819 ();
 sg13g2_decap_4 FILLER_13_858 ();
 sg13g2_fill_2 FILLER_13_862 ();
 sg13g2_fill_2 FILLER_13_914 ();
 sg13g2_fill_1 FILLER_13_916 ();
 sg13g2_fill_2 FILLER_13_948 ();
 sg13g2_fill_1 FILLER_13_950 ();
 sg13g2_fill_2 FILLER_13_1031 ();
 sg13g2_decap_8 FILLER_13_1059 ();
 sg13g2_fill_2 FILLER_13_1083 ();
 sg13g2_fill_1 FILLER_13_1085 ();
 sg13g2_fill_2 FILLER_13_1097 ();
 sg13g2_fill_1 FILLER_13_1099 ();
 sg13g2_fill_2 FILLER_13_1115 ();
 sg13g2_fill_2 FILLER_13_1164 ();
 sg13g2_fill_1 FILLER_13_1166 ();
 sg13g2_fill_2 FILLER_13_1181 ();
 sg13g2_fill_1 FILLER_13_1183 ();
 sg13g2_fill_2 FILLER_13_1198 ();
 sg13g2_fill_1 FILLER_13_1259 ();
 sg13g2_decap_8 FILLER_13_1304 ();
 sg13g2_decap_8 FILLER_13_1311 ();
 sg13g2_decap_8 FILLER_13_1318 ();
 sg13g2_decap_8 FILLER_13_1325 ();
 sg13g2_decap_8 FILLER_13_1332 ();
 sg13g2_decap_8 FILLER_13_1339 ();
 sg13g2_decap_8 FILLER_13_1346 ();
 sg13g2_decap_8 FILLER_13_1353 ();
 sg13g2_decap_8 FILLER_13_1360 ();
 sg13g2_decap_8 FILLER_13_1367 ();
 sg13g2_decap_8 FILLER_13_1374 ();
 sg13g2_decap_8 FILLER_13_1381 ();
 sg13g2_decap_8 FILLER_13_1388 ();
 sg13g2_decap_8 FILLER_13_1395 ();
 sg13g2_decap_8 FILLER_13_1402 ();
 sg13g2_decap_8 FILLER_13_1409 ();
 sg13g2_decap_8 FILLER_13_1416 ();
 sg13g2_decap_8 FILLER_13_1423 ();
 sg13g2_decap_8 FILLER_13_1430 ();
 sg13g2_decap_8 FILLER_13_1437 ();
 sg13g2_decap_8 FILLER_13_1444 ();
 sg13g2_decap_8 FILLER_13_1451 ();
 sg13g2_decap_8 FILLER_13_1458 ();
 sg13g2_decap_8 FILLER_13_1465 ();
 sg13g2_decap_8 FILLER_13_1472 ();
 sg13g2_decap_8 FILLER_13_1479 ();
 sg13g2_decap_8 FILLER_13_1486 ();
 sg13g2_decap_8 FILLER_13_1493 ();
 sg13g2_decap_8 FILLER_13_1500 ();
 sg13g2_decap_8 FILLER_13_1507 ();
 sg13g2_decap_8 FILLER_13_1514 ();
 sg13g2_decap_8 FILLER_13_1521 ();
 sg13g2_decap_8 FILLER_13_1528 ();
 sg13g2_decap_8 FILLER_13_1535 ();
 sg13g2_decap_8 FILLER_13_1542 ();
 sg13g2_decap_8 FILLER_13_1549 ();
 sg13g2_decap_8 FILLER_13_1556 ();
 sg13g2_decap_8 FILLER_13_1563 ();
 sg13g2_decap_8 FILLER_13_1570 ();
 sg13g2_decap_8 FILLER_13_1577 ();
 sg13g2_decap_8 FILLER_13_1584 ();
 sg13g2_decap_8 FILLER_13_1591 ();
 sg13g2_decap_8 FILLER_13_1598 ();
 sg13g2_decap_8 FILLER_13_1605 ();
 sg13g2_decap_8 FILLER_13_1612 ();
 sg13g2_decap_8 FILLER_13_1619 ();
 sg13g2_decap_8 FILLER_13_1626 ();
 sg13g2_decap_8 FILLER_13_1633 ();
 sg13g2_decap_8 FILLER_13_1640 ();
 sg13g2_decap_8 FILLER_13_1647 ();
 sg13g2_decap_8 FILLER_13_1654 ();
 sg13g2_decap_8 FILLER_13_1661 ();
 sg13g2_decap_8 FILLER_13_1668 ();
 sg13g2_decap_8 FILLER_13_1675 ();
 sg13g2_decap_8 FILLER_13_1682 ();
 sg13g2_decap_8 FILLER_13_1689 ();
 sg13g2_decap_8 FILLER_13_1696 ();
 sg13g2_decap_8 FILLER_13_1703 ();
 sg13g2_decap_8 FILLER_13_1710 ();
 sg13g2_decap_8 FILLER_13_1717 ();
 sg13g2_decap_8 FILLER_13_1724 ();
 sg13g2_decap_8 FILLER_13_1731 ();
 sg13g2_decap_8 FILLER_13_1738 ();
 sg13g2_decap_8 FILLER_13_1745 ();
 sg13g2_decap_8 FILLER_13_1752 ();
 sg13g2_decap_8 FILLER_13_1759 ();
 sg13g2_fill_2 FILLER_13_1766 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_fill_2 FILLER_14_42 ();
 sg13g2_fill_1 FILLER_14_88 ();
 sg13g2_fill_2 FILLER_14_109 ();
 sg13g2_fill_1 FILLER_14_111 ();
 sg13g2_fill_2 FILLER_14_143 ();
 sg13g2_fill_1 FILLER_14_180 ();
 sg13g2_fill_2 FILLER_14_233 ();
 sg13g2_fill_2 FILLER_14_245 ();
 sg13g2_fill_2 FILLER_14_317 ();
 sg13g2_fill_1 FILLER_14_319 ();
 sg13g2_fill_2 FILLER_14_370 ();
 sg13g2_fill_1 FILLER_14_384 ();
 sg13g2_fill_2 FILLER_14_393 ();
 sg13g2_fill_2 FILLER_14_403 ();
 sg13g2_fill_2 FILLER_14_428 ();
 sg13g2_fill_1 FILLER_14_430 ();
 sg13g2_fill_1 FILLER_14_457 ();
 sg13g2_fill_2 FILLER_14_471 ();
 sg13g2_fill_1 FILLER_14_504 ();
 sg13g2_fill_2 FILLER_14_529 ();
 sg13g2_fill_1 FILLER_14_696 ();
 sg13g2_fill_2 FILLER_14_707 ();
 sg13g2_decap_8 FILLER_14_740 ();
 sg13g2_fill_2 FILLER_14_747 ();
 sg13g2_fill_1 FILLER_14_749 ();
 sg13g2_fill_2 FILLER_14_772 ();
 sg13g2_fill_1 FILLER_14_774 ();
 sg13g2_fill_1 FILLER_14_793 ();
 sg13g2_fill_2 FILLER_14_798 ();
 sg13g2_fill_2 FILLER_14_814 ();
 sg13g2_fill_1 FILLER_14_816 ();
 sg13g2_fill_2 FILLER_14_827 ();
 sg13g2_fill_1 FILLER_14_847 ();
 sg13g2_fill_1 FILLER_14_863 ();
 sg13g2_fill_2 FILLER_14_872 ();
 sg13g2_decap_8 FILLER_14_886 ();
 sg13g2_decap_4 FILLER_14_893 ();
 sg13g2_fill_1 FILLER_14_897 ();
 sg13g2_fill_1 FILLER_14_949 ();
 sg13g2_fill_2 FILLER_14_974 ();
 sg13g2_decap_4 FILLER_14_989 ();
 sg13g2_fill_1 FILLER_14_993 ();
 sg13g2_fill_1 FILLER_14_1019 ();
 sg13g2_fill_2 FILLER_14_1061 ();
 sg13g2_fill_1 FILLER_14_1098 ();
 sg13g2_fill_2 FILLER_14_1204 ();
 sg13g2_fill_1 FILLER_14_1206 ();
 sg13g2_fill_2 FILLER_14_1234 ();
 sg13g2_fill_1 FILLER_14_1236 ();
 sg13g2_decap_8 FILLER_14_1304 ();
 sg13g2_decap_8 FILLER_14_1311 ();
 sg13g2_decap_8 FILLER_14_1318 ();
 sg13g2_decap_8 FILLER_14_1325 ();
 sg13g2_decap_8 FILLER_14_1332 ();
 sg13g2_decap_8 FILLER_14_1339 ();
 sg13g2_decap_8 FILLER_14_1346 ();
 sg13g2_decap_8 FILLER_14_1353 ();
 sg13g2_decap_8 FILLER_14_1360 ();
 sg13g2_decap_8 FILLER_14_1367 ();
 sg13g2_decap_8 FILLER_14_1374 ();
 sg13g2_decap_8 FILLER_14_1381 ();
 sg13g2_decap_8 FILLER_14_1388 ();
 sg13g2_decap_8 FILLER_14_1395 ();
 sg13g2_decap_8 FILLER_14_1402 ();
 sg13g2_decap_8 FILLER_14_1409 ();
 sg13g2_decap_8 FILLER_14_1416 ();
 sg13g2_decap_8 FILLER_14_1423 ();
 sg13g2_decap_8 FILLER_14_1430 ();
 sg13g2_decap_8 FILLER_14_1437 ();
 sg13g2_decap_8 FILLER_14_1444 ();
 sg13g2_decap_8 FILLER_14_1451 ();
 sg13g2_decap_8 FILLER_14_1458 ();
 sg13g2_decap_8 FILLER_14_1465 ();
 sg13g2_decap_8 FILLER_14_1472 ();
 sg13g2_decap_8 FILLER_14_1479 ();
 sg13g2_decap_8 FILLER_14_1486 ();
 sg13g2_decap_8 FILLER_14_1493 ();
 sg13g2_decap_8 FILLER_14_1500 ();
 sg13g2_decap_8 FILLER_14_1507 ();
 sg13g2_decap_8 FILLER_14_1514 ();
 sg13g2_decap_8 FILLER_14_1521 ();
 sg13g2_decap_8 FILLER_14_1528 ();
 sg13g2_decap_8 FILLER_14_1535 ();
 sg13g2_decap_8 FILLER_14_1542 ();
 sg13g2_decap_8 FILLER_14_1549 ();
 sg13g2_decap_8 FILLER_14_1556 ();
 sg13g2_decap_8 FILLER_14_1563 ();
 sg13g2_decap_8 FILLER_14_1570 ();
 sg13g2_decap_8 FILLER_14_1577 ();
 sg13g2_decap_8 FILLER_14_1584 ();
 sg13g2_decap_8 FILLER_14_1591 ();
 sg13g2_decap_8 FILLER_14_1598 ();
 sg13g2_decap_8 FILLER_14_1605 ();
 sg13g2_decap_8 FILLER_14_1612 ();
 sg13g2_decap_8 FILLER_14_1619 ();
 sg13g2_decap_8 FILLER_14_1626 ();
 sg13g2_decap_8 FILLER_14_1633 ();
 sg13g2_decap_8 FILLER_14_1640 ();
 sg13g2_decap_8 FILLER_14_1647 ();
 sg13g2_decap_8 FILLER_14_1654 ();
 sg13g2_decap_8 FILLER_14_1661 ();
 sg13g2_decap_8 FILLER_14_1668 ();
 sg13g2_decap_8 FILLER_14_1675 ();
 sg13g2_decap_8 FILLER_14_1682 ();
 sg13g2_decap_8 FILLER_14_1689 ();
 sg13g2_decap_8 FILLER_14_1696 ();
 sg13g2_decap_8 FILLER_14_1703 ();
 sg13g2_decap_8 FILLER_14_1710 ();
 sg13g2_decap_8 FILLER_14_1717 ();
 sg13g2_decap_8 FILLER_14_1724 ();
 sg13g2_decap_8 FILLER_14_1731 ();
 sg13g2_decap_8 FILLER_14_1738 ();
 sg13g2_decap_8 FILLER_14_1745 ();
 sg13g2_decap_8 FILLER_14_1752 ();
 sg13g2_decap_8 FILLER_14_1759 ();
 sg13g2_fill_2 FILLER_14_1766 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_4 FILLER_15_28 ();
 sg13g2_fill_1 FILLER_15_32 ();
 sg13g2_fill_2 FILLER_15_86 ();
 sg13g2_decap_8 FILLER_15_120 ();
 sg13g2_fill_2 FILLER_15_150 ();
 sg13g2_fill_1 FILLER_15_152 ();
 sg13g2_fill_1 FILLER_15_167 ();
 sg13g2_fill_1 FILLER_15_187 ();
 sg13g2_fill_1 FILLER_15_196 ();
 sg13g2_fill_2 FILLER_15_216 ();
 sg13g2_fill_2 FILLER_15_242 ();
 sg13g2_decap_8 FILLER_15_280 ();
 sg13g2_decap_4 FILLER_15_292 ();
 sg13g2_fill_2 FILLER_15_296 ();
 sg13g2_fill_2 FILLER_15_314 ();
 sg13g2_fill_1 FILLER_15_388 ();
 sg13g2_fill_1 FILLER_15_419 ();
 sg13g2_decap_8 FILLER_15_424 ();
 sg13g2_fill_2 FILLER_15_431 ();
 sg13g2_decap_8 FILLER_15_444 ();
 sg13g2_decap_4 FILLER_15_456 ();
 sg13g2_fill_2 FILLER_15_460 ();
 sg13g2_fill_2 FILLER_15_514 ();
 sg13g2_fill_1 FILLER_15_528 ();
 sg13g2_fill_1 FILLER_15_568 ();
 sg13g2_fill_2 FILLER_15_579 ();
 sg13g2_fill_2 FILLER_15_633 ();
 sg13g2_fill_1 FILLER_15_635 ();
 sg13g2_fill_2 FILLER_15_664 ();
 sg13g2_fill_2 FILLER_15_674 ();
 sg13g2_fill_1 FILLER_15_690 ();
 sg13g2_fill_2 FILLER_15_794 ();
 sg13g2_fill_2 FILLER_15_824 ();
 sg13g2_fill_1 FILLER_15_826 ();
 sg13g2_fill_2 FILLER_15_872 ();
 sg13g2_fill_2 FILLER_15_919 ();
 sg13g2_fill_2 FILLER_15_926 ();
 sg13g2_fill_2 FILLER_15_940 ();
 sg13g2_fill_1 FILLER_15_942 ();
 sg13g2_fill_2 FILLER_15_964 ();
 sg13g2_fill_1 FILLER_15_992 ();
 sg13g2_fill_2 FILLER_15_1012 ();
 sg13g2_fill_1 FILLER_15_1014 ();
 sg13g2_fill_2 FILLER_15_1037 ();
 sg13g2_decap_4 FILLER_15_1081 ();
 sg13g2_fill_2 FILLER_15_1095 ();
 sg13g2_fill_2 FILLER_15_1106 ();
 sg13g2_fill_1 FILLER_15_1108 ();
 sg13g2_fill_2 FILLER_15_1146 ();
 sg13g2_fill_1 FILLER_15_1148 ();
 sg13g2_fill_1 FILLER_15_1235 ();
 sg13g2_fill_1 FILLER_15_1273 ();
 sg13g2_decap_8 FILLER_15_1295 ();
 sg13g2_decap_8 FILLER_15_1302 ();
 sg13g2_decap_8 FILLER_15_1309 ();
 sg13g2_decap_8 FILLER_15_1316 ();
 sg13g2_decap_8 FILLER_15_1323 ();
 sg13g2_decap_8 FILLER_15_1330 ();
 sg13g2_decap_8 FILLER_15_1337 ();
 sg13g2_decap_8 FILLER_15_1344 ();
 sg13g2_decap_8 FILLER_15_1351 ();
 sg13g2_decap_8 FILLER_15_1358 ();
 sg13g2_decap_8 FILLER_15_1365 ();
 sg13g2_decap_8 FILLER_15_1372 ();
 sg13g2_decap_8 FILLER_15_1379 ();
 sg13g2_decap_8 FILLER_15_1386 ();
 sg13g2_decap_8 FILLER_15_1393 ();
 sg13g2_decap_8 FILLER_15_1400 ();
 sg13g2_decap_8 FILLER_15_1407 ();
 sg13g2_decap_8 FILLER_15_1414 ();
 sg13g2_decap_8 FILLER_15_1421 ();
 sg13g2_decap_8 FILLER_15_1428 ();
 sg13g2_decap_8 FILLER_15_1435 ();
 sg13g2_decap_8 FILLER_15_1442 ();
 sg13g2_decap_8 FILLER_15_1449 ();
 sg13g2_decap_8 FILLER_15_1456 ();
 sg13g2_decap_8 FILLER_15_1463 ();
 sg13g2_decap_8 FILLER_15_1470 ();
 sg13g2_decap_8 FILLER_15_1477 ();
 sg13g2_decap_8 FILLER_15_1484 ();
 sg13g2_decap_8 FILLER_15_1491 ();
 sg13g2_decap_8 FILLER_15_1498 ();
 sg13g2_decap_8 FILLER_15_1505 ();
 sg13g2_decap_8 FILLER_15_1512 ();
 sg13g2_decap_8 FILLER_15_1519 ();
 sg13g2_decap_8 FILLER_15_1526 ();
 sg13g2_decap_8 FILLER_15_1533 ();
 sg13g2_decap_8 FILLER_15_1540 ();
 sg13g2_decap_8 FILLER_15_1547 ();
 sg13g2_decap_8 FILLER_15_1554 ();
 sg13g2_decap_8 FILLER_15_1561 ();
 sg13g2_decap_8 FILLER_15_1568 ();
 sg13g2_decap_8 FILLER_15_1575 ();
 sg13g2_decap_8 FILLER_15_1582 ();
 sg13g2_decap_8 FILLER_15_1589 ();
 sg13g2_decap_8 FILLER_15_1596 ();
 sg13g2_decap_8 FILLER_15_1603 ();
 sg13g2_decap_8 FILLER_15_1610 ();
 sg13g2_decap_8 FILLER_15_1617 ();
 sg13g2_decap_8 FILLER_15_1624 ();
 sg13g2_decap_8 FILLER_15_1631 ();
 sg13g2_decap_8 FILLER_15_1638 ();
 sg13g2_decap_8 FILLER_15_1645 ();
 sg13g2_decap_8 FILLER_15_1652 ();
 sg13g2_decap_8 FILLER_15_1659 ();
 sg13g2_decap_8 FILLER_15_1666 ();
 sg13g2_decap_8 FILLER_15_1673 ();
 sg13g2_decap_8 FILLER_15_1680 ();
 sg13g2_decap_8 FILLER_15_1687 ();
 sg13g2_decap_8 FILLER_15_1694 ();
 sg13g2_decap_8 FILLER_15_1701 ();
 sg13g2_decap_8 FILLER_15_1708 ();
 sg13g2_decap_8 FILLER_15_1715 ();
 sg13g2_decap_8 FILLER_15_1722 ();
 sg13g2_decap_8 FILLER_15_1729 ();
 sg13g2_decap_8 FILLER_15_1736 ();
 sg13g2_decap_8 FILLER_15_1743 ();
 sg13g2_decap_8 FILLER_15_1750 ();
 sg13g2_decap_8 FILLER_15_1757 ();
 sg13g2_decap_4 FILLER_15_1764 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_fill_2 FILLER_16_28 ();
 sg13g2_fill_1 FILLER_16_30 ();
 sg13g2_fill_1 FILLER_16_76 ();
 sg13g2_fill_1 FILLER_16_108 ();
 sg13g2_decap_8 FILLER_16_139 ();
 sg13g2_fill_1 FILLER_16_146 ();
 sg13g2_fill_2 FILLER_16_221 ();
 sg13g2_fill_1 FILLER_16_230 ();
 sg13g2_fill_1 FILLER_16_269 ();
 sg13g2_decap_4 FILLER_16_289 ();
 sg13g2_fill_1 FILLER_16_293 ();
 sg13g2_decap_8 FILLER_16_299 ();
 sg13g2_fill_2 FILLER_16_306 ();
 sg13g2_fill_1 FILLER_16_323 ();
 sg13g2_decap_4 FILLER_16_338 ();
 sg13g2_decap_4 FILLER_16_357 ();
 sg13g2_fill_1 FILLER_16_361 ();
 sg13g2_fill_1 FILLER_16_366 ();
 sg13g2_fill_2 FILLER_16_378 ();
 sg13g2_fill_2 FILLER_16_385 ();
 sg13g2_fill_1 FILLER_16_387 ();
 sg13g2_fill_2 FILLER_16_420 ();
 sg13g2_decap_4 FILLER_16_427 ();
 sg13g2_fill_2 FILLER_16_431 ();
 sg13g2_fill_2 FILLER_16_470 ();
 sg13g2_fill_1 FILLER_16_472 ();
 sg13g2_fill_2 FILLER_16_481 ();
 sg13g2_fill_1 FILLER_16_483 ();
 sg13g2_fill_1 FILLER_16_535 ();
 sg13g2_fill_2 FILLER_16_619 ();
 sg13g2_fill_1 FILLER_16_621 ();
 sg13g2_fill_1 FILLER_16_652 ();
 sg13g2_fill_2 FILLER_16_714 ();
 sg13g2_fill_1 FILLER_16_716 ();
 sg13g2_fill_2 FILLER_16_726 ();
 sg13g2_fill_2 FILLER_16_741 ();
 sg13g2_fill_1 FILLER_16_743 ();
 sg13g2_decap_8 FILLER_16_752 ();
 sg13g2_fill_1 FILLER_16_759 ();
 sg13g2_fill_2 FILLER_16_765 ();
 sg13g2_fill_2 FILLER_16_772 ();
 sg13g2_fill_1 FILLER_16_774 ();
 sg13g2_fill_1 FILLER_16_863 ();
 sg13g2_decap_8 FILLER_16_883 ();
 sg13g2_decap_8 FILLER_16_890 ();
 sg13g2_fill_2 FILLER_16_897 ();
 sg13g2_fill_1 FILLER_16_899 ();
 sg13g2_decap_4 FILLER_16_905 ();
 sg13g2_fill_2 FILLER_16_952 ();
 sg13g2_fill_1 FILLER_16_954 ();
 sg13g2_fill_2 FILLER_16_991 ();
 sg13g2_decap_4 FILLER_16_1056 ();
 sg13g2_fill_1 FILLER_16_1060 ();
 sg13g2_fill_1 FILLER_16_1088 ();
 sg13g2_fill_1 FILLER_16_1139 ();
 sg13g2_fill_2 FILLER_16_1149 ();
 sg13g2_fill_1 FILLER_16_1151 ();
 sg13g2_fill_1 FILLER_16_1157 ();
 sg13g2_fill_2 FILLER_16_1168 ();
 sg13g2_fill_2 FILLER_16_1175 ();
 sg13g2_fill_1 FILLER_16_1177 ();
 sg13g2_fill_2 FILLER_16_1215 ();
 sg13g2_fill_2 FILLER_16_1271 ();
 sg13g2_decap_8 FILLER_16_1299 ();
 sg13g2_decap_8 FILLER_16_1306 ();
 sg13g2_decap_8 FILLER_16_1313 ();
 sg13g2_decap_8 FILLER_16_1320 ();
 sg13g2_decap_8 FILLER_16_1327 ();
 sg13g2_decap_8 FILLER_16_1334 ();
 sg13g2_decap_8 FILLER_16_1341 ();
 sg13g2_decap_8 FILLER_16_1348 ();
 sg13g2_decap_8 FILLER_16_1355 ();
 sg13g2_decap_8 FILLER_16_1362 ();
 sg13g2_decap_8 FILLER_16_1369 ();
 sg13g2_decap_8 FILLER_16_1376 ();
 sg13g2_decap_8 FILLER_16_1383 ();
 sg13g2_decap_8 FILLER_16_1390 ();
 sg13g2_decap_8 FILLER_16_1397 ();
 sg13g2_decap_8 FILLER_16_1404 ();
 sg13g2_decap_8 FILLER_16_1411 ();
 sg13g2_decap_8 FILLER_16_1418 ();
 sg13g2_decap_8 FILLER_16_1425 ();
 sg13g2_decap_8 FILLER_16_1432 ();
 sg13g2_decap_8 FILLER_16_1439 ();
 sg13g2_decap_8 FILLER_16_1446 ();
 sg13g2_decap_8 FILLER_16_1453 ();
 sg13g2_decap_8 FILLER_16_1460 ();
 sg13g2_decap_8 FILLER_16_1467 ();
 sg13g2_decap_8 FILLER_16_1474 ();
 sg13g2_decap_8 FILLER_16_1481 ();
 sg13g2_decap_8 FILLER_16_1488 ();
 sg13g2_decap_8 FILLER_16_1495 ();
 sg13g2_decap_8 FILLER_16_1502 ();
 sg13g2_decap_8 FILLER_16_1509 ();
 sg13g2_decap_8 FILLER_16_1516 ();
 sg13g2_decap_8 FILLER_16_1523 ();
 sg13g2_decap_8 FILLER_16_1530 ();
 sg13g2_decap_8 FILLER_16_1537 ();
 sg13g2_decap_8 FILLER_16_1544 ();
 sg13g2_decap_8 FILLER_16_1551 ();
 sg13g2_decap_8 FILLER_16_1558 ();
 sg13g2_decap_8 FILLER_16_1565 ();
 sg13g2_decap_8 FILLER_16_1572 ();
 sg13g2_decap_8 FILLER_16_1579 ();
 sg13g2_decap_8 FILLER_16_1586 ();
 sg13g2_decap_8 FILLER_16_1593 ();
 sg13g2_decap_8 FILLER_16_1600 ();
 sg13g2_decap_8 FILLER_16_1607 ();
 sg13g2_decap_8 FILLER_16_1614 ();
 sg13g2_decap_8 FILLER_16_1621 ();
 sg13g2_decap_8 FILLER_16_1628 ();
 sg13g2_decap_8 FILLER_16_1635 ();
 sg13g2_decap_8 FILLER_16_1642 ();
 sg13g2_decap_8 FILLER_16_1649 ();
 sg13g2_decap_8 FILLER_16_1656 ();
 sg13g2_decap_8 FILLER_16_1663 ();
 sg13g2_decap_8 FILLER_16_1670 ();
 sg13g2_decap_8 FILLER_16_1677 ();
 sg13g2_decap_8 FILLER_16_1684 ();
 sg13g2_decap_8 FILLER_16_1691 ();
 sg13g2_decap_8 FILLER_16_1698 ();
 sg13g2_decap_8 FILLER_16_1705 ();
 sg13g2_decap_8 FILLER_16_1712 ();
 sg13g2_decap_8 FILLER_16_1719 ();
 sg13g2_decap_8 FILLER_16_1726 ();
 sg13g2_decap_8 FILLER_16_1733 ();
 sg13g2_decap_8 FILLER_16_1740 ();
 sg13g2_decap_8 FILLER_16_1747 ();
 sg13g2_decap_8 FILLER_16_1754 ();
 sg13g2_decap_8 FILLER_16_1761 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_fill_2 FILLER_17_28 ();
 sg13g2_fill_2 FILLER_17_56 ();
 sg13g2_fill_1 FILLER_17_58 ();
 sg13g2_fill_2 FILLER_17_73 ();
 sg13g2_fill_1 FILLER_17_75 ();
 sg13g2_fill_2 FILLER_17_86 ();
 sg13g2_fill_1 FILLER_17_98 ();
 sg13g2_fill_2 FILLER_17_104 ();
 sg13g2_fill_1 FILLER_17_106 ();
 sg13g2_fill_1 FILLER_17_117 ();
 sg13g2_fill_2 FILLER_17_123 ();
 sg13g2_fill_2 FILLER_17_165 ();
 sg13g2_fill_1 FILLER_17_181 ();
 sg13g2_fill_1 FILLER_17_217 ();
 sg13g2_fill_1 FILLER_17_237 ();
 sg13g2_fill_2 FILLER_17_322 ();
 sg13g2_fill_1 FILLER_17_324 ();
 sg13g2_decap_4 FILLER_17_335 ();
 sg13g2_decap_4 FILLER_17_360 ();
 sg13g2_fill_1 FILLER_17_364 ();
 sg13g2_fill_1 FILLER_17_380 ();
 sg13g2_decap_4 FILLER_17_387 ();
 sg13g2_fill_2 FILLER_17_422 ();
 sg13g2_fill_2 FILLER_17_434 ();
 sg13g2_fill_1 FILLER_17_436 ();
 sg13g2_fill_2 FILLER_17_468 ();
 sg13g2_fill_1 FILLER_17_470 ();
 sg13g2_fill_2 FILLER_17_490 ();
 sg13g2_fill_2 FILLER_17_501 ();
 sg13g2_fill_2 FILLER_17_512 ();
 sg13g2_fill_2 FILLER_17_520 ();
 sg13g2_fill_1 FILLER_17_522 ();
 sg13g2_fill_2 FILLER_17_555 ();
 sg13g2_fill_1 FILLER_17_574 ();
 sg13g2_fill_1 FILLER_17_589 ();
 sg13g2_fill_1 FILLER_17_609 ();
 sg13g2_fill_1 FILLER_17_656 ();
 sg13g2_fill_2 FILLER_17_675 ();
 sg13g2_fill_1 FILLER_17_726 ();
 sg13g2_fill_1 FILLER_17_815 ();
 sg13g2_fill_2 FILLER_17_834 ();
 sg13g2_fill_2 FILLER_17_919 ();
 sg13g2_fill_1 FILLER_17_921 ();
 sg13g2_decap_8 FILLER_17_987 ();
 sg13g2_decap_4 FILLER_17_994 ();
 sg13g2_decap_8 FILLER_17_1007 ();
 sg13g2_decap_4 FILLER_17_1019 ();
 sg13g2_decap_8 FILLER_17_1048 ();
 sg13g2_decap_4 FILLER_17_1055 ();
 sg13g2_fill_1 FILLER_17_1112 ();
 sg13g2_fill_2 FILLER_17_1122 ();
 sg13g2_fill_2 FILLER_17_1150 ();
 sg13g2_fill_1 FILLER_17_1152 ();
 sg13g2_fill_2 FILLER_17_1236 ();
 sg13g2_fill_1 FILLER_17_1238 ();
 sg13g2_decap_8 FILLER_17_1291 ();
 sg13g2_decap_8 FILLER_17_1298 ();
 sg13g2_decap_8 FILLER_17_1305 ();
 sg13g2_decap_8 FILLER_17_1312 ();
 sg13g2_decap_8 FILLER_17_1319 ();
 sg13g2_decap_8 FILLER_17_1326 ();
 sg13g2_decap_8 FILLER_17_1333 ();
 sg13g2_decap_8 FILLER_17_1340 ();
 sg13g2_decap_8 FILLER_17_1347 ();
 sg13g2_decap_8 FILLER_17_1354 ();
 sg13g2_decap_8 FILLER_17_1361 ();
 sg13g2_decap_8 FILLER_17_1368 ();
 sg13g2_decap_8 FILLER_17_1375 ();
 sg13g2_decap_8 FILLER_17_1382 ();
 sg13g2_decap_8 FILLER_17_1389 ();
 sg13g2_decap_8 FILLER_17_1396 ();
 sg13g2_decap_8 FILLER_17_1403 ();
 sg13g2_decap_8 FILLER_17_1410 ();
 sg13g2_decap_8 FILLER_17_1417 ();
 sg13g2_decap_8 FILLER_17_1424 ();
 sg13g2_decap_8 FILLER_17_1431 ();
 sg13g2_decap_8 FILLER_17_1438 ();
 sg13g2_decap_8 FILLER_17_1445 ();
 sg13g2_decap_8 FILLER_17_1452 ();
 sg13g2_decap_8 FILLER_17_1459 ();
 sg13g2_decap_8 FILLER_17_1466 ();
 sg13g2_decap_8 FILLER_17_1473 ();
 sg13g2_decap_8 FILLER_17_1480 ();
 sg13g2_decap_8 FILLER_17_1487 ();
 sg13g2_decap_8 FILLER_17_1494 ();
 sg13g2_decap_8 FILLER_17_1501 ();
 sg13g2_decap_8 FILLER_17_1508 ();
 sg13g2_decap_8 FILLER_17_1515 ();
 sg13g2_decap_8 FILLER_17_1522 ();
 sg13g2_decap_8 FILLER_17_1529 ();
 sg13g2_decap_8 FILLER_17_1536 ();
 sg13g2_decap_8 FILLER_17_1543 ();
 sg13g2_decap_8 FILLER_17_1550 ();
 sg13g2_decap_8 FILLER_17_1557 ();
 sg13g2_decap_8 FILLER_17_1564 ();
 sg13g2_decap_8 FILLER_17_1571 ();
 sg13g2_decap_8 FILLER_17_1578 ();
 sg13g2_decap_8 FILLER_17_1585 ();
 sg13g2_decap_8 FILLER_17_1592 ();
 sg13g2_decap_8 FILLER_17_1599 ();
 sg13g2_decap_8 FILLER_17_1606 ();
 sg13g2_decap_8 FILLER_17_1613 ();
 sg13g2_decap_8 FILLER_17_1620 ();
 sg13g2_decap_8 FILLER_17_1627 ();
 sg13g2_decap_8 FILLER_17_1634 ();
 sg13g2_decap_8 FILLER_17_1641 ();
 sg13g2_decap_8 FILLER_17_1648 ();
 sg13g2_decap_8 FILLER_17_1655 ();
 sg13g2_decap_8 FILLER_17_1662 ();
 sg13g2_decap_8 FILLER_17_1669 ();
 sg13g2_decap_8 FILLER_17_1676 ();
 sg13g2_decap_8 FILLER_17_1683 ();
 sg13g2_decap_8 FILLER_17_1690 ();
 sg13g2_decap_8 FILLER_17_1697 ();
 sg13g2_decap_8 FILLER_17_1704 ();
 sg13g2_decap_8 FILLER_17_1711 ();
 sg13g2_decap_8 FILLER_17_1718 ();
 sg13g2_decap_8 FILLER_17_1725 ();
 sg13g2_decap_8 FILLER_17_1732 ();
 sg13g2_decap_8 FILLER_17_1739 ();
 sg13g2_decap_8 FILLER_17_1746 ();
 sg13g2_decap_8 FILLER_17_1753 ();
 sg13g2_decap_8 FILLER_17_1760 ();
 sg13g2_fill_1 FILLER_17_1767 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_4 FILLER_18_35 ();
 sg13g2_fill_2 FILLER_18_70 ();
 sg13g2_fill_2 FILLER_18_91 ();
 sg13g2_fill_1 FILLER_18_93 ();
 sg13g2_fill_2 FILLER_18_104 ();
 sg13g2_fill_2 FILLER_18_148 ();
 sg13g2_fill_2 FILLER_18_155 ();
 sg13g2_fill_1 FILLER_18_157 ();
 sg13g2_fill_2 FILLER_18_162 ();
 sg13g2_fill_1 FILLER_18_181 ();
 sg13g2_fill_2 FILLER_18_216 ();
 sg13g2_fill_1 FILLER_18_218 ();
 sg13g2_fill_1 FILLER_18_238 ();
 sg13g2_fill_2 FILLER_18_265 ();
 sg13g2_fill_1 FILLER_18_276 ();
 sg13g2_fill_1 FILLER_18_282 ();
 sg13g2_fill_2 FILLER_18_288 ();
 sg13g2_decap_4 FILLER_18_305 ();
 sg13g2_decap_8 FILLER_18_335 ();
 sg13g2_fill_1 FILLER_18_342 ();
 sg13g2_decap_4 FILLER_18_358 ();
 sg13g2_fill_1 FILLER_18_385 ();
 sg13g2_decap_8 FILLER_18_410 ();
 sg13g2_fill_2 FILLER_18_422 ();
 sg13g2_fill_2 FILLER_18_439 ();
 sg13g2_decap_8 FILLER_18_447 ();
 sg13g2_fill_1 FILLER_18_477 ();
 sg13g2_fill_1 FILLER_18_502 ();
 sg13g2_fill_2 FILLER_18_515 ();
 sg13g2_fill_2 FILLER_18_531 ();
 sg13g2_fill_2 FILLER_18_541 ();
 sg13g2_fill_1 FILLER_18_556 ();
 sg13g2_fill_1 FILLER_18_562 ();
 sg13g2_fill_2 FILLER_18_573 ();
 sg13g2_fill_1 FILLER_18_575 ();
 sg13g2_fill_2 FILLER_18_584 ();
 sg13g2_fill_2 FILLER_18_626 ();
 sg13g2_fill_1 FILLER_18_646 ();
 sg13g2_fill_2 FILLER_18_728 ();
 sg13g2_fill_2 FILLER_18_738 ();
 sg13g2_fill_1 FILLER_18_740 ();
 sg13g2_fill_2 FILLER_18_759 ();
 sg13g2_fill_1 FILLER_18_761 ();
 sg13g2_decap_8 FILLER_18_766 ();
 sg13g2_decap_4 FILLER_18_773 ();
 sg13g2_fill_2 FILLER_18_777 ();
 sg13g2_fill_1 FILLER_18_791 ();
 sg13g2_fill_2 FILLER_18_827 ();
 sg13g2_fill_1 FILLER_18_848 ();
 sg13g2_decap_4 FILLER_18_860 ();
 sg13g2_fill_2 FILLER_18_874 ();
 sg13g2_fill_2 FILLER_18_915 ();
 sg13g2_fill_1 FILLER_18_917 ();
 sg13g2_fill_2 FILLER_18_988 ();
 sg13g2_fill_1 FILLER_18_990 ();
 sg13g2_fill_2 FILLER_18_1017 ();
 sg13g2_fill_1 FILLER_18_1019 ();
 sg13g2_decap_4 FILLER_18_1069 ();
 sg13g2_fill_1 FILLER_18_1095 ();
 sg13g2_decap_8 FILLER_18_1149 ();
 sg13g2_decap_8 FILLER_18_1156 ();
 sg13g2_fill_2 FILLER_18_1163 ();
 sg13g2_decap_4 FILLER_18_1169 ();
 sg13g2_fill_2 FILLER_18_1186 ();
 sg13g2_fill_1 FILLER_18_1217 ();
 sg13g2_fill_2 FILLER_18_1253 ();
 sg13g2_decap_8 FILLER_18_1304 ();
 sg13g2_decap_8 FILLER_18_1311 ();
 sg13g2_decap_8 FILLER_18_1318 ();
 sg13g2_decap_8 FILLER_18_1325 ();
 sg13g2_decap_8 FILLER_18_1332 ();
 sg13g2_decap_8 FILLER_18_1339 ();
 sg13g2_decap_8 FILLER_18_1346 ();
 sg13g2_decap_8 FILLER_18_1353 ();
 sg13g2_decap_8 FILLER_18_1360 ();
 sg13g2_decap_8 FILLER_18_1367 ();
 sg13g2_decap_8 FILLER_18_1374 ();
 sg13g2_decap_8 FILLER_18_1381 ();
 sg13g2_decap_8 FILLER_18_1388 ();
 sg13g2_decap_8 FILLER_18_1395 ();
 sg13g2_decap_8 FILLER_18_1402 ();
 sg13g2_decap_8 FILLER_18_1409 ();
 sg13g2_decap_8 FILLER_18_1416 ();
 sg13g2_decap_8 FILLER_18_1423 ();
 sg13g2_decap_8 FILLER_18_1430 ();
 sg13g2_decap_8 FILLER_18_1437 ();
 sg13g2_decap_8 FILLER_18_1444 ();
 sg13g2_decap_8 FILLER_18_1451 ();
 sg13g2_decap_8 FILLER_18_1458 ();
 sg13g2_decap_8 FILLER_18_1465 ();
 sg13g2_decap_8 FILLER_18_1472 ();
 sg13g2_decap_8 FILLER_18_1479 ();
 sg13g2_decap_8 FILLER_18_1486 ();
 sg13g2_decap_8 FILLER_18_1493 ();
 sg13g2_decap_8 FILLER_18_1500 ();
 sg13g2_decap_8 FILLER_18_1507 ();
 sg13g2_decap_8 FILLER_18_1514 ();
 sg13g2_decap_8 FILLER_18_1521 ();
 sg13g2_decap_8 FILLER_18_1528 ();
 sg13g2_decap_8 FILLER_18_1535 ();
 sg13g2_decap_8 FILLER_18_1542 ();
 sg13g2_decap_8 FILLER_18_1549 ();
 sg13g2_decap_8 FILLER_18_1556 ();
 sg13g2_decap_8 FILLER_18_1563 ();
 sg13g2_decap_8 FILLER_18_1570 ();
 sg13g2_decap_8 FILLER_18_1577 ();
 sg13g2_decap_8 FILLER_18_1584 ();
 sg13g2_decap_8 FILLER_18_1591 ();
 sg13g2_decap_8 FILLER_18_1598 ();
 sg13g2_decap_8 FILLER_18_1605 ();
 sg13g2_decap_8 FILLER_18_1612 ();
 sg13g2_decap_8 FILLER_18_1619 ();
 sg13g2_decap_8 FILLER_18_1626 ();
 sg13g2_decap_8 FILLER_18_1633 ();
 sg13g2_decap_8 FILLER_18_1640 ();
 sg13g2_decap_8 FILLER_18_1647 ();
 sg13g2_decap_8 FILLER_18_1654 ();
 sg13g2_decap_8 FILLER_18_1661 ();
 sg13g2_decap_8 FILLER_18_1668 ();
 sg13g2_decap_8 FILLER_18_1675 ();
 sg13g2_decap_8 FILLER_18_1682 ();
 sg13g2_decap_8 FILLER_18_1689 ();
 sg13g2_decap_8 FILLER_18_1696 ();
 sg13g2_decap_8 FILLER_18_1703 ();
 sg13g2_decap_8 FILLER_18_1710 ();
 sg13g2_decap_8 FILLER_18_1717 ();
 sg13g2_decap_8 FILLER_18_1724 ();
 sg13g2_decap_8 FILLER_18_1731 ();
 sg13g2_decap_8 FILLER_18_1738 ();
 sg13g2_decap_8 FILLER_18_1745 ();
 sg13g2_decap_8 FILLER_18_1752 ();
 sg13g2_decap_8 FILLER_18_1759 ();
 sg13g2_fill_2 FILLER_18_1766 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_fill_2 FILLER_19_35 ();
 sg13g2_fill_1 FILLER_19_63 ();
 sg13g2_fill_2 FILLER_19_79 ();
 sg13g2_fill_2 FILLER_19_138 ();
 sg13g2_fill_1 FILLER_19_145 ();
 sg13g2_fill_2 FILLER_19_196 ();
 sg13g2_fill_1 FILLER_19_198 ();
 sg13g2_fill_2 FILLER_19_212 ();
 sg13g2_fill_1 FILLER_19_214 ();
 sg13g2_fill_2 FILLER_19_223 ();
 sg13g2_fill_2 FILLER_19_286 ();
 sg13g2_decap_4 FILLER_19_330 ();
 sg13g2_decap_8 FILLER_19_380 ();
 sg13g2_decap_8 FILLER_19_387 ();
 sg13g2_fill_2 FILLER_19_394 ();
 sg13g2_fill_1 FILLER_19_396 ();
 sg13g2_decap_8 FILLER_19_405 ();
 sg13g2_decap_4 FILLER_19_412 ();
 sg13g2_fill_2 FILLER_19_416 ();
 sg13g2_fill_2 FILLER_19_435 ();
 sg13g2_fill_1 FILLER_19_457 ();
 sg13g2_fill_1 FILLER_19_468 ();
 sg13g2_fill_2 FILLER_19_485 ();
 sg13g2_fill_1 FILLER_19_487 ();
 sg13g2_fill_1 FILLER_19_497 ();
 sg13g2_fill_2 FILLER_19_529 ();
 sg13g2_fill_1 FILLER_19_565 ();
 sg13g2_fill_2 FILLER_19_571 ();
 sg13g2_fill_2 FILLER_19_599 ();
 sg13g2_fill_2 FILLER_19_609 ();
 sg13g2_fill_1 FILLER_19_611 ();
 sg13g2_fill_1 FILLER_19_657 ();
 sg13g2_fill_2 FILLER_19_756 ();
 sg13g2_fill_2 FILLER_19_784 ();
 sg13g2_fill_1 FILLER_19_786 ();
 sg13g2_fill_2 FILLER_19_824 ();
 sg13g2_fill_2 FILLER_19_831 ();
 sg13g2_fill_1 FILLER_19_833 ();
 sg13g2_fill_1 FILLER_19_840 ();
 sg13g2_decap_8 FILLER_19_856 ();
 sg13g2_fill_2 FILLER_19_889 ();
 sg13g2_decap_8 FILLER_19_925 ();
 sg13g2_fill_2 FILLER_19_932 ();
 sg13g2_fill_2 FILLER_19_939 ();
 sg13g2_fill_1 FILLER_19_941 ();
 sg13g2_fill_2 FILLER_19_970 ();
 sg13g2_fill_2 FILLER_19_996 ();
 sg13g2_fill_2 FILLER_19_1015 ();
 sg13g2_fill_1 FILLER_19_1017 ();
 sg13g2_decap_8 FILLER_19_1034 ();
 sg13g2_decap_8 FILLER_19_1041 ();
 sg13g2_fill_2 FILLER_19_1048 ();
 sg13g2_decap_4 FILLER_19_1074 ();
 sg13g2_fill_2 FILLER_19_1078 ();
 sg13g2_decap_4 FILLER_19_1130 ();
 sg13g2_decap_8 FILLER_19_1140 ();
 sg13g2_fill_1 FILLER_19_1147 ();
 sg13g2_fill_2 FILLER_19_1174 ();
 sg13g2_fill_2 FILLER_19_1207 ();
 sg13g2_fill_1 FILLER_19_1209 ();
 sg13g2_decap_8 FILLER_19_1306 ();
 sg13g2_decap_8 FILLER_19_1313 ();
 sg13g2_decap_8 FILLER_19_1320 ();
 sg13g2_decap_8 FILLER_19_1327 ();
 sg13g2_decap_8 FILLER_19_1334 ();
 sg13g2_decap_8 FILLER_19_1341 ();
 sg13g2_decap_8 FILLER_19_1348 ();
 sg13g2_decap_8 FILLER_19_1355 ();
 sg13g2_decap_8 FILLER_19_1362 ();
 sg13g2_decap_8 FILLER_19_1369 ();
 sg13g2_decap_8 FILLER_19_1376 ();
 sg13g2_decap_8 FILLER_19_1383 ();
 sg13g2_decap_8 FILLER_19_1390 ();
 sg13g2_decap_8 FILLER_19_1397 ();
 sg13g2_decap_8 FILLER_19_1404 ();
 sg13g2_decap_8 FILLER_19_1411 ();
 sg13g2_decap_8 FILLER_19_1418 ();
 sg13g2_decap_8 FILLER_19_1425 ();
 sg13g2_decap_8 FILLER_19_1432 ();
 sg13g2_decap_8 FILLER_19_1439 ();
 sg13g2_decap_8 FILLER_19_1446 ();
 sg13g2_decap_8 FILLER_19_1453 ();
 sg13g2_decap_8 FILLER_19_1460 ();
 sg13g2_decap_8 FILLER_19_1467 ();
 sg13g2_decap_8 FILLER_19_1474 ();
 sg13g2_decap_8 FILLER_19_1481 ();
 sg13g2_decap_8 FILLER_19_1488 ();
 sg13g2_decap_8 FILLER_19_1495 ();
 sg13g2_decap_8 FILLER_19_1502 ();
 sg13g2_decap_8 FILLER_19_1509 ();
 sg13g2_decap_8 FILLER_19_1516 ();
 sg13g2_decap_8 FILLER_19_1523 ();
 sg13g2_decap_8 FILLER_19_1530 ();
 sg13g2_decap_8 FILLER_19_1537 ();
 sg13g2_decap_8 FILLER_19_1544 ();
 sg13g2_decap_8 FILLER_19_1551 ();
 sg13g2_decap_8 FILLER_19_1558 ();
 sg13g2_decap_8 FILLER_19_1565 ();
 sg13g2_decap_8 FILLER_19_1572 ();
 sg13g2_decap_8 FILLER_19_1579 ();
 sg13g2_decap_8 FILLER_19_1586 ();
 sg13g2_decap_8 FILLER_19_1593 ();
 sg13g2_decap_8 FILLER_19_1600 ();
 sg13g2_decap_8 FILLER_19_1607 ();
 sg13g2_decap_8 FILLER_19_1614 ();
 sg13g2_decap_8 FILLER_19_1621 ();
 sg13g2_decap_8 FILLER_19_1628 ();
 sg13g2_decap_8 FILLER_19_1635 ();
 sg13g2_decap_8 FILLER_19_1642 ();
 sg13g2_decap_8 FILLER_19_1649 ();
 sg13g2_decap_8 FILLER_19_1656 ();
 sg13g2_decap_8 FILLER_19_1663 ();
 sg13g2_decap_8 FILLER_19_1670 ();
 sg13g2_decap_8 FILLER_19_1677 ();
 sg13g2_decap_8 FILLER_19_1684 ();
 sg13g2_decap_8 FILLER_19_1691 ();
 sg13g2_decap_8 FILLER_19_1698 ();
 sg13g2_decap_8 FILLER_19_1705 ();
 sg13g2_decap_8 FILLER_19_1712 ();
 sg13g2_decap_8 FILLER_19_1719 ();
 sg13g2_decap_8 FILLER_19_1726 ();
 sg13g2_decap_8 FILLER_19_1733 ();
 sg13g2_decap_8 FILLER_19_1740 ();
 sg13g2_decap_8 FILLER_19_1747 ();
 sg13g2_decap_8 FILLER_19_1754 ();
 sg13g2_decap_8 FILLER_19_1761 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_fill_1 FILLER_20_35 ();
 sg13g2_fill_2 FILLER_20_89 ();
 sg13g2_fill_1 FILLER_20_91 ();
 sg13g2_fill_2 FILLER_20_97 ();
 sg13g2_fill_1 FILLER_20_99 ();
 sg13g2_fill_2 FILLER_20_118 ();
 sg13g2_fill_1 FILLER_20_120 ();
 sg13g2_decap_4 FILLER_20_145 ();
 sg13g2_decap_8 FILLER_20_163 ();
 sg13g2_fill_1 FILLER_20_170 ();
 sg13g2_fill_1 FILLER_20_177 ();
 sg13g2_fill_1 FILLER_20_228 ();
 sg13g2_fill_1 FILLER_20_234 ();
 sg13g2_fill_1 FILLER_20_240 ();
 sg13g2_fill_1 FILLER_20_246 ();
 sg13g2_fill_1 FILLER_20_258 ();
 sg13g2_fill_1 FILLER_20_315 ();
 sg13g2_decap_4 FILLER_20_324 ();
 sg13g2_fill_2 FILLER_20_328 ();
 sg13g2_decap_4 FILLER_20_338 ();
 sg13g2_fill_1 FILLER_20_357 ();
 sg13g2_fill_2 FILLER_20_376 ();
 sg13g2_decap_4 FILLER_20_407 ();
 sg13g2_fill_1 FILLER_20_411 ();
 sg13g2_fill_2 FILLER_20_425 ();
 sg13g2_decap_4 FILLER_20_445 ();
 sg13g2_fill_2 FILLER_20_449 ();
 sg13g2_fill_2 FILLER_20_479 ();
 sg13g2_fill_2 FILLER_20_528 ();
 sg13g2_fill_2 FILLER_20_575 ();
 sg13g2_fill_1 FILLER_20_586 ();
 sg13g2_fill_2 FILLER_20_593 ();
 sg13g2_fill_2 FILLER_20_699 ();
 sg13g2_fill_1 FILLER_20_701 ();
 sg13g2_fill_2 FILLER_20_726 ();
 sg13g2_fill_1 FILLER_20_728 ();
 sg13g2_fill_1 FILLER_20_874 ();
 sg13g2_fill_2 FILLER_20_879 ();
 sg13g2_fill_1 FILLER_20_881 ();
 sg13g2_decap_4 FILLER_20_886 ();
 sg13g2_fill_2 FILLER_20_900 ();
 sg13g2_fill_2 FILLER_20_927 ();
 sg13g2_fill_1 FILLER_20_929 ();
 sg13g2_fill_2 FILLER_20_971 ();
 sg13g2_fill_1 FILLER_20_1009 ();
 sg13g2_decap_8 FILLER_20_1038 ();
 sg13g2_decap_8 FILLER_20_1045 ();
 sg13g2_decap_8 FILLER_20_1052 ();
 sg13g2_fill_1 FILLER_20_1059 ();
 sg13g2_decap_4 FILLER_20_1071 ();
 sg13g2_fill_1 FILLER_20_1097 ();
 sg13g2_fill_2 FILLER_20_1158 ();
 sg13g2_fill_1 FILLER_20_1160 ();
 sg13g2_fill_1 FILLER_20_1177 ();
 sg13g2_decap_8 FILLER_20_1210 ();
 sg13g2_fill_2 FILLER_20_1238 ();
 sg13g2_fill_2 FILLER_20_1249 ();
 sg13g2_fill_1 FILLER_20_1251 ();
 sg13g2_fill_2 FILLER_20_1274 ();
 sg13g2_fill_1 FILLER_20_1276 ();
 sg13g2_fill_2 FILLER_20_1282 ();
 sg13g2_fill_1 FILLER_20_1284 ();
 sg13g2_decap_8 FILLER_20_1315 ();
 sg13g2_decap_8 FILLER_20_1322 ();
 sg13g2_decap_8 FILLER_20_1329 ();
 sg13g2_decap_8 FILLER_20_1336 ();
 sg13g2_decap_8 FILLER_20_1343 ();
 sg13g2_decap_8 FILLER_20_1350 ();
 sg13g2_decap_8 FILLER_20_1357 ();
 sg13g2_decap_8 FILLER_20_1364 ();
 sg13g2_decap_8 FILLER_20_1371 ();
 sg13g2_decap_8 FILLER_20_1378 ();
 sg13g2_decap_8 FILLER_20_1385 ();
 sg13g2_decap_8 FILLER_20_1392 ();
 sg13g2_decap_8 FILLER_20_1399 ();
 sg13g2_decap_8 FILLER_20_1406 ();
 sg13g2_decap_8 FILLER_20_1413 ();
 sg13g2_decap_8 FILLER_20_1420 ();
 sg13g2_decap_8 FILLER_20_1427 ();
 sg13g2_decap_8 FILLER_20_1434 ();
 sg13g2_decap_8 FILLER_20_1441 ();
 sg13g2_decap_8 FILLER_20_1448 ();
 sg13g2_decap_8 FILLER_20_1455 ();
 sg13g2_decap_8 FILLER_20_1462 ();
 sg13g2_decap_8 FILLER_20_1469 ();
 sg13g2_decap_8 FILLER_20_1476 ();
 sg13g2_decap_8 FILLER_20_1483 ();
 sg13g2_decap_8 FILLER_20_1490 ();
 sg13g2_decap_8 FILLER_20_1497 ();
 sg13g2_decap_8 FILLER_20_1504 ();
 sg13g2_decap_8 FILLER_20_1511 ();
 sg13g2_decap_8 FILLER_20_1518 ();
 sg13g2_decap_8 FILLER_20_1525 ();
 sg13g2_decap_8 FILLER_20_1532 ();
 sg13g2_decap_8 FILLER_20_1539 ();
 sg13g2_decap_8 FILLER_20_1546 ();
 sg13g2_decap_8 FILLER_20_1553 ();
 sg13g2_decap_8 FILLER_20_1560 ();
 sg13g2_decap_8 FILLER_20_1567 ();
 sg13g2_decap_8 FILLER_20_1574 ();
 sg13g2_decap_8 FILLER_20_1581 ();
 sg13g2_decap_8 FILLER_20_1588 ();
 sg13g2_decap_8 FILLER_20_1595 ();
 sg13g2_decap_8 FILLER_20_1602 ();
 sg13g2_decap_8 FILLER_20_1609 ();
 sg13g2_decap_8 FILLER_20_1616 ();
 sg13g2_decap_8 FILLER_20_1623 ();
 sg13g2_decap_8 FILLER_20_1630 ();
 sg13g2_decap_8 FILLER_20_1637 ();
 sg13g2_decap_8 FILLER_20_1644 ();
 sg13g2_decap_8 FILLER_20_1651 ();
 sg13g2_decap_8 FILLER_20_1658 ();
 sg13g2_decap_8 FILLER_20_1665 ();
 sg13g2_decap_8 FILLER_20_1672 ();
 sg13g2_decap_8 FILLER_20_1679 ();
 sg13g2_decap_8 FILLER_20_1686 ();
 sg13g2_decap_8 FILLER_20_1693 ();
 sg13g2_decap_8 FILLER_20_1700 ();
 sg13g2_decap_8 FILLER_20_1707 ();
 sg13g2_decap_8 FILLER_20_1714 ();
 sg13g2_decap_8 FILLER_20_1721 ();
 sg13g2_decap_8 FILLER_20_1728 ();
 sg13g2_decap_8 FILLER_20_1735 ();
 sg13g2_decap_8 FILLER_20_1742 ();
 sg13g2_decap_8 FILLER_20_1749 ();
 sg13g2_decap_8 FILLER_20_1756 ();
 sg13g2_decap_4 FILLER_20_1763 ();
 sg13g2_fill_1 FILLER_20_1767 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_fill_2 FILLER_21_56 ();
 sg13g2_fill_1 FILLER_21_58 ();
 sg13g2_fill_2 FILLER_21_94 ();
 sg13g2_fill_1 FILLER_21_96 ();
 sg13g2_fill_1 FILLER_21_133 ();
 sg13g2_fill_1 FILLER_21_140 ();
 sg13g2_fill_2 FILLER_21_188 ();
 sg13g2_fill_1 FILLER_21_225 ();
 sg13g2_fill_2 FILLER_21_267 ();
 sg13g2_decap_8 FILLER_21_281 ();
 sg13g2_decap_4 FILLER_21_288 ();
 sg13g2_decap_8 FILLER_21_296 ();
 sg13g2_fill_1 FILLER_21_315 ();
 sg13g2_decap_4 FILLER_21_321 ();
 sg13g2_fill_2 FILLER_21_335 ();
 sg13g2_fill_1 FILLER_21_337 ();
 sg13g2_fill_2 FILLER_21_344 ();
 sg13g2_fill_1 FILLER_21_352 ();
 sg13g2_decap_4 FILLER_21_385 ();
 sg13g2_fill_2 FILLER_21_407 ();
 sg13g2_fill_1 FILLER_21_409 ();
 sg13g2_decap_4 FILLER_21_438 ();
 sg13g2_fill_1 FILLER_21_442 ();
 sg13g2_fill_1 FILLER_21_467 ();
 sg13g2_fill_1 FILLER_21_473 ();
 sg13g2_fill_2 FILLER_21_488 ();
 sg13g2_fill_1 FILLER_21_490 ();
 sg13g2_fill_1 FILLER_21_574 ();
 sg13g2_fill_2 FILLER_21_618 ();
 sg13g2_fill_1 FILLER_21_620 ();
 sg13g2_fill_2 FILLER_21_656 ();
 sg13g2_fill_1 FILLER_21_673 ();
 sg13g2_fill_2 FILLER_21_712 ();
 sg13g2_fill_1 FILLER_21_714 ();
 sg13g2_fill_1 FILLER_21_756 ();
 sg13g2_fill_2 FILLER_21_778 ();
 sg13g2_fill_1 FILLER_21_780 ();
 sg13g2_fill_2 FILLER_21_816 ();
 sg13g2_fill_2 FILLER_21_844 ();
 sg13g2_fill_1 FILLER_21_846 ();
 sg13g2_fill_2 FILLER_21_879 ();
 sg13g2_fill_1 FILLER_21_881 ();
 sg13g2_fill_2 FILLER_21_896 ();
 sg13g2_fill_1 FILLER_21_898 ();
 sg13g2_fill_1 FILLER_21_922 ();
 sg13g2_decap_8 FILLER_21_932 ();
 sg13g2_fill_1 FILLER_21_939 ();
 sg13g2_fill_1 FILLER_21_944 ();
 sg13g2_decap_8 FILLER_21_971 ();
 sg13g2_decap_8 FILLER_21_978 ();
 sg13g2_fill_2 FILLER_21_985 ();
 sg13g2_fill_1 FILLER_21_987 ();
 sg13g2_fill_2 FILLER_21_997 ();
 sg13g2_fill_1 FILLER_21_999 ();
 sg13g2_fill_2 FILLER_21_1016 ();
 sg13g2_fill_1 FILLER_21_1018 ();
 sg13g2_fill_2 FILLER_21_1099 ();
 sg13g2_fill_1 FILLER_21_1101 ();
 sg13g2_fill_2 FILLER_21_1111 ();
 sg13g2_fill_2 FILLER_21_1117 ();
 sg13g2_decap_8 FILLER_21_1128 ();
 sg13g2_fill_2 FILLER_21_1174 ();
 sg13g2_fill_2 FILLER_21_1202 ();
 sg13g2_fill_2 FILLER_21_1245 ();
 sg13g2_fill_1 FILLER_21_1252 ();
 sg13g2_fill_2 FILLER_21_1283 ();
 sg13g2_decap_8 FILLER_21_1320 ();
 sg13g2_decap_8 FILLER_21_1327 ();
 sg13g2_decap_8 FILLER_21_1334 ();
 sg13g2_decap_8 FILLER_21_1341 ();
 sg13g2_decap_8 FILLER_21_1348 ();
 sg13g2_decap_8 FILLER_21_1355 ();
 sg13g2_decap_8 FILLER_21_1362 ();
 sg13g2_decap_8 FILLER_21_1369 ();
 sg13g2_decap_8 FILLER_21_1376 ();
 sg13g2_decap_8 FILLER_21_1383 ();
 sg13g2_decap_8 FILLER_21_1390 ();
 sg13g2_decap_8 FILLER_21_1397 ();
 sg13g2_decap_8 FILLER_21_1404 ();
 sg13g2_decap_8 FILLER_21_1411 ();
 sg13g2_decap_8 FILLER_21_1418 ();
 sg13g2_decap_8 FILLER_21_1425 ();
 sg13g2_decap_8 FILLER_21_1432 ();
 sg13g2_decap_8 FILLER_21_1439 ();
 sg13g2_decap_8 FILLER_21_1446 ();
 sg13g2_decap_8 FILLER_21_1453 ();
 sg13g2_decap_8 FILLER_21_1460 ();
 sg13g2_decap_8 FILLER_21_1467 ();
 sg13g2_decap_8 FILLER_21_1474 ();
 sg13g2_decap_8 FILLER_21_1481 ();
 sg13g2_decap_8 FILLER_21_1488 ();
 sg13g2_decap_8 FILLER_21_1495 ();
 sg13g2_decap_8 FILLER_21_1502 ();
 sg13g2_decap_8 FILLER_21_1509 ();
 sg13g2_decap_8 FILLER_21_1516 ();
 sg13g2_decap_8 FILLER_21_1523 ();
 sg13g2_decap_8 FILLER_21_1530 ();
 sg13g2_decap_8 FILLER_21_1537 ();
 sg13g2_decap_8 FILLER_21_1544 ();
 sg13g2_decap_8 FILLER_21_1551 ();
 sg13g2_decap_8 FILLER_21_1558 ();
 sg13g2_decap_8 FILLER_21_1565 ();
 sg13g2_decap_8 FILLER_21_1572 ();
 sg13g2_decap_8 FILLER_21_1579 ();
 sg13g2_decap_8 FILLER_21_1586 ();
 sg13g2_decap_8 FILLER_21_1593 ();
 sg13g2_decap_8 FILLER_21_1600 ();
 sg13g2_decap_8 FILLER_21_1607 ();
 sg13g2_decap_8 FILLER_21_1614 ();
 sg13g2_decap_8 FILLER_21_1621 ();
 sg13g2_decap_8 FILLER_21_1628 ();
 sg13g2_decap_8 FILLER_21_1635 ();
 sg13g2_decap_8 FILLER_21_1642 ();
 sg13g2_decap_8 FILLER_21_1649 ();
 sg13g2_decap_8 FILLER_21_1656 ();
 sg13g2_decap_8 FILLER_21_1663 ();
 sg13g2_decap_8 FILLER_21_1670 ();
 sg13g2_decap_8 FILLER_21_1677 ();
 sg13g2_decap_8 FILLER_21_1684 ();
 sg13g2_decap_8 FILLER_21_1691 ();
 sg13g2_decap_8 FILLER_21_1698 ();
 sg13g2_decap_8 FILLER_21_1705 ();
 sg13g2_decap_8 FILLER_21_1712 ();
 sg13g2_decap_8 FILLER_21_1719 ();
 sg13g2_decap_8 FILLER_21_1726 ();
 sg13g2_decap_8 FILLER_21_1733 ();
 sg13g2_decap_8 FILLER_21_1740 ();
 sg13g2_decap_8 FILLER_21_1747 ();
 sg13g2_decap_8 FILLER_21_1754 ();
 sg13g2_decap_8 FILLER_21_1761 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_4 FILLER_22_35 ();
 sg13g2_fill_2 FILLER_22_39 ();
 sg13g2_decap_4 FILLER_22_101 ();
 sg13g2_fill_2 FILLER_22_105 ();
 sg13g2_decap_4 FILLER_22_112 ();
 sg13g2_fill_2 FILLER_22_116 ();
 sg13g2_decap_4 FILLER_22_122 ();
 sg13g2_fill_2 FILLER_22_166 ();
 sg13g2_fill_1 FILLER_22_174 ();
 sg13g2_fill_2 FILLER_22_180 ();
 sg13g2_fill_1 FILLER_22_187 ();
 sg13g2_fill_2 FILLER_22_193 ();
 sg13g2_fill_1 FILLER_22_195 ();
 sg13g2_decap_4 FILLER_22_259 ();
 sg13g2_fill_2 FILLER_22_263 ();
 sg13g2_decap_4 FILLER_22_275 ();
 sg13g2_fill_2 FILLER_22_331 ();
 sg13g2_fill_2 FILLER_22_394 ();
 sg13g2_fill_1 FILLER_22_396 ();
 sg13g2_fill_2 FILLER_22_405 ();
 sg13g2_fill_1 FILLER_22_420 ();
 sg13g2_decap_4 FILLER_22_428 ();
 sg13g2_fill_1 FILLER_22_432 ();
 sg13g2_fill_2 FILLER_22_485 ();
 sg13g2_fill_1 FILLER_22_487 ();
 sg13g2_fill_1 FILLER_22_519 ();
 sg13g2_fill_2 FILLER_22_529 ();
 sg13g2_fill_2 FILLER_22_541 ();
 sg13g2_fill_1 FILLER_22_543 ();
 sg13g2_fill_2 FILLER_22_608 ();
 sg13g2_fill_1 FILLER_22_610 ();
 sg13g2_fill_2 FILLER_22_661 ();
 sg13g2_fill_2 FILLER_22_689 ();
 sg13g2_decap_8 FILLER_22_780 ();
 sg13g2_fill_1 FILLER_22_787 ();
 sg13g2_fill_2 FILLER_22_832 ();
 sg13g2_fill_1 FILLER_22_834 ();
 sg13g2_fill_2 FILLER_22_922 ();
 sg13g2_fill_1 FILLER_22_930 ();
 sg13g2_decap_8 FILLER_22_949 ();
 sg13g2_decap_8 FILLER_22_965 ();
 sg13g2_fill_1 FILLER_22_972 ();
 sg13g2_decap_8 FILLER_22_981 ();
 sg13g2_fill_1 FILLER_22_988 ();
 sg13g2_fill_2 FILLER_22_994 ();
 sg13g2_fill_2 FILLER_22_1001 ();
 sg13g2_fill_1 FILLER_22_1003 ();
 sg13g2_decap_8 FILLER_22_1009 ();
 sg13g2_decap_8 FILLER_22_1016 ();
 sg13g2_fill_2 FILLER_22_1042 ();
 sg13g2_fill_1 FILLER_22_1044 ();
 sg13g2_fill_2 FILLER_22_1071 ();
 sg13g2_fill_2 FILLER_22_1087 ();
 sg13g2_fill_1 FILLER_22_1089 ();
 sg13g2_decap_4 FILLER_22_1116 ();
 sg13g2_fill_2 FILLER_22_1120 ();
 sg13g2_fill_2 FILLER_22_1127 ();
 sg13g2_fill_1 FILLER_22_1129 ();
 sg13g2_fill_1 FILLER_22_1156 ();
 sg13g2_fill_2 FILLER_22_1185 ();
 sg13g2_fill_1 FILLER_22_1187 ();
 sg13g2_fill_2 FILLER_22_1211 ();
 sg13g2_fill_1 FILLER_22_1213 ();
 sg13g2_fill_2 FILLER_22_1218 ();
 sg13g2_fill_1 FILLER_22_1234 ();
 sg13g2_fill_2 FILLER_22_1269 ();
 sg13g2_fill_2 FILLER_22_1292 ();
 sg13g2_decap_8 FILLER_22_1333 ();
 sg13g2_decap_8 FILLER_22_1340 ();
 sg13g2_decap_8 FILLER_22_1347 ();
 sg13g2_decap_8 FILLER_22_1354 ();
 sg13g2_decap_8 FILLER_22_1361 ();
 sg13g2_decap_8 FILLER_22_1368 ();
 sg13g2_decap_8 FILLER_22_1375 ();
 sg13g2_decap_8 FILLER_22_1382 ();
 sg13g2_decap_8 FILLER_22_1389 ();
 sg13g2_decap_8 FILLER_22_1396 ();
 sg13g2_decap_8 FILLER_22_1403 ();
 sg13g2_decap_8 FILLER_22_1410 ();
 sg13g2_decap_8 FILLER_22_1417 ();
 sg13g2_decap_8 FILLER_22_1424 ();
 sg13g2_decap_8 FILLER_22_1431 ();
 sg13g2_decap_8 FILLER_22_1438 ();
 sg13g2_decap_8 FILLER_22_1445 ();
 sg13g2_decap_8 FILLER_22_1452 ();
 sg13g2_decap_8 FILLER_22_1459 ();
 sg13g2_decap_8 FILLER_22_1466 ();
 sg13g2_decap_8 FILLER_22_1473 ();
 sg13g2_decap_8 FILLER_22_1480 ();
 sg13g2_decap_8 FILLER_22_1487 ();
 sg13g2_decap_8 FILLER_22_1494 ();
 sg13g2_decap_8 FILLER_22_1501 ();
 sg13g2_decap_8 FILLER_22_1508 ();
 sg13g2_decap_8 FILLER_22_1515 ();
 sg13g2_decap_8 FILLER_22_1522 ();
 sg13g2_decap_8 FILLER_22_1529 ();
 sg13g2_decap_8 FILLER_22_1536 ();
 sg13g2_decap_8 FILLER_22_1543 ();
 sg13g2_decap_8 FILLER_22_1550 ();
 sg13g2_decap_8 FILLER_22_1557 ();
 sg13g2_decap_8 FILLER_22_1564 ();
 sg13g2_decap_8 FILLER_22_1571 ();
 sg13g2_decap_8 FILLER_22_1578 ();
 sg13g2_decap_8 FILLER_22_1585 ();
 sg13g2_decap_8 FILLER_22_1592 ();
 sg13g2_decap_8 FILLER_22_1599 ();
 sg13g2_decap_8 FILLER_22_1606 ();
 sg13g2_decap_8 FILLER_22_1613 ();
 sg13g2_decap_8 FILLER_22_1620 ();
 sg13g2_decap_8 FILLER_22_1627 ();
 sg13g2_decap_8 FILLER_22_1634 ();
 sg13g2_decap_8 FILLER_22_1641 ();
 sg13g2_decap_8 FILLER_22_1648 ();
 sg13g2_decap_8 FILLER_22_1655 ();
 sg13g2_decap_8 FILLER_22_1662 ();
 sg13g2_decap_8 FILLER_22_1669 ();
 sg13g2_decap_8 FILLER_22_1676 ();
 sg13g2_decap_8 FILLER_22_1683 ();
 sg13g2_decap_8 FILLER_22_1690 ();
 sg13g2_decap_8 FILLER_22_1697 ();
 sg13g2_decap_8 FILLER_22_1704 ();
 sg13g2_decap_8 FILLER_22_1711 ();
 sg13g2_decap_8 FILLER_22_1718 ();
 sg13g2_decap_8 FILLER_22_1725 ();
 sg13g2_decap_8 FILLER_22_1732 ();
 sg13g2_decap_8 FILLER_22_1739 ();
 sg13g2_decap_8 FILLER_22_1746 ();
 sg13g2_decap_8 FILLER_22_1753 ();
 sg13g2_decap_8 FILLER_22_1760 ();
 sg13g2_fill_1 FILLER_22_1767 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_fill_2 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_85 ();
 sg13g2_decap_8 FILLER_23_92 ();
 sg13g2_fill_2 FILLER_23_99 ();
 sg13g2_fill_1 FILLER_23_107 ();
 sg13g2_fill_2 FILLER_23_123 ();
 sg13g2_decap_8 FILLER_23_129 ();
 sg13g2_fill_2 FILLER_23_136 ();
 sg13g2_fill_1 FILLER_23_138 ();
 sg13g2_fill_2 FILLER_23_180 ();
 sg13g2_decap_4 FILLER_23_213 ();
 sg13g2_fill_2 FILLER_23_223 ();
 sg13g2_decap_4 FILLER_23_235 ();
 sg13g2_fill_2 FILLER_23_239 ();
 sg13g2_fill_2 FILLER_23_276 ();
 sg13g2_fill_1 FILLER_23_340 ();
 sg13g2_fill_2 FILLER_23_346 ();
 sg13g2_fill_2 FILLER_23_357 ();
 sg13g2_fill_2 FILLER_23_368 ();
 sg13g2_fill_1 FILLER_23_375 ();
 sg13g2_fill_2 FILLER_23_390 ();
 sg13g2_fill_1 FILLER_23_397 ();
 sg13g2_decap_8 FILLER_23_407 ();
 sg13g2_fill_2 FILLER_23_423 ();
 sg13g2_fill_1 FILLER_23_425 ();
 sg13g2_decap_8 FILLER_23_434 ();
 sg13g2_fill_1 FILLER_23_441 ();
 sg13g2_fill_2 FILLER_23_530 ();
 sg13g2_fill_1 FILLER_23_567 ();
 sg13g2_fill_2 FILLER_23_627 ();
 sg13g2_fill_1 FILLER_23_629 ();
 sg13g2_fill_1 FILLER_23_691 ();
 sg13g2_fill_2 FILLER_23_703 ();
 sg13g2_fill_1 FILLER_23_705 ();
 sg13g2_fill_2 FILLER_23_730 ();
 sg13g2_fill_1 FILLER_23_732 ();
 sg13g2_decap_8 FILLER_23_786 ();
 sg13g2_fill_1 FILLER_23_793 ();
 sg13g2_decap_8 FILLER_23_799 ();
 sg13g2_decap_8 FILLER_23_806 ();
 sg13g2_decap_8 FILLER_23_813 ();
 sg13g2_fill_2 FILLER_23_820 ();
 sg13g2_fill_1 FILLER_23_822 ();
 sg13g2_fill_2 FILLER_23_842 ();
 sg13g2_fill_2 FILLER_23_853 ();
 sg13g2_fill_1 FILLER_23_855 ();
 sg13g2_decap_4 FILLER_23_864 ();
 sg13g2_fill_2 FILLER_23_883 ();
 sg13g2_fill_1 FILLER_23_885 ();
 sg13g2_fill_2 FILLER_23_891 ();
 sg13g2_fill_2 FILLER_23_919 ();
 sg13g2_fill_1 FILLER_23_921 ();
 sg13g2_fill_1 FILLER_23_936 ();
 sg13g2_decap_8 FILLER_23_997 ();
 sg13g2_fill_2 FILLER_23_1051 ();
 sg13g2_fill_1 FILLER_23_1053 ();
 sg13g2_fill_2 FILLER_23_1058 ();
 sg13g2_fill_2 FILLER_23_1115 ();
 sg13g2_fill_1 FILLER_23_1117 ();
 sg13g2_fill_1 FILLER_23_1152 ();
 sg13g2_decap_8 FILLER_23_1187 ();
 sg13g2_fill_1 FILLER_23_1199 ();
 sg13g2_fill_1 FILLER_23_1248 ();
 sg13g2_fill_1 FILLER_23_1264 ();
 sg13g2_fill_1 FILLER_23_1284 ();
 sg13g2_decap_8 FILLER_23_1338 ();
 sg13g2_decap_8 FILLER_23_1345 ();
 sg13g2_decap_8 FILLER_23_1352 ();
 sg13g2_decap_8 FILLER_23_1359 ();
 sg13g2_decap_8 FILLER_23_1366 ();
 sg13g2_decap_8 FILLER_23_1373 ();
 sg13g2_decap_8 FILLER_23_1380 ();
 sg13g2_decap_8 FILLER_23_1387 ();
 sg13g2_decap_8 FILLER_23_1394 ();
 sg13g2_decap_8 FILLER_23_1401 ();
 sg13g2_decap_8 FILLER_23_1408 ();
 sg13g2_decap_8 FILLER_23_1415 ();
 sg13g2_decap_8 FILLER_23_1422 ();
 sg13g2_decap_8 FILLER_23_1429 ();
 sg13g2_decap_8 FILLER_23_1436 ();
 sg13g2_decap_8 FILLER_23_1443 ();
 sg13g2_decap_8 FILLER_23_1450 ();
 sg13g2_decap_8 FILLER_23_1457 ();
 sg13g2_decap_8 FILLER_23_1464 ();
 sg13g2_decap_8 FILLER_23_1471 ();
 sg13g2_decap_8 FILLER_23_1478 ();
 sg13g2_decap_8 FILLER_23_1485 ();
 sg13g2_decap_8 FILLER_23_1492 ();
 sg13g2_decap_8 FILLER_23_1499 ();
 sg13g2_decap_8 FILLER_23_1506 ();
 sg13g2_decap_8 FILLER_23_1513 ();
 sg13g2_decap_8 FILLER_23_1520 ();
 sg13g2_decap_8 FILLER_23_1527 ();
 sg13g2_decap_8 FILLER_23_1534 ();
 sg13g2_decap_8 FILLER_23_1541 ();
 sg13g2_decap_8 FILLER_23_1548 ();
 sg13g2_decap_8 FILLER_23_1555 ();
 sg13g2_decap_8 FILLER_23_1562 ();
 sg13g2_decap_8 FILLER_23_1569 ();
 sg13g2_decap_8 FILLER_23_1576 ();
 sg13g2_decap_8 FILLER_23_1583 ();
 sg13g2_decap_8 FILLER_23_1590 ();
 sg13g2_decap_8 FILLER_23_1597 ();
 sg13g2_decap_8 FILLER_23_1604 ();
 sg13g2_decap_8 FILLER_23_1611 ();
 sg13g2_decap_8 FILLER_23_1618 ();
 sg13g2_decap_8 FILLER_23_1625 ();
 sg13g2_decap_8 FILLER_23_1632 ();
 sg13g2_decap_8 FILLER_23_1639 ();
 sg13g2_decap_8 FILLER_23_1646 ();
 sg13g2_decap_8 FILLER_23_1653 ();
 sg13g2_decap_8 FILLER_23_1660 ();
 sg13g2_decap_8 FILLER_23_1667 ();
 sg13g2_decap_8 FILLER_23_1674 ();
 sg13g2_decap_8 FILLER_23_1681 ();
 sg13g2_decap_8 FILLER_23_1688 ();
 sg13g2_decap_8 FILLER_23_1695 ();
 sg13g2_decap_8 FILLER_23_1702 ();
 sg13g2_decap_8 FILLER_23_1709 ();
 sg13g2_decap_8 FILLER_23_1716 ();
 sg13g2_decap_8 FILLER_23_1723 ();
 sg13g2_decap_8 FILLER_23_1730 ();
 sg13g2_decap_8 FILLER_23_1737 ();
 sg13g2_decap_8 FILLER_23_1744 ();
 sg13g2_decap_8 FILLER_23_1751 ();
 sg13g2_decap_8 FILLER_23_1758 ();
 sg13g2_fill_2 FILLER_23_1765 ();
 sg13g2_fill_1 FILLER_23_1767 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_fill_2 FILLER_24_49 ();
 sg13g2_fill_2 FILLER_24_73 ();
 sg13g2_fill_1 FILLER_24_75 ();
 sg13g2_fill_2 FILLER_24_147 ();
 sg13g2_fill_1 FILLER_24_149 ();
 sg13g2_fill_2 FILLER_24_156 ();
 sg13g2_fill_1 FILLER_24_184 ();
 sg13g2_decap_8 FILLER_24_204 ();
 sg13g2_fill_1 FILLER_24_216 ();
 sg13g2_fill_1 FILLER_24_228 ();
 sg13g2_fill_2 FILLER_24_243 ();
 sg13g2_fill_2 FILLER_24_260 ();
 sg13g2_fill_2 FILLER_24_317 ();
 sg13g2_fill_1 FILLER_24_319 ();
 sg13g2_fill_2 FILLER_24_394 ();
 sg13g2_fill_1 FILLER_24_396 ();
 sg13g2_fill_1 FILLER_24_423 ();
 sg13g2_fill_2 FILLER_24_442 ();
 sg13g2_fill_1 FILLER_24_444 ();
 sg13g2_decap_4 FILLER_24_454 ();
 sg13g2_decap_8 FILLER_24_501 ();
 sg13g2_fill_1 FILLER_24_508 ();
 sg13g2_fill_2 FILLER_24_525 ();
 sg13g2_fill_1 FILLER_24_527 ();
 sg13g2_fill_2 FILLER_24_559 ();
 sg13g2_fill_2 FILLER_24_587 ();
 sg13g2_fill_2 FILLER_24_603 ();
 sg13g2_fill_1 FILLER_24_605 ();
 sg13g2_decap_8 FILLER_24_640 ();
 sg13g2_decap_4 FILLER_24_679 ();
 sg13g2_fill_1 FILLER_24_726 ();
 sg13g2_fill_1 FILLER_24_744 ();
 sg13g2_fill_2 FILLER_24_774 ();
 sg13g2_decap_8 FILLER_24_792 ();
 sg13g2_fill_1 FILLER_24_799 ();
 sg13g2_fill_2 FILLER_24_826 ();
 sg13g2_fill_2 FILLER_24_871 ();
 sg13g2_fill_2 FILLER_24_964 ();
 sg13g2_fill_1 FILLER_24_966 ();
 sg13g2_fill_1 FILLER_24_994 ();
 sg13g2_decap_8 FILLER_24_1013 ();
 sg13g2_decap_4 FILLER_24_1020 ();
 sg13g2_fill_1 FILLER_24_1024 ();
 sg13g2_fill_2 FILLER_24_1042 ();
 sg13g2_fill_1 FILLER_24_1044 ();
 sg13g2_fill_2 FILLER_24_1120 ();
 sg13g2_fill_2 FILLER_24_1126 ();
 sg13g2_fill_2 FILLER_24_1133 ();
 sg13g2_fill_2 FILLER_24_1153 ();
 sg13g2_fill_1 FILLER_24_1155 ();
 sg13g2_fill_2 FILLER_24_1201 ();
 sg13g2_fill_1 FILLER_24_1203 ();
 sg13g2_fill_2 FILLER_24_1212 ();
 sg13g2_fill_2 FILLER_24_1218 ();
 sg13g2_fill_1 FILLER_24_1220 ();
 sg13g2_fill_1 FILLER_24_1255 ();
 sg13g2_decap_8 FILLER_24_1340 ();
 sg13g2_decap_8 FILLER_24_1347 ();
 sg13g2_decap_8 FILLER_24_1354 ();
 sg13g2_decap_8 FILLER_24_1361 ();
 sg13g2_decap_8 FILLER_24_1368 ();
 sg13g2_decap_8 FILLER_24_1375 ();
 sg13g2_decap_8 FILLER_24_1382 ();
 sg13g2_decap_8 FILLER_24_1389 ();
 sg13g2_decap_8 FILLER_24_1396 ();
 sg13g2_decap_8 FILLER_24_1403 ();
 sg13g2_decap_8 FILLER_24_1410 ();
 sg13g2_decap_8 FILLER_24_1417 ();
 sg13g2_decap_8 FILLER_24_1424 ();
 sg13g2_decap_8 FILLER_24_1431 ();
 sg13g2_decap_8 FILLER_24_1438 ();
 sg13g2_decap_8 FILLER_24_1445 ();
 sg13g2_decap_8 FILLER_24_1452 ();
 sg13g2_decap_8 FILLER_24_1459 ();
 sg13g2_decap_8 FILLER_24_1466 ();
 sg13g2_decap_8 FILLER_24_1473 ();
 sg13g2_decap_8 FILLER_24_1480 ();
 sg13g2_decap_8 FILLER_24_1487 ();
 sg13g2_decap_8 FILLER_24_1494 ();
 sg13g2_decap_8 FILLER_24_1501 ();
 sg13g2_decap_8 FILLER_24_1508 ();
 sg13g2_decap_8 FILLER_24_1515 ();
 sg13g2_decap_8 FILLER_24_1522 ();
 sg13g2_decap_8 FILLER_24_1529 ();
 sg13g2_decap_8 FILLER_24_1536 ();
 sg13g2_decap_8 FILLER_24_1543 ();
 sg13g2_decap_8 FILLER_24_1550 ();
 sg13g2_decap_8 FILLER_24_1557 ();
 sg13g2_decap_8 FILLER_24_1564 ();
 sg13g2_decap_8 FILLER_24_1571 ();
 sg13g2_decap_8 FILLER_24_1578 ();
 sg13g2_decap_8 FILLER_24_1585 ();
 sg13g2_decap_8 FILLER_24_1592 ();
 sg13g2_decap_8 FILLER_24_1599 ();
 sg13g2_decap_8 FILLER_24_1606 ();
 sg13g2_decap_8 FILLER_24_1613 ();
 sg13g2_decap_8 FILLER_24_1620 ();
 sg13g2_decap_8 FILLER_24_1627 ();
 sg13g2_decap_8 FILLER_24_1634 ();
 sg13g2_decap_8 FILLER_24_1641 ();
 sg13g2_decap_8 FILLER_24_1648 ();
 sg13g2_decap_8 FILLER_24_1655 ();
 sg13g2_decap_8 FILLER_24_1662 ();
 sg13g2_decap_8 FILLER_24_1669 ();
 sg13g2_decap_8 FILLER_24_1676 ();
 sg13g2_decap_8 FILLER_24_1683 ();
 sg13g2_decap_8 FILLER_24_1690 ();
 sg13g2_decap_8 FILLER_24_1697 ();
 sg13g2_decap_8 FILLER_24_1704 ();
 sg13g2_decap_8 FILLER_24_1711 ();
 sg13g2_decap_8 FILLER_24_1718 ();
 sg13g2_decap_8 FILLER_24_1725 ();
 sg13g2_decap_8 FILLER_24_1732 ();
 sg13g2_decap_8 FILLER_24_1739 ();
 sg13g2_decap_8 FILLER_24_1746 ();
 sg13g2_decap_8 FILLER_24_1753 ();
 sg13g2_decap_8 FILLER_24_1760 ();
 sg13g2_fill_1 FILLER_24_1767 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_fill_2 FILLER_25_42 ();
 sg13g2_fill_1 FILLER_25_44 ();
 sg13g2_decap_4 FILLER_25_93 ();
 sg13g2_fill_1 FILLER_25_108 ();
 sg13g2_fill_1 FILLER_25_114 ();
 sg13g2_decap_8 FILLER_25_126 ();
 sg13g2_fill_2 FILLER_25_133 ();
 sg13g2_decap_8 FILLER_25_140 ();
 sg13g2_decap_4 FILLER_25_147 ();
 sg13g2_fill_2 FILLER_25_160 ();
 sg13g2_fill_2 FILLER_25_167 ();
 sg13g2_fill_2 FILLER_25_218 ();
 sg13g2_fill_2 FILLER_25_223 ();
 sg13g2_fill_1 FILLER_25_225 ();
 sg13g2_fill_2 FILLER_25_255 ();
 sg13g2_fill_2 FILLER_25_357 ();
 sg13g2_fill_1 FILLER_25_359 ();
 sg13g2_fill_2 FILLER_25_375 ();
 sg13g2_fill_1 FILLER_25_387 ();
 sg13g2_fill_2 FILLER_25_433 ();
 sg13g2_fill_2 FILLER_25_458 ();
 sg13g2_decap_8 FILLER_25_475 ();
 sg13g2_fill_1 FILLER_25_482 ();
 sg13g2_decap_4 FILLER_25_487 ();
 sg13g2_fill_1 FILLER_25_491 ();
 sg13g2_fill_1 FILLER_25_505 ();
 sg13g2_decap_4 FILLER_25_510 ();
 sg13g2_decap_8 FILLER_25_517 ();
 sg13g2_decap_4 FILLER_25_524 ();
 sg13g2_fill_2 FILLER_25_564 ();
 sg13g2_fill_2 FILLER_25_571 ();
 sg13g2_fill_1 FILLER_25_573 ();
 sg13g2_decap_8 FILLER_25_582 ();
 sg13g2_decap_4 FILLER_25_589 ();
 sg13g2_fill_2 FILLER_25_593 ();
 sg13g2_fill_2 FILLER_25_630 ();
 sg13g2_decap_4 FILLER_25_645 ();
 sg13g2_fill_2 FILLER_25_649 ();
 sg13g2_decap_4 FILLER_25_691 ();
 sg13g2_fill_2 FILLER_25_723 ();
 sg13g2_fill_2 FILLER_25_755 ();
 sg13g2_decap_4 FILLER_25_796 ();
 sg13g2_fill_2 FILLER_25_814 ();
 sg13g2_fill_2 FILLER_25_850 ();
 sg13g2_fill_1 FILLER_25_871 ();
 sg13g2_fill_2 FILLER_25_885 ();
 sg13g2_fill_1 FILLER_25_887 ();
 sg13g2_fill_2 FILLER_25_892 ();
 sg13g2_fill_1 FILLER_25_894 ();
 sg13g2_fill_2 FILLER_25_899 ();
 sg13g2_fill_1 FILLER_25_914 ();
 sg13g2_fill_1 FILLER_25_933 ();
 sg13g2_fill_2 FILLER_25_965 ();
 sg13g2_fill_1 FILLER_25_967 ();
 sg13g2_fill_1 FILLER_25_974 ();
 sg13g2_fill_1 FILLER_25_989 ();
 sg13g2_fill_1 FILLER_25_999 ();
 sg13g2_decap_8 FILLER_25_1015 ();
 sg13g2_fill_1 FILLER_25_1022 ();
 sg13g2_fill_1 FILLER_25_1028 ();
 sg13g2_fill_2 FILLER_25_1034 ();
 sg13g2_fill_2 FILLER_25_1041 ();
 sg13g2_fill_1 FILLER_25_1043 ();
 sg13g2_fill_2 FILLER_25_1049 ();
 sg13g2_fill_1 FILLER_25_1051 ();
 sg13g2_fill_1 FILLER_25_1069 ();
 sg13g2_fill_2 FILLER_25_1118 ();
 sg13g2_decap_4 FILLER_25_1161 ();
 sg13g2_fill_1 FILLER_25_1205 ();
 sg13g2_fill_2 FILLER_25_1251 ();
 sg13g2_fill_1 FILLER_25_1293 ();
 sg13g2_fill_2 FILLER_25_1304 ();
 sg13g2_decap_8 FILLER_25_1336 ();
 sg13g2_decap_8 FILLER_25_1343 ();
 sg13g2_decap_8 FILLER_25_1350 ();
 sg13g2_decap_8 FILLER_25_1357 ();
 sg13g2_decap_8 FILLER_25_1364 ();
 sg13g2_decap_8 FILLER_25_1371 ();
 sg13g2_decap_8 FILLER_25_1378 ();
 sg13g2_decap_8 FILLER_25_1385 ();
 sg13g2_decap_8 FILLER_25_1392 ();
 sg13g2_decap_8 FILLER_25_1399 ();
 sg13g2_decap_8 FILLER_25_1406 ();
 sg13g2_decap_8 FILLER_25_1413 ();
 sg13g2_decap_8 FILLER_25_1420 ();
 sg13g2_decap_8 FILLER_25_1427 ();
 sg13g2_decap_8 FILLER_25_1434 ();
 sg13g2_decap_8 FILLER_25_1441 ();
 sg13g2_decap_8 FILLER_25_1448 ();
 sg13g2_decap_8 FILLER_25_1455 ();
 sg13g2_decap_8 FILLER_25_1462 ();
 sg13g2_decap_8 FILLER_25_1469 ();
 sg13g2_decap_8 FILLER_25_1476 ();
 sg13g2_decap_8 FILLER_25_1483 ();
 sg13g2_decap_8 FILLER_25_1490 ();
 sg13g2_decap_8 FILLER_25_1497 ();
 sg13g2_decap_8 FILLER_25_1504 ();
 sg13g2_decap_8 FILLER_25_1511 ();
 sg13g2_decap_8 FILLER_25_1518 ();
 sg13g2_decap_8 FILLER_25_1525 ();
 sg13g2_decap_8 FILLER_25_1532 ();
 sg13g2_decap_8 FILLER_25_1539 ();
 sg13g2_decap_8 FILLER_25_1546 ();
 sg13g2_decap_8 FILLER_25_1553 ();
 sg13g2_decap_8 FILLER_25_1560 ();
 sg13g2_decap_8 FILLER_25_1567 ();
 sg13g2_decap_8 FILLER_25_1574 ();
 sg13g2_decap_8 FILLER_25_1581 ();
 sg13g2_decap_8 FILLER_25_1588 ();
 sg13g2_decap_8 FILLER_25_1595 ();
 sg13g2_decap_8 FILLER_25_1602 ();
 sg13g2_decap_8 FILLER_25_1609 ();
 sg13g2_decap_8 FILLER_25_1616 ();
 sg13g2_decap_8 FILLER_25_1623 ();
 sg13g2_decap_8 FILLER_25_1630 ();
 sg13g2_decap_8 FILLER_25_1637 ();
 sg13g2_decap_8 FILLER_25_1644 ();
 sg13g2_decap_8 FILLER_25_1651 ();
 sg13g2_decap_8 FILLER_25_1658 ();
 sg13g2_decap_8 FILLER_25_1665 ();
 sg13g2_decap_8 FILLER_25_1672 ();
 sg13g2_decap_8 FILLER_25_1679 ();
 sg13g2_decap_8 FILLER_25_1686 ();
 sg13g2_decap_8 FILLER_25_1693 ();
 sg13g2_decap_8 FILLER_25_1700 ();
 sg13g2_decap_8 FILLER_25_1707 ();
 sg13g2_decap_8 FILLER_25_1714 ();
 sg13g2_decap_8 FILLER_25_1721 ();
 sg13g2_decap_8 FILLER_25_1728 ();
 sg13g2_decap_8 FILLER_25_1735 ();
 sg13g2_decap_8 FILLER_25_1742 ();
 sg13g2_decap_8 FILLER_25_1749 ();
 sg13g2_decap_8 FILLER_25_1756 ();
 sg13g2_decap_4 FILLER_25_1763 ();
 sg13g2_fill_1 FILLER_25_1767 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_4 FILLER_26_49 ();
 sg13g2_fill_2 FILLER_26_79 ();
 sg13g2_fill_1 FILLER_26_81 ();
 sg13g2_fill_2 FILLER_26_92 ();
 sg13g2_fill_1 FILLER_26_94 ();
 sg13g2_fill_1 FILLER_26_139 ();
 sg13g2_fill_1 FILLER_26_148 ();
 sg13g2_fill_2 FILLER_26_399 ();
 sg13g2_decap_4 FILLER_26_424 ();
 sg13g2_fill_1 FILLER_26_433 ();
 sg13g2_fill_2 FILLER_26_500 ();
 sg13g2_fill_2 FILLER_26_542 ();
 sg13g2_fill_1 FILLER_26_570 ();
 sg13g2_fill_2 FILLER_26_579 ();
 sg13g2_decap_4 FILLER_26_642 ();
 sg13g2_fill_2 FILLER_26_646 ();
 sg13g2_fill_1 FILLER_26_666 ();
 sg13g2_decap_4 FILLER_26_670 ();
 sg13g2_fill_2 FILLER_26_689 ();
 sg13g2_fill_1 FILLER_26_691 ();
 sg13g2_fill_2 FILLER_26_700 ();
 sg13g2_fill_1 FILLER_26_702 ();
 sg13g2_fill_2 FILLER_26_715 ();
 sg13g2_fill_2 FILLER_26_740 ();
 sg13g2_fill_2 FILLER_26_780 ();
 sg13g2_fill_1 FILLER_26_782 ();
 sg13g2_decap_4 FILLER_26_793 ();
 sg13g2_decap_8 FILLER_26_823 ();
 sg13g2_decap_4 FILLER_26_835 ();
 sg13g2_decap_8 FILLER_26_883 ();
 sg13g2_fill_1 FILLER_26_890 ();
 sg13g2_fill_2 FILLER_26_960 ();
 sg13g2_fill_2 FILLER_26_1003 ();
 sg13g2_fill_1 FILLER_26_1005 ();
 sg13g2_fill_1 FILLER_26_1032 ();
 sg13g2_decap_4 FILLER_26_1039 ();
 sg13g2_fill_1 FILLER_26_1114 ();
 sg13g2_fill_1 FILLER_26_1183 ();
 sg13g2_fill_2 FILLER_26_1256 ();
 sg13g2_fill_1 FILLER_26_1284 ();
 sg13g2_fill_1 FILLER_26_1300 ();
 sg13g2_decap_8 FILLER_26_1336 ();
 sg13g2_decap_8 FILLER_26_1343 ();
 sg13g2_decap_8 FILLER_26_1350 ();
 sg13g2_decap_8 FILLER_26_1357 ();
 sg13g2_decap_8 FILLER_26_1364 ();
 sg13g2_decap_8 FILLER_26_1371 ();
 sg13g2_decap_8 FILLER_26_1378 ();
 sg13g2_decap_8 FILLER_26_1385 ();
 sg13g2_decap_8 FILLER_26_1392 ();
 sg13g2_decap_8 FILLER_26_1399 ();
 sg13g2_decap_8 FILLER_26_1406 ();
 sg13g2_decap_8 FILLER_26_1413 ();
 sg13g2_decap_8 FILLER_26_1420 ();
 sg13g2_decap_8 FILLER_26_1427 ();
 sg13g2_decap_8 FILLER_26_1434 ();
 sg13g2_decap_8 FILLER_26_1441 ();
 sg13g2_decap_8 FILLER_26_1448 ();
 sg13g2_decap_8 FILLER_26_1455 ();
 sg13g2_decap_8 FILLER_26_1462 ();
 sg13g2_decap_8 FILLER_26_1469 ();
 sg13g2_decap_8 FILLER_26_1476 ();
 sg13g2_decap_8 FILLER_26_1483 ();
 sg13g2_decap_8 FILLER_26_1490 ();
 sg13g2_decap_8 FILLER_26_1497 ();
 sg13g2_decap_8 FILLER_26_1504 ();
 sg13g2_decap_8 FILLER_26_1511 ();
 sg13g2_decap_8 FILLER_26_1518 ();
 sg13g2_decap_8 FILLER_26_1525 ();
 sg13g2_decap_8 FILLER_26_1532 ();
 sg13g2_decap_8 FILLER_26_1539 ();
 sg13g2_decap_8 FILLER_26_1546 ();
 sg13g2_decap_8 FILLER_26_1553 ();
 sg13g2_decap_8 FILLER_26_1560 ();
 sg13g2_decap_8 FILLER_26_1567 ();
 sg13g2_decap_8 FILLER_26_1574 ();
 sg13g2_decap_8 FILLER_26_1581 ();
 sg13g2_decap_8 FILLER_26_1588 ();
 sg13g2_decap_8 FILLER_26_1595 ();
 sg13g2_decap_8 FILLER_26_1602 ();
 sg13g2_decap_8 FILLER_26_1609 ();
 sg13g2_decap_8 FILLER_26_1616 ();
 sg13g2_decap_8 FILLER_26_1623 ();
 sg13g2_decap_8 FILLER_26_1630 ();
 sg13g2_decap_8 FILLER_26_1637 ();
 sg13g2_decap_8 FILLER_26_1644 ();
 sg13g2_decap_8 FILLER_26_1651 ();
 sg13g2_decap_8 FILLER_26_1658 ();
 sg13g2_decap_8 FILLER_26_1665 ();
 sg13g2_decap_8 FILLER_26_1672 ();
 sg13g2_decap_8 FILLER_26_1679 ();
 sg13g2_decap_8 FILLER_26_1686 ();
 sg13g2_decap_8 FILLER_26_1693 ();
 sg13g2_decap_8 FILLER_26_1700 ();
 sg13g2_decap_8 FILLER_26_1707 ();
 sg13g2_decap_8 FILLER_26_1714 ();
 sg13g2_decap_8 FILLER_26_1721 ();
 sg13g2_decap_8 FILLER_26_1728 ();
 sg13g2_decap_8 FILLER_26_1735 ();
 sg13g2_decap_8 FILLER_26_1742 ();
 sg13g2_decap_8 FILLER_26_1749 ();
 sg13g2_decap_8 FILLER_26_1756 ();
 sg13g2_decap_4 FILLER_26_1763 ();
 sg13g2_fill_1 FILLER_26_1767 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_fill_2 FILLER_27_49 ();
 sg13g2_decap_4 FILLER_27_89 ();
 sg13g2_fill_1 FILLER_27_108 ();
 sg13g2_fill_1 FILLER_27_114 ();
 sg13g2_decap_4 FILLER_27_119 ();
 sg13g2_fill_2 FILLER_27_123 ();
 sg13g2_fill_2 FILLER_27_177 ();
 sg13g2_fill_1 FILLER_27_179 ();
 sg13g2_fill_1 FILLER_27_200 ();
 sg13g2_decap_8 FILLER_27_206 ();
 sg13g2_decap_8 FILLER_27_213 ();
 sg13g2_fill_1 FILLER_27_220 ();
 sg13g2_fill_2 FILLER_27_234 ();
 sg13g2_fill_2 FILLER_27_241 ();
 sg13g2_fill_2 FILLER_27_248 ();
 sg13g2_fill_1 FILLER_27_254 ();
 sg13g2_fill_2 FILLER_27_272 ();
 sg13g2_fill_1 FILLER_27_274 ();
 sg13g2_fill_2 FILLER_27_284 ();
 sg13g2_fill_2 FILLER_27_310 ();
 sg13g2_fill_1 FILLER_27_312 ();
 sg13g2_fill_2 FILLER_27_351 ();
 sg13g2_fill_1 FILLER_27_353 ();
 sg13g2_fill_1 FILLER_27_390 ();
 sg13g2_fill_2 FILLER_27_400 ();
 sg13g2_fill_2 FILLER_27_428 ();
 sg13g2_fill_1 FILLER_27_430 ();
 sg13g2_fill_1 FILLER_27_450 ();
 sg13g2_fill_2 FILLER_27_466 ();
 sg13g2_fill_1 FILLER_27_473 ();
 sg13g2_fill_1 FILLER_27_486 ();
 sg13g2_decap_4 FILLER_27_511 ();
 sg13g2_fill_2 FILLER_27_515 ();
 sg13g2_decap_8 FILLER_27_526 ();
 sg13g2_decap_8 FILLER_27_544 ();
 sg13g2_fill_2 FILLER_27_551 ();
 sg13g2_decap_4 FILLER_27_584 ();
 sg13g2_fill_1 FILLER_27_588 ();
 sg13g2_fill_2 FILLER_27_612 ();
 sg13g2_fill_2 FILLER_27_622 ();
 sg13g2_fill_1 FILLER_27_624 ();
 sg13g2_fill_1 FILLER_27_651 ();
 sg13g2_fill_2 FILLER_27_660 ();
 sg13g2_fill_1 FILLER_27_662 ();
 sg13g2_decap_4 FILLER_27_672 ();
 sg13g2_fill_2 FILLER_27_676 ();
 sg13g2_decap_8 FILLER_27_707 ();
 sg13g2_decap_8 FILLER_27_714 ();
 sg13g2_fill_1 FILLER_27_746 ();
 sg13g2_decap_4 FILLER_27_755 ();
 sg13g2_decap_8 FILLER_27_805 ();
 sg13g2_fill_1 FILLER_27_812 ();
 sg13g2_fill_2 FILLER_27_822 ();
 sg13g2_fill_2 FILLER_27_850 ();
 sg13g2_fill_2 FILLER_27_905 ();
 sg13g2_fill_2 FILLER_27_913 ();
 sg13g2_fill_1 FILLER_27_915 ();
 sg13g2_fill_1 FILLER_27_959 ();
 sg13g2_decap_8 FILLER_27_964 ();
 sg13g2_decap_4 FILLER_27_971 ();
 sg13g2_fill_1 FILLER_27_975 ();
 sg13g2_fill_1 FILLER_27_981 ();
 sg13g2_fill_2 FILLER_27_994 ();
 sg13g2_fill_1 FILLER_27_996 ();
 sg13g2_fill_2 FILLER_27_1017 ();
 sg13g2_fill_1 FILLER_27_1037 ();
 sg13g2_fill_1 FILLER_27_1043 ();
 sg13g2_fill_2 FILLER_27_1126 ();
 sg13g2_fill_1 FILLER_27_1185 ();
 sg13g2_fill_2 FILLER_27_1221 ();
 sg13g2_fill_2 FILLER_27_1231 ();
 sg13g2_fill_1 FILLER_27_1253 ();
 sg13g2_fill_2 FILLER_27_1280 ();
 sg13g2_decap_8 FILLER_27_1334 ();
 sg13g2_decap_8 FILLER_27_1341 ();
 sg13g2_decap_8 FILLER_27_1348 ();
 sg13g2_decap_8 FILLER_27_1355 ();
 sg13g2_decap_8 FILLER_27_1362 ();
 sg13g2_decap_8 FILLER_27_1369 ();
 sg13g2_decap_8 FILLER_27_1376 ();
 sg13g2_decap_8 FILLER_27_1383 ();
 sg13g2_decap_8 FILLER_27_1390 ();
 sg13g2_decap_8 FILLER_27_1397 ();
 sg13g2_decap_8 FILLER_27_1404 ();
 sg13g2_decap_8 FILLER_27_1411 ();
 sg13g2_decap_8 FILLER_27_1418 ();
 sg13g2_decap_8 FILLER_27_1425 ();
 sg13g2_decap_8 FILLER_27_1432 ();
 sg13g2_decap_8 FILLER_27_1439 ();
 sg13g2_decap_8 FILLER_27_1446 ();
 sg13g2_decap_8 FILLER_27_1453 ();
 sg13g2_decap_8 FILLER_27_1460 ();
 sg13g2_decap_8 FILLER_27_1467 ();
 sg13g2_decap_8 FILLER_27_1474 ();
 sg13g2_decap_8 FILLER_27_1481 ();
 sg13g2_decap_8 FILLER_27_1488 ();
 sg13g2_decap_8 FILLER_27_1495 ();
 sg13g2_decap_8 FILLER_27_1502 ();
 sg13g2_decap_8 FILLER_27_1509 ();
 sg13g2_decap_8 FILLER_27_1516 ();
 sg13g2_decap_8 FILLER_27_1523 ();
 sg13g2_decap_8 FILLER_27_1530 ();
 sg13g2_decap_8 FILLER_27_1537 ();
 sg13g2_decap_8 FILLER_27_1544 ();
 sg13g2_decap_8 FILLER_27_1551 ();
 sg13g2_decap_8 FILLER_27_1558 ();
 sg13g2_decap_8 FILLER_27_1565 ();
 sg13g2_decap_8 FILLER_27_1572 ();
 sg13g2_decap_8 FILLER_27_1579 ();
 sg13g2_decap_8 FILLER_27_1586 ();
 sg13g2_decap_8 FILLER_27_1593 ();
 sg13g2_decap_8 FILLER_27_1600 ();
 sg13g2_decap_8 FILLER_27_1607 ();
 sg13g2_decap_8 FILLER_27_1614 ();
 sg13g2_decap_8 FILLER_27_1621 ();
 sg13g2_decap_8 FILLER_27_1628 ();
 sg13g2_decap_8 FILLER_27_1635 ();
 sg13g2_decap_8 FILLER_27_1642 ();
 sg13g2_decap_8 FILLER_27_1649 ();
 sg13g2_decap_8 FILLER_27_1656 ();
 sg13g2_decap_8 FILLER_27_1663 ();
 sg13g2_decap_8 FILLER_27_1670 ();
 sg13g2_decap_8 FILLER_27_1677 ();
 sg13g2_decap_8 FILLER_27_1684 ();
 sg13g2_decap_8 FILLER_27_1691 ();
 sg13g2_decap_8 FILLER_27_1698 ();
 sg13g2_decap_8 FILLER_27_1705 ();
 sg13g2_decap_8 FILLER_27_1712 ();
 sg13g2_decap_8 FILLER_27_1719 ();
 sg13g2_decap_8 FILLER_27_1726 ();
 sg13g2_decap_8 FILLER_27_1733 ();
 sg13g2_decap_8 FILLER_27_1740 ();
 sg13g2_decap_8 FILLER_27_1747 ();
 sg13g2_decap_8 FILLER_27_1754 ();
 sg13g2_decap_8 FILLER_27_1761 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_4 FILLER_28_42 ();
 sg13g2_fill_1 FILLER_28_46 ();
 sg13g2_decap_4 FILLER_28_103 ();
 sg13g2_decap_8 FILLER_28_142 ();
 sg13g2_decap_4 FILLER_28_149 ();
 sg13g2_fill_1 FILLER_28_153 ();
 sg13g2_fill_2 FILLER_28_204 ();
 sg13g2_fill_1 FILLER_28_206 ();
 sg13g2_fill_2 FILLER_28_239 ();
 sg13g2_fill_1 FILLER_28_241 ();
 sg13g2_fill_2 FILLER_28_268 ();
 sg13g2_fill_2 FILLER_28_341 ();
 sg13g2_fill_2 FILLER_28_348 ();
 sg13g2_fill_1 FILLER_28_350 ();
 sg13g2_fill_2 FILLER_28_377 ();
 sg13g2_fill_1 FILLER_28_379 ();
 sg13g2_fill_2 FILLER_28_428 ();
 sg13g2_fill_1 FILLER_28_470 ();
 sg13g2_fill_1 FILLER_28_494 ();
 sg13g2_decap_4 FILLER_28_547 ();
 sg13g2_decap_8 FILLER_28_559 ();
 sg13g2_decap_8 FILLER_28_566 ();
 sg13g2_decap_8 FILLER_28_573 ();
 sg13g2_decap_4 FILLER_28_580 ();
 sg13g2_fill_1 FILLER_28_614 ();
 sg13g2_fill_1 FILLER_28_621 ();
 sg13g2_decap_4 FILLER_28_641 ();
 sg13g2_fill_1 FILLER_28_645 ();
 sg13g2_fill_2 FILLER_28_660 ();
 sg13g2_fill_2 FILLER_28_680 ();
 sg13g2_fill_1 FILLER_28_691 ();
 sg13g2_decap_8 FILLER_28_696 ();
 sg13g2_decap_4 FILLER_28_703 ();
 sg13g2_decap_4 FILLER_28_712 ();
 sg13g2_decap_8 FILLER_28_721 ();
 sg13g2_fill_2 FILLER_28_728 ();
 sg13g2_fill_1 FILLER_28_730 ();
 sg13g2_decap_4 FILLER_28_762 ();
 sg13g2_fill_2 FILLER_28_766 ();
 sg13g2_fill_2 FILLER_28_787 ();
 sg13g2_fill_1 FILLER_28_789 ();
 sg13g2_decap_4 FILLER_28_826 ();
 sg13g2_fill_2 FILLER_28_933 ();
 sg13g2_fill_2 FILLER_28_943 ();
 sg13g2_fill_2 FILLER_28_985 ();
 sg13g2_fill_1 FILLER_28_987 ();
 sg13g2_fill_2 FILLER_28_999 ();
 sg13g2_fill_1 FILLER_28_1001 ();
 sg13g2_fill_2 FILLER_28_1015 ();
 sg13g2_fill_2 FILLER_28_1025 ();
 sg13g2_fill_1 FILLER_28_1027 ();
 sg13g2_decap_4 FILLER_28_1034 ();
 sg13g2_decap_8 FILLER_28_1042 ();
 sg13g2_fill_1 FILLER_28_1049 ();
 sg13g2_fill_1 FILLER_28_1076 ();
 sg13g2_decap_4 FILLER_28_1147 ();
 sg13g2_decap_4 FILLER_28_1164 ();
 sg13g2_fill_2 FILLER_28_1168 ();
 sg13g2_decap_4 FILLER_28_1197 ();
 sg13g2_fill_1 FILLER_28_1201 ();
 sg13g2_fill_1 FILLER_28_1251 ();
 sg13g2_fill_1 FILLER_28_1261 ();
 sg13g2_fill_1 FILLER_28_1271 ();
 sg13g2_fill_1 FILLER_28_1306 ();
 sg13g2_decap_8 FILLER_28_1333 ();
 sg13g2_decap_8 FILLER_28_1340 ();
 sg13g2_decap_8 FILLER_28_1347 ();
 sg13g2_decap_8 FILLER_28_1354 ();
 sg13g2_decap_8 FILLER_28_1361 ();
 sg13g2_decap_8 FILLER_28_1368 ();
 sg13g2_decap_8 FILLER_28_1375 ();
 sg13g2_decap_8 FILLER_28_1382 ();
 sg13g2_decap_8 FILLER_28_1389 ();
 sg13g2_decap_8 FILLER_28_1396 ();
 sg13g2_decap_8 FILLER_28_1403 ();
 sg13g2_decap_8 FILLER_28_1410 ();
 sg13g2_decap_8 FILLER_28_1417 ();
 sg13g2_decap_8 FILLER_28_1424 ();
 sg13g2_decap_8 FILLER_28_1431 ();
 sg13g2_decap_8 FILLER_28_1438 ();
 sg13g2_decap_8 FILLER_28_1445 ();
 sg13g2_decap_8 FILLER_28_1452 ();
 sg13g2_decap_8 FILLER_28_1459 ();
 sg13g2_decap_8 FILLER_28_1466 ();
 sg13g2_decap_8 FILLER_28_1473 ();
 sg13g2_decap_8 FILLER_28_1480 ();
 sg13g2_decap_8 FILLER_28_1487 ();
 sg13g2_decap_8 FILLER_28_1494 ();
 sg13g2_decap_8 FILLER_28_1501 ();
 sg13g2_decap_8 FILLER_28_1508 ();
 sg13g2_decap_8 FILLER_28_1515 ();
 sg13g2_decap_8 FILLER_28_1522 ();
 sg13g2_decap_8 FILLER_28_1529 ();
 sg13g2_decap_8 FILLER_28_1536 ();
 sg13g2_decap_8 FILLER_28_1543 ();
 sg13g2_decap_8 FILLER_28_1550 ();
 sg13g2_decap_8 FILLER_28_1557 ();
 sg13g2_decap_8 FILLER_28_1564 ();
 sg13g2_decap_8 FILLER_28_1571 ();
 sg13g2_decap_8 FILLER_28_1578 ();
 sg13g2_decap_8 FILLER_28_1585 ();
 sg13g2_decap_8 FILLER_28_1592 ();
 sg13g2_decap_8 FILLER_28_1599 ();
 sg13g2_decap_8 FILLER_28_1606 ();
 sg13g2_decap_8 FILLER_28_1613 ();
 sg13g2_decap_8 FILLER_28_1620 ();
 sg13g2_decap_8 FILLER_28_1627 ();
 sg13g2_decap_8 FILLER_28_1634 ();
 sg13g2_decap_8 FILLER_28_1641 ();
 sg13g2_decap_8 FILLER_28_1648 ();
 sg13g2_decap_8 FILLER_28_1655 ();
 sg13g2_decap_8 FILLER_28_1662 ();
 sg13g2_decap_8 FILLER_28_1669 ();
 sg13g2_decap_8 FILLER_28_1676 ();
 sg13g2_decap_8 FILLER_28_1683 ();
 sg13g2_decap_8 FILLER_28_1690 ();
 sg13g2_decap_8 FILLER_28_1697 ();
 sg13g2_decap_8 FILLER_28_1704 ();
 sg13g2_decap_8 FILLER_28_1711 ();
 sg13g2_decap_8 FILLER_28_1718 ();
 sg13g2_decap_8 FILLER_28_1725 ();
 sg13g2_decap_8 FILLER_28_1732 ();
 sg13g2_decap_8 FILLER_28_1739 ();
 sg13g2_decap_8 FILLER_28_1746 ();
 sg13g2_decap_8 FILLER_28_1753 ();
 sg13g2_decap_8 FILLER_28_1760 ();
 sg13g2_fill_1 FILLER_28_1767 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_fill_2 FILLER_29_70 ();
 sg13g2_fill_1 FILLER_29_135 ();
 sg13g2_fill_1 FILLER_29_162 ();
 sg13g2_decap_4 FILLER_29_225 ();
 sg13g2_fill_2 FILLER_29_314 ();
 sg13g2_fill_1 FILLER_29_316 ();
 sg13g2_fill_1 FILLER_29_326 ();
 sg13g2_fill_2 FILLER_29_332 ();
 sg13g2_fill_1 FILLER_29_334 ();
 sg13g2_fill_2 FILLER_29_380 ();
 sg13g2_fill_1 FILLER_29_382 ();
 sg13g2_fill_2 FILLER_29_411 ();
 sg13g2_fill_1 FILLER_29_423 ();
 sg13g2_decap_4 FILLER_29_429 ();
 sg13g2_fill_1 FILLER_29_433 ();
 sg13g2_fill_2 FILLER_29_470 ();
 sg13g2_fill_1 FILLER_29_472 ();
 sg13g2_fill_2 FILLER_29_504 ();
 sg13g2_decap_4 FILLER_29_563 ();
 sg13g2_fill_2 FILLER_29_583 ();
 sg13g2_fill_1 FILLER_29_585 ();
 sg13g2_fill_1 FILLER_29_600 ();
 sg13g2_decap_4 FILLER_29_618 ();
 sg13g2_fill_1 FILLER_29_622 ();
 sg13g2_decap_4 FILLER_29_626 ();
 sg13g2_fill_1 FILLER_29_630 ();
 sg13g2_decap_4 FILLER_29_640 ();
 sg13g2_fill_2 FILLER_29_644 ();
 sg13g2_decap_8 FILLER_29_672 ();
 sg13g2_fill_2 FILLER_29_679 ();
 sg13g2_fill_2 FILLER_29_694 ();
 sg13g2_fill_1 FILLER_29_696 ();
 sg13g2_fill_2 FILLER_29_716 ();
 sg13g2_fill_2 FILLER_29_723 ();
 sg13g2_fill_2 FILLER_29_730 ();
 sg13g2_fill_1 FILLER_29_732 ();
 sg13g2_decap_4 FILLER_29_753 ();
 sg13g2_fill_1 FILLER_29_757 ();
 sg13g2_fill_1 FILLER_29_766 ();
 sg13g2_fill_2 FILLER_29_793 ();
 sg13g2_fill_1 FILLER_29_795 ();
 sg13g2_fill_2 FILLER_29_810 ();
 sg13g2_fill_1 FILLER_29_812 ();
 sg13g2_decap_8 FILLER_29_824 ();
 sg13g2_decap_8 FILLER_29_831 ();
 sg13g2_decap_8 FILLER_29_838 ();
 sg13g2_decap_8 FILLER_29_845 ();
 sg13g2_fill_2 FILLER_29_852 ();
 sg13g2_fill_2 FILLER_29_895 ();
 sg13g2_fill_2 FILLER_29_906 ();
 sg13g2_fill_1 FILLER_29_908 ();
 sg13g2_fill_2 FILLER_29_945 ();
 sg13g2_fill_1 FILLER_29_947 ();
 sg13g2_decap_4 FILLER_29_978 ();
 sg13g2_decap_4 FILLER_29_999 ();
 sg13g2_fill_1 FILLER_29_1003 ();
 sg13g2_fill_2 FILLER_29_1052 ();
 sg13g2_fill_1 FILLER_29_1054 ();
 sg13g2_fill_1 FILLER_29_1086 ();
 sg13g2_fill_2 FILLER_29_1255 ();
 sg13g2_fill_1 FILLER_29_1257 ();
 sg13g2_fill_2 FILLER_29_1293 ();
 sg13g2_fill_1 FILLER_29_1295 ();
 sg13g2_decap_8 FILLER_29_1340 ();
 sg13g2_decap_8 FILLER_29_1347 ();
 sg13g2_decap_8 FILLER_29_1354 ();
 sg13g2_decap_8 FILLER_29_1361 ();
 sg13g2_decap_8 FILLER_29_1368 ();
 sg13g2_decap_8 FILLER_29_1375 ();
 sg13g2_decap_8 FILLER_29_1382 ();
 sg13g2_decap_8 FILLER_29_1389 ();
 sg13g2_decap_8 FILLER_29_1396 ();
 sg13g2_decap_8 FILLER_29_1403 ();
 sg13g2_decap_8 FILLER_29_1410 ();
 sg13g2_decap_8 FILLER_29_1417 ();
 sg13g2_decap_8 FILLER_29_1424 ();
 sg13g2_decap_8 FILLER_29_1431 ();
 sg13g2_decap_8 FILLER_29_1438 ();
 sg13g2_decap_8 FILLER_29_1445 ();
 sg13g2_decap_8 FILLER_29_1452 ();
 sg13g2_decap_8 FILLER_29_1459 ();
 sg13g2_decap_8 FILLER_29_1466 ();
 sg13g2_decap_8 FILLER_29_1473 ();
 sg13g2_decap_8 FILLER_29_1480 ();
 sg13g2_decap_8 FILLER_29_1487 ();
 sg13g2_decap_8 FILLER_29_1494 ();
 sg13g2_decap_8 FILLER_29_1501 ();
 sg13g2_decap_8 FILLER_29_1508 ();
 sg13g2_decap_8 FILLER_29_1515 ();
 sg13g2_decap_8 FILLER_29_1522 ();
 sg13g2_decap_8 FILLER_29_1529 ();
 sg13g2_decap_8 FILLER_29_1536 ();
 sg13g2_decap_8 FILLER_29_1543 ();
 sg13g2_decap_8 FILLER_29_1550 ();
 sg13g2_decap_8 FILLER_29_1557 ();
 sg13g2_decap_8 FILLER_29_1564 ();
 sg13g2_decap_8 FILLER_29_1571 ();
 sg13g2_decap_8 FILLER_29_1578 ();
 sg13g2_decap_8 FILLER_29_1585 ();
 sg13g2_decap_8 FILLER_29_1592 ();
 sg13g2_decap_8 FILLER_29_1599 ();
 sg13g2_decap_8 FILLER_29_1606 ();
 sg13g2_decap_8 FILLER_29_1613 ();
 sg13g2_decap_8 FILLER_29_1620 ();
 sg13g2_decap_8 FILLER_29_1627 ();
 sg13g2_decap_8 FILLER_29_1634 ();
 sg13g2_decap_8 FILLER_29_1641 ();
 sg13g2_decap_8 FILLER_29_1648 ();
 sg13g2_decap_8 FILLER_29_1655 ();
 sg13g2_decap_8 FILLER_29_1662 ();
 sg13g2_decap_8 FILLER_29_1669 ();
 sg13g2_decap_8 FILLER_29_1676 ();
 sg13g2_decap_8 FILLER_29_1683 ();
 sg13g2_decap_8 FILLER_29_1690 ();
 sg13g2_decap_8 FILLER_29_1697 ();
 sg13g2_decap_8 FILLER_29_1704 ();
 sg13g2_decap_8 FILLER_29_1711 ();
 sg13g2_decap_8 FILLER_29_1718 ();
 sg13g2_decap_8 FILLER_29_1725 ();
 sg13g2_decap_8 FILLER_29_1732 ();
 sg13g2_decap_8 FILLER_29_1739 ();
 sg13g2_decap_8 FILLER_29_1746 ();
 sg13g2_decap_8 FILLER_29_1753 ();
 sg13g2_decap_8 FILLER_29_1760 ();
 sg13g2_fill_1 FILLER_29_1767 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_4 FILLER_30_49 ();
 sg13g2_fill_1 FILLER_30_53 ();
 sg13g2_fill_2 FILLER_30_80 ();
 sg13g2_fill_1 FILLER_30_113 ();
 sg13g2_fill_2 FILLER_30_149 ();
 sg13g2_fill_2 FILLER_30_170 ();
 sg13g2_fill_1 FILLER_30_172 ();
 sg13g2_fill_1 FILLER_30_184 ();
 sg13g2_fill_2 FILLER_30_190 ();
 sg13g2_fill_1 FILLER_30_197 ();
 sg13g2_fill_2 FILLER_30_207 ();
 sg13g2_fill_1 FILLER_30_209 ();
 sg13g2_fill_1 FILLER_30_223 ();
 sg13g2_fill_2 FILLER_30_264 ();
 sg13g2_fill_2 FILLER_30_271 ();
 sg13g2_fill_2 FILLER_30_296 ();
 sg13g2_fill_1 FILLER_30_298 ();
 sg13g2_decap_4 FILLER_30_304 ();
 sg13g2_fill_2 FILLER_30_308 ();
 sg13g2_fill_2 FILLER_30_341 ();
 sg13g2_fill_2 FILLER_30_428 ();
 sg13g2_fill_2 FILLER_30_509 ();
 sg13g2_decap_8 FILLER_30_537 ();
 sg13g2_decap_8 FILLER_30_544 ();
 sg13g2_decap_8 FILLER_30_551 ();
 sg13g2_decap_8 FILLER_30_558 ();
 sg13g2_fill_2 FILLER_30_565 ();
 sg13g2_decap_8 FILLER_30_575 ();
 sg13g2_decap_4 FILLER_30_582 ();
 sg13g2_fill_2 FILLER_30_647 ();
 sg13g2_decap_4 FILLER_30_670 ();
 sg13g2_fill_2 FILLER_30_709 ();
 sg13g2_decap_4 FILLER_30_723 ();
 sg13g2_fill_2 FILLER_30_766 ();
 sg13g2_fill_1 FILLER_30_768 ();
 sg13g2_decap_4 FILLER_30_781 ();
 sg13g2_fill_2 FILLER_30_801 ();
 sg13g2_fill_1 FILLER_30_803 ();
 sg13g2_fill_1 FILLER_30_813 ();
 sg13g2_fill_2 FILLER_30_927 ();
 sg13g2_fill_1 FILLER_30_929 ();
 sg13g2_fill_1 FILLER_30_944 ();
 sg13g2_fill_2 FILLER_30_959 ();
 sg13g2_decap_4 FILLER_30_984 ();
 sg13g2_fill_2 FILLER_30_988 ();
 sg13g2_fill_2 FILLER_30_1020 ();
 sg13g2_fill_2 FILLER_30_1027 ();
 sg13g2_fill_2 FILLER_30_1039 ();
 sg13g2_fill_2 FILLER_30_1081 ();
 sg13g2_fill_2 FILLER_30_1094 ();
 sg13g2_decap_4 FILLER_30_1163 ();
 sg13g2_decap_4 FILLER_30_1176 ();
 sg13g2_fill_1 FILLER_30_1210 ();
 sg13g2_decap_8 FILLER_30_1336 ();
 sg13g2_decap_8 FILLER_30_1343 ();
 sg13g2_decap_8 FILLER_30_1350 ();
 sg13g2_decap_8 FILLER_30_1357 ();
 sg13g2_decap_8 FILLER_30_1364 ();
 sg13g2_decap_8 FILLER_30_1371 ();
 sg13g2_decap_8 FILLER_30_1378 ();
 sg13g2_decap_8 FILLER_30_1385 ();
 sg13g2_decap_8 FILLER_30_1392 ();
 sg13g2_decap_8 FILLER_30_1399 ();
 sg13g2_decap_8 FILLER_30_1406 ();
 sg13g2_decap_8 FILLER_30_1413 ();
 sg13g2_decap_8 FILLER_30_1420 ();
 sg13g2_decap_8 FILLER_30_1427 ();
 sg13g2_decap_8 FILLER_30_1434 ();
 sg13g2_decap_8 FILLER_30_1441 ();
 sg13g2_decap_8 FILLER_30_1448 ();
 sg13g2_decap_8 FILLER_30_1455 ();
 sg13g2_decap_8 FILLER_30_1462 ();
 sg13g2_decap_8 FILLER_30_1469 ();
 sg13g2_decap_8 FILLER_30_1476 ();
 sg13g2_decap_8 FILLER_30_1483 ();
 sg13g2_decap_8 FILLER_30_1490 ();
 sg13g2_decap_8 FILLER_30_1497 ();
 sg13g2_decap_8 FILLER_30_1504 ();
 sg13g2_decap_8 FILLER_30_1511 ();
 sg13g2_decap_8 FILLER_30_1518 ();
 sg13g2_decap_8 FILLER_30_1525 ();
 sg13g2_decap_8 FILLER_30_1532 ();
 sg13g2_decap_8 FILLER_30_1539 ();
 sg13g2_decap_8 FILLER_30_1546 ();
 sg13g2_decap_8 FILLER_30_1553 ();
 sg13g2_decap_8 FILLER_30_1560 ();
 sg13g2_decap_8 FILLER_30_1567 ();
 sg13g2_decap_8 FILLER_30_1574 ();
 sg13g2_decap_8 FILLER_30_1581 ();
 sg13g2_decap_8 FILLER_30_1588 ();
 sg13g2_decap_8 FILLER_30_1595 ();
 sg13g2_decap_8 FILLER_30_1602 ();
 sg13g2_decap_8 FILLER_30_1609 ();
 sg13g2_decap_8 FILLER_30_1616 ();
 sg13g2_decap_8 FILLER_30_1623 ();
 sg13g2_decap_8 FILLER_30_1630 ();
 sg13g2_decap_8 FILLER_30_1637 ();
 sg13g2_decap_8 FILLER_30_1644 ();
 sg13g2_decap_8 FILLER_30_1651 ();
 sg13g2_decap_8 FILLER_30_1658 ();
 sg13g2_decap_8 FILLER_30_1665 ();
 sg13g2_decap_8 FILLER_30_1672 ();
 sg13g2_decap_8 FILLER_30_1679 ();
 sg13g2_decap_8 FILLER_30_1686 ();
 sg13g2_decap_8 FILLER_30_1693 ();
 sg13g2_decap_8 FILLER_30_1700 ();
 sg13g2_decap_8 FILLER_30_1707 ();
 sg13g2_decap_8 FILLER_30_1714 ();
 sg13g2_decap_8 FILLER_30_1721 ();
 sg13g2_decap_8 FILLER_30_1728 ();
 sg13g2_decap_8 FILLER_30_1735 ();
 sg13g2_decap_8 FILLER_30_1742 ();
 sg13g2_decap_8 FILLER_30_1749 ();
 sg13g2_decap_8 FILLER_30_1756 ();
 sg13g2_decap_4 FILLER_30_1763 ();
 sg13g2_fill_1 FILLER_30_1767 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_fill_2 FILLER_31_77 ();
 sg13g2_fill_2 FILLER_31_124 ();
 sg13g2_decap_8 FILLER_31_130 ();
 sg13g2_fill_1 FILLER_31_163 ();
 sg13g2_fill_2 FILLER_31_225 ();
 sg13g2_fill_2 FILLER_31_269 ();
 sg13g2_decap_4 FILLER_31_312 ();
 sg13g2_fill_2 FILLER_31_373 ();
 sg13g2_fill_2 FILLER_31_406 ();
 sg13g2_fill_1 FILLER_31_408 ();
 sg13g2_decap_4 FILLER_31_421 ();
 sg13g2_fill_1 FILLER_31_425 ();
 sg13g2_fill_2 FILLER_31_431 ();
 sg13g2_fill_2 FILLER_31_477 ();
 sg13g2_decap_4 FILLER_31_518 ();
 sg13g2_fill_1 FILLER_31_525 ();
 sg13g2_fill_2 FILLER_31_578 ();
 sg13g2_fill_1 FILLER_31_580 ();
 sg13g2_fill_1 FILLER_31_603 ();
 sg13g2_fill_1 FILLER_31_609 ();
 sg13g2_fill_1 FILLER_31_620 ();
 sg13g2_decap_8 FILLER_31_630 ();
 sg13g2_decap_8 FILLER_31_637 ();
 sg13g2_fill_1 FILLER_31_669 ();
 sg13g2_fill_2 FILLER_31_682 ();
 sg13g2_decap_4 FILLER_31_701 ();
 sg13g2_decap_8 FILLER_31_718 ();
 sg13g2_decap_8 FILLER_31_725 ();
 sg13g2_fill_2 FILLER_31_732 ();
 sg13g2_fill_1 FILLER_31_734 ();
 sg13g2_decap_8 FILLER_31_746 ();
 sg13g2_fill_2 FILLER_31_753 ();
 sg13g2_fill_1 FILLER_31_755 ();
 sg13g2_fill_1 FILLER_31_767 ();
 sg13g2_decap_4 FILLER_31_777 ();
 sg13g2_fill_1 FILLER_31_781 ();
 sg13g2_fill_1 FILLER_31_793 ();
 sg13g2_decap_8 FILLER_31_824 ();
 sg13g2_decap_8 FILLER_31_831 ();
 sg13g2_decap_8 FILLER_31_838 ();
 sg13g2_decap_8 FILLER_31_845 ();
 sg13g2_decap_8 FILLER_31_852 ();
 sg13g2_fill_2 FILLER_31_859 ();
 sg13g2_fill_1 FILLER_31_861 ();
 sg13g2_decap_4 FILLER_31_866 ();
 sg13g2_fill_1 FILLER_31_870 ();
 sg13g2_fill_1 FILLER_31_908 ();
 sg13g2_fill_1 FILLER_31_914 ();
 sg13g2_fill_2 FILLER_31_928 ();
 sg13g2_fill_1 FILLER_31_930 ();
 sg13g2_decap_8 FILLER_31_985 ();
 sg13g2_fill_2 FILLER_31_992 ();
 sg13g2_fill_2 FILLER_31_999 ();
 sg13g2_fill_1 FILLER_31_1006 ();
 sg13g2_decap_4 FILLER_31_1012 ();
 sg13g2_fill_2 FILLER_31_1092 ();
 sg13g2_fill_1 FILLER_31_1128 ();
 sg13g2_fill_1 FILLER_31_1143 ();
 sg13g2_fill_2 FILLER_31_1170 ();
 sg13g2_fill_2 FILLER_31_1180 ();
 sg13g2_fill_2 FILLER_31_1241 ();
 sg13g2_fill_1 FILLER_31_1243 ();
 sg13g2_fill_2 FILLER_31_1258 ();
 sg13g2_fill_2 FILLER_31_1277 ();
 sg13g2_fill_1 FILLER_31_1279 ();
 sg13g2_fill_2 FILLER_31_1295 ();
 sg13g2_decap_8 FILLER_31_1332 ();
 sg13g2_decap_8 FILLER_31_1339 ();
 sg13g2_decap_8 FILLER_31_1346 ();
 sg13g2_decap_8 FILLER_31_1353 ();
 sg13g2_decap_8 FILLER_31_1360 ();
 sg13g2_decap_8 FILLER_31_1367 ();
 sg13g2_decap_8 FILLER_31_1374 ();
 sg13g2_decap_8 FILLER_31_1381 ();
 sg13g2_decap_8 FILLER_31_1388 ();
 sg13g2_decap_8 FILLER_31_1395 ();
 sg13g2_decap_8 FILLER_31_1402 ();
 sg13g2_decap_8 FILLER_31_1409 ();
 sg13g2_decap_8 FILLER_31_1416 ();
 sg13g2_decap_8 FILLER_31_1423 ();
 sg13g2_decap_8 FILLER_31_1430 ();
 sg13g2_decap_8 FILLER_31_1437 ();
 sg13g2_decap_8 FILLER_31_1444 ();
 sg13g2_decap_8 FILLER_31_1451 ();
 sg13g2_decap_8 FILLER_31_1458 ();
 sg13g2_decap_8 FILLER_31_1465 ();
 sg13g2_decap_8 FILLER_31_1472 ();
 sg13g2_decap_8 FILLER_31_1479 ();
 sg13g2_decap_8 FILLER_31_1486 ();
 sg13g2_decap_8 FILLER_31_1493 ();
 sg13g2_decap_8 FILLER_31_1500 ();
 sg13g2_decap_8 FILLER_31_1507 ();
 sg13g2_decap_8 FILLER_31_1514 ();
 sg13g2_decap_8 FILLER_31_1521 ();
 sg13g2_decap_8 FILLER_31_1528 ();
 sg13g2_decap_8 FILLER_31_1535 ();
 sg13g2_decap_8 FILLER_31_1542 ();
 sg13g2_decap_8 FILLER_31_1549 ();
 sg13g2_decap_8 FILLER_31_1556 ();
 sg13g2_decap_8 FILLER_31_1563 ();
 sg13g2_decap_8 FILLER_31_1570 ();
 sg13g2_decap_8 FILLER_31_1577 ();
 sg13g2_decap_8 FILLER_31_1584 ();
 sg13g2_decap_8 FILLER_31_1591 ();
 sg13g2_decap_8 FILLER_31_1598 ();
 sg13g2_decap_8 FILLER_31_1605 ();
 sg13g2_decap_8 FILLER_31_1612 ();
 sg13g2_decap_8 FILLER_31_1619 ();
 sg13g2_decap_8 FILLER_31_1626 ();
 sg13g2_decap_8 FILLER_31_1633 ();
 sg13g2_decap_8 FILLER_31_1640 ();
 sg13g2_decap_8 FILLER_31_1647 ();
 sg13g2_decap_8 FILLER_31_1654 ();
 sg13g2_decap_8 FILLER_31_1661 ();
 sg13g2_decap_8 FILLER_31_1668 ();
 sg13g2_decap_8 FILLER_31_1675 ();
 sg13g2_decap_8 FILLER_31_1682 ();
 sg13g2_decap_8 FILLER_31_1689 ();
 sg13g2_decap_8 FILLER_31_1696 ();
 sg13g2_decap_8 FILLER_31_1703 ();
 sg13g2_decap_8 FILLER_31_1710 ();
 sg13g2_decap_8 FILLER_31_1717 ();
 sg13g2_decap_8 FILLER_31_1724 ();
 sg13g2_decap_8 FILLER_31_1731 ();
 sg13g2_decap_8 FILLER_31_1738 ();
 sg13g2_decap_8 FILLER_31_1745 ();
 sg13g2_decap_8 FILLER_31_1752 ();
 sg13g2_decap_8 FILLER_31_1759 ();
 sg13g2_fill_2 FILLER_31_1766 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_8 FILLER_32_84 ();
 sg13g2_decap_8 FILLER_32_91 ();
 sg13g2_decap_8 FILLER_32_98 ();
 sg13g2_decap_8 FILLER_32_105 ();
 sg13g2_decap_8 FILLER_32_112 ();
 sg13g2_fill_2 FILLER_32_119 ();
 sg13g2_fill_1 FILLER_32_121 ();
 sg13g2_decap_8 FILLER_32_130 ();
 sg13g2_fill_2 FILLER_32_163 ();
 sg13g2_fill_2 FILLER_32_174 ();
 sg13g2_fill_2 FILLER_32_230 ();
 sg13g2_fill_1 FILLER_32_232 ();
 sg13g2_fill_2 FILLER_32_243 ();
 sg13g2_fill_1 FILLER_32_245 ();
 sg13g2_fill_2 FILLER_32_251 ();
 sg13g2_fill_1 FILLER_32_294 ();
 sg13g2_fill_2 FILLER_32_371 ();
 sg13g2_decap_4 FILLER_32_378 ();
 sg13g2_fill_1 FILLER_32_382 ();
 sg13g2_decap_4 FILLER_32_387 ();
 sg13g2_fill_2 FILLER_32_391 ();
 sg13g2_fill_2 FILLER_32_397 ();
 sg13g2_fill_2 FILLER_32_404 ();
 sg13g2_fill_1 FILLER_32_411 ();
 sg13g2_fill_2 FILLER_32_435 ();
 sg13g2_fill_2 FILLER_32_478 ();
 sg13g2_fill_1 FILLER_32_486 ();
 sg13g2_decap_8 FILLER_32_513 ();
 sg13g2_decap_8 FILLER_32_520 ();
 sg13g2_decap_4 FILLER_32_527 ();
 sg13g2_fill_1 FILLER_32_531 ();
 sg13g2_fill_1 FILLER_32_542 ();
 sg13g2_decap_4 FILLER_32_548 ();
 sg13g2_fill_1 FILLER_32_552 ();
 sg13g2_decap_4 FILLER_32_557 ();
 sg13g2_fill_2 FILLER_32_561 ();
 sg13g2_decap_4 FILLER_32_589 ();
 sg13g2_fill_2 FILLER_32_593 ();
 sg13g2_fill_2 FILLER_32_599 ();
 sg13g2_decap_4 FILLER_32_650 ();
 sg13g2_fill_2 FILLER_32_676 ();
 sg13g2_fill_1 FILLER_32_690 ();
 sg13g2_decap_8 FILLER_32_696 ();
 sg13g2_fill_2 FILLER_32_703 ();
 sg13g2_decap_8 FILLER_32_723 ();
 sg13g2_decap_4 FILLER_32_730 ();
 sg13g2_decap_4 FILLER_32_748 ();
 sg13g2_fill_2 FILLER_32_752 ();
 sg13g2_decap_4 FILLER_32_791 ();
 sg13g2_decap_4 FILLER_32_888 ();
 sg13g2_decap_4 FILLER_32_905 ();
 sg13g2_fill_1 FILLER_32_909 ();
 sg13g2_fill_1 FILLER_32_958 ();
 sg13g2_fill_1 FILLER_32_1004 ();
 sg13g2_decap_4 FILLER_32_1023 ();
 sg13g2_fill_2 FILLER_32_1027 ();
 sg13g2_fill_2 FILLER_32_1067 ();
 sg13g2_fill_1 FILLER_32_1139 ();
 sg13g2_fill_1 FILLER_32_1169 ();
 sg13g2_fill_1 FILLER_32_1183 ();
 sg13g2_fill_1 FILLER_32_1197 ();
 sg13g2_decap_8 FILLER_32_1263 ();
 sg13g2_fill_1 FILLER_32_1270 ();
 sg13g2_fill_2 FILLER_32_1285 ();
 sg13g2_fill_1 FILLER_32_1287 ();
 sg13g2_decap_8 FILLER_32_1324 ();
 sg13g2_decap_8 FILLER_32_1331 ();
 sg13g2_decap_8 FILLER_32_1338 ();
 sg13g2_decap_8 FILLER_32_1345 ();
 sg13g2_decap_8 FILLER_32_1352 ();
 sg13g2_decap_8 FILLER_32_1359 ();
 sg13g2_decap_8 FILLER_32_1366 ();
 sg13g2_decap_8 FILLER_32_1373 ();
 sg13g2_decap_8 FILLER_32_1380 ();
 sg13g2_decap_8 FILLER_32_1387 ();
 sg13g2_decap_8 FILLER_32_1394 ();
 sg13g2_decap_8 FILLER_32_1401 ();
 sg13g2_decap_8 FILLER_32_1408 ();
 sg13g2_decap_8 FILLER_32_1415 ();
 sg13g2_decap_8 FILLER_32_1422 ();
 sg13g2_decap_8 FILLER_32_1429 ();
 sg13g2_decap_8 FILLER_32_1436 ();
 sg13g2_decap_8 FILLER_32_1443 ();
 sg13g2_decap_8 FILLER_32_1450 ();
 sg13g2_decap_8 FILLER_32_1457 ();
 sg13g2_decap_8 FILLER_32_1464 ();
 sg13g2_decap_8 FILLER_32_1471 ();
 sg13g2_decap_8 FILLER_32_1478 ();
 sg13g2_decap_8 FILLER_32_1485 ();
 sg13g2_decap_8 FILLER_32_1492 ();
 sg13g2_decap_8 FILLER_32_1499 ();
 sg13g2_decap_8 FILLER_32_1506 ();
 sg13g2_decap_8 FILLER_32_1513 ();
 sg13g2_decap_8 FILLER_32_1520 ();
 sg13g2_decap_8 FILLER_32_1527 ();
 sg13g2_decap_8 FILLER_32_1534 ();
 sg13g2_decap_8 FILLER_32_1541 ();
 sg13g2_decap_8 FILLER_32_1548 ();
 sg13g2_decap_8 FILLER_32_1555 ();
 sg13g2_decap_8 FILLER_32_1562 ();
 sg13g2_decap_8 FILLER_32_1569 ();
 sg13g2_decap_8 FILLER_32_1576 ();
 sg13g2_decap_8 FILLER_32_1583 ();
 sg13g2_decap_8 FILLER_32_1590 ();
 sg13g2_decap_8 FILLER_32_1597 ();
 sg13g2_decap_8 FILLER_32_1604 ();
 sg13g2_decap_8 FILLER_32_1611 ();
 sg13g2_decap_8 FILLER_32_1618 ();
 sg13g2_decap_8 FILLER_32_1625 ();
 sg13g2_decap_8 FILLER_32_1632 ();
 sg13g2_decap_8 FILLER_32_1639 ();
 sg13g2_decap_8 FILLER_32_1646 ();
 sg13g2_decap_8 FILLER_32_1653 ();
 sg13g2_decap_8 FILLER_32_1660 ();
 sg13g2_decap_8 FILLER_32_1667 ();
 sg13g2_decap_8 FILLER_32_1674 ();
 sg13g2_decap_8 FILLER_32_1681 ();
 sg13g2_decap_8 FILLER_32_1688 ();
 sg13g2_decap_8 FILLER_32_1695 ();
 sg13g2_decap_8 FILLER_32_1702 ();
 sg13g2_decap_8 FILLER_32_1709 ();
 sg13g2_decap_8 FILLER_32_1716 ();
 sg13g2_decap_8 FILLER_32_1723 ();
 sg13g2_decap_8 FILLER_32_1730 ();
 sg13g2_decap_8 FILLER_32_1737 ();
 sg13g2_decap_8 FILLER_32_1744 ();
 sg13g2_decap_8 FILLER_32_1751 ();
 sg13g2_decap_8 FILLER_32_1758 ();
 sg13g2_fill_2 FILLER_32_1765 ();
 sg13g2_fill_1 FILLER_32_1767 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_decap_8 FILLER_33_91 ();
 sg13g2_decap_8 FILLER_33_98 ();
 sg13g2_decap_8 FILLER_33_105 ();
 sg13g2_decap_8 FILLER_33_112 ();
 sg13g2_decap_8 FILLER_33_119 ();
 sg13g2_decap_8 FILLER_33_126 ();
 sg13g2_decap_8 FILLER_33_133 ();
 sg13g2_decap_8 FILLER_33_140 ();
 sg13g2_fill_2 FILLER_33_147 ();
 sg13g2_fill_1 FILLER_33_149 ();
 sg13g2_fill_2 FILLER_33_185 ();
 sg13g2_fill_1 FILLER_33_187 ();
 sg13g2_fill_2 FILLER_33_268 ();
 sg13g2_decap_4 FILLER_33_328 ();
 sg13g2_fill_1 FILLER_33_351 ();
 sg13g2_fill_1 FILLER_33_360 ();
 sg13g2_decap_8 FILLER_33_391 ();
 sg13g2_fill_1 FILLER_33_398 ();
 sg13g2_fill_1 FILLER_33_434 ();
 sg13g2_fill_2 FILLER_33_494 ();
 sg13g2_fill_2 FILLER_33_577 ();
 sg13g2_fill_2 FILLER_33_613 ();
 sg13g2_decap_8 FILLER_33_630 ();
 sg13g2_fill_2 FILLER_33_637 ();
 sg13g2_fill_1 FILLER_33_639 ();
 sg13g2_fill_1 FILLER_33_653 ();
 sg13g2_fill_2 FILLER_33_659 ();
 sg13g2_fill_1 FILLER_33_661 ();
 sg13g2_fill_1 FILLER_33_693 ();
 sg13g2_fill_2 FILLER_33_729 ();
 sg13g2_fill_2 FILLER_33_749 ();
 sg13g2_fill_1 FILLER_33_790 ();
 sg13g2_fill_1 FILLER_33_796 ();
 sg13g2_decap_8 FILLER_33_841 ();
 sg13g2_decap_8 FILLER_33_848 ();
 sg13g2_decap_4 FILLER_33_855 ();
 sg13g2_fill_2 FILLER_33_868 ();
 sg13g2_fill_1 FILLER_33_870 ();
 sg13g2_fill_2 FILLER_33_925 ();
 sg13g2_fill_1 FILLER_33_962 ();
 sg13g2_decap_8 FILLER_33_982 ();
 sg13g2_decap_4 FILLER_33_989 ();
 sg13g2_fill_2 FILLER_33_1026 ();
 sg13g2_fill_1 FILLER_33_1033 ();
 sg13g2_fill_1 FILLER_33_1094 ();
 sg13g2_fill_1 FILLER_33_1135 ();
 sg13g2_fill_1 FILLER_33_1146 ();
 sg13g2_fill_1 FILLER_33_1175 ();
 sg13g2_fill_1 FILLER_33_1204 ();
 sg13g2_fill_2 FILLER_33_1215 ();
 sg13g2_fill_1 FILLER_33_1217 ();
 sg13g2_decap_4 FILLER_33_1231 ();
 sg13g2_fill_1 FILLER_33_1235 ();
 sg13g2_fill_2 FILLER_33_1246 ();
 sg13g2_fill_1 FILLER_33_1248 ();
 sg13g2_decap_8 FILLER_33_1323 ();
 sg13g2_decap_8 FILLER_33_1330 ();
 sg13g2_decap_8 FILLER_33_1337 ();
 sg13g2_decap_8 FILLER_33_1344 ();
 sg13g2_decap_8 FILLER_33_1351 ();
 sg13g2_decap_8 FILLER_33_1358 ();
 sg13g2_decap_8 FILLER_33_1365 ();
 sg13g2_decap_8 FILLER_33_1372 ();
 sg13g2_decap_8 FILLER_33_1379 ();
 sg13g2_decap_8 FILLER_33_1386 ();
 sg13g2_decap_8 FILLER_33_1393 ();
 sg13g2_decap_8 FILLER_33_1400 ();
 sg13g2_decap_8 FILLER_33_1407 ();
 sg13g2_decap_8 FILLER_33_1414 ();
 sg13g2_decap_8 FILLER_33_1421 ();
 sg13g2_decap_8 FILLER_33_1428 ();
 sg13g2_decap_8 FILLER_33_1435 ();
 sg13g2_decap_8 FILLER_33_1442 ();
 sg13g2_decap_8 FILLER_33_1449 ();
 sg13g2_decap_8 FILLER_33_1456 ();
 sg13g2_decap_8 FILLER_33_1463 ();
 sg13g2_decap_8 FILLER_33_1470 ();
 sg13g2_decap_8 FILLER_33_1477 ();
 sg13g2_decap_8 FILLER_33_1484 ();
 sg13g2_decap_8 FILLER_33_1491 ();
 sg13g2_decap_8 FILLER_33_1498 ();
 sg13g2_decap_8 FILLER_33_1505 ();
 sg13g2_decap_8 FILLER_33_1512 ();
 sg13g2_decap_8 FILLER_33_1519 ();
 sg13g2_decap_8 FILLER_33_1526 ();
 sg13g2_decap_8 FILLER_33_1533 ();
 sg13g2_decap_8 FILLER_33_1540 ();
 sg13g2_decap_8 FILLER_33_1547 ();
 sg13g2_decap_8 FILLER_33_1554 ();
 sg13g2_decap_8 FILLER_33_1561 ();
 sg13g2_decap_8 FILLER_33_1568 ();
 sg13g2_decap_8 FILLER_33_1575 ();
 sg13g2_decap_8 FILLER_33_1582 ();
 sg13g2_decap_8 FILLER_33_1589 ();
 sg13g2_decap_8 FILLER_33_1596 ();
 sg13g2_decap_8 FILLER_33_1603 ();
 sg13g2_decap_8 FILLER_33_1610 ();
 sg13g2_decap_8 FILLER_33_1617 ();
 sg13g2_decap_8 FILLER_33_1624 ();
 sg13g2_decap_8 FILLER_33_1631 ();
 sg13g2_decap_8 FILLER_33_1638 ();
 sg13g2_decap_8 FILLER_33_1645 ();
 sg13g2_decap_8 FILLER_33_1652 ();
 sg13g2_decap_8 FILLER_33_1659 ();
 sg13g2_decap_8 FILLER_33_1666 ();
 sg13g2_decap_8 FILLER_33_1673 ();
 sg13g2_decap_8 FILLER_33_1680 ();
 sg13g2_decap_8 FILLER_33_1687 ();
 sg13g2_decap_8 FILLER_33_1694 ();
 sg13g2_decap_8 FILLER_33_1701 ();
 sg13g2_decap_8 FILLER_33_1708 ();
 sg13g2_decap_8 FILLER_33_1715 ();
 sg13g2_decap_8 FILLER_33_1722 ();
 sg13g2_decap_8 FILLER_33_1729 ();
 sg13g2_decap_8 FILLER_33_1736 ();
 sg13g2_decap_8 FILLER_33_1743 ();
 sg13g2_decap_8 FILLER_33_1750 ();
 sg13g2_decap_8 FILLER_33_1757 ();
 sg13g2_decap_4 FILLER_33_1764 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_decap_8 FILLER_34_91 ();
 sg13g2_decap_8 FILLER_34_98 ();
 sg13g2_decap_8 FILLER_34_105 ();
 sg13g2_decap_8 FILLER_34_112 ();
 sg13g2_decap_8 FILLER_34_119 ();
 sg13g2_decap_8 FILLER_34_126 ();
 sg13g2_decap_8 FILLER_34_133 ();
 sg13g2_decap_8 FILLER_34_140 ();
 sg13g2_decap_8 FILLER_34_147 ();
 sg13g2_decap_8 FILLER_34_154 ();
 sg13g2_fill_2 FILLER_34_161 ();
 sg13g2_fill_1 FILLER_34_163 ();
 sg13g2_decap_8 FILLER_34_177 ();
 sg13g2_decap_8 FILLER_34_184 ();
 sg13g2_decap_8 FILLER_34_191 ();
 sg13g2_decap_8 FILLER_34_198 ();
 sg13g2_fill_2 FILLER_34_205 ();
 sg13g2_fill_1 FILLER_34_207 ();
 sg13g2_fill_2 FILLER_34_229 ();
 sg13g2_fill_1 FILLER_34_266 ();
 sg13g2_fill_2 FILLER_34_316 ();
 sg13g2_fill_2 FILLER_34_342 ();
 sg13g2_fill_1 FILLER_34_344 ();
 sg13g2_fill_1 FILLER_34_350 ();
 sg13g2_decap_4 FILLER_34_377 ();
 sg13g2_fill_1 FILLER_34_381 ();
 sg13g2_decap_8 FILLER_34_408 ();
 sg13g2_decap_4 FILLER_34_415 ();
 sg13g2_fill_1 FILLER_34_419 ();
 sg13g2_fill_2 FILLER_34_466 ();
 sg13g2_fill_1 FILLER_34_468 ();
 sg13g2_fill_2 FILLER_34_478 ();
 sg13g2_fill_2 FILLER_34_552 ();
 sg13g2_fill_1 FILLER_34_554 ();
 sg13g2_fill_2 FILLER_34_602 ();
 sg13g2_fill_1 FILLER_34_618 ();
 sg13g2_fill_2 FILLER_34_634 ();
 sg13g2_fill_1 FILLER_34_682 ();
 sg13g2_decap_8 FILLER_34_722 ();
 sg13g2_fill_1 FILLER_34_729 ();
 sg13g2_decap_4 FILLER_34_765 ();
 sg13g2_fill_1 FILLER_34_795 ();
 sg13g2_fill_2 FILLER_34_808 ();
 sg13g2_fill_2 FILLER_34_826 ();
 sg13g2_fill_1 FILLER_34_828 ();
 sg13g2_fill_2 FILLER_34_838 ();
 sg13g2_decap_4 FILLER_34_893 ();
 sg13g2_fill_2 FILLER_34_903 ();
 sg13g2_fill_1 FILLER_34_905 ();
 sg13g2_fill_1 FILLER_34_944 ();
 sg13g2_fill_1 FILLER_34_954 ();
 sg13g2_fill_1 FILLER_34_959 ();
 sg13g2_fill_2 FILLER_34_1001 ();
 sg13g2_fill_1 FILLER_34_1018 ();
 sg13g2_fill_2 FILLER_34_1054 ();
 sg13g2_fill_1 FILLER_34_1056 ();
 sg13g2_fill_1 FILLER_34_1074 ();
 sg13g2_fill_1 FILLER_34_1080 ();
 sg13g2_fill_1 FILLER_34_1226 ();
 sg13g2_fill_2 FILLER_34_1241 ();
 sg13g2_fill_1 FILLER_34_1243 ();
 sg13g2_fill_1 FILLER_34_1253 ();
 sg13g2_fill_2 FILLER_34_1258 ();
 sg13g2_fill_1 FILLER_34_1278 ();
 sg13g2_fill_1 FILLER_34_1301 ();
 sg13g2_decap_8 FILLER_34_1320 ();
 sg13g2_decap_8 FILLER_34_1327 ();
 sg13g2_decap_8 FILLER_34_1334 ();
 sg13g2_decap_8 FILLER_34_1341 ();
 sg13g2_decap_8 FILLER_34_1348 ();
 sg13g2_decap_8 FILLER_34_1355 ();
 sg13g2_decap_8 FILLER_34_1362 ();
 sg13g2_decap_8 FILLER_34_1369 ();
 sg13g2_decap_8 FILLER_34_1376 ();
 sg13g2_decap_8 FILLER_34_1383 ();
 sg13g2_decap_8 FILLER_34_1390 ();
 sg13g2_decap_8 FILLER_34_1397 ();
 sg13g2_decap_8 FILLER_34_1404 ();
 sg13g2_decap_8 FILLER_34_1411 ();
 sg13g2_decap_8 FILLER_34_1418 ();
 sg13g2_decap_8 FILLER_34_1425 ();
 sg13g2_decap_8 FILLER_34_1432 ();
 sg13g2_decap_8 FILLER_34_1439 ();
 sg13g2_decap_8 FILLER_34_1446 ();
 sg13g2_decap_8 FILLER_34_1453 ();
 sg13g2_decap_8 FILLER_34_1460 ();
 sg13g2_decap_8 FILLER_34_1467 ();
 sg13g2_decap_8 FILLER_34_1474 ();
 sg13g2_decap_8 FILLER_34_1481 ();
 sg13g2_decap_8 FILLER_34_1488 ();
 sg13g2_decap_8 FILLER_34_1495 ();
 sg13g2_decap_8 FILLER_34_1502 ();
 sg13g2_decap_8 FILLER_34_1509 ();
 sg13g2_decap_8 FILLER_34_1516 ();
 sg13g2_decap_8 FILLER_34_1523 ();
 sg13g2_decap_8 FILLER_34_1530 ();
 sg13g2_decap_8 FILLER_34_1537 ();
 sg13g2_decap_8 FILLER_34_1544 ();
 sg13g2_decap_8 FILLER_34_1551 ();
 sg13g2_decap_8 FILLER_34_1558 ();
 sg13g2_decap_8 FILLER_34_1565 ();
 sg13g2_decap_8 FILLER_34_1572 ();
 sg13g2_decap_8 FILLER_34_1579 ();
 sg13g2_decap_8 FILLER_34_1586 ();
 sg13g2_decap_8 FILLER_34_1593 ();
 sg13g2_decap_8 FILLER_34_1600 ();
 sg13g2_decap_8 FILLER_34_1607 ();
 sg13g2_decap_8 FILLER_34_1614 ();
 sg13g2_decap_8 FILLER_34_1621 ();
 sg13g2_decap_8 FILLER_34_1628 ();
 sg13g2_decap_8 FILLER_34_1635 ();
 sg13g2_decap_8 FILLER_34_1642 ();
 sg13g2_decap_8 FILLER_34_1649 ();
 sg13g2_decap_8 FILLER_34_1656 ();
 sg13g2_decap_8 FILLER_34_1663 ();
 sg13g2_decap_8 FILLER_34_1670 ();
 sg13g2_decap_8 FILLER_34_1677 ();
 sg13g2_decap_8 FILLER_34_1684 ();
 sg13g2_decap_8 FILLER_34_1691 ();
 sg13g2_decap_8 FILLER_34_1698 ();
 sg13g2_decap_8 FILLER_34_1705 ();
 sg13g2_decap_8 FILLER_34_1712 ();
 sg13g2_decap_8 FILLER_34_1719 ();
 sg13g2_decap_8 FILLER_34_1726 ();
 sg13g2_decap_8 FILLER_34_1733 ();
 sg13g2_decap_8 FILLER_34_1740 ();
 sg13g2_decap_8 FILLER_34_1747 ();
 sg13g2_decap_8 FILLER_34_1754 ();
 sg13g2_decap_8 FILLER_34_1761 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_decap_8 FILLER_35_98 ();
 sg13g2_decap_8 FILLER_35_105 ();
 sg13g2_decap_8 FILLER_35_112 ();
 sg13g2_decap_8 FILLER_35_119 ();
 sg13g2_decap_8 FILLER_35_126 ();
 sg13g2_decap_8 FILLER_35_133 ();
 sg13g2_decap_8 FILLER_35_140 ();
 sg13g2_decap_8 FILLER_35_147 ();
 sg13g2_decap_8 FILLER_35_154 ();
 sg13g2_decap_8 FILLER_35_161 ();
 sg13g2_decap_8 FILLER_35_168 ();
 sg13g2_decap_8 FILLER_35_175 ();
 sg13g2_decap_8 FILLER_35_182 ();
 sg13g2_decap_8 FILLER_35_189 ();
 sg13g2_decap_8 FILLER_35_196 ();
 sg13g2_decap_8 FILLER_35_203 ();
 sg13g2_fill_1 FILLER_35_218 ();
 sg13g2_fill_2 FILLER_35_282 ();
 sg13g2_fill_1 FILLER_35_369 ();
 sg13g2_fill_2 FILLER_35_379 ();
 sg13g2_fill_1 FILLER_35_381 ();
 sg13g2_fill_2 FILLER_35_391 ();
 sg13g2_fill_2 FILLER_35_495 ();
 sg13g2_fill_1 FILLER_35_497 ();
 sg13g2_decap_4 FILLER_35_533 ();
 sg13g2_fill_1 FILLER_35_572 ();
 sg13g2_fill_2 FILLER_35_582 ();
 sg13g2_fill_2 FILLER_35_610 ();
 sg13g2_fill_1 FILLER_35_628 ();
 sg13g2_fill_1 FILLER_35_654 ();
 sg13g2_fill_2 FILLER_35_675 ();
 sg13g2_fill_1 FILLER_35_709 ();
 sg13g2_fill_1 FILLER_35_714 ();
 sg13g2_decap_8 FILLER_35_720 ();
 sg13g2_fill_2 FILLER_35_727 ();
 sg13g2_fill_1 FILLER_35_729 ();
 sg13g2_decap_8 FILLER_35_782 ();
 sg13g2_decap_8 FILLER_35_789 ();
 sg13g2_fill_2 FILLER_35_980 ();
 sg13g2_decap_8 FILLER_35_987 ();
 sg13g2_decap_4 FILLER_35_994 ();
 sg13g2_fill_2 FILLER_35_1018 ();
 sg13g2_fill_2 FILLER_35_1034 ();
 sg13g2_fill_1 FILLER_35_1044 ();
 sg13g2_fill_2 FILLER_35_1053 ();
 sg13g2_fill_2 FILLER_35_1126 ();
 sg13g2_decap_4 FILLER_35_1201 ();
 sg13g2_fill_1 FILLER_35_1205 ();
 sg13g2_fill_2 FILLER_35_1254 ();
 sg13g2_fill_1 FILLER_35_1286 ();
 sg13g2_decap_8 FILLER_35_1313 ();
 sg13g2_decap_8 FILLER_35_1320 ();
 sg13g2_decap_8 FILLER_35_1327 ();
 sg13g2_decap_8 FILLER_35_1334 ();
 sg13g2_decap_8 FILLER_35_1341 ();
 sg13g2_decap_8 FILLER_35_1348 ();
 sg13g2_decap_8 FILLER_35_1355 ();
 sg13g2_decap_8 FILLER_35_1362 ();
 sg13g2_decap_8 FILLER_35_1369 ();
 sg13g2_decap_8 FILLER_35_1376 ();
 sg13g2_decap_8 FILLER_35_1383 ();
 sg13g2_decap_8 FILLER_35_1390 ();
 sg13g2_decap_8 FILLER_35_1397 ();
 sg13g2_decap_8 FILLER_35_1404 ();
 sg13g2_decap_8 FILLER_35_1411 ();
 sg13g2_decap_8 FILLER_35_1418 ();
 sg13g2_decap_8 FILLER_35_1425 ();
 sg13g2_decap_8 FILLER_35_1432 ();
 sg13g2_decap_8 FILLER_35_1439 ();
 sg13g2_decap_8 FILLER_35_1446 ();
 sg13g2_decap_8 FILLER_35_1453 ();
 sg13g2_decap_8 FILLER_35_1460 ();
 sg13g2_decap_8 FILLER_35_1467 ();
 sg13g2_decap_8 FILLER_35_1474 ();
 sg13g2_decap_8 FILLER_35_1481 ();
 sg13g2_decap_8 FILLER_35_1488 ();
 sg13g2_decap_8 FILLER_35_1495 ();
 sg13g2_decap_8 FILLER_35_1502 ();
 sg13g2_decap_8 FILLER_35_1509 ();
 sg13g2_decap_8 FILLER_35_1516 ();
 sg13g2_decap_8 FILLER_35_1523 ();
 sg13g2_decap_8 FILLER_35_1530 ();
 sg13g2_decap_8 FILLER_35_1537 ();
 sg13g2_decap_8 FILLER_35_1544 ();
 sg13g2_decap_8 FILLER_35_1551 ();
 sg13g2_decap_8 FILLER_35_1558 ();
 sg13g2_decap_8 FILLER_35_1565 ();
 sg13g2_decap_8 FILLER_35_1572 ();
 sg13g2_decap_8 FILLER_35_1579 ();
 sg13g2_decap_8 FILLER_35_1586 ();
 sg13g2_decap_8 FILLER_35_1593 ();
 sg13g2_decap_8 FILLER_35_1600 ();
 sg13g2_decap_8 FILLER_35_1607 ();
 sg13g2_decap_8 FILLER_35_1614 ();
 sg13g2_decap_8 FILLER_35_1621 ();
 sg13g2_decap_8 FILLER_35_1628 ();
 sg13g2_decap_8 FILLER_35_1635 ();
 sg13g2_decap_8 FILLER_35_1642 ();
 sg13g2_decap_8 FILLER_35_1649 ();
 sg13g2_decap_8 FILLER_35_1656 ();
 sg13g2_decap_8 FILLER_35_1663 ();
 sg13g2_decap_8 FILLER_35_1670 ();
 sg13g2_decap_8 FILLER_35_1677 ();
 sg13g2_decap_8 FILLER_35_1684 ();
 sg13g2_decap_8 FILLER_35_1691 ();
 sg13g2_decap_8 FILLER_35_1698 ();
 sg13g2_decap_8 FILLER_35_1705 ();
 sg13g2_decap_8 FILLER_35_1712 ();
 sg13g2_decap_8 FILLER_35_1719 ();
 sg13g2_decap_8 FILLER_35_1726 ();
 sg13g2_decap_8 FILLER_35_1733 ();
 sg13g2_decap_8 FILLER_35_1740 ();
 sg13g2_decap_8 FILLER_35_1747 ();
 sg13g2_decap_8 FILLER_35_1754 ();
 sg13g2_decap_8 FILLER_35_1761 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_decap_8 FILLER_36_112 ();
 sg13g2_decap_8 FILLER_36_119 ();
 sg13g2_decap_8 FILLER_36_126 ();
 sg13g2_decap_8 FILLER_36_133 ();
 sg13g2_decap_8 FILLER_36_140 ();
 sg13g2_decap_8 FILLER_36_147 ();
 sg13g2_decap_8 FILLER_36_154 ();
 sg13g2_decap_8 FILLER_36_161 ();
 sg13g2_decap_8 FILLER_36_168 ();
 sg13g2_decap_8 FILLER_36_175 ();
 sg13g2_decap_8 FILLER_36_182 ();
 sg13g2_decap_8 FILLER_36_189 ();
 sg13g2_decap_8 FILLER_36_196 ();
 sg13g2_decap_8 FILLER_36_203 ();
 sg13g2_decap_4 FILLER_36_210 ();
 sg13g2_fill_1 FILLER_36_235 ();
 sg13g2_fill_1 FILLER_36_302 ();
 sg13g2_decap_8 FILLER_36_307 ();
 sg13g2_fill_2 FILLER_36_314 ();
 sg13g2_fill_1 FILLER_36_316 ();
 sg13g2_decap_8 FILLER_36_335 ();
 sg13g2_decap_8 FILLER_36_342 ();
 sg13g2_fill_1 FILLER_36_349 ();
 sg13g2_decap_8 FILLER_36_409 ();
 sg13g2_fill_1 FILLER_36_416 ();
 sg13g2_fill_2 FILLER_36_443 ();
 sg13g2_decap_8 FILLER_36_450 ();
 sg13g2_decap_8 FILLER_36_457 ();
 sg13g2_decap_4 FILLER_36_464 ();
 sg13g2_fill_2 FILLER_36_468 ();
 sg13g2_fill_1 FILLER_36_478 ();
 sg13g2_fill_1 FILLER_36_487 ();
 sg13g2_fill_2 FILLER_36_498 ();
 sg13g2_fill_1 FILLER_36_500 ();
 sg13g2_fill_2 FILLER_36_513 ();
 sg13g2_fill_1 FILLER_36_515 ();
 sg13g2_decap_4 FILLER_36_546 ();
 sg13g2_fill_1 FILLER_36_576 ();
 sg13g2_fill_1 FILLER_36_607 ();
 sg13g2_fill_2 FILLER_36_612 ();
 sg13g2_decap_8 FILLER_36_625 ();
 sg13g2_fill_2 FILLER_36_654 ();
 sg13g2_fill_1 FILLER_36_656 ();
 sg13g2_fill_2 FILLER_36_673 ();
 sg13g2_fill_2 FILLER_36_685 ();
 sg13g2_decap_8 FILLER_36_700 ();
 sg13g2_fill_1 FILLER_36_707 ();
 sg13g2_fill_2 FILLER_36_732 ();
 sg13g2_fill_1 FILLER_36_734 ();
 sg13g2_fill_1 FILLER_36_748 ();
 sg13g2_decap_4 FILLER_36_758 ();
 sg13g2_fill_2 FILLER_36_762 ();
 sg13g2_decap_4 FILLER_36_839 ();
 sg13g2_fill_1 FILLER_36_848 ();
 sg13g2_fill_1 FILLER_36_883 ();
 sg13g2_decap_4 FILLER_36_892 ();
 sg13g2_fill_2 FILLER_36_930 ();
 sg13g2_decap_8 FILLER_36_993 ();
 sg13g2_fill_2 FILLER_36_1031 ();
 sg13g2_fill_1 FILLER_36_1033 ();
 sg13g2_fill_2 FILLER_36_1100 ();
 sg13g2_fill_2 FILLER_36_1231 ();
 sg13g2_decap_8 FILLER_36_1298 ();
 sg13g2_decap_8 FILLER_36_1305 ();
 sg13g2_decap_8 FILLER_36_1312 ();
 sg13g2_decap_8 FILLER_36_1319 ();
 sg13g2_decap_8 FILLER_36_1326 ();
 sg13g2_decap_8 FILLER_36_1333 ();
 sg13g2_decap_8 FILLER_36_1340 ();
 sg13g2_decap_8 FILLER_36_1347 ();
 sg13g2_decap_8 FILLER_36_1354 ();
 sg13g2_decap_8 FILLER_36_1361 ();
 sg13g2_decap_8 FILLER_36_1368 ();
 sg13g2_decap_8 FILLER_36_1375 ();
 sg13g2_decap_8 FILLER_36_1382 ();
 sg13g2_decap_8 FILLER_36_1389 ();
 sg13g2_decap_8 FILLER_36_1396 ();
 sg13g2_decap_8 FILLER_36_1403 ();
 sg13g2_decap_8 FILLER_36_1410 ();
 sg13g2_decap_8 FILLER_36_1417 ();
 sg13g2_decap_8 FILLER_36_1424 ();
 sg13g2_decap_8 FILLER_36_1431 ();
 sg13g2_decap_8 FILLER_36_1438 ();
 sg13g2_decap_8 FILLER_36_1445 ();
 sg13g2_decap_8 FILLER_36_1452 ();
 sg13g2_decap_8 FILLER_36_1459 ();
 sg13g2_decap_8 FILLER_36_1466 ();
 sg13g2_decap_8 FILLER_36_1473 ();
 sg13g2_decap_8 FILLER_36_1480 ();
 sg13g2_decap_8 FILLER_36_1487 ();
 sg13g2_decap_8 FILLER_36_1494 ();
 sg13g2_decap_8 FILLER_36_1501 ();
 sg13g2_decap_8 FILLER_36_1508 ();
 sg13g2_decap_8 FILLER_36_1515 ();
 sg13g2_decap_8 FILLER_36_1522 ();
 sg13g2_decap_8 FILLER_36_1529 ();
 sg13g2_decap_8 FILLER_36_1536 ();
 sg13g2_decap_8 FILLER_36_1543 ();
 sg13g2_decap_8 FILLER_36_1550 ();
 sg13g2_decap_8 FILLER_36_1557 ();
 sg13g2_decap_8 FILLER_36_1564 ();
 sg13g2_decap_8 FILLER_36_1571 ();
 sg13g2_decap_8 FILLER_36_1578 ();
 sg13g2_decap_8 FILLER_36_1585 ();
 sg13g2_decap_8 FILLER_36_1592 ();
 sg13g2_decap_8 FILLER_36_1599 ();
 sg13g2_decap_8 FILLER_36_1606 ();
 sg13g2_decap_8 FILLER_36_1613 ();
 sg13g2_decap_8 FILLER_36_1620 ();
 sg13g2_decap_8 FILLER_36_1627 ();
 sg13g2_decap_8 FILLER_36_1634 ();
 sg13g2_decap_8 FILLER_36_1641 ();
 sg13g2_decap_8 FILLER_36_1648 ();
 sg13g2_decap_8 FILLER_36_1655 ();
 sg13g2_decap_8 FILLER_36_1662 ();
 sg13g2_decap_8 FILLER_36_1669 ();
 sg13g2_decap_8 FILLER_36_1676 ();
 sg13g2_decap_8 FILLER_36_1683 ();
 sg13g2_decap_8 FILLER_36_1690 ();
 sg13g2_decap_8 FILLER_36_1697 ();
 sg13g2_decap_8 FILLER_36_1704 ();
 sg13g2_decap_8 FILLER_36_1711 ();
 sg13g2_decap_8 FILLER_36_1718 ();
 sg13g2_decap_8 FILLER_36_1725 ();
 sg13g2_decap_8 FILLER_36_1732 ();
 sg13g2_decap_8 FILLER_36_1739 ();
 sg13g2_decap_8 FILLER_36_1746 ();
 sg13g2_decap_8 FILLER_36_1753 ();
 sg13g2_decap_8 FILLER_36_1760 ();
 sg13g2_fill_1 FILLER_36_1767 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_8 FILLER_37_112 ();
 sg13g2_decap_8 FILLER_37_119 ();
 sg13g2_decap_8 FILLER_37_126 ();
 sg13g2_decap_8 FILLER_37_133 ();
 sg13g2_decap_8 FILLER_37_140 ();
 sg13g2_decap_8 FILLER_37_147 ();
 sg13g2_decap_8 FILLER_37_154 ();
 sg13g2_decap_8 FILLER_37_161 ();
 sg13g2_decap_8 FILLER_37_168 ();
 sg13g2_decap_8 FILLER_37_175 ();
 sg13g2_decap_8 FILLER_37_182 ();
 sg13g2_decap_8 FILLER_37_189 ();
 sg13g2_fill_2 FILLER_37_199 ();
 sg13g2_fill_1 FILLER_37_201 ();
 sg13g2_fill_2 FILLER_37_228 ();
 sg13g2_fill_1 FILLER_37_230 ();
 sg13g2_fill_1 FILLER_37_258 ();
 sg13g2_fill_1 FILLER_37_273 ();
 sg13g2_fill_1 FILLER_37_283 ();
 sg13g2_decap_8 FILLER_37_292 ();
 sg13g2_decap_4 FILLER_37_299 ();
 sg13g2_fill_2 FILLER_37_303 ();
 sg13g2_fill_2 FILLER_37_321 ();
 sg13g2_fill_1 FILLER_37_323 ();
 sg13g2_decap_4 FILLER_37_340 ();
 sg13g2_fill_1 FILLER_37_344 ();
 sg13g2_fill_1 FILLER_37_358 ();
 sg13g2_decap_8 FILLER_37_380 ();
 sg13g2_fill_1 FILLER_37_387 ();
 sg13g2_decap_8 FILLER_37_412 ();
 sg13g2_decap_8 FILLER_37_426 ();
 sg13g2_fill_2 FILLER_37_433 ();
 sg13g2_fill_1 FILLER_37_466 ();
 sg13g2_fill_1 FILLER_37_477 ();
 sg13g2_decap_4 FILLER_37_483 ();
 sg13g2_fill_1 FILLER_37_487 ();
 sg13g2_fill_1 FILLER_37_507 ();
 sg13g2_fill_1 FILLER_37_541 ();
 sg13g2_fill_2 FILLER_37_547 ();
 sg13g2_fill_1 FILLER_37_549 ();
 sg13g2_decap_4 FILLER_37_559 ();
 sg13g2_fill_2 FILLER_37_567 ();
 sg13g2_decap_4 FILLER_37_573 ();
 sg13g2_fill_2 FILLER_37_577 ();
 sg13g2_decap_4 FILLER_37_589 ();
 sg13g2_fill_2 FILLER_37_593 ();
 sg13g2_fill_2 FILLER_37_605 ();
 sg13g2_fill_1 FILLER_37_607 ();
 sg13g2_decap_8 FILLER_37_694 ();
 sg13g2_decap_8 FILLER_37_701 ();
 sg13g2_decap_4 FILLER_37_708 ();
 sg13g2_fill_1 FILLER_37_712 ();
 sg13g2_decap_8 FILLER_37_737 ();
 sg13g2_decap_4 FILLER_37_744 ();
 sg13g2_fill_1 FILLER_37_748 ();
 sg13g2_fill_2 FILLER_37_762 ();
 sg13g2_fill_1 FILLER_37_764 ();
 sg13g2_fill_1 FILLER_37_776 ();
 sg13g2_fill_2 FILLER_37_797 ();
 sg13g2_fill_1 FILLER_37_799 ();
 sg13g2_decap_4 FILLER_37_835 ();
 sg13g2_decap_4 FILLER_37_899 ();
 sg13g2_decap_8 FILLER_37_911 ();
 sg13g2_fill_1 FILLER_37_921 ();
 sg13g2_fill_2 FILLER_37_926 ();
 sg13g2_fill_1 FILLER_37_928 ();
 sg13g2_decap_8 FILLER_37_1007 ();
 sg13g2_decap_8 FILLER_37_1014 ();
 sg13g2_fill_1 FILLER_37_1021 ();
 sg13g2_fill_1 FILLER_37_1071 ();
 sg13g2_fill_2 FILLER_37_1152 ();
 sg13g2_fill_1 FILLER_37_1154 ();
 sg13g2_fill_2 FILLER_37_1198 ();
 sg13g2_fill_1 FILLER_37_1200 ();
 sg13g2_decap_8 FILLER_37_1262 ();
 sg13g2_decap_8 FILLER_37_1269 ();
 sg13g2_decap_4 FILLER_37_1276 ();
 sg13g2_fill_1 FILLER_37_1284 ();
 sg13g2_fill_2 FILLER_37_1298 ();
 sg13g2_decap_8 FILLER_37_1309 ();
 sg13g2_decap_8 FILLER_37_1316 ();
 sg13g2_decap_8 FILLER_37_1323 ();
 sg13g2_decap_8 FILLER_37_1330 ();
 sg13g2_decap_8 FILLER_37_1337 ();
 sg13g2_decap_8 FILLER_37_1344 ();
 sg13g2_decap_8 FILLER_37_1351 ();
 sg13g2_decap_8 FILLER_37_1358 ();
 sg13g2_decap_8 FILLER_37_1365 ();
 sg13g2_decap_8 FILLER_37_1372 ();
 sg13g2_decap_8 FILLER_37_1379 ();
 sg13g2_decap_8 FILLER_37_1386 ();
 sg13g2_decap_8 FILLER_37_1393 ();
 sg13g2_decap_8 FILLER_37_1400 ();
 sg13g2_decap_8 FILLER_37_1407 ();
 sg13g2_decap_8 FILLER_37_1414 ();
 sg13g2_decap_8 FILLER_37_1421 ();
 sg13g2_decap_8 FILLER_37_1428 ();
 sg13g2_decap_8 FILLER_37_1435 ();
 sg13g2_decap_8 FILLER_37_1442 ();
 sg13g2_decap_8 FILLER_37_1449 ();
 sg13g2_decap_8 FILLER_37_1456 ();
 sg13g2_decap_8 FILLER_37_1463 ();
 sg13g2_decap_8 FILLER_37_1470 ();
 sg13g2_decap_8 FILLER_37_1477 ();
 sg13g2_decap_8 FILLER_37_1484 ();
 sg13g2_decap_8 FILLER_37_1491 ();
 sg13g2_decap_8 FILLER_37_1498 ();
 sg13g2_decap_8 FILLER_37_1505 ();
 sg13g2_decap_8 FILLER_37_1512 ();
 sg13g2_decap_8 FILLER_37_1519 ();
 sg13g2_decap_8 FILLER_37_1526 ();
 sg13g2_decap_8 FILLER_37_1533 ();
 sg13g2_decap_8 FILLER_37_1540 ();
 sg13g2_decap_8 FILLER_37_1547 ();
 sg13g2_decap_8 FILLER_37_1554 ();
 sg13g2_decap_8 FILLER_37_1561 ();
 sg13g2_decap_8 FILLER_37_1568 ();
 sg13g2_decap_8 FILLER_37_1575 ();
 sg13g2_decap_8 FILLER_37_1582 ();
 sg13g2_decap_8 FILLER_37_1589 ();
 sg13g2_decap_8 FILLER_37_1596 ();
 sg13g2_decap_8 FILLER_37_1603 ();
 sg13g2_decap_8 FILLER_37_1610 ();
 sg13g2_decap_8 FILLER_37_1617 ();
 sg13g2_decap_8 FILLER_37_1624 ();
 sg13g2_decap_8 FILLER_37_1631 ();
 sg13g2_decap_8 FILLER_37_1638 ();
 sg13g2_decap_8 FILLER_37_1645 ();
 sg13g2_decap_8 FILLER_37_1652 ();
 sg13g2_decap_8 FILLER_37_1659 ();
 sg13g2_decap_8 FILLER_37_1666 ();
 sg13g2_decap_8 FILLER_37_1673 ();
 sg13g2_decap_8 FILLER_37_1680 ();
 sg13g2_decap_8 FILLER_37_1687 ();
 sg13g2_decap_8 FILLER_37_1694 ();
 sg13g2_decap_8 FILLER_37_1701 ();
 sg13g2_decap_8 FILLER_37_1708 ();
 sg13g2_decap_8 FILLER_37_1715 ();
 sg13g2_decap_8 FILLER_37_1722 ();
 sg13g2_decap_8 FILLER_37_1729 ();
 sg13g2_decap_8 FILLER_37_1736 ();
 sg13g2_decap_8 FILLER_37_1743 ();
 sg13g2_decap_8 FILLER_37_1750 ();
 sg13g2_decap_8 FILLER_37_1757 ();
 sg13g2_decap_4 FILLER_37_1764 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_8 FILLER_38_56 ();
 sg13g2_decap_8 FILLER_38_63 ();
 sg13g2_decap_8 FILLER_38_70 ();
 sg13g2_decap_8 FILLER_38_77 ();
 sg13g2_decap_8 FILLER_38_84 ();
 sg13g2_decap_8 FILLER_38_91 ();
 sg13g2_decap_8 FILLER_38_98 ();
 sg13g2_decap_8 FILLER_38_105 ();
 sg13g2_decap_8 FILLER_38_112 ();
 sg13g2_decap_8 FILLER_38_119 ();
 sg13g2_decap_8 FILLER_38_126 ();
 sg13g2_decap_8 FILLER_38_133 ();
 sg13g2_decap_8 FILLER_38_140 ();
 sg13g2_decap_8 FILLER_38_147 ();
 sg13g2_decap_8 FILLER_38_154 ();
 sg13g2_decap_8 FILLER_38_161 ();
 sg13g2_decap_8 FILLER_38_168 ();
 sg13g2_fill_2 FILLER_38_175 ();
 sg13g2_decap_8 FILLER_38_181 ();
 sg13g2_fill_2 FILLER_38_197 ();
 sg13g2_fill_1 FILLER_38_228 ();
 sg13g2_fill_1 FILLER_38_247 ();
 sg13g2_decap_4 FILLER_38_291 ();
 sg13g2_fill_2 FILLER_38_295 ();
 sg13g2_fill_2 FILLER_38_313 ();
 sg13g2_fill_2 FILLER_38_334 ();
 sg13g2_fill_1 FILLER_38_336 ();
 sg13g2_fill_2 FILLER_38_345 ();
 sg13g2_fill_1 FILLER_38_347 ();
 sg13g2_fill_1 FILLER_38_361 ();
 sg13g2_decap_8 FILLER_38_374 ();
 sg13g2_fill_1 FILLER_38_381 ();
 sg13g2_fill_1 FILLER_38_407 ();
 sg13g2_decap_4 FILLER_38_433 ();
 sg13g2_decap_4 FILLER_38_450 ();
 sg13g2_fill_1 FILLER_38_454 ();
 sg13g2_fill_2 FILLER_38_462 ();
 sg13g2_fill_1 FILLER_38_477 ();
 sg13g2_decap_4 FILLER_38_508 ();
 sg13g2_fill_1 FILLER_38_528 ();
 sg13g2_decap_8 FILLER_38_547 ();
 sg13g2_decap_4 FILLER_38_554 ();
 sg13g2_decap_8 FILLER_38_566 ();
 sg13g2_fill_2 FILLER_38_573 ();
 sg13g2_fill_1 FILLER_38_575 ();
 sg13g2_fill_2 FILLER_38_683 ();
 sg13g2_decap_8 FILLER_38_711 ();
 sg13g2_decap_4 FILLER_38_734 ();
 sg13g2_fill_2 FILLER_38_738 ();
 sg13g2_fill_2 FILLER_38_769 ();
 sg13g2_fill_1 FILLER_38_771 ();
 sg13g2_fill_2 FILLER_38_840 ();
 sg13g2_fill_1 FILLER_38_842 ();
 sg13g2_decap_8 FILLER_38_847 ();
 sg13g2_decap_8 FILLER_38_854 ();
 sg13g2_decap_8 FILLER_38_861 ();
 sg13g2_decap_8 FILLER_38_868 ();
 sg13g2_decap_4 FILLER_38_875 ();
 sg13g2_decap_8 FILLER_38_884 ();
 sg13g2_decap_8 FILLER_38_891 ();
 sg13g2_fill_2 FILLER_38_898 ();
 sg13g2_fill_1 FILLER_38_900 ();
 sg13g2_fill_2 FILLER_38_919 ();
 sg13g2_fill_1 FILLER_38_955 ();
 sg13g2_fill_2 FILLER_38_1061 ();
 sg13g2_fill_1 FILLER_38_1072 ();
 sg13g2_fill_2 FILLER_38_1129 ();
 sg13g2_fill_1 FILLER_38_1131 ();
 sg13g2_decap_4 FILLER_38_1140 ();
 sg13g2_fill_2 FILLER_38_1144 ();
 sg13g2_fill_2 FILLER_38_1185 ();
 sg13g2_fill_1 FILLER_38_1187 ();
 sg13g2_decap_8 FILLER_38_1197 ();
 sg13g2_fill_2 FILLER_38_1240 ();
 sg13g2_decap_8 FILLER_38_1251 ();
 sg13g2_decap_8 FILLER_38_1258 ();
 sg13g2_decap_8 FILLER_38_1265 ();
 sg13g2_decap_8 FILLER_38_1272 ();
 sg13g2_decap_8 FILLER_38_1279 ();
 sg13g2_decap_8 FILLER_38_1286 ();
 sg13g2_decap_8 FILLER_38_1293 ();
 sg13g2_decap_8 FILLER_38_1300 ();
 sg13g2_decap_8 FILLER_38_1307 ();
 sg13g2_decap_8 FILLER_38_1314 ();
 sg13g2_decap_8 FILLER_38_1321 ();
 sg13g2_decap_8 FILLER_38_1328 ();
 sg13g2_decap_8 FILLER_38_1335 ();
 sg13g2_decap_8 FILLER_38_1342 ();
 sg13g2_decap_8 FILLER_38_1349 ();
 sg13g2_decap_8 FILLER_38_1356 ();
 sg13g2_decap_8 FILLER_38_1363 ();
 sg13g2_decap_8 FILLER_38_1370 ();
 sg13g2_decap_8 FILLER_38_1377 ();
 sg13g2_decap_8 FILLER_38_1384 ();
 sg13g2_decap_8 FILLER_38_1391 ();
 sg13g2_decap_8 FILLER_38_1398 ();
 sg13g2_decap_8 FILLER_38_1405 ();
 sg13g2_decap_8 FILLER_38_1412 ();
 sg13g2_decap_8 FILLER_38_1419 ();
 sg13g2_decap_8 FILLER_38_1426 ();
 sg13g2_decap_8 FILLER_38_1433 ();
 sg13g2_decap_8 FILLER_38_1440 ();
 sg13g2_decap_8 FILLER_38_1447 ();
 sg13g2_decap_8 FILLER_38_1454 ();
 sg13g2_decap_8 FILLER_38_1461 ();
 sg13g2_decap_8 FILLER_38_1468 ();
 sg13g2_decap_8 FILLER_38_1475 ();
 sg13g2_decap_8 FILLER_38_1482 ();
 sg13g2_decap_8 FILLER_38_1489 ();
 sg13g2_decap_8 FILLER_38_1496 ();
 sg13g2_decap_8 FILLER_38_1503 ();
 sg13g2_decap_8 FILLER_38_1510 ();
 sg13g2_decap_8 FILLER_38_1517 ();
 sg13g2_decap_8 FILLER_38_1524 ();
 sg13g2_decap_8 FILLER_38_1531 ();
 sg13g2_decap_8 FILLER_38_1538 ();
 sg13g2_decap_8 FILLER_38_1545 ();
 sg13g2_decap_8 FILLER_38_1552 ();
 sg13g2_decap_8 FILLER_38_1559 ();
 sg13g2_decap_8 FILLER_38_1566 ();
 sg13g2_decap_8 FILLER_38_1573 ();
 sg13g2_decap_8 FILLER_38_1580 ();
 sg13g2_decap_8 FILLER_38_1587 ();
 sg13g2_decap_8 FILLER_38_1594 ();
 sg13g2_decap_8 FILLER_38_1601 ();
 sg13g2_decap_8 FILLER_38_1608 ();
 sg13g2_decap_8 FILLER_38_1615 ();
 sg13g2_decap_8 FILLER_38_1622 ();
 sg13g2_decap_8 FILLER_38_1629 ();
 sg13g2_decap_8 FILLER_38_1636 ();
 sg13g2_decap_8 FILLER_38_1643 ();
 sg13g2_decap_8 FILLER_38_1650 ();
 sg13g2_decap_8 FILLER_38_1657 ();
 sg13g2_decap_8 FILLER_38_1664 ();
 sg13g2_decap_8 FILLER_38_1671 ();
 sg13g2_decap_8 FILLER_38_1678 ();
 sg13g2_decap_8 FILLER_38_1685 ();
 sg13g2_decap_8 FILLER_38_1692 ();
 sg13g2_decap_8 FILLER_38_1699 ();
 sg13g2_decap_8 FILLER_38_1706 ();
 sg13g2_decap_8 FILLER_38_1713 ();
 sg13g2_decap_8 FILLER_38_1720 ();
 sg13g2_decap_8 FILLER_38_1727 ();
 sg13g2_decap_8 FILLER_38_1734 ();
 sg13g2_decap_8 FILLER_38_1741 ();
 sg13g2_decap_8 FILLER_38_1748 ();
 sg13g2_decap_8 FILLER_38_1755 ();
 sg13g2_decap_4 FILLER_38_1762 ();
 sg13g2_fill_2 FILLER_38_1766 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_14 ();
 sg13g2_decap_8 FILLER_39_21 ();
 sg13g2_decap_8 FILLER_39_28 ();
 sg13g2_decap_8 FILLER_39_35 ();
 sg13g2_decap_8 FILLER_39_42 ();
 sg13g2_decap_8 FILLER_39_49 ();
 sg13g2_decap_8 FILLER_39_56 ();
 sg13g2_decap_8 FILLER_39_63 ();
 sg13g2_decap_8 FILLER_39_70 ();
 sg13g2_decap_8 FILLER_39_77 ();
 sg13g2_decap_8 FILLER_39_84 ();
 sg13g2_decap_8 FILLER_39_91 ();
 sg13g2_decap_8 FILLER_39_98 ();
 sg13g2_decap_8 FILLER_39_105 ();
 sg13g2_decap_8 FILLER_39_112 ();
 sg13g2_decap_8 FILLER_39_119 ();
 sg13g2_decap_8 FILLER_39_126 ();
 sg13g2_decap_8 FILLER_39_133 ();
 sg13g2_decap_8 FILLER_39_140 ();
 sg13g2_decap_8 FILLER_39_147 ();
 sg13g2_decap_8 FILLER_39_154 ();
 sg13g2_decap_8 FILLER_39_161 ();
 sg13g2_fill_2 FILLER_39_168 ();
 sg13g2_fill_1 FILLER_39_170 ();
 sg13g2_fill_2 FILLER_39_197 ();
 sg13g2_fill_1 FILLER_39_241 ();
 sg13g2_decap_8 FILLER_39_285 ();
 sg13g2_decap_8 FILLER_39_292 ();
 sg13g2_decap_4 FILLER_39_299 ();
 sg13g2_fill_1 FILLER_39_303 ();
 sg13g2_decap_4 FILLER_39_331 ();
 sg13g2_fill_2 FILLER_39_335 ();
 sg13g2_decap_8 FILLER_39_342 ();
 sg13g2_fill_2 FILLER_39_349 ();
 sg13g2_fill_1 FILLER_39_351 ();
 sg13g2_fill_1 FILLER_39_357 ();
 sg13g2_decap_8 FILLER_39_371 ();
 sg13g2_decap_4 FILLER_39_378 ();
 sg13g2_fill_1 FILLER_39_382 ();
 sg13g2_decap_8 FILLER_39_404 ();
 sg13g2_fill_2 FILLER_39_411 ();
 sg13g2_fill_1 FILLER_39_413 ();
 sg13g2_fill_2 FILLER_39_434 ();
 sg13g2_fill_2 FILLER_39_446 ();
 sg13g2_fill_1 FILLER_39_448 ();
 sg13g2_decap_8 FILLER_39_469 ();
 sg13g2_decap_4 FILLER_39_476 ();
 sg13g2_fill_1 FILLER_39_480 ();
 sg13g2_fill_1 FILLER_39_497 ();
 sg13g2_decap_4 FILLER_39_502 ();
 sg13g2_decap_4 FILLER_39_526 ();
 sg13g2_fill_1 FILLER_39_546 ();
 sg13g2_fill_2 FILLER_39_555 ();
 sg13g2_fill_1 FILLER_39_557 ();
 sg13g2_fill_2 FILLER_39_563 ();
 sg13g2_fill_1 FILLER_39_565 ();
 sg13g2_fill_1 FILLER_39_578 ();
 sg13g2_decap_8 FILLER_39_584 ();
 sg13g2_fill_2 FILLER_39_591 ();
 sg13g2_fill_2 FILLER_39_606 ();
 sg13g2_fill_1 FILLER_39_608 ();
 sg13g2_fill_1 FILLER_39_613 ();
 sg13g2_fill_2 FILLER_39_619 ();
 sg13g2_fill_1 FILLER_39_621 ();
 sg13g2_fill_2 FILLER_39_625 ();
 sg13g2_fill_1 FILLER_39_635 ();
 sg13g2_fill_2 FILLER_39_654 ();
 sg13g2_fill_1 FILLER_39_663 ();
 sg13g2_fill_2 FILLER_39_671 ();
 sg13g2_decap_8 FILLER_39_677 ();
 sg13g2_fill_2 FILLER_39_684 ();
 sg13g2_fill_1 FILLER_39_686 ();
 sg13g2_fill_2 FILLER_39_692 ();
 sg13g2_decap_8 FILLER_39_735 ();
 sg13g2_decap_4 FILLER_39_742 ();
 sg13g2_fill_2 FILLER_39_772 ();
 sg13g2_fill_1 FILLER_39_774 ();
 sg13g2_fill_1 FILLER_39_809 ();
 sg13g2_decap_8 FILLER_39_845 ();
 sg13g2_decap_8 FILLER_39_852 ();
 sg13g2_decap_8 FILLER_39_859 ();
 sg13g2_decap_8 FILLER_39_866 ();
 sg13g2_decap_8 FILLER_39_873 ();
 sg13g2_decap_8 FILLER_39_880 ();
 sg13g2_fill_2 FILLER_39_948 ();
 sg13g2_fill_2 FILLER_39_966 ();
 sg13g2_fill_1 FILLER_39_991 ();
 sg13g2_decap_8 FILLER_39_1001 ();
 sg13g2_decap_4 FILLER_39_1008 ();
 sg13g2_fill_1 FILLER_39_1012 ();
 sg13g2_decap_8 FILLER_39_1016 ();
 sg13g2_decap_8 FILLER_39_1023 ();
 sg13g2_fill_1 FILLER_39_1030 ();
 sg13g2_fill_2 FILLER_39_1069 ();
 sg13g2_decap_8 FILLER_39_1123 ();
 sg13g2_decap_8 FILLER_39_1130 ();
 sg13g2_decap_8 FILLER_39_1137 ();
 sg13g2_decap_4 FILLER_39_1144 ();
 sg13g2_fill_2 FILLER_39_1148 ();
 sg13g2_decap_8 FILLER_39_1172 ();
 sg13g2_decap_8 FILLER_39_1179 ();
 sg13g2_decap_8 FILLER_39_1186 ();
 sg13g2_fill_2 FILLER_39_1193 ();
 sg13g2_fill_1 FILLER_39_1195 ();
 sg13g2_decap_8 FILLER_39_1204 ();
 sg13g2_fill_1 FILLER_39_1211 ();
 sg13g2_decap_8 FILLER_39_1216 ();
 sg13g2_decap_8 FILLER_39_1223 ();
 sg13g2_decap_8 FILLER_39_1230 ();
 sg13g2_decap_8 FILLER_39_1237 ();
 sg13g2_decap_8 FILLER_39_1244 ();
 sg13g2_decap_8 FILLER_39_1251 ();
 sg13g2_decap_8 FILLER_39_1258 ();
 sg13g2_decap_8 FILLER_39_1265 ();
 sg13g2_decap_8 FILLER_39_1272 ();
 sg13g2_decap_8 FILLER_39_1279 ();
 sg13g2_decap_8 FILLER_39_1286 ();
 sg13g2_decap_8 FILLER_39_1293 ();
 sg13g2_decap_8 FILLER_39_1300 ();
 sg13g2_decap_8 FILLER_39_1307 ();
 sg13g2_decap_8 FILLER_39_1314 ();
 sg13g2_decap_8 FILLER_39_1321 ();
 sg13g2_decap_8 FILLER_39_1328 ();
 sg13g2_decap_8 FILLER_39_1335 ();
 sg13g2_decap_8 FILLER_39_1342 ();
 sg13g2_decap_8 FILLER_39_1349 ();
 sg13g2_decap_8 FILLER_39_1356 ();
 sg13g2_decap_8 FILLER_39_1363 ();
 sg13g2_decap_8 FILLER_39_1370 ();
 sg13g2_decap_8 FILLER_39_1377 ();
 sg13g2_decap_8 FILLER_39_1384 ();
 sg13g2_decap_8 FILLER_39_1391 ();
 sg13g2_decap_8 FILLER_39_1398 ();
 sg13g2_decap_8 FILLER_39_1405 ();
 sg13g2_decap_8 FILLER_39_1412 ();
 sg13g2_decap_8 FILLER_39_1419 ();
 sg13g2_decap_8 FILLER_39_1426 ();
 sg13g2_decap_8 FILLER_39_1433 ();
 sg13g2_decap_8 FILLER_39_1440 ();
 sg13g2_decap_8 FILLER_39_1447 ();
 sg13g2_decap_8 FILLER_39_1454 ();
 sg13g2_decap_8 FILLER_39_1461 ();
 sg13g2_decap_8 FILLER_39_1468 ();
 sg13g2_decap_8 FILLER_39_1475 ();
 sg13g2_decap_8 FILLER_39_1482 ();
 sg13g2_decap_8 FILLER_39_1489 ();
 sg13g2_decap_8 FILLER_39_1496 ();
 sg13g2_decap_8 FILLER_39_1503 ();
 sg13g2_decap_8 FILLER_39_1510 ();
 sg13g2_decap_8 FILLER_39_1517 ();
 sg13g2_decap_8 FILLER_39_1524 ();
 sg13g2_decap_8 FILLER_39_1531 ();
 sg13g2_decap_8 FILLER_39_1538 ();
 sg13g2_decap_8 FILLER_39_1545 ();
 sg13g2_decap_8 FILLER_39_1552 ();
 sg13g2_decap_8 FILLER_39_1559 ();
 sg13g2_decap_8 FILLER_39_1566 ();
 sg13g2_decap_8 FILLER_39_1573 ();
 sg13g2_decap_8 FILLER_39_1580 ();
 sg13g2_decap_8 FILLER_39_1587 ();
 sg13g2_decap_8 FILLER_39_1594 ();
 sg13g2_decap_8 FILLER_39_1601 ();
 sg13g2_decap_8 FILLER_39_1608 ();
 sg13g2_decap_8 FILLER_39_1615 ();
 sg13g2_decap_8 FILLER_39_1622 ();
 sg13g2_decap_8 FILLER_39_1629 ();
 sg13g2_decap_8 FILLER_39_1636 ();
 sg13g2_decap_8 FILLER_39_1643 ();
 sg13g2_decap_8 FILLER_39_1650 ();
 sg13g2_decap_8 FILLER_39_1657 ();
 sg13g2_decap_8 FILLER_39_1664 ();
 sg13g2_decap_8 FILLER_39_1671 ();
 sg13g2_decap_8 FILLER_39_1678 ();
 sg13g2_decap_8 FILLER_39_1685 ();
 sg13g2_decap_8 FILLER_39_1692 ();
 sg13g2_decap_8 FILLER_39_1699 ();
 sg13g2_decap_8 FILLER_39_1706 ();
 sg13g2_decap_8 FILLER_39_1713 ();
 sg13g2_decap_8 FILLER_39_1720 ();
 sg13g2_decap_8 FILLER_39_1727 ();
 sg13g2_decap_8 FILLER_39_1734 ();
 sg13g2_decap_8 FILLER_39_1741 ();
 sg13g2_decap_8 FILLER_39_1748 ();
 sg13g2_decap_8 FILLER_39_1755 ();
 sg13g2_decap_4 FILLER_39_1762 ();
 sg13g2_fill_2 FILLER_39_1766 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_14 ();
 sg13g2_decap_8 FILLER_40_21 ();
 sg13g2_decap_8 FILLER_40_28 ();
 sg13g2_decap_8 FILLER_40_35 ();
 sg13g2_decap_8 FILLER_40_42 ();
 sg13g2_decap_8 FILLER_40_49 ();
 sg13g2_decap_8 FILLER_40_56 ();
 sg13g2_decap_8 FILLER_40_63 ();
 sg13g2_decap_8 FILLER_40_70 ();
 sg13g2_decap_8 FILLER_40_77 ();
 sg13g2_decap_8 FILLER_40_84 ();
 sg13g2_decap_8 FILLER_40_91 ();
 sg13g2_decap_8 FILLER_40_98 ();
 sg13g2_decap_8 FILLER_40_105 ();
 sg13g2_decap_8 FILLER_40_112 ();
 sg13g2_decap_8 FILLER_40_119 ();
 sg13g2_decap_8 FILLER_40_126 ();
 sg13g2_decap_8 FILLER_40_133 ();
 sg13g2_decap_8 FILLER_40_140 ();
 sg13g2_decap_8 FILLER_40_147 ();
 sg13g2_decap_8 FILLER_40_154 ();
 sg13g2_decap_4 FILLER_40_161 ();
 sg13g2_fill_2 FILLER_40_165 ();
 sg13g2_decap_4 FILLER_40_171 ();
 sg13g2_fill_1 FILLER_40_175 ();
 sg13g2_fill_1 FILLER_40_188 ();
 sg13g2_fill_2 FILLER_40_201 ();
 sg13g2_decap_4 FILLER_40_304 ();
 sg13g2_decap_4 FILLER_40_336 ();
 sg13g2_fill_1 FILLER_40_340 ();
 sg13g2_fill_2 FILLER_40_346 ();
 sg13g2_fill_1 FILLER_40_348 ();
 sg13g2_fill_1 FILLER_40_354 ();
 sg13g2_fill_2 FILLER_40_360 ();
 sg13g2_decap_8 FILLER_40_375 ();
 sg13g2_decap_4 FILLER_40_382 ();
 sg13g2_fill_2 FILLER_40_386 ();
 sg13g2_fill_2 FILLER_40_400 ();
 sg13g2_fill_1 FILLER_40_402 ();
 sg13g2_fill_2 FILLER_40_429 ();
 sg13g2_decap_8 FILLER_40_491 ();
 sg13g2_decap_8 FILLER_40_498 ();
 sg13g2_fill_2 FILLER_40_505 ();
 sg13g2_decap_8 FILLER_40_527 ();
 sg13g2_fill_2 FILLER_40_534 ();
 sg13g2_fill_2 FILLER_40_558 ();
 sg13g2_fill_1 FILLER_40_560 ();
 sg13g2_fill_1 FILLER_40_586 ();
 sg13g2_decap_4 FILLER_40_604 ();
 sg13g2_fill_2 FILLER_40_630 ();
 sg13g2_fill_1 FILLER_40_678 ();
 sg13g2_fill_1 FILLER_40_722 ();
 sg13g2_decap_8 FILLER_40_743 ();
 sg13g2_fill_2 FILLER_40_750 ();
 sg13g2_fill_1 FILLER_40_752 ();
 sg13g2_decap_4 FILLER_40_768 ();
 sg13g2_fill_1 FILLER_40_772 ();
 sg13g2_fill_2 FILLER_40_805 ();
 sg13g2_decap_4 FILLER_40_810 ();
 sg13g2_decap_4 FILLER_40_828 ();
 sg13g2_fill_2 FILLER_40_832 ();
 sg13g2_decap_8 FILLER_40_839 ();
 sg13g2_decap_8 FILLER_40_846 ();
 sg13g2_decap_8 FILLER_40_853 ();
 sg13g2_decap_8 FILLER_40_860 ();
 sg13g2_fill_2 FILLER_40_867 ();
 sg13g2_decap_8 FILLER_40_874 ();
 sg13g2_fill_2 FILLER_40_881 ();
 sg13g2_decap_8 FILLER_40_893 ();
 sg13g2_fill_2 FILLER_40_900 ();
 sg13g2_fill_1 FILLER_40_902 ();
 sg13g2_fill_1 FILLER_40_967 ();
 sg13g2_fill_1 FILLER_40_973 ();
 sg13g2_fill_1 FILLER_40_1025 ();
 sg13g2_fill_2 FILLER_40_1048 ();
 sg13g2_fill_1 FILLER_40_1050 ();
 sg13g2_decap_8 FILLER_40_1086 ();
 sg13g2_fill_2 FILLER_40_1093 ();
 sg13g2_fill_1 FILLER_40_1095 ();
 sg13g2_decap_8 FILLER_40_1105 ();
 sg13g2_decap_8 FILLER_40_1112 ();
 sg13g2_decap_8 FILLER_40_1119 ();
 sg13g2_decap_8 FILLER_40_1126 ();
 sg13g2_decap_8 FILLER_40_1133 ();
 sg13g2_decap_8 FILLER_40_1140 ();
 sg13g2_decap_8 FILLER_40_1147 ();
 sg13g2_decap_8 FILLER_40_1154 ();
 sg13g2_decap_8 FILLER_40_1161 ();
 sg13g2_decap_8 FILLER_40_1168 ();
 sg13g2_decap_8 FILLER_40_1175 ();
 sg13g2_decap_8 FILLER_40_1182 ();
 sg13g2_decap_8 FILLER_40_1189 ();
 sg13g2_decap_8 FILLER_40_1196 ();
 sg13g2_decap_8 FILLER_40_1203 ();
 sg13g2_decap_8 FILLER_40_1210 ();
 sg13g2_decap_8 FILLER_40_1217 ();
 sg13g2_decap_8 FILLER_40_1224 ();
 sg13g2_decap_8 FILLER_40_1231 ();
 sg13g2_decap_8 FILLER_40_1238 ();
 sg13g2_decap_8 FILLER_40_1245 ();
 sg13g2_decap_8 FILLER_40_1252 ();
 sg13g2_decap_8 FILLER_40_1259 ();
 sg13g2_decap_8 FILLER_40_1266 ();
 sg13g2_decap_8 FILLER_40_1273 ();
 sg13g2_decap_8 FILLER_40_1280 ();
 sg13g2_decap_8 FILLER_40_1287 ();
 sg13g2_decap_8 FILLER_40_1294 ();
 sg13g2_decap_8 FILLER_40_1301 ();
 sg13g2_decap_8 FILLER_40_1308 ();
 sg13g2_decap_8 FILLER_40_1315 ();
 sg13g2_decap_8 FILLER_40_1322 ();
 sg13g2_decap_8 FILLER_40_1329 ();
 sg13g2_decap_8 FILLER_40_1336 ();
 sg13g2_decap_8 FILLER_40_1343 ();
 sg13g2_decap_8 FILLER_40_1350 ();
 sg13g2_decap_8 FILLER_40_1357 ();
 sg13g2_decap_8 FILLER_40_1364 ();
 sg13g2_decap_8 FILLER_40_1371 ();
 sg13g2_decap_8 FILLER_40_1378 ();
 sg13g2_decap_8 FILLER_40_1385 ();
 sg13g2_decap_8 FILLER_40_1392 ();
 sg13g2_decap_8 FILLER_40_1399 ();
 sg13g2_decap_8 FILLER_40_1406 ();
 sg13g2_decap_8 FILLER_40_1413 ();
 sg13g2_decap_8 FILLER_40_1420 ();
 sg13g2_decap_8 FILLER_40_1427 ();
 sg13g2_decap_8 FILLER_40_1434 ();
 sg13g2_decap_8 FILLER_40_1441 ();
 sg13g2_decap_8 FILLER_40_1448 ();
 sg13g2_decap_8 FILLER_40_1455 ();
 sg13g2_decap_8 FILLER_40_1462 ();
 sg13g2_decap_8 FILLER_40_1469 ();
 sg13g2_decap_8 FILLER_40_1476 ();
 sg13g2_decap_8 FILLER_40_1483 ();
 sg13g2_decap_8 FILLER_40_1490 ();
 sg13g2_decap_8 FILLER_40_1497 ();
 sg13g2_decap_8 FILLER_40_1504 ();
 sg13g2_decap_8 FILLER_40_1511 ();
 sg13g2_decap_8 FILLER_40_1518 ();
 sg13g2_decap_8 FILLER_40_1525 ();
 sg13g2_decap_8 FILLER_40_1532 ();
 sg13g2_decap_8 FILLER_40_1539 ();
 sg13g2_decap_8 FILLER_40_1546 ();
 sg13g2_decap_8 FILLER_40_1553 ();
 sg13g2_decap_8 FILLER_40_1560 ();
 sg13g2_decap_8 FILLER_40_1567 ();
 sg13g2_decap_8 FILLER_40_1574 ();
 sg13g2_decap_8 FILLER_40_1581 ();
 sg13g2_decap_8 FILLER_40_1588 ();
 sg13g2_decap_8 FILLER_40_1595 ();
 sg13g2_decap_8 FILLER_40_1602 ();
 sg13g2_decap_8 FILLER_40_1609 ();
 sg13g2_decap_8 FILLER_40_1616 ();
 sg13g2_decap_8 FILLER_40_1623 ();
 sg13g2_decap_8 FILLER_40_1630 ();
 sg13g2_decap_8 FILLER_40_1637 ();
 sg13g2_decap_8 FILLER_40_1644 ();
 sg13g2_decap_8 FILLER_40_1651 ();
 sg13g2_decap_8 FILLER_40_1658 ();
 sg13g2_decap_8 FILLER_40_1665 ();
 sg13g2_decap_8 FILLER_40_1672 ();
 sg13g2_decap_8 FILLER_40_1679 ();
 sg13g2_decap_8 FILLER_40_1686 ();
 sg13g2_decap_8 FILLER_40_1693 ();
 sg13g2_decap_8 FILLER_40_1700 ();
 sg13g2_decap_8 FILLER_40_1707 ();
 sg13g2_decap_8 FILLER_40_1714 ();
 sg13g2_decap_8 FILLER_40_1721 ();
 sg13g2_decap_8 FILLER_40_1728 ();
 sg13g2_decap_8 FILLER_40_1735 ();
 sg13g2_decap_8 FILLER_40_1742 ();
 sg13g2_decap_8 FILLER_40_1749 ();
 sg13g2_decap_8 FILLER_40_1756 ();
 sg13g2_decap_4 FILLER_40_1763 ();
 sg13g2_fill_1 FILLER_40_1767 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_8 FILLER_41_14 ();
 sg13g2_decap_8 FILLER_41_21 ();
 sg13g2_decap_8 FILLER_41_28 ();
 sg13g2_decap_8 FILLER_41_35 ();
 sg13g2_decap_8 FILLER_41_42 ();
 sg13g2_decap_8 FILLER_41_49 ();
 sg13g2_decap_8 FILLER_41_56 ();
 sg13g2_decap_8 FILLER_41_63 ();
 sg13g2_decap_8 FILLER_41_70 ();
 sg13g2_decap_8 FILLER_41_77 ();
 sg13g2_decap_8 FILLER_41_84 ();
 sg13g2_decap_8 FILLER_41_91 ();
 sg13g2_decap_8 FILLER_41_98 ();
 sg13g2_decap_8 FILLER_41_105 ();
 sg13g2_decap_8 FILLER_41_112 ();
 sg13g2_decap_8 FILLER_41_119 ();
 sg13g2_decap_8 FILLER_41_126 ();
 sg13g2_decap_8 FILLER_41_133 ();
 sg13g2_decap_8 FILLER_41_140 ();
 sg13g2_decap_8 FILLER_41_147 ();
 sg13g2_decap_8 FILLER_41_154 ();
 sg13g2_fill_2 FILLER_41_161 ();
 sg13g2_fill_1 FILLER_41_189 ();
 sg13g2_fill_2 FILLER_41_199 ();
 sg13g2_fill_2 FILLER_41_210 ();
 sg13g2_fill_1 FILLER_41_215 ();
 sg13g2_fill_2 FILLER_41_243 ();
 sg13g2_fill_1 FILLER_41_245 ();
 sg13g2_fill_2 FILLER_41_255 ();
 sg13g2_decap_4 FILLER_41_306 ();
 sg13g2_fill_2 FILLER_41_310 ();
 sg13g2_fill_1 FILLER_41_334 ();
 sg13g2_fill_2 FILLER_41_364 ();
 sg13g2_fill_2 FILLER_41_378 ();
 sg13g2_fill_2 FILLER_41_405 ();
 sg13g2_decap_8 FILLER_41_424 ();
 sg13g2_decap_4 FILLER_41_431 ();
 sg13g2_fill_2 FILLER_41_447 ();
 sg13g2_decap_8 FILLER_41_462 ();
 sg13g2_decap_4 FILLER_41_482 ();
 sg13g2_fill_1 FILLER_41_536 ();
 sg13g2_decap_8 FILLER_41_561 ();
 sg13g2_decap_4 FILLER_41_568 ();
 sg13g2_decap_4 FILLER_41_580 ();
 sg13g2_decap_8 FILLER_41_601 ();
 sg13g2_decap_8 FILLER_41_608 ();
 sg13g2_fill_2 FILLER_41_615 ();
 sg13g2_fill_1 FILLER_41_617 ();
 sg13g2_decap_4 FILLER_41_630 ();
 sg13g2_fill_2 FILLER_41_634 ();
 sg13g2_fill_1 FILLER_41_665 ();
 sg13g2_fill_2 FILLER_41_719 ();
 sg13g2_fill_1 FILLER_41_742 ();
 sg13g2_fill_2 FILLER_41_748 ();
 sg13g2_fill_1 FILLER_41_755 ();
 sg13g2_fill_2 FILLER_41_764 ();
 sg13g2_fill_1 FILLER_41_766 ();
 sg13g2_fill_2 FILLER_41_783 ();
 sg13g2_fill_2 FILLER_41_845 ();
 sg13g2_fill_1 FILLER_41_847 ();
 sg13g2_decap_8 FILLER_41_853 ();
 sg13g2_fill_2 FILLER_41_860 ();
 sg13g2_fill_1 FILLER_41_862 ();
 sg13g2_fill_2 FILLER_41_912 ();
 sg13g2_fill_1 FILLER_41_955 ();
 sg13g2_fill_2 FILLER_41_992 ();
 sg13g2_decap_8 FILLER_41_1064 ();
 sg13g2_decap_8 FILLER_41_1071 ();
 sg13g2_decap_8 FILLER_41_1078 ();
 sg13g2_decap_8 FILLER_41_1085 ();
 sg13g2_decap_8 FILLER_41_1092 ();
 sg13g2_decap_8 FILLER_41_1099 ();
 sg13g2_decap_8 FILLER_41_1106 ();
 sg13g2_decap_8 FILLER_41_1113 ();
 sg13g2_decap_8 FILLER_41_1120 ();
 sg13g2_decap_8 FILLER_41_1127 ();
 sg13g2_decap_8 FILLER_41_1134 ();
 sg13g2_decap_8 FILLER_41_1141 ();
 sg13g2_decap_8 FILLER_41_1148 ();
 sg13g2_decap_8 FILLER_41_1155 ();
 sg13g2_decap_8 FILLER_41_1162 ();
 sg13g2_decap_8 FILLER_41_1169 ();
 sg13g2_decap_8 FILLER_41_1176 ();
 sg13g2_decap_8 FILLER_41_1183 ();
 sg13g2_decap_8 FILLER_41_1190 ();
 sg13g2_decap_8 FILLER_41_1197 ();
 sg13g2_decap_8 FILLER_41_1204 ();
 sg13g2_decap_8 FILLER_41_1211 ();
 sg13g2_decap_8 FILLER_41_1218 ();
 sg13g2_decap_8 FILLER_41_1225 ();
 sg13g2_decap_8 FILLER_41_1232 ();
 sg13g2_decap_8 FILLER_41_1239 ();
 sg13g2_decap_8 FILLER_41_1246 ();
 sg13g2_decap_8 FILLER_41_1253 ();
 sg13g2_decap_8 FILLER_41_1260 ();
 sg13g2_decap_8 FILLER_41_1267 ();
 sg13g2_decap_8 FILLER_41_1274 ();
 sg13g2_decap_8 FILLER_41_1281 ();
 sg13g2_decap_8 FILLER_41_1288 ();
 sg13g2_decap_8 FILLER_41_1295 ();
 sg13g2_decap_8 FILLER_41_1302 ();
 sg13g2_decap_8 FILLER_41_1309 ();
 sg13g2_decap_8 FILLER_41_1316 ();
 sg13g2_decap_8 FILLER_41_1323 ();
 sg13g2_decap_8 FILLER_41_1330 ();
 sg13g2_decap_8 FILLER_41_1337 ();
 sg13g2_decap_8 FILLER_41_1344 ();
 sg13g2_decap_8 FILLER_41_1351 ();
 sg13g2_decap_8 FILLER_41_1358 ();
 sg13g2_decap_8 FILLER_41_1365 ();
 sg13g2_decap_8 FILLER_41_1372 ();
 sg13g2_decap_8 FILLER_41_1379 ();
 sg13g2_decap_8 FILLER_41_1386 ();
 sg13g2_decap_8 FILLER_41_1393 ();
 sg13g2_decap_8 FILLER_41_1400 ();
 sg13g2_decap_8 FILLER_41_1407 ();
 sg13g2_decap_8 FILLER_41_1414 ();
 sg13g2_decap_8 FILLER_41_1421 ();
 sg13g2_decap_8 FILLER_41_1428 ();
 sg13g2_decap_8 FILLER_41_1435 ();
 sg13g2_decap_8 FILLER_41_1442 ();
 sg13g2_decap_8 FILLER_41_1449 ();
 sg13g2_decap_8 FILLER_41_1456 ();
 sg13g2_decap_8 FILLER_41_1463 ();
 sg13g2_decap_8 FILLER_41_1470 ();
 sg13g2_decap_8 FILLER_41_1477 ();
 sg13g2_decap_8 FILLER_41_1484 ();
 sg13g2_decap_8 FILLER_41_1491 ();
 sg13g2_decap_8 FILLER_41_1498 ();
 sg13g2_decap_8 FILLER_41_1505 ();
 sg13g2_decap_8 FILLER_41_1512 ();
 sg13g2_decap_8 FILLER_41_1519 ();
 sg13g2_decap_8 FILLER_41_1526 ();
 sg13g2_decap_8 FILLER_41_1533 ();
 sg13g2_decap_8 FILLER_41_1540 ();
 sg13g2_decap_8 FILLER_41_1547 ();
 sg13g2_decap_8 FILLER_41_1554 ();
 sg13g2_decap_8 FILLER_41_1561 ();
 sg13g2_decap_8 FILLER_41_1568 ();
 sg13g2_decap_8 FILLER_41_1575 ();
 sg13g2_decap_8 FILLER_41_1582 ();
 sg13g2_decap_8 FILLER_41_1589 ();
 sg13g2_decap_8 FILLER_41_1596 ();
 sg13g2_decap_8 FILLER_41_1603 ();
 sg13g2_decap_8 FILLER_41_1610 ();
 sg13g2_decap_8 FILLER_41_1617 ();
 sg13g2_decap_8 FILLER_41_1624 ();
 sg13g2_decap_8 FILLER_41_1631 ();
 sg13g2_decap_8 FILLER_41_1638 ();
 sg13g2_decap_8 FILLER_41_1645 ();
 sg13g2_decap_8 FILLER_41_1652 ();
 sg13g2_decap_8 FILLER_41_1659 ();
 sg13g2_decap_8 FILLER_41_1666 ();
 sg13g2_decap_8 FILLER_41_1673 ();
 sg13g2_decap_8 FILLER_41_1680 ();
 sg13g2_decap_8 FILLER_41_1687 ();
 sg13g2_decap_8 FILLER_41_1694 ();
 sg13g2_decap_8 FILLER_41_1701 ();
 sg13g2_decap_8 FILLER_41_1708 ();
 sg13g2_decap_8 FILLER_41_1715 ();
 sg13g2_decap_8 FILLER_41_1722 ();
 sg13g2_decap_8 FILLER_41_1729 ();
 sg13g2_decap_8 FILLER_41_1736 ();
 sg13g2_decap_8 FILLER_41_1743 ();
 sg13g2_decap_8 FILLER_41_1750 ();
 sg13g2_decap_8 FILLER_41_1757 ();
 sg13g2_decap_4 FILLER_41_1764 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_decap_8 FILLER_42_14 ();
 sg13g2_decap_8 FILLER_42_21 ();
 sg13g2_decap_8 FILLER_42_28 ();
 sg13g2_decap_8 FILLER_42_35 ();
 sg13g2_decap_8 FILLER_42_42 ();
 sg13g2_decap_8 FILLER_42_49 ();
 sg13g2_decap_8 FILLER_42_56 ();
 sg13g2_decap_8 FILLER_42_63 ();
 sg13g2_decap_8 FILLER_42_70 ();
 sg13g2_decap_8 FILLER_42_77 ();
 sg13g2_decap_8 FILLER_42_84 ();
 sg13g2_decap_8 FILLER_42_91 ();
 sg13g2_decap_8 FILLER_42_98 ();
 sg13g2_decap_8 FILLER_42_105 ();
 sg13g2_decap_8 FILLER_42_112 ();
 sg13g2_decap_8 FILLER_42_119 ();
 sg13g2_decap_8 FILLER_42_126 ();
 sg13g2_decap_8 FILLER_42_133 ();
 sg13g2_decap_8 FILLER_42_140 ();
 sg13g2_decap_8 FILLER_42_147 ();
 sg13g2_decap_8 FILLER_42_154 ();
 sg13g2_decap_8 FILLER_42_161 ();
 sg13g2_decap_8 FILLER_42_171 ();
 sg13g2_fill_1 FILLER_42_178 ();
 sg13g2_decap_4 FILLER_42_212 ();
 sg13g2_fill_1 FILLER_42_289 ();
 sg13g2_decap_8 FILLER_42_328 ();
 sg13g2_decap_4 FILLER_42_335 ();
 sg13g2_fill_2 FILLER_42_339 ();
 sg13g2_decap_4 FILLER_42_357 ();
 sg13g2_fill_1 FILLER_42_361 ();
 sg13g2_decap_8 FILLER_42_374 ();
 sg13g2_decap_8 FILLER_42_381 ();
 sg13g2_fill_2 FILLER_42_388 ();
 sg13g2_decap_4 FILLER_42_428 ();
 sg13g2_fill_2 FILLER_42_432 ();
 sg13g2_decap_4 FILLER_42_443 ();
 sg13g2_fill_2 FILLER_42_447 ();
 sg13g2_decap_4 FILLER_42_465 ();
 sg13g2_fill_2 FILLER_42_469 ();
 sg13g2_decap_8 FILLER_42_483 ();
 sg13g2_decap_8 FILLER_42_490 ();
 sg13g2_decap_4 FILLER_42_497 ();
 sg13g2_decap_4 FILLER_42_505 ();
 sg13g2_decap_8 FILLER_42_526 ();
 sg13g2_decap_8 FILLER_42_533 ();
 sg13g2_fill_1 FILLER_42_540 ();
 sg13g2_fill_1 FILLER_42_546 ();
 sg13g2_decap_4 FILLER_42_559 ();
 sg13g2_fill_2 FILLER_42_563 ();
 sg13g2_fill_1 FILLER_42_584 ();
 sg13g2_fill_2 FILLER_42_599 ();
 sg13g2_decap_8 FILLER_42_609 ();
 sg13g2_fill_2 FILLER_42_616 ();
 sg13g2_fill_1 FILLER_42_618 ();
 sg13g2_fill_2 FILLER_42_640 ();
 sg13g2_fill_1 FILLER_42_642 ();
 sg13g2_fill_1 FILLER_42_656 ();
 sg13g2_fill_2 FILLER_42_739 ();
 sg13g2_fill_2 FILLER_42_764 ();
 sg13g2_fill_1 FILLER_42_766 ();
 sg13g2_decap_4 FILLER_42_779 ();
 sg13g2_decap_8 FILLER_42_808 ();
 sg13g2_fill_2 FILLER_42_815 ();
 sg13g2_fill_1 FILLER_42_817 ();
 sg13g2_decap_8 FILLER_42_823 ();
 sg13g2_decap_4 FILLER_42_830 ();
 sg13g2_fill_2 FILLER_42_837 ();
 sg13g2_fill_1 FILLER_42_839 ();
 sg13g2_decap_4 FILLER_42_849 ();
 sg13g2_fill_1 FILLER_42_876 ();
 sg13g2_decap_8 FILLER_42_898 ();
 sg13g2_decap_4 FILLER_42_905 ();
 sg13g2_fill_2 FILLER_42_931 ();
 sg13g2_fill_1 FILLER_42_960 ();
 sg13g2_fill_2 FILLER_42_974 ();
 sg13g2_fill_1 FILLER_42_976 ();
 sg13g2_decap_4 FILLER_42_997 ();
 sg13g2_decap_8 FILLER_42_1028 ();
 sg13g2_decap_8 FILLER_42_1035 ();
 sg13g2_decap_8 FILLER_42_1042 ();
 sg13g2_decap_8 FILLER_42_1049 ();
 sg13g2_decap_8 FILLER_42_1056 ();
 sg13g2_decap_8 FILLER_42_1063 ();
 sg13g2_decap_8 FILLER_42_1070 ();
 sg13g2_decap_8 FILLER_42_1077 ();
 sg13g2_decap_8 FILLER_42_1084 ();
 sg13g2_decap_8 FILLER_42_1091 ();
 sg13g2_decap_8 FILLER_42_1098 ();
 sg13g2_decap_8 FILLER_42_1105 ();
 sg13g2_decap_8 FILLER_42_1112 ();
 sg13g2_decap_8 FILLER_42_1119 ();
 sg13g2_decap_8 FILLER_42_1126 ();
 sg13g2_decap_8 FILLER_42_1133 ();
 sg13g2_decap_8 FILLER_42_1140 ();
 sg13g2_decap_8 FILLER_42_1147 ();
 sg13g2_decap_8 FILLER_42_1154 ();
 sg13g2_decap_8 FILLER_42_1161 ();
 sg13g2_decap_8 FILLER_42_1168 ();
 sg13g2_decap_8 FILLER_42_1175 ();
 sg13g2_decap_8 FILLER_42_1182 ();
 sg13g2_decap_8 FILLER_42_1189 ();
 sg13g2_decap_8 FILLER_42_1196 ();
 sg13g2_decap_8 FILLER_42_1203 ();
 sg13g2_decap_8 FILLER_42_1210 ();
 sg13g2_decap_8 FILLER_42_1217 ();
 sg13g2_decap_8 FILLER_42_1224 ();
 sg13g2_decap_8 FILLER_42_1231 ();
 sg13g2_decap_8 FILLER_42_1238 ();
 sg13g2_decap_8 FILLER_42_1245 ();
 sg13g2_decap_8 FILLER_42_1252 ();
 sg13g2_decap_8 FILLER_42_1259 ();
 sg13g2_decap_8 FILLER_42_1266 ();
 sg13g2_decap_8 FILLER_42_1273 ();
 sg13g2_decap_8 FILLER_42_1280 ();
 sg13g2_decap_8 FILLER_42_1287 ();
 sg13g2_decap_8 FILLER_42_1294 ();
 sg13g2_decap_8 FILLER_42_1301 ();
 sg13g2_decap_8 FILLER_42_1308 ();
 sg13g2_decap_8 FILLER_42_1315 ();
 sg13g2_decap_8 FILLER_42_1322 ();
 sg13g2_decap_8 FILLER_42_1329 ();
 sg13g2_decap_8 FILLER_42_1336 ();
 sg13g2_decap_8 FILLER_42_1343 ();
 sg13g2_decap_8 FILLER_42_1350 ();
 sg13g2_decap_8 FILLER_42_1357 ();
 sg13g2_decap_8 FILLER_42_1364 ();
 sg13g2_decap_8 FILLER_42_1371 ();
 sg13g2_decap_8 FILLER_42_1378 ();
 sg13g2_decap_8 FILLER_42_1385 ();
 sg13g2_decap_8 FILLER_42_1392 ();
 sg13g2_decap_8 FILLER_42_1399 ();
 sg13g2_decap_8 FILLER_42_1406 ();
 sg13g2_decap_8 FILLER_42_1413 ();
 sg13g2_decap_8 FILLER_42_1420 ();
 sg13g2_decap_8 FILLER_42_1427 ();
 sg13g2_decap_8 FILLER_42_1434 ();
 sg13g2_decap_8 FILLER_42_1441 ();
 sg13g2_decap_8 FILLER_42_1448 ();
 sg13g2_decap_8 FILLER_42_1455 ();
 sg13g2_decap_8 FILLER_42_1462 ();
 sg13g2_decap_8 FILLER_42_1469 ();
 sg13g2_decap_8 FILLER_42_1476 ();
 sg13g2_decap_8 FILLER_42_1483 ();
 sg13g2_decap_8 FILLER_42_1490 ();
 sg13g2_decap_8 FILLER_42_1497 ();
 sg13g2_decap_8 FILLER_42_1504 ();
 sg13g2_decap_8 FILLER_42_1511 ();
 sg13g2_decap_8 FILLER_42_1518 ();
 sg13g2_decap_8 FILLER_42_1525 ();
 sg13g2_decap_8 FILLER_42_1532 ();
 sg13g2_decap_8 FILLER_42_1539 ();
 sg13g2_decap_8 FILLER_42_1546 ();
 sg13g2_decap_8 FILLER_42_1553 ();
 sg13g2_decap_8 FILLER_42_1560 ();
 sg13g2_decap_8 FILLER_42_1567 ();
 sg13g2_decap_8 FILLER_42_1574 ();
 sg13g2_decap_8 FILLER_42_1581 ();
 sg13g2_decap_8 FILLER_42_1588 ();
 sg13g2_decap_8 FILLER_42_1595 ();
 sg13g2_decap_8 FILLER_42_1602 ();
 sg13g2_decap_8 FILLER_42_1609 ();
 sg13g2_decap_8 FILLER_42_1616 ();
 sg13g2_decap_8 FILLER_42_1623 ();
 sg13g2_decap_8 FILLER_42_1630 ();
 sg13g2_decap_8 FILLER_42_1637 ();
 sg13g2_decap_8 FILLER_42_1644 ();
 sg13g2_decap_8 FILLER_42_1651 ();
 sg13g2_decap_8 FILLER_42_1658 ();
 sg13g2_decap_8 FILLER_42_1665 ();
 sg13g2_decap_8 FILLER_42_1672 ();
 sg13g2_decap_8 FILLER_42_1679 ();
 sg13g2_decap_8 FILLER_42_1686 ();
 sg13g2_decap_8 FILLER_42_1693 ();
 sg13g2_decap_8 FILLER_42_1700 ();
 sg13g2_decap_8 FILLER_42_1707 ();
 sg13g2_decap_8 FILLER_42_1714 ();
 sg13g2_decap_8 FILLER_42_1721 ();
 sg13g2_decap_8 FILLER_42_1728 ();
 sg13g2_decap_8 FILLER_42_1735 ();
 sg13g2_decap_8 FILLER_42_1742 ();
 sg13g2_decap_8 FILLER_42_1749 ();
 sg13g2_decap_8 FILLER_42_1756 ();
 sg13g2_decap_4 FILLER_42_1763 ();
 sg13g2_fill_1 FILLER_42_1767 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_decap_8 FILLER_43_14 ();
 sg13g2_decap_8 FILLER_43_21 ();
 sg13g2_decap_8 FILLER_43_28 ();
 sg13g2_decap_8 FILLER_43_35 ();
 sg13g2_decap_8 FILLER_43_42 ();
 sg13g2_decap_8 FILLER_43_49 ();
 sg13g2_decap_8 FILLER_43_56 ();
 sg13g2_decap_8 FILLER_43_63 ();
 sg13g2_decap_8 FILLER_43_70 ();
 sg13g2_decap_8 FILLER_43_77 ();
 sg13g2_decap_8 FILLER_43_84 ();
 sg13g2_decap_8 FILLER_43_91 ();
 sg13g2_decap_8 FILLER_43_98 ();
 sg13g2_decap_8 FILLER_43_105 ();
 sg13g2_decap_8 FILLER_43_112 ();
 sg13g2_decap_8 FILLER_43_119 ();
 sg13g2_decap_8 FILLER_43_126 ();
 sg13g2_decap_8 FILLER_43_133 ();
 sg13g2_decap_8 FILLER_43_140 ();
 sg13g2_decap_8 FILLER_43_147 ();
 sg13g2_decap_8 FILLER_43_154 ();
 sg13g2_decap_4 FILLER_43_161 ();
 sg13g2_fill_2 FILLER_43_252 ();
 sg13g2_decap_8 FILLER_43_308 ();
 sg13g2_fill_2 FILLER_43_336 ();
 sg13g2_fill_1 FILLER_43_338 ();
 sg13g2_fill_2 FILLER_43_351 ();
 sg13g2_fill_1 FILLER_43_353 ();
 sg13g2_fill_2 FILLER_43_376 ();
 sg13g2_fill_1 FILLER_43_378 ();
 sg13g2_decap_4 FILLER_43_384 ();
 sg13g2_decap_8 FILLER_43_400 ();
 sg13g2_decap_4 FILLER_43_407 ();
 sg13g2_fill_1 FILLER_43_424 ();
 sg13g2_fill_2 FILLER_43_446 ();
 sg13g2_fill_1 FILLER_43_463 ();
 sg13g2_decap_4 FILLER_43_514 ();
 sg13g2_fill_1 FILLER_43_518 ();
 sg13g2_decap_8 FILLER_43_527 ();
 sg13g2_fill_1 FILLER_43_534 ();
 sg13g2_decap_8 FILLER_43_560 ();
 sg13g2_fill_1 FILLER_43_567 ();
 sg13g2_decap_4 FILLER_43_573 ();
 sg13g2_fill_2 FILLER_43_577 ();
 sg13g2_fill_1 FILLER_43_591 ();
 sg13g2_fill_2 FILLER_43_600 ();
 sg13g2_fill_1 FILLER_43_602 ();
 sg13g2_decap_8 FILLER_43_610 ();
 sg13g2_fill_2 FILLER_43_617 ();
 sg13g2_decap_4 FILLER_43_660 ();
 sg13g2_fill_1 FILLER_43_664 ();
 sg13g2_decap_8 FILLER_43_670 ();
 sg13g2_fill_2 FILLER_43_677 ();
 sg13g2_fill_1 FILLER_43_679 ();
 sg13g2_decap_4 FILLER_43_686 ();
 sg13g2_decap_4 FILLER_43_723 ();
 sg13g2_fill_1 FILLER_43_732 ();
 sg13g2_fill_1 FILLER_43_746 ();
 sg13g2_decap_4 FILLER_43_761 ();
 sg13g2_fill_1 FILLER_43_765 ();
 sg13g2_fill_1 FILLER_43_771 ();
 sg13g2_fill_1 FILLER_43_778 ();
 sg13g2_fill_2 FILLER_43_794 ();
 sg13g2_fill_1 FILLER_43_796 ();
 sg13g2_fill_1 FILLER_43_805 ();
 sg13g2_fill_2 FILLER_43_819 ();
 sg13g2_fill_1 FILLER_43_833 ();
 sg13g2_decap_8 FILLER_43_861 ();
 sg13g2_decap_8 FILLER_43_868 ();
 sg13g2_decap_8 FILLER_43_875 ();
 sg13g2_fill_2 FILLER_43_882 ();
 sg13g2_decap_4 FILLER_43_896 ();
 sg13g2_decap_4 FILLER_43_912 ();
 sg13g2_fill_1 FILLER_43_916 ();
 sg13g2_fill_1 FILLER_43_923 ();
 sg13g2_decap_8 FILLER_43_936 ();
 sg13g2_decap_8 FILLER_43_943 ();
 sg13g2_decap_8 FILLER_43_950 ();
 sg13g2_fill_2 FILLER_43_957 ();
 sg13g2_fill_1 FILLER_43_968 ();
 sg13g2_decap_4 FILLER_43_977 ();
 sg13g2_fill_1 FILLER_43_981 ();
 sg13g2_decap_8 FILLER_43_1034 ();
 sg13g2_decap_8 FILLER_43_1041 ();
 sg13g2_decap_8 FILLER_43_1048 ();
 sg13g2_decap_8 FILLER_43_1055 ();
 sg13g2_decap_8 FILLER_43_1062 ();
 sg13g2_decap_8 FILLER_43_1069 ();
 sg13g2_decap_8 FILLER_43_1076 ();
 sg13g2_decap_8 FILLER_43_1083 ();
 sg13g2_decap_8 FILLER_43_1090 ();
 sg13g2_decap_8 FILLER_43_1097 ();
 sg13g2_decap_8 FILLER_43_1104 ();
 sg13g2_decap_8 FILLER_43_1111 ();
 sg13g2_decap_8 FILLER_43_1118 ();
 sg13g2_decap_8 FILLER_43_1125 ();
 sg13g2_decap_8 FILLER_43_1132 ();
 sg13g2_decap_8 FILLER_43_1139 ();
 sg13g2_decap_8 FILLER_43_1146 ();
 sg13g2_decap_8 FILLER_43_1153 ();
 sg13g2_decap_8 FILLER_43_1160 ();
 sg13g2_decap_8 FILLER_43_1167 ();
 sg13g2_decap_8 FILLER_43_1174 ();
 sg13g2_decap_8 FILLER_43_1181 ();
 sg13g2_decap_8 FILLER_43_1188 ();
 sg13g2_decap_8 FILLER_43_1195 ();
 sg13g2_decap_8 FILLER_43_1202 ();
 sg13g2_decap_8 FILLER_43_1209 ();
 sg13g2_decap_8 FILLER_43_1216 ();
 sg13g2_decap_8 FILLER_43_1223 ();
 sg13g2_decap_8 FILLER_43_1230 ();
 sg13g2_decap_8 FILLER_43_1237 ();
 sg13g2_decap_8 FILLER_43_1244 ();
 sg13g2_decap_8 FILLER_43_1251 ();
 sg13g2_decap_8 FILLER_43_1258 ();
 sg13g2_decap_8 FILLER_43_1265 ();
 sg13g2_decap_8 FILLER_43_1272 ();
 sg13g2_decap_8 FILLER_43_1279 ();
 sg13g2_decap_8 FILLER_43_1286 ();
 sg13g2_decap_8 FILLER_43_1293 ();
 sg13g2_decap_8 FILLER_43_1300 ();
 sg13g2_decap_8 FILLER_43_1307 ();
 sg13g2_decap_8 FILLER_43_1314 ();
 sg13g2_decap_8 FILLER_43_1321 ();
 sg13g2_decap_8 FILLER_43_1328 ();
 sg13g2_decap_8 FILLER_43_1335 ();
 sg13g2_decap_8 FILLER_43_1342 ();
 sg13g2_decap_8 FILLER_43_1349 ();
 sg13g2_decap_8 FILLER_43_1356 ();
 sg13g2_decap_8 FILLER_43_1363 ();
 sg13g2_decap_8 FILLER_43_1370 ();
 sg13g2_decap_8 FILLER_43_1377 ();
 sg13g2_decap_8 FILLER_43_1384 ();
 sg13g2_decap_8 FILLER_43_1391 ();
 sg13g2_decap_8 FILLER_43_1398 ();
 sg13g2_decap_8 FILLER_43_1405 ();
 sg13g2_decap_8 FILLER_43_1412 ();
 sg13g2_decap_8 FILLER_43_1419 ();
 sg13g2_decap_8 FILLER_43_1426 ();
 sg13g2_decap_8 FILLER_43_1433 ();
 sg13g2_decap_8 FILLER_43_1440 ();
 sg13g2_decap_8 FILLER_43_1447 ();
 sg13g2_decap_8 FILLER_43_1454 ();
 sg13g2_decap_8 FILLER_43_1461 ();
 sg13g2_decap_8 FILLER_43_1468 ();
 sg13g2_decap_8 FILLER_43_1475 ();
 sg13g2_decap_8 FILLER_43_1482 ();
 sg13g2_decap_8 FILLER_43_1489 ();
 sg13g2_decap_8 FILLER_43_1496 ();
 sg13g2_decap_8 FILLER_43_1503 ();
 sg13g2_decap_8 FILLER_43_1510 ();
 sg13g2_decap_8 FILLER_43_1517 ();
 sg13g2_decap_8 FILLER_43_1524 ();
 sg13g2_decap_8 FILLER_43_1531 ();
 sg13g2_decap_8 FILLER_43_1538 ();
 sg13g2_decap_8 FILLER_43_1545 ();
 sg13g2_decap_8 FILLER_43_1552 ();
 sg13g2_decap_8 FILLER_43_1559 ();
 sg13g2_decap_8 FILLER_43_1566 ();
 sg13g2_decap_8 FILLER_43_1573 ();
 sg13g2_decap_8 FILLER_43_1580 ();
 sg13g2_decap_8 FILLER_43_1587 ();
 sg13g2_decap_8 FILLER_43_1594 ();
 sg13g2_decap_8 FILLER_43_1601 ();
 sg13g2_decap_8 FILLER_43_1608 ();
 sg13g2_decap_8 FILLER_43_1615 ();
 sg13g2_decap_8 FILLER_43_1622 ();
 sg13g2_decap_8 FILLER_43_1629 ();
 sg13g2_decap_8 FILLER_43_1636 ();
 sg13g2_decap_8 FILLER_43_1643 ();
 sg13g2_decap_8 FILLER_43_1650 ();
 sg13g2_decap_8 FILLER_43_1657 ();
 sg13g2_decap_8 FILLER_43_1664 ();
 sg13g2_decap_8 FILLER_43_1671 ();
 sg13g2_decap_8 FILLER_43_1678 ();
 sg13g2_decap_8 FILLER_43_1685 ();
 sg13g2_decap_8 FILLER_43_1692 ();
 sg13g2_decap_8 FILLER_43_1699 ();
 sg13g2_decap_8 FILLER_43_1706 ();
 sg13g2_decap_8 FILLER_43_1713 ();
 sg13g2_decap_8 FILLER_43_1720 ();
 sg13g2_decap_8 FILLER_43_1727 ();
 sg13g2_decap_8 FILLER_43_1734 ();
 sg13g2_decap_8 FILLER_43_1741 ();
 sg13g2_decap_8 FILLER_43_1748 ();
 sg13g2_decap_8 FILLER_43_1755 ();
 sg13g2_decap_4 FILLER_43_1762 ();
 sg13g2_fill_2 FILLER_43_1766 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_decap_8 FILLER_44_14 ();
 sg13g2_decap_8 FILLER_44_21 ();
 sg13g2_decap_8 FILLER_44_28 ();
 sg13g2_decap_8 FILLER_44_35 ();
 sg13g2_decap_8 FILLER_44_42 ();
 sg13g2_decap_8 FILLER_44_49 ();
 sg13g2_decap_8 FILLER_44_56 ();
 sg13g2_decap_8 FILLER_44_63 ();
 sg13g2_decap_8 FILLER_44_70 ();
 sg13g2_decap_8 FILLER_44_77 ();
 sg13g2_decap_8 FILLER_44_84 ();
 sg13g2_decap_8 FILLER_44_91 ();
 sg13g2_decap_8 FILLER_44_98 ();
 sg13g2_decap_8 FILLER_44_105 ();
 sg13g2_decap_8 FILLER_44_112 ();
 sg13g2_decap_8 FILLER_44_119 ();
 sg13g2_decap_8 FILLER_44_126 ();
 sg13g2_decap_8 FILLER_44_133 ();
 sg13g2_decap_8 FILLER_44_140 ();
 sg13g2_decap_8 FILLER_44_147 ();
 sg13g2_decap_8 FILLER_44_154 ();
 sg13g2_decap_8 FILLER_44_161 ();
 sg13g2_decap_8 FILLER_44_168 ();
 sg13g2_fill_2 FILLER_44_175 ();
 sg13g2_decap_8 FILLER_44_207 ();
 sg13g2_fill_1 FILLER_44_248 ();
 sg13g2_decap_8 FILLER_44_311 ();
 sg13g2_decap_8 FILLER_44_318 ();
 sg13g2_decap_4 FILLER_44_325 ();
 sg13g2_fill_1 FILLER_44_364 ();
 sg13g2_fill_2 FILLER_44_370 ();
 sg13g2_decap_8 FILLER_44_394 ();
 sg13g2_fill_2 FILLER_44_401 ();
 sg13g2_fill_1 FILLER_44_403 ();
 sg13g2_fill_2 FILLER_44_409 ();
 sg13g2_fill_1 FILLER_44_411 ();
 sg13g2_decap_8 FILLER_44_424 ();
 sg13g2_fill_2 FILLER_44_431 ();
 sg13g2_fill_1 FILLER_44_433 ();
 sg13g2_decap_8 FILLER_44_452 ();
 sg13g2_fill_2 FILLER_44_459 ();
 sg13g2_fill_1 FILLER_44_461 ();
 sg13g2_fill_2 FILLER_44_471 ();
 sg13g2_fill_2 FILLER_44_483 ();
 sg13g2_decap_8 FILLER_44_489 ();
 sg13g2_fill_2 FILLER_44_496 ();
 sg13g2_decap_4 FILLER_44_502 ();
 sg13g2_fill_2 FILLER_44_506 ();
 sg13g2_fill_2 FILLER_44_532 ();
 sg13g2_fill_2 FILLER_44_554 ();
 sg13g2_fill_1 FILLER_44_556 ();
 sg13g2_decap_4 FILLER_44_569 ();
 sg13g2_fill_2 FILLER_44_588 ();
 sg13g2_fill_2 FILLER_44_616 ();
 sg13g2_fill_1 FILLER_44_618 ();
 sg13g2_fill_2 FILLER_44_631 ();
 sg13g2_decap_8 FILLER_44_642 ();
 sg13g2_decap_8 FILLER_44_649 ();
 sg13g2_decap_4 FILLER_44_656 ();
 sg13g2_fill_1 FILLER_44_660 ();
 sg13g2_decap_4 FILLER_44_672 ();
 sg13g2_decap_8 FILLER_44_695 ();
 sg13g2_decap_8 FILLER_44_716 ();
 sg13g2_fill_2 FILLER_44_732 ();
 sg13g2_fill_1 FILLER_44_741 ();
 sg13g2_decap_8 FILLER_44_747 ();
 sg13g2_decap_8 FILLER_44_754 ();
 sg13g2_fill_2 FILLER_44_761 ();
 sg13g2_decap_8 FILLER_44_789 ();
 sg13g2_fill_2 FILLER_44_796 ();
 sg13g2_fill_1 FILLER_44_798 ();
 sg13g2_decap_4 FILLER_44_833 ();
 sg13g2_fill_1 FILLER_44_837 ();
 sg13g2_fill_2 FILLER_44_845 ();
 sg13g2_fill_1 FILLER_44_857 ();
 sg13g2_fill_2 FILLER_44_863 ();
 sg13g2_fill_1 FILLER_44_888 ();
 sg13g2_fill_1 FILLER_44_898 ();
 sg13g2_fill_2 FILLER_44_918 ();
 sg13g2_decap_4 FILLER_44_942 ();
 sg13g2_decap_4 FILLER_44_978 ();
 sg13g2_fill_1 FILLER_44_982 ();
 sg13g2_decap_8 FILLER_44_987 ();
 sg13g2_decap_8 FILLER_44_994 ();
 sg13g2_decap_8 FILLER_44_1001 ();
 sg13g2_decap_8 FILLER_44_1008 ();
 sg13g2_fill_2 FILLER_44_1028 ();
 sg13g2_decap_8 FILLER_44_1039 ();
 sg13g2_decap_8 FILLER_44_1046 ();
 sg13g2_decap_8 FILLER_44_1053 ();
 sg13g2_decap_8 FILLER_44_1060 ();
 sg13g2_decap_8 FILLER_44_1067 ();
 sg13g2_decap_8 FILLER_44_1074 ();
 sg13g2_decap_8 FILLER_44_1081 ();
 sg13g2_decap_8 FILLER_44_1088 ();
 sg13g2_decap_8 FILLER_44_1095 ();
 sg13g2_decap_8 FILLER_44_1102 ();
 sg13g2_decap_8 FILLER_44_1109 ();
 sg13g2_decap_8 FILLER_44_1116 ();
 sg13g2_decap_8 FILLER_44_1123 ();
 sg13g2_decap_8 FILLER_44_1130 ();
 sg13g2_decap_8 FILLER_44_1137 ();
 sg13g2_decap_8 FILLER_44_1144 ();
 sg13g2_decap_8 FILLER_44_1151 ();
 sg13g2_decap_8 FILLER_44_1158 ();
 sg13g2_decap_8 FILLER_44_1165 ();
 sg13g2_decap_8 FILLER_44_1172 ();
 sg13g2_decap_8 FILLER_44_1179 ();
 sg13g2_decap_8 FILLER_44_1186 ();
 sg13g2_decap_8 FILLER_44_1193 ();
 sg13g2_decap_8 FILLER_44_1200 ();
 sg13g2_decap_8 FILLER_44_1207 ();
 sg13g2_decap_8 FILLER_44_1214 ();
 sg13g2_decap_8 FILLER_44_1221 ();
 sg13g2_decap_8 FILLER_44_1228 ();
 sg13g2_decap_8 FILLER_44_1235 ();
 sg13g2_decap_8 FILLER_44_1242 ();
 sg13g2_decap_8 FILLER_44_1249 ();
 sg13g2_decap_8 FILLER_44_1256 ();
 sg13g2_decap_8 FILLER_44_1263 ();
 sg13g2_decap_8 FILLER_44_1270 ();
 sg13g2_decap_8 FILLER_44_1277 ();
 sg13g2_decap_8 FILLER_44_1284 ();
 sg13g2_decap_8 FILLER_44_1291 ();
 sg13g2_decap_8 FILLER_44_1298 ();
 sg13g2_decap_8 FILLER_44_1305 ();
 sg13g2_decap_8 FILLER_44_1312 ();
 sg13g2_decap_8 FILLER_44_1319 ();
 sg13g2_decap_8 FILLER_44_1326 ();
 sg13g2_decap_8 FILLER_44_1333 ();
 sg13g2_decap_8 FILLER_44_1340 ();
 sg13g2_decap_8 FILLER_44_1347 ();
 sg13g2_decap_8 FILLER_44_1354 ();
 sg13g2_decap_8 FILLER_44_1361 ();
 sg13g2_decap_8 FILLER_44_1368 ();
 sg13g2_decap_8 FILLER_44_1375 ();
 sg13g2_decap_8 FILLER_44_1382 ();
 sg13g2_decap_8 FILLER_44_1389 ();
 sg13g2_decap_8 FILLER_44_1396 ();
 sg13g2_decap_8 FILLER_44_1403 ();
 sg13g2_decap_8 FILLER_44_1410 ();
 sg13g2_decap_8 FILLER_44_1417 ();
 sg13g2_decap_8 FILLER_44_1424 ();
 sg13g2_decap_8 FILLER_44_1431 ();
 sg13g2_decap_8 FILLER_44_1438 ();
 sg13g2_decap_8 FILLER_44_1445 ();
 sg13g2_decap_8 FILLER_44_1452 ();
 sg13g2_decap_8 FILLER_44_1459 ();
 sg13g2_decap_8 FILLER_44_1466 ();
 sg13g2_decap_8 FILLER_44_1473 ();
 sg13g2_decap_8 FILLER_44_1480 ();
 sg13g2_decap_8 FILLER_44_1487 ();
 sg13g2_decap_8 FILLER_44_1494 ();
 sg13g2_decap_8 FILLER_44_1501 ();
 sg13g2_decap_8 FILLER_44_1508 ();
 sg13g2_decap_8 FILLER_44_1515 ();
 sg13g2_decap_8 FILLER_44_1522 ();
 sg13g2_decap_8 FILLER_44_1529 ();
 sg13g2_decap_8 FILLER_44_1536 ();
 sg13g2_decap_8 FILLER_44_1543 ();
 sg13g2_decap_8 FILLER_44_1550 ();
 sg13g2_decap_8 FILLER_44_1557 ();
 sg13g2_decap_8 FILLER_44_1564 ();
 sg13g2_decap_8 FILLER_44_1571 ();
 sg13g2_decap_8 FILLER_44_1578 ();
 sg13g2_decap_8 FILLER_44_1585 ();
 sg13g2_decap_8 FILLER_44_1592 ();
 sg13g2_decap_8 FILLER_44_1599 ();
 sg13g2_decap_8 FILLER_44_1606 ();
 sg13g2_decap_8 FILLER_44_1613 ();
 sg13g2_decap_8 FILLER_44_1620 ();
 sg13g2_decap_8 FILLER_44_1627 ();
 sg13g2_decap_8 FILLER_44_1634 ();
 sg13g2_decap_8 FILLER_44_1641 ();
 sg13g2_decap_8 FILLER_44_1648 ();
 sg13g2_decap_8 FILLER_44_1655 ();
 sg13g2_decap_8 FILLER_44_1662 ();
 sg13g2_decap_8 FILLER_44_1669 ();
 sg13g2_decap_8 FILLER_44_1676 ();
 sg13g2_decap_8 FILLER_44_1683 ();
 sg13g2_decap_8 FILLER_44_1690 ();
 sg13g2_decap_8 FILLER_44_1697 ();
 sg13g2_decap_8 FILLER_44_1704 ();
 sg13g2_decap_8 FILLER_44_1711 ();
 sg13g2_decap_8 FILLER_44_1718 ();
 sg13g2_decap_8 FILLER_44_1725 ();
 sg13g2_decap_8 FILLER_44_1732 ();
 sg13g2_decap_8 FILLER_44_1739 ();
 sg13g2_decap_8 FILLER_44_1746 ();
 sg13g2_decap_8 FILLER_44_1753 ();
 sg13g2_decap_8 FILLER_44_1760 ();
 sg13g2_fill_1 FILLER_44_1767 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_7 ();
 sg13g2_decap_8 FILLER_45_14 ();
 sg13g2_decap_8 FILLER_45_21 ();
 sg13g2_decap_8 FILLER_45_28 ();
 sg13g2_decap_8 FILLER_45_35 ();
 sg13g2_decap_8 FILLER_45_42 ();
 sg13g2_decap_8 FILLER_45_49 ();
 sg13g2_decap_8 FILLER_45_56 ();
 sg13g2_decap_8 FILLER_45_63 ();
 sg13g2_decap_8 FILLER_45_70 ();
 sg13g2_decap_8 FILLER_45_77 ();
 sg13g2_decap_8 FILLER_45_84 ();
 sg13g2_decap_8 FILLER_45_91 ();
 sg13g2_decap_8 FILLER_45_98 ();
 sg13g2_decap_8 FILLER_45_105 ();
 sg13g2_decap_8 FILLER_45_112 ();
 sg13g2_decap_8 FILLER_45_119 ();
 sg13g2_decap_8 FILLER_45_126 ();
 sg13g2_decap_8 FILLER_45_133 ();
 sg13g2_decap_8 FILLER_45_140 ();
 sg13g2_fill_1 FILLER_45_147 ();
 sg13g2_decap_4 FILLER_45_158 ();
 sg13g2_fill_1 FILLER_45_162 ();
 sg13g2_decap_4 FILLER_45_210 ();
 sg13g2_fill_1 FILLER_45_214 ();
 sg13g2_fill_1 FILLER_45_256 ();
 sg13g2_fill_1 FILLER_45_266 ();
 sg13g2_decap_8 FILLER_45_308 ();
 sg13g2_decap_8 FILLER_45_318 ();
 sg13g2_decap_4 FILLER_45_325 ();
 sg13g2_fill_2 FILLER_45_329 ();
 sg13g2_fill_1 FILLER_45_358 ();
 sg13g2_decap_8 FILLER_45_362 ();
 sg13g2_decap_4 FILLER_45_369 ();
 sg13g2_fill_1 FILLER_45_373 ();
 sg13g2_fill_2 FILLER_45_395 ();
 sg13g2_fill_2 FILLER_45_426 ();
 sg13g2_fill_1 FILLER_45_428 ();
 sg13g2_fill_2 FILLER_45_451 ();
 sg13g2_fill_1 FILLER_45_453 ();
 sg13g2_fill_1 FILLER_45_473 ();
 sg13g2_fill_1 FILLER_45_482 ();
 sg13g2_fill_2 FILLER_45_489 ();
 sg13g2_decap_8 FILLER_45_504 ();
 sg13g2_decap_8 FILLER_45_511 ();
 sg13g2_decap_8 FILLER_45_535 ();
 sg13g2_fill_2 FILLER_45_542 ();
 sg13g2_fill_1 FILLER_45_544 ();
 sg13g2_fill_1 FILLER_45_565 ();
 sg13g2_decap_8 FILLER_45_607 ();
 sg13g2_decap_8 FILLER_45_619 ();
 sg13g2_decap_4 FILLER_45_635 ();
 sg13g2_fill_1 FILLER_45_639 ();
 sg13g2_fill_2 FILLER_45_663 ();
 sg13g2_fill_2 FILLER_45_676 ();
 sg13g2_fill_1 FILLER_45_682 ();
 sg13g2_fill_1 FILLER_45_700 ();
 sg13g2_fill_1 FILLER_45_715 ();
 sg13g2_fill_2 FILLER_45_732 ();
 sg13g2_fill_1 FILLER_45_734 ();
 sg13g2_decap_8 FILLER_45_756 ();
 sg13g2_decap_8 FILLER_45_763 ();
 sg13g2_decap_4 FILLER_45_770 ();
 sg13g2_fill_1 FILLER_45_774 ();
 sg13g2_decap_4 FILLER_45_787 ();
 sg13g2_decap_8 FILLER_45_796 ();
 sg13g2_decap_4 FILLER_45_822 ();
 sg13g2_decap_8 FILLER_45_831 ();
 sg13g2_decap_8 FILLER_45_882 ();
 sg13g2_decap_4 FILLER_45_889 ();
 sg13g2_fill_2 FILLER_45_893 ();
 sg13g2_fill_1 FILLER_45_899 ();
 sg13g2_fill_1 FILLER_45_904 ();
 sg13g2_fill_1 FILLER_45_910 ();
 sg13g2_decap_4 FILLER_45_916 ();
 sg13g2_fill_2 FILLER_45_920 ();
 sg13g2_fill_2 FILLER_45_948 ();
 sg13g2_fill_1 FILLER_45_972 ();
 sg13g2_fill_2 FILLER_45_981 ();
 sg13g2_decap_8 FILLER_45_996 ();
 sg13g2_fill_2 FILLER_45_1003 ();
 sg13g2_decap_8 FILLER_45_1012 ();
 sg13g2_decap_8 FILLER_45_1019 ();
 sg13g2_decap_8 FILLER_45_1026 ();
 sg13g2_decap_8 FILLER_45_1033 ();
 sg13g2_decap_8 FILLER_45_1040 ();
 sg13g2_decap_8 FILLER_45_1047 ();
 sg13g2_decap_8 FILLER_45_1054 ();
 sg13g2_decap_8 FILLER_45_1061 ();
 sg13g2_decap_8 FILLER_45_1068 ();
 sg13g2_decap_8 FILLER_45_1075 ();
 sg13g2_decap_8 FILLER_45_1082 ();
 sg13g2_decap_8 FILLER_45_1089 ();
 sg13g2_decap_8 FILLER_45_1096 ();
 sg13g2_decap_8 FILLER_45_1103 ();
 sg13g2_decap_8 FILLER_45_1110 ();
 sg13g2_decap_8 FILLER_45_1117 ();
 sg13g2_decap_8 FILLER_45_1124 ();
 sg13g2_decap_8 FILLER_45_1131 ();
 sg13g2_decap_8 FILLER_45_1138 ();
 sg13g2_decap_8 FILLER_45_1145 ();
 sg13g2_decap_8 FILLER_45_1152 ();
 sg13g2_decap_8 FILLER_45_1159 ();
 sg13g2_decap_8 FILLER_45_1166 ();
 sg13g2_decap_8 FILLER_45_1173 ();
 sg13g2_decap_8 FILLER_45_1180 ();
 sg13g2_decap_8 FILLER_45_1187 ();
 sg13g2_decap_8 FILLER_45_1194 ();
 sg13g2_decap_8 FILLER_45_1201 ();
 sg13g2_decap_8 FILLER_45_1208 ();
 sg13g2_decap_8 FILLER_45_1215 ();
 sg13g2_decap_8 FILLER_45_1222 ();
 sg13g2_decap_8 FILLER_45_1229 ();
 sg13g2_decap_8 FILLER_45_1236 ();
 sg13g2_decap_8 FILLER_45_1243 ();
 sg13g2_decap_8 FILLER_45_1250 ();
 sg13g2_decap_8 FILLER_45_1257 ();
 sg13g2_decap_8 FILLER_45_1264 ();
 sg13g2_decap_8 FILLER_45_1271 ();
 sg13g2_decap_8 FILLER_45_1278 ();
 sg13g2_decap_8 FILLER_45_1285 ();
 sg13g2_decap_8 FILLER_45_1292 ();
 sg13g2_decap_8 FILLER_45_1299 ();
 sg13g2_decap_8 FILLER_45_1306 ();
 sg13g2_decap_8 FILLER_45_1313 ();
 sg13g2_decap_8 FILLER_45_1320 ();
 sg13g2_decap_8 FILLER_45_1327 ();
 sg13g2_decap_8 FILLER_45_1334 ();
 sg13g2_decap_8 FILLER_45_1341 ();
 sg13g2_decap_8 FILLER_45_1348 ();
 sg13g2_decap_8 FILLER_45_1355 ();
 sg13g2_decap_8 FILLER_45_1362 ();
 sg13g2_decap_8 FILLER_45_1369 ();
 sg13g2_decap_8 FILLER_45_1376 ();
 sg13g2_decap_8 FILLER_45_1383 ();
 sg13g2_decap_8 FILLER_45_1390 ();
 sg13g2_decap_8 FILLER_45_1397 ();
 sg13g2_decap_8 FILLER_45_1404 ();
 sg13g2_decap_8 FILLER_45_1411 ();
 sg13g2_decap_8 FILLER_45_1418 ();
 sg13g2_decap_8 FILLER_45_1425 ();
 sg13g2_decap_8 FILLER_45_1432 ();
 sg13g2_decap_8 FILLER_45_1439 ();
 sg13g2_decap_8 FILLER_45_1446 ();
 sg13g2_decap_8 FILLER_45_1453 ();
 sg13g2_decap_8 FILLER_45_1460 ();
 sg13g2_decap_8 FILLER_45_1467 ();
 sg13g2_decap_8 FILLER_45_1474 ();
 sg13g2_decap_8 FILLER_45_1481 ();
 sg13g2_decap_8 FILLER_45_1488 ();
 sg13g2_decap_8 FILLER_45_1495 ();
 sg13g2_decap_8 FILLER_45_1502 ();
 sg13g2_decap_8 FILLER_45_1509 ();
 sg13g2_decap_8 FILLER_45_1516 ();
 sg13g2_decap_8 FILLER_45_1523 ();
 sg13g2_decap_8 FILLER_45_1530 ();
 sg13g2_decap_8 FILLER_45_1537 ();
 sg13g2_decap_8 FILLER_45_1544 ();
 sg13g2_decap_8 FILLER_45_1551 ();
 sg13g2_decap_8 FILLER_45_1558 ();
 sg13g2_decap_8 FILLER_45_1565 ();
 sg13g2_decap_8 FILLER_45_1572 ();
 sg13g2_decap_8 FILLER_45_1579 ();
 sg13g2_decap_8 FILLER_45_1586 ();
 sg13g2_decap_8 FILLER_45_1593 ();
 sg13g2_decap_8 FILLER_45_1600 ();
 sg13g2_decap_8 FILLER_45_1607 ();
 sg13g2_decap_8 FILLER_45_1614 ();
 sg13g2_decap_8 FILLER_45_1621 ();
 sg13g2_decap_8 FILLER_45_1628 ();
 sg13g2_decap_8 FILLER_45_1635 ();
 sg13g2_decap_8 FILLER_45_1642 ();
 sg13g2_decap_8 FILLER_45_1649 ();
 sg13g2_decap_8 FILLER_45_1656 ();
 sg13g2_decap_8 FILLER_45_1663 ();
 sg13g2_decap_8 FILLER_45_1670 ();
 sg13g2_decap_8 FILLER_45_1677 ();
 sg13g2_decap_8 FILLER_45_1684 ();
 sg13g2_decap_8 FILLER_45_1691 ();
 sg13g2_decap_8 FILLER_45_1698 ();
 sg13g2_decap_8 FILLER_45_1705 ();
 sg13g2_decap_8 FILLER_45_1712 ();
 sg13g2_decap_8 FILLER_45_1719 ();
 sg13g2_decap_8 FILLER_45_1726 ();
 sg13g2_decap_8 FILLER_45_1733 ();
 sg13g2_decap_8 FILLER_45_1740 ();
 sg13g2_decap_8 FILLER_45_1747 ();
 sg13g2_decap_8 FILLER_45_1754 ();
 sg13g2_decap_8 FILLER_45_1761 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_7 ();
 sg13g2_decap_8 FILLER_46_14 ();
 sg13g2_decap_8 FILLER_46_21 ();
 sg13g2_decap_8 FILLER_46_28 ();
 sg13g2_decap_8 FILLER_46_35 ();
 sg13g2_decap_8 FILLER_46_42 ();
 sg13g2_decap_8 FILLER_46_49 ();
 sg13g2_decap_8 FILLER_46_56 ();
 sg13g2_decap_8 FILLER_46_63 ();
 sg13g2_decap_8 FILLER_46_70 ();
 sg13g2_decap_8 FILLER_46_77 ();
 sg13g2_decap_8 FILLER_46_84 ();
 sg13g2_decap_8 FILLER_46_91 ();
 sg13g2_fill_2 FILLER_46_98 ();
 sg13g2_fill_1 FILLER_46_100 ();
 sg13g2_decap_4 FILLER_46_104 ();
 sg13g2_fill_2 FILLER_46_108 ();
 sg13g2_decap_4 FILLER_46_115 ();
 sg13g2_fill_1 FILLER_46_119 ();
 sg13g2_decap_8 FILLER_46_124 ();
 sg13g2_decap_8 FILLER_46_140 ();
 sg13g2_fill_1 FILLER_46_176 ();
 sg13g2_fill_1 FILLER_46_180 ();
 sg13g2_fill_2 FILLER_46_268 ();
 sg13g2_decap_4 FILLER_46_305 ();
 sg13g2_fill_1 FILLER_46_309 ();
 sg13g2_fill_2 FILLER_46_336 ();
 sg13g2_fill_2 FILLER_46_364 ();
 sg13g2_decap_4 FILLER_46_386 ();
 sg13g2_fill_1 FILLER_46_400 ();
 sg13g2_decap_4 FILLER_46_410 ();
 sg13g2_fill_1 FILLER_46_414 ();
 sg13g2_decap_4 FILLER_46_420 ();
 sg13g2_fill_1 FILLER_46_424 ();
 sg13g2_fill_1 FILLER_46_469 ();
 sg13g2_fill_1 FILLER_46_475 ();
 sg13g2_fill_2 FILLER_46_481 ();
 sg13g2_fill_1 FILLER_46_506 ();
 sg13g2_decap_8 FILLER_46_530 ();
 sg13g2_fill_2 FILLER_46_537 ();
 sg13g2_fill_2 FILLER_46_561 ();
 sg13g2_decap_8 FILLER_46_568 ();
 sg13g2_fill_1 FILLER_46_575 ();
 sg13g2_decap_4 FILLER_46_581 ();
 sg13g2_fill_1 FILLER_46_585 ();
 sg13g2_fill_1 FILLER_46_615 ();
 sg13g2_decap_8 FILLER_46_643 ();
 sg13g2_decap_8 FILLER_46_650 ();
 sg13g2_fill_2 FILLER_46_657 ();
 sg13g2_fill_1 FILLER_46_663 ();
 sg13g2_decap_4 FILLER_46_675 ();
 sg13g2_fill_1 FILLER_46_679 ();
 sg13g2_fill_2 FILLER_46_697 ();
 sg13g2_fill_2 FILLER_46_709 ();
 sg13g2_fill_2 FILLER_46_717 ();
 sg13g2_fill_1 FILLER_46_719 ();
 sg13g2_decap_4 FILLER_46_732 ();
 sg13g2_fill_1 FILLER_46_736 ();
 sg13g2_fill_2 FILLER_46_742 ();
 sg13g2_fill_1 FILLER_46_744 ();
 sg13g2_decap_4 FILLER_46_762 ();
 sg13g2_fill_2 FILLER_46_771 ();
 sg13g2_decap_4 FILLER_46_790 ();
 sg13g2_fill_2 FILLER_46_794 ();
 sg13g2_fill_2 FILLER_46_800 ();
 sg13g2_decap_8 FILLER_46_817 ();
 sg13g2_fill_1 FILLER_46_824 ();
 sg13g2_fill_1 FILLER_46_829 ();
 sg13g2_fill_2 FILLER_46_846 ();
 sg13g2_decap_8 FILLER_46_857 ();
 sg13g2_fill_1 FILLER_46_864 ();
 sg13g2_fill_2 FILLER_46_888 ();
 sg13g2_fill_1 FILLER_46_890 ();
 sg13g2_fill_2 FILLER_46_899 ();
 sg13g2_fill_1 FILLER_46_901 ();
 sg13g2_fill_1 FILLER_46_915 ();
 sg13g2_fill_2 FILLER_46_947 ();
 sg13g2_fill_2 FILLER_46_975 ();
 sg13g2_fill_2 FILLER_46_1003 ();
 sg13g2_decap_8 FILLER_46_1045 ();
 sg13g2_decap_8 FILLER_46_1052 ();
 sg13g2_decap_8 FILLER_46_1059 ();
 sg13g2_decap_8 FILLER_46_1066 ();
 sg13g2_decap_8 FILLER_46_1073 ();
 sg13g2_decap_8 FILLER_46_1080 ();
 sg13g2_decap_8 FILLER_46_1087 ();
 sg13g2_decap_8 FILLER_46_1094 ();
 sg13g2_decap_8 FILLER_46_1101 ();
 sg13g2_decap_8 FILLER_46_1108 ();
 sg13g2_decap_8 FILLER_46_1115 ();
 sg13g2_decap_8 FILLER_46_1122 ();
 sg13g2_decap_8 FILLER_46_1129 ();
 sg13g2_decap_8 FILLER_46_1136 ();
 sg13g2_decap_8 FILLER_46_1143 ();
 sg13g2_decap_8 FILLER_46_1150 ();
 sg13g2_decap_8 FILLER_46_1157 ();
 sg13g2_decap_8 FILLER_46_1164 ();
 sg13g2_decap_8 FILLER_46_1171 ();
 sg13g2_decap_8 FILLER_46_1178 ();
 sg13g2_decap_8 FILLER_46_1185 ();
 sg13g2_decap_8 FILLER_46_1192 ();
 sg13g2_decap_8 FILLER_46_1199 ();
 sg13g2_decap_8 FILLER_46_1206 ();
 sg13g2_decap_8 FILLER_46_1213 ();
 sg13g2_decap_8 FILLER_46_1220 ();
 sg13g2_decap_8 FILLER_46_1227 ();
 sg13g2_decap_8 FILLER_46_1234 ();
 sg13g2_decap_8 FILLER_46_1241 ();
 sg13g2_decap_8 FILLER_46_1248 ();
 sg13g2_decap_8 FILLER_46_1255 ();
 sg13g2_decap_8 FILLER_46_1262 ();
 sg13g2_decap_8 FILLER_46_1269 ();
 sg13g2_decap_8 FILLER_46_1276 ();
 sg13g2_decap_8 FILLER_46_1283 ();
 sg13g2_decap_8 FILLER_46_1290 ();
 sg13g2_decap_8 FILLER_46_1297 ();
 sg13g2_decap_8 FILLER_46_1304 ();
 sg13g2_decap_8 FILLER_46_1311 ();
 sg13g2_decap_8 FILLER_46_1318 ();
 sg13g2_decap_8 FILLER_46_1325 ();
 sg13g2_decap_8 FILLER_46_1332 ();
 sg13g2_decap_8 FILLER_46_1339 ();
 sg13g2_decap_8 FILLER_46_1346 ();
 sg13g2_decap_8 FILLER_46_1353 ();
 sg13g2_decap_8 FILLER_46_1360 ();
 sg13g2_decap_8 FILLER_46_1367 ();
 sg13g2_decap_8 FILLER_46_1374 ();
 sg13g2_decap_8 FILLER_46_1381 ();
 sg13g2_decap_8 FILLER_46_1388 ();
 sg13g2_decap_8 FILLER_46_1395 ();
 sg13g2_decap_8 FILLER_46_1402 ();
 sg13g2_decap_8 FILLER_46_1409 ();
 sg13g2_decap_8 FILLER_46_1416 ();
 sg13g2_decap_8 FILLER_46_1423 ();
 sg13g2_decap_8 FILLER_46_1430 ();
 sg13g2_decap_8 FILLER_46_1437 ();
 sg13g2_decap_8 FILLER_46_1444 ();
 sg13g2_decap_8 FILLER_46_1451 ();
 sg13g2_decap_8 FILLER_46_1458 ();
 sg13g2_decap_8 FILLER_46_1465 ();
 sg13g2_decap_8 FILLER_46_1472 ();
 sg13g2_decap_8 FILLER_46_1479 ();
 sg13g2_decap_8 FILLER_46_1486 ();
 sg13g2_decap_8 FILLER_46_1493 ();
 sg13g2_decap_8 FILLER_46_1500 ();
 sg13g2_decap_8 FILLER_46_1507 ();
 sg13g2_decap_8 FILLER_46_1514 ();
 sg13g2_decap_8 FILLER_46_1521 ();
 sg13g2_decap_8 FILLER_46_1528 ();
 sg13g2_decap_8 FILLER_46_1535 ();
 sg13g2_decap_8 FILLER_46_1542 ();
 sg13g2_decap_8 FILLER_46_1549 ();
 sg13g2_decap_8 FILLER_46_1556 ();
 sg13g2_decap_8 FILLER_46_1563 ();
 sg13g2_decap_8 FILLER_46_1570 ();
 sg13g2_decap_8 FILLER_46_1577 ();
 sg13g2_decap_8 FILLER_46_1584 ();
 sg13g2_decap_8 FILLER_46_1591 ();
 sg13g2_decap_8 FILLER_46_1598 ();
 sg13g2_decap_8 FILLER_46_1605 ();
 sg13g2_decap_8 FILLER_46_1612 ();
 sg13g2_decap_8 FILLER_46_1619 ();
 sg13g2_decap_8 FILLER_46_1626 ();
 sg13g2_decap_8 FILLER_46_1633 ();
 sg13g2_decap_8 FILLER_46_1640 ();
 sg13g2_decap_8 FILLER_46_1647 ();
 sg13g2_decap_8 FILLER_46_1654 ();
 sg13g2_decap_8 FILLER_46_1661 ();
 sg13g2_decap_8 FILLER_46_1668 ();
 sg13g2_decap_8 FILLER_46_1675 ();
 sg13g2_decap_8 FILLER_46_1682 ();
 sg13g2_decap_8 FILLER_46_1689 ();
 sg13g2_decap_8 FILLER_46_1696 ();
 sg13g2_decap_8 FILLER_46_1703 ();
 sg13g2_decap_8 FILLER_46_1710 ();
 sg13g2_decap_8 FILLER_46_1717 ();
 sg13g2_decap_8 FILLER_46_1724 ();
 sg13g2_decap_8 FILLER_46_1731 ();
 sg13g2_decap_8 FILLER_46_1738 ();
 sg13g2_decap_8 FILLER_46_1745 ();
 sg13g2_decap_8 FILLER_46_1752 ();
 sg13g2_decap_8 FILLER_46_1759 ();
 sg13g2_fill_2 FILLER_46_1766 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_7 ();
 sg13g2_decap_8 FILLER_47_14 ();
 sg13g2_decap_8 FILLER_47_21 ();
 sg13g2_decap_8 FILLER_47_28 ();
 sg13g2_decap_8 FILLER_47_35 ();
 sg13g2_decap_8 FILLER_47_42 ();
 sg13g2_decap_8 FILLER_47_49 ();
 sg13g2_decap_8 FILLER_47_56 ();
 sg13g2_decap_8 FILLER_47_63 ();
 sg13g2_decap_4 FILLER_47_70 ();
 sg13g2_fill_1 FILLER_47_74 ();
 sg13g2_decap_8 FILLER_47_78 ();
 sg13g2_decap_4 FILLER_47_85 ();
 sg13g2_fill_2 FILLER_47_144 ();
 sg13g2_fill_1 FILLER_47_146 ();
 sg13g2_fill_1 FILLER_47_183 ();
 sg13g2_fill_1 FILLER_47_203 ();
 sg13g2_fill_1 FILLER_47_248 ();
 sg13g2_decap_4 FILLER_47_291 ();
 sg13g2_fill_1 FILLER_47_325 ();
 sg13g2_fill_1 FILLER_47_348 ();
 sg13g2_fill_2 FILLER_47_391 ();
 sg13g2_fill_1 FILLER_47_393 ();
 sg13g2_fill_1 FILLER_47_446 ();
 sg13g2_fill_2 FILLER_47_452 ();
 sg13g2_fill_2 FILLER_47_479 ();
 sg13g2_fill_1 FILLER_47_481 ();
 sg13g2_fill_2 FILLER_47_487 ();
 sg13g2_fill_1 FILLER_47_489 ();
 sg13g2_fill_2 FILLER_47_497 ();
 sg13g2_decap_4 FILLER_47_509 ();
 sg13g2_fill_1 FILLER_47_513 ();
 sg13g2_decap_8 FILLER_47_526 ();
 sg13g2_decap_8 FILLER_47_533 ();
 sg13g2_decap_4 FILLER_47_540 ();
 sg13g2_decap_8 FILLER_47_549 ();
 sg13g2_fill_1 FILLER_47_556 ();
 sg13g2_fill_1 FILLER_47_583 ();
 sg13g2_decap_8 FILLER_47_637 ();
 sg13g2_fill_2 FILLER_47_644 ();
 sg13g2_decap_8 FILLER_47_680 ();
 sg13g2_fill_2 FILLER_47_699 ();
 sg13g2_fill_1 FILLER_47_706 ();
 sg13g2_decap_8 FILLER_47_738 ();
 sg13g2_fill_1 FILLER_47_770 ();
 sg13g2_fill_2 FILLER_47_794 ();
 sg13g2_fill_1 FILLER_47_796 ();
 sg13g2_decap_4 FILLER_47_814 ();
 sg13g2_fill_1 FILLER_47_818 ();
 sg13g2_fill_2 FILLER_47_846 ();
 sg13g2_decap_4 FILLER_47_865 ();
 sg13g2_fill_1 FILLER_47_869 ();
 sg13g2_fill_2 FILLER_47_875 ();
 sg13g2_fill_2 FILLER_47_890 ();
 sg13g2_decap_4 FILLER_47_896 ();
 sg13g2_fill_1 FILLER_47_900 ();
 sg13g2_fill_1 FILLER_47_923 ();
 sg13g2_decap_8 FILLER_47_940 ();
 sg13g2_decap_8 FILLER_47_947 ();
 sg13g2_fill_2 FILLER_47_954 ();
 sg13g2_fill_2 FILLER_47_972 ();
 sg13g2_fill_1 FILLER_47_974 ();
 sg13g2_fill_1 FILLER_47_982 ();
 sg13g2_decap_8 FILLER_47_995 ();
 sg13g2_decap_8 FILLER_47_1002 ();
 sg13g2_decap_8 FILLER_47_1009 ();
 sg13g2_decap_8 FILLER_47_1016 ();
 sg13g2_decap_8 FILLER_47_1023 ();
 sg13g2_decap_8 FILLER_47_1030 ();
 sg13g2_decap_8 FILLER_47_1037 ();
 sg13g2_decap_8 FILLER_47_1044 ();
 sg13g2_decap_8 FILLER_47_1051 ();
 sg13g2_decap_8 FILLER_47_1058 ();
 sg13g2_decap_8 FILLER_47_1065 ();
 sg13g2_decap_8 FILLER_47_1072 ();
 sg13g2_decap_8 FILLER_47_1079 ();
 sg13g2_decap_8 FILLER_47_1086 ();
 sg13g2_decap_8 FILLER_47_1093 ();
 sg13g2_decap_8 FILLER_47_1100 ();
 sg13g2_decap_8 FILLER_47_1107 ();
 sg13g2_decap_8 FILLER_47_1114 ();
 sg13g2_decap_8 FILLER_47_1121 ();
 sg13g2_decap_8 FILLER_47_1128 ();
 sg13g2_decap_8 FILLER_47_1135 ();
 sg13g2_decap_8 FILLER_47_1142 ();
 sg13g2_decap_8 FILLER_47_1149 ();
 sg13g2_decap_8 FILLER_47_1156 ();
 sg13g2_decap_8 FILLER_47_1163 ();
 sg13g2_decap_8 FILLER_47_1170 ();
 sg13g2_decap_8 FILLER_47_1177 ();
 sg13g2_decap_8 FILLER_47_1184 ();
 sg13g2_decap_8 FILLER_47_1191 ();
 sg13g2_decap_8 FILLER_47_1198 ();
 sg13g2_decap_8 FILLER_47_1205 ();
 sg13g2_decap_8 FILLER_47_1212 ();
 sg13g2_decap_8 FILLER_47_1219 ();
 sg13g2_decap_8 FILLER_47_1226 ();
 sg13g2_decap_8 FILLER_47_1233 ();
 sg13g2_decap_8 FILLER_47_1240 ();
 sg13g2_decap_8 FILLER_47_1247 ();
 sg13g2_decap_8 FILLER_47_1254 ();
 sg13g2_decap_8 FILLER_47_1261 ();
 sg13g2_decap_8 FILLER_47_1268 ();
 sg13g2_decap_8 FILLER_47_1275 ();
 sg13g2_decap_8 FILLER_47_1282 ();
 sg13g2_decap_8 FILLER_47_1289 ();
 sg13g2_decap_8 FILLER_47_1296 ();
 sg13g2_decap_8 FILLER_47_1303 ();
 sg13g2_decap_8 FILLER_47_1310 ();
 sg13g2_decap_8 FILLER_47_1317 ();
 sg13g2_decap_8 FILLER_47_1324 ();
 sg13g2_decap_8 FILLER_47_1331 ();
 sg13g2_decap_8 FILLER_47_1338 ();
 sg13g2_decap_8 FILLER_47_1345 ();
 sg13g2_decap_8 FILLER_47_1352 ();
 sg13g2_decap_8 FILLER_47_1359 ();
 sg13g2_decap_8 FILLER_47_1366 ();
 sg13g2_decap_8 FILLER_47_1373 ();
 sg13g2_decap_8 FILLER_47_1380 ();
 sg13g2_decap_8 FILLER_47_1387 ();
 sg13g2_decap_8 FILLER_47_1394 ();
 sg13g2_decap_8 FILLER_47_1401 ();
 sg13g2_decap_8 FILLER_47_1408 ();
 sg13g2_decap_8 FILLER_47_1415 ();
 sg13g2_decap_8 FILLER_47_1422 ();
 sg13g2_decap_8 FILLER_47_1429 ();
 sg13g2_decap_8 FILLER_47_1436 ();
 sg13g2_decap_8 FILLER_47_1443 ();
 sg13g2_decap_8 FILLER_47_1450 ();
 sg13g2_decap_8 FILLER_47_1457 ();
 sg13g2_decap_8 FILLER_47_1464 ();
 sg13g2_decap_8 FILLER_47_1471 ();
 sg13g2_decap_8 FILLER_47_1478 ();
 sg13g2_decap_8 FILLER_47_1485 ();
 sg13g2_decap_8 FILLER_47_1492 ();
 sg13g2_decap_8 FILLER_47_1499 ();
 sg13g2_decap_8 FILLER_47_1506 ();
 sg13g2_decap_8 FILLER_47_1513 ();
 sg13g2_decap_8 FILLER_47_1520 ();
 sg13g2_decap_8 FILLER_47_1527 ();
 sg13g2_decap_8 FILLER_47_1534 ();
 sg13g2_decap_8 FILLER_47_1541 ();
 sg13g2_decap_8 FILLER_47_1548 ();
 sg13g2_decap_8 FILLER_47_1555 ();
 sg13g2_decap_8 FILLER_47_1562 ();
 sg13g2_decap_8 FILLER_47_1569 ();
 sg13g2_decap_8 FILLER_47_1576 ();
 sg13g2_decap_8 FILLER_47_1583 ();
 sg13g2_decap_8 FILLER_47_1590 ();
 sg13g2_decap_8 FILLER_47_1597 ();
 sg13g2_decap_8 FILLER_47_1604 ();
 sg13g2_decap_8 FILLER_47_1611 ();
 sg13g2_decap_8 FILLER_47_1618 ();
 sg13g2_decap_8 FILLER_47_1625 ();
 sg13g2_decap_8 FILLER_47_1632 ();
 sg13g2_decap_8 FILLER_47_1639 ();
 sg13g2_decap_8 FILLER_47_1646 ();
 sg13g2_decap_8 FILLER_47_1653 ();
 sg13g2_decap_8 FILLER_47_1660 ();
 sg13g2_decap_8 FILLER_47_1667 ();
 sg13g2_decap_8 FILLER_47_1674 ();
 sg13g2_decap_8 FILLER_47_1681 ();
 sg13g2_decap_8 FILLER_47_1688 ();
 sg13g2_decap_8 FILLER_47_1695 ();
 sg13g2_decap_8 FILLER_47_1702 ();
 sg13g2_decap_8 FILLER_47_1709 ();
 sg13g2_decap_8 FILLER_47_1716 ();
 sg13g2_decap_8 FILLER_47_1723 ();
 sg13g2_decap_8 FILLER_47_1730 ();
 sg13g2_decap_8 FILLER_47_1737 ();
 sg13g2_decap_8 FILLER_47_1744 ();
 sg13g2_decap_8 FILLER_47_1751 ();
 sg13g2_decap_8 FILLER_47_1758 ();
 sg13g2_fill_2 FILLER_47_1765 ();
 sg13g2_fill_1 FILLER_47_1767 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_decap_8 FILLER_48_14 ();
 sg13g2_decap_8 FILLER_48_21 ();
 sg13g2_decap_8 FILLER_48_28 ();
 sg13g2_decap_8 FILLER_48_35 ();
 sg13g2_decap_8 FILLER_48_42 ();
 sg13g2_decap_8 FILLER_48_49 ();
 sg13g2_decap_8 FILLER_48_56 ();
 sg13g2_decap_8 FILLER_48_63 ();
 sg13g2_fill_2 FILLER_48_101 ();
 sg13g2_fill_1 FILLER_48_111 ();
 sg13g2_fill_2 FILLER_48_176 ();
 sg13g2_fill_1 FILLER_48_178 ();
 sg13g2_fill_2 FILLER_48_205 ();
 sg13g2_fill_2 FILLER_48_213 ();
 sg13g2_fill_1 FILLER_48_215 ();
 sg13g2_fill_2 FILLER_48_241 ();
 sg13g2_fill_1 FILLER_48_267 ();
 sg13g2_fill_1 FILLER_48_272 ();
 sg13g2_decap_8 FILLER_48_291 ();
 sg13g2_fill_1 FILLER_48_298 ();
 sg13g2_fill_2 FILLER_48_343 ();
 sg13g2_fill_1 FILLER_48_376 ();
 sg13g2_fill_2 FILLER_48_392 ();
 sg13g2_fill_1 FILLER_48_394 ();
 sg13g2_fill_2 FILLER_48_413 ();
 sg13g2_fill_1 FILLER_48_418 ();
 sg13g2_decap_8 FILLER_48_427 ();
 sg13g2_fill_2 FILLER_48_434 ();
 sg13g2_fill_1 FILLER_48_462 ();
 sg13g2_decap_4 FILLER_48_557 ();
 sg13g2_fill_2 FILLER_48_561 ();
 sg13g2_fill_2 FILLER_48_598 ();
 sg13g2_fill_1 FILLER_48_609 ();
 sg13g2_fill_1 FILLER_48_619 ();
 sg13g2_fill_2 FILLER_48_639 ();
 sg13g2_fill_2 FILLER_48_646 ();
 sg13g2_decap_4 FILLER_48_656 ();
 sg13g2_decap_8 FILLER_48_669 ();
 sg13g2_fill_1 FILLER_48_676 ();
 sg13g2_decap_4 FILLER_48_694 ();
 sg13g2_fill_2 FILLER_48_698 ();
 sg13g2_decap_8 FILLER_48_734 ();
 sg13g2_decap_4 FILLER_48_741 ();
 sg13g2_fill_2 FILLER_48_745 ();
 sg13g2_decap_8 FILLER_48_759 ();
 sg13g2_fill_1 FILLER_48_770 ();
 sg13g2_fill_2 FILLER_48_776 ();
 sg13g2_fill_1 FILLER_48_778 ();
 sg13g2_decap_4 FILLER_48_792 ();
 sg13g2_fill_2 FILLER_48_803 ();
 sg13g2_fill_1 FILLER_48_816 ();
 sg13g2_decap_4 FILLER_48_825 ();
 sg13g2_fill_2 FILLER_48_838 ();
 sg13g2_fill_1 FILLER_48_840 ();
 sg13g2_decap_8 FILLER_48_866 ();
 sg13g2_decap_4 FILLER_48_873 ();
 sg13g2_decap_8 FILLER_48_895 ();
 sg13g2_decap_8 FILLER_48_919 ();
 sg13g2_decap_4 FILLER_48_926 ();
 sg13g2_decap_8 FILLER_48_943 ();
 sg13g2_fill_2 FILLER_48_950 ();
 sg13g2_fill_1 FILLER_48_952 ();
 sg13g2_fill_2 FILLER_48_976 ();
 sg13g2_decap_8 FILLER_48_1007 ();
 sg13g2_decap_8 FILLER_48_1014 ();
 sg13g2_decap_8 FILLER_48_1021 ();
 sg13g2_decap_8 FILLER_48_1028 ();
 sg13g2_decap_8 FILLER_48_1035 ();
 sg13g2_decap_8 FILLER_48_1042 ();
 sg13g2_decap_8 FILLER_48_1049 ();
 sg13g2_decap_8 FILLER_48_1056 ();
 sg13g2_decap_8 FILLER_48_1063 ();
 sg13g2_decap_8 FILLER_48_1070 ();
 sg13g2_decap_8 FILLER_48_1077 ();
 sg13g2_decap_8 FILLER_48_1084 ();
 sg13g2_decap_8 FILLER_48_1091 ();
 sg13g2_decap_8 FILLER_48_1098 ();
 sg13g2_decap_8 FILLER_48_1105 ();
 sg13g2_decap_8 FILLER_48_1112 ();
 sg13g2_decap_8 FILLER_48_1119 ();
 sg13g2_decap_8 FILLER_48_1126 ();
 sg13g2_decap_8 FILLER_48_1133 ();
 sg13g2_decap_8 FILLER_48_1140 ();
 sg13g2_decap_8 FILLER_48_1147 ();
 sg13g2_decap_8 FILLER_48_1154 ();
 sg13g2_decap_8 FILLER_48_1161 ();
 sg13g2_decap_8 FILLER_48_1168 ();
 sg13g2_decap_8 FILLER_48_1175 ();
 sg13g2_decap_8 FILLER_48_1182 ();
 sg13g2_decap_8 FILLER_48_1189 ();
 sg13g2_decap_8 FILLER_48_1196 ();
 sg13g2_decap_8 FILLER_48_1203 ();
 sg13g2_decap_8 FILLER_48_1210 ();
 sg13g2_decap_8 FILLER_48_1217 ();
 sg13g2_decap_8 FILLER_48_1224 ();
 sg13g2_decap_8 FILLER_48_1231 ();
 sg13g2_decap_8 FILLER_48_1238 ();
 sg13g2_decap_8 FILLER_48_1245 ();
 sg13g2_decap_8 FILLER_48_1252 ();
 sg13g2_decap_8 FILLER_48_1259 ();
 sg13g2_decap_8 FILLER_48_1266 ();
 sg13g2_decap_8 FILLER_48_1273 ();
 sg13g2_decap_8 FILLER_48_1280 ();
 sg13g2_decap_8 FILLER_48_1287 ();
 sg13g2_decap_8 FILLER_48_1294 ();
 sg13g2_decap_8 FILLER_48_1301 ();
 sg13g2_decap_8 FILLER_48_1308 ();
 sg13g2_decap_8 FILLER_48_1315 ();
 sg13g2_decap_8 FILLER_48_1322 ();
 sg13g2_decap_8 FILLER_48_1329 ();
 sg13g2_decap_8 FILLER_48_1336 ();
 sg13g2_decap_8 FILLER_48_1343 ();
 sg13g2_decap_8 FILLER_48_1350 ();
 sg13g2_decap_8 FILLER_48_1357 ();
 sg13g2_decap_8 FILLER_48_1364 ();
 sg13g2_decap_8 FILLER_48_1371 ();
 sg13g2_decap_8 FILLER_48_1378 ();
 sg13g2_decap_8 FILLER_48_1385 ();
 sg13g2_decap_8 FILLER_48_1392 ();
 sg13g2_decap_8 FILLER_48_1399 ();
 sg13g2_decap_8 FILLER_48_1406 ();
 sg13g2_decap_8 FILLER_48_1413 ();
 sg13g2_decap_8 FILLER_48_1420 ();
 sg13g2_decap_8 FILLER_48_1427 ();
 sg13g2_decap_8 FILLER_48_1434 ();
 sg13g2_decap_8 FILLER_48_1441 ();
 sg13g2_decap_8 FILLER_48_1448 ();
 sg13g2_decap_8 FILLER_48_1455 ();
 sg13g2_decap_8 FILLER_48_1462 ();
 sg13g2_decap_8 FILLER_48_1469 ();
 sg13g2_decap_8 FILLER_48_1476 ();
 sg13g2_decap_8 FILLER_48_1483 ();
 sg13g2_decap_8 FILLER_48_1490 ();
 sg13g2_decap_8 FILLER_48_1497 ();
 sg13g2_decap_8 FILLER_48_1504 ();
 sg13g2_decap_8 FILLER_48_1511 ();
 sg13g2_decap_8 FILLER_48_1518 ();
 sg13g2_decap_8 FILLER_48_1525 ();
 sg13g2_decap_8 FILLER_48_1532 ();
 sg13g2_decap_8 FILLER_48_1539 ();
 sg13g2_decap_8 FILLER_48_1546 ();
 sg13g2_decap_8 FILLER_48_1553 ();
 sg13g2_decap_8 FILLER_48_1560 ();
 sg13g2_decap_8 FILLER_48_1567 ();
 sg13g2_decap_8 FILLER_48_1574 ();
 sg13g2_decap_8 FILLER_48_1581 ();
 sg13g2_decap_8 FILLER_48_1588 ();
 sg13g2_decap_8 FILLER_48_1595 ();
 sg13g2_decap_8 FILLER_48_1602 ();
 sg13g2_decap_8 FILLER_48_1609 ();
 sg13g2_decap_8 FILLER_48_1616 ();
 sg13g2_decap_8 FILLER_48_1623 ();
 sg13g2_decap_8 FILLER_48_1630 ();
 sg13g2_decap_8 FILLER_48_1637 ();
 sg13g2_decap_8 FILLER_48_1644 ();
 sg13g2_decap_8 FILLER_48_1651 ();
 sg13g2_decap_8 FILLER_48_1658 ();
 sg13g2_decap_8 FILLER_48_1665 ();
 sg13g2_decap_8 FILLER_48_1672 ();
 sg13g2_decap_8 FILLER_48_1679 ();
 sg13g2_decap_8 FILLER_48_1686 ();
 sg13g2_decap_8 FILLER_48_1693 ();
 sg13g2_decap_8 FILLER_48_1700 ();
 sg13g2_decap_8 FILLER_48_1707 ();
 sg13g2_decap_8 FILLER_48_1714 ();
 sg13g2_decap_8 FILLER_48_1721 ();
 sg13g2_decap_8 FILLER_48_1728 ();
 sg13g2_decap_8 FILLER_48_1735 ();
 sg13g2_decap_8 FILLER_48_1742 ();
 sg13g2_decap_8 FILLER_48_1749 ();
 sg13g2_decap_8 FILLER_48_1756 ();
 sg13g2_decap_4 FILLER_48_1763 ();
 sg13g2_fill_1 FILLER_48_1767 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_7 ();
 sg13g2_decap_8 FILLER_49_14 ();
 sg13g2_decap_8 FILLER_49_21 ();
 sg13g2_decap_8 FILLER_49_28 ();
 sg13g2_decap_8 FILLER_49_35 ();
 sg13g2_decap_8 FILLER_49_42 ();
 sg13g2_decap_8 FILLER_49_49 ();
 sg13g2_decap_8 FILLER_49_56 ();
 sg13g2_decap_8 FILLER_49_63 ();
 sg13g2_decap_8 FILLER_49_70 ();
 sg13g2_fill_1 FILLER_49_116 ();
 sg13g2_fill_1 FILLER_49_145 ();
 sg13g2_fill_2 FILLER_49_151 ();
 sg13g2_fill_1 FILLER_49_192 ();
 sg13g2_fill_2 FILLER_49_243 ();
 sg13g2_fill_2 FILLER_49_251 ();
 sg13g2_fill_1 FILLER_49_268 ();
 sg13g2_decap_4 FILLER_49_300 ();
 sg13g2_fill_1 FILLER_49_304 ();
 sg13g2_fill_2 FILLER_49_330 ();
 sg13g2_decap_4 FILLER_49_358 ();
 sg13g2_fill_2 FILLER_49_380 ();
 sg13g2_decap_8 FILLER_49_418 ();
 sg13g2_fill_1 FILLER_49_425 ();
 sg13g2_fill_1 FILLER_49_454 ();
 sg13g2_fill_1 FILLER_49_479 ();
 sg13g2_fill_1 FILLER_49_502 ();
 sg13g2_fill_2 FILLER_49_517 ();
 sg13g2_fill_1 FILLER_49_519 ();
 sg13g2_fill_1 FILLER_49_533 ();
 sg13g2_fill_2 FILLER_49_551 ();
 sg13g2_decap_4 FILLER_49_558 ();
 sg13g2_fill_1 FILLER_49_562 ();
 sg13g2_decap_8 FILLER_49_571 ();
 sg13g2_decap_4 FILLER_49_587 ();
 sg13g2_fill_2 FILLER_49_620 ();
 sg13g2_fill_1 FILLER_49_652 ();
 sg13g2_decap_4 FILLER_49_658 ();
 sg13g2_fill_2 FILLER_49_662 ();
 sg13g2_fill_2 FILLER_49_669 ();
 sg13g2_decap_8 FILLER_49_679 ();
 sg13g2_fill_2 FILLER_49_686 ();
 sg13g2_decap_8 FILLER_49_705 ();
 sg13g2_decap_4 FILLER_49_712 ();
 sg13g2_fill_2 FILLER_49_716 ();
 sg13g2_fill_2 FILLER_49_732 ();
 sg13g2_fill_1 FILLER_49_734 ();
 sg13g2_decap_4 FILLER_49_758 ();
 sg13g2_decap_4 FILLER_49_791 ();
 sg13g2_fill_1 FILLER_49_795 ();
 sg13g2_fill_2 FILLER_49_805 ();
 sg13g2_fill_1 FILLER_49_807 ();
 sg13g2_fill_1 FILLER_49_825 ();
 sg13g2_decap_8 FILLER_49_831 ();
 sg13g2_decap_8 FILLER_49_838 ();
 sg13g2_decap_4 FILLER_49_845 ();
 sg13g2_fill_1 FILLER_49_849 ();
 sg13g2_decap_4 FILLER_49_866 ();
 sg13g2_fill_2 FILLER_49_870 ();
 sg13g2_fill_1 FILLER_49_898 ();
 sg13g2_fill_2 FILLER_49_925 ();
 sg13g2_fill_1 FILLER_49_927 ();
 sg13g2_decap_8 FILLER_49_951 ();
 sg13g2_fill_1 FILLER_49_958 ();
 sg13g2_decap_4 FILLER_49_970 ();
 sg13g2_fill_2 FILLER_49_974 ();
 sg13g2_decap_8 FILLER_49_1003 ();
 sg13g2_decap_8 FILLER_49_1010 ();
 sg13g2_decap_8 FILLER_49_1017 ();
 sg13g2_decap_8 FILLER_49_1024 ();
 sg13g2_decap_8 FILLER_49_1031 ();
 sg13g2_decap_8 FILLER_49_1038 ();
 sg13g2_decap_8 FILLER_49_1045 ();
 sg13g2_decap_8 FILLER_49_1052 ();
 sg13g2_decap_8 FILLER_49_1059 ();
 sg13g2_decap_8 FILLER_49_1066 ();
 sg13g2_decap_8 FILLER_49_1073 ();
 sg13g2_decap_8 FILLER_49_1080 ();
 sg13g2_decap_8 FILLER_49_1087 ();
 sg13g2_decap_8 FILLER_49_1094 ();
 sg13g2_decap_8 FILLER_49_1101 ();
 sg13g2_decap_8 FILLER_49_1108 ();
 sg13g2_decap_8 FILLER_49_1115 ();
 sg13g2_decap_8 FILLER_49_1122 ();
 sg13g2_decap_8 FILLER_49_1129 ();
 sg13g2_decap_8 FILLER_49_1136 ();
 sg13g2_decap_8 FILLER_49_1143 ();
 sg13g2_decap_8 FILLER_49_1150 ();
 sg13g2_decap_8 FILLER_49_1157 ();
 sg13g2_decap_8 FILLER_49_1164 ();
 sg13g2_decap_8 FILLER_49_1171 ();
 sg13g2_decap_8 FILLER_49_1178 ();
 sg13g2_decap_8 FILLER_49_1185 ();
 sg13g2_decap_8 FILLER_49_1192 ();
 sg13g2_decap_8 FILLER_49_1199 ();
 sg13g2_decap_8 FILLER_49_1206 ();
 sg13g2_decap_8 FILLER_49_1213 ();
 sg13g2_decap_8 FILLER_49_1220 ();
 sg13g2_decap_8 FILLER_49_1227 ();
 sg13g2_decap_8 FILLER_49_1234 ();
 sg13g2_decap_8 FILLER_49_1241 ();
 sg13g2_decap_8 FILLER_49_1248 ();
 sg13g2_decap_8 FILLER_49_1255 ();
 sg13g2_decap_8 FILLER_49_1262 ();
 sg13g2_decap_8 FILLER_49_1269 ();
 sg13g2_decap_8 FILLER_49_1276 ();
 sg13g2_decap_8 FILLER_49_1283 ();
 sg13g2_decap_8 FILLER_49_1290 ();
 sg13g2_decap_8 FILLER_49_1297 ();
 sg13g2_decap_8 FILLER_49_1304 ();
 sg13g2_decap_8 FILLER_49_1311 ();
 sg13g2_decap_8 FILLER_49_1318 ();
 sg13g2_decap_8 FILLER_49_1325 ();
 sg13g2_decap_8 FILLER_49_1332 ();
 sg13g2_decap_8 FILLER_49_1339 ();
 sg13g2_decap_8 FILLER_49_1346 ();
 sg13g2_decap_8 FILLER_49_1353 ();
 sg13g2_decap_8 FILLER_49_1360 ();
 sg13g2_decap_8 FILLER_49_1367 ();
 sg13g2_decap_8 FILLER_49_1374 ();
 sg13g2_decap_8 FILLER_49_1381 ();
 sg13g2_decap_8 FILLER_49_1388 ();
 sg13g2_decap_8 FILLER_49_1395 ();
 sg13g2_decap_8 FILLER_49_1402 ();
 sg13g2_decap_8 FILLER_49_1409 ();
 sg13g2_decap_8 FILLER_49_1416 ();
 sg13g2_decap_8 FILLER_49_1423 ();
 sg13g2_decap_8 FILLER_49_1430 ();
 sg13g2_decap_8 FILLER_49_1437 ();
 sg13g2_decap_8 FILLER_49_1444 ();
 sg13g2_decap_8 FILLER_49_1451 ();
 sg13g2_decap_8 FILLER_49_1458 ();
 sg13g2_decap_8 FILLER_49_1465 ();
 sg13g2_decap_8 FILLER_49_1472 ();
 sg13g2_decap_8 FILLER_49_1479 ();
 sg13g2_decap_8 FILLER_49_1486 ();
 sg13g2_decap_8 FILLER_49_1493 ();
 sg13g2_decap_8 FILLER_49_1500 ();
 sg13g2_decap_8 FILLER_49_1507 ();
 sg13g2_decap_8 FILLER_49_1514 ();
 sg13g2_decap_8 FILLER_49_1521 ();
 sg13g2_decap_8 FILLER_49_1528 ();
 sg13g2_decap_8 FILLER_49_1535 ();
 sg13g2_decap_8 FILLER_49_1542 ();
 sg13g2_decap_8 FILLER_49_1549 ();
 sg13g2_decap_8 FILLER_49_1556 ();
 sg13g2_decap_8 FILLER_49_1563 ();
 sg13g2_decap_8 FILLER_49_1570 ();
 sg13g2_decap_8 FILLER_49_1577 ();
 sg13g2_decap_8 FILLER_49_1584 ();
 sg13g2_decap_8 FILLER_49_1591 ();
 sg13g2_decap_8 FILLER_49_1598 ();
 sg13g2_decap_8 FILLER_49_1605 ();
 sg13g2_decap_8 FILLER_49_1612 ();
 sg13g2_decap_8 FILLER_49_1619 ();
 sg13g2_decap_8 FILLER_49_1626 ();
 sg13g2_decap_8 FILLER_49_1633 ();
 sg13g2_decap_8 FILLER_49_1640 ();
 sg13g2_decap_8 FILLER_49_1647 ();
 sg13g2_decap_8 FILLER_49_1654 ();
 sg13g2_decap_8 FILLER_49_1661 ();
 sg13g2_decap_8 FILLER_49_1668 ();
 sg13g2_decap_8 FILLER_49_1675 ();
 sg13g2_decap_8 FILLER_49_1682 ();
 sg13g2_decap_8 FILLER_49_1689 ();
 sg13g2_decap_8 FILLER_49_1696 ();
 sg13g2_decap_8 FILLER_49_1703 ();
 sg13g2_decap_8 FILLER_49_1710 ();
 sg13g2_decap_8 FILLER_49_1717 ();
 sg13g2_decap_8 FILLER_49_1724 ();
 sg13g2_decap_8 FILLER_49_1731 ();
 sg13g2_decap_8 FILLER_49_1738 ();
 sg13g2_decap_8 FILLER_49_1745 ();
 sg13g2_decap_8 FILLER_49_1752 ();
 sg13g2_decap_8 FILLER_49_1759 ();
 sg13g2_fill_2 FILLER_49_1766 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_8 FILLER_50_7 ();
 sg13g2_decap_8 FILLER_50_14 ();
 sg13g2_decap_8 FILLER_50_21 ();
 sg13g2_decap_8 FILLER_50_28 ();
 sg13g2_decap_8 FILLER_50_35 ();
 sg13g2_decap_8 FILLER_50_42 ();
 sg13g2_decap_8 FILLER_50_49 ();
 sg13g2_decap_8 FILLER_50_56 ();
 sg13g2_decap_8 FILLER_50_63 ();
 sg13g2_decap_4 FILLER_50_70 ();
 sg13g2_fill_2 FILLER_50_74 ();
 sg13g2_fill_2 FILLER_50_92 ();
 sg13g2_fill_1 FILLER_50_111 ();
 sg13g2_fill_1 FILLER_50_160 ();
 sg13g2_fill_1 FILLER_50_166 ();
 sg13g2_fill_2 FILLER_50_186 ();
 sg13g2_fill_2 FILLER_50_200 ();
 sg13g2_fill_1 FILLER_50_202 ();
 sg13g2_fill_1 FILLER_50_208 ();
 sg13g2_fill_2 FILLER_50_266 ();
 sg13g2_fill_1 FILLER_50_268 ();
 sg13g2_fill_2 FILLER_50_277 ();
 sg13g2_fill_1 FILLER_50_282 ();
 sg13g2_fill_1 FILLER_50_293 ();
 sg13g2_decap_8 FILLER_50_303 ();
 sg13g2_decap_4 FILLER_50_310 ();
 sg13g2_decap_4 FILLER_50_334 ();
 sg13g2_fill_1 FILLER_50_355 ();
 sg13g2_decap_8 FILLER_50_390 ();
 sg13g2_fill_2 FILLER_50_400 ();
 sg13g2_decap_4 FILLER_50_411 ();
 sg13g2_fill_2 FILLER_50_415 ();
 sg13g2_fill_2 FILLER_50_447 ();
 sg13g2_fill_1 FILLER_50_449 ();
 sg13g2_decap_8 FILLER_50_459 ();
 sg13g2_fill_1 FILLER_50_466 ();
 sg13g2_fill_2 FILLER_50_505 ();
 sg13g2_fill_1 FILLER_50_507 ();
 sg13g2_fill_2 FILLER_50_521 ();
 sg13g2_fill_1 FILLER_50_547 ();
 sg13g2_fill_1 FILLER_50_577 ();
 sg13g2_fill_2 FILLER_50_586 ();
 sg13g2_fill_1 FILLER_50_588 ();
 sg13g2_fill_1 FILLER_50_593 ();
 sg13g2_fill_1 FILLER_50_620 ();
 sg13g2_fill_2 FILLER_50_625 ();
 sg13g2_decap_4 FILLER_50_653 ();
 sg13g2_fill_1 FILLER_50_683 ();
 sg13g2_decap_4 FILLER_50_714 ();
 sg13g2_decap_4 FILLER_50_741 ();
 sg13g2_fill_1 FILLER_50_745 ();
 sg13g2_fill_2 FILLER_50_751 ();
 sg13g2_decap_4 FILLER_50_771 ();
 sg13g2_decap_8 FILLER_50_785 ();
 sg13g2_decap_4 FILLER_50_792 ();
 sg13g2_fill_2 FILLER_50_796 ();
 sg13g2_decap_4 FILLER_50_806 ();
 sg13g2_fill_2 FILLER_50_810 ();
 sg13g2_decap_4 FILLER_50_833 ();
 sg13g2_fill_2 FILLER_50_837 ();
 sg13g2_fill_1 FILLER_50_847 ();
 sg13g2_decap_8 FILLER_50_865 ();
 sg13g2_fill_2 FILLER_50_872 ();
 sg13g2_fill_1 FILLER_50_874 ();
 sg13g2_decap_4 FILLER_50_900 ();
 sg13g2_fill_1 FILLER_50_904 ();
 sg13g2_fill_1 FILLER_50_925 ();
 sg13g2_decap_4 FILLER_50_931 ();
 sg13g2_fill_2 FILLER_50_935 ();
 sg13g2_decap_4 FILLER_50_946 ();
 sg13g2_fill_1 FILLER_50_950 ();
 sg13g2_decap_4 FILLER_50_977 ();
 sg13g2_fill_2 FILLER_50_985 ();
 sg13g2_decap_8 FILLER_50_1000 ();
 sg13g2_decap_8 FILLER_50_1007 ();
 sg13g2_decap_8 FILLER_50_1014 ();
 sg13g2_decap_8 FILLER_50_1021 ();
 sg13g2_decap_8 FILLER_50_1028 ();
 sg13g2_decap_8 FILLER_50_1035 ();
 sg13g2_decap_8 FILLER_50_1042 ();
 sg13g2_decap_8 FILLER_50_1049 ();
 sg13g2_decap_8 FILLER_50_1056 ();
 sg13g2_decap_8 FILLER_50_1063 ();
 sg13g2_decap_8 FILLER_50_1070 ();
 sg13g2_decap_8 FILLER_50_1077 ();
 sg13g2_decap_8 FILLER_50_1084 ();
 sg13g2_decap_8 FILLER_50_1091 ();
 sg13g2_decap_8 FILLER_50_1098 ();
 sg13g2_decap_8 FILLER_50_1105 ();
 sg13g2_decap_8 FILLER_50_1112 ();
 sg13g2_decap_8 FILLER_50_1119 ();
 sg13g2_decap_8 FILLER_50_1126 ();
 sg13g2_decap_8 FILLER_50_1133 ();
 sg13g2_decap_8 FILLER_50_1140 ();
 sg13g2_decap_8 FILLER_50_1147 ();
 sg13g2_decap_8 FILLER_50_1154 ();
 sg13g2_decap_8 FILLER_50_1161 ();
 sg13g2_decap_8 FILLER_50_1168 ();
 sg13g2_decap_8 FILLER_50_1175 ();
 sg13g2_decap_8 FILLER_50_1182 ();
 sg13g2_decap_8 FILLER_50_1189 ();
 sg13g2_decap_8 FILLER_50_1196 ();
 sg13g2_decap_8 FILLER_50_1203 ();
 sg13g2_decap_8 FILLER_50_1210 ();
 sg13g2_decap_8 FILLER_50_1217 ();
 sg13g2_decap_8 FILLER_50_1224 ();
 sg13g2_decap_8 FILLER_50_1231 ();
 sg13g2_decap_8 FILLER_50_1238 ();
 sg13g2_decap_8 FILLER_50_1245 ();
 sg13g2_decap_8 FILLER_50_1252 ();
 sg13g2_decap_8 FILLER_50_1259 ();
 sg13g2_decap_8 FILLER_50_1266 ();
 sg13g2_decap_8 FILLER_50_1273 ();
 sg13g2_decap_8 FILLER_50_1280 ();
 sg13g2_decap_8 FILLER_50_1287 ();
 sg13g2_decap_8 FILLER_50_1294 ();
 sg13g2_decap_8 FILLER_50_1301 ();
 sg13g2_decap_8 FILLER_50_1308 ();
 sg13g2_decap_8 FILLER_50_1315 ();
 sg13g2_decap_8 FILLER_50_1322 ();
 sg13g2_decap_8 FILLER_50_1329 ();
 sg13g2_decap_8 FILLER_50_1336 ();
 sg13g2_decap_8 FILLER_50_1343 ();
 sg13g2_decap_8 FILLER_50_1350 ();
 sg13g2_decap_8 FILLER_50_1357 ();
 sg13g2_decap_8 FILLER_50_1364 ();
 sg13g2_decap_8 FILLER_50_1371 ();
 sg13g2_decap_8 FILLER_50_1378 ();
 sg13g2_decap_8 FILLER_50_1385 ();
 sg13g2_decap_8 FILLER_50_1392 ();
 sg13g2_decap_8 FILLER_50_1399 ();
 sg13g2_decap_8 FILLER_50_1406 ();
 sg13g2_decap_8 FILLER_50_1413 ();
 sg13g2_decap_8 FILLER_50_1420 ();
 sg13g2_decap_8 FILLER_50_1427 ();
 sg13g2_decap_8 FILLER_50_1434 ();
 sg13g2_decap_8 FILLER_50_1441 ();
 sg13g2_decap_8 FILLER_50_1448 ();
 sg13g2_decap_8 FILLER_50_1455 ();
 sg13g2_decap_8 FILLER_50_1462 ();
 sg13g2_decap_8 FILLER_50_1469 ();
 sg13g2_decap_8 FILLER_50_1476 ();
 sg13g2_decap_8 FILLER_50_1483 ();
 sg13g2_decap_8 FILLER_50_1490 ();
 sg13g2_decap_8 FILLER_50_1497 ();
 sg13g2_decap_8 FILLER_50_1504 ();
 sg13g2_decap_8 FILLER_50_1511 ();
 sg13g2_decap_8 FILLER_50_1518 ();
 sg13g2_decap_8 FILLER_50_1525 ();
 sg13g2_decap_8 FILLER_50_1532 ();
 sg13g2_decap_8 FILLER_50_1539 ();
 sg13g2_decap_8 FILLER_50_1546 ();
 sg13g2_decap_8 FILLER_50_1553 ();
 sg13g2_decap_8 FILLER_50_1560 ();
 sg13g2_decap_8 FILLER_50_1567 ();
 sg13g2_decap_8 FILLER_50_1574 ();
 sg13g2_decap_8 FILLER_50_1581 ();
 sg13g2_decap_8 FILLER_50_1588 ();
 sg13g2_decap_8 FILLER_50_1595 ();
 sg13g2_decap_8 FILLER_50_1602 ();
 sg13g2_decap_8 FILLER_50_1609 ();
 sg13g2_decap_8 FILLER_50_1616 ();
 sg13g2_decap_8 FILLER_50_1623 ();
 sg13g2_decap_8 FILLER_50_1630 ();
 sg13g2_decap_8 FILLER_50_1637 ();
 sg13g2_decap_8 FILLER_50_1644 ();
 sg13g2_decap_8 FILLER_50_1651 ();
 sg13g2_decap_8 FILLER_50_1658 ();
 sg13g2_decap_8 FILLER_50_1665 ();
 sg13g2_decap_8 FILLER_50_1672 ();
 sg13g2_decap_8 FILLER_50_1679 ();
 sg13g2_decap_8 FILLER_50_1686 ();
 sg13g2_decap_8 FILLER_50_1693 ();
 sg13g2_decap_8 FILLER_50_1700 ();
 sg13g2_decap_8 FILLER_50_1707 ();
 sg13g2_decap_8 FILLER_50_1714 ();
 sg13g2_decap_8 FILLER_50_1721 ();
 sg13g2_decap_8 FILLER_50_1728 ();
 sg13g2_decap_8 FILLER_50_1735 ();
 sg13g2_decap_8 FILLER_50_1742 ();
 sg13g2_decap_8 FILLER_50_1749 ();
 sg13g2_decap_8 FILLER_50_1756 ();
 sg13g2_decap_4 FILLER_50_1763 ();
 sg13g2_fill_1 FILLER_50_1767 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_decap_8 FILLER_51_7 ();
 sg13g2_decap_8 FILLER_51_14 ();
 sg13g2_decap_8 FILLER_51_21 ();
 sg13g2_decap_8 FILLER_51_28 ();
 sg13g2_decap_8 FILLER_51_35 ();
 sg13g2_decap_8 FILLER_51_42 ();
 sg13g2_decap_8 FILLER_51_49 ();
 sg13g2_decap_8 FILLER_51_56 ();
 sg13g2_decap_4 FILLER_51_63 ();
 sg13g2_fill_2 FILLER_51_67 ();
 sg13g2_fill_2 FILLER_51_98 ();
 sg13g2_fill_1 FILLER_51_135 ();
 sg13g2_fill_2 FILLER_51_161 ();
 sg13g2_decap_4 FILLER_51_191 ();
 sg13g2_fill_1 FILLER_51_251 ();
 sg13g2_fill_2 FILLER_51_271 ();
 sg13g2_fill_1 FILLER_51_301 ();
 sg13g2_fill_2 FILLER_51_352 ();
 sg13g2_fill_1 FILLER_51_423 ();
 sg13g2_fill_2 FILLER_51_456 ();
 sg13g2_fill_2 FILLER_51_472 ();
 sg13g2_fill_1 FILLER_51_474 ();
 sg13g2_fill_2 FILLER_51_489 ();
 sg13g2_fill_1 FILLER_51_491 ();
 sg13g2_fill_2 FILLER_51_514 ();
 sg13g2_fill_1 FILLER_51_516 ();
 sg13g2_decap_4 FILLER_51_529 ();
 sg13g2_decap_8 FILLER_51_547 ();
 sg13g2_decap_4 FILLER_51_554 ();
 sg13g2_fill_1 FILLER_51_579 ();
 sg13g2_fill_2 FILLER_51_596 ();
 sg13g2_fill_1 FILLER_51_608 ();
 sg13g2_fill_2 FILLER_51_614 ();
 sg13g2_fill_2 FILLER_51_656 ();
 sg13g2_decap_4 FILLER_51_689 ();
 sg13g2_decap_4 FILLER_51_698 ();
 sg13g2_fill_2 FILLER_51_702 ();
 sg13g2_decap_8 FILLER_51_708 ();
 sg13g2_decap_4 FILLER_51_715 ();
 sg13g2_fill_2 FILLER_51_749 ();
 sg13g2_fill_1 FILLER_51_751 ();
 sg13g2_fill_1 FILLER_51_766 ();
 sg13g2_fill_1 FILLER_51_772 ();
 sg13g2_decap_4 FILLER_51_782 ();
 sg13g2_fill_1 FILLER_51_786 ();
 sg13g2_decap_4 FILLER_51_813 ();
 sg13g2_decap_8 FILLER_51_822 ();
 sg13g2_fill_2 FILLER_51_829 ();
 sg13g2_fill_2 FILLER_51_841 ();
 sg13g2_fill_1 FILLER_51_859 ();
 sg13g2_decap_8 FILLER_51_870 ();
 sg13g2_fill_2 FILLER_51_877 ();
 sg13g2_fill_1 FILLER_51_879 ();
 sg13g2_decap_8 FILLER_51_892 ();
 sg13g2_decap_4 FILLER_51_899 ();
 sg13g2_fill_1 FILLER_51_903 ();
 sg13g2_decap_4 FILLER_51_917 ();
 sg13g2_fill_1 FILLER_51_921 ();
 sg13g2_decap_4 FILLER_51_954 ();
 sg13g2_decap_8 FILLER_51_991 ();
 sg13g2_decap_8 FILLER_51_998 ();
 sg13g2_decap_8 FILLER_51_1005 ();
 sg13g2_decap_8 FILLER_51_1012 ();
 sg13g2_decap_8 FILLER_51_1019 ();
 sg13g2_decap_8 FILLER_51_1026 ();
 sg13g2_decap_8 FILLER_51_1033 ();
 sg13g2_decap_8 FILLER_51_1040 ();
 sg13g2_decap_8 FILLER_51_1047 ();
 sg13g2_decap_8 FILLER_51_1054 ();
 sg13g2_decap_8 FILLER_51_1061 ();
 sg13g2_decap_8 FILLER_51_1068 ();
 sg13g2_decap_8 FILLER_51_1075 ();
 sg13g2_decap_8 FILLER_51_1082 ();
 sg13g2_decap_8 FILLER_51_1089 ();
 sg13g2_decap_8 FILLER_51_1096 ();
 sg13g2_decap_8 FILLER_51_1103 ();
 sg13g2_decap_8 FILLER_51_1110 ();
 sg13g2_decap_8 FILLER_51_1117 ();
 sg13g2_decap_8 FILLER_51_1124 ();
 sg13g2_decap_8 FILLER_51_1131 ();
 sg13g2_decap_8 FILLER_51_1138 ();
 sg13g2_decap_8 FILLER_51_1145 ();
 sg13g2_decap_8 FILLER_51_1152 ();
 sg13g2_decap_8 FILLER_51_1159 ();
 sg13g2_decap_8 FILLER_51_1166 ();
 sg13g2_decap_8 FILLER_51_1173 ();
 sg13g2_decap_8 FILLER_51_1180 ();
 sg13g2_decap_8 FILLER_51_1187 ();
 sg13g2_decap_8 FILLER_51_1194 ();
 sg13g2_decap_8 FILLER_51_1201 ();
 sg13g2_decap_8 FILLER_51_1208 ();
 sg13g2_decap_8 FILLER_51_1215 ();
 sg13g2_decap_8 FILLER_51_1222 ();
 sg13g2_decap_8 FILLER_51_1229 ();
 sg13g2_decap_8 FILLER_51_1236 ();
 sg13g2_decap_8 FILLER_51_1243 ();
 sg13g2_decap_8 FILLER_51_1250 ();
 sg13g2_decap_8 FILLER_51_1257 ();
 sg13g2_decap_8 FILLER_51_1264 ();
 sg13g2_decap_8 FILLER_51_1271 ();
 sg13g2_decap_8 FILLER_51_1278 ();
 sg13g2_decap_8 FILLER_51_1285 ();
 sg13g2_decap_8 FILLER_51_1292 ();
 sg13g2_decap_8 FILLER_51_1299 ();
 sg13g2_decap_8 FILLER_51_1306 ();
 sg13g2_decap_8 FILLER_51_1313 ();
 sg13g2_decap_8 FILLER_51_1320 ();
 sg13g2_decap_8 FILLER_51_1327 ();
 sg13g2_decap_8 FILLER_51_1334 ();
 sg13g2_decap_8 FILLER_51_1341 ();
 sg13g2_decap_8 FILLER_51_1348 ();
 sg13g2_decap_8 FILLER_51_1355 ();
 sg13g2_decap_8 FILLER_51_1362 ();
 sg13g2_decap_8 FILLER_51_1369 ();
 sg13g2_decap_8 FILLER_51_1376 ();
 sg13g2_decap_8 FILLER_51_1383 ();
 sg13g2_decap_8 FILLER_51_1390 ();
 sg13g2_decap_8 FILLER_51_1397 ();
 sg13g2_decap_8 FILLER_51_1404 ();
 sg13g2_decap_8 FILLER_51_1411 ();
 sg13g2_decap_8 FILLER_51_1418 ();
 sg13g2_decap_8 FILLER_51_1425 ();
 sg13g2_decap_8 FILLER_51_1432 ();
 sg13g2_decap_8 FILLER_51_1439 ();
 sg13g2_decap_8 FILLER_51_1446 ();
 sg13g2_decap_8 FILLER_51_1453 ();
 sg13g2_decap_8 FILLER_51_1460 ();
 sg13g2_decap_8 FILLER_51_1467 ();
 sg13g2_decap_8 FILLER_51_1474 ();
 sg13g2_decap_8 FILLER_51_1481 ();
 sg13g2_decap_8 FILLER_51_1488 ();
 sg13g2_decap_8 FILLER_51_1495 ();
 sg13g2_decap_8 FILLER_51_1502 ();
 sg13g2_decap_8 FILLER_51_1509 ();
 sg13g2_decap_8 FILLER_51_1516 ();
 sg13g2_decap_8 FILLER_51_1523 ();
 sg13g2_decap_8 FILLER_51_1530 ();
 sg13g2_decap_8 FILLER_51_1537 ();
 sg13g2_decap_8 FILLER_51_1544 ();
 sg13g2_decap_8 FILLER_51_1551 ();
 sg13g2_decap_8 FILLER_51_1558 ();
 sg13g2_decap_8 FILLER_51_1565 ();
 sg13g2_decap_8 FILLER_51_1572 ();
 sg13g2_decap_8 FILLER_51_1579 ();
 sg13g2_decap_8 FILLER_51_1586 ();
 sg13g2_decap_8 FILLER_51_1593 ();
 sg13g2_decap_8 FILLER_51_1600 ();
 sg13g2_decap_8 FILLER_51_1607 ();
 sg13g2_decap_8 FILLER_51_1614 ();
 sg13g2_decap_8 FILLER_51_1621 ();
 sg13g2_decap_8 FILLER_51_1628 ();
 sg13g2_decap_8 FILLER_51_1635 ();
 sg13g2_decap_8 FILLER_51_1642 ();
 sg13g2_decap_8 FILLER_51_1649 ();
 sg13g2_decap_8 FILLER_51_1656 ();
 sg13g2_decap_8 FILLER_51_1663 ();
 sg13g2_decap_8 FILLER_51_1670 ();
 sg13g2_decap_8 FILLER_51_1677 ();
 sg13g2_decap_8 FILLER_51_1684 ();
 sg13g2_decap_8 FILLER_51_1691 ();
 sg13g2_decap_8 FILLER_51_1698 ();
 sg13g2_decap_8 FILLER_51_1705 ();
 sg13g2_decap_8 FILLER_51_1712 ();
 sg13g2_decap_8 FILLER_51_1719 ();
 sg13g2_decap_8 FILLER_51_1726 ();
 sg13g2_decap_8 FILLER_51_1733 ();
 sg13g2_decap_8 FILLER_51_1740 ();
 sg13g2_decap_8 FILLER_51_1747 ();
 sg13g2_decap_8 FILLER_51_1754 ();
 sg13g2_decap_8 FILLER_51_1761 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_decap_8 FILLER_52_7 ();
 sg13g2_decap_8 FILLER_52_14 ();
 sg13g2_decap_8 FILLER_52_21 ();
 sg13g2_decap_8 FILLER_52_28 ();
 sg13g2_decap_8 FILLER_52_35 ();
 sg13g2_decap_8 FILLER_52_42 ();
 sg13g2_decap_8 FILLER_52_49 ();
 sg13g2_decap_8 FILLER_52_56 ();
 sg13g2_fill_1 FILLER_52_63 ();
 sg13g2_fill_1 FILLER_52_117 ();
 sg13g2_fill_2 FILLER_52_199 ();
 sg13g2_fill_1 FILLER_52_224 ();
 sg13g2_fill_2 FILLER_52_240 ();
 sg13g2_fill_1 FILLER_52_245 ();
 sg13g2_fill_1 FILLER_52_254 ();
 sg13g2_fill_2 FILLER_52_286 ();
 sg13g2_fill_1 FILLER_52_327 ();
 sg13g2_decap_8 FILLER_52_337 ();
 sg13g2_decap_4 FILLER_52_344 ();
 sg13g2_fill_1 FILLER_52_394 ();
 sg13g2_fill_2 FILLER_52_493 ();
 sg13g2_fill_1 FILLER_52_495 ();
 sg13g2_fill_2 FILLER_52_514 ();
 sg13g2_fill_2 FILLER_52_552 ();
 sg13g2_decap_8 FILLER_52_577 ();
 sg13g2_fill_2 FILLER_52_584 ();
 sg13g2_fill_1 FILLER_52_601 ();
 sg13g2_fill_2 FILLER_52_606 ();
 sg13g2_fill_1 FILLER_52_608 ();
 sg13g2_decap_4 FILLER_52_614 ();
 sg13g2_fill_1 FILLER_52_618 ();
 sg13g2_fill_2 FILLER_52_624 ();
 sg13g2_fill_1 FILLER_52_640 ();
 sg13g2_fill_2 FILLER_52_650 ();
 sg13g2_fill_2 FILLER_52_684 ();
 sg13g2_fill_1 FILLER_52_686 ();
 sg13g2_decap_4 FILLER_52_709 ();
 sg13g2_decap_4 FILLER_52_734 ();
 sg13g2_fill_2 FILLER_52_810 ();
 sg13g2_fill_1 FILLER_52_819 ();
 sg13g2_fill_1 FILLER_52_840 ();
 sg13g2_fill_1 FILLER_52_871 ();
 sg13g2_fill_1 FILLER_52_876 ();
 sg13g2_fill_2 FILLER_52_881 ();
 sg13g2_fill_1 FILLER_52_883 ();
 sg13g2_fill_2 FILLER_52_894 ();
 sg13g2_fill_2 FILLER_52_903 ();
 sg13g2_fill_1 FILLER_52_905 ();
 sg13g2_fill_2 FILLER_52_924 ();
 sg13g2_fill_1 FILLER_52_926 ();
 sg13g2_fill_2 FILLER_52_931 ();
 sg13g2_decap_4 FILLER_52_946 ();
 sg13g2_fill_1 FILLER_52_950 ();
 sg13g2_decap_8 FILLER_52_961 ();
 sg13g2_fill_2 FILLER_52_968 ();
 sg13g2_fill_1 FILLER_52_970 ();
 sg13g2_decap_8 FILLER_52_975 ();
 sg13g2_decap_8 FILLER_52_982 ();
 sg13g2_decap_8 FILLER_52_989 ();
 sg13g2_decap_8 FILLER_52_996 ();
 sg13g2_decap_8 FILLER_52_1003 ();
 sg13g2_decap_8 FILLER_52_1010 ();
 sg13g2_decap_8 FILLER_52_1017 ();
 sg13g2_decap_8 FILLER_52_1024 ();
 sg13g2_decap_8 FILLER_52_1031 ();
 sg13g2_decap_8 FILLER_52_1038 ();
 sg13g2_decap_8 FILLER_52_1045 ();
 sg13g2_decap_8 FILLER_52_1052 ();
 sg13g2_decap_8 FILLER_52_1059 ();
 sg13g2_decap_8 FILLER_52_1066 ();
 sg13g2_decap_8 FILLER_52_1073 ();
 sg13g2_decap_8 FILLER_52_1080 ();
 sg13g2_decap_8 FILLER_52_1087 ();
 sg13g2_decap_8 FILLER_52_1094 ();
 sg13g2_decap_8 FILLER_52_1101 ();
 sg13g2_decap_8 FILLER_52_1108 ();
 sg13g2_decap_8 FILLER_52_1115 ();
 sg13g2_decap_8 FILLER_52_1122 ();
 sg13g2_decap_8 FILLER_52_1129 ();
 sg13g2_decap_8 FILLER_52_1136 ();
 sg13g2_decap_8 FILLER_52_1143 ();
 sg13g2_decap_8 FILLER_52_1150 ();
 sg13g2_decap_8 FILLER_52_1157 ();
 sg13g2_decap_8 FILLER_52_1164 ();
 sg13g2_decap_8 FILLER_52_1171 ();
 sg13g2_decap_8 FILLER_52_1178 ();
 sg13g2_decap_8 FILLER_52_1185 ();
 sg13g2_decap_8 FILLER_52_1192 ();
 sg13g2_decap_8 FILLER_52_1199 ();
 sg13g2_decap_8 FILLER_52_1206 ();
 sg13g2_decap_8 FILLER_52_1213 ();
 sg13g2_decap_8 FILLER_52_1220 ();
 sg13g2_decap_8 FILLER_52_1227 ();
 sg13g2_decap_8 FILLER_52_1234 ();
 sg13g2_decap_8 FILLER_52_1241 ();
 sg13g2_decap_8 FILLER_52_1248 ();
 sg13g2_decap_8 FILLER_52_1255 ();
 sg13g2_decap_8 FILLER_52_1262 ();
 sg13g2_decap_8 FILLER_52_1269 ();
 sg13g2_decap_8 FILLER_52_1276 ();
 sg13g2_decap_8 FILLER_52_1283 ();
 sg13g2_decap_8 FILLER_52_1290 ();
 sg13g2_decap_8 FILLER_52_1297 ();
 sg13g2_decap_8 FILLER_52_1304 ();
 sg13g2_decap_8 FILLER_52_1311 ();
 sg13g2_decap_8 FILLER_52_1318 ();
 sg13g2_decap_8 FILLER_52_1325 ();
 sg13g2_decap_8 FILLER_52_1332 ();
 sg13g2_decap_8 FILLER_52_1339 ();
 sg13g2_decap_8 FILLER_52_1346 ();
 sg13g2_decap_8 FILLER_52_1353 ();
 sg13g2_decap_8 FILLER_52_1360 ();
 sg13g2_decap_8 FILLER_52_1367 ();
 sg13g2_decap_8 FILLER_52_1374 ();
 sg13g2_decap_8 FILLER_52_1381 ();
 sg13g2_decap_8 FILLER_52_1388 ();
 sg13g2_decap_8 FILLER_52_1395 ();
 sg13g2_decap_8 FILLER_52_1402 ();
 sg13g2_decap_8 FILLER_52_1409 ();
 sg13g2_decap_8 FILLER_52_1416 ();
 sg13g2_decap_8 FILLER_52_1423 ();
 sg13g2_decap_8 FILLER_52_1430 ();
 sg13g2_decap_8 FILLER_52_1437 ();
 sg13g2_decap_8 FILLER_52_1444 ();
 sg13g2_decap_8 FILLER_52_1451 ();
 sg13g2_decap_8 FILLER_52_1458 ();
 sg13g2_decap_8 FILLER_52_1465 ();
 sg13g2_decap_8 FILLER_52_1472 ();
 sg13g2_decap_8 FILLER_52_1479 ();
 sg13g2_decap_8 FILLER_52_1486 ();
 sg13g2_decap_8 FILLER_52_1493 ();
 sg13g2_decap_8 FILLER_52_1500 ();
 sg13g2_decap_8 FILLER_52_1507 ();
 sg13g2_decap_8 FILLER_52_1514 ();
 sg13g2_decap_8 FILLER_52_1521 ();
 sg13g2_decap_8 FILLER_52_1528 ();
 sg13g2_decap_8 FILLER_52_1535 ();
 sg13g2_decap_8 FILLER_52_1542 ();
 sg13g2_decap_8 FILLER_52_1549 ();
 sg13g2_decap_8 FILLER_52_1556 ();
 sg13g2_decap_8 FILLER_52_1563 ();
 sg13g2_decap_8 FILLER_52_1570 ();
 sg13g2_decap_8 FILLER_52_1577 ();
 sg13g2_decap_8 FILLER_52_1584 ();
 sg13g2_decap_8 FILLER_52_1591 ();
 sg13g2_decap_8 FILLER_52_1598 ();
 sg13g2_decap_8 FILLER_52_1605 ();
 sg13g2_decap_8 FILLER_52_1612 ();
 sg13g2_decap_8 FILLER_52_1619 ();
 sg13g2_decap_8 FILLER_52_1626 ();
 sg13g2_decap_8 FILLER_52_1633 ();
 sg13g2_decap_8 FILLER_52_1640 ();
 sg13g2_decap_8 FILLER_52_1647 ();
 sg13g2_decap_8 FILLER_52_1654 ();
 sg13g2_decap_8 FILLER_52_1661 ();
 sg13g2_decap_8 FILLER_52_1668 ();
 sg13g2_decap_8 FILLER_52_1675 ();
 sg13g2_decap_8 FILLER_52_1682 ();
 sg13g2_decap_8 FILLER_52_1689 ();
 sg13g2_decap_8 FILLER_52_1696 ();
 sg13g2_decap_8 FILLER_52_1703 ();
 sg13g2_decap_8 FILLER_52_1710 ();
 sg13g2_decap_8 FILLER_52_1717 ();
 sg13g2_decap_8 FILLER_52_1724 ();
 sg13g2_decap_8 FILLER_52_1731 ();
 sg13g2_decap_8 FILLER_52_1738 ();
 sg13g2_decap_8 FILLER_52_1745 ();
 sg13g2_decap_8 FILLER_52_1752 ();
 sg13g2_decap_8 FILLER_52_1759 ();
 sg13g2_fill_2 FILLER_52_1766 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_decap_8 FILLER_53_7 ();
 sg13g2_decap_8 FILLER_53_14 ();
 sg13g2_decap_8 FILLER_53_21 ();
 sg13g2_decap_8 FILLER_53_28 ();
 sg13g2_decap_8 FILLER_53_35 ();
 sg13g2_decap_8 FILLER_53_42 ();
 sg13g2_decap_8 FILLER_53_49 ();
 sg13g2_decap_8 FILLER_53_56 ();
 sg13g2_decap_8 FILLER_53_63 ();
 sg13g2_decap_4 FILLER_53_70 ();
 sg13g2_fill_2 FILLER_53_74 ();
 sg13g2_fill_1 FILLER_53_117 ();
 sg13g2_fill_1 FILLER_53_154 ();
 sg13g2_fill_2 FILLER_53_163 ();
 sg13g2_fill_2 FILLER_53_220 ();
 sg13g2_fill_1 FILLER_53_256 ();
 sg13g2_fill_1 FILLER_53_270 ();
 sg13g2_fill_2 FILLER_53_276 ();
 sg13g2_fill_1 FILLER_53_313 ();
 sg13g2_fill_1 FILLER_53_386 ();
 sg13g2_fill_1 FILLER_53_406 ();
 sg13g2_fill_1 FILLER_53_473 ();
 sg13g2_fill_2 FILLER_53_539 ();
 sg13g2_fill_1 FILLER_53_541 ();
 sg13g2_fill_1 FILLER_53_574 ();
 sg13g2_decap_8 FILLER_53_583 ();
 sg13g2_fill_1 FILLER_53_590 ();
 sg13g2_decap_4 FILLER_53_601 ();
 sg13g2_decap_4 FILLER_53_620 ();
 sg13g2_decap_8 FILLER_53_627 ();
 sg13g2_fill_2 FILLER_53_634 ();
 sg13g2_fill_1 FILLER_53_636 ();
 sg13g2_fill_2 FILLER_53_644 ();
 sg13g2_decap_4 FILLER_53_679 ();
 sg13g2_fill_1 FILLER_53_683 ();
 sg13g2_fill_1 FILLER_53_688 ();
 sg13g2_decap_4 FILLER_53_715 ();
 sg13g2_fill_2 FILLER_53_719 ();
 sg13g2_decap_8 FILLER_53_726 ();
 sg13g2_decap_4 FILLER_53_733 ();
 sg13g2_fill_1 FILLER_53_752 ();
 sg13g2_fill_2 FILLER_53_762 ();
 sg13g2_fill_1 FILLER_53_764 ();
 sg13g2_fill_1 FILLER_53_774 ();
 sg13g2_fill_2 FILLER_53_780 ();
 sg13g2_fill_2 FILLER_53_791 ();
 sg13g2_fill_1 FILLER_53_793 ();
 sg13g2_fill_1 FILLER_53_811 ();
 sg13g2_fill_2 FILLER_53_833 ();
 sg13g2_fill_2 FILLER_53_855 ();
 sg13g2_decap_8 FILLER_53_866 ();
 sg13g2_decap_8 FILLER_53_873 ();
 sg13g2_fill_2 FILLER_53_890 ();
 sg13g2_fill_1 FILLER_53_892 ();
 sg13g2_fill_2 FILLER_53_898 ();
 sg13g2_decap_8 FILLER_53_915 ();
 sg13g2_decap_8 FILLER_53_922 ();
 sg13g2_decap_8 FILLER_53_929 ();
 sg13g2_decap_4 FILLER_53_936 ();
 sg13g2_fill_2 FILLER_53_971 ();
 sg13g2_decap_8 FILLER_53_996 ();
 sg13g2_decap_8 FILLER_53_1003 ();
 sg13g2_decap_8 FILLER_53_1010 ();
 sg13g2_decap_8 FILLER_53_1017 ();
 sg13g2_decap_8 FILLER_53_1024 ();
 sg13g2_decap_8 FILLER_53_1031 ();
 sg13g2_decap_8 FILLER_53_1038 ();
 sg13g2_decap_8 FILLER_53_1045 ();
 sg13g2_decap_8 FILLER_53_1052 ();
 sg13g2_decap_8 FILLER_53_1059 ();
 sg13g2_decap_8 FILLER_53_1066 ();
 sg13g2_decap_8 FILLER_53_1073 ();
 sg13g2_decap_8 FILLER_53_1080 ();
 sg13g2_decap_8 FILLER_53_1087 ();
 sg13g2_decap_8 FILLER_53_1094 ();
 sg13g2_decap_8 FILLER_53_1101 ();
 sg13g2_decap_8 FILLER_53_1108 ();
 sg13g2_decap_8 FILLER_53_1115 ();
 sg13g2_decap_8 FILLER_53_1122 ();
 sg13g2_decap_8 FILLER_53_1129 ();
 sg13g2_decap_8 FILLER_53_1136 ();
 sg13g2_decap_8 FILLER_53_1143 ();
 sg13g2_decap_8 FILLER_53_1150 ();
 sg13g2_decap_8 FILLER_53_1157 ();
 sg13g2_decap_8 FILLER_53_1164 ();
 sg13g2_decap_8 FILLER_53_1171 ();
 sg13g2_decap_8 FILLER_53_1178 ();
 sg13g2_decap_8 FILLER_53_1185 ();
 sg13g2_decap_8 FILLER_53_1192 ();
 sg13g2_decap_8 FILLER_53_1199 ();
 sg13g2_decap_8 FILLER_53_1206 ();
 sg13g2_decap_8 FILLER_53_1213 ();
 sg13g2_decap_8 FILLER_53_1220 ();
 sg13g2_decap_8 FILLER_53_1227 ();
 sg13g2_decap_8 FILLER_53_1234 ();
 sg13g2_decap_8 FILLER_53_1241 ();
 sg13g2_decap_8 FILLER_53_1248 ();
 sg13g2_decap_8 FILLER_53_1255 ();
 sg13g2_decap_8 FILLER_53_1262 ();
 sg13g2_decap_8 FILLER_53_1269 ();
 sg13g2_decap_8 FILLER_53_1276 ();
 sg13g2_decap_8 FILLER_53_1283 ();
 sg13g2_decap_8 FILLER_53_1290 ();
 sg13g2_decap_8 FILLER_53_1297 ();
 sg13g2_decap_8 FILLER_53_1304 ();
 sg13g2_decap_8 FILLER_53_1311 ();
 sg13g2_decap_8 FILLER_53_1318 ();
 sg13g2_decap_8 FILLER_53_1325 ();
 sg13g2_decap_8 FILLER_53_1332 ();
 sg13g2_decap_8 FILLER_53_1339 ();
 sg13g2_decap_8 FILLER_53_1346 ();
 sg13g2_decap_8 FILLER_53_1353 ();
 sg13g2_decap_8 FILLER_53_1360 ();
 sg13g2_decap_8 FILLER_53_1367 ();
 sg13g2_decap_8 FILLER_53_1374 ();
 sg13g2_decap_8 FILLER_53_1381 ();
 sg13g2_decap_8 FILLER_53_1388 ();
 sg13g2_decap_8 FILLER_53_1395 ();
 sg13g2_decap_8 FILLER_53_1402 ();
 sg13g2_decap_8 FILLER_53_1409 ();
 sg13g2_decap_8 FILLER_53_1416 ();
 sg13g2_decap_8 FILLER_53_1423 ();
 sg13g2_decap_8 FILLER_53_1430 ();
 sg13g2_decap_8 FILLER_53_1437 ();
 sg13g2_decap_8 FILLER_53_1444 ();
 sg13g2_decap_8 FILLER_53_1451 ();
 sg13g2_decap_8 FILLER_53_1458 ();
 sg13g2_decap_8 FILLER_53_1465 ();
 sg13g2_decap_8 FILLER_53_1472 ();
 sg13g2_decap_8 FILLER_53_1479 ();
 sg13g2_decap_8 FILLER_53_1486 ();
 sg13g2_decap_8 FILLER_53_1493 ();
 sg13g2_decap_8 FILLER_53_1500 ();
 sg13g2_decap_8 FILLER_53_1507 ();
 sg13g2_decap_8 FILLER_53_1514 ();
 sg13g2_decap_8 FILLER_53_1521 ();
 sg13g2_decap_8 FILLER_53_1528 ();
 sg13g2_decap_8 FILLER_53_1535 ();
 sg13g2_decap_8 FILLER_53_1542 ();
 sg13g2_decap_8 FILLER_53_1549 ();
 sg13g2_decap_8 FILLER_53_1556 ();
 sg13g2_decap_8 FILLER_53_1563 ();
 sg13g2_decap_8 FILLER_53_1570 ();
 sg13g2_decap_8 FILLER_53_1577 ();
 sg13g2_decap_8 FILLER_53_1584 ();
 sg13g2_decap_8 FILLER_53_1591 ();
 sg13g2_decap_8 FILLER_53_1598 ();
 sg13g2_decap_8 FILLER_53_1605 ();
 sg13g2_decap_8 FILLER_53_1612 ();
 sg13g2_decap_8 FILLER_53_1619 ();
 sg13g2_decap_8 FILLER_53_1626 ();
 sg13g2_decap_8 FILLER_53_1633 ();
 sg13g2_decap_8 FILLER_53_1640 ();
 sg13g2_decap_8 FILLER_53_1647 ();
 sg13g2_decap_8 FILLER_53_1654 ();
 sg13g2_decap_8 FILLER_53_1661 ();
 sg13g2_decap_8 FILLER_53_1668 ();
 sg13g2_decap_8 FILLER_53_1675 ();
 sg13g2_decap_8 FILLER_53_1682 ();
 sg13g2_decap_8 FILLER_53_1689 ();
 sg13g2_decap_8 FILLER_53_1696 ();
 sg13g2_decap_8 FILLER_53_1703 ();
 sg13g2_decap_8 FILLER_53_1710 ();
 sg13g2_decap_8 FILLER_53_1717 ();
 sg13g2_decap_8 FILLER_53_1724 ();
 sg13g2_decap_8 FILLER_53_1731 ();
 sg13g2_decap_8 FILLER_53_1738 ();
 sg13g2_decap_8 FILLER_53_1745 ();
 sg13g2_decap_8 FILLER_53_1752 ();
 sg13g2_decap_8 FILLER_53_1759 ();
 sg13g2_fill_2 FILLER_53_1766 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_decap_8 FILLER_54_7 ();
 sg13g2_decap_8 FILLER_54_14 ();
 sg13g2_decap_8 FILLER_54_21 ();
 sg13g2_decap_8 FILLER_54_28 ();
 sg13g2_decap_8 FILLER_54_35 ();
 sg13g2_decap_8 FILLER_54_42 ();
 sg13g2_decap_8 FILLER_54_49 ();
 sg13g2_decap_8 FILLER_54_56 ();
 sg13g2_decap_8 FILLER_54_63 ();
 sg13g2_decap_8 FILLER_54_70 ();
 sg13g2_fill_1 FILLER_54_77 ();
 sg13g2_fill_1 FILLER_54_112 ();
 sg13g2_fill_2 FILLER_54_140 ();
 sg13g2_fill_1 FILLER_54_155 ();
 sg13g2_fill_1 FILLER_54_192 ();
 sg13g2_fill_2 FILLER_54_207 ();
 sg13g2_fill_1 FILLER_54_223 ();
 sg13g2_fill_2 FILLER_54_242 ();
 sg13g2_decap_8 FILLER_54_320 ();
 sg13g2_fill_2 FILLER_54_501 ();
 sg13g2_decap_4 FILLER_54_542 ();
 sg13g2_fill_2 FILLER_54_546 ();
 sg13g2_decap_8 FILLER_54_551 ();
 sg13g2_decap_8 FILLER_54_578 ();
 sg13g2_decap_4 FILLER_54_585 ();
 sg13g2_fill_1 FILLER_54_589 ();
 sg13g2_fill_2 FILLER_54_603 ();
 sg13g2_fill_1 FILLER_54_605 ();
 sg13g2_fill_1 FILLER_54_613 ();
 sg13g2_fill_1 FILLER_54_621 ();
 sg13g2_fill_1 FILLER_54_648 ();
 sg13g2_decap_8 FILLER_54_662 ();
 sg13g2_fill_1 FILLER_54_688 ();
 sg13g2_fill_2 FILLER_54_717 ();
 sg13g2_fill_2 FILLER_54_753 ();
 sg13g2_fill_2 FILLER_54_763 ();
 sg13g2_fill_2 FILLER_54_789 ();
 sg13g2_fill_1 FILLER_54_791 ();
 sg13g2_decap_8 FILLER_54_910 ();
 sg13g2_fill_2 FILLER_54_950 ();
 sg13g2_fill_1 FILLER_54_966 ();
 sg13g2_decap_8 FILLER_54_1012 ();
 sg13g2_decap_8 FILLER_54_1019 ();
 sg13g2_decap_8 FILLER_54_1026 ();
 sg13g2_decap_8 FILLER_54_1033 ();
 sg13g2_decap_8 FILLER_54_1040 ();
 sg13g2_decap_8 FILLER_54_1047 ();
 sg13g2_decap_8 FILLER_54_1054 ();
 sg13g2_decap_8 FILLER_54_1061 ();
 sg13g2_decap_8 FILLER_54_1068 ();
 sg13g2_decap_8 FILLER_54_1075 ();
 sg13g2_decap_8 FILLER_54_1082 ();
 sg13g2_decap_8 FILLER_54_1089 ();
 sg13g2_decap_8 FILLER_54_1096 ();
 sg13g2_decap_8 FILLER_54_1103 ();
 sg13g2_decap_8 FILLER_54_1110 ();
 sg13g2_decap_8 FILLER_54_1117 ();
 sg13g2_decap_8 FILLER_54_1124 ();
 sg13g2_decap_8 FILLER_54_1131 ();
 sg13g2_decap_8 FILLER_54_1138 ();
 sg13g2_decap_8 FILLER_54_1145 ();
 sg13g2_decap_8 FILLER_54_1152 ();
 sg13g2_decap_8 FILLER_54_1159 ();
 sg13g2_decap_8 FILLER_54_1166 ();
 sg13g2_decap_8 FILLER_54_1173 ();
 sg13g2_decap_8 FILLER_54_1180 ();
 sg13g2_decap_8 FILLER_54_1187 ();
 sg13g2_decap_8 FILLER_54_1194 ();
 sg13g2_decap_8 FILLER_54_1201 ();
 sg13g2_decap_8 FILLER_54_1208 ();
 sg13g2_decap_8 FILLER_54_1215 ();
 sg13g2_decap_8 FILLER_54_1222 ();
 sg13g2_decap_8 FILLER_54_1229 ();
 sg13g2_decap_8 FILLER_54_1236 ();
 sg13g2_decap_8 FILLER_54_1243 ();
 sg13g2_decap_8 FILLER_54_1250 ();
 sg13g2_decap_8 FILLER_54_1257 ();
 sg13g2_decap_8 FILLER_54_1264 ();
 sg13g2_decap_8 FILLER_54_1271 ();
 sg13g2_decap_8 FILLER_54_1278 ();
 sg13g2_decap_8 FILLER_54_1285 ();
 sg13g2_decap_8 FILLER_54_1292 ();
 sg13g2_decap_8 FILLER_54_1299 ();
 sg13g2_decap_8 FILLER_54_1306 ();
 sg13g2_decap_8 FILLER_54_1313 ();
 sg13g2_decap_8 FILLER_54_1320 ();
 sg13g2_decap_8 FILLER_54_1327 ();
 sg13g2_decap_8 FILLER_54_1334 ();
 sg13g2_decap_8 FILLER_54_1341 ();
 sg13g2_decap_8 FILLER_54_1348 ();
 sg13g2_decap_8 FILLER_54_1355 ();
 sg13g2_decap_8 FILLER_54_1362 ();
 sg13g2_decap_8 FILLER_54_1369 ();
 sg13g2_decap_8 FILLER_54_1376 ();
 sg13g2_decap_8 FILLER_54_1383 ();
 sg13g2_decap_8 FILLER_54_1390 ();
 sg13g2_decap_8 FILLER_54_1397 ();
 sg13g2_decap_8 FILLER_54_1404 ();
 sg13g2_decap_8 FILLER_54_1411 ();
 sg13g2_decap_8 FILLER_54_1418 ();
 sg13g2_decap_8 FILLER_54_1425 ();
 sg13g2_decap_8 FILLER_54_1432 ();
 sg13g2_decap_8 FILLER_54_1439 ();
 sg13g2_decap_8 FILLER_54_1446 ();
 sg13g2_decap_8 FILLER_54_1453 ();
 sg13g2_decap_8 FILLER_54_1460 ();
 sg13g2_decap_8 FILLER_54_1467 ();
 sg13g2_decap_8 FILLER_54_1474 ();
 sg13g2_decap_8 FILLER_54_1481 ();
 sg13g2_decap_8 FILLER_54_1488 ();
 sg13g2_decap_8 FILLER_54_1495 ();
 sg13g2_decap_8 FILLER_54_1502 ();
 sg13g2_decap_8 FILLER_54_1509 ();
 sg13g2_decap_8 FILLER_54_1516 ();
 sg13g2_decap_8 FILLER_54_1523 ();
 sg13g2_decap_8 FILLER_54_1530 ();
 sg13g2_decap_8 FILLER_54_1537 ();
 sg13g2_decap_8 FILLER_54_1544 ();
 sg13g2_decap_8 FILLER_54_1551 ();
 sg13g2_decap_8 FILLER_54_1558 ();
 sg13g2_decap_8 FILLER_54_1565 ();
 sg13g2_decap_8 FILLER_54_1572 ();
 sg13g2_decap_8 FILLER_54_1579 ();
 sg13g2_decap_8 FILLER_54_1586 ();
 sg13g2_decap_8 FILLER_54_1593 ();
 sg13g2_decap_8 FILLER_54_1600 ();
 sg13g2_decap_8 FILLER_54_1607 ();
 sg13g2_decap_8 FILLER_54_1614 ();
 sg13g2_decap_8 FILLER_54_1621 ();
 sg13g2_decap_8 FILLER_54_1628 ();
 sg13g2_decap_8 FILLER_54_1635 ();
 sg13g2_decap_8 FILLER_54_1642 ();
 sg13g2_decap_8 FILLER_54_1649 ();
 sg13g2_decap_8 FILLER_54_1656 ();
 sg13g2_decap_8 FILLER_54_1663 ();
 sg13g2_decap_8 FILLER_54_1670 ();
 sg13g2_decap_8 FILLER_54_1677 ();
 sg13g2_decap_8 FILLER_54_1684 ();
 sg13g2_decap_8 FILLER_54_1691 ();
 sg13g2_decap_8 FILLER_54_1698 ();
 sg13g2_decap_8 FILLER_54_1705 ();
 sg13g2_decap_8 FILLER_54_1712 ();
 sg13g2_decap_8 FILLER_54_1719 ();
 sg13g2_decap_8 FILLER_54_1726 ();
 sg13g2_decap_8 FILLER_54_1733 ();
 sg13g2_decap_8 FILLER_54_1740 ();
 sg13g2_decap_8 FILLER_54_1747 ();
 sg13g2_decap_8 FILLER_54_1754 ();
 sg13g2_decap_8 FILLER_54_1761 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_decap_8 FILLER_55_7 ();
 sg13g2_decap_8 FILLER_55_14 ();
 sg13g2_decap_8 FILLER_55_21 ();
 sg13g2_decap_8 FILLER_55_28 ();
 sg13g2_decap_8 FILLER_55_35 ();
 sg13g2_decap_8 FILLER_55_42 ();
 sg13g2_decap_8 FILLER_55_49 ();
 sg13g2_decap_8 FILLER_55_56 ();
 sg13g2_fill_2 FILLER_55_63 ();
 sg13g2_fill_1 FILLER_55_65 ();
 sg13g2_fill_1 FILLER_55_92 ();
 sg13g2_fill_1 FILLER_55_106 ();
 sg13g2_fill_1 FILLER_55_147 ();
 sg13g2_fill_1 FILLER_55_174 ();
 sg13g2_fill_2 FILLER_55_236 ();
 sg13g2_fill_1 FILLER_55_261 ();
 sg13g2_fill_2 FILLER_55_284 ();
 sg13g2_fill_1 FILLER_55_286 ();
 sg13g2_decap_4 FILLER_55_327 ();
 sg13g2_fill_1 FILLER_55_331 ();
 sg13g2_fill_2 FILLER_55_375 ();
 sg13g2_fill_2 FILLER_55_425 ();
 sg13g2_fill_1 FILLER_55_427 ();
 sg13g2_fill_2 FILLER_55_463 ();
 sg13g2_fill_2 FILLER_55_491 ();
 sg13g2_fill_1 FILLER_55_493 ();
 sg13g2_fill_2 FILLER_55_507 ();
 sg13g2_fill_1 FILLER_55_523 ();
 sg13g2_fill_2 FILLER_55_547 ();
 sg13g2_fill_1 FILLER_55_549 ();
 sg13g2_decap_4 FILLER_55_574 ();
 sg13g2_fill_1 FILLER_55_578 ();
 sg13g2_fill_2 FILLER_55_591 ();
 sg13g2_fill_1 FILLER_55_601 ();
 sg13g2_fill_2 FILLER_55_630 ();
 sg13g2_fill_1 FILLER_55_640 ();
 sg13g2_decap_4 FILLER_55_677 ();
 sg13g2_fill_2 FILLER_55_681 ();
 sg13g2_fill_2 FILLER_55_705 ();
 sg13g2_fill_2 FILLER_55_715 ();
 sg13g2_fill_2 FILLER_55_762 ();
 sg13g2_fill_1 FILLER_55_764 ();
 sg13g2_decap_4 FILLER_55_787 ();
 sg13g2_fill_1 FILLER_55_791 ();
 sg13g2_fill_1 FILLER_55_818 ();
 sg13g2_fill_1 FILLER_55_837 ();
 sg13g2_fill_2 FILLER_55_880 ();
 sg13g2_decap_8 FILLER_55_890 ();
 sg13g2_fill_2 FILLER_55_897 ();
 sg13g2_decap_8 FILLER_55_908 ();
 sg13g2_decap_8 FILLER_55_915 ();
 sg13g2_fill_2 FILLER_55_922 ();
 sg13g2_fill_2 FILLER_55_938 ();
 sg13g2_fill_1 FILLER_55_940 ();
 sg13g2_fill_2 FILLER_55_973 ();
 sg13g2_fill_1 FILLER_55_975 ();
 sg13g2_fill_2 FILLER_55_987 ();
 sg13g2_decap_8 FILLER_55_1023 ();
 sg13g2_decap_8 FILLER_55_1030 ();
 sg13g2_decap_8 FILLER_55_1037 ();
 sg13g2_decap_8 FILLER_55_1044 ();
 sg13g2_decap_8 FILLER_55_1051 ();
 sg13g2_decap_8 FILLER_55_1058 ();
 sg13g2_decap_8 FILLER_55_1065 ();
 sg13g2_decap_8 FILLER_55_1072 ();
 sg13g2_decap_8 FILLER_55_1079 ();
 sg13g2_decap_8 FILLER_55_1086 ();
 sg13g2_decap_8 FILLER_55_1093 ();
 sg13g2_decap_8 FILLER_55_1100 ();
 sg13g2_decap_8 FILLER_55_1107 ();
 sg13g2_decap_8 FILLER_55_1114 ();
 sg13g2_decap_8 FILLER_55_1121 ();
 sg13g2_decap_8 FILLER_55_1128 ();
 sg13g2_decap_8 FILLER_55_1135 ();
 sg13g2_decap_8 FILLER_55_1142 ();
 sg13g2_decap_8 FILLER_55_1149 ();
 sg13g2_decap_8 FILLER_55_1156 ();
 sg13g2_decap_8 FILLER_55_1163 ();
 sg13g2_decap_8 FILLER_55_1170 ();
 sg13g2_decap_8 FILLER_55_1177 ();
 sg13g2_decap_8 FILLER_55_1184 ();
 sg13g2_decap_8 FILLER_55_1191 ();
 sg13g2_decap_8 FILLER_55_1198 ();
 sg13g2_decap_8 FILLER_55_1205 ();
 sg13g2_decap_8 FILLER_55_1212 ();
 sg13g2_decap_8 FILLER_55_1219 ();
 sg13g2_decap_8 FILLER_55_1226 ();
 sg13g2_decap_8 FILLER_55_1233 ();
 sg13g2_decap_8 FILLER_55_1240 ();
 sg13g2_decap_8 FILLER_55_1247 ();
 sg13g2_decap_8 FILLER_55_1254 ();
 sg13g2_decap_8 FILLER_55_1261 ();
 sg13g2_decap_8 FILLER_55_1268 ();
 sg13g2_decap_8 FILLER_55_1275 ();
 sg13g2_decap_8 FILLER_55_1282 ();
 sg13g2_decap_8 FILLER_55_1289 ();
 sg13g2_decap_8 FILLER_55_1296 ();
 sg13g2_decap_8 FILLER_55_1303 ();
 sg13g2_decap_8 FILLER_55_1310 ();
 sg13g2_decap_8 FILLER_55_1317 ();
 sg13g2_decap_8 FILLER_55_1324 ();
 sg13g2_decap_8 FILLER_55_1331 ();
 sg13g2_decap_8 FILLER_55_1338 ();
 sg13g2_decap_8 FILLER_55_1345 ();
 sg13g2_decap_8 FILLER_55_1352 ();
 sg13g2_decap_8 FILLER_55_1359 ();
 sg13g2_decap_8 FILLER_55_1366 ();
 sg13g2_decap_8 FILLER_55_1373 ();
 sg13g2_decap_8 FILLER_55_1380 ();
 sg13g2_decap_8 FILLER_55_1387 ();
 sg13g2_decap_8 FILLER_55_1394 ();
 sg13g2_decap_8 FILLER_55_1401 ();
 sg13g2_decap_8 FILLER_55_1408 ();
 sg13g2_decap_8 FILLER_55_1415 ();
 sg13g2_decap_8 FILLER_55_1422 ();
 sg13g2_decap_8 FILLER_55_1429 ();
 sg13g2_decap_8 FILLER_55_1436 ();
 sg13g2_decap_8 FILLER_55_1443 ();
 sg13g2_decap_8 FILLER_55_1450 ();
 sg13g2_decap_8 FILLER_55_1457 ();
 sg13g2_decap_8 FILLER_55_1464 ();
 sg13g2_decap_8 FILLER_55_1471 ();
 sg13g2_decap_8 FILLER_55_1478 ();
 sg13g2_decap_8 FILLER_55_1485 ();
 sg13g2_decap_8 FILLER_55_1492 ();
 sg13g2_decap_8 FILLER_55_1499 ();
 sg13g2_decap_8 FILLER_55_1506 ();
 sg13g2_decap_8 FILLER_55_1513 ();
 sg13g2_decap_8 FILLER_55_1520 ();
 sg13g2_decap_8 FILLER_55_1527 ();
 sg13g2_decap_8 FILLER_55_1534 ();
 sg13g2_decap_8 FILLER_55_1541 ();
 sg13g2_decap_8 FILLER_55_1548 ();
 sg13g2_decap_8 FILLER_55_1555 ();
 sg13g2_decap_8 FILLER_55_1562 ();
 sg13g2_decap_8 FILLER_55_1569 ();
 sg13g2_decap_8 FILLER_55_1576 ();
 sg13g2_decap_8 FILLER_55_1583 ();
 sg13g2_decap_8 FILLER_55_1590 ();
 sg13g2_decap_8 FILLER_55_1597 ();
 sg13g2_decap_8 FILLER_55_1604 ();
 sg13g2_decap_8 FILLER_55_1611 ();
 sg13g2_decap_8 FILLER_55_1618 ();
 sg13g2_decap_8 FILLER_55_1625 ();
 sg13g2_decap_8 FILLER_55_1632 ();
 sg13g2_decap_8 FILLER_55_1639 ();
 sg13g2_decap_8 FILLER_55_1646 ();
 sg13g2_decap_8 FILLER_55_1653 ();
 sg13g2_decap_8 FILLER_55_1660 ();
 sg13g2_decap_8 FILLER_55_1667 ();
 sg13g2_decap_8 FILLER_55_1674 ();
 sg13g2_decap_8 FILLER_55_1681 ();
 sg13g2_decap_8 FILLER_55_1688 ();
 sg13g2_decap_8 FILLER_55_1695 ();
 sg13g2_decap_8 FILLER_55_1702 ();
 sg13g2_decap_8 FILLER_55_1709 ();
 sg13g2_decap_8 FILLER_55_1716 ();
 sg13g2_decap_8 FILLER_55_1723 ();
 sg13g2_decap_8 FILLER_55_1730 ();
 sg13g2_decap_8 FILLER_55_1737 ();
 sg13g2_decap_8 FILLER_55_1744 ();
 sg13g2_decap_8 FILLER_55_1751 ();
 sg13g2_decap_8 FILLER_55_1758 ();
 sg13g2_fill_2 FILLER_55_1765 ();
 sg13g2_fill_1 FILLER_55_1767 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_decap_8 FILLER_56_7 ();
 sg13g2_decap_8 FILLER_56_14 ();
 sg13g2_decap_8 FILLER_56_21 ();
 sg13g2_decap_8 FILLER_56_28 ();
 sg13g2_decap_8 FILLER_56_35 ();
 sg13g2_decap_8 FILLER_56_42 ();
 sg13g2_decap_8 FILLER_56_49 ();
 sg13g2_decap_8 FILLER_56_56 ();
 sg13g2_fill_1 FILLER_56_63 ();
 sg13g2_fill_1 FILLER_56_186 ();
 sg13g2_fill_1 FILLER_56_213 ();
 sg13g2_fill_2 FILLER_56_287 ();
 sg13g2_fill_1 FILLER_56_289 ();
 sg13g2_fill_1 FILLER_56_349 ();
 sg13g2_fill_2 FILLER_56_410 ();
 sg13g2_fill_1 FILLER_56_464 ();
 sg13g2_fill_1 FILLER_56_526 ();
 sg13g2_fill_1 FILLER_56_570 ();
 sg13g2_fill_1 FILLER_56_577 ();
 sg13g2_decap_8 FILLER_56_585 ();
 sg13g2_fill_2 FILLER_56_592 ();
 sg13g2_decap_4 FILLER_56_603 ();
 sg13g2_fill_2 FILLER_56_607 ();
 sg13g2_fill_2 FILLER_56_619 ();
 sg13g2_fill_1 FILLER_56_621 ();
 sg13g2_fill_1 FILLER_56_628 ();
 sg13g2_fill_2 FILLER_56_678 ();
 sg13g2_fill_1 FILLER_56_680 ();
 sg13g2_fill_2 FILLER_56_686 ();
 sg13g2_fill_1 FILLER_56_692 ();
 sg13g2_decap_4 FILLER_56_716 ();
 sg13g2_fill_1 FILLER_56_720 ();
 sg13g2_fill_2 FILLER_56_734 ();
 sg13g2_fill_2 FILLER_56_741 ();
 sg13g2_fill_2 FILLER_56_748 ();
 sg13g2_fill_2 FILLER_56_756 ();
 sg13g2_fill_1 FILLER_56_762 ();
 sg13g2_fill_2 FILLER_56_775 ();
 sg13g2_decap_8 FILLER_56_802 ();
 sg13g2_fill_1 FILLER_56_809 ();
 sg13g2_decap_8 FILLER_56_879 ();
 sg13g2_decap_8 FILLER_56_886 ();
 sg13g2_decap_8 FILLER_56_893 ();
 sg13g2_decap_8 FILLER_56_900 ();
 sg13g2_fill_2 FILLER_56_907 ();
 sg13g2_fill_1 FILLER_56_909 ();
 sg13g2_fill_1 FILLER_56_941 ();
 sg13g2_decap_8 FILLER_56_1027 ();
 sg13g2_decap_8 FILLER_56_1034 ();
 sg13g2_decap_8 FILLER_56_1041 ();
 sg13g2_decap_8 FILLER_56_1048 ();
 sg13g2_decap_8 FILLER_56_1055 ();
 sg13g2_decap_8 FILLER_56_1062 ();
 sg13g2_decap_8 FILLER_56_1069 ();
 sg13g2_decap_8 FILLER_56_1076 ();
 sg13g2_decap_8 FILLER_56_1083 ();
 sg13g2_decap_8 FILLER_56_1090 ();
 sg13g2_decap_8 FILLER_56_1097 ();
 sg13g2_decap_8 FILLER_56_1104 ();
 sg13g2_decap_8 FILLER_56_1111 ();
 sg13g2_decap_8 FILLER_56_1118 ();
 sg13g2_decap_8 FILLER_56_1125 ();
 sg13g2_decap_8 FILLER_56_1132 ();
 sg13g2_decap_8 FILLER_56_1139 ();
 sg13g2_decap_8 FILLER_56_1146 ();
 sg13g2_decap_8 FILLER_56_1153 ();
 sg13g2_decap_8 FILLER_56_1160 ();
 sg13g2_decap_8 FILLER_56_1167 ();
 sg13g2_decap_8 FILLER_56_1174 ();
 sg13g2_decap_8 FILLER_56_1181 ();
 sg13g2_decap_8 FILLER_56_1188 ();
 sg13g2_decap_8 FILLER_56_1195 ();
 sg13g2_decap_8 FILLER_56_1202 ();
 sg13g2_decap_8 FILLER_56_1209 ();
 sg13g2_decap_8 FILLER_56_1216 ();
 sg13g2_decap_8 FILLER_56_1223 ();
 sg13g2_decap_8 FILLER_56_1230 ();
 sg13g2_decap_8 FILLER_56_1237 ();
 sg13g2_decap_8 FILLER_56_1244 ();
 sg13g2_decap_8 FILLER_56_1251 ();
 sg13g2_decap_8 FILLER_56_1258 ();
 sg13g2_decap_8 FILLER_56_1265 ();
 sg13g2_decap_8 FILLER_56_1272 ();
 sg13g2_decap_8 FILLER_56_1279 ();
 sg13g2_decap_8 FILLER_56_1286 ();
 sg13g2_decap_8 FILLER_56_1293 ();
 sg13g2_decap_8 FILLER_56_1300 ();
 sg13g2_decap_8 FILLER_56_1307 ();
 sg13g2_decap_8 FILLER_56_1314 ();
 sg13g2_decap_8 FILLER_56_1321 ();
 sg13g2_decap_8 FILLER_56_1328 ();
 sg13g2_decap_8 FILLER_56_1335 ();
 sg13g2_decap_8 FILLER_56_1342 ();
 sg13g2_decap_8 FILLER_56_1349 ();
 sg13g2_decap_8 FILLER_56_1356 ();
 sg13g2_decap_8 FILLER_56_1363 ();
 sg13g2_decap_8 FILLER_56_1370 ();
 sg13g2_decap_8 FILLER_56_1377 ();
 sg13g2_decap_8 FILLER_56_1384 ();
 sg13g2_decap_8 FILLER_56_1391 ();
 sg13g2_decap_8 FILLER_56_1398 ();
 sg13g2_decap_8 FILLER_56_1405 ();
 sg13g2_decap_8 FILLER_56_1412 ();
 sg13g2_decap_8 FILLER_56_1419 ();
 sg13g2_decap_8 FILLER_56_1426 ();
 sg13g2_decap_8 FILLER_56_1433 ();
 sg13g2_decap_8 FILLER_56_1440 ();
 sg13g2_decap_8 FILLER_56_1447 ();
 sg13g2_decap_8 FILLER_56_1454 ();
 sg13g2_decap_8 FILLER_56_1461 ();
 sg13g2_decap_8 FILLER_56_1468 ();
 sg13g2_decap_8 FILLER_56_1475 ();
 sg13g2_decap_8 FILLER_56_1482 ();
 sg13g2_decap_8 FILLER_56_1489 ();
 sg13g2_decap_8 FILLER_56_1496 ();
 sg13g2_decap_8 FILLER_56_1503 ();
 sg13g2_decap_8 FILLER_56_1510 ();
 sg13g2_decap_8 FILLER_56_1517 ();
 sg13g2_decap_8 FILLER_56_1524 ();
 sg13g2_decap_8 FILLER_56_1531 ();
 sg13g2_decap_8 FILLER_56_1538 ();
 sg13g2_decap_8 FILLER_56_1545 ();
 sg13g2_decap_8 FILLER_56_1552 ();
 sg13g2_decap_8 FILLER_56_1559 ();
 sg13g2_decap_8 FILLER_56_1566 ();
 sg13g2_decap_8 FILLER_56_1573 ();
 sg13g2_decap_8 FILLER_56_1580 ();
 sg13g2_decap_8 FILLER_56_1587 ();
 sg13g2_decap_8 FILLER_56_1594 ();
 sg13g2_decap_8 FILLER_56_1601 ();
 sg13g2_decap_8 FILLER_56_1608 ();
 sg13g2_decap_8 FILLER_56_1615 ();
 sg13g2_decap_8 FILLER_56_1622 ();
 sg13g2_decap_8 FILLER_56_1629 ();
 sg13g2_decap_8 FILLER_56_1636 ();
 sg13g2_decap_8 FILLER_56_1643 ();
 sg13g2_decap_8 FILLER_56_1650 ();
 sg13g2_decap_8 FILLER_56_1657 ();
 sg13g2_decap_8 FILLER_56_1664 ();
 sg13g2_decap_8 FILLER_56_1671 ();
 sg13g2_decap_8 FILLER_56_1678 ();
 sg13g2_decap_8 FILLER_56_1685 ();
 sg13g2_decap_8 FILLER_56_1692 ();
 sg13g2_decap_8 FILLER_56_1699 ();
 sg13g2_decap_8 FILLER_56_1706 ();
 sg13g2_decap_8 FILLER_56_1713 ();
 sg13g2_decap_8 FILLER_56_1720 ();
 sg13g2_decap_8 FILLER_56_1727 ();
 sg13g2_decap_8 FILLER_56_1734 ();
 sg13g2_decap_8 FILLER_56_1741 ();
 sg13g2_decap_8 FILLER_56_1748 ();
 sg13g2_decap_8 FILLER_56_1755 ();
 sg13g2_decap_4 FILLER_56_1762 ();
 sg13g2_fill_2 FILLER_56_1766 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_decap_8 FILLER_57_7 ();
 sg13g2_decap_8 FILLER_57_14 ();
 sg13g2_decap_8 FILLER_57_21 ();
 sg13g2_decap_8 FILLER_57_28 ();
 sg13g2_decap_8 FILLER_57_35 ();
 sg13g2_decap_8 FILLER_57_42 ();
 sg13g2_decap_8 FILLER_57_49 ();
 sg13g2_decap_8 FILLER_57_56 ();
 sg13g2_decap_8 FILLER_57_63 ();
 sg13g2_fill_2 FILLER_57_70 ();
 sg13g2_decap_4 FILLER_57_75 ();
 sg13g2_fill_1 FILLER_57_79 ();
 sg13g2_fill_1 FILLER_57_92 ();
 sg13g2_fill_1 FILLER_57_98 ();
 sg13g2_fill_1 FILLER_57_107 ();
 sg13g2_fill_2 FILLER_57_116 ();
 sg13g2_fill_1 FILLER_57_152 ();
 sg13g2_fill_2 FILLER_57_158 ();
 sg13g2_fill_2 FILLER_57_165 ();
 sg13g2_fill_1 FILLER_57_202 ();
 sg13g2_fill_2 FILLER_57_213 ();
 sg13g2_fill_1 FILLER_57_229 ();
 sg13g2_fill_2 FILLER_57_253 ();
 sg13g2_fill_2 FILLER_57_321 ();
 sg13g2_fill_1 FILLER_57_323 ();
 sg13g2_fill_2 FILLER_57_377 ();
 sg13g2_fill_1 FILLER_57_399 ();
 sg13g2_decap_8 FILLER_57_440 ();
 sg13g2_fill_1 FILLER_57_447 ();
 sg13g2_decap_8 FILLER_57_453 ();
 sg13g2_fill_2 FILLER_57_460 ();
 sg13g2_decap_4 FILLER_57_480 ();
 sg13g2_fill_2 FILLER_57_528 ();
 sg13g2_fill_1 FILLER_57_530 ();
 sg13g2_decap_8 FILLER_57_543 ();
 sg13g2_fill_1 FILLER_57_550 ();
 sg13g2_fill_1 FILLER_57_559 ();
 sg13g2_fill_1 FILLER_57_565 ();
 sg13g2_decap_4 FILLER_57_571 ();
 sg13g2_fill_2 FILLER_57_575 ();
 sg13g2_fill_2 FILLER_57_593 ();
 sg13g2_fill_2 FILLER_57_600 ();
 sg13g2_fill_1 FILLER_57_602 ();
 sg13g2_fill_2 FILLER_57_615 ();
 sg13g2_fill_2 FILLER_57_627 ();
 sg13g2_fill_2 FILLER_57_634 ();
 sg13g2_decap_4 FILLER_57_655 ();
 sg13g2_decap_4 FILLER_57_664 ();
 sg13g2_decap_4 FILLER_57_692 ();
 sg13g2_fill_2 FILLER_57_696 ();
 sg13g2_decap_4 FILLER_57_710 ();
 sg13g2_fill_2 FILLER_57_714 ();
 sg13g2_fill_1 FILLER_57_721 ();
 sg13g2_fill_2 FILLER_57_730 ();
 sg13g2_fill_2 FILLER_57_767 ();
 sg13g2_fill_1 FILLER_57_769 ();
 sg13g2_decap_8 FILLER_57_788 ();
 sg13g2_decap_4 FILLER_57_805 ();
 sg13g2_fill_1 FILLER_57_809 ();
 sg13g2_decap_4 FILLER_57_836 ();
 sg13g2_fill_1 FILLER_57_840 ();
 sg13g2_decap_4 FILLER_57_856 ();
 sg13g2_decap_8 FILLER_57_869 ();
 sg13g2_decap_8 FILLER_57_876 ();
 sg13g2_decap_8 FILLER_57_883 ();
 sg13g2_decap_4 FILLER_57_890 ();
 sg13g2_decap_8 FILLER_57_899 ();
 sg13g2_decap_8 FILLER_57_906 ();
 sg13g2_decap_4 FILLER_57_913 ();
 sg13g2_fill_2 FILLER_57_917 ();
 sg13g2_fill_1 FILLER_57_944 ();
 sg13g2_fill_1 FILLER_57_954 ();
 sg13g2_decap_8 FILLER_57_1032 ();
 sg13g2_decap_8 FILLER_57_1039 ();
 sg13g2_decap_8 FILLER_57_1046 ();
 sg13g2_decap_8 FILLER_57_1053 ();
 sg13g2_decap_8 FILLER_57_1060 ();
 sg13g2_decap_8 FILLER_57_1067 ();
 sg13g2_decap_8 FILLER_57_1074 ();
 sg13g2_decap_8 FILLER_57_1081 ();
 sg13g2_decap_8 FILLER_57_1088 ();
 sg13g2_decap_8 FILLER_57_1095 ();
 sg13g2_decap_8 FILLER_57_1102 ();
 sg13g2_decap_8 FILLER_57_1109 ();
 sg13g2_decap_8 FILLER_57_1116 ();
 sg13g2_decap_8 FILLER_57_1123 ();
 sg13g2_decap_8 FILLER_57_1130 ();
 sg13g2_decap_8 FILLER_57_1137 ();
 sg13g2_decap_8 FILLER_57_1144 ();
 sg13g2_decap_8 FILLER_57_1151 ();
 sg13g2_decap_8 FILLER_57_1158 ();
 sg13g2_decap_8 FILLER_57_1165 ();
 sg13g2_decap_8 FILLER_57_1172 ();
 sg13g2_decap_8 FILLER_57_1179 ();
 sg13g2_decap_8 FILLER_57_1186 ();
 sg13g2_decap_8 FILLER_57_1193 ();
 sg13g2_decap_8 FILLER_57_1200 ();
 sg13g2_decap_8 FILLER_57_1207 ();
 sg13g2_decap_8 FILLER_57_1214 ();
 sg13g2_decap_8 FILLER_57_1221 ();
 sg13g2_decap_8 FILLER_57_1228 ();
 sg13g2_decap_8 FILLER_57_1235 ();
 sg13g2_decap_8 FILLER_57_1242 ();
 sg13g2_decap_8 FILLER_57_1249 ();
 sg13g2_decap_8 FILLER_57_1256 ();
 sg13g2_decap_8 FILLER_57_1263 ();
 sg13g2_decap_8 FILLER_57_1270 ();
 sg13g2_decap_8 FILLER_57_1277 ();
 sg13g2_decap_8 FILLER_57_1284 ();
 sg13g2_decap_8 FILLER_57_1291 ();
 sg13g2_decap_8 FILLER_57_1298 ();
 sg13g2_decap_8 FILLER_57_1305 ();
 sg13g2_decap_8 FILLER_57_1312 ();
 sg13g2_decap_8 FILLER_57_1319 ();
 sg13g2_decap_8 FILLER_57_1326 ();
 sg13g2_decap_8 FILLER_57_1333 ();
 sg13g2_decap_8 FILLER_57_1340 ();
 sg13g2_decap_8 FILLER_57_1347 ();
 sg13g2_decap_8 FILLER_57_1354 ();
 sg13g2_decap_8 FILLER_57_1361 ();
 sg13g2_decap_8 FILLER_57_1368 ();
 sg13g2_decap_8 FILLER_57_1375 ();
 sg13g2_decap_8 FILLER_57_1382 ();
 sg13g2_decap_8 FILLER_57_1389 ();
 sg13g2_decap_8 FILLER_57_1396 ();
 sg13g2_decap_8 FILLER_57_1403 ();
 sg13g2_decap_8 FILLER_57_1410 ();
 sg13g2_decap_8 FILLER_57_1417 ();
 sg13g2_decap_8 FILLER_57_1424 ();
 sg13g2_decap_8 FILLER_57_1431 ();
 sg13g2_decap_8 FILLER_57_1438 ();
 sg13g2_decap_8 FILLER_57_1445 ();
 sg13g2_decap_8 FILLER_57_1452 ();
 sg13g2_decap_8 FILLER_57_1459 ();
 sg13g2_decap_8 FILLER_57_1466 ();
 sg13g2_decap_8 FILLER_57_1473 ();
 sg13g2_decap_8 FILLER_57_1480 ();
 sg13g2_decap_8 FILLER_57_1487 ();
 sg13g2_decap_8 FILLER_57_1494 ();
 sg13g2_decap_8 FILLER_57_1501 ();
 sg13g2_decap_8 FILLER_57_1508 ();
 sg13g2_decap_8 FILLER_57_1515 ();
 sg13g2_decap_8 FILLER_57_1522 ();
 sg13g2_decap_8 FILLER_57_1529 ();
 sg13g2_decap_8 FILLER_57_1536 ();
 sg13g2_decap_8 FILLER_57_1543 ();
 sg13g2_decap_8 FILLER_57_1550 ();
 sg13g2_decap_8 FILLER_57_1557 ();
 sg13g2_decap_8 FILLER_57_1564 ();
 sg13g2_decap_8 FILLER_57_1571 ();
 sg13g2_decap_8 FILLER_57_1578 ();
 sg13g2_decap_8 FILLER_57_1585 ();
 sg13g2_decap_8 FILLER_57_1592 ();
 sg13g2_decap_8 FILLER_57_1599 ();
 sg13g2_decap_8 FILLER_57_1606 ();
 sg13g2_decap_8 FILLER_57_1613 ();
 sg13g2_decap_8 FILLER_57_1620 ();
 sg13g2_decap_8 FILLER_57_1627 ();
 sg13g2_decap_8 FILLER_57_1634 ();
 sg13g2_decap_8 FILLER_57_1641 ();
 sg13g2_decap_8 FILLER_57_1648 ();
 sg13g2_decap_8 FILLER_57_1655 ();
 sg13g2_decap_8 FILLER_57_1662 ();
 sg13g2_decap_8 FILLER_57_1669 ();
 sg13g2_decap_8 FILLER_57_1676 ();
 sg13g2_decap_8 FILLER_57_1683 ();
 sg13g2_decap_8 FILLER_57_1690 ();
 sg13g2_decap_8 FILLER_57_1697 ();
 sg13g2_decap_8 FILLER_57_1704 ();
 sg13g2_decap_8 FILLER_57_1711 ();
 sg13g2_decap_8 FILLER_57_1718 ();
 sg13g2_decap_8 FILLER_57_1725 ();
 sg13g2_decap_8 FILLER_57_1732 ();
 sg13g2_decap_8 FILLER_57_1739 ();
 sg13g2_decap_8 FILLER_57_1746 ();
 sg13g2_decap_8 FILLER_57_1753 ();
 sg13g2_decap_8 FILLER_57_1760 ();
 sg13g2_fill_1 FILLER_57_1767 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_decap_8 FILLER_58_7 ();
 sg13g2_decap_8 FILLER_58_14 ();
 sg13g2_decap_8 FILLER_58_21 ();
 sg13g2_decap_8 FILLER_58_28 ();
 sg13g2_decap_8 FILLER_58_35 ();
 sg13g2_decap_8 FILLER_58_42 ();
 sg13g2_decap_8 FILLER_58_49 ();
 sg13g2_decap_8 FILLER_58_56 ();
 sg13g2_decap_8 FILLER_58_63 ();
 sg13g2_decap_4 FILLER_58_70 ();
 sg13g2_fill_1 FILLER_58_74 ();
 sg13g2_fill_1 FILLER_58_130 ();
 sg13g2_fill_2 FILLER_58_140 ();
 sg13g2_fill_1 FILLER_58_181 ();
 sg13g2_fill_2 FILLER_58_192 ();
 sg13g2_fill_2 FILLER_58_257 ();
 sg13g2_fill_2 FILLER_58_273 ();
 sg13g2_fill_1 FILLER_58_383 ();
 sg13g2_decap_8 FILLER_58_397 ();
 sg13g2_decap_4 FILLER_58_443 ();
 sg13g2_fill_1 FILLER_58_447 ();
 sg13g2_decap_8 FILLER_58_461 ();
 sg13g2_decap_8 FILLER_58_468 ();
 sg13g2_decap_8 FILLER_58_475 ();
 sg13g2_decap_4 FILLER_58_482 ();
 sg13g2_fill_1 FILLER_58_525 ();
 sg13g2_fill_1 FILLER_58_583 ();
 sg13g2_fill_2 FILLER_58_595 ();
 sg13g2_fill_1 FILLER_58_597 ();
 sg13g2_decap_8 FILLER_58_631 ();
 sg13g2_fill_2 FILLER_58_662 ();
 sg13g2_fill_1 FILLER_58_664 ();
 sg13g2_fill_1 FILLER_58_692 ();
 sg13g2_fill_2 FILLER_58_702 ();
 sg13g2_fill_2 FILLER_58_721 ();
 sg13g2_fill_1 FILLER_58_723 ();
 sg13g2_fill_2 FILLER_58_729 ();
 sg13g2_fill_1 FILLER_58_731 ();
 sg13g2_fill_1 FILLER_58_778 ();
 sg13g2_decap_4 FILLER_58_792 ();
 sg13g2_fill_2 FILLER_58_806 ();
 sg13g2_fill_1 FILLER_58_808 ();
 sg13g2_fill_2 FILLER_58_819 ();
 sg13g2_fill_1 FILLER_58_821 ();
 sg13g2_decap_8 FILLER_58_904 ();
 sg13g2_decap_8 FILLER_58_911 ();
 sg13g2_decap_8 FILLER_58_918 ();
 sg13g2_decap_4 FILLER_58_925 ();
 sg13g2_fill_2 FILLER_58_970 ();
 sg13g2_fill_1 FILLER_58_989 ();
 sg13g2_decap_4 FILLER_58_1028 ();
 sg13g2_decap_8 FILLER_58_1044 ();
 sg13g2_decap_4 FILLER_58_1051 ();
 sg13g2_decap_8 FILLER_58_1064 ();
 sg13g2_decap_8 FILLER_58_1071 ();
 sg13g2_decap_8 FILLER_58_1078 ();
 sg13g2_decap_8 FILLER_58_1085 ();
 sg13g2_decap_8 FILLER_58_1092 ();
 sg13g2_decap_8 FILLER_58_1099 ();
 sg13g2_decap_8 FILLER_58_1106 ();
 sg13g2_decap_8 FILLER_58_1113 ();
 sg13g2_decap_8 FILLER_58_1120 ();
 sg13g2_decap_8 FILLER_58_1127 ();
 sg13g2_decap_8 FILLER_58_1134 ();
 sg13g2_decap_8 FILLER_58_1141 ();
 sg13g2_decap_8 FILLER_58_1148 ();
 sg13g2_decap_8 FILLER_58_1155 ();
 sg13g2_decap_8 FILLER_58_1162 ();
 sg13g2_decap_8 FILLER_58_1169 ();
 sg13g2_decap_8 FILLER_58_1176 ();
 sg13g2_decap_8 FILLER_58_1183 ();
 sg13g2_decap_8 FILLER_58_1190 ();
 sg13g2_decap_8 FILLER_58_1197 ();
 sg13g2_decap_8 FILLER_58_1204 ();
 sg13g2_decap_8 FILLER_58_1211 ();
 sg13g2_decap_8 FILLER_58_1218 ();
 sg13g2_decap_8 FILLER_58_1225 ();
 sg13g2_decap_8 FILLER_58_1232 ();
 sg13g2_decap_8 FILLER_58_1239 ();
 sg13g2_decap_8 FILLER_58_1246 ();
 sg13g2_decap_8 FILLER_58_1253 ();
 sg13g2_decap_8 FILLER_58_1260 ();
 sg13g2_decap_8 FILLER_58_1267 ();
 sg13g2_decap_8 FILLER_58_1274 ();
 sg13g2_decap_8 FILLER_58_1281 ();
 sg13g2_decap_8 FILLER_58_1288 ();
 sg13g2_decap_8 FILLER_58_1295 ();
 sg13g2_decap_8 FILLER_58_1302 ();
 sg13g2_decap_8 FILLER_58_1309 ();
 sg13g2_decap_8 FILLER_58_1316 ();
 sg13g2_decap_8 FILLER_58_1323 ();
 sg13g2_decap_8 FILLER_58_1330 ();
 sg13g2_decap_8 FILLER_58_1337 ();
 sg13g2_decap_8 FILLER_58_1344 ();
 sg13g2_decap_8 FILLER_58_1351 ();
 sg13g2_decap_8 FILLER_58_1358 ();
 sg13g2_decap_8 FILLER_58_1365 ();
 sg13g2_decap_8 FILLER_58_1372 ();
 sg13g2_decap_8 FILLER_58_1379 ();
 sg13g2_decap_8 FILLER_58_1386 ();
 sg13g2_decap_8 FILLER_58_1393 ();
 sg13g2_decap_8 FILLER_58_1400 ();
 sg13g2_decap_8 FILLER_58_1407 ();
 sg13g2_decap_8 FILLER_58_1414 ();
 sg13g2_decap_8 FILLER_58_1421 ();
 sg13g2_decap_8 FILLER_58_1428 ();
 sg13g2_decap_8 FILLER_58_1435 ();
 sg13g2_decap_8 FILLER_58_1442 ();
 sg13g2_decap_8 FILLER_58_1449 ();
 sg13g2_decap_8 FILLER_58_1456 ();
 sg13g2_decap_8 FILLER_58_1463 ();
 sg13g2_decap_8 FILLER_58_1470 ();
 sg13g2_decap_8 FILLER_58_1477 ();
 sg13g2_decap_8 FILLER_58_1484 ();
 sg13g2_decap_8 FILLER_58_1491 ();
 sg13g2_decap_8 FILLER_58_1498 ();
 sg13g2_decap_8 FILLER_58_1505 ();
 sg13g2_decap_8 FILLER_58_1512 ();
 sg13g2_decap_8 FILLER_58_1519 ();
 sg13g2_decap_8 FILLER_58_1526 ();
 sg13g2_decap_8 FILLER_58_1533 ();
 sg13g2_decap_8 FILLER_58_1540 ();
 sg13g2_decap_8 FILLER_58_1547 ();
 sg13g2_decap_8 FILLER_58_1554 ();
 sg13g2_decap_8 FILLER_58_1561 ();
 sg13g2_decap_8 FILLER_58_1568 ();
 sg13g2_decap_8 FILLER_58_1575 ();
 sg13g2_decap_8 FILLER_58_1582 ();
 sg13g2_decap_8 FILLER_58_1589 ();
 sg13g2_decap_8 FILLER_58_1596 ();
 sg13g2_decap_8 FILLER_58_1603 ();
 sg13g2_decap_8 FILLER_58_1610 ();
 sg13g2_decap_8 FILLER_58_1617 ();
 sg13g2_decap_8 FILLER_58_1624 ();
 sg13g2_decap_8 FILLER_58_1631 ();
 sg13g2_decap_8 FILLER_58_1638 ();
 sg13g2_decap_8 FILLER_58_1645 ();
 sg13g2_decap_8 FILLER_58_1652 ();
 sg13g2_decap_8 FILLER_58_1659 ();
 sg13g2_decap_8 FILLER_58_1666 ();
 sg13g2_decap_8 FILLER_58_1673 ();
 sg13g2_decap_8 FILLER_58_1680 ();
 sg13g2_decap_8 FILLER_58_1687 ();
 sg13g2_decap_8 FILLER_58_1694 ();
 sg13g2_decap_8 FILLER_58_1701 ();
 sg13g2_decap_8 FILLER_58_1708 ();
 sg13g2_decap_8 FILLER_58_1715 ();
 sg13g2_decap_8 FILLER_58_1722 ();
 sg13g2_decap_8 FILLER_58_1729 ();
 sg13g2_decap_8 FILLER_58_1736 ();
 sg13g2_decap_8 FILLER_58_1743 ();
 sg13g2_decap_8 FILLER_58_1750 ();
 sg13g2_decap_8 FILLER_58_1757 ();
 sg13g2_decap_4 FILLER_58_1764 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_decap_8 FILLER_59_7 ();
 sg13g2_decap_8 FILLER_59_14 ();
 sg13g2_decap_8 FILLER_59_21 ();
 sg13g2_decap_8 FILLER_59_28 ();
 sg13g2_decap_8 FILLER_59_35 ();
 sg13g2_decap_8 FILLER_59_42 ();
 sg13g2_decap_8 FILLER_59_49 ();
 sg13g2_decap_8 FILLER_59_56 ();
 sg13g2_decap_8 FILLER_59_63 ();
 sg13g2_decap_4 FILLER_59_70 ();
 sg13g2_decap_4 FILLER_59_109 ();
 sg13g2_fill_2 FILLER_59_148 ();
 sg13g2_fill_2 FILLER_59_178 ();
 sg13g2_fill_1 FILLER_59_242 ();
 sg13g2_fill_1 FILLER_59_252 ();
 sg13g2_fill_2 FILLER_59_330 ();
 sg13g2_fill_2 FILLER_59_360 ();
 sg13g2_fill_1 FILLER_59_362 ();
 sg13g2_fill_2 FILLER_59_372 ();
 sg13g2_decap_8 FILLER_59_410 ();
 sg13g2_decap_8 FILLER_59_417 ();
 sg13g2_decap_8 FILLER_59_424 ();
 sg13g2_fill_2 FILLER_59_462 ();
 sg13g2_fill_1 FILLER_59_464 ();
 sg13g2_fill_2 FILLER_59_506 ();
 sg13g2_fill_2 FILLER_59_514 ();
 sg13g2_fill_1 FILLER_59_516 ();
 sg13g2_fill_2 FILLER_59_532 ();
 sg13g2_decap_4 FILLER_59_543 ();
 sg13g2_fill_1 FILLER_59_547 ();
 sg13g2_decap_8 FILLER_59_570 ();
 sg13g2_fill_2 FILLER_59_577 ();
 sg13g2_fill_1 FILLER_59_587 ();
 sg13g2_decap_4 FILLER_59_598 ();
 sg13g2_decap_4 FILLER_59_608 ();
 sg13g2_fill_1 FILLER_59_612 ();
 sg13g2_fill_1 FILLER_59_642 ();
 sg13g2_fill_2 FILLER_59_672 ();
 sg13g2_fill_1 FILLER_59_674 ();
 sg13g2_fill_2 FILLER_59_685 ();
 sg13g2_fill_1 FILLER_59_687 ();
 sg13g2_decap_8 FILLER_59_702 ();
 sg13g2_fill_1 FILLER_59_709 ();
 sg13g2_fill_2 FILLER_59_726 ();
 sg13g2_decap_8 FILLER_59_745 ();
 sg13g2_decap_4 FILLER_59_752 ();
 sg13g2_fill_2 FILLER_59_790 ();
 sg13g2_decap_4 FILLER_59_818 ();
 sg13g2_fill_2 FILLER_59_822 ();
 sg13g2_fill_1 FILLER_59_833 ();
 sg13g2_decap_4 FILLER_59_843 ();
 sg13g2_fill_1 FILLER_59_847 ();
 sg13g2_decap_4 FILLER_59_855 ();
 sg13g2_fill_2 FILLER_59_873 ();
 sg13g2_fill_2 FILLER_59_885 ();
 sg13g2_fill_1 FILLER_59_887 ();
 sg13g2_fill_2 FILLER_59_968 ();
 sg13g2_decap_8 FILLER_59_1071 ();
 sg13g2_decap_8 FILLER_59_1078 ();
 sg13g2_decap_8 FILLER_59_1085 ();
 sg13g2_decap_8 FILLER_59_1092 ();
 sg13g2_decap_8 FILLER_59_1099 ();
 sg13g2_decap_8 FILLER_59_1106 ();
 sg13g2_decap_8 FILLER_59_1113 ();
 sg13g2_decap_8 FILLER_59_1120 ();
 sg13g2_decap_8 FILLER_59_1127 ();
 sg13g2_decap_8 FILLER_59_1134 ();
 sg13g2_decap_8 FILLER_59_1141 ();
 sg13g2_decap_8 FILLER_59_1148 ();
 sg13g2_decap_8 FILLER_59_1155 ();
 sg13g2_decap_8 FILLER_59_1162 ();
 sg13g2_decap_8 FILLER_59_1169 ();
 sg13g2_decap_8 FILLER_59_1176 ();
 sg13g2_decap_8 FILLER_59_1183 ();
 sg13g2_decap_8 FILLER_59_1190 ();
 sg13g2_decap_8 FILLER_59_1197 ();
 sg13g2_decap_8 FILLER_59_1204 ();
 sg13g2_decap_8 FILLER_59_1211 ();
 sg13g2_decap_8 FILLER_59_1218 ();
 sg13g2_decap_8 FILLER_59_1225 ();
 sg13g2_decap_8 FILLER_59_1232 ();
 sg13g2_decap_8 FILLER_59_1239 ();
 sg13g2_decap_8 FILLER_59_1246 ();
 sg13g2_decap_8 FILLER_59_1253 ();
 sg13g2_decap_8 FILLER_59_1260 ();
 sg13g2_decap_8 FILLER_59_1267 ();
 sg13g2_decap_8 FILLER_59_1274 ();
 sg13g2_decap_8 FILLER_59_1281 ();
 sg13g2_decap_8 FILLER_59_1288 ();
 sg13g2_decap_8 FILLER_59_1295 ();
 sg13g2_decap_8 FILLER_59_1302 ();
 sg13g2_decap_8 FILLER_59_1309 ();
 sg13g2_decap_8 FILLER_59_1316 ();
 sg13g2_decap_8 FILLER_59_1323 ();
 sg13g2_decap_8 FILLER_59_1330 ();
 sg13g2_decap_8 FILLER_59_1337 ();
 sg13g2_decap_8 FILLER_59_1344 ();
 sg13g2_decap_8 FILLER_59_1351 ();
 sg13g2_decap_8 FILLER_59_1358 ();
 sg13g2_decap_8 FILLER_59_1365 ();
 sg13g2_decap_8 FILLER_59_1372 ();
 sg13g2_decap_8 FILLER_59_1379 ();
 sg13g2_decap_8 FILLER_59_1386 ();
 sg13g2_decap_8 FILLER_59_1393 ();
 sg13g2_decap_8 FILLER_59_1400 ();
 sg13g2_decap_8 FILLER_59_1407 ();
 sg13g2_decap_8 FILLER_59_1414 ();
 sg13g2_decap_8 FILLER_59_1421 ();
 sg13g2_decap_8 FILLER_59_1428 ();
 sg13g2_decap_8 FILLER_59_1435 ();
 sg13g2_decap_8 FILLER_59_1442 ();
 sg13g2_decap_8 FILLER_59_1449 ();
 sg13g2_decap_8 FILLER_59_1456 ();
 sg13g2_decap_8 FILLER_59_1463 ();
 sg13g2_decap_8 FILLER_59_1470 ();
 sg13g2_decap_8 FILLER_59_1477 ();
 sg13g2_decap_8 FILLER_59_1484 ();
 sg13g2_decap_8 FILLER_59_1491 ();
 sg13g2_decap_8 FILLER_59_1498 ();
 sg13g2_decap_8 FILLER_59_1505 ();
 sg13g2_decap_8 FILLER_59_1512 ();
 sg13g2_decap_8 FILLER_59_1519 ();
 sg13g2_decap_8 FILLER_59_1526 ();
 sg13g2_decap_8 FILLER_59_1533 ();
 sg13g2_decap_8 FILLER_59_1540 ();
 sg13g2_decap_8 FILLER_59_1547 ();
 sg13g2_decap_8 FILLER_59_1554 ();
 sg13g2_decap_8 FILLER_59_1561 ();
 sg13g2_decap_8 FILLER_59_1568 ();
 sg13g2_decap_8 FILLER_59_1575 ();
 sg13g2_decap_8 FILLER_59_1582 ();
 sg13g2_decap_8 FILLER_59_1589 ();
 sg13g2_decap_8 FILLER_59_1596 ();
 sg13g2_decap_8 FILLER_59_1603 ();
 sg13g2_decap_8 FILLER_59_1610 ();
 sg13g2_decap_8 FILLER_59_1617 ();
 sg13g2_decap_8 FILLER_59_1624 ();
 sg13g2_decap_8 FILLER_59_1631 ();
 sg13g2_decap_8 FILLER_59_1638 ();
 sg13g2_decap_8 FILLER_59_1645 ();
 sg13g2_decap_8 FILLER_59_1652 ();
 sg13g2_decap_8 FILLER_59_1659 ();
 sg13g2_decap_8 FILLER_59_1666 ();
 sg13g2_decap_8 FILLER_59_1673 ();
 sg13g2_decap_8 FILLER_59_1680 ();
 sg13g2_decap_8 FILLER_59_1687 ();
 sg13g2_decap_8 FILLER_59_1694 ();
 sg13g2_decap_8 FILLER_59_1701 ();
 sg13g2_decap_8 FILLER_59_1708 ();
 sg13g2_decap_8 FILLER_59_1715 ();
 sg13g2_decap_8 FILLER_59_1722 ();
 sg13g2_decap_8 FILLER_59_1729 ();
 sg13g2_decap_8 FILLER_59_1736 ();
 sg13g2_decap_8 FILLER_59_1743 ();
 sg13g2_decap_8 FILLER_59_1750 ();
 sg13g2_decap_8 FILLER_59_1757 ();
 sg13g2_decap_4 FILLER_59_1764 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_decap_8 FILLER_60_7 ();
 sg13g2_decap_8 FILLER_60_14 ();
 sg13g2_decap_8 FILLER_60_21 ();
 sg13g2_decap_8 FILLER_60_28 ();
 sg13g2_decap_8 FILLER_60_35 ();
 sg13g2_decap_8 FILLER_60_42 ();
 sg13g2_decap_8 FILLER_60_49 ();
 sg13g2_decap_8 FILLER_60_56 ();
 sg13g2_decap_8 FILLER_60_63 ();
 sg13g2_decap_8 FILLER_60_70 ();
 sg13g2_fill_2 FILLER_60_77 ();
 sg13g2_decap_8 FILLER_60_82 ();
 sg13g2_fill_2 FILLER_60_89 ();
 sg13g2_fill_1 FILLER_60_91 ();
 sg13g2_fill_1 FILLER_60_97 ();
 sg13g2_fill_2 FILLER_60_134 ();
 sg13g2_fill_1 FILLER_60_170 ();
 sg13g2_decap_8 FILLER_60_254 ();
 sg13g2_fill_1 FILLER_60_274 ();
 sg13g2_fill_1 FILLER_60_284 ();
 sg13g2_fill_1 FILLER_60_299 ();
 sg13g2_fill_1 FILLER_60_310 ();
 sg13g2_fill_2 FILLER_60_363 ();
 sg13g2_fill_2 FILLER_60_376 ();
 sg13g2_fill_1 FILLER_60_449 ();
 sg13g2_decap_4 FILLER_60_482 ();
 sg13g2_fill_1 FILLER_60_486 ();
 sg13g2_fill_1 FILLER_60_523 ();
 sg13g2_decap_4 FILLER_60_536 ();
 sg13g2_fill_1 FILLER_60_568 ();
 sg13g2_decap_8 FILLER_60_630 ();
 sg13g2_fill_2 FILLER_60_637 ();
 sg13g2_fill_1 FILLER_60_639 ();
 sg13g2_decap_8 FILLER_60_657 ();
 sg13g2_decap_8 FILLER_60_664 ();
 sg13g2_fill_2 FILLER_60_697 ();
 sg13g2_decap_8 FILLER_60_709 ();
 sg13g2_decap_8 FILLER_60_716 ();
 sg13g2_decap_8 FILLER_60_759 ();
 sg13g2_fill_2 FILLER_60_766 ();
 sg13g2_fill_1 FILLER_60_768 ();
 sg13g2_decap_4 FILLER_60_792 ();
 sg13g2_decap_8 FILLER_60_800 ();
 sg13g2_decap_4 FILLER_60_807 ();
 sg13g2_fill_1 FILLER_60_811 ();
 sg13g2_decap_4 FILLER_60_815 ();
 sg13g2_fill_2 FILLER_60_819 ();
 sg13g2_fill_2 FILLER_60_830 ();
 sg13g2_fill_2 FILLER_60_841 ();
 sg13g2_decap_8 FILLER_60_848 ();
 sg13g2_decap_8 FILLER_60_855 ();
 sg13g2_fill_2 FILLER_60_862 ();
 sg13g2_fill_2 FILLER_60_872 ();
 sg13g2_decap_4 FILLER_60_918 ();
 sg13g2_fill_1 FILLER_60_922 ();
 sg13g2_fill_2 FILLER_60_928 ();
 sg13g2_fill_2 FILLER_60_940 ();
 sg13g2_fill_2 FILLER_60_960 ();
 sg13g2_fill_2 FILLER_60_967 ();
 sg13g2_fill_1 FILLER_60_1003 ();
 sg13g2_fill_1 FILLER_60_1012 ();
 sg13g2_decap_8 FILLER_60_1063 ();
 sg13g2_decap_8 FILLER_60_1070 ();
 sg13g2_decap_8 FILLER_60_1077 ();
 sg13g2_decap_8 FILLER_60_1084 ();
 sg13g2_decap_8 FILLER_60_1091 ();
 sg13g2_decap_8 FILLER_60_1098 ();
 sg13g2_decap_8 FILLER_60_1105 ();
 sg13g2_decap_8 FILLER_60_1112 ();
 sg13g2_decap_8 FILLER_60_1119 ();
 sg13g2_decap_8 FILLER_60_1126 ();
 sg13g2_decap_8 FILLER_60_1133 ();
 sg13g2_decap_8 FILLER_60_1140 ();
 sg13g2_decap_8 FILLER_60_1147 ();
 sg13g2_decap_8 FILLER_60_1154 ();
 sg13g2_decap_8 FILLER_60_1161 ();
 sg13g2_decap_8 FILLER_60_1168 ();
 sg13g2_decap_8 FILLER_60_1175 ();
 sg13g2_decap_8 FILLER_60_1182 ();
 sg13g2_decap_8 FILLER_60_1189 ();
 sg13g2_decap_8 FILLER_60_1196 ();
 sg13g2_decap_8 FILLER_60_1203 ();
 sg13g2_decap_8 FILLER_60_1210 ();
 sg13g2_decap_8 FILLER_60_1217 ();
 sg13g2_decap_8 FILLER_60_1224 ();
 sg13g2_decap_8 FILLER_60_1231 ();
 sg13g2_decap_8 FILLER_60_1238 ();
 sg13g2_decap_8 FILLER_60_1245 ();
 sg13g2_decap_8 FILLER_60_1252 ();
 sg13g2_decap_8 FILLER_60_1259 ();
 sg13g2_decap_8 FILLER_60_1266 ();
 sg13g2_decap_8 FILLER_60_1273 ();
 sg13g2_decap_8 FILLER_60_1280 ();
 sg13g2_decap_8 FILLER_60_1287 ();
 sg13g2_decap_8 FILLER_60_1294 ();
 sg13g2_decap_8 FILLER_60_1301 ();
 sg13g2_decap_8 FILLER_60_1308 ();
 sg13g2_decap_8 FILLER_60_1315 ();
 sg13g2_decap_8 FILLER_60_1322 ();
 sg13g2_decap_8 FILLER_60_1329 ();
 sg13g2_decap_8 FILLER_60_1336 ();
 sg13g2_decap_8 FILLER_60_1343 ();
 sg13g2_decap_8 FILLER_60_1350 ();
 sg13g2_decap_8 FILLER_60_1357 ();
 sg13g2_decap_8 FILLER_60_1364 ();
 sg13g2_decap_8 FILLER_60_1371 ();
 sg13g2_decap_8 FILLER_60_1378 ();
 sg13g2_decap_8 FILLER_60_1385 ();
 sg13g2_decap_8 FILLER_60_1392 ();
 sg13g2_decap_8 FILLER_60_1399 ();
 sg13g2_decap_8 FILLER_60_1406 ();
 sg13g2_decap_8 FILLER_60_1413 ();
 sg13g2_decap_8 FILLER_60_1420 ();
 sg13g2_decap_8 FILLER_60_1427 ();
 sg13g2_decap_8 FILLER_60_1434 ();
 sg13g2_decap_8 FILLER_60_1441 ();
 sg13g2_decap_8 FILLER_60_1448 ();
 sg13g2_decap_8 FILLER_60_1455 ();
 sg13g2_decap_8 FILLER_60_1462 ();
 sg13g2_decap_8 FILLER_60_1469 ();
 sg13g2_decap_8 FILLER_60_1476 ();
 sg13g2_decap_8 FILLER_60_1483 ();
 sg13g2_decap_8 FILLER_60_1490 ();
 sg13g2_decap_8 FILLER_60_1497 ();
 sg13g2_decap_8 FILLER_60_1504 ();
 sg13g2_decap_8 FILLER_60_1511 ();
 sg13g2_decap_8 FILLER_60_1518 ();
 sg13g2_decap_8 FILLER_60_1525 ();
 sg13g2_decap_8 FILLER_60_1532 ();
 sg13g2_decap_8 FILLER_60_1539 ();
 sg13g2_decap_8 FILLER_60_1546 ();
 sg13g2_decap_8 FILLER_60_1553 ();
 sg13g2_decap_8 FILLER_60_1560 ();
 sg13g2_decap_8 FILLER_60_1567 ();
 sg13g2_decap_8 FILLER_60_1574 ();
 sg13g2_decap_8 FILLER_60_1581 ();
 sg13g2_decap_8 FILLER_60_1588 ();
 sg13g2_decap_8 FILLER_60_1595 ();
 sg13g2_decap_8 FILLER_60_1602 ();
 sg13g2_decap_8 FILLER_60_1609 ();
 sg13g2_decap_8 FILLER_60_1616 ();
 sg13g2_decap_8 FILLER_60_1623 ();
 sg13g2_decap_8 FILLER_60_1630 ();
 sg13g2_decap_8 FILLER_60_1637 ();
 sg13g2_decap_8 FILLER_60_1644 ();
 sg13g2_decap_8 FILLER_60_1651 ();
 sg13g2_decap_8 FILLER_60_1658 ();
 sg13g2_decap_8 FILLER_60_1665 ();
 sg13g2_decap_8 FILLER_60_1672 ();
 sg13g2_decap_8 FILLER_60_1679 ();
 sg13g2_decap_8 FILLER_60_1686 ();
 sg13g2_decap_8 FILLER_60_1693 ();
 sg13g2_decap_8 FILLER_60_1700 ();
 sg13g2_decap_8 FILLER_60_1707 ();
 sg13g2_decap_8 FILLER_60_1714 ();
 sg13g2_decap_8 FILLER_60_1721 ();
 sg13g2_decap_8 FILLER_60_1728 ();
 sg13g2_decap_8 FILLER_60_1735 ();
 sg13g2_decap_8 FILLER_60_1742 ();
 sg13g2_decap_8 FILLER_60_1749 ();
 sg13g2_decap_8 FILLER_60_1756 ();
 sg13g2_decap_4 FILLER_60_1763 ();
 sg13g2_fill_1 FILLER_60_1767 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_decap_8 FILLER_61_7 ();
 sg13g2_decap_8 FILLER_61_14 ();
 sg13g2_decap_8 FILLER_61_21 ();
 sg13g2_decap_8 FILLER_61_28 ();
 sg13g2_decap_8 FILLER_61_35 ();
 sg13g2_decap_8 FILLER_61_42 ();
 sg13g2_decap_8 FILLER_61_49 ();
 sg13g2_decap_8 FILLER_61_56 ();
 sg13g2_decap_8 FILLER_61_63 ();
 sg13g2_decap_8 FILLER_61_70 ();
 sg13g2_decap_8 FILLER_61_77 ();
 sg13g2_decap_8 FILLER_61_84 ();
 sg13g2_decap_8 FILLER_61_91 ();
 sg13g2_decap_8 FILLER_61_98 ();
 sg13g2_decap_8 FILLER_61_105 ();
 sg13g2_fill_1 FILLER_61_112 ();
 sg13g2_fill_2 FILLER_61_116 ();
 sg13g2_fill_2 FILLER_61_126 ();
 sg13g2_decap_8 FILLER_61_139 ();
 sg13g2_fill_2 FILLER_61_146 ();
 sg13g2_fill_1 FILLER_61_148 ();
 sg13g2_decap_4 FILLER_61_152 ();
 sg13g2_fill_1 FILLER_61_156 ();
 sg13g2_fill_1 FILLER_61_179 ();
 sg13g2_fill_1 FILLER_61_189 ();
 sg13g2_fill_2 FILLER_61_206 ();
 sg13g2_decap_4 FILLER_61_245 ();
 sg13g2_decap_8 FILLER_61_254 ();
 sg13g2_fill_2 FILLER_61_261 ();
 sg13g2_fill_2 FILLER_61_295 ();
 sg13g2_fill_1 FILLER_61_305 ();
 sg13g2_fill_2 FILLER_61_324 ();
 sg13g2_fill_1 FILLER_61_326 ();
 sg13g2_decap_8 FILLER_61_434 ();
 sg13g2_decap_8 FILLER_61_441 ();
 sg13g2_fill_2 FILLER_61_448 ();
 sg13g2_decap_8 FILLER_61_462 ();
 sg13g2_fill_2 FILLER_61_484 ();
 sg13g2_fill_1 FILLER_61_486 ();
 sg13g2_decap_8 FILLER_61_500 ();
 sg13g2_fill_1 FILLER_61_507 ();
 sg13g2_decap_4 FILLER_61_524 ();
 sg13g2_decap_8 FILLER_61_533 ();
 sg13g2_decap_8 FILLER_61_540 ();
 sg13g2_decap_4 FILLER_61_547 ();
 sg13g2_fill_1 FILLER_61_570 ();
 sg13g2_fill_2 FILLER_61_590 ();
 sg13g2_decap_4 FILLER_61_602 ();
 sg13g2_fill_2 FILLER_61_606 ();
 sg13g2_fill_2 FILLER_61_643 ();
 sg13g2_fill_1 FILLER_61_645 ();
 sg13g2_decap_8 FILLER_61_651 ();
 sg13g2_fill_2 FILLER_61_658 ();
 sg13g2_fill_1 FILLER_61_660 ();
 sg13g2_decap_8 FILLER_61_679 ();
 sg13g2_decap_8 FILLER_61_686 ();
 sg13g2_decap_4 FILLER_61_693 ();
 sg13g2_fill_1 FILLER_61_697 ();
 sg13g2_decap_4 FILLER_61_729 ();
 sg13g2_fill_2 FILLER_61_736 ();
 sg13g2_fill_1 FILLER_61_738 ();
 sg13g2_decap_4 FILLER_61_773 ();
 sg13g2_fill_1 FILLER_61_777 ();
 sg13g2_fill_2 FILLER_61_786 ();
 sg13g2_fill_1 FILLER_61_826 ();
 sg13g2_fill_2 FILLER_61_889 ();
 sg13g2_fill_1 FILLER_61_891 ();
 sg13g2_fill_2 FILLER_61_1033 ();
 sg13g2_fill_1 FILLER_61_1035 ();
 sg13g2_decap_8 FILLER_61_1074 ();
 sg13g2_decap_8 FILLER_61_1081 ();
 sg13g2_decap_8 FILLER_61_1088 ();
 sg13g2_decap_8 FILLER_61_1095 ();
 sg13g2_decap_8 FILLER_61_1102 ();
 sg13g2_decap_8 FILLER_61_1109 ();
 sg13g2_decap_8 FILLER_61_1116 ();
 sg13g2_decap_8 FILLER_61_1123 ();
 sg13g2_decap_8 FILLER_61_1130 ();
 sg13g2_decap_8 FILLER_61_1137 ();
 sg13g2_decap_8 FILLER_61_1144 ();
 sg13g2_decap_8 FILLER_61_1151 ();
 sg13g2_decap_8 FILLER_61_1158 ();
 sg13g2_decap_8 FILLER_61_1165 ();
 sg13g2_decap_8 FILLER_61_1172 ();
 sg13g2_decap_8 FILLER_61_1179 ();
 sg13g2_decap_8 FILLER_61_1186 ();
 sg13g2_decap_8 FILLER_61_1193 ();
 sg13g2_decap_8 FILLER_61_1200 ();
 sg13g2_decap_8 FILLER_61_1207 ();
 sg13g2_decap_8 FILLER_61_1214 ();
 sg13g2_decap_8 FILLER_61_1221 ();
 sg13g2_decap_8 FILLER_61_1228 ();
 sg13g2_decap_8 FILLER_61_1235 ();
 sg13g2_decap_8 FILLER_61_1242 ();
 sg13g2_decap_8 FILLER_61_1249 ();
 sg13g2_decap_8 FILLER_61_1256 ();
 sg13g2_decap_8 FILLER_61_1263 ();
 sg13g2_decap_8 FILLER_61_1270 ();
 sg13g2_decap_8 FILLER_61_1277 ();
 sg13g2_decap_8 FILLER_61_1284 ();
 sg13g2_decap_8 FILLER_61_1291 ();
 sg13g2_decap_8 FILLER_61_1298 ();
 sg13g2_decap_8 FILLER_61_1305 ();
 sg13g2_decap_8 FILLER_61_1312 ();
 sg13g2_decap_8 FILLER_61_1319 ();
 sg13g2_decap_8 FILLER_61_1326 ();
 sg13g2_decap_8 FILLER_61_1333 ();
 sg13g2_decap_8 FILLER_61_1340 ();
 sg13g2_decap_8 FILLER_61_1347 ();
 sg13g2_decap_8 FILLER_61_1354 ();
 sg13g2_decap_8 FILLER_61_1361 ();
 sg13g2_decap_8 FILLER_61_1368 ();
 sg13g2_decap_8 FILLER_61_1375 ();
 sg13g2_decap_8 FILLER_61_1382 ();
 sg13g2_decap_8 FILLER_61_1389 ();
 sg13g2_decap_8 FILLER_61_1396 ();
 sg13g2_decap_8 FILLER_61_1403 ();
 sg13g2_decap_8 FILLER_61_1410 ();
 sg13g2_decap_8 FILLER_61_1417 ();
 sg13g2_decap_8 FILLER_61_1424 ();
 sg13g2_decap_8 FILLER_61_1431 ();
 sg13g2_decap_8 FILLER_61_1438 ();
 sg13g2_decap_8 FILLER_61_1445 ();
 sg13g2_decap_8 FILLER_61_1452 ();
 sg13g2_decap_8 FILLER_61_1459 ();
 sg13g2_decap_8 FILLER_61_1466 ();
 sg13g2_decap_8 FILLER_61_1473 ();
 sg13g2_decap_8 FILLER_61_1480 ();
 sg13g2_decap_8 FILLER_61_1487 ();
 sg13g2_decap_8 FILLER_61_1494 ();
 sg13g2_decap_8 FILLER_61_1501 ();
 sg13g2_decap_8 FILLER_61_1508 ();
 sg13g2_decap_8 FILLER_61_1515 ();
 sg13g2_decap_8 FILLER_61_1522 ();
 sg13g2_decap_8 FILLER_61_1529 ();
 sg13g2_decap_8 FILLER_61_1536 ();
 sg13g2_decap_8 FILLER_61_1543 ();
 sg13g2_decap_8 FILLER_61_1550 ();
 sg13g2_decap_8 FILLER_61_1557 ();
 sg13g2_decap_8 FILLER_61_1564 ();
 sg13g2_decap_8 FILLER_61_1571 ();
 sg13g2_decap_8 FILLER_61_1578 ();
 sg13g2_decap_8 FILLER_61_1585 ();
 sg13g2_decap_8 FILLER_61_1592 ();
 sg13g2_decap_8 FILLER_61_1599 ();
 sg13g2_decap_8 FILLER_61_1606 ();
 sg13g2_decap_8 FILLER_61_1613 ();
 sg13g2_decap_8 FILLER_61_1620 ();
 sg13g2_decap_8 FILLER_61_1627 ();
 sg13g2_decap_8 FILLER_61_1634 ();
 sg13g2_decap_8 FILLER_61_1641 ();
 sg13g2_decap_8 FILLER_61_1648 ();
 sg13g2_decap_8 FILLER_61_1655 ();
 sg13g2_decap_8 FILLER_61_1662 ();
 sg13g2_decap_8 FILLER_61_1669 ();
 sg13g2_decap_8 FILLER_61_1676 ();
 sg13g2_decap_8 FILLER_61_1683 ();
 sg13g2_decap_8 FILLER_61_1690 ();
 sg13g2_decap_8 FILLER_61_1697 ();
 sg13g2_decap_8 FILLER_61_1704 ();
 sg13g2_decap_8 FILLER_61_1711 ();
 sg13g2_decap_8 FILLER_61_1718 ();
 sg13g2_decap_8 FILLER_61_1725 ();
 sg13g2_decap_8 FILLER_61_1732 ();
 sg13g2_decap_8 FILLER_61_1739 ();
 sg13g2_decap_8 FILLER_61_1746 ();
 sg13g2_decap_8 FILLER_61_1753 ();
 sg13g2_decap_8 FILLER_61_1760 ();
 sg13g2_fill_1 FILLER_61_1767 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_decap_8 FILLER_62_7 ();
 sg13g2_decap_8 FILLER_62_14 ();
 sg13g2_decap_8 FILLER_62_21 ();
 sg13g2_decap_8 FILLER_62_28 ();
 sg13g2_decap_8 FILLER_62_35 ();
 sg13g2_decap_8 FILLER_62_42 ();
 sg13g2_decap_8 FILLER_62_49 ();
 sg13g2_decap_8 FILLER_62_56 ();
 sg13g2_decap_8 FILLER_62_63 ();
 sg13g2_decap_8 FILLER_62_70 ();
 sg13g2_decap_8 FILLER_62_77 ();
 sg13g2_decap_8 FILLER_62_84 ();
 sg13g2_decap_8 FILLER_62_91 ();
 sg13g2_decap_8 FILLER_62_98 ();
 sg13g2_decap_8 FILLER_62_105 ();
 sg13g2_decap_8 FILLER_62_112 ();
 sg13g2_decap_8 FILLER_62_119 ();
 sg13g2_fill_2 FILLER_62_126 ();
 sg13g2_fill_2 FILLER_62_249 ();
 sg13g2_fill_1 FILLER_62_251 ();
 sg13g2_fill_2 FILLER_62_268 ();
 sg13g2_fill_2 FILLER_62_361 ();
 sg13g2_fill_1 FILLER_62_363 ();
 sg13g2_fill_1 FILLER_62_376 ();
 sg13g2_fill_1 FILLER_62_414 ();
 sg13g2_fill_1 FILLER_62_440 ();
 sg13g2_decap_4 FILLER_62_457 ();
 sg13g2_decap_8 FILLER_62_466 ();
 sg13g2_fill_1 FILLER_62_473 ();
 sg13g2_fill_1 FILLER_62_480 ();
 sg13g2_decap_4 FILLER_62_492 ();
 sg13g2_fill_2 FILLER_62_496 ();
 sg13g2_decap_4 FILLER_62_503 ();
 sg13g2_fill_1 FILLER_62_507 ();
 sg13g2_fill_2 FILLER_62_516 ();
 sg13g2_fill_1 FILLER_62_518 ();
 sg13g2_decap_4 FILLER_62_531 ();
 sg13g2_fill_2 FILLER_62_540 ();
 sg13g2_fill_1 FILLER_62_542 ();
 sg13g2_decap_4 FILLER_62_548 ();
 sg13g2_fill_1 FILLER_62_552 ();
 sg13g2_decap_4 FILLER_62_624 ();
 sg13g2_fill_1 FILLER_62_628 ();
 sg13g2_decap_8 FILLER_62_669 ();
 sg13g2_decap_4 FILLER_62_676 ();
 sg13g2_fill_2 FILLER_62_680 ();
 sg13g2_fill_2 FILLER_62_699 ();
 sg13g2_fill_2 FILLER_62_710 ();
 sg13g2_fill_1 FILLER_62_712 ();
 sg13g2_decap_4 FILLER_62_726 ();
 sg13g2_fill_2 FILLER_62_730 ();
 sg13g2_fill_1 FILLER_62_738 ();
 sg13g2_fill_2 FILLER_62_744 ();
 sg13g2_fill_2 FILLER_62_755 ();
 sg13g2_fill_1 FILLER_62_757 ();
 sg13g2_fill_1 FILLER_62_812 ();
 sg13g2_fill_1 FILLER_62_827 ();
 sg13g2_decap_8 FILLER_62_846 ();
 sg13g2_decap_8 FILLER_62_916 ();
 sg13g2_decap_8 FILLER_62_923 ();
 sg13g2_fill_2 FILLER_62_930 ();
 sg13g2_decap_8 FILLER_62_937 ();
 sg13g2_decap_4 FILLER_62_944 ();
 sg13g2_fill_2 FILLER_62_948 ();
 sg13g2_decap_8 FILLER_62_958 ();
 sg13g2_fill_1 FILLER_62_965 ();
 sg13g2_fill_2 FILLER_62_985 ();
 sg13g2_fill_1 FILLER_62_1018 ();
 sg13g2_fill_2 FILLER_62_1038 ();
 sg13g2_fill_2 FILLER_62_1045 ();
 sg13g2_decap_8 FILLER_62_1090 ();
 sg13g2_decap_8 FILLER_62_1097 ();
 sg13g2_decap_8 FILLER_62_1104 ();
 sg13g2_decap_8 FILLER_62_1111 ();
 sg13g2_decap_8 FILLER_62_1118 ();
 sg13g2_decap_8 FILLER_62_1125 ();
 sg13g2_decap_8 FILLER_62_1132 ();
 sg13g2_decap_8 FILLER_62_1139 ();
 sg13g2_decap_8 FILLER_62_1146 ();
 sg13g2_decap_8 FILLER_62_1153 ();
 sg13g2_decap_8 FILLER_62_1160 ();
 sg13g2_decap_8 FILLER_62_1167 ();
 sg13g2_decap_8 FILLER_62_1174 ();
 sg13g2_decap_8 FILLER_62_1181 ();
 sg13g2_decap_8 FILLER_62_1188 ();
 sg13g2_decap_8 FILLER_62_1195 ();
 sg13g2_decap_8 FILLER_62_1202 ();
 sg13g2_decap_8 FILLER_62_1209 ();
 sg13g2_decap_8 FILLER_62_1216 ();
 sg13g2_decap_8 FILLER_62_1223 ();
 sg13g2_decap_8 FILLER_62_1230 ();
 sg13g2_decap_8 FILLER_62_1237 ();
 sg13g2_decap_8 FILLER_62_1244 ();
 sg13g2_decap_8 FILLER_62_1251 ();
 sg13g2_decap_8 FILLER_62_1258 ();
 sg13g2_decap_8 FILLER_62_1265 ();
 sg13g2_decap_8 FILLER_62_1272 ();
 sg13g2_decap_8 FILLER_62_1279 ();
 sg13g2_decap_8 FILLER_62_1286 ();
 sg13g2_decap_8 FILLER_62_1293 ();
 sg13g2_decap_8 FILLER_62_1300 ();
 sg13g2_decap_8 FILLER_62_1307 ();
 sg13g2_decap_8 FILLER_62_1314 ();
 sg13g2_decap_8 FILLER_62_1321 ();
 sg13g2_decap_8 FILLER_62_1328 ();
 sg13g2_decap_8 FILLER_62_1335 ();
 sg13g2_decap_8 FILLER_62_1342 ();
 sg13g2_decap_8 FILLER_62_1349 ();
 sg13g2_decap_8 FILLER_62_1356 ();
 sg13g2_decap_8 FILLER_62_1363 ();
 sg13g2_decap_8 FILLER_62_1370 ();
 sg13g2_decap_8 FILLER_62_1377 ();
 sg13g2_decap_8 FILLER_62_1384 ();
 sg13g2_decap_8 FILLER_62_1391 ();
 sg13g2_decap_8 FILLER_62_1398 ();
 sg13g2_decap_8 FILLER_62_1405 ();
 sg13g2_decap_8 FILLER_62_1412 ();
 sg13g2_decap_8 FILLER_62_1419 ();
 sg13g2_decap_8 FILLER_62_1426 ();
 sg13g2_decap_8 FILLER_62_1433 ();
 sg13g2_decap_8 FILLER_62_1440 ();
 sg13g2_decap_8 FILLER_62_1447 ();
 sg13g2_decap_8 FILLER_62_1454 ();
 sg13g2_decap_8 FILLER_62_1461 ();
 sg13g2_decap_8 FILLER_62_1468 ();
 sg13g2_decap_8 FILLER_62_1475 ();
 sg13g2_decap_8 FILLER_62_1482 ();
 sg13g2_decap_8 FILLER_62_1489 ();
 sg13g2_decap_8 FILLER_62_1496 ();
 sg13g2_decap_8 FILLER_62_1503 ();
 sg13g2_decap_8 FILLER_62_1510 ();
 sg13g2_decap_8 FILLER_62_1517 ();
 sg13g2_decap_8 FILLER_62_1524 ();
 sg13g2_decap_8 FILLER_62_1531 ();
 sg13g2_decap_8 FILLER_62_1538 ();
 sg13g2_decap_8 FILLER_62_1545 ();
 sg13g2_decap_8 FILLER_62_1552 ();
 sg13g2_decap_8 FILLER_62_1559 ();
 sg13g2_decap_8 FILLER_62_1566 ();
 sg13g2_decap_8 FILLER_62_1573 ();
 sg13g2_decap_8 FILLER_62_1580 ();
 sg13g2_decap_8 FILLER_62_1587 ();
 sg13g2_decap_8 FILLER_62_1594 ();
 sg13g2_decap_8 FILLER_62_1601 ();
 sg13g2_decap_8 FILLER_62_1608 ();
 sg13g2_decap_8 FILLER_62_1615 ();
 sg13g2_decap_8 FILLER_62_1622 ();
 sg13g2_decap_8 FILLER_62_1629 ();
 sg13g2_decap_8 FILLER_62_1636 ();
 sg13g2_decap_8 FILLER_62_1643 ();
 sg13g2_decap_8 FILLER_62_1650 ();
 sg13g2_decap_8 FILLER_62_1657 ();
 sg13g2_decap_8 FILLER_62_1664 ();
 sg13g2_decap_8 FILLER_62_1671 ();
 sg13g2_decap_8 FILLER_62_1678 ();
 sg13g2_decap_8 FILLER_62_1685 ();
 sg13g2_decap_8 FILLER_62_1692 ();
 sg13g2_decap_8 FILLER_62_1699 ();
 sg13g2_decap_8 FILLER_62_1706 ();
 sg13g2_decap_8 FILLER_62_1713 ();
 sg13g2_decap_8 FILLER_62_1720 ();
 sg13g2_decap_8 FILLER_62_1727 ();
 sg13g2_decap_8 FILLER_62_1734 ();
 sg13g2_decap_8 FILLER_62_1741 ();
 sg13g2_decap_8 FILLER_62_1748 ();
 sg13g2_decap_8 FILLER_62_1755 ();
 sg13g2_decap_4 FILLER_62_1762 ();
 sg13g2_fill_2 FILLER_62_1766 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_decap_8 FILLER_63_7 ();
 sg13g2_decap_8 FILLER_63_14 ();
 sg13g2_decap_8 FILLER_63_21 ();
 sg13g2_decap_8 FILLER_63_28 ();
 sg13g2_decap_8 FILLER_63_35 ();
 sg13g2_decap_8 FILLER_63_42 ();
 sg13g2_decap_8 FILLER_63_49 ();
 sg13g2_decap_8 FILLER_63_56 ();
 sg13g2_decap_8 FILLER_63_63 ();
 sg13g2_decap_8 FILLER_63_70 ();
 sg13g2_decap_8 FILLER_63_77 ();
 sg13g2_decap_8 FILLER_63_84 ();
 sg13g2_decap_4 FILLER_63_91 ();
 sg13g2_fill_2 FILLER_63_95 ();
 sg13g2_fill_2 FILLER_63_123 ();
 sg13g2_fill_1 FILLER_63_125 ();
 sg13g2_fill_1 FILLER_63_132 ();
 sg13g2_decap_4 FILLER_63_136 ();
 sg13g2_decap_8 FILLER_63_144 ();
 sg13g2_decap_4 FILLER_63_151 ();
 sg13g2_fill_1 FILLER_63_155 ();
 sg13g2_decap_8 FILLER_63_173 ();
 sg13g2_decap_8 FILLER_63_180 ();
 sg13g2_fill_1 FILLER_63_187 ();
 sg13g2_decap_8 FILLER_63_203 ();
 sg13g2_decap_4 FILLER_63_210 ();
 sg13g2_fill_1 FILLER_63_214 ();
 sg13g2_fill_2 FILLER_63_247 ();
 sg13g2_fill_1 FILLER_63_249 ();
 sg13g2_fill_2 FILLER_63_338 ();
 sg13g2_fill_1 FILLER_63_376 ();
 sg13g2_fill_2 FILLER_63_382 ();
 sg13g2_fill_1 FILLER_63_389 ();
 sg13g2_decap_4 FILLER_63_402 ();
 sg13g2_fill_2 FILLER_63_406 ();
 sg13g2_fill_2 FILLER_63_418 ();
 sg13g2_fill_2 FILLER_63_425 ();
 sg13g2_decap_8 FILLER_63_443 ();
 sg13g2_fill_2 FILLER_63_450 ();
 sg13g2_fill_2 FILLER_63_473 ();
 sg13g2_fill_1 FILLER_63_475 ();
 sg13g2_fill_2 FILLER_63_481 ();
 sg13g2_fill_1 FILLER_63_483 ();
 sg13g2_fill_2 FILLER_63_512 ();
 sg13g2_fill_1 FILLER_63_514 ();
 sg13g2_fill_2 FILLER_63_527 ();
 sg13g2_fill_1 FILLER_63_529 ();
 sg13g2_fill_1 FILLER_63_549 ();
 sg13g2_decap_8 FILLER_63_555 ();
 sg13g2_decap_8 FILLER_63_562 ();
 sg13g2_decap_8 FILLER_63_569 ();
 sg13g2_decap_8 FILLER_63_576 ();
 sg13g2_fill_2 FILLER_63_583 ();
 sg13g2_decap_8 FILLER_63_593 ();
 sg13g2_fill_1 FILLER_63_600 ();
 sg13g2_decap_8 FILLER_63_617 ();
 sg13g2_fill_2 FILLER_63_624 ();
 sg13g2_decap_8 FILLER_63_631 ();
 sg13g2_decap_4 FILLER_63_638 ();
 sg13g2_fill_2 FILLER_63_642 ();
 sg13g2_fill_2 FILLER_63_649 ();
 sg13g2_fill_1 FILLER_63_651 ();
 sg13g2_decap_4 FILLER_63_657 ();
 sg13g2_fill_1 FILLER_63_661 ();
 sg13g2_decap_8 FILLER_63_667 ();
 sg13g2_fill_2 FILLER_63_674 ();
 sg13g2_fill_1 FILLER_63_686 ();
 sg13g2_decap_4 FILLER_63_699 ();
 sg13g2_fill_2 FILLER_63_703 ();
 sg13g2_fill_2 FILLER_63_741 ();
 sg13g2_fill_1 FILLER_63_750 ();
 sg13g2_fill_1 FILLER_63_767 ();
 sg13g2_fill_2 FILLER_63_777 ();
 sg13g2_fill_1 FILLER_63_779 ();
 sg13g2_decap_8 FILLER_63_805 ();
 sg13g2_fill_2 FILLER_63_817 ();
 sg13g2_decap_4 FILLER_63_837 ();
 sg13g2_fill_1 FILLER_63_885 ();
 sg13g2_fill_2 FILLER_63_899 ();
 sg13g2_fill_2 FILLER_63_910 ();
 sg13g2_fill_2 FILLER_63_929 ();
 sg13g2_decap_8 FILLER_63_944 ();
 sg13g2_decap_8 FILLER_63_951 ();
 sg13g2_decap_4 FILLER_63_958 ();
 sg13g2_fill_1 FILLER_63_962 ();
 sg13g2_fill_2 FILLER_63_993 ();
 sg13g2_fill_2 FILLER_63_1011 ();
 sg13g2_fill_2 FILLER_63_1055 ();
 sg13g2_decap_8 FILLER_63_1077 ();
 sg13g2_decap_8 FILLER_63_1084 ();
 sg13g2_decap_8 FILLER_63_1091 ();
 sg13g2_decap_8 FILLER_63_1098 ();
 sg13g2_decap_8 FILLER_63_1105 ();
 sg13g2_decap_8 FILLER_63_1112 ();
 sg13g2_decap_8 FILLER_63_1119 ();
 sg13g2_decap_8 FILLER_63_1126 ();
 sg13g2_decap_8 FILLER_63_1133 ();
 sg13g2_decap_8 FILLER_63_1140 ();
 sg13g2_decap_8 FILLER_63_1147 ();
 sg13g2_decap_8 FILLER_63_1154 ();
 sg13g2_decap_8 FILLER_63_1161 ();
 sg13g2_decap_8 FILLER_63_1168 ();
 sg13g2_decap_8 FILLER_63_1175 ();
 sg13g2_decap_8 FILLER_63_1182 ();
 sg13g2_decap_8 FILLER_63_1189 ();
 sg13g2_decap_8 FILLER_63_1196 ();
 sg13g2_decap_8 FILLER_63_1203 ();
 sg13g2_decap_8 FILLER_63_1210 ();
 sg13g2_decap_8 FILLER_63_1217 ();
 sg13g2_decap_8 FILLER_63_1224 ();
 sg13g2_decap_8 FILLER_63_1231 ();
 sg13g2_decap_8 FILLER_63_1238 ();
 sg13g2_decap_8 FILLER_63_1245 ();
 sg13g2_decap_8 FILLER_63_1252 ();
 sg13g2_decap_8 FILLER_63_1259 ();
 sg13g2_decap_8 FILLER_63_1266 ();
 sg13g2_decap_8 FILLER_63_1273 ();
 sg13g2_decap_8 FILLER_63_1280 ();
 sg13g2_decap_8 FILLER_63_1287 ();
 sg13g2_decap_8 FILLER_63_1294 ();
 sg13g2_decap_8 FILLER_63_1301 ();
 sg13g2_decap_8 FILLER_63_1308 ();
 sg13g2_decap_8 FILLER_63_1315 ();
 sg13g2_decap_8 FILLER_63_1322 ();
 sg13g2_decap_8 FILLER_63_1329 ();
 sg13g2_decap_8 FILLER_63_1336 ();
 sg13g2_decap_8 FILLER_63_1343 ();
 sg13g2_decap_8 FILLER_63_1350 ();
 sg13g2_decap_8 FILLER_63_1357 ();
 sg13g2_decap_8 FILLER_63_1364 ();
 sg13g2_decap_8 FILLER_63_1371 ();
 sg13g2_decap_8 FILLER_63_1378 ();
 sg13g2_decap_8 FILLER_63_1385 ();
 sg13g2_decap_8 FILLER_63_1392 ();
 sg13g2_decap_8 FILLER_63_1399 ();
 sg13g2_decap_8 FILLER_63_1406 ();
 sg13g2_decap_8 FILLER_63_1413 ();
 sg13g2_decap_8 FILLER_63_1420 ();
 sg13g2_decap_8 FILLER_63_1427 ();
 sg13g2_decap_8 FILLER_63_1434 ();
 sg13g2_decap_8 FILLER_63_1441 ();
 sg13g2_decap_8 FILLER_63_1448 ();
 sg13g2_decap_8 FILLER_63_1455 ();
 sg13g2_decap_8 FILLER_63_1462 ();
 sg13g2_decap_8 FILLER_63_1469 ();
 sg13g2_decap_8 FILLER_63_1476 ();
 sg13g2_decap_8 FILLER_63_1483 ();
 sg13g2_decap_8 FILLER_63_1490 ();
 sg13g2_decap_8 FILLER_63_1497 ();
 sg13g2_decap_8 FILLER_63_1504 ();
 sg13g2_decap_8 FILLER_63_1511 ();
 sg13g2_decap_8 FILLER_63_1518 ();
 sg13g2_decap_8 FILLER_63_1525 ();
 sg13g2_decap_8 FILLER_63_1532 ();
 sg13g2_decap_8 FILLER_63_1539 ();
 sg13g2_decap_8 FILLER_63_1546 ();
 sg13g2_decap_8 FILLER_63_1553 ();
 sg13g2_decap_8 FILLER_63_1560 ();
 sg13g2_decap_8 FILLER_63_1567 ();
 sg13g2_decap_8 FILLER_63_1574 ();
 sg13g2_decap_8 FILLER_63_1581 ();
 sg13g2_decap_8 FILLER_63_1588 ();
 sg13g2_decap_8 FILLER_63_1595 ();
 sg13g2_decap_8 FILLER_63_1602 ();
 sg13g2_decap_8 FILLER_63_1609 ();
 sg13g2_decap_8 FILLER_63_1616 ();
 sg13g2_decap_8 FILLER_63_1623 ();
 sg13g2_decap_8 FILLER_63_1630 ();
 sg13g2_decap_8 FILLER_63_1637 ();
 sg13g2_decap_8 FILLER_63_1644 ();
 sg13g2_decap_8 FILLER_63_1651 ();
 sg13g2_decap_8 FILLER_63_1658 ();
 sg13g2_decap_8 FILLER_63_1665 ();
 sg13g2_decap_8 FILLER_63_1672 ();
 sg13g2_decap_8 FILLER_63_1679 ();
 sg13g2_decap_8 FILLER_63_1686 ();
 sg13g2_decap_8 FILLER_63_1693 ();
 sg13g2_decap_8 FILLER_63_1700 ();
 sg13g2_decap_8 FILLER_63_1707 ();
 sg13g2_decap_8 FILLER_63_1714 ();
 sg13g2_decap_8 FILLER_63_1721 ();
 sg13g2_decap_8 FILLER_63_1728 ();
 sg13g2_decap_8 FILLER_63_1735 ();
 sg13g2_decap_8 FILLER_63_1742 ();
 sg13g2_decap_8 FILLER_63_1749 ();
 sg13g2_decap_8 FILLER_63_1756 ();
 sg13g2_decap_4 FILLER_63_1763 ();
 sg13g2_fill_1 FILLER_63_1767 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_8 FILLER_64_7 ();
 sg13g2_decap_8 FILLER_64_14 ();
 sg13g2_decap_8 FILLER_64_21 ();
 sg13g2_decap_8 FILLER_64_28 ();
 sg13g2_decap_8 FILLER_64_35 ();
 sg13g2_decap_8 FILLER_64_42 ();
 sg13g2_decap_8 FILLER_64_49 ();
 sg13g2_decap_8 FILLER_64_56 ();
 sg13g2_decap_8 FILLER_64_63 ();
 sg13g2_decap_8 FILLER_64_70 ();
 sg13g2_decap_8 FILLER_64_77 ();
 sg13g2_decap_8 FILLER_64_84 ();
 sg13g2_decap_8 FILLER_64_91 ();
 sg13g2_decap_8 FILLER_64_98 ();
 sg13g2_decap_8 FILLER_64_105 ();
 sg13g2_fill_2 FILLER_64_164 ();
 sg13g2_fill_2 FILLER_64_170 ();
 sg13g2_decap_8 FILLER_64_198 ();
 sg13g2_decap_8 FILLER_64_213 ();
 sg13g2_fill_1 FILLER_64_223 ();
 sg13g2_fill_2 FILLER_64_250 ();
 sg13g2_fill_1 FILLER_64_312 ();
 sg13g2_fill_2 FILLER_64_326 ();
 sg13g2_fill_1 FILLER_64_346 ();
 sg13g2_fill_2 FILLER_64_373 ();
 sg13g2_fill_1 FILLER_64_399 ();
 sg13g2_fill_2 FILLER_64_419 ();
 sg13g2_fill_1 FILLER_64_448 ();
 sg13g2_fill_2 FILLER_64_461 ();
 sg13g2_decap_8 FILLER_64_468 ();
 sg13g2_decap_8 FILLER_64_475 ();
 sg13g2_fill_2 FILLER_64_495 ();
 sg13g2_decap_4 FILLER_64_502 ();
 sg13g2_fill_2 FILLER_64_506 ();
 sg13g2_fill_2 FILLER_64_513 ();
 sg13g2_decap_8 FILLER_64_524 ();
 sg13g2_fill_2 FILLER_64_531 ();
 sg13g2_fill_1 FILLER_64_537 ();
 sg13g2_fill_2 FILLER_64_548 ();
 sg13g2_fill_1 FILLER_64_550 ();
 sg13g2_decap_8 FILLER_64_560 ();
 sg13g2_decap_8 FILLER_64_567 ();
 sg13g2_decap_8 FILLER_64_574 ();
 sg13g2_decap_8 FILLER_64_581 ();
 sg13g2_decap_8 FILLER_64_588 ();
 sg13g2_decap_8 FILLER_64_595 ();
 sg13g2_decap_8 FILLER_64_602 ();
 sg13g2_decap_8 FILLER_64_609 ();
 sg13g2_fill_1 FILLER_64_616 ();
 sg13g2_decap_8 FILLER_64_628 ();
 sg13g2_decap_8 FILLER_64_635 ();
 sg13g2_fill_2 FILLER_64_647 ();
 sg13g2_fill_1 FILLER_64_649 ();
 sg13g2_fill_2 FILLER_64_655 ();
 sg13g2_fill_1 FILLER_64_657 ();
 sg13g2_decap_8 FILLER_64_667 ();
 sg13g2_fill_1 FILLER_64_674 ();
 sg13g2_fill_1 FILLER_64_690 ();
 sg13g2_decap_4 FILLER_64_709 ();
 sg13g2_fill_2 FILLER_64_726 ();
 sg13g2_fill_1 FILLER_64_728 ();
 sg13g2_fill_2 FILLER_64_790 ();
 sg13g2_fill_2 FILLER_64_805 ();
 sg13g2_fill_2 FILLER_64_820 ();
 sg13g2_decap_8 FILLER_64_847 ();
 sg13g2_decap_4 FILLER_64_854 ();
 sg13g2_fill_1 FILLER_64_863 ();
 sg13g2_fill_2 FILLER_64_877 ();
 sg13g2_fill_2 FILLER_64_889 ();
 sg13g2_fill_1 FILLER_64_891 ();
 sg13g2_decap_8 FILLER_64_915 ();
 sg13g2_fill_1 FILLER_64_922 ();
 sg13g2_decap_4 FILLER_64_975 ();
 sg13g2_fill_1 FILLER_64_979 ();
 sg13g2_fill_1 FILLER_64_1001 ();
 sg13g2_fill_2 FILLER_64_1031 ();
 sg13g2_fill_2 FILLER_64_1064 ();
 sg13g2_decap_8 FILLER_64_1101 ();
 sg13g2_decap_8 FILLER_64_1108 ();
 sg13g2_decap_8 FILLER_64_1115 ();
 sg13g2_decap_8 FILLER_64_1122 ();
 sg13g2_decap_8 FILLER_64_1129 ();
 sg13g2_decap_8 FILLER_64_1136 ();
 sg13g2_decap_8 FILLER_64_1143 ();
 sg13g2_decap_8 FILLER_64_1150 ();
 sg13g2_decap_8 FILLER_64_1157 ();
 sg13g2_decap_8 FILLER_64_1164 ();
 sg13g2_decap_8 FILLER_64_1171 ();
 sg13g2_decap_8 FILLER_64_1178 ();
 sg13g2_decap_8 FILLER_64_1185 ();
 sg13g2_decap_8 FILLER_64_1192 ();
 sg13g2_decap_8 FILLER_64_1199 ();
 sg13g2_decap_8 FILLER_64_1206 ();
 sg13g2_decap_8 FILLER_64_1213 ();
 sg13g2_decap_8 FILLER_64_1220 ();
 sg13g2_decap_8 FILLER_64_1227 ();
 sg13g2_decap_8 FILLER_64_1234 ();
 sg13g2_decap_8 FILLER_64_1241 ();
 sg13g2_decap_8 FILLER_64_1248 ();
 sg13g2_decap_8 FILLER_64_1255 ();
 sg13g2_decap_8 FILLER_64_1262 ();
 sg13g2_decap_8 FILLER_64_1269 ();
 sg13g2_decap_8 FILLER_64_1276 ();
 sg13g2_decap_8 FILLER_64_1283 ();
 sg13g2_decap_8 FILLER_64_1290 ();
 sg13g2_decap_8 FILLER_64_1297 ();
 sg13g2_decap_8 FILLER_64_1304 ();
 sg13g2_decap_8 FILLER_64_1311 ();
 sg13g2_decap_8 FILLER_64_1318 ();
 sg13g2_decap_8 FILLER_64_1325 ();
 sg13g2_decap_8 FILLER_64_1332 ();
 sg13g2_decap_8 FILLER_64_1339 ();
 sg13g2_decap_8 FILLER_64_1346 ();
 sg13g2_decap_8 FILLER_64_1353 ();
 sg13g2_decap_8 FILLER_64_1360 ();
 sg13g2_decap_8 FILLER_64_1367 ();
 sg13g2_decap_8 FILLER_64_1374 ();
 sg13g2_decap_8 FILLER_64_1381 ();
 sg13g2_decap_8 FILLER_64_1388 ();
 sg13g2_decap_8 FILLER_64_1395 ();
 sg13g2_decap_8 FILLER_64_1402 ();
 sg13g2_decap_8 FILLER_64_1409 ();
 sg13g2_decap_8 FILLER_64_1416 ();
 sg13g2_decap_8 FILLER_64_1423 ();
 sg13g2_decap_8 FILLER_64_1430 ();
 sg13g2_decap_8 FILLER_64_1437 ();
 sg13g2_decap_8 FILLER_64_1444 ();
 sg13g2_decap_8 FILLER_64_1451 ();
 sg13g2_decap_8 FILLER_64_1458 ();
 sg13g2_decap_8 FILLER_64_1465 ();
 sg13g2_decap_8 FILLER_64_1472 ();
 sg13g2_decap_8 FILLER_64_1479 ();
 sg13g2_decap_8 FILLER_64_1486 ();
 sg13g2_decap_8 FILLER_64_1493 ();
 sg13g2_decap_8 FILLER_64_1500 ();
 sg13g2_decap_8 FILLER_64_1507 ();
 sg13g2_decap_8 FILLER_64_1514 ();
 sg13g2_decap_8 FILLER_64_1521 ();
 sg13g2_decap_8 FILLER_64_1528 ();
 sg13g2_decap_8 FILLER_64_1535 ();
 sg13g2_decap_8 FILLER_64_1542 ();
 sg13g2_decap_8 FILLER_64_1549 ();
 sg13g2_decap_8 FILLER_64_1556 ();
 sg13g2_decap_8 FILLER_64_1563 ();
 sg13g2_decap_8 FILLER_64_1570 ();
 sg13g2_decap_8 FILLER_64_1577 ();
 sg13g2_decap_8 FILLER_64_1584 ();
 sg13g2_decap_8 FILLER_64_1591 ();
 sg13g2_decap_8 FILLER_64_1598 ();
 sg13g2_decap_8 FILLER_64_1605 ();
 sg13g2_decap_8 FILLER_64_1612 ();
 sg13g2_decap_8 FILLER_64_1619 ();
 sg13g2_decap_8 FILLER_64_1626 ();
 sg13g2_decap_8 FILLER_64_1633 ();
 sg13g2_decap_8 FILLER_64_1640 ();
 sg13g2_decap_8 FILLER_64_1647 ();
 sg13g2_decap_8 FILLER_64_1654 ();
 sg13g2_decap_8 FILLER_64_1661 ();
 sg13g2_decap_8 FILLER_64_1668 ();
 sg13g2_decap_8 FILLER_64_1675 ();
 sg13g2_decap_8 FILLER_64_1682 ();
 sg13g2_decap_8 FILLER_64_1689 ();
 sg13g2_decap_8 FILLER_64_1696 ();
 sg13g2_decap_8 FILLER_64_1703 ();
 sg13g2_decap_8 FILLER_64_1710 ();
 sg13g2_decap_8 FILLER_64_1717 ();
 sg13g2_decap_8 FILLER_64_1724 ();
 sg13g2_decap_8 FILLER_64_1731 ();
 sg13g2_decap_8 FILLER_64_1738 ();
 sg13g2_decap_8 FILLER_64_1745 ();
 sg13g2_decap_8 FILLER_64_1752 ();
 sg13g2_decap_8 FILLER_64_1759 ();
 sg13g2_fill_2 FILLER_64_1766 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_8 FILLER_65_7 ();
 sg13g2_decap_8 FILLER_65_14 ();
 sg13g2_decap_8 FILLER_65_21 ();
 sg13g2_decap_8 FILLER_65_28 ();
 sg13g2_decap_8 FILLER_65_35 ();
 sg13g2_decap_8 FILLER_65_42 ();
 sg13g2_decap_8 FILLER_65_49 ();
 sg13g2_decap_8 FILLER_65_56 ();
 sg13g2_fill_2 FILLER_65_63 ();
 sg13g2_fill_2 FILLER_65_94 ();
 sg13g2_fill_1 FILLER_65_96 ();
 sg13g2_decap_8 FILLER_65_106 ();
 sg13g2_fill_2 FILLER_65_113 ();
 sg13g2_fill_1 FILLER_65_120 ();
 sg13g2_fill_2 FILLER_65_138 ();
 sg13g2_fill_1 FILLER_65_140 ();
 sg13g2_fill_2 FILLER_65_151 ();
 sg13g2_decap_4 FILLER_65_180 ();
 sg13g2_fill_1 FILLER_65_184 ();
 sg13g2_decap_4 FILLER_65_236 ();
 sg13g2_fill_1 FILLER_65_240 ();
 sg13g2_decap_8 FILLER_65_259 ();
 sg13g2_decap_8 FILLER_65_266 ();
 sg13g2_fill_1 FILLER_65_273 ();
 sg13g2_fill_1 FILLER_65_277 ();
 sg13g2_fill_2 FILLER_65_283 ();
 sg13g2_fill_1 FILLER_65_317 ();
 sg13g2_fill_2 FILLER_65_332 ();
 sg13g2_decap_4 FILLER_65_343 ();
 sg13g2_fill_2 FILLER_65_374 ();
 sg13g2_fill_2 FILLER_65_384 ();
 sg13g2_decap_4 FILLER_65_400 ();
 sg13g2_decap_8 FILLER_65_416 ();
 sg13g2_decap_4 FILLER_65_427 ();
 sg13g2_fill_2 FILLER_65_453 ();
 sg13g2_fill_1 FILLER_65_455 ();
 sg13g2_decap_4 FILLER_65_477 ();
 sg13g2_fill_2 FILLER_65_481 ();
 sg13g2_fill_2 FILLER_65_512 ();
 sg13g2_fill_1 FILLER_65_514 ();
 sg13g2_fill_1 FILLER_65_523 ();
 sg13g2_fill_1 FILLER_65_543 ();
 sg13g2_fill_2 FILLER_65_549 ();
 sg13g2_decap_8 FILLER_65_556 ();
 sg13g2_fill_2 FILLER_65_563 ();
 sg13g2_fill_1 FILLER_65_565 ();
 sg13g2_decap_4 FILLER_65_571 ();
 sg13g2_fill_1 FILLER_65_575 ();
 sg13g2_decap_8 FILLER_65_584 ();
 sg13g2_decap_8 FILLER_65_591 ();
 sg13g2_decap_8 FILLER_65_598 ();
 sg13g2_fill_2 FILLER_65_605 ();
 sg13g2_decap_4 FILLER_65_632 ();
 sg13g2_fill_2 FILLER_65_643 ();
 sg13g2_fill_1 FILLER_65_660 ();
 sg13g2_fill_1 FILLER_65_667 ();
 sg13g2_fill_2 FILLER_65_683 ();
 sg13g2_fill_1 FILLER_65_685 ();
 sg13g2_fill_2 FILLER_65_698 ();
 sg13g2_fill_2 FILLER_65_708 ();
 sg13g2_fill_1 FILLER_65_710 ();
 sg13g2_decap_4 FILLER_65_719 ();
 sg13g2_fill_2 FILLER_65_778 ();
 sg13g2_fill_1 FILLER_65_780 ();
 sg13g2_fill_2 FILLER_65_790 ();
 sg13g2_decap_8 FILLER_65_808 ();
 sg13g2_decap_4 FILLER_65_815 ();
 sg13g2_fill_2 FILLER_65_840 ();
 sg13g2_fill_1 FILLER_65_842 ();
 sg13g2_decap_8 FILLER_65_857 ();
 sg13g2_decap_4 FILLER_65_864 ();
 sg13g2_fill_2 FILLER_65_868 ();
 sg13g2_decap_4 FILLER_65_878 ();
 sg13g2_fill_2 FILLER_65_893 ();
 sg13g2_decap_4 FILLER_65_921 ();
 sg13g2_fill_1 FILLER_65_968 ();
 sg13g2_fill_2 FILLER_65_979 ();
 sg13g2_decap_8 FILLER_65_986 ();
 sg13g2_decap_8 FILLER_65_993 ();
 sg13g2_decap_8 FILLER_65_1000 ();
 sg13g2_fill_1 FILLER_65_1012 ();
 sg13g2_fill_2 FILLER_65_1045 ();
 sg13g2_fill_1 FILLER_65_1047 ();
 sg13g2_fill_1 FILLER_65_1053 ();
 sg13g2_decap_8 FILLER_65_1081 ();
 sg13g2_decap_8 FILLER_65_1088 ();
 sg13g2_decap_8 FILLER_65_1095 ();
 sg13g2_decap_8 FILLER_65_1102 ();
 sg13g2_decap_8 FILLER_65_1109 ();
 sg13g2_decap_8 FILLER_65_1116 ();
 sg13g2_decap_8 FILLER_65_1123 ();
 sg13g2_decap_8 FILLER_65_1130 ();
 sg13g2_decap_8 FILLER_65_1137 ();
 sg13g2_decap_8 FILLER_65_1144 ();
 sg13g2_decap_8 FILLER_65_1151 ();
 sg13g2_decap_8 FILLER_65_1158 ();
 sg13g2_decap_8 FILLER_65_1165 ();
 sg13g2_decap_8 FILLER_65_1172 ();
 sg13g2_decap_8 FILLER_65_1179 ();
 sg13g2_decap_8 FILLER_65_1186 ();
 sg13g2_decap_8 FILLER_65_1193 ();
 sg13g2_decap_8 FILLER_65_1200 ();
 sg13g2_decap_8 FILLER_65_1207 ();
 sg13g2_decap_8 FILLER_65_1214 ();
 sg13g2_decap_8 FILLER_65_1221 ();
 sg13g2_decap_8 FILLER_65_1228 ();
 sg13g2_decap_8 FILLER_65_1235 ();
 sg13g2_decap_8 FILLER_65_1242 ();
 sg13g2_decap_8 FILLER_65_1249 ();
 sg13g2_decap_8 FILLER_65_1256 ();
 sg13g2_decap_8 FILLER_65_1263 ();
 sg13g2_decap_8 FILLER_65_1270 ();
 sg13g2_decap_8 FILLER_65_1277 ();
 sg13g2_decap_8 FILLER_65_1284 ();
 sg13g2_decap_8 FILLER_65_1291 ();
 sg13g2_decap_8 FILLER_65_1298 ();
 sg13g2_decap_8 FILLER_65_1305 ();
 sg13g2_decap_8 FILLER_65_1312 ();
 sg13g2_decap_8 FILLER_65_1319 ();
 sg13g2_decap_8 FILLER_65_1326 ();
 sg13g2_decap_8 FILLER_65_1333 ();
 sg13g2_decap_8 FILLER_65_1340 ();
 sg13g2_decap_8 FILLER_65_1347 ();
 sg13g2_decap_8 FILLER_65_1354 ();
 sg13g2_decap_8 FILLER_65_1361 ();
 sg13g2_decap_8 FILLER_65_1368 ();
 sg13g2_decap_8 FILLER_65_1375 ();
 sg13g2_decap_8 FILLER_65_1382 ();
 sg13g2_decap_8 FILLER_65_1389 ();
 sg13g2_decap_8 FILLER_65_1396 ();
 sg13g2_decap_8 FILLER_65_1403 ();
 sg13g2_decap_8 FILLER_65_1410 ();
 sg13g2_decap_8 FILLER_65_1417 ();
 sg13g2_decap_8 FILLER_65_1424 ();
 sg13g2_decap_8 FILLER_65_1431 ();
 sg13g2_decap_8 FILLER_65_1438 ();
 sg13g2_decap_8 FILLER_65_1445 ();
 sg13g2_decap_8 FILLER_65_1452 ();
 sg13g2_decap_8 FILLER_65_1459 ();
 sg13g2_decap_8 FILLER_65_1466 ();
 sg13g2_decap_8 FILLER_65_1473 ();
 sg13g2_decap_8 FILLER_65_1480 ();
 sg13g2_decap_8 FILLER_65_1487 ();
 sg13g2_decap_8 FILLER_65_1494 ();
 sg13g2_decap_8 FILLER_65_1501 ();
 sg13g2_decap_8 FILLER_65_1508 ();
 sg13g2_decap_8 FILLER_65_1515 ();
 sg13g2_decap_8 FILLER_65_1522 ();
 sg13g2_decap_8 FILLER_65_1529 ();
 sg13g2_decap_8 FILLER_65_1536 ();
 sg13g2_decap_8 FILLER_65_1543 ();
 sg13g2_decap_8 FILLER_65_1550 ();
 sg13g2_decap_8 FILLER_65_1557 ();
 sg13g2_decap_8 FILLER_65_1564 ();
 sg13g2_decap_8 FILLER_65_1571 ();
 sg13g2_decap_8 FILLER_65_1578 ();
 sg13g2_decap_8 FILLER_65_1585 ();
 sg13g2_decap_8 FILLER_65_1592 ();
 sg13g2_decap_8 FILLER_65_1599 ();
 sg13g2_decap_8 FILLER_65_1606 ();
 sg13g2_decap_8 FILLER_65_1613 ();
 sg13g2_decap_8 FILLER_65_1620 ();
 sg13g2_decap_8 FILLER_65_1627 ();
 sg13g2_decap_8 FILLER_65_1634 ();
 sg13g2_decap_8 FILLER_65_1641 ();
 sg13g2_decap_8 FILLER_65_1648 ();
 sg13g2_decap_8 FILLER_65_1655 ();
 sg13g2_decap_8 FILLER_65_1662 ();
 sg13g2_decap_8 FILLER_65_1669 ();
 sg13g2_decap_8 FILLER_65_1676 ();
 sg13g2_decap_8 FILLER_65_1683 ();
 sg13g2_decap_8 FILLER_65_1690 ();
 sg13g2_decap_8 FILLER_65_1697 ();
 sg13g2_decap_8 FILLER_65_1704 ();
 sg13g2_decap_8 FILLER_65_1711 ();
 sg13g2_decap_8 FILLER_65_1718 ();
 sg13g2_decap_8 FILLER_65_1725 ();
 sg13g2_decap_8 FILLER_65_1732 ();
 sg13g2_decap_8 FILLER_65_1739 ();
 sg13g2_decap_8 FILLER_65_1746 ();
 sg13g2_decap_8 FILLER_65_1753 ();
 sg13g2_decap_8 FILLER_65_1760 ();
 sg13g2_fill_1 FILLER_65_1767 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_8 FILLER_66_7 ();
 sg13g2_decap_8 FILLER_66_14 ();
 sg13g2_decap_8 FILLER_66_21 ();
 sg13g2_decap_8 FILLER_66_28 ();
 sg13g2_decap_8 FILLER_66_35 ();
 sg13g2_decap_8 FILLER_66_42 ();
 sg13g2_decap_4 FILLER_66_49 ();
 sg13g2_fill_1 FILLER_66_53 ();
 sg13g2_decap_4 FILLER_66_83 ();
 sg13g2_fill_2 FILLER_66_109 ();
 sg13g2_fill_2 FILLER_66_123 ();
 sg13g2_fill_2 FILLER_66_148 ();
 sg13g2_fill_2 FILLER_66_154 ();
 sg13g2_fill_1 FILLER_66_156 ();
 sg13g2_fill_1 FILLER_66_166 ();
 sg13g2_decap_8 FILLER_66_177 ();
 sg13g2_fill_1 FILLER_66_184 ();
 sg13g2_fill_1 FILLER_66_194 ();
 sg13g2_fill_2 FILLER_66_202 ();
 sg13g2_decap_8 FILLER_66_218 ();
 sg13g2_decap_4 FILLER_66_225 ();
 sg13g2_fill_2 FILLER_66_238 ();
 sg13g2_fill_2 FILLER_66_254 ();
 sg13g2_fill_1 FILLER_66_256 ();
 sg13g2_fill_2 FILLER_66_296 ();
 sg13g2_fill_2 FILLER_66_340 ();
 sg13g2_fill_1 FILLER_66_342 ();
 sg13g2_fill_2 FILLER_66_356 ();
 sg13g2_fill_1 FILLER_66_371 ();
 sg13g2_decap_8 FILLER_66_384 ();
 sg13g2_fill_2 FILLER_66_391 ();
 sg13g2_fill_1 FILLER_66_393 ();
 sg13g2_decap_4 FILLER_66_412 ();
 sg13g2_fill_1 FILLER_66_416 ();
 sg13g2_fill_1 FILLER_66_434 ();
 sg13g2_fill_1 FILLER_66_443 ();
 sg13g2_decap_4 FILLER_66_456 ();
 sg13g2_fill_2 FILLER_66_460 ();
 sg13g2_fill_2 FILLER_66_471 ();
 sg13g2_fill_1 FILLER_66_473 ();
 sg13g2_fill_2 FILLER_66_482 ();
 sg13g2_fill_1 FILLER_66_484 ();
 sg13g2_fill_1 FILLER_66_490 ();
 sg13g2_decap_4 FILLER_66_517 ();
 sg13g2_decap_4 FILLER_66_534 ();
 sg13g2_fill_2 FILLER_66_553 ();
 sg13g2_decap_8 FILLER_66_560 ();
 sg13g2_fill_2 FILLER_66_567 ();
 sg13g2_decap_4 FILLER_66_574 ();
 sg13g2_fill_2 FILLER_66_578 ();
 sg13g2_decap_8 FILLER_66_590 ();
 sg13g2_decap_4 FILLER_66_597 ();
 sg13g2_fill_1 FILLER_66_601 ();
 sg13g2_decap_8 FILLER_66_608 ();
 sg13g2_fill_2 FILLER_66_615 ();
 sg13g2_fill_1 FILLER_66_622 ();
 sg13g2_decap_8 FILLER_66_628 ();
 sg13g2_fill_2 FILLER_66_635 ();
 sg13g2_fill_1 FILLER_66_637 ();
 sg13g2_fill_1 FILLER_66_652 ();
 sg13g2_decap_4 FILLER_66_669 ();
 sg13g2_fill_1 FILLER_66_673 ();
 sg13g2_decap_8 FILLER_66_684 ();
 sg13g2_fill_2 FILLER_66_691 ();
 sg13g2_fill_1 FILLER_66_698 ();
 sg13g2_fill_1 FILLER_66_709 ();
 sg13g2_fill_2 FILLER_66_738 ();
 sg13g2_fill_2 FILLER_66_753 ();
 sg13g2_fill_2 FILLER_66_763 ();
 sg13g2_fill_2 FILLER_66_796 ();
 sg13g2_fill_1 FILLER_66_798 ();
 sg13g2_fill_2 FILLER_66_814 ();
 sg13g2_fill_1 FILLER_66_833 ();
 sg13g2_fill_2 FILLER_66_874 ();
 sg13g2_fill_1 FILLER_66_876 ();
 sg13g2_fill_1 FILLER_66_889 ();
 sg13g2_fill_2 FILLER_66_916 ();
 sg13g2_fill_1 FILLER_66_918 ();
 sg13g2_fill_1 FILLER_66_924 ();
 sg13g2_fill_2 FILLER_66_931 ();
 sg13g2_fill_2 FILLER_66_964 ();
 sg13g2_fill_1 FILLER_66_966 ();
 sg13g2_fill_2 FILLER_66_989 ();
 sg13g2_fill_1 FILLER_66_991 ();
 sg13g2_fill_1 FILLER_66_1004 ();
 sg13g2_decap_8 FILLER_66_1033 ();
 sg13g2_fill_2 FILLER_66_1049 ();
 sg13g2_fill_1 FILLER_66_1051 ();
 sg13g2_decap_8 FILLER_66_1078 ();
 sg13g2_decap_8 FILLER_66_1085 ();
 sg13g2_decap_8 FILLER_66_1092 ();
 sg13g2_decap_8 FILLER_66_1099 ();
 sg13g2_decap_8 FILLER_66_1106 ();
 sg13g2_decap_8 FILLER_66_1113 ();
 sg13g2_decap_8 FILLER_66_1120 ();
 sg13g2_decap_8 FILLER_66_1127 ();
 sg13g2_decap_8 FILLER_66_1134 ();
 sg13g2_decap_8 FILLER_66_1141 ();
 sg13g2_decap_8 FILLER_66_1148 ();
 sg13g2_decap_8 FILLER_66_1155 ();
 sg13g2_decap_8 FILLER_66_1162 ();
 sg13g2_decap_8 FILLER_66_1169 ();
 sg13g2_decap_8 FILLER_66_1176 ();
 sg13g2_decap_8 FILLER_66_1183 ();
 sg13g2_decap_8 FILLER_66_1190 ();
 sg13g2_decap_8 FILLER_66_1197 ();
 sg13g2_decap_8 FILLER_66_1204 ();
 sg13g2_decap_8 FILLER_66_1211 ();
 sg13g2_decap_8 FILLER_66_1218 ();
 sg13g2_decap_8 FILLER_66_1225 ();
 sg13g2_decap_8 FILLER_66_1232 ();
 sg13g2_decap_8 FILLER_66_1239 ();
 sg13g2_decap_8 FILLER_66_1246 ();
 sg13g2_decap_8 FILLER_66_1253 ();
 sg13g2_decap_8 FILLER_66_1260 ();
 sg13g2_decap_8 FILLER_66_1267 ();
 sg13g2_decap_8 FILLER_66_1274 ();
 sg13g2_decap_8 FILLER_66_1281 ();
 sg13g2_decap_8 FILLER_66_1288 ();
 sg13g2_decap_8 FILLER_66_1295 ();
 sg13g2_decap_8 FILLER_66_1302 ();
 sg13g2_decap_8 FILLER_66_1309 ();
 sg13g2_decap_8 FILLER_66_1316 ();
 sg13g2_decap_8 FILLER_66_1323 ();
 sg13g2_decap_8 FILLER_66_1330 ();
 sg13g2_decap_8 FILLER_66_1337 ();
 sg13g2_decap_8 FILLER_66_1344 ();
 sg13g2_decap_8 FILLER_66_1351 ();
 sg13g2_decap_8 FILLER_66_1358 ();
 sg13g2_decap_8 FILLER_66_1365 ();
 sg13g2_decap_8 FILLER_66_1372 ();
 sg13g2_decap_8 FILLER_66_1379 ();
 sg13g2_decap_8 FILLER_66_1386 ();
 sg13g2_decap_8 FILLER_66_1393 ();
 sg13g2_decap_8 FILLER_66_1400 ();
 sg13g2_decap_8 FILLER_66_1407 ();
 sg13g2_decap_8 FILLER_66_1414 ();
 sg13g2_decap_8 FILLER_66_1421 ();
 sg13g2_decap_8 FILLER_66_1428 ();
 sg13g2_decap_8 FILLER_66_1435 ();
 sg13g2_decap_8 FILLER_66_1442 ();
 sg13g2_decap_8 FILLER_66_1449 ();
 sg13g2_decap_8 FILLER_66_1456 ();
 sg13g2_decap_8 FILLER_66_1463 ();
 sg13g2_decap_8 FILLER_66_1470 ();
 sg13g2_decap_8 FILLER_66_1477 ();
 sg13g2_decap_8 FILLER_66_1484 ();
 sg13g2_decap_8 FILLER_66_1491 ();
 sg13g2_decap_8 FILLER_66_1498 ();
 sg13g2_decap_8 FILLER_66_1505 ();
 sg13g2_decap_8 FILLER_66_1512 ();
 sg13g2_decap_8 FILLER_66_1519 ();
 sg13g2_decap_8 FILLER_66_1526 ();
 sg13g2_decap_8 FILLER_66_1533 ();
 sg13g2_decap_8 FILLER_66_1540 ();
 sg13g2_decap_8 FILLER_66_1547 ();
 sg13g2_decap_8 FILLER_66_1554 ();
 sg13g2_decap_8 FILLER_66_1561 ();
 sg13g2_decap_8 FILLER_66_1568 ();
 sg13g2_decap_8 FILLER_66_1575 ();
 sg13g2_decap_8 FILLER_66_1582 ();
 sg13g2_decap_8 FILLER_66_1589 ();
 sg13g2_decap_8 FILLER_66_1596 ();
 sg13g2_decap_8 FILLER_66_1603 ();
 sg13g2_decap_8 FILLER_66_1610 ();
 sg13g2_decap_8 FILLER_66_1617 ();
 sg13g2_decap_8 FILLER_66_1624 ();
 sg13g2_decap_8 FILLER_66_1631 ();
 sg13g2_decap_8 FILLER_66_1638 ();
 sg13g2_decap_8 FILLER_66_1645 ();
 sg13g2_decap_8 FILLER_66_1652 ();
 sg13g2_decap_8 FILLER_66_1659 ();
 sg13g2_decap_8 FILLER_66_1666 ();
 sg13g2_decap_8 FILLER_66_1673 ();
 sg13g2_decap_8 FILLER_66_1680 ();
 sg13g2_decap_8 FILLER_66_1687 ();
 sg13g2_decap_8 FILLER_66_1694 ();
 sg13g2_decap_8 FILLER_66_1701 ();
 sg13g2_decap_8 FILLER_66_1708 ();
 sg13g2_decap_8 FILLER_66_1715 ();
 sg13g2_decap_8 FILLER_66_1722 ();
 sg13g2_decap_8 FILLER_66_1729 ();
 sg13g2_decap_8 FILLER_66_1736 ();
 sg13g2_decap_8 FILLER_66_1743 ();
 sg13g2_decap_8 FILLER_66_1750 ();
 sg13g2_decap_8 FILLER_66_1757 ();
 sg13g2_decap_4 FILLER_66_1764 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_8 FILLER_67_7 ();
 sg13g2_decap_8 FILLER_67_14 ();
 sg13g2_decap_8 FILLER_67_21 ();
 sg13g2_decap_8 FILLER_67_28 ();
 sg13g2_decap_8 FILLER_67_35 ();
 sg13g2_decap_8 FILLER_67_42 ();
 sg13g2_decap_8 FILLER_67_49 ();
 sg13g2_decap_4 FILLER_67_56 ();
 sg13g2_fill_2 FILLER_67_60 ();
 sg13g2_fill_1 FILLER_67_87 ();
 sg13g2_decap_4 FILLER_67_111 ();
 sg13g2_fill_2 FILLER_67_121 ();
 sg13g2_fill_1 FILLER_67_183 ();
 sg13g2_fill_2 FILLER_67_210 ();
 sg13g2_fill_1 FILLER_67_212 ();
 sg13g2_fill_2 FILLER_67_222 ();
 sg13g2_decap_4 FILLER_67_271 ();
 sg13g2_fill_1 FILLER_67_275 ();
 sg13g2_fill_2 FILLER_67_306 ();
 sg13g2_fill_1 FILLER_67_308 ();
 sg13g2_fill_2 FILLER_67_340 ();
 sg13g2_fill_1 FILLER_67_342 ();
 sg13g2_fill_1 FILLER_67_356 ();
 sg13g2_fill_2 FILLER_67_365 ();
 sg13g2_fill_1 FILLER_67_367 ();
 sg13g2_fill_2 FILLER_67_395 ();
 sg13g2_decap_4 FILLER_67_420 ();
 sg13g2_decap_4 FILLER_67_429 ();
 sg13g2_fill_2 FILLER_67_433 ();
 sg13g2_fill_2 FILLER_67_439 ();
 sg13g2_fill_1 FILLER_67_446 ();
 sg13g2_fill_2 FILLER_67_450 ();
 sg13g2_fill_1 FILLER_67_452 ();
 sg13g2_decap_4 FILLER_67_458 ();
 sg13g2_decap_4 FILLER_67_475 ();
 sg13g2_fill_1 FILLER_67_479 ();
 sg13g2_decap_8 FILLER_67_497 ();
 sg13g2_fill_2 FILLER_67_504 ();
 sg13g2_fill_1 FILLER_67_506 ();
 sg13g2_decap_4 FILLER_67_524 ();
 sg13g2_fill_1 FILLER_67_528 ();
 sg13g2_decap_4 FILLER_67_548 ();
 sg13g2_fill_2 FILLER_67_562 ();
 sg13g2_fill_1 FILLER_67_564 ();
 sg13g2_decap_4 FILLER_67_594 ();
 sg13g2_fill_1 FILLER_67_637 ();
 sg13g2_fill_2 FILLER_67_656 ();
 sg13g2_fill_2 FILLER_67_666 ();
 sg13g2_fill_1 FILLER_67_668 ();
 sg13g2_fill_2 FILLER_67_692 ();
 sg13g2_fill_2 FILLER_67_702 ();
 sg13g2_decap_8 FILLER_67_713 ();
 sg13g2_fill_2 FILLER_67_720 ();
 sg13g2_decap_4 FILLER_67_730 ();
 sg13g2_decap_8 FILLER_67_759 ();
 sg13g2_fill_2 FILLER_67_831 ();
 sg13g2_fill_1 FILLER_67_833 ();
 sg13g2_fill_2 FILLER_67_856 ();
 sg13g2_fill_2 FILLER_67_875 ();
 sg13g2_fill_2 FILLER_67_886 ();
 sg13g2_fill_1 FILLER_67_888 ();
 sg13g2_decap_4 FILLER_67_936 ();
 sg13g2_fill_2 FILLER_67_940 ();
 sg13g2_decap_8 FILLER_67_960 ();
 sg13g2_fill_1 FILLER_67_967 ();
 sg13g2_fill_1 FILLER_67_972 ();
 sg13g2_fill_1 FILLER_67_984 ();
 sg13g2_decap_8 FILLER_67_990 ();
 sg13g2_decap_8 FILLER_67_997 ();
 sg13g2_decap_4 FILLER_67_1004 ();
 sg13g2_decap_8 FILLER_67_1033 ();
 sg13g2_fill_1 FILLER_67_1040 ();
 sg13g2_decap_4 FILLER_67_1046 ();
 sg13g2_decap_8 FILLER_67_1073 ();
 sg13g2_decap_8 FILLER_67_1080 ();
 sg13g2_decap_8 FILLER_67_1087 ();
 sg13g2_decap_8 FILLER_67_1094 ();
 sg13g2_decap_8 FILLER_67_1101 ();
 sg13g2_decap_8 FILLER_67_1108 ();
 sg13g2_decap_8 FILLER_67_1115 ();
 sg13g2_decap_8 FILLER_67_1122 ();
 sg13g2_decap_8 FILLER_67_1129 ();
 sg13g2_decap_8 FILLER_67_1136 ();
 sg13g2_decap_8 FILLER_67_1143 ();
 sg13g2_decap_8 FILLER_67_1150 ();
 sg13g2_decap_8 FILLER_67_1157 ();
 sg13g2_decap_8 FILLER_67_1164 ();
 sg13g2_decap_8 FILLER_67_1171 ();
 sg13g2_decap_8 FILLER_67_1178 ();
 sg13g2_decap_8 FILLER_67_1185 ();
 sg13g2_decap_8 FILLER_67_1192 ();
 sg13g2_decap_8 FILLER_67_1199 ();
 sg13g2_decap_8 FILLER_67_1206 ();
 sg13g2_decap_8 FILLER_67_1213 ();
 sg13g2_decap_8 FILLER_67_1220 ();
 sg13g2_decap_8 FILLER_67_1227 ();
 sg13g2_decap_8 FILLER_67_1234 ();
 sg13g2_decap_8 FILLER_67_1241 ();
 sg13g2_decap_8 FILLER_67_1248 ();
 sg13g2_decap_8 FILLER_67_1255 ();
 sg13g2_decap_8 FILLER_67_1262 ();
 sg13g2_decap_8 FILLER_67_1269 ();
 sg13g2_decap_8 FILLER_67_1276 ();
 sg13g2_decap_8 FILLER_67_1283 ();
 sg13g2_decap_8 FILLER_67_1290 ();
 sg13g2_decap_8 FILLER_67_1297 ();
 sg13g2_decap_8 FILLER_67_1304 ();
 sg13g2_decap_8 FILLER_67_1311 ();
 sg13g2_decap_8 FILLER_67_1318 ();
 sg13g2_decap_8 FILLER_67_1325 ();
 sg13g2_decap_8 FILLER_67_1332 ();
 sg13g2_decap_8 FILLER_67_1339 ();
 sg13g2_decap_8 FILLER_67_1346 ();
 sg13g2_decap_8 FILLER_67_1353 ();
 sg13g2_decap_8 FILLER_67_1360 ();
 sg13g2_decap_8 FILLER_67_1367 ();
 sg13g2_decap_8 FILLER_67_1374 ();
 sg13g2_decap_8 FILLER_67_1381 ();
 sg13g2_decap_8 FILLER_67_1388 ();
 sg13g2_decap_8 FILLER_67_1395 ();
 sg13g2_decap_8 FILLER_67_1402 ();
 sg13g2_decap_8 FILLER_67_1409 ();
 sg13g2_decap_8 FILLER_67_1416 ();
 sg13g2_decap_8 FILLER_67_1423 ();
 sg13g2_decap_8 FILLER_67_1430 ();
 sg13g2_decap_8 FILLER_67_1437 ();
 sg13g2_decap_8 FILLER_67_1444 ();
 sg13g2_decap_8 FILLER_67_1451 ();
 sg13g2_decap_8 FILLER_67_1458 ();
 sg13g2_decap_8 FILLER_67_1465 ();
 sg13g2_decap_8 FILLER_67_1472 ();
 sg13g2_decap_8 FILLER_67_1479 ();
 sg13g2_decap_8 FILLER_67_1486 ();
 sg13g2_decap_8 FILLER_67_1493 ();
 sg13g2_decap_8 FILLER_67_1500 ();
 sg13g2_decap_8 FILLER_67_1507 ();
 sg13g2_decap_8 FILLER_67_1514 ();
 sg13g2_decap_8 FILLER_67_1521 ();
 sg13g2_decap_8 FILLER_67_1528 ();
 sg13g2_decap_8 FILLER_67_1535 ();
 sg13g2_decap_8 FILLER_67_1542 ();
 sg13g2_decap_8 FILLER_67_1549 ();
 sg13g2_decap_8 FILLER_67_1556 ();
 sg13g2_decap_8 FILLER_67_1563 ();
 sg13g2_decap_8 FILLER_67_1570 ();
 sg13g2_decap_8 FILLER_67_1577 ();
 sg13g2_decap_8 FILLER_67_1584 ();
 sg13g2_decap_8 FILLER_67_1591 ();
 sg13g2_decap_8 FILLER_67_1598 ();
 sg13g2_decap_8 FILLER_67_1605 ();
 sg13g2_decap_8 FILLER_67_1612 ();
 sg13g2_decap_8 FILLER_67_1619 ();
 sg13g2_decap_8 FILLER_67_1626 ();
 sg13g2_decap_8 FILLER_67_1633 ();
 sg13g2_decap_8 FILLER_67_1640 ();
 sg13g2_decap_8 FILLER_67_1647 ();
 sg13g2_decap_8 FILLER_67_1654 ();
 sg13g2_decap_8 FILLER_67_1661 ();
 sg13g2_decap_8 FILLER_67_1668 ();
 sg13g2_decap_8 FILLER_67_1675 ();
 sg13g2_decap_8 FILLER_67_1682 ();
 sg13g2_decap_8 FILLER_67_1689 ();
 sg13g2_decap_8 FILLER_67_1696 ();
 sg13g2_decap_8 FILLER_67_1703 ();
 sg13g2_decap_8 FILLER_67_1710 ();
 sg13g2_decap_8 FILLER_67_1717 ();
 sg13g2_decap_8 FILLER_67_1724 ();
 sg13g2_decap_8 FILLER_67_1731 ();
 sg13g2_decap_8 FILLER_67_1738 ();
 sg13g2_decap_8 FILLER_67_1745 ();
 sg13g2_decap_8 FILLER_67_1752 ();
 sg13g2_decap_8 FILLER_67_1759 ();
 sg13g2_fill_2 FILLER_67_1766 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_8 FILLER_68_7 ();
 sg13g2_decap_8 FILLER_68_14 ();
 sg13g2_decap_8 FILLER_68_21 ();
 sg13g2_decap_8 FILLER_68_28 ();
 sg13g2_decap_8 FILLER_68_35 ();
 sg13g2_decap_8 FILLER_68_42 ();
 sg13g2_fill_1 FILLER_68_49 ();
 sg13g2_fill_2 FILLER_68_76 ();
 sg13g2_fill_1 FILLER_68_78 ();
 sg13g2_fill_2 FILLER_68_101 ();
 sg13g2_fill_1 FILLER_68_111 ();
 sg13g2_decap_8 FILLER_68_130 ();
 sg13g2_decap_4 FILLER_68_159 ();
 sg13g2_fill_1 FILLER_68_163 ();
 sg13g2_fill_2 FILLER_68_184 ();
 sg13g2_fill_1 FILLER_68_232 ();
 sg13g2_fill_2 FILLER_68_238 ();
 sg13g2_fill_1 FILLER_68_240 ();
 sg13g2_fill_2 FILLER_68_302 ();
 sg13g2_fill_1 FILLER_68_304 ();
 sg13g2_fill_2 FILLER_68_310 ();
 sg13g2_fill_1 FILLER_68_312 ();
 sg13g2_fill_1 FILLER_68_318 ();
 sg13g2_fill_1 FILLER_68_323 ();
 sg13g2_fill_2 FILLER_68_332 ();
 sg13g2_fill_1 FILLER_68_334 ();
 sg13g2_decap_8 FILLER_68_340 ();
 sg13g2_decap_8 FILLER_68_347 ();
 sg13g2_fill_1 FILLER_68_354 ();
 sg13g2_fill_1 FILLER_68_360 ();
 sg13g2_fill_2 FILLER_68_371 ();
 sg13g2_fill_2 FILLER_68_377 ();
 sg13g2_decap_8 FILLER_68_386 ();
 sg13g2_fill_2 FILLER_68_397 ();
 sg13g2_fill_1 FILLER_68_411 ();
 sg13g2_fill_2 FILLER_68_459 ();
 sg13g2_fill_1 FILLER_68_474 ();
 sg13g2_fill_2 FILLER_68_495 ();
 sg13g2_decap_4 FILLER_68_502 ();
 sg13g2_fill_2 FILLER_68_506 ();
 sg13g2_decap_8 FILLER_68_530 ();
 sg13g2_decap_4 FILLER_68_537 ();
 sg13g2_fill_2 FILLER_68_541 ();
 sg13g2_decap_8 FILLER_68_568 ();
 sg13g2_decap_4 FILLER_68_575 ();
 sg13g2_fill_2 FILLER_68_579 ();
 sg13g2_fill_2 FILLER_68_591 ();
 sg13g2_fill_1 FILLER_68_593 ();
 sg13g2_fill_2 FILLER_68_605 ();
 sg13g2_decap_4 FILLER_68_612 ();
 sg13g2_decap_8 FILLER_68_643 ();
 sg13g2_fill_2 FILLER_68_650 ();
 sg13g2_fill_1 FILLER_68_652 ();
 sg13g2_decap_8 FILLER_68_663 ();
 sg13g2_decap_8 FILLER_68_670 ();
 sg13g2_fill_2 FILLER_68_677 ();
 sg13g2_fill_1 FILLER_68_679 ();
 sg13g2_decap_4 FILLER_68_717 ();
 sg13g2_fill_2 FILLER_68_721 ();
 sg13g2_decap_4 FILLER_68_740 ();
 sg13g2_decap_4 FILLER_68_753 ();
 sg13g2_fill_2 FILLER_68_793 ();
 sg13g2_decap_4 FILLER_68_827 ();
 sg13g2_fill_1 FILLER_68_831 ();
 sg13g2_fill_2 FILLER_68_835 ();
 sg13g2_fill_2 FILLER_68_863 ();
 sg13g2_fill_1 FILLER_68_865 ();
 sg13g2_decap_8 FILLER_68_884 ();
 sg13g2_fill_2 FILLER_68_891 ();
 sg13g2_fill_1 FILLER_68_919 ();
 sg13g2_fill_1 FILLER_68_923 ();
 sg13g2_decap_8 FILLER_68_933 ();
 sg13g2_decap_4 FILLER_68_940 ();
 sg13g2_fill_1 FILLER_68_944 ();
 sg13g2_decap_4 FILLER_68_967 ();
 sg13g2_decap_4 FILLER_68_984 ();
 sg13g2_fill_2 FILLER_68_996 ();
 sg13g2_decap_4 FILLER_68_1034 ();
 sg13g2_fill_2 FILLER_68_1038 ();
 sg13g2_decap_8 FILLER_68_1066 ();
 sg13g2_decap_8 FILLER_68_1073 ();
 sg13g2_decap_8 FILLER_68_1080 ();
 sg13g2_decap_8 FILLER_68_1087 ();
 sg13g2_decap_8 FILLER_68_1094 ();
 sg13g2_decap_8 FILLER_68_1101 ();
 sg13g2_decap_8 FILLER_68_1108 ();
 sg13g2_decap_8 FILLER_68_1115 ();
 sg13g2_decap_8 FILLER_68_1122 ();
 sg13g2_decap_8 FILLER_68_1129 ();
 sg13g2_decap_8 FILLER_68_1136 ();
 sg13g2_decap_8 FILLER_68_1143 ();
 sg13g2_decap_8 FILLER_68_1150 ();
 sg13g2_decap_8 FILLER_68_1157 ();
 sg13g2_decap_8 FILLER_68_1164 ();
 sg13g2_decap_8 FILLER_68_1171 ();
 sg13g2_decap_8 FILLER_68_1178 ();
 sg13g2_decap_8 FILLER_68_1185 ();
 sg13g2_decap_8 FILLER_68_1192 ();
 sg13g2_decap_8 FILLER_68_1199 ();
 sg13g2_decap_8 FILLER_68_1206 ();
 sg13g2_decap_8 FILLER_68_1213 ();
 sg13g2_decap_8 FILLER_68_1220 ();
 sg13g2_decap_8 FILLER_68_1227 ();
 sg13g2_decap_8 FILLER_68_1234 ();
 sg13g2_decap_8 FILLER_68_1241 ();
 sg13g2_decap_8 FILLER_68_1248 ();
 sg13g2_decap_8 FILLER_68_1255 ();
 sg13g2_decap_8 FILLER_68_1262 ();
 sg13g2_decap_8 FILLER_68_1269 ();
 sg13g2_decap_8 FILLER_68_1276 ();
 sg13g2_decap_8 FILLER_68_1283 ();
 sg13g2_decap_8 FILLER_68_1290 ();
 sg13g2_decap_8 FILLER_68_1297 ();
 sg13g2_decap_8 FILLER_68_1304 ();
 sg13g2_decap_8 FILLER_68_1311 ();
 sg13g2_decap_8 FILLER_68_1318 ();
 sg13g2_decap_8 FILLER_68_1325 ();
 sg13g2_decap_8 FILLER_68_1332 ();
 sg13g2_decap_8 FILLER_68_1339 ();
 sg13g2_decap_8 FILLER_68_1346 ();
 sg13g2_decap_8 FILLER_68_1353 ();
 sg13g2_decap_8 FILLER_68_1360 ();
 sg13g2_decap_8 FILLER_68_1367 ();
 sg13g2_decap_8 FILLER_68_1374 ();
 sg13g2_decap_8 FILLER_68_1381 ();
 sg13g2_decap_8 FILLER_68_1388 ();
 sg13g2_decap_8 FILLER_68_1395 ();
 sg13g2_decap_8 FILLER_68_1402 ();
 sg13g2_decap_8 FILLER_68_1409 ();
 sg13g2_decap_8 FILLER_68_1416 ();
 sg13g2_decap_8 FILLER_68_1423 ();
 sg13g2_decap_8 FILLER_68_1430 ();
 sg13g2_decap_8 FILLER_68_1437 ();
 sg13g2_decap_8 FILLER_68_1444 ();
 sg13g2_decap_8 FILLER_68_1451 ();
 sg13g2_decap_8 FILLER_68_1458 ();
 sg13g2_decap_8 FILLER_68_1465 ();
 sg13g2_decap_8 FILLER_68_1472 ();
 sg13g2_decap_8 FILLER_68_1479 ();
 sg13g2_decap_8 FILLER_68_1486 ();
 sg13g2_decap_8 FILLER_68_1493 ();
 sg13g2_decap_8 FILLER_68_1500 ();
 sg13g2_decap_8 FILLER_68_1507 ();
 sg13g2_decap_8 FILLER_68_1514 ();
 sg13g2_decap_8 FILLER_68_1521 ();
 sg13g2_decap_8 FILLER_68_1528 ();
 sg13g2_decap_8 FILLER_68_1535 ();
 sg13g2_decap_8 FILLER_68_1542 ();
 sg13g2_decap_8 FILLER_68_1549 ();
 sg13g2_decap_8 FILLER_68_1556 ();
 sg13g2_decap_8 FILLER_68_1563 ();
 sg13g2_decap_8 FILLER_68_1570 ();
 sg13g2_decap_8 FILLER_68_1577 ();
 sg13g2_decap_8 FILLER_68_1584 ();
 sg13g2_decap_8 FILLER_68_1591 ();
 sg13g2_decap_8 FILLER_68_1598 ();
 sg13g2_decap_8 FILLER_68_1605 ();
 sg13g2_decap_8 FILLER_68_1612 ();
 sg13g2_decap_8 FILLER_68_1619 ();
 sg13g2_decap_8 FILLER_68_1626 ();
 sg13g2_decap_8 FILLER_68_1633 ();
 sg13g2_decap_8 FILLER_68_1640 ();
 sg13g2_decap_8 FILLER_68_1647 ();
 sg13g2_decap_8 FILLER_68_1654 ();
 sg13g2_decap_8 FILLER_68_1661 ();
 sg13g2_decap_8 FILLER_68_1668 ();
 sg13g2_decap_8 FILLER_68_1675 ();
 sg13g2_decap_8 FILLER_68_1682 ();
 sg13g2_decap_8 FILLER_68_1689 ();
 sg13g2_decap_8 FILLER_68_1696 ();
 sg13g2_decap_8 FILLER_68_1703 ();
 sg13g2_decap_8 FILLER_68_1710 ();
 sg13g2_decap_8 FILLER_68_1717 ();
 sg13g2_decap_8 FILLER_68_1724 ();
 sg13g2_decap_8 FILLER_68_1731 ();
 sg13g2_decap_8 FILLER_68_1738 ();
 sg13g2_decap_8 FILLER_68_1745 ();
 sg13g2_decap_8 FILLER_68_1752 ();
 sg13g2_decap_8 FILLER_68_1759 ();
 sg13g2_fill_2 FILLER_68_1766 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_8 FILLER_69_7 ();
 sg13g2_decap_8 FILLER_69_14 ();
 sg13g2_decap_8 FILLER_69_21 ();
 sg13g2_decap_8 FILLER_69_28 ();
 sg13g2_decap_8 FILLER_69_35 ();
 sg13g2_fill_2 FILLER_69_42 ();
 sg13g2_fill_2 FILLER_69_53 ();
 sg13g2_fill_1 FILLER_69_60 ();
 sg13g2_fill_2 FILLER_69_89 ();
 sg13g2_fill_1 FILLER_69_118 ();
 sg13g2_decap_8 FILLER_69_127 ();
 sg13g2_fill_2 FILLER_69_134 ();
 sg13g2_decap_4 FILLER_69_165 ();
 sg13g2_fill_2 FILLER_69_179 ();
 sg13g2_fill_1 FILLER_69_181 ();
 sg13g2_decap_8 FILLER_69_187 ();
 sg13g2_fill_2 FILLER_69_194 ();
 sg13g2_decap_4 FILLER_69_200 ();
 sg13g2_decap_4 FILLER_69_217 ();
 sg13g2_decap_4 FILLER_69_266 ();
 sg13g2_fill_2 FILLER_69_270 ();
 sg13g2_fill_2 FILLER_69_342 ();
 sg13g2_fill_1 FILLER_69_344 ();
 sg13g2_fill_2 FILLER_69_350 ();
 sg13g2_fill_1 FILLER_69_352 ();
 sg13g2_fill_2 FILLER_69_370 ();
 sg13g2_fill_2 FILLER_69_389 ();
 sg13g2_fill_2 FILLER_69_406 ();
 sg13g2_fill_1 FILLER_69_408 ();
 sg13g2_decap_4 FILLER_69_423 ();
 sg13g2_decap_4 FILLER_69_435 ();
 sg13g2_fill_1 FILLER_69_439 ();
 sg13g2_fill_2 FILLER_69_456 ();
 sg13g2_fill_1 FILLER_69_458 ();
 sg13g2_decap_8 FILLER_69_474 ();
 sg13g2_decap_4 FILLER_69_513 ();
 sg13g2_fill_1 FILLER_69_529 ();
 sg13g2_decap_4 FILLER_69_547 ();
 sg13g2_decap_8 FILLER_69_563 ();
 sg13g2_decap_8 FILLER_69_585 ();
 sg13g2_decap_4 FILLER_69_592 ();
 sg13g2_fill_1 FILLER_69_596 ();
 sg13g2_fill_2 FILLER_69_602 ();
 sg13g2_fill_1 FILLER_69_604 ();
 sg13g2_decap_8 FILLER_69_617 ();
 sg13g2_fill_1 FILLER_69_624 ();
 sg13g2_fill_1 FILLER_69_641 ();
 sg13g2_fill_2 FILLER_69_668 ();
 sg13g2_fill_2 FILLER_69_696 ();
 sg13g2_fill_1 FILLER_69_698 ();
 sg13g2_decap_8 FILLER_69_725 ();
 sg13g2_fill_2 FILLER_69_732 ();
 sg13g2_fill_1 FILLER_69_734 ();
 sg13g2_fill_2 FILLER_69_740 ();
 sg13g2_decap_4 FILLER_69_755 ();
 sg13g2_fill_1 FILLER_69_759 ();
 sg13g2_fill_1 FILLER_69_766 ();
 sg13g2_decap_4 FILLER_69_786 ();
 sg13g2_fill_1 FILLER_69_800 ();
 sg13g2_decap_4 FILLER_69_827 ();
 sg13g2_fill_1 FILLER_69_831 ();
 sg13g2_decap_8 FILLER_69_858 ();
 sg13g2_decap_4 FILLER_69_865 ();
 sg13g2_fill_1 FILLER_69_869 ();
 sg13g2_fill_1 FILLER_69_912 ();
 sg13g2_decap_4 FILLER_69_963 ();
 sg13g2_fill_2 FILLER_69_967 ();
 sg13g2_fill_2 FILLER_69_979 ();
 sg13g2_decap_8 FILLER_69_994 ();
 sg13g2_decap_4 FILLER_69_1001 ();
 sg13g2_fill_1 FILLER_69_1005 ();
 sg13g2_decap_8 FILLER_69_1032 ();
 sg13g2_fill_1 FILLER_69_1039 ();
 sg13g2_fill_1 FILLER_69_1050 ();
 sg13g2_fill_2 FILLER_69_1061 ();
 sg13g2_fill_1 FILLER_69_1063 ();
 sg13g2_decap_8 FILLER_69_1072 ();
 sg13g2_decap_8 FILLER_69_1079 ();
 sg13g2_decap_8 FILLER_69_1086 ();
 sg13g2_decap_8 FILLER_69_1093 ();
 sg13g2_decap_8 FILLER_69_1100 ();
 sg13g2_decap_8 FILLER_69_1107 ();
 sg13g2_decap_8 FILLER_69_1114 ();
 sg13g2_decap_8 FILLER_69_1121 ();
 sg13g2_decap_8 FILLER_69_1128 ();
 sg13g2_decap_8 FILLER_69_1135 ();
 sg13g2_decap_8 FILLER_69_1142 ();
 sg13g2_decap_8 FILLER_69_1149 ();
 sg13g2_decap_8 FILLER_69_1156 ();
 sg13g2_decap_8 FILLER_69_1163 ();
 sg13g2_decap_8 FILLER_69_1170 ();
 sg13g2_decap_8 FILLER_69_1177 ();
 sg13g2_decap_8 FILLER_69_1184 ();
 sg13g2_decap_8 FILLER_69_1191 ();
 sg13g2_decap_8 FILLER_69_1198 ();
 sg13g2_decap_8 FILLER_69_1205 ();
 sg13g2_decap_8 FILLER_69_1212 ();
 sg13g2_decap_8 FILLER_69_1219 ();
 sg13g2_decap_8 FILLER_69_1226 ();
 sg13g2_decap_8 FILLER_69_1233 ();
 sg13g2_decap_8 FILLER_69_1240 ();
 sg13g2_decap_8 FILLER_69_1247 ();
 sg13g2_decap_8 FILLER_69_1254 ();
 sg13g2_decap_8 FILLER_69_1261 ();
 sg13g2_decap_8 FILLER_69_1268 ();
 sg13g2_decap_8 FILLER_69_1275 ();
 sg13g2_decap_8 FILLER_69_1282 ();
 sg13g2_decap_8 FILLER_69_1289 ();
 sg13g2_decap_8 FILLER_69_1296 ();
 sg13g2_decap_8 FILLER_69_1303 ();
 sg13g2_decap_8 FILLER_69_1310 ();
 sg13g2_decap_8 FILLER_69_1317 ();
 sg13g2_decap_8 FILLER_69_1324 ();
 sg13g2_decap_8 FILLER_69_1331 ();
 sg13g2_decap_8 FILLER_69_1338 ();
 sg13g2_decap_8 FILLER_69_1345 ();
 sg13g2_decap_8 FILLER_69_1352 ();
 sg13g2_decap_8 FILLER_69_1359 ();
 sg13g2_decap_8 FILLER_69_1366 ();
 sg13g2_decap_8 FILLER_69_1373 ();
 sg13g2_decap_8 FILLER_69_1380 ();
 sg13g2_decap_8 FILLER_69_1387 ();
 sg13g2_decap_8 FILLER_69_1394 ();
 sg13g2_decap_8 FILLER_69_1401 ();
 sg13g2_decap_8 FILLER_69_1408 ();
 sg13g2_decap_8 FILLER_69_1415 ();
 sg13g2_decap_8 FILLER_69_1422 ();
 sg13g2_decap_8 FILLER_69_1429 ();
 sg13g2_decap_8 FILLER_69_1436 ();
 sg13g2_decap_8 FILLER_69_1443 ();
 sg13g2_decap_8 FILLER_69_1450 ();
 sg13g2_decap_8 FILLER_69_1457 ();
 sg13g2_decap_8 FILLER_69_1464 ();
 sg13g2_decap_8 FILLER_69_1471 ();
 sg13g2_decap_8 FILLER_69_1478 ();
 sg13g2_decap_8 FILLER_69_1485 ();
 sg13g2_decap_8 FILLER_69_1492 ();
 sg13g2_decap_8 FILLER_69_1499 ();
 sg13g2_decap_8 FILLER_69_1506 ();
 sg13g2_decap_8 FILLER_69_1513 ();
 sg13g2_decap_8 FILLER_69_1520 ();
 sg13g2_decap_8 FILLER_69_1527 ();
 sg13g2_decap_8 FILLER_69_1534 ();
 sg13g2_decap_8 FILLER_69_1541 ();
 sg13g2_decap_8 FILLER_69_1548 ();
 sg13g2_decap_8 FILLER_69_1555 ();
 sg13g2_decap_8 FILLER_69_1562 ();
 sg13g2_decap_8 FILLER_69_1569 ();
 sg13g2_decap_8 FILLER_69_1576 ();
 sg13g2_decap_8 FILLER_69_1583 ();
 sg13g2_decap_8 FILLER_69_1590 ();
 sg13g2_decap_8 FILLER_69_1597 ();
 sg13g2_decap_8 FILLER_69_1604 ();
 sg13g2_decap_8 FILLER_69_1611 ();
 sg13g2_decap_8 FILLER_69_1618 ();
 sg13g2_decap_8 FILLER_69_1625 ();
 sg13g2_decap_8 FILLER_69_1632 ();
 sg13g2_decap_8 FILLER_69_1639 ();
 sg13g2_decap_8 FILLER_69_1646 ();
 sg13g2_decap_8 FILLER_69_1653 ();
 sg13g2_decap_8 FILLER_69_1660 ();
 sg13g2_decap_8 FILLER_69_1667 ();
 sg13g2_decap_8 FILLER_69_1674 ();
 sg13g2_decap_8 FILLER_69_1681 ();
 sg13g2_decap_8 FILLER_69_1688 ();
 sg13g2_decap_8 FILLER_69_1695 ();
 sg13g2_decap_8 FILLER_69_1702 ();
 sg13g2_decap_8 FILLER_69_1709 ();
 sg13g2_decap_8 FILLER_69_1716 ();
 sg13g2_decap_8 FILLER_69_1723 ();
 sg13g2_decap_8 FILLER_69_1730 ();
 sg13g2_decap_8 FILLER_69_1737 ();
 sg13g2_decap_8 FILLER_69_1744 ();
 sg13g2_decap_8 FILLER_69_1751 ();
 sg13g2_decap_8 FILLER_69_1758 ();
 sg13g2_fill_2 FILLER_69_1765 ();
 sg13g2_fill_1 FILLER_69_1767 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_decap_8 FILLER_70_14 ();
 sg13g2_decap_8 FILLER_70_21 ();
 sg13g2_decap_8 FILLER_70_28 ();
 sg13g2_fill_2 FILLER_70_61 ();
 sg13g2_fill_1 FILLER_70_63 ();
 sg13g2_fill_2 FILLER_70_90 ();
 sg13g2_fill_1 FILLER_70_92 ();
 sg13g2_decap_4 FILLER_70_120 ();
 sg13g2_fill_1 FILLER_70_124 ();
 sg13g2_fill_2 FILLER_70_137 ();
 sg13g2_decap_8 FILLER_70_151 ();
 sg13g2_decap_8 FILLER_70_158 ();
 sg13g2_decap_8 FILLER_70_165 ();
 sg13g2_fill_2 FILLER_70_172 ();
 sg13g2_fill_1 FILLER_70_174 ();
 sg13g2_fill_2 FILLER_70_216 ();
 sg13g2_fill_1 FILLER_70_218 ();
 sg13g2_fill_2 FILLER_70_235 ();
 sg13g2_fill_1 FILLER_70_237 ();
 sg13g2_decap_8 FILLER_70_242 ();
 sg13g2_decap_8 FILLER_70_249 ();
 sg13g2_decap_4 FILLER_70_256 ();
 sg13g2_fill_1 FILLER_70_260 ();
 sg13g2_decap_8 FILLER_70_269 ();
 sg13g2_fill_2 FILLER_70_320 ();
 sg13g2_fill_1 FILLER_70_322 ();
 sg13g2_fill_2 FILLER_70_334 ();
 sg13g2_fill_2 FILLER_70_341 ();
 sg13g2_decap_8 FILLER_70_364 ();
 sg13g2_fill_2 FILLER_70_387 ();
 sg13g2_fill_2 FILLER_70_399 ();
 sg13g2_fill_1 FILLER_70_401 ();
 sg13g2_decap_8 FILLER_70_421 ();
 sg13g2_decap_4 FILLER_70_428 ();
 sg13g2_fill_2 FILLER_70_432 ();
 sg13g2_fill_2 FILLER_70_442 ();
 sg13g2_fill_2 FILLER_70_465 ();
 sg13g2_decap_8 FILLER_70_475 ();
 sg13g2_decap_8 FILLER_70_482 ();
 sg13g2_fill_2 FILLER_70_489 ();
 sg13g2_fill_2 FILLER_70_495 ();
 sg13g2_decap_4 FILLER_70_505 ();
 sg13g2_fill_1 FILLER_70_509 ();
 sg13g2_fill_2 FILLER_70_516 ();
 sg13g2_fill_2 FILLER_70_522 ();
 sg13g2_fill_1 FILLER_70_524 ();
 sg13g2_decap_4 FILLER_70_530 ();
 sg13g2_fill_1 FILLER_70_534 ();
 sg13g2_fill_2 FILLER_70_561 ();
 sg13g2_fill_1 FILLER_70_586 ();
 sg13g2_fill_1 FILLER_70_617 ();
 sg13g2_decap_8 FILLER_70_623 ();
 sg13g2_decap_4 FILLER_70_630 ();
 sg13g2_fill_1 FILLER_70_634 ();
 sg13g2_fill_2 FILLER_70_647 ();
 sg13g2_fill_1 FILLER_70_649 ();
 sg13g2_fill_1 FILLER_70_659 ();
 sg13g2_fill_2 FILLER_70_676 ();
 sg13g2_decap_8 FILLER_70_686 ();
 sg13g2_decap_8 FILLER_70_699 ();
 sg13g2_fill_1 FILLER_70_706 ();
 sg13g2_decap_8 FILLER_70_711 ();
 sg13g2_fill_2 FILLER_70_728 ();
 sg13g2_decap_4 FILLER_70_740 ();
 sg13g2_fill_2 FILLER_70_744 ();
 sg13g2_fill_2 FILLER_70_772 ();
 sg13g2_fill_1 FILLER_70_774 ();
 sg13g2_fill_1 FILLER_70_793 ();
 sg13g2_decap_8 FILLER_70_799 ();
 sg13g2_fill_1 FILLER_70_806 ();
 sg13g2_decap_8 FILLER_70_840 ();
 sg13g2_decap_8 FILLER_70_861 ();
 sg13g2_decap_4 FILLER_70_868 ();
 sg13g2_fill_1 FILLER_70_872 ();
 sg13g2_fill_1 FILLER_70_896 ();
 sg13g2_fill_2 FILLER_70_902 ();
 sg13g2_fill_2 FILLER_70_930 ();
 sg13g2_fill_1 FILLER_70_932 ();
 sg13g2_fill_2 FILLER_70_942 ();
 sg13g2_fill_1 FILLER_70_944 ();
 sg13g2_fill_2 FILLER_70_964 ();
 sg13g2_fill_2 FILLER_70_989 ();
 sg13g2_decap_4 FILLER_70_1002 ();
 sg13g2_fill_1 FILLER_70_1046 ();
 sg13g2_decap_8 FILLER_70_1082 ();
 sg13g2_decap_8 FILLER_70_1089 ();
 sg13g2_decap_8 FILLER_70_1096 ();
 sg13g2_decap_8 FILLER_70_1103 ();
 sg13g2_decap_8 FILLER_70_1110 ();
 sg13g2_decap_8 FILLER_70_1117 ();
 sg13g2_decap_8 FILLER_70_1124 ();
 sg13g2_decap_8 FILLER_70_1131 ();
 sg13g2_decap_8 FILLER_70_1138 ();
 sg13g2_decap_8 FILLER_70_1145 ();
 sg13g2_decap_8 FILLER_70_1152 ();
 sg13g2_decap_8 FILLER_70_1159 ();
 sg13g2_decap_8 FILLER_70_1166 ();
 sg13g2_decap_8 FILLER_70_1173 ();
 sg13g2_decap_8 FILLER_70_1180 ();
 sg13g2_decap_8 FILLER_70_1187 ();
 sg13g2_decap_8 FILLER_70_1194 ();
 sg13g2_decap_8 FILLER_70_1201 ();
 sg13g2_decap_8 FILLER_70_1208 ();
 sg13g2_decap_8 FILLER_70_1215 ();
 sg13g2_decap_8 FILLER_70_1222 ();
 sg13g2_decap_8 FILLER_70_1229 ();
 sg13g2_decap_8 FILLER_70_1236 ();
 sg13g2_decap_8 FILLER_70_1243 ();
 sg13g2_decap_8 FILLER_70_1250 ();
 sg13g2_decap_8 FILLER_70_1257 ();
 sg13g2_decap_8 FILLER_70_1264 ();
 sg13g2_decap_8 FILLER_70_1271 ();
 sg13g2_decap_8 FILLER_70_1278 ();
 sg13g2_decap_8 FILLER_70_1285 ();
 sg13g2_decap_8 FILLER_70_1292 ();
 sg13g2_decap_8 FILLER_70_1299 ();
 sg13g2_decap_8 FILLER_70_1306 ();
 sg13g2_decap_8 FILLER_70_1313 ();
 sg13g2_decap_8 FILLER_70_1320 ();
 sg13g2_decap_8 FILLER_70_1327 ();
 sg13g2_decap_8 FILLER_70_1334 ();
 sg13g2_decap_8 FILLER_70_1341 ();
 sg13g2_decap_8 FILLER_70_1348 ();
 sg13g2_decap_8 FILLER_70_1355 ();
 sg13g2_decap_8 FILLER_70_1362 ();
 sg13g2_decap_8 FILLER_70_1369 ();
 sg13g2_decap_8 FILLER_70_1376 ();
 sg13g2_decap_8 FILLER_70_1383 ();
 sg13g2_decap_8 FILLER_70_1390 ();
 sg13g2_decap_8 FILLER_70_1397 ();
 sg13g2_decap_8 FILLER_70_1404 ();
 sg13g2_decap_8 FILLER_70_1411 ();
 sg13g2_decap_8 FILLER_70_1418 ();
 sg13g2_decap_8 FILLER_70_1425 ();
 sg13g2_decap_8 FILLER_70_1432 ();
 sg13g2_decap_8 FILLER_70_1439 ();
 sg13g2_decap_8 FILLER_70_1446 ();
 sg13g2_decap_8 FILLER_70_1453 ();
 sg13g2_decap_8 FILLER_70_1460 ();
 sg13g2_decap_8 FILLER_70_1467 ();
 sg13g2_decap_8 FILLER_70_1474 ();
 sg13g2_decap_8 FILLER_70_1481 ();
 sg13g2_decap_8 FILLER_70_1488 ();
 sg13g2_decap_8 FILLER_70_1495 ();
 sg13g2_decap_8 FILLER_70_1502 ();
 sg13g2_decap_8 FILLER_70_1509 ();
 sg13g2_decap_8 FILLER_70_1516 ();
 sg13g2_decap_8 FILLER_70_1523 ();
 sg13g2_decap_8 FILLER_70_1530 ();
 sg13g2_decap_8 FILLER_70_1537 ();
 sg13g2_decap_8 FILLER_70_1544 ();
 sg13g2_decap_8 FILLER_70_1551 ();
 sg13g2_decap_8 FILLER_70_1558 ();
 sg13g2_decap_8 FILLER_70_1565 ();
 sg13g2_decap_8 FILLER_70_1572 ();
 sg13g2_decap_8 FILLER_70_1579 ();
 sg13g2_decap_8 FILLER_70_1586 ();
 sg13g2_decap_8 FILLER_70_1593 ();
 sg13g2_decap_8 FILLER_70_1600 ();
 sg13g2_decap_8 FILLER_70_1607 ();
 sg13g2_decap_8 FILLER_70_1614 ();
 sg13g2_decap_8 FILLER_70_1621 ();
 sg13g2_decap_8 FILLER_70_1628 ();
 sg13g2_decap_8 FILLER_70_1635 ();
 sg13g2_decap_8 FILLER_70_1642 ();
 sg13g2_decap_8 FILLER_70_1649 ();
 sg13g2_decap_8 FILLER_70_1656 ();
 sg13g2_decap_8 FILLER_70_1663 ();
 sg13g2_decap_8 FILLER_70_1670 ();
 sg13g2_decap_8 FILLER_70_1677 ();
 sg13g2_decap_8 FILLER_70_1684 ();
 sg13g2_decap_8 FILLER_70_1691 ();
 sg13g2_decap_8 FILLER_70_1698 ();
 sg13g2_decap_8 FILLER_70_1705 ();
 sg13g2_decap_8 FILLER_70_1712 ();
 sg13g2_decap_8 FILLER_70_1719 ();
 sg13g2_decap_8 FILLER_70_1726 ();
 sg13g2_decap_8 FILLER_70_1733 ();
 sg13g2_decap_8 FILLER_70_1740 ();
 sg13g2_decap_8 FILLER_70_1747 ();
 sg13g2_decap_8 FILLER_70_1754 ();
 sg13g2_decap_8 FILLER_70_1761 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_decap_8 FILLER_71_7 ();
 sg13g2_decap_8 FILLER_71_14 ();
 sg13g2_decap_8 FILLER_71_21 ();
 sg13g2_decap_4 FILLER_71_28 ();
 sg13g2_fill_2 FILLER_71_32 ();
 sg13g2_fill_1 FILLER_71_60 ();
 sg13g2_fill_2 FILLER_71_69 ();
 sg13g2_fill_1 FILLER_71_75 ();
 sg13g2_decap_8 FILLER_71_81 ();
 sg13g2_decap_8 FILLER_71_88 ();
 sg13g2_fill_1 FILLER_71_95 ();
 sg13g2_fill_2 FILLER_71_109 ();
 sg13g2_decap_8 FILLER_71_116 ();
 sg13g2_fill_2 FILLER_71_123 ();
 sg13g2_decap_4 FILLER_71_145 ();
 sg13g2_fill_2 FILLER_71_149 ();
 sg13g2_fill_1 FILLER_71_164 ();
 sg13g2_fill_2 FILLER_71_198 ();
 sg13g2_fill_2 FILLER_71_217 ();
 sg13g2_fill_1 FILLER_71_219 ();
 sg13g2_fill_2 FILLER_71_226 ();
 sg13g2_fill_1 FILLER_71_228 ();
 sg13g2_fill_1 FILLER_71_245 ();
 sg13g2_fill_1 FILLER_71_256 ();
 sg13g2_decap_4 FILLER_71_282 ();
 sg13g2_fill_1 FILLER_71_286 ();
 sg13g2_fill_2 FILLER_71_329 ();
 sg13g2_decap_8 FILLER_71_340 ();
 sg13g2_decap_4 FILLER_71_374 ();
 sg13g2_fill_1 FILLER_71_378 ();
 sg13g2_decap_8 FILLER_71_394 ();
 sg13g2_decap_8 FILLER_71_401 ();
 sg13g2_decap_4 FILLER_71_408 ();
 sg13g2_fill_1 FILLER_71_412 ();
 sg13g2_fill_2 FILLER_71_434 ();
 sg13g2_fill_2 FILLER_71_466 ();
 sg13g2_decap_8 FILLER_71_486 ();
 sg13g2_fill_1 FILLER_71_520 ();
 sg13g2_decap_8 FILLER_71_526 ();
 sg13g2_fill_1 FILLER_71_533 ();
 sg13g2_decap_8 FILLER_71_549 ();
 sg13g2_decap_8 FILLER_71_556 ();
 sg13g2_fill_1 FILLER_71_563 ();
 sg13g2_decap_8 FILLER_71_577 ();
 sg13g2_decap_8 FILLER_71_584 ();
 sg13g2_decap_4 FILLER_71_591 ();
 sg13g2_fill_1 FILLER_71_595 ();
 sg13g2_fill_1 FILLER_71_601 ();
 sg13g2_fill_1 FILLER_71_606 ();
 sg13g2_decap_4 FILLER_71_618 ();
 sg13g2_fill_2 FILLER_71_622 ();
 sg13g2_decap_4 FILLER_71_640 ();
 sg13g2_fill_2 FILLER_71_644 ();
 sg13g2_fill_1 FILLER_71_664 ();
 sg13g2_decap_4 FILLER_71_681 ();
 sg13g2_fill_1 FILLER_71_699 ();
 sg13g2_fill_2 FILLER_71_750 ();
 sg13g2_fill_1 FILLER_71_752 ();
 sg13g2_decap_8 FILLER_71_767 ();
 sg13g2_decap_4 FILLER_71_774 ();
 sg13g2_fill_2 FILLER_71_778 ();
 sg13g2_fill_2 FILLER_71_794 ();
 sg13g2_fill_1 FILLER_71_804 ();
 sg13g2_decap_4 FILLER_71_819 ();
 sg13g2_fill_2 FILLER_71_823 ();
 sg13g2_fill_2 FILLER_71_894 ();
 sg13g2_fill_1 FILLER_71_896 ();
 sg13g2_decap_8 FILLER_71_912 ();
 sg13g2_fill_1 FILLER_71_927 ();
 sg13g2_fill_1 FILLER_71_959 ();
 sg13g2_fill_2 FILLER_71_974 ();
 sg13g2_fill_1 FILLER_71_976 ();
 sg13g2_fill_2 FILLER_71_1020 ();
 sg13g2_fill_1 FILLER_71_1022 ();
 sg13g2_decap_8 FILLER_71_1026 ();
 sg13g2_fill_2 FILLER_71_1033 ();
 sg13g2_fill_2 FILLER_71_1044 ();
 sg13g2_decap_8 FILLER_71_1056 ();
 sg13g2_decap_8 FILLER_71_1063 ();
 sg13g2_decap_8 FILLER_71_1070 ();
 sg13g2_decap_8 FILLER_71_1077 ();
 sg13g2_decap_8 FILLER_71_1084 ();
 sg13g2_decap_8 FILLER_71_1091 ();
 sg13g2_decap_8 FILLER_71_1098 ();
 sg13g2_decap_8 FILLER_71_1105 ();
 sg13g2_decap_8 FILLER_71_1112 ();
 sg13g2_decap_8 FILLER_71_1119 ();
 sg13g2_decap_8 FILLER_71_1126 ();
 sg13g2_decap_8 FILLER_71_1133 ();
 sg13g2_decap_8 FILLER_71_1140 ();
 sg13g2_decap_8 FILLER_71_1147 ();
 sg13g2_decap_8 FILLER_71_1154 ();
 sg13g2_decap_8 FILLER_71_1161 ();
 sg13g2_decap_8 FILLER_71_1168 ();
 sg13g2_decap_8 FILLER_71_1175 ();
 sg13g2_decap_8 FILLER_71_1182 ();
 sg13g2_decap_8 FILLER_71_1189 ();
 sg13g2_decap_8 FILLER_71_1196 ();
 sg13g2_decap_8 FILLER_71_1203 ();
 sg13g2_decap_8 FILLER_71_1210 ();
 sg13g2_decap_8 FILLER_71_1217 ();
 sg13g2_decap_8 FILLER_71_1224 ();
 sg13g2_decap_8 FILLER_71_1231 ();
 sg13g2_decap_8 FILLER_71_1238 ();
 sg13g2_decap_8 FILLER_71_1245 ();
 sg13g2_decap_8 FILLER_71_1252 ();
 sg13g2_decap_8 FILLER_71_1259 ();
 sg13g2_decap_8 FILLER_71_1266 ();
 sg13g2_decap_8 FILLER_71_1273 ();
 sg13g2_decap_8 FILLER_71_1280 ();
 sg13g2_decap_8 FILLER_71_1287 ();
 sg13g2_decap_8 FILLER_71_1294 ();
 sg13g2_decap_8 FILLER_71_1301 ();
 sg13g2_decap_8 FILLER_71_1308 ();
 sg13g2_decap_8 FILLER_71_1315 ();
 sg13g2_decap_8 FILLER_71_1322 ();
 sg13g2_decap_8 FILLER_71_1329 ();
 sg13g2_decap_8 FILLER_71_1336 ();
 sg13g2_decap_8 FILLER_71_1343 ();
 sg13g2_decap_8 FILLER_71_1350 ();
 sg13g2_decap_8 FILLER_71_1357 ();
 sg13g2_decap_8 FILLER_71_1364 ();
 sg13g2_decap_8 FILLER_71_1371 ();
 sg13g2_decap_8 FILLER_71_1378 ();
 sg13g2_decap_8 FILLER_71_1385 ();
 sg13g2_decap_8 FILLER_71_1392 ();
 sg13g2_decap_8 FILLER_71_1399 ();
 sg13g2_decap_8 FILLER_71_1406 ();
 sg13g2_decap_8 FILLER_71_1413 ();
 sg13g2_decap_8 FILLER_71_1420 ();
 sg13g2_decap_8 FILLER_71_1427 ();
 sg13g2_decap_8 FILLER_71_1434 ();
 sg13g2_decap_8 FILLER_71_1441 ();
 sg13g2_decap_8 FILLER_71_1448 ();
 sg13g2_decap_8 FILLER_71_1455 ();
 sg13g2_decap_8 FILLER_71_1462 ();
 sg13g2_decap_8 FILLER_71_1469 ();
 sg13g2_decap_8 FILLER_71_1476 ();
 sg13g2_decap_8 FILLER_71_1483 ();
 sg13g2_decap_8 FILLER_71_1490 ();
 sg13g2_decap_8 FILLER_71_1497 ();
 sg13g2_decap_8 FILLER_71_1504 ();
 sg13g2_decap_8 FILLER_71_1511 ();
 sg13g2_decap_8 FILLER_71_1518 ();
 sg13g2_decap_8 FILLER_71_1525 ();
 sg13g2_decap_8 FILLER_71_1532 ();
 sg13g2_decap_8 FILLER_71_1539 ();
 sg13g2_decap_8 FILLER_71_1546 ();
 sg13g2_decap_8 FILLER_71_1553 ();
 sg13g2_decap_8 FILLER_71_1560 ();
 sg13g2_decap_8 FILLER_71_1567 ();
 sg13g2_decap_8 FILLER_71_1574 ();
 sg13g2_decap_8 FILLER_71_1581 ();
 sg13g2_decap_8 FILLER_71_1588 ();
 sg13g2_decap_8 FILLER_71_1595 ();
 sg13g2_decap_8 FILLER_71_1602 ();
 sg13g2_decap_8 FILLER_71_1609 ();
 sg13g2_decap_8 FILLER_71_1616 ();
 sg13g2_decap_8 FILLER_71_1623 ();
 sg13g2_decap_8 FILLER_71_1630 ();
 sg13g2_decap_8 FILLER_71_1637 ();
 sg13g2_decap_8 FILLER_71_1644 ();
 sg13g2_decap_8 FILLER_71_1651 ();
 sg13g2_decap_8 FILLER_71_1658 ();
 sg13g2_decap_8 FILLER_71_1665 ();
 sg13g2_decap_8 FILLER_71_1672 ();
 sg13g2_decap_8 FILLER_71_1679 ();
 sg13g2_decap_8 FILLER_71_1686 ();
 sg13g2_decap_8 FILLER_71_1693 ();
 sg13g2_decap_8 FILLER_71_1700 ();
 sg13g2_decap_8 FILLER_71_1707 ();
 sg13g2_decap_8 FILLER_71_1714 ();
 sg13g2_decap_8 FILLER_71_1721 ();
 sg13g2_decap_8 FILLER_71_1728 ();
 sg13g2_decap_8 FILLER_71_1735 ();
 sg13g2_decap_8 FILLER_71_1742 ();
 sg13g2_decap_8 FILLER_71_1749 ();
 sg13g2_decap_8 FILLER_71_1756 ();
 sg13g2_decap_4 FILLER_71_1763 ();
 sg13g2_fill_1 FILLER_71_1767 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_decap_8 FILLER_72_14 ();
 sg13g2_decap_8 FILLER_72_21 ();
 sg13g2_decap_8 FILLER_72_28 ();
 sg13g2_decap_8 FILLER_72_35 ();
 sg13g2_decap_4 FILLER_72_42 ();
 sg13g2_fill_2 FILLER_72_46 ();
 sg13g2_fill_2 FILLER_72_57 ();
 sg13g2_fill_1 FILLER_72_59 ();
 sg13g2_fill_1 FILLER_72_76 ();
 sg13g2_fill_2 FILLER_72_82 ();
 sg13g2_fill_1 FILLER_72_84 ();
 sg13g2_fill_2 FILLER_72_107 ();
 sg13g2_decap_4 FILLER_72_114 ();
 sg13g2_fill_2 FILLER_72_118 ();
 sg13g2_fill_2 FILLER_72_132 ();
 sg13g2_fill_2 FILLER_72_146 ();
 sg13g2_decap_4 FILLER_72_174 ();
 sg13g2_fill_2 FILLER_72_190 ();
 sg13g2_fill_1 FILLER_72_192 ();
 sg13g2_fill_1 FILLER_72_246 ();
 sg13g2_decap_4 FILLER_72_255 ();
 sg13g2_fill_2 FILLER_72_272 ();
 sg13g2_fill_2 FILLER_72_287 ();
 sg13g2_fill_1 FILLER_72_289 ();
 sg13g2_fill_2 FILLER_72_296 ();
 sg13g2_fill_1 FILLER_72_298 ();
 sg13g2_fill_1 FILLER_72_312 ();
 sg13g2_fill_2 FILLER_72_347 ();
 sg13g2_fill_1 FILLER_72_349 ();
 sg13g2_fill_2 FILLER_72_358 ();
 sg13g2_fill_1 FILLER_72_417 ();
 sg13g2_decap_8 FILLER_72_433 ();
 sg13g2_fill_2 FILLER_72_440 ();
 sg13g2_decap_8 FILLER_72_455 ();
 sg13g2_fill_1 FILLER_72_462 ();
 sg13g2_fill_1 FILLER_72_481 ();
 sg13g2_fill_1 FILLER_72_498 ();
 sg13g2_fill_2 FILLER_72_504 ();
 sg13g2_fill_1 FILLER_72_506 ();
 sg13g2_decap_4 FILLER_72_537 ();
 sg13g2_fill_2 FILLER_72_546 ();
 sg13g2_fill_1 FILLER_72_552 ();
 sg13g2_decap_8 FILLER_72_557 ();
 sg13g2_fill_2 FILLER_72_564 ();
 sg13g2_fill_1 FILLER_72_566 ();
 sg13g2_fill_2 FILLER_72_577 ();
 sg13g2_fill_1 FILLER_72_579 ();
 sg13g2_fill_1 FILLER_72_588 ();
 sg13g2_fill_1 FILLER_72_611 ();
 sg13g2_fill_2 FILLER_72_644 ();
 sg13g2_decap_8 FILLER_72_684 ();
 sg13g2_fill_2 FILLER_72_691 ();
 sg13g2_decap_4 FILLER_72_698 ();
 sg13g2_decap_4 FILLER_72_714 ();
 sg13g2_fill_2 FILLER_72_718 ();
 sg13g2_decap_8 FILLER_72_732 ();
 sg13g2_fill_1 FILLER_72_739 ();
 sg13g2_fill_1 FILLER_72_743 ();
 sg13g2_decap_4 FILLER_72_778 ();
 sg13g2_fill_1 FILLER_72_798 ();
 sg13g2_fill_2 FILLER_72_820 ();
 sg13g2_fill_1 FILLER_72_822 ();
 sg13g2_fill_1 FILLER_72_845 ();
 sg13g2_decap_4 FILLER_72_863 ();
 sg13g2_fill_1 FILLER_72_867 ();
 sg13g2_decap_4 FILLER_72_873 ();
 sg13g2_fill_1 FILLER_72_877 ();
 sg13g2_fill_1 FILLER_72_895 ();
 sg13g2_decap_8 FILLER_72_922 ();
 sg13g2_decap_4 FILLER_72_929 ();
 sg13g2_fill_2 FILLER_72_933 ();
 sg13g2_fill_2 FILLER_72_957 ();
 sg13g2_decap_8 FILLER_72_962 ();
 sg13g2_fill_2 FILLER_72_969 ();
 sg13g2_fill_1 FILLER_72_971 ();
 sg13g2_decap_4 FILLER_72_982 ();
 sg13g2_fill_1 FILLER_72_986 ();
 sg13g2_fill_2 FILLER_72_991 ();
 sg13g2_decap_4 FILLER_72_1001 ();
 sg13g2_decap_8 FILLER_72_1013 ();
 sg13g2_decap_8 FILLER_72_1020 ();
 sg13g2_decap_8 FILLER_72_1027 ();
 sg13g2_decap_8 FILLER_72_1034 ();
 sg13g2_decap_8 FILLER_72_1041 ();
 sg13g2_decap_8 FILLER_72_1048 ();
 sg13g2_decap_8 FILLER_72_1055 ();
 sg13g2_decap_8 FILLER_72_1062 ();
 sg13g2_decap_8 FILLER_72_1069 ();
 sg13g2_decap_8 FILLER_72_1076 ();
 sg13g2_decap_8 FILLER_72_1083 ();
 sg13g2_decap_8 FILLER_72_1090 ();
 sg13g2_decap_8 FILLER_72_1097 ();
 sg13g2_decap_8 FILLER_72_1104 ();
 sg13g2_decap_8 FILLER_72_1111 ();
 sg13g2_decap_8 FILLER_72_1118 ();
 sg13g2_decap_8 FILLER_72_1125 ();
 sg13g2_decap_8 FILLER_72_1132 ();
 sg13g2_decap_8 FILLER_72_1139 ();
 sg13g2_decap_8 FILLER_72_1146 ();
 sg13g2_decap_8 FILLER_72_1153 ();
 sg13g2_decap_8 FILLER_72_1160 ();
 sg13g2_decap_8 FILLER_72_1167 ();
 sg13g2_decap_8 FILLER_72_1174 ();
 sg13g2_decap_8 FILLER_72_1181 ();
 sg13g2_decap_8 FILLER_72_1188 ();
 sg13g2_decap_8 FILLER_72_1195 ();
 sg13g2_decap_8 FILLER_72_1202 ();
 sg13g2_decap_8 FILLER_72_1209 ();
 sg13g2_decap_8 FILLER_72_1216 ();
 sg13g2_decap_8 FILLER_72_1223 ();
 sg13g2_decap_8 FILLER_72_1230 ();
 sg13g2_decap_8 FILLER_72_1237 ();
 sg13g2_decap_8 FILLER_72_1244 ();
 sg13g2_decap_8 FILLER_72_1251 ();
 sg13g2_decap_8 FILLER_72_1258 ();
 sg13g2_decap_8 FILLER_72_1265 ();
 sg13g2_decap_8 FILLER_72_1272 ();
 sg13g2_decap_8 FILLER_72_1279 ();
 sg13g2_decap_8 FILLER_72_1286 ();
 sg13g2_decap_8 FILLER_72_1293 ();
 sg13g2_decap_8 FILLER_72_1300 ();
 sg13g2_decap_8 FILLER_72_1307 ();
 sg13g2_decap_8 FILLER_72_1314 ();
 sg13g2_decap_8 FILLER_72_1321 ();
 sg13g2_decap_8 FILLER_72_1328 ();
 sg13g2_decap_8 FILLER_72_1335 ();
 sg13g2_decap_8 FILLER_72_1342 ();
 sg13g2_decap_8 FILLER_72_1349 ();
 sg13g2_decap_8 FILLER_72_1356 ();
 sg13g2_decap_8 FILLER_72_1363 ();
 sg13g2_decap_8 FILLER_72_1370 ();
 sg13g2_decap_8 FILLER_72_1377 ();
 sg13g2_decap_8 FILLER_72_1384 ();
 sg13g2_decap_8 FILLER_72_1391 ();
 sg13g2_decap_8 FILLER_72_1398 ();
 sg13g2_decap_8 FILLER_72_1405 ();
 sg13g2_decap_8 FILLER_72_1412 ();
 sg13g2_decap_8 FILLER_72_1419 ();
 sg13g2_decap_8 FILLER_72_1426 ();
 sg13g2_decap_8 FILLER_72_1433 ();
 sg13g2_decap_8 FILLER_72_1440 ();
 sg13g2_decap_8 FILLER_72_1447 ();
 sg13g2_decap_8 FILLER_72_1454 ();
 sg13g2_decap_8 FILLER_72_1461 ();
 sg13g2_decap_8 FILLER_72_1468 ();
 sg13g2_decap_8 FILLER_72_1475 ();
 sg13g2_decap_8 FILLER_72_1482 ();
 sg13g2_decap_8 FILLER_72_1489 ();
 sg13g2_decap_8 FILLER_72_1496 ();
 sg13g2_decap_8 FILLER_72_1503 ();
 sg13g2_decap_8 FILLER_72_1510 ();
 sg13g2_decap_8 FILLER_72_1517 ();
 sg13g2_decap_8 FILLER_72_1524 ();
 sg13g2_decap_8 FILLER_72_1531 ();
 sg13g2_decap_8 FILLER_72_1538 ();
 sg13g2_decap_8 FILLER_72_1545 ();
 sg13g2_decap_8 FILLER_72_1552 ();
 sg13g2_decap_8 FILLER_72_1559 ();
 sg13g2_decap_8 FILLER_72_1566 ();
 sg13g2_decap_8 FILLER_72_1573 ();
 sg13g2_decap_8 FILLER_72_1580 ();
 sg13g2_decap_8 FILLER_72_1587 ();
 sg13g2_decap_8 FILLER_72_1594 ();
 sg13g2_decap_8 FILLER_72_1601 ();
 sg13g2_decap_8 FILLER_72_1608 ();
 sg13g2_decap_8 FILLER_72_1615 ();
 sg13g2_decap_8 FILLER_72_1622 ();
 sg13g2_decap_8 FILLER_72_1629 ();
 sg13g2_decap_8 FILLER_72_1636 ();
 sg13g2_decap_8 FILLER_72_1643 ();
 sg13g2_decap_8 FILLER_72_1650 ();
 sg13g2_decap_8 FILLER_72_1657 ();
 sg13g2_decap_8 FILLER_72_1664 ();
 sg13g2_decap_8 FILLER_72_1671 ();
 sg13g2_decap_8 FILLER_72_1678 ();
 sg13g2_decap_8 FILLER_72_1685 ();
 sg13g2_decap_8 FILLER_72_1692 ();
 sg13g2_decap_8 FILLER_72_1699 ();
 sg13g2_decap_8 FILLER_72_1706 ();
 sg13g2_decap_8 FILLER_72_1713 ();
 sg13g2_decap_8 FILLER_72_1720 ();
 sg13g2_decap_8 FILLER_72_1727 ();
 sg13g2_decap_8 FILLER_72_1734 ();
 sg13g2_decap_8 FILLER_72_1741 ();
 sg13g2_decap_8 FILLER_72_1748 ();
 sg13g2_decap_8 FILLER_72_1755 ();
 sg13g2_decap_4 FILLER_72_1762 ();
 sg13g2_fill_2 FILLER_72_1766 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_decap_8 FILLER_73_14 ();
 sg13g2_decap_8 FILLER_73_21 ();
 sg13g2_fill_2 FILLER_73_28 ();
 sg13g2_fill_1 FILLER_73_30 ();
 sg13g2_fill_2 FILLER_73_65 ();
 sg13g2_fill_1 FILLER_73_67 ();
 sg13g2_fill_1 FILLER_73_85 ();
 sg13g2_fill_2 FILLER_73_97 ();
 sg13g2_decap_8 FILLER_73_115 ();
 sg13g2_decap_4 FILLER_73_122 ();
 sg13g2_fill_2 FILLER_73_139 ();
 sg13g2_fill_1 FILLER_73_141 ();
 sg13g2_fill_1 FILLER_73_159 ();
 sg13g2_decap_8 FILLER_73_168 ();
 sg13g2_decap_8 FILLER_73_175 ();
 sg13g2_fill_1 FILLER_73_182 ();
 sg13g2_fill_1 FILLER_73_213 ();
 sg13g2_decap_4 FILLER_73_219 ();
 sg13g2_fill_1 FILLER_73_223 ();
 sg13g2_fill_1 FILLER_73_242 ();
 sg13g2_fill_1 FILLER_73_249 ();
 sg13g2_decap_8 FILLER_73_264 ();
 sg13g2_fill_2 FILLER_73_291 ();
 sg13g2_fill_1 FILLER_73_293 ();
 sg13g2_fill_2 FILLER_73_299 ();
 sg13g2_fill_1 FILLER_73_301 ();
 sg13g2_decap_8 FILLER_73_346 ();
 sg13g2_fill_2 FILLER_73_353 ();
 sg13g2_fill_1 FILLER_73_355 ();
 sg13g2_fill_1 FILLER_73_382 ();
 sg13g2_decap_8 FILLER_73_387 ();
 sg13g2_decap_8 FILLER_73_394 ();
 sg13g2_fill_2 FILLER_73_401 ();
 sg13g2_fill_1 FILLER_73_403 ();
 sg13g2_fill_2 FILLER_73_413 ();
 sg13g2_fill_1 FILLER_73_415 ();
 sg13g2_fill_1 FILLER_73_434 ();
 sg13g2_decap_8 FILLER_73_450 ();
 sg13g2_fill_2 FILLER_73_457 ();
 sg13g2_fill_1 FILLER_73_459 ();
 sg13g2_decap_8 FILLER_73_481 ();
 sg13g2_fill_1 FILLER_73_493 ();
 sg13g2_fill_2 FILLER_73_507 ();
 sg13g2_decap_4 FILLER_73_517 ();
 sg13g2_fill_1 FILLER_73_521 ();
 sg13g2_decap_4 FILLER_73_546 ();
 sg13g2_decap_8 FILLER_73_568 ();
 sg13g2_decap_4 FILLER_73_575 ();
 sg13g2_fill_2 FILLER_73_579 ();
 sg13g2_decap_8 FILLER_73_589 ();
 sg13g2_fill_1 FILLER_73_596 ();
 sg13g2_fill_2 FILLER_73_616 ();
 sg13g2_fill_1 FILLER_73_618 ();
 sg13g2_decap_8 FILLER_73_628 ();
 sg13g2_fill_2 FILLER_73_635 ();
 sg13g2_decap_8 FILLER_73_641 ();
 sg13g2_fill_1 FILLER_73_648 ();
 sg13g2_decap_4 FILLER_73_657 ();
 sg13g2_fill_2 FILLER_73_667 ();
 sg13g2_fill_1 FILLER_73_669 ();
 sg13g2_decap_4 FILLER_73_690 ();
 sg13g2_fill_1 FILLER_73_694 ();
 sg13g2_decap_4 FILLER_73_730 ();
 sg13g2_fill_1 FILLER_73_734 ();
 sg13g2_fill_2 FILLER_73_751 ();
 sg13g2_fill_1 FILLER_73_753 ();
 sg13g2_decap_8 FILLER_73_768 ();
 sg13g2_decap_4 FILLER_73_775 ();
 sg13g2_fill_2 FILLER_73_779 ();
 sg13g2_fill_2 FILLER_73_788 ();
 sg13g2_fill_1 FILLER_73_790 ();
 sg13g2_fill_1 FILLER_73_804 ();
 sg13g2_decap_4 FILLER_73_813 ();
 sg13g2_fill_2 FILLER_73_830 ();
 sg13g2_fill_1 FILLER_73_849 ();
 sg13g2_decap_4 FILLER_73_921 ();
 sg13g2_fill_2 FILLER_73_938 ();
 sg13g2_fill_1 FILLER_73_948 ();
 sg13g2_fill_2 FILLER_73_984 ();
 sg13g2_fill_1 FILLER_73_1003 ();
 sg13g2_decap_8 FILLER_73_1035 ();
 sg13g2_decap_8 FILLER_73_1042 ();
 sg13g2_decap_8 FILLER_73_1049 ();
 sg13g2_decap_8 FILLER_73_1056 ();
 sg13g2_decap_8 FILLER_73_1063 ();
 sg13g2_decap_8 FILLER_73_1070 ();
 sg13g2_decap_8 FILLER_73_1077 ();
 sg13g2_decap_8 FILLER_73_1084 ();
 sg13g2_decap_8 FILLER_73_1091 ();
 sg13g2_decap_8 FILLER_73_1098 ();
 sg13g2_decap_8 FILLER_73_1105 ();
 sg13g2_decap_8 FILLER_73_1112 ();
 sg13g2_decap_8 FILLER_73_1119 ();
 sg13g2_decap_8 FILLER_73_1126 ();
 sg13g2_decap_8 FILLER_73_1133 ();
 sg13g2_decap_8 FILLER_73_1140 ();
 sg13g2_decap_8 FILLER_73_1147 ();
 sg13g2_decap_8 FILLER_73_1154 ();
 sg13g2_decap_8 FILLER_73_1161 ();
 sg13g2_decap_8 FILLER_73_1168 ();
 sg13g2_decap_8 FILLER_73_1175 ();
 sg13g2_decap_8 FILLER_73_1182 ();
 sg13g2_decap_8 FILLER_73_1189 ();
 sg13g2_decap_8 FILLER_73_1196 ();
 sg13g2_decap_8 FILLER_73_1203 ();
 sg13g2_decap_8 FILLER_73_1210 ();
 sg13g2_decap_8 FILLER_73_1217 ();
 sg13g2_decap_8 FILLER_73_1224 ();
 sg13g2_decap_8 FILLER_73_1231 ();
 sg13g2_decap_8 FILLER_73_1238 ();
 sg13g2_decap_8 FILLER_73_1245 ();
 sg13g2_decap_8 FILLER_73_1252 ();
 sg13g2_decap_8 FILLER_73_1259 ();
 sg13g2_decap_8 FILLER_73_1266 ();
 sg13g2_decap_8 FILLER_73_1273 ();
 sg13g2_decap_8 FILLER_73_1280 ();
 sg13g2_decap_8 FILLER_73_1287 ();
 sg13g2_decap_8 FILLER_73_1294 ();
 sg13g2_decap_8 FILLER_73_1301 ();
 sg13g2_decap_8 FILLER_73_1308 ();
 sg13g2_decap_8 FILLER_73_1315 ();
 sg13g2_decap_8 FILLER_73_1322 ();
 sg13g2_decap_8 FILLER_73_1329 ();
 sg13g2_decap_8 FILLER_73_1336 ();
 sg13g2_decap_8 FILLER_73_1343 ();
 sg13g2_decap_8 FILLER_73_1350 ();
 sg13g2_decap_8 FILLER_73_1357 ();
 sg13g2_decap_8 FILLER_73_1364 ();
 sg13g2_decap_8 FILLER_73_1371 ();
 sg13g2_decap_8 FILLER_73_1378 ();
 sg13g2_decap_8 FILLER_73_1385 ();
 sg13g2_decap_8 FILLER_73_1392 ();
 sg13g2_decap_8 FILLER_73_1399 ();
 sg13g2_decap_8 FILLER_73_1406 ();
 sg13g2_decap_8 FILLER_73_1413 ();
 sg13g2_decap_8 FILLER_73_1420 ();
 sg13g2_decap_8 FILLER_73_1427 ();
 sg13g2_decap_8 FILLER_73_1434 ();
 sg13g2_decap_8 FILLER_73_1441 ();
 sg13g2_decap_8 FILLER_73_1448 ();
 sg13g2_decap_8 FILLER_73_1455 ();
 sg13g2_decap_8 FILLER_73_1462 ();
 sg13g2_decap_8 FILLER_73_1469 ();
 sg13g2_decap_8 FILLER_73_1476 ();
 sg13g2_decap_8 FILLER_73_1483 ();
 sg13g2_decap_8 FILLER_73_1490 ();
 sg13g2_decap_8 FILLER_73_1497 ();
 sg13g2_decap_8 FILLER_73_1504 ();
 sg13g2_decap_8 FILLER_73_1511 ();
 sg13g2_decap_8 FILLER_73_1518 ();
 sg13g2_decap_8 FILLER_73_1525 ();
 sg13g2_decap_8 FILLER_73_1532 ();
 sg13g2_decap_8 FILLER_73_1539 ();
 sg13g2_decap_8 FILLER_73_1546 ();
 sg13g2_decap_8 FILLER_73_1553 ();
 sg13g2_decap_8 FILLER_73_1560 ();
 sg13g2_decap_8 FILLER_73_1567 ();
 sg13g2_decap_8 FILLER_73_1574 ();
 sg13g2_decap_8 FILLER_73_1581 ();
 sg13g2_decap_8 FILLER_73_1588 ();
 sg13g2_decap_8 FILLER_73_1595 ();
 sg13g2_decap_8 FILLER_73_1602 ();
 sg13g2_decap_8 FILLER_73_1609 ();
 sg13g2_decap_8 FILLER_73_1616 ();
 sg13g2_decap_8 FILLER_73_1623 ();
 sg13g2_decap_8 FILLER_73_1630 ();
 sg13g2_decap_8 FILLER_73_1637 ();
 sg13g2_decap_8 FILLER_73_1644 ();
 sg13g2_decap_8 FILLER_73_1651 ();
 sg13g2_decap_8 FILLER_73_1658 ();
 sg13g2_decap_8 FILLER_73_1665 ();
 sg13g2_decap_8 FILLER_73_1672 ();
 sg13g2_decap_8 FILLER_73_1679 ();
 sg13g2_decap_8 FILLER_73_1686 ();
 sg13g2_decap_8 FILLER_73_1693 ();
 sg13g2_decap_8 FILLER_73_1700 ();
 sg13g2_decap_8 FILLER_73_1707 ();
 sg13g2_decap_8 FILLER_73_1714 ();
 sg13g2_decap_8 FILLER_73_1721 ();
 sg13g2_decap_8 FILLER_73_1728 ();
 sg13g2_decap_8 FILLER_73_1735 ();
 sg13g2_decap_8 FILLER_73_1742 ();
 sg13g2_decap_8 FILLER_73_1749 ();
 sg13g2_decap_8 FILLER_73_1756 ();
 sg13g2_decap_4 FILLER_73_1763 ();
 sg13g2_fill_1 FILLER_73_1767 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_decap_8 FILLER_74_14 ();
 sg13g2_decap_8 FILLER_74_21 ();
 sg13g2_decap_8 FILLER_74_28 ();
 sg13g2_decap_8 FILLER_74_35 ();
 sg13g2_decap_4 FILLER_74_42 ();
 sg13g2_fill_2 FILLER_74_46 ();
 sg13g2_fill_2 FILLER_74_70 ();
 sg13g2_fill_2 FILLER_74_101 ();
 sg13g2_fill_1 FILLER_74_103 ();
 sg13g2_fill_2 FILLER_74_121 ();
 sg13g2_fill_1 FILLER_74_146 ();
 sg13g2_decap_4 FILLER_74_171 ();
 sg13g2_fill_1 FILLER_74_191 ();
 sg13g2_fill_2 FILLER_74_209 ();
 sg13g2_fill_1 FILLER_74_211 ();
 sg13g2_decap_4 FILLER_74_229 ();
 sg13g2_fill_2 FILLER_74_357 ();
 sg13g2_fill_2 FILLER_74_371 ();
 sg13g2_fill_2 FILLER_74_387 ();
 sg13g2_fill_1 FILLER_74_389 ();
 sg13g2_fill_1 FILLER_74_436 ();
 sg13g2_fill_2 FILLER_74_450 ();
 sg13g2_fill_1 FILLER_74_452 ();
 sg13g2_decap_8 FILLER_74_477 ();
 sg13g2_decap_8 FILLER_74_484 ();
 sg13g2_fill_1 FILLER_74_491 ();
 sg13g2_decap_4 FILLER_74_505 ();
 sg13g2_decap_8 FILLER_74_517 ();
 sg13g2_fill_2 FILLER_74_552 ();
 sg13g2_decap_4 FILLER_74_578 ();
 sg13g2_decap_8 FILLER_74_587 ();
 sg13g2_decap_4 FILLER_74_594 ();
 sg13g2_fill_2 FILLER_74_603 ();
 sg13g2_fill_1 FILLER_74_605 ();
 sg13g2_fill_1 FILLER_74_611 ();
 sg13g2_decap_4 FILLER_74_627 ();
 sg13g2_fill_2 FILLER_74_652 ();
 sg13g2_decap_4 FILLER_74_666 ();
 sg13g2_decap_8 FILLER_74_684 ();
 sg13g2_fill_2 FILLER_74_703 ();
 sg13g2_fill_2 FILLER_74_715 ();
 sg13g2_fill_1 FILLER_74_717 ();
 sg13g2_decap_8 FILLER_74_724 ();
 sg13g2_fill_1 FILLER_74_731 ();
 sg13g2_fill_2 FILLER_74_736 ();
 sg13g2_fill_1 FILLER_74_738 ();
 sg13g2_decap_4 FILLER_74_743 ();
 sg13g2_fill_1 FILLER_74_747 ();
 sg13g2_fill_2 FILLER_74_773 ();
 sg13g2_fill_2 FILLER_74_792 ();
 sg13g2_fill_1 FILLER_74_794 ();
 sg13g2_decap_4 FILLER_74_807 ();
 sg13g2_fill_2 FILLER_74_811 ();
 sg13g2_fill_2 FILLER_74_821 ();
 sg13g2_fill_2 FILLER_74_828 ();
 sg13g2_decap_4 FILLER_74_835 ();
 sg13g2_fill_2 FILLER_74_839 ();
 sg13g2_fill_2 FILLER_74_856 ();
 sg13g2_fill_1 FILLER_74_858 ();
 sg13g2_fill_2 FILLER_74_894 ();
 sg13g2_decap_4 FILLER_74_911 ();
 sg13g2_fill_1 FILLER_74_944 ();
 sg13g2_fill_2 FILLER_74_957 ();
 sg13g2_decap_4 FILLER_74_965 ();
 sg13g2_decap_8 FILLER_74_1000 ();
 sg13g2_fill_2 FILLER_74_1007 ();
 sg13g2_fill_2 FILLER_74_1021 ();
 sg13g2_decap_8 FILLER_74_1032 ();
 sg13g2_decap_8 FILLER_74_1039 ();
 sg13g2_decap_8 FILLER_74_1046 ();
 sg13g2_decap_8 FILLER_74_1053 ();
 sg13g2_decap_8 FILLER_74_1060 ();
 sg13g2_decap_8 FILLER_74_1067 ();
 sg13g2_decap_8 FILLER_74_1074 ();
 sg13g2_decap_8 FILLER_74_1081 ();
 sg13g2_decap_8 FILLER_74_1088 ();
 sg13g2_decap_8 FILLER_74_1095 ();
 sg13g2_decap_8 FILLER_74_1102 ();
 sg13g2_decap_8 FILLER_74_1109 ();
 sg13g2_decap_8 FILLER_74_1116 ();
 sg13g2_decap_8 FILLER_74_1123 ();
 sg13g2_decap_8 FILLER_74_1130 ();
 sg13g2_decap_8 FILLER_74_1137 ();
 sg13g2_decap_8 FILLER_74_1144 ();
 sg13g2_decap_8 FILLER_74_1151 ();
 sg13g2_decap_8 FILLER_74_1158 ();
 sg13g2_decap_8 FILLER_74_1165 ();
 sg13g2_decap_8 FILLER_74_1172 ();
 sg13g2_decap_8 FILLER_74_1179 ();
 sg13g2_decap_8 FILLER_74_1186 ();
 sg13g2_decap_8 FILLER_74_1193 ();
 sg13g2_decap_8 FILLER_74_1200 ();
 sg13g2_decap_8 FILLER_74_1207 ();
 sg13g2_decap_8 FILLER_74_1214 ();
 sg13g2_decap_8 FILLER_74_1221 ();
 sg13g2_decap_8 FILLER_74_1228 ();
 sg13g2_decap_8 FILLER_74_1235 ();
 sg13g2_decap_8 FILLER_74_1242 ();
 sg13g2_decap_8 FILLER_74_1249 ();
 sg13g2_decap_8 FILLER_74_1256 ();
 sg13g2_decap_8 FILLER_74_1263 ();
 sg13g2_decap_8 FILLER_74_1270 ();
 sg13g2_decap_8 FILLER_74_1277 ();
 sg13g2_decap_8 FILLER_74_1284 ();
 sg13g2_decap_8 FILLER_74_1291 ();
 sg13g2_decap_8 FILLER_74_1298 ();
 sg13g2_decap_8 FILLER_74_1305 ();
 sg13g2_decap_8 FILLER_74_1312 ();
 sg13g2_decap_8 FILLER_74_1319 ();
 sg13g2_decap_8 FILLER_74_1326 ();
 sg13g2_decap_8 FILLER_74_1333 ();
 sg13g2_decap_8 FILLER_74_1340 ();
 sg13g2_decap_8 FILLER_74_1347 ();
 sg13g2_decap_8 FILLER_74_1354 ();
 sg13g2_decap_8 FILLER_74_1361 ();
 sg13g2_decap_8 FILLER_74_1368 ();
 sg13g2_decap_8 FILLER_74_1375 ();
 sg13g2_decap_8 FILLER_74_1382 ();
 sg13g2_decap_8 FILLER_74_1389 ();
 sg13g2_decap_8 FILLER_74_1396 ();
 sg13g2_decap_8 FILLER_74_1403 ();
 sg13g2_decap_8 FILLER_74_1410 ();
 sg13g2_decap_8 FILLER_74_1417 ();
 sg13g2_decap_8 FILLER_74_1424 ();
 sg13g2_decap_8 FILLER_74_1431 ();
 sg13g2_decap_8 FILLER_74_1438 ();
 sg13g2_decap_8 FILLER_74_1445 ();
 sg13g2_decap_8 FILLER_74_1452 ();
 sg13g2_decap_8 FILLER_74_1459 ();
 sg13g2_decap_8 FILLER_74_1466 ();
 sg13g2_decap_8 FILLER_74_1473 ();
 sg13g2_decap_8 FILLER_74_1480 ();
 sg13g2_decap_8 FILLER_74_1487 ();
 sg13g2_decap_8 FILLER_74_1494 ();
 sg13g2_decap_8 FILLER_74_1501 ();
 sg13g2_decap_8 FILLER_74_1508 ();
 sg13g2_decap_8 FILLER_74_1515 ();
 sg13g2_decap_8 FILLER_74_1522 ();
 sg13g2_decap_8 FILLER_74_1529 ();
 sg13g2_decap_8 FILLER_74_1536 ();
 sg13g2_decap_8 FILLER_74_1543 ();
 sg13g2_decap_8 FILLER_74_1550 ();
 sg13g2_decap_8 FILLER_74_1557 ();
 sg13g2_decap_8 FILLER_74_1564 ();
 sg13g2_decap_8 FILLER_74_1571 ();
 sg13g2_decap_8 FILLER_74_1578 ();
 sg13g2_decap_8 FILLER_74_1585 ();
 sg13g2_decap_8 FILLER_74_1592 ();
 sg13g2_decap_8 FILLER_74_1599 ();
 sg13g2_decap_8 FILLER_74_1606 ();
 sg13g2_decap_8 FILLER_74_1613 ();
 sg13g2_decap_8 FILLER_74_1620 ();
 sg13g2_decap_8 FILLER_74_1627 ();
 sg13g2_decap_8 FILLER_74_1634 ();
 sg13g2_decap_8 FILLER_74_1641 ();
 sg13g2_decap_8 FILLER_74_1648 ();
 sg13g2_decap_8 FILLER_74_1655 ();
 sg13g2_decap_8 FILLER_74_1662 ();
 sg13g2_decap_8 FILLER_74_1669 ();
 sg13g2_decap_8 FILLER_74_1676 ();
 sg13g2_decap_8 FILLER_74_1683 ();
 sg13g2_decap_8 FILLER_74_1690 ();
 sg13g2_decap_8 FILLER_74_1697 ();
 sg13g2_decap_8 FILLER_74_1704 ();
 sg13g2_decap_8 FILLER_74_1711 ();
 sg13g2_decap_8 FILLER_74_1718 ();
 sg13g2_decap_8 FILLER_74_1725 ();
 sg13g2_decap_8 FILLER_74_1732 ();
 sg13g2_decap_8 FILLER_74_1739 ();
 sg13g2_decap_8 FILLER_74_1746 ();
 sg13g2_decap_8 FILLER_74_1753 ();
 sg13g2_decap_8 FILLER_74_1760 ();
 sg13g2_fill_1 FILLER_74_1767 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_14 ();
 sg13g2_decap_8 FILLER_75_21 ();
 sg13g2_decap_8 FILLER_75_28 ();
 sg13g2_decap_8 FILLER_75_35 ();
 sg13g2_decap_8 FILLER_75_42 ();
 sg13g2_decap_8 FILLER_75_49 ();
 sg13g2_fill_2 FILLER_75_56 ();
 sg13g2_fill_1 FILLER_75_58 ();
 sg13g2_fill_2 FILLER_75_75 ();
 sg13g2_fill_1 FILLER_75_77 ();
 sg13g2_fill_1 FILLER_75_91 ();
 sg13g2_fill_1 FILLER_75_102 ();
 sg13g2_fill_1 FILLER_75_134 ();
 sg13g2_fill_2 FILLER_75_147 ();
 sg13g2_decap_8 FILLER_75_165 ();
 sg13g2_decap_4 FILLER_75_172 ();
 sg13g2_fill_2 FILLER_75_184 ();
 sg13g2_fill_1 FILLER_75_249 ();
 sg13g2_fill_2 FILLER_75_264 ();
 sg13g2_fill_2 FILLER_75_280 ();
 sg13g2_fill_2 FILLER_75_290 ();
 sg13g2_fill_1 FILLER_75_292 ();
 sg13g2_fill_2 FILLER_75_316 ();
 sg13g2_fill_1 FILLER_75_318 ();
 sg13g2_decap_8 FILLER_75_332 ();
 sg13g2_fill_1 FILLER_75_339 ();
 sg13g2_decap_4 FILLER_75_350 ();
 sg13g2_fill_2 FILLER_75_359 ();
 sg13g2_fill_1 FILLER_75_411 ();
 sg13g2_fill_2 FILLER_75_417 ();
 sg13g2_fill_1 FILLER_75_419 ();
 sg13g2_fill_1 FILLER_75_425 ();
 sg13g2_fill_2 FILLER_75_445 ();
 sg13g2_fill_1 FILLER_75_447 ();
 sg13g2_fill_2 FILLER_75_460 ();
 sg13g2_decap_8 FILLER_75_475 ();
 sg13g2_fill_1 FILLER_75_490 ();
 sg13g2_fill_2 FILLER_75_503 ();
 sg13g2_fill_1 FILLER_75_505 ();
 sg13g2_decap_4 FILLER_75_524 ();
 sg13g2_decap_8 FILLER_75_544 ();
 sg13g2_fill_1 FILLER_75_551 ();
 sg13g2_decap_8 FILLER_75_585 ();
 sg13g2_decap_8 FILLER_75_592 ();
 sg13g2_decap_8 FILLER_75_599 ();
 sg13g2_decap_8 FILLER_75_606 ();
 sg13g2_fill_1 FILLER_75_613 ();
 sg13g2_decap_8 FILLER_75_643 ();
 sg13g2_decap_4 FILLER_75_658 ();
 sg13g2_fill_2 FILLER_75_662 ();
 sg13g2_fill_2 FILLER_75_689 ();
 sg13g2_fill_1 FILLER_75_691 ();
 sg13g2_decap_8 FILLER_75_717 ();
 sg13g2_decap_4 FILLER_75_724 ();
 sg13g2_fill_2 FILLER_75_742 ();
 sg13g2_fill_1 FILLER_75_744 ();
 sg13g2_decap_4 FILLER_75_762 ();
 sg13g2_fill_1 FILLER_75_766 ();
 sg13g2_fill_2 FILLER_75_780 ();
 sg13g2_fill_1 FILLER_75_782 ();
 sg13g2_decap_4 FILLER_75_791 ();
 sg13g2_fill_2 FILLER_75_795 ();
 sg13g2_fill_2 FILLER_75_818 ();
 sg13g2_fill_1 FILLER_75_820 ();
 sg13g2_decap_4 FILLER_75_857 ();
 sg13g2_decap_8 FILLER_75_870 ();
 sg13g2_fill_1 FILLER_75_886 ();
 sg13g2_fill_2 FILLER_75_932 ();
 sg13g2_fill_1 FILLER_75_960 ();
 sg13g2_fill_1 FILLER_75_970 ();
 sg13g2_fill_2 FILLER_75_984 ();
 sg13g2_fill_1 FILLER_75_996 ();
 sg13g2_decap_8 FILLER_75_1023 ();
 sg13g2_decap_8 FILLER_75_1030 ();
 sg13g2_decap_8 FILLER_75_1037 ();
 sg13g2_decap_8 FILLER_75_1044 ();
 sg13g2_decap_8 FILLER_75_1051 ();
 sg13g2_decap_8 FILLER_75_1058 ();
 sg13g2_decap_8 FILLER_75_1065 ();
 sg13g2_decap_8 FILLER_75_1072 ();
 sg13g2_decap_8 FILLER_75_1079 ();
 sg13g2_decap_8 FILLER_75_1086 ();
 sg13g2_decap_8 FILLER_75_1093 ();
 sg13g2_decap_8 FILLER_75_1100 ();
 sg13g2_decap_8 FILLER_75_1107 ();
 sg13g2_decap_8 FILLER_75_1114 ();
 sg13g2_decap_8 FILLER_75_1121 ();
 sg13g2_decap_8 FILLER_75_1128 ();
 sg13g2_decap_8 FILLER_75_1135 ();
 sg13g2_decap_8 FILLER_75_1142 ();
 sg13g2_decap_8 FILLER_75_1149 ();
 sg13g2_decap_8 FILLER_75_1156 ();
 sg13g2_decap_8 FILLER_75_1163 ();
 sg13g2_decap_8 FILLER_75_1170 ();
 sg13g2_decap_8 FILLER_75_1177 ();
 sg13g2_decap_8 FILLER_75_1184 ();
 sg13g2_decap_8 FILLER_75_1191 ();
 sg13g2_decap_8 FILLER_75_1198 ();
 sg13g2_decap_8 FILLER_75_1205 ();
 sg13g2_decap_8 FILLER_75_1212 ();
 sg13g2_decap_8 FILLER_75_1219 ();
 sg13g2_decap_8 FILLER_75_1226 ();
 sg13g2_decap_8 FILLER_75_1233 ();
 sg13g2_decap_8 FILLER_75_1240 ();
 sg13g2_decap_8 FILLER_75_1247 ();
 sg13g2_decap_8 FILLER_75_1254 ();
 sg13g2_decap_8 FILLER_75_1261 ();
 sg13g2_decap_8 FILLER_75_1268 ();
 sg13g2_decap_8 FILLER_75_1275 ();
 sg13g2_decap_8 FILLER_75_1282 ();
 sg13g2_decap_8 FILLER_75_1289 ();
 sg13g2_decap_8 FILLER_75_1296 ();
 sg13g2_decap_8 FILLER_75_1303 ();
 sg13g2_decap_8 FILLER_75_1310 ();
 sg13g2_decap_8 FILLER_75_1317 ();
 sg13g2_decap_8 FILLER_75_1324 ();
 sg13g2_decap_8 FILLER_75_1331 ();
 sg13g2_decap_8 FILLER_75_1338 ();
 sg13g2_decap_8 FILLER_75_1345 ();
 sg13g2_decap_8 FILLER_75_1352 ();
 sg13g2_decap_8 FILLER_75_1359 ();
 sg13g2_decap_8 FILLER_75_1366 ();
 sg13g2_decap_8 FILLER_75_1373 ();
 sg13g2_decap_8 FILLER_75_1380 ();
 sg13g2_decap_8 FILLER_75_1387 ();
 sg13g2_decap_8 FILLER_75_1394 ();
 sg13g2_decap_8 FILLER_75_1401 ();
 sg13g2_decap_8 FILLER_75_1408 ();
 sg13g2_decap_8 FILLER_75_1415 ();
 sg13g2_decap_8 FILLER_75_1422 ();
 sg13g2_decap_8 FILLER_75_1429 ();
 sg13g2_decap_8 FILLER_75_1436 ();
 sg13g2_decap_8 FILLER_75_1443 ();
 sg13g2_decap_8 FILLER_75_1450 ();
 sg13g2_decap_8 FILLER_75_1457 ();
 sg13g2_decap_8 FILLER_75_1464 ();
 sg13g2_decap_8 FILLER_75_1471 ();
 sg13g2_decap_8 FILLER_75_1478 ();
 sg13g2_decap_8 FILLER_75_1485 ();
 sg13g2_decap_8 FILLER_75_1492 ();
 sg13g2_decap_8 FILLER_75_1499 ();
 sg13g2_decap_8 FILLER_75_1506 ();
 sg13g2_decap_8 FILLER_75_1513 ();
 sg13g2_decap_8 FILLER_75_1520 ();
 sg13g2_decap_8 FILLER_75_1527 ();
 sg13g2_decap_8 FILLER_75_1534 ();
 sg13g2_decap_8 FILLER_75_1541 ();
 sg13g2_decap_8 FILLER_75_1548 ();
 sg13g2_decap_8 FILLER_75_1555 ();
 sg13g2_decap_8 FILLER_75_1562 ();
 sg13g2_decap_8 FILLER_75_1569 ();
 sg13g2_decap_8 FILLER_75_1576 ();
 sg13g2_decap_8 FILLER_75_1583 ();
 sg13g2_decap_8 FILLER_75_1590 ();
 sg13g2_decap_8 FILLER_75_1597 ();
 sg13g2_decap_8 FILLER_75_1604 ();
 sg13g2_decap_8 FILLER_75_1611 ();
 sg13g2_decap_8 FILLER_75_1618 ();
 sg13g2_decap_8 FILLER_75_1625 ();
 sg13g2_decap_8 FILLER_75_1632 ();
 sg13g2_decap_8 FILLER_75_1639 ();
 sg13g2_decap_8 FILLER_75_1646 ();
 sg13g2_decap_8 FILLER_75_1653 ();
 sg13g2_decap_8 FILLER_75_1660 ();
 sg13g2_decap_8 FILLER_75_1667 ();
 sg13g2_decap_8 FILLER_75_1674 ();
 sg13g2_decap_8 FILLER_75_1681 ();
 sg13g2_decap_8 FILLER_75_1688 ();
 sg13g2_decap_8 FILLER_75_1695 ();
 sg13g2_decap_8 FILLER_75_1702 ();
 sg13g2_decap_8 FILLER_75_1709 ();
 sg13g2_decap_8 FILLER_75_1716 ();
 sg13g2_decap_8 FILLER_75_1723 ();
 sg13g2_decap_8 FILLER_75_1730 ();
 sg13g2_decap_8 FILLER_75_1737 ();
 sg13g2_decap_8 FILLER_75_1744 ();
 sg13g2_decap_8 FILLER_75_1751 ();
 sg13g2_decap_8 FILLER_75_1758 ();
 sg13g2_fill_2 FILLER_75_1765 ();
 sg13g2_fill_1 FILLER_75_1767 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_8 FILLER_76_21 ();
 sg13g2_decap_8 FILLER_76_28 ();
 sg13g2_decap_8 FILLER_76_35 ();
 sg13g2_decap_8 FILLER_76_42 ();
 sg13g2_decap_4 FILLER_76_49 ();
 sg13g2_fill_1 FILLER_76_66 ();
 sg13g2_fill_2 FILLER_76_72 ();
 sg13g2_fill_1 FILLER_76_74 ();
 sg13g2_fill_1 FILLER_76_89 ();
 sg13g2_decap_8 FILLER_76_97 ();
 sg13g2_decap_4 FILLER_76_104 ();
 sg13g2_fill_2 FILLER_76_108 ();
 sg13g2_decap_8 FILLER_76_127 ();
 sg13g2_decap_8 FILLER_76_134 ();
 sg13g2_fill_1 FILLER_76_141 ();
 sg13g2_fill_2 FILLER_76_161 ();
 sg13g2_fill_1 FILLER_76_163 ();
 sg13g2_fill_1 FILLER_76_248 ();
 sg13g2_fill_2 FILLER_76_280 ();
 sg13g2_fill_1 FILLER_76_282 ();
 sg13g2_fill_2 FILLER_76_319 ();
 sg13g2_fill_1 FILLER_76_321 ();
 sg13g2_fill_2 FILLER_76_330 ();
 sg13g2_fill_2 FILLER_76_355 ();
 sg13g2_fill_1 FILLER_76_357 ();
 sg13g2_fill_1 FILLER_76_365 ();
 sg13g2_fill_1 FILLER_76_375 ();
 sg13g2_fill_2 FILLER_76_392 ();
 sg13g2_fill_1 FILLER_76_416 ();
 sg13g2_fill_1 FILLER_76_424 ();
 sg13g2_decap_4 FILLER_76_451 ();
 sg13g2_decap_8 FILLER_76_468 ();
 sg13g2_fill_1 FILLER_76_475 ();
 sg13g2_fill_1 FILLER_76_484 ();
 sg13g2_fill_2 FILLER_76_498 ();
 sg13g2_fill_1 FILLER_76_500 ();
 sg13g2_decap_8 FILLER_76_517 ();
 sg13g2_decap_4 FILLER_76_550 ();
 sg13g2_fill_2 FILLER_76_554 ();
 sg13g2_decap_8 FILLER_76_574 ();
 sg13g2_decap_8 FILLER_76_581 ();
 sg13g2_decap_8 FILLER_76_588 ();
 sg13g2_fill_2 FILLER_76_595 ();
 sg13g2_fill_1 FILLER_76_597 ();
 sg13g2_decap_8 FILLER_76_606 ();
 sg13g2_decap_4 FILLER_76_613 ();
 sg13g2_decap_4 FILLER_76_642 ();
 sg13g2_fill_1 FILLER_76_646 ();
 sg13g2_fill_2 FILLER_76_664 ();
 sg13g2_decap_4 FILLER_76_683 ();
 sg13g2_fill_1 FILLER_76_687 ();
 sg13g2_decap_8 FILLER_76_691 ();
 sg13g2_fill_2 FILLER_76_698 ();
 sg13g2_decap_4 FILLER_76_709 ();
 sg13g2_fill_1 FILLER_76_713 ();
 sg13g2_fill_2 FILLER_76_726 ();
 sg13g2_fill_2 FILLER_76_741 ();
 sg13g2_fill_1 FILLER_76_743 ();
 sg13g2_fill_2 FILLER_76_762 ();
 sg13g2_fill_1 FILLER_76_764 ();
 sg13g2_fill_2 FILLER_76_770 ();
 sg13g2_fill_1 FILLER_76_777 ();
 sg13g2_decap_8 FILLER_76_785 ();
 sg13g2_decap_8 FILLER_76_792 ();
 sg13g2_fill_1 FILLER_76_799 ();
 sg13g2_decap_8 FILLER_76_813 ();
 sg13g2_decap_4 FILLER_76_820 ();
 sg13g2_fill_1 FILLER_76_824 ();
 sg13g2_fill_1 FILLER_76_830 ();
 sg13g2_fill_1 FILLER_76_839 ();
 sg13g2_fill_1 FILLER_76_849 ();
 sg13g2_fill_2 FILLER_76_863 ();
 sg13g2_fill_1 FILLER_76_865 ();
 sg13g2_fill_1 FILLER_76_917 ();
 sg13g2_decap_8 FILLER_76_961 ();
 sg13g2_decap_8 FILLER_76_968 ();
 sg13g2_fill_2 FILLER_76_975 ();
 sg13g2_fill_1 FILLER_76_977 ();
 sg13g2_decap_8 FILLER_76_982 ();
 sg13g2_fill_2 FILLER_76_989 ();
 sg13g2_decap_8 FILLER_76_996 ();
 sg13g2_decap_8 FILLER_76_1003 ();
 sg13g2_decap_8 FILLER_76_1010 ();
 sg13g2_decap_8 FILLER_76_1017 ();
 sg13g2_decap_8 FILLER_76_1024 ();
 sg13g2_decap_8 FILLER_76_1031 ();
 sg13g2_decap_8 FILLER_76_1038 ();
 sg13g2_decap_8 FILLER_76_1045 ();
 sg13g2_decap_8 FILLER_76_1052 ();
 sg13g2_decap_8 FILLER_76_1059 ();
 sg13g2_decap_8 FILLER_76_1066 ();
 sg13g2_decap_8 FILLER_76_1073 ();
 sg13g2_decap_8 FILLER_76_1080 ();
 sg13g2_decap_8 FILLER_76_1087 ();
 sg13g2_decap_8 FILLER_76_1094 ();
 sg13g2_decap_8 FILLER_76_1101 ();
 sg13g2_decap_8 FILLER_76_1108 ();
 sg13g2_decap_8 FILLER_76_1115 ();
 sg13g2_decap_8 FILLER_76_1122 ();
 sg13g2_decap_8 FILLER_76_1129 ();
 sg13g2_decap_8 FILLER_76_1136 ();
 sg13g2_decap_8 FILLER_76_1143 ();
 sg13g2_decap_8 FILLER_76_1150 ();
 sg13g2_decap_8 FILLER_76_1157 ();
 sg13g2_decap_8 FILLER_76_1164 ();
 sg13g2_decap_8 FILLER_76_1171 ();
 sg13g2_decap_8 FILLER_76_1178 ();
 sg13g2_decap_8 FILLER_76_1185 ();
 sg13g2_decap_8 FILLER_76_1192 ();
 sg13g2_decap_8 FILLER_76_1199 ();
 sg13g2_decap_8 FILLER_76_1206 ();
 sg13g2_decap_8 FILLER_76_1213 ();
 sg13g2_decap_8 FILLER_76_1220 ();
 sg13g2_decap_8 FILLER_76_1227 ();
 sg13g2_decap_8 FILLER_76_1234 ();
 sg13g2_decap_8 FILLER_76_1241 ();
 sg13g2_decap_8 FILLER_76_1248 ();
 sg13g2_decap_8 FILLER_76_1255 ();
 sg13g2_decap_8 FILLER_76_1262 ();
 sg13g2_decap_8 FILLER_76_1269 ();
 sg13g2_decap_8 FILLER_76_1276 ();
 sg13g2_decap_8 FILLER_76_1283 ();
 sg13g2_decap_8 FILLER_76_1290 ();
 sg13g2_decap_8 FILLER_76_1297 ();
 sg13g2_decap_8 FILLER_76_1304 ();
 sg13g2_decap_8 FILLER_76_1311 ();
 sg13g2_decap_8 FILLER_76_1318 ();
 sg13g2_decap_8 FILLER_76_1325 ();
 sg13g2_decap_8 FILLER_76_1332 ();
 sg13g2_decap_8 FILLER_76_1339 ();
 sg13g2_decap_8 FILLER_76_1346 ();
 sg13g2_decap_8 FILLER_76_1353 ();
 sg13g2_decap_8 FILLER_76_1360 ();
 sg13g2_decap_8 FILLER_76_1367 ();
 sg13g2_decap_8 FILLER_76_1374 ();
 sg13g2_decap_8 FILLER_76_1381 ();
 sg13g2_decap_8 FILLER_76_1388 ();
 sg13g2_decap_8 FILLER_76_1395 ();
 sg13g2_decap_8 FILLER_76_1402 ();
 sg13g2_decap_8 FILLER_76_1409 ();
 sg13g2_decap_8 FILLER_76_1416 ();
 sg13g2_decap_8 FILLER_76_1423 ();
 sg13g2_decap_8 FILLER_76_1430 ();
 sg13g2_decap_8 FILLER_76_1437 ();
 sg13g2_decap_8 FILLER_76_1444 ();
 sg13g2_decap_8 FILLER_76_1451 ();
 sg13g2_decap_8 FILLER_76_1458 ();
 sg13g2_decap_8 FILLER_76_1465 ();
 sg13g2_decap_8 FILLER_76_1472 ();
 sg13g2_decap_8 FILLER_76_1479 ();
 sg13g2_decap_8 FILLER_76_1486 ();
 sg13g2_decap_8 FILLER_76_1493 ();
 sg13g2_decap_8 FILLER_76_1500 ();
 sg13g2_decap_8 FILLER_76_1507 ();
 sg13g2_decap_8 FILLER_76_1514 ();
 sg13g2_decap_8 FILLER_76_1521 ();
 sg13g2_decap_8 FILLER_76_1528 ();
 sg13g2_decap_8 FILLER_76_1535 ();
 sg13g2_decap_8 FILLER_76_1542 ();
 sg13g2_decap_8 FILLER_76_1549 ();
 sg13g2_decap_8 FILLER_76_1556 ();
 sg13g2_decap_8 FILLER_76_1563 ();
 sg13g2_decap_8 FILLER_76_1570 ();
 sg13g2_decap_8 FILLER_76_1577 ();
 sg13g2_decap_8 FILLER_76_1584 ();
 sg13g2_decap_8 FILLER_76_1591 ();
 sg13g2_decap_8 FILLER_76_1598 ();
 sg13g2_decap_8 FILLER_76_1605 ();
 sg13g2_decap_8 FILLER_76_1612 ();
 sg13g2_decap_8 FILLER_76_1619 ();
 sg13g2_decap_8 FILLER_76_1626 ();
 sg13g2_decap_8 FILLER_76_1633 ();
 sg13g2_decap_8 FILLER_76_1640 ();
 sg13g2_decap_8 FILLER_76_1647 ();
 sg13g2_decap_8 FILLER_76_1654 ();
 sg13g2_decap_8 FILLER_76_1661 ();
 sg13g2_decap_8 FILLER_76_1668 ();
 sg13g2_decap_8 FILLER_76_1675 ();
 sg13g2_decap_8 FILLER_76_1682 ();
 sg13g2_decap_8 FILLER_76_1689 ();
 sg13g2_decap_8 FILLER_76_1696 ();
 sg13g2_decap_8 FILLER_76_1703 ();
 sg13g2_decap_8 FILLER_76_1710 ();
 sg13g2_decap_8 FILLER_76_1717 ();
 sg13g2_decap_8 FILLER_76_1724 ();
 sg13g2_decap_8 FILLER_76_1731 ();
 sg13g2_decap_8 FILLER_76_1738 ();
 sg13g2_decap_8 FILLER_76_1745 ();
 sg13g2_decap_8 FILLER_76_1752 ();
 sg13g2_decap_8 FILLER_76_1759 ();
 sg13g2_fill_2 FILLER_76_1766 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_fill_2 FILLER_77_28 ();
 sg13g2_fill_1 FILLER_77_56 ();
 sg13g2_fill_2 FILLER_77_70 ();
 sg13g2_fill_1 FILLER_77_72 ();
 sg13g2_fill_1 FILLER_77_79 ();
 sg13g2_fill_2 FILLER_77_85 ();
 sg13g2_decap_4 FILLER_77_113 ();
 sg13g2_fill_1 FILLER_77_136 ();
 sg13g2_fill_2 FILLER_77_151 ();
 sg13g2_fill_1 FILLER_77_153 ();
 sg13g2_decap_8 FILLER_77_180 ();
 sg13g2_fill_1 FILLER_77_232 ();
 sg13g2_fill_2 FILLER_77_238 ();
 sg13g2_fill_1 FILLER_77_240 ();
 sg13g2_fill_1 FILLER_77_272 ();
 sg13g2_decap_8 FILLER_77_313 ();
 sg13g2_fill_1 FILLER_77_326 ();
 sg13g2_decap_4 FILLER_77_332 ();
 sg13g2_fill_2 FILLER_77_336 ();
 sg13g2_fill_2 FILLER_77_354 ();
 sg13g2_fill_1 FILLER_77_356 ();
 sg13g2_fill_1 FILLER_77_373 ();
 sg13g2_fill_2 FILLER_77_426 ();
 sg13g2_decap_8 FILLER_77_454 ();
 sg13g2_decap_8 FILLER_77_461 ();
 sg13g2_decap_8 FILLER_77_468 ();
 sg13g2_fill_2 FILLER_77_475 ();
 sg13g2_fill_2 FILLER_77_485 ();
 sg13g2_decap_8 FILLER_77_492 ();
 sg13g2_decap_8 FILLER_77_499 ();
 sg13g2_decap_8 FILLER_77_506 ();
 sg13g2_decap_8 FILLER_77_513 ();
 sg13g2_decap_8 FILLER_77_520 ();
 sg13g2_fill_2 FILLER_77_527 ();
 sg13g2_fill_1 FILLER_77_529 ();
 sg13g2_decap_8 FILLER_77_543 ();
 sg13g2_decap_8 FILLER_77_550 ();
 sg13g2_decap_8 FILLER_77_557 ();
 sg13g2_decap_8 FILLER_77_564 ();
 sg13g2_decap_8 FILLER_77_571 ();
 sg13g2_decap_8 FILLER_77_578 ();
 sg13g2_decap_8 FILLER_77_585 ();
 sg13g2_decap_8 FILLER_77_592 ();
 sg13g2_decap_8 FILLER_77_599 ();
 sg13g2_decap_8 FILLER_77_606 ();
 sg13g2_decap_8 FILLER_77_613 ();
 sg13g2_decap_4 FILLER_77_620 ();
 sg13g2_fill_1 FILLER_77_624 ();
 sg13g2_decap_4 FILLER_77_634 ();
 sg13g2_fill_1 FILLER_77_638 ();
 sg13g2_fill_2 FILLER_77_661 ();
 sg13g2_fill_2 FILLER_77_680 ();
 sg13g2_fill_2 FILLER_77_713 ();
 sg13g2_fill_1 FILLER_77_741 ();
 sg13g2_decap_4 FILLER_77_746 ();
 sg13g2_fill_1 FILLER_77_750 ();
 sg13g2_fill_1 FILLER_77_791 ();
 sg13g2_fill_2 FILLER_77_813 ();
 sg13g2_fill_1 FILLER_77_815 ();
 sg13g2_decap_8 FILLER_77_851 ();
 sg13g2_fill_1 FILLER_77_858 ();
 sg13g2_decap_8 FILLER_77_869 ();
 sg13g2_decap_8 FILLER_77_876 ();
 sg13g2_decap_8 FILLER_77_883 ();
 sg13g2_decap_8 FILLER_77_895 ();
 sg13g2_fill_2 FILLER_77_902 ();
 sg13g2_fill_1 FILLER_77_904 ();
 sg13g2_decap_8 FILLER_77_914 ();
 sg13g2_decap_8 FILLER_77_921 ();
 sg13g2_decap_8 FILLER_77_928 ();
 sg13g2_decap_8 FILLER_77_944 ();
 sg13g2_decap_8 FILLER_77_951 ();
 sg13g2_decap_8 FILLER_77_958 ();
 sg13g2_decap_8 FILLER_77_965 ();
 sg13g2_decap_8 FILLER_77_972 ();
 sg13g2_decap_8 FILLER_77_979 ();
 sg13g2_decap_8 FILLER_77_986 ();
 sg13g2_decap_8 FILLER_77_993 ();
 sg13g2_decap_8 FILLER_77_1000 ();
 sg13g2_decap_8 FILLER_77_1007 ();
 sg13g2_decap_8 FILLER_77_1014 ();
 sg13g2_decap_8 FILLER_77_1021 ();
 sg13g2_decap_8 FILLER_77_1028 ();
 sg13g2_decap_8 FILLER_77_1035 ();
 sg13g2_decap_8 FILLER_77_1042 ();
 sg13g2_decap_8 FILLER_77_1049 ();
 sg13g2_decap_8 FILLER_77_1056 ();
 sg13g2_decap_8 FILLER_77_1063 ();
 sg13g2_decap_8 FILLER_77_1070 ();
 sg13g2_decap_8 FILLER_77_1077 ();
 sg13g2_decap_8 FILLER_77_1084 ();
 sg13g2_decap_8 FILLER_77_1091 ();
 sg13g2_decap_8 FILLER_77_1098 ();
 sg13g2_decap_8 FILLER_77_1105 ();
 sg13g2_decap_8 FILLER_77_1112 ();
 sg13g2_decap_8 FILLER_77_1119 ();
 sg13g2_decap_8 FILLER_77_1126 ();
 sg13g2_decap_8 FILLER_77_1133 ();
 sg13g2_decap_8 FILLER_77_1140 ();
 sg13g2_decap_8 FILLER_77_1147 ();
 sg13g2_decap_8 FILLER_77_1154 ();
 sg13g2_decap_8 FILLER_77_1161 ();
 sg13g2_decap_8 FILLER_77_1168 ();
 sg13g2_decap_8 FILLER_77_1175 ();
 sg13g2_decap_8 FILLER_77_1182 ();
 sg13g2_decap_8 FILLER_77_1189 ();
 sg13g2_decap_8 FILLER_77_1196 ();
 sg13g2_decap_8 FILLER_77_1203 ();
 sg13g2_decap_8 FILLER_77_1210 ();
 sg13g2_decap_8 FILLER_77_1217 ();
 sg13g2_decap_8 FILLER_77_1224 ();
 sg13g2_decap_8 FILLER_77_1231 ();
 sg13g2_decap_8 FILLER_77_1238 ();
 sg13g2_decap_8 FILLER_77_1245 ();
 sg13g2_decap_8 FILLER_77_1252 ();
 sg13g2_decap_8 FILLER_77_1259 ();
 sg13g2_decap_8 FILLER_77_1266 ();
 sg13g2_decap_8 FILLER_77_1273 ();
 sg13g2_decap_8 FILLER_77_1280 ();
 sg13g2_decap_8 FILLER_77_1287 ();
 sg13g2_decap_8 FILLER_77_1294 ();
 sg13g2_decap_8 FILLER_77_1301 ();
 sg13g2_decap_8 FILLER_77_1308 ();
 sg13g2_decap_8 FILLER_77_1315 ();
 sg13g2_decap_8 FILLER_77_1322 ();
 sg13g2_decap_8 FILLER_77_1329 ();
 sg13g2_decap_8 FILLER_77_1336 ();
 sg13g2_decap_8 FILLER_77_1343 ();
 sg13g2_decap_8 FILLER_77_1350 ();
 sg13g2_decap_8 FILLER_77_1357 ();
 sg13g2_decap_8 FILLER_77_1364 ();
 sg13g2_decap_8 FILLER_77_1371 ();
 sg13g2_decap_8 FILLER_77_1378 ();
 sg13g2_decap_8 FILLER_77_1385 ();
 sg13g2_decap_8 FILLER_77_1392 ();
 sg13g2_decap_8 FILLER_77_1399 ();
 sg13g2_decap_8 FILLER_77_1406 ();
 sg13g2_decap_8 FILLER_77_1413 ();
 sg13g2_decap_8 FILLER_77_1420 ();
 sg13g2_decap_8 FILLER_77_1427 ();
 sg13g2_decap_8 FILLER_77_1434 ();
 sg13g2_decap_8 FILLER_77_1441 ();
 sg13g2_decap_8 FILLER_77_1448 ();
 sg13g2_decap_8 FILLER_77_1455 ();
 sg13g2_decap_8 FILLER_77_1462 ();
 sg13g2_decap_8 FILLER_77_1469 ();
 sg13g2_decap_8 FILLER_77_1476 ();
 sg13g2_decap_8 FILLER_77_1483 ();
 sg13g2_decap_8 FILLER_77_1490 ();
 sg13g2_decap_8 FILLER_77_1497 ();
 sg13g2_decap_8 FILLER_77_1504 ();
 sg13g2_decap_8 FILLER_77_1511 ();
 sg13g2_decap_8 FILLER_77_1518 ();
 sg13g2_decap_8 FILLER_77_1525 ();
 sg13g2_decap_8 FILLER_77_1532 ();
 sg13g2_decap_8 FILLER_77_1539 ();
 sg13g2_decap_8 FILLER_77_1546 ();
 sg13g2_decap_8 FILLER_77_1553 ();
 sg13g2_decap_8 FILLER_77_1560 ();
 sg13g2_decap_8 FILLER_77_1567 ();
 sg13g2_decap_8 FILLER_77_1574 ();
 sg13g2_decap_8 FILLER_77_1581 ();
 sg13g2_decap_8 FILLER_77_1588 ();
 sg13g2_decap_8 FILLER_77_1595 ();
 sg13g2_decap_8 FILLER_77_1602 ();
 sg13g2_decap_8 FILLER_77_1609 ();
 sg13g2_decap_8 FILLER_77_1616 ();
 sg13g2_decap_8 FILLER_77_1623 ();
 sg13g2_decap_8 FILLER_77_1630 ();
 sg13g2_decap_8 FILLER_77_1637 ();
 sg13g2_decap_8 FILLER_77_1644 ();
 sg13g2_decap_8 FILLER_77_1651 ();
 sg13g2_decap_8 FILLER_77_1658 ();
 sg13g2_decap_8 FILLER_77_1665 ();
 sg13g2_decap_8 FILLER_77_1672 ();
 sg13g2_decap_8 FILLER_77_1679 ();
 sg13g2_decap_8 FILLER_77_1686 ();
 sg13g2_decap_8 FILLER_77_1693 ();
 sg13g2_decap_8 FILLER_77_1700 ();
 sg13g2_decap_8 FILLER_77_1707 ();
 sg13g2_decap_8 FILLER_77_1714 ();
 sg13g2_decap_8 FILLER_77_1721 ();
 sg13g2_decap_8 FILLER_77_1728 ();
 sg13g2_decap_8 FILLER_77_1735 ();
 sg13g2_decap_8 FILLER_77_1742 ();
 sg13g2_decap_8 FILLER_77_1749 ();
 sg13g2_decap_8 FILLER_77_1756 ();
 sg13g2_decap_4 FILLER_77_1763 ();
 sg13g2_fill_1 FILLER_77_1767 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_decap_8 FILLER_78_28 ();
 sg13g2_decap_4 FILLER_78_35 ();
 sg13g2_fill_2 FILLER_78_39 ();
 sg13g2_fill_2 FILLER_78_59 ();
 sg13g2_fill_1 FILLER_78_61 ();
 sg13g2_fill_2 FILLER_78_67 ();
 sg13g2_fill_2 FILLER_78_78 ();
 sg13g2_fill_1 FILLER_78_80 ();
 sg13g2_fill_2 FILLER_78_95 ();
 sg13g2_fill_1 FILLER_78_118 ();
 sg13g2_decap_4 FILLER_78_170 ();
 sg13g2_fill_1 FILLER_78_174 ();
 sg13g2_fill_2 FILLER_78_201 ();
 sg13g2_fill_2 FILLER_78_212 ();
 sg13g2_fill_1 FILLER_78_214 ();
 sg13g2_fill_2 FILLER_78_238 ();
 sg13g2_fill_1 FILLER_78_240 ();
 sg13g2_fill_2 FILLER_78_250 ();
 sg13g2_decap_8 FILLER_78_283 ();
 sg13g2_fill_2 FILLER_78_290 ();
 sg13g2_fill_1 FILLER_78_292 ();
 sg13g2_decap_4 FILLER_78_302 ();
 sg13g2_fill_2 FILLER_78_337 ();
 sg13g2_fill_1 FILLER_78_339 ();
 sg13g2_decap_4 FILLER_78_375 ();
 sg13g2_fill_1 FILLER_78_379 ();
 sg13g2_decap_8 FILLER_78_389 ();
 sg13g2_decap_8 FILLER_78_396 ();
 sg13g2_decap_8 FILLER_78_403 ();
 sg13g2_decap_8 FILLER_78_410 ();
 sg13g2_decap_8 FILLER_78_417 ();
 sg13g2_decap_8 FILLER_78_424 ();
 sg13g2_decap_8 FILLER_78_431 ();
 sg13g2_decap_8 FILLER_78_438 ();
 sg13g2_decap_8 FILLER_78_445 ();
 sg13g2_decap_8 FILLER_78_452 ();
 sg13g2_decap_8 FILLER_78_459 ();
 sg13g2_decap_8 FILLER_78_466 ();
 sg13g2_decap_8 FILLER_78_473 ();
 sg13g2_decap_8 FILLER_78_480 ();
 sg13g2_decap_8 FILLER_78_487 ();
 sg13g2_decap_8 FILLER_78_494 ();
 sg13g2_decap_8 FILLER_78_501 ();
 sg13g2_decap_8 FILLER_78_508 ();
 sg13g2_decap_8 FILLER_78_515 ();
 sg13g2_decap_8 FILLER_78_522 ();
 sg13g2_decap_8 FILLER_78_529 ();
 sg13g2_decap_8 FILLER_78_536 ();
 sg13g2_decap_8 FILLER_78_543 ();
 sg13g2_decap_8 FILLER_78_550 ();
 sg13g2_decap_8 FILLER_78_557 ();
 sg13g2_decap_8 FILLER_78_564 ();
 sg13g2_decap_8 FILLER_78_571 ();
 sg13g2_decap_8 FILLER_78_578 ();
 sg13g2_decap_8 FILLER_78_585 ();
 sg13g2_decap_8 FILLER_78_592 ();
 sg13g2_decap_8 FILLER_78_599 ();
 sg13g2_decap_8 FILLER_78_606 ();
 sg13g2_decap_8 FILLER_78_613 ();
 sg13g2_decap_8 FILLER_78_620 ();
 sg13g2_decap_8 FILLER_78_627 ();
 sg13g2_decap_8 FILLER_78_634 ();
 sg13g2_decap_4 FILLER_78_641 ();
 sg13g2_fill_2 FILLER_78_645 ();
 sg13g2_fill_2 FILLER_78_659 ();
 sg13g2_fill_1 FILLER_78_661 ();
 sg13g2_decap_8 FILLER_78_679 ();
 sg13g2_decap_8 FILLER_78_686 ();
 sg13g2_decap_4 FILLER_78_693 ();
 sg13g2_decap_8 FILLER_78_702 ();
 sg13g2_decap_8 FILLER_78_709 ();
 sg13g2_fill_2 FILLER_78_716 ();
 sg13g2_decap_4 FILLER_78_723 ();
 sg13g2_fill_1 FILLER_78_727 ();
 sg13g2_fill_2 FILLER_78_736 ();
 sg13g2_fill_1 FILLER_78_738 ();
 sg13g2_decap_8 FILLER_78_760 ();
 sg13g2_fill_2 FILLER_78_767 ();
 sg13g2_decap_8 FILLER_78_772 ();
 sg13g2_fill_2 FILLER_78_779 ();
 sg13g2_decap_8 FILLER_78_786 ();
 sg13g2_decap_8 FILLER_78_793 ();
 sg13g2_fill_2 FILLER_78_800 ();
 sg13g2_decap_8 FILLER_78_807 ();
 sg13g2_decap_8 FILLER_78_814 ();
 sg13g2_fill_2 FILLER_78_821 ();
 sg13g2_fill_1 FILLER_78_823 ();
 sg13g2_decap_8 FILLER_78_829 ();
 sg13g2_decap_8 FILLER_78_836 ();
 sg13g2_decap_8 FILLER_78_843 ();
 sg13g2_decap_8 FILLER_78_850 ();
 sg13g2_decap_8 FILLER_78_857 ();
 sg13g2_decap_8 FILLER_78_864 ();
 sg13g2_decap_8 FILLER_78_871 ();
 sg13g2_decap_8 FILLER_78_878 ();
 sg13g2_decap_8 FILLER_78_885 ();
 sg13g2_decap_8 FILLER_78_892 ();
 sg13g2_decap_8 FILLER_78_899 ();
 sg13g2_decap_8 FILLER_78_906 ();
 sg13g2_decap_8 FILLER_78_913 ();
 sg13g2_decap_8 FILLER_78_920 ();
 sg13g2_decap_8 FILLER_78_927 ();
 sg13g2_decap_8 FILLER_78_934 ();
 sg13g2_decap_8 FILLER_78_941 ();
 sg13g2_decap_8 FILLER_78_948 ();
 sg13g2_decap_8 FILLER_78_955 ();
 sg13g2_decap_8 FILLER_78_962 ();
 sg13g2_decap_8 FILLER_78_969 ();
 sg13g2_decap_8 FILLER_78_976 ();
 sg13g2_decap_8 FILLER_78_983 ();
 sg13g2_decap_8 FILLER_78_990 ();
 sg13g2_decap_8 FILLER_78_997 ();
 sg13g2_decap_8 FILLER_78_1004 ();
 sg13g2_decap_8 FILLER_78_1011 ();
 sg13g2_decap_8 FILLER_78_1018 ();
 sg13g2_decap_8 FILLER_78_1025 ();
 sg13g2_decap_8 FILLER_78_1032 ();
 sg13g2_decap_8 FILLER_78_1039 ();
 sg13g2_decap_8 FILLER_78_1046 ();
 sg13g2_decap_8 FILLER_78_1053 ();
 sg13g2_decap_8 FILLER_78_1060 ();
 sg13g2_decap_8 FILLER_78_1067 ();
 sg13g2_decap_8 FILLER_78_1074 ();
 sg13g2_decap_8 FILLER_78_1081 ();
 sg13g2_decap_8 FILLER_78_1088 ();
 sg13g2_decap_8 FILLER_78_1095 ();
 sg13g2_decap_8 FILLER_78_1102 ();
 sg13g2_decap_8 FILLER_78_1109 ();
 sg13g2_decap_8 FILLER_78_1116 ();
 sg13g2_decap_8 FILLER_78_1123 ();
 sg13g2_decap_8 FILLER_78_1130 ();
 sg13g2_decap_8 FILLER_78_1137 ();
 sg13g2_decap_8 FILLER_78_1144 ();
 sg13g2_decap_8 FILLER_78_1151 ();
 sg13g2_decap_8 FILLER_78_1158 ();
 sg13g2_decap_8 FILLER_78_1165 ();
 sg13g2_decap_8 FILLER_78_1172 ();
 sg13g2_decap_8 FILLER_78_1179 ();
 sg13g2_decap_8 FILLER_78_1186 ();
 sg13g2_decap_8 FILLER_78_1193 ();
 sg13g2_decap_8 FILLER_78_1200 ();
 sg13g2_decap_8 FILLER_78_1207 ();
 sg13g2_decap_8 FILLER_78_1214 ();
 sg13g2_decap_8 FILLER_78_1221 ();
 sg13g2_decap_8 FILLER_78_1228 ();
 sg13g2_decap_8 FILLER_78_1235 ();
 sg13g2_decap_8 FILLER_78_1242 ();
 sg13g2_decap_8 FILLER_78_1249 ();
 sg13g2_decap_8 FILLER_78_1256 ();
 sg13g2_decap_8 FILLER_78_1263 ();
 sg13g2_decap_8 FILLER_78_1270 ();
 sg13g2_decap_8 FILLER_78_1277 ();
 sg13g2_decap_8 FILLER_78_1284 ();
 sg13g2_decap_8 FILLER_78_1291 ();
 sg13g2_decap_8 FILLER_78_1298 ();
 sg13g2_decap_8 FILLER_78_1305 ();
 sg13g2_decap_8 FILLER_78_1312 ();
 sg13g2_decap_8 FILLER_78_1319 ();
 sg13g2_decap_8 FILLER_78_1326 ();
 sg13g2_decap_8 FILLER_78_1333 ();
 sg13g2_decap_8 FILLER_78_1340 ();
 sg13g2_decap_8 FILLER_78_1347 ();
 sg13g2_decap_8 FILLER_78_1354 ();
 sg13g2_decap_8 FILLER_78_1361 ();
 sg13g2_decap_8 FILLER_78_1368 ();
 sg13g2_decap_8 FILLER_78_1375 ();
 sg13g2_decap_8 FILLER_78_1382 ();
 sg13g2_decap_8 FILLER_78_1389 ();
 sg13g2_decap_8 FILLER_78_1396 ();
 sg13g2_decap_8 FILLER_78_1403 ();
 sg13g2_decap_8 FILLER_78_1410 ();
 sg13g2_decap_8 FILLER_78_1417 ();
 sg13g2_decap_8 FILLER_78_1424 ();
 sg13g2_decap_8 FILLER_78_1431 ();
 sg13g2_decap_8 FILLER_78_1438 ();
 sg13g2_decap_8 FILLER_78_1445 ();
 sg13g2_decap_8 FILLER_78_1452 ();
 sg13g2_decap_8 FILLER_78_1459 ();
 sg13g2_decap_8 FILLER_78_1466 ();
 sg13g2_decap_8 FILLER_78_1473 ();
 sg13g2_decap_8 FILLER_78_1480 ();
 sg13g2_decap_8 FILLER_78_1487 ();
 sg13g2_decap_8 FILLER_78_1494 ();
 sg13g2_decap_8 FILLER_78_1501 ();
 sg13g2_decap_8 FILLER_78_1508 ();
 sg13g2_decap_8 FILLER_78_1515 ();
 sg13g2_decap_8 FILLER_78_1522 ();
 sg13g2_decap_8 FILLER_78_1529 ();
 sg13g2_decap_8 FILLER_78_1536 ();
 sg13g2_decap_8 FILLER_78_1543 ();
 sg13g2_decap_8 FILLER_78_1550 ();
 sg13g2_decap_8 FILLER_78_1557 ();
 sg13g2_decap_8 FILLER_78_1564 ();
 sg13g2_decap_8 FILLER_78_1571 ();
 sg13g2_decap_8 FILLER_78_1578 ();
 sg13g2_decap_8 FILLER_78_1585 ();
 sg13g2_decap_8 FILLER_78_1592 ();
 sg13g2_decap_8 FILLER_78_1599 ();
 sg13g2_decap_8 FILLER_78_1606 ();
 sg13g2_decap_8 FILLER_78_1613 ();
 sg13g2_decap_8 FILLER_78_1620 ();
 sg13g2_decap_8 FILLER_78_1627 ();
 sg13g2_decap_8 FILLER_78_1634 ();
 sg13g2_decap_8 FILLER_78_1641 ();
 sg13g2_decap_8 FILLER_78_1648 ();
 sg13g2_decap_8 FILLER_78_1655 ();
 sg13g2_decap_8 FILLER_78_1662 ();
 sg13g2_decap_8 FILLER_78_1669 ();
 sg13g2_decap_8 FILLER_78_1676 ();
 sg13g2_decap_8 FILLER_78_1683 ();
 sg13g2_decap_8 FILLER_78_1690 ();
 sg13g2_decap_8 FILLER_78_1697 ();
 sg13g2_decap_8 FILLER_78_1704 ();
 sg13g2_decap_8 FILLER_78_1711 ();
 sg13g2_decap_8 FILLER_78_1718 ();
 sg13g2_decap_8 FILLER_78_1725 ();
 sg13g2_decap_8 FILLER_78_1732 ();
 sg13g2_decap_8 FILLER_78_1739 ();
 sg13g2_decap_8 FILLER_78_1746 ();
 sg13g2_decap_8 FILLER_78_1753 ();
 sg13g2_decap_8 FILLER_78_1760 ();
 sg13g2_fill_1 FILLER_78_1767 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_decap_8 FILLER_79_35 ();
 sg13g2_decap_8 FILLER_79_42 ();
 sg13g2_decap_8 FILLER_79_49 ();
 sg13g2_decap_4 FILLER_79_56 ();
 sg13g2_fill_2 FILLER_79_60 ();
 sg13g2_fill_2 FILLER_79_104 ();
 sg13g2_fill_1 FILLER_79_123 ();
 sg13g2_decap_8 FILLER_79_147 ();
 sg13g2_decap_8 FILLER_79_154 ();
 sg13g2_decap_8 FILLER_79_161 ();
 sg13g2_decap_8 FILLER_79_168 ();
 sg13g2_decap_8 FILLER_79_175 ();
 sg13g2_fill_2 FILLER_79_182 ();
 sg13g2_fill_2 FILLER_79_193 ();
 sg13g2_fill_1 FILLER_79_195 ();
 sg13g2_fill_2 FILLER_79_257 ();
 sg13g2_decap_8 FILLER_79_268 ();
 sg13g2_decap_8 FILLER_79_275 ();
 sg13g2_decap_8 FILLER_79_282 ();
 sg13g2_decap_8 FILLER_79_289 ();
 sg13g2_decap_8 FILLER_79_304 ();
 sg13g2_decap_8 FILLER_79_311 ();
 sg13g2_decap_8 FILLER_79_318 ();
 sg13g2_fill_2 FILLER_79_325 ();
 sg13g2_fill_2 FILLER_79_340 ();
 sg13g2_fill_1 FILLER_79_342 ();
 sg13g2_decap_8 FILLER_79_347 ();
 sg13g2_decap_4 FILLER_79_354 ();
 sg13g2_decap_8 FILLER_79_367 ();
 sg13g2_decap_8 FILLER_79_374 ();
 sg13g2_decap_8 FILLER_79_381 ();
 sg13g2_decap_8 FILLER_79_388 ();
 sg13g2_decap_8 FILLER_79_395 ();
 sg13g2_decap_8 FILLER_79_402 ();
 sg13g2_decap_8 FILLER_79_409 ();
 sg13g2_decap_8 FILLER_79_416 ();
 sg13g2_decap_8 FILLER_79_423 ();
 sg13g2_decap_8 FILLER_79_430 ();
 sg13g2_decap_8 FILLER_79_437 ();
 sg13g2_decap_8 FILLER_79_444 ();
 sg13g2_decap_8 FILLER_79_451 ();
 sg13g2_decap_8 FILLER_79_458 ();
 sg13g2_decap_8 FILLER_79_465 ();
 sg13g2_decap_8 FILLER_79_472 ();
 sg13g2_decap_8 FILLER_79_479 ();
 sg13g2_decap_8 FILLER_79_486 ();
 sg13g2_decap_8 FILLER_79_493 ();
 sg13g2_decap_8 FILLER_79_500 ();
 sg13g2_decap_8 FILLER_79_507 ();
 sg13g2_decap_8 FILLER_79_514 ();
 sg13g2_decap_8 FILLER_79_521 ();
 sg13g2_decap_8 FILLER_79_528 ();
 sg13g2_decap_8 FILLER_79_535 ();
 sg13g2_decap_8 FILLER_79_542 ();
 sg13g2_decap_8 FILLER_79_549 ();
 sg13g2_decap_8 FILLER_79_556 ();
 sg13g2_decap_8 FILLER_79_563 ();
 sg13g2_decap_8 FILLER_79_570 ();
 sg13g2_decap_8 FILLER_79_577 ();
 sg13g2_decap_8 FILLER_79_584 ();
 sg13g2_decap_8 FILLER_79_591 ();
 sg13g2_decap_8 FILLER_79_598 ();
 sg13g2_decap_8 FILLER_79_605 ();
 sg13g2_decap_8 FILLER_79_612 ();
 sg13g2_decap_8 FILLER_79_619 ();
 sg13g2_decap_8 FILLER_79_626 ();
 sg13g2_decap_8 FILLER_79_633 ();
 sg13g2_decap_8 FILLER_79_640 ();
 sg13g2_decap_8 FILLER_79_647 ();
 sg13g2_decap_8 FILLER_79_654 ();
 sg13g2_decap_8 FILLER_79_661 ();
 sg13g2_decap_8 FILLER_79_668 ();
 sg13g2_decap_8 FILLER_79_675 ();
 sg13g2_decap_8 FILLER_79_682 ();
 sg13g2_decap_8 FILLER_79_689 ();
 sg13g2_decap_8 FILLER_79_696 ();
 sg13g2_decap_8 FILLER_79_703 ();
 sg13g2_decap_8 FILLER_79_710 ();
 sg13g2_decap_8 FILLER_79_717 ();
 sg13g2_decap_8 FILLER_79_724 ();
 sg13g2_decap_8 FILLER_79_731 ();
 sg13g2_decap_8 FILLER_79_738 ();
 sg13g2_decap_8 FILLER_79_745 ();
 sg13g2_decap_8 FILLER_79_752 ();
 sg13g2_decap_8 FILLER_79_759 ();
 sg13g2_decap_8 FILLER_79_766 ();
 sg13g2_decap_8 FILLER_79_773 ();
 sg13g2_decap_8 FILLER_79_780 ();
 sg13g2_decap_8 FILLER_79_787 ();
 sg13g2_decap_8 FILLER_79_794 ();
 sg13g2_decap_8 FILLER_79_801 ();
 sg13g2_decap_8 FILLER_79_808 ();
 sg13g2_decap_8 FILLER_79_815 ();
 sg13g2_decap_8 FILLER_79_822 ();
 sg13g2_decap_8 FILLER_79_829 ();
 sg13g2_decap_8 FILLER_79_836 ();
 sg13g2_decap_8 FILLER_79_843 ();
 sg13g2_decap_8 FILLER_79_850 ();
 sg13g2_decap_8 FILLER_79_857 ();
 sg13g2_decap_8 FILLER_79_864 ();
 sg13g2_decap_8 FILLER_79_871 ();
 sg13g2_decap_8 FILLER_79_878 ();
 sg13g2_decap_8 FILLER_79_885 ();
 sg13g2_decap_8 FILLER_79_892 ();
 sg13g2_decap_8 FILLER_79_899 ();
 sg13g2_decap_8 FILLER_79_906 ();
 sg13g2_decap_8 FILLER_79_913 ();
 sg13g2_decap_8 FILLER_79_920 ();
 sg13g2_decap_8 FILLER_79_927 ();
 sg13g2_decap_8 FILLER_79_934 ();
 sg13g2_decap_8 FILLER_79_941 ();
 sg13g2_decap_8 FILLER_79_948 ();
 sg13g2_decap_8 FILLER_79_955 ();
 sg13g2_decap_8 FILLER_79_962 ();
 sg13g2_decap_8 FILLER_79_969 ();
 sg13g2_decap_8 FILLER_79_976 ();
 sg13g2_decap_8 FILLER_79_983 ();
 sg13g2_decap_8 FILLER_79_990 ();
 sg13g2_decap_8 FILLER_79_997 ();
 sg13g2_decap_8 FILLER_79_1004 ();
 sg13g2_decap_8 FILLER_79_1011 ();
 sg13g2_decap_8 FILLER_79_1018 ();
 sg13g2_decap_8 FILLER_79_1025 ();
 sg13g2_decap_8 FILLER_79_1032 ();
 sg13g2_decap_8 FILLER_79_1039 ();
 sg13g2_decap_8 FILLER_79_1046 ();
 sg13g2_decap_8 FILLER_79_1053 ();
 sg13g2_decap_8 FILLER_79_1060 ();
 sg13g2_decap_8 FILLER_79_1067 ();
 sg13g2_decap_8 FILLER_79_1074 ();
 sg13g2_decap_8 FILLER_79_1081 ();
 sg13g2_decap_8 FILLER_79_1088 ();
 sg13g2_decap_8 FILLER_79_1095 ();
 sg13g2_decap_8 FILLER_79_1102 ();
 sg13g2_decap_8 FILLER_79_1109 ();
 sg13g2_decap_8 FILLER_79_1116 ();
 sg13g2_decap_8 FILLER_79_1123 ();
 sg13g2_decap_8 FILLER_79_1130 ();
 sg13g2_decap_8 FILLER_79_1137 ();
 sg13g2_decap_8 FILLER_79_1144 ();
 sg13g2_decap_8 FILLER_79_1151 ();
 sg13g2_decap_8 FILLER_79_1158 ();
 sg13g2_decap_8 FILLER_79_1165 ();
 sg13g2_decap_8 FILLER_79_1172 ();
 sg13g2_decap_8 FILLER_79_1179 ();
 sg13g2_decap_8 FILLER_79_1186 ();
 sg13g2_decap_8 FILLER_79_1193 ();
 sg13g2_decap_8 FILLER_79_1200 ();
 sg13g2_decap_8 FILLER_79_1207 ();
 sg13g2_decap_8 FILLER_79_1214 ();
 sg13g2_decap_8 FILLER_79_1221 ();
 sg13g2_decap_8 FILLER_79_1228 ();
 sg13g2_decap_8 FILLER_79_1235 ();
 sg13g2_decap_8 FILLER_79_1242 ();
 sg13g2_decap_8 FILLER_79_1249 ();
 sg13g2_decap_8 FILLER_79_1256 ();
 sg13g2_decap_8 FILLER_79_1263 ();
 sg13g2_decap_8 FILLER_79_1270 ();
 sg13g2_decap_8 FILLER_79_1277 ();
 sg13g2_decap_8 FILLER_79_1284 ();
 sg13g2_decap_8 FILLER_79_1291 ();
 sg13g2_decap_8 FILLER_79_1298 ();
 sg13g2_decap_8 FILLER_79_1305 ();
 sg13g2_decap_8 FILLER_79_1312 ();
 sg13g2_decap_8 FILLER_79_1319 ();
 sg13g2_decap_8 FILLER_79_1326 ();
 sg13g2_decap_8 FILLER_79_1333 ();
 sg13g2_decap_8 FILLER_79_1340 ();
 sg13g2_decap_8 FILLER_79_1347 ();
 sg13g2_decap_8 FILLER_79_1354 ();
 sg13g2_decap_8 FILLER_79_1361 ();
 sg13g2_decap_8 FILLER_79_1368 ();
 sg13g2_decap_8 FILLER_79_1375 ();
 sg13g2_decap_8 FILLER_79_1382 ();
 sg13g2_decap_8 FILLER_79_1389 ();
 sg13g2_decap_8 FILLER_79_1396 ();
 sg13g2_decap_8 FILLER_79_1403 ();
 sg13g2_decap_8 FILLER_79_1410 ();
 sg13g2_decap_8 FILLER_79_1417 ();
 sg13g2_decap_8 FILLER_79_1424 ();
 sg13g2_decap_8 FILLER_79_1431 ();
 sg13g2_decap_8 FILLER_79_1438 ();
 sg13g2_decap_8 FILLER_79_1445 ();
 sg13g2_decap_8 FILLER_79_1452 ();
 sg13g2_decap_8 FILLER_79_1459 ();
 sg13g2_decap_8 FILLER_79_1466 ();
 sg13g2_decap_8 FILLER_79_1473 ();
 sg13g2_decap_8 FILLER_79_1480 ();
 sg13g2_decap_8 FILLER_79_1487 ();
 sg13g2_decap_8 FILLER_79_1494 ();
 sg13g2_decap_8 FILLER_79_1501 ();
 sg13g2_decap_8 FILLER_79_1508 ();
 sg13g2_decap_8 FILLER_79_1515 ();
 sg13g2_decap_8 FILLER_79_1522 ();
 sg13g2_decap_8 FILLER_79_1529 ();
 sg13g2_decap_8 FILLER_79_1536 ();
 sg13g2_decap_8 FILLER_79_1543 ();
 sg13g2_decap_8 FILLER_79_1550 ();
 sg13g2_decap_8 FILLER_79_1557 ();
 sg13g2_decap_8 FILLER_79_1564 ();
 sg13g2_decap_8 FILLER_79_1571 ();
 sg13g2_decap_8 FILLER_79_1578 ();
 sg13g2_decap_8 FILLER_79_1585 ();
 sg13g2_decap_8 FILLER_79_1592 ();
 sg13g2_decap_8 FILLER_79_1599 ();
 sg13g2_decap_8 FILLER_79_1606 ();
 sg13g2_decap_8 FILLER_79_1613 ();
 sg13g2_decap_8 FILLER_79_1620 ();
 sg13g2_decap_8 FILLER_79_1627 ();
 sg13g2_decap_8 FILLER_79_1634 ();
 sg13g2_decap_8 FILLER_79_1641 ();
 sg13g2_decap_8 FILLER_79_1648 ();
 sg13g2_decap_8 FILLER_79_1655 ();
 sg13g2_decap_8 FILLER_79_1662 ();
 sg13g2_decap_8 FILLER_79_1669 ();
 sg13g2_decap_8 FILLER_79_1676 ();
 sg13g2_decap_8 FILLER_79_1683 ();
 sg13g2_decap_8 FILLER_79_1690 ();
 sg13g2_decap_8 FILLER_79_1697 ();
 sg13g2_decap_8 FILLER_79_1704 ();
 sg13g2_decap_8 FILLER_79_1711 ();
 sg13g2_decap_8 FILLER_79_1718 ();
 sg13g2_decap_8 FILLER_79_1725 ();
 sg13g2_decap_8 FILLER_79_1732 ();
 sg13g2_decap_8 FILLER_79_1739 ();
 sg13g2_decap_8 FILLER_79_1746 ();
 sg13g2_decap_8 FILLER_79_1753 ();
 sg13g2_decap_8 FILLER_79_1760 ();
 sg13g2_fill_1 FILLER_79_1767 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_42 ();
 sg13g2_decap_8 FILLER_80_49 ();
 sg13g2_decap_4 FILLER_80_60 ();
 sg13g2_fill_2 FILLER_80_76 ();
 sg13g2_fill_2 FILLER_80_100 ();
 sg13g2_fill_1 FILLER_80_102 ();
 sg13g2_fill_2 FILLER_80_141 ();
 sg13g2_fill_1 FILLER_80_143 ();
 sg13g2_decap_4 FILLER_80_148 ();
 sg13g2_decap_4 FILLER_80_156 ();
 sg13g2_decap_4 FILLER_80_164 ();
 sg13g2_decap_4 FILLER_80_172 ();
 sg13g2_decap_8 FILLER_80_180 ();
 sg13g2_decap_8 FILLER_80_187 ();
 sg13g2_decap_8 FILLER_80_194 ();
 sg13g2_decap_4 FILLER_80_201 ();
 sg13g2_fill_2 FILLER_80_205 ();
 sg13g2_decap_8 FILLER_80_212 ();
 sg13g2_decap_8 FILLER_80_219 ();
 sg13g2_fill_2 FILLER_80_226 ();
 sg13g2_fill_1 FILLER_80_228 ();
 sg13g2_decap_8 FILLER_80_263 ();
 sg13g2_decap_8 FILLER_80_270 ();
 sg13g2_decap_8 FILLER_80_277 ();
 sg13g2_decap_8 FILLER_80_284 ();
 sg13g2_decap_8 FILLER_80_291 ();
 sg13g2_decap_4 FILLER_80_298 ();
 sg13g2_fill_2 FILLER_80_302 ();
 sg13g2_fill_2 FILLER_80_309 ();
 sg13g2_fill_1 FILLER_80_311 ();
 sg13g2_decap_8 FILLER_80_325 ();
 sg13g2_decap_8 FILLER_80_332 ();
 sg13g2_decap_8 FILLER_80_339 ();
 sg13g2_decap_8 FILLER_80_346 ();
 sg13g2_decap_8 FILLER_80_353 ();
 sg13g2_decap_8 FILLER_80_360 ();
 sg13g2_decap_8 FILLER_80_367 ();
 sg13g2_decap_8 FILLER_80_374 ();
 sg13g2_decap_8 FILLER_80_381 ();
 sg13g2_decap_8 FILLER_80_388 ();
 sg13g2_decap_8 FILLER_80_395 ();
 sg13g2_decap_8 FILLER_80_402 ();
 sg13g2_decap_8 FILLER_80_409 ();
 sg13g2_decap_8 FILLER_80_416 ();
 sg13g2_decap_8 FILLER_80_423 ();
 sg13g2_decap_8 FILLER_80_430 ();
 sg13g2_decap_8 FILLER_80_437 ();
 sg13g2_decap_8 FILLER_80_444 ();
 sg13g2_decap_8 FILLER_80_451 ();
 sg13g2_decap_8 FILLER_80_458 ();
 sg13g2_decap_8 FILLER_80_465 ();
 sg13g2_decap_8 FILLER_80_472 ();
 sg13g2_decap_8 FILLER_80_479 ();
 sg13g2_decap_8 FILLER_80_486 ();
 sg13g2_decap_8 FILLER_80_493 ();
 sg13g2_decap_8 FILLER_80_500 ();
 sg13g2_decap_8 FILLER_80_507 ();
 sg13g2_decap_8 FILLER_80_514 ();
 sg13g2_decap_8 FILLER_80_521 ();
 sg13g2_decap_8 FILLER_80_528 ();
 sg13g2_decap_8 FILLER_80_535 ();
 sg13g2_decap_8 FILLER_80_542 ();
 sg13g2_decap_8 FILLER_80_549 ();
 sg13g2_decap_8 FILLER_80_556 ();
 sg13g2_decap_8 FILLER_80_563 ();
 sg13g2_decap_8 FILLER_80_570 ();
 sg13g2_decap_8 FILLER_80_577 ();
 sg13g2_decap_8 FILLER_80_584 ();
 sg13g2_decap_8 FILLER_80_591 ();
 sg13g2_decap_8 FILLER_80_598 ();
 sg13g2_decap_8 FILLER_80_605 ();
 sg13g2_decap_8 FILLER_80_612 ();
 sg13g2_decap_8 FILLER_80_619 ();
 sg13g2_decap_8 FILLER_80_626 ();
 sg13g2_decap_8 FILLER_80_633 ();
 sg13g2_decap_8 FILLER_80_640 ();
 sg13g2_decap_8 FILLER_80_647 ();
 sg13g2_decap_8 FILLER_80_654 ();
 sg13g2_decap_8 FILLER_80_661 ();
 sg13g2_decap_8 FILLER_80_668 ();
 sg13g2_decap_8 FILLER_80_675 ();
 sg13g2_decap_8 FILLER_80_682 ();
 sg13g2_decap_8 FILLER_80_689 ();
 sg13g2_decap_8 FILLER_80_696 ();
 sg13g2_decap_8 FILLER_80_703 ();
 sg13g2_decap_8 FILLER_80_710 ();
 sg13g2_decap_8 FILLER_80_717 ();
 sg13g2_decap_8 FILLER_80_724 ();
 sg13g2_decap_8 FILLER_80_731 ();
 sg13g2_decap_8 FILLER_80_738 ();
 sg13g2_decap_8 FILLER_80_745 ();
 sg13g2_decap_8 FILLER_80_752 ();
 sg13g2_decap_8 FILLER_80_759 ();
 sg13g2_decap_8 FILLER_80_766 ();
 sg13g2_decap_8 FILLER_80_773 ();
 sg13g2_decap_8 FILLER_80_780 ();
 sg13g2_decap_8 FILLER_80_787 ();
 sg13g2_decap_8 FILLER_80_794 ();
 sg13g2_decap_8 FILLER_80_801 ();
 sg13g2_decap_8 FILLER_80_808 ();
 sg13g2_decap_8 FILLER_80_815 ();
 sg13g2_decap_8 FILLER_80_822 ();
 sg13g2_decap_8 FILLER_80_829 ();
 sg13g2_decap_8 FILLER_80_836 ();
 sg13g2_decap_8 FILLER_80_843 ();
 sg13g2_decap_8 FILLER_80_850 ();
 sg13g2_decap_8 FILLER_80_857 ();
 sg13g2_decap_8 FILLER_80_864 ();
 sg13g2_decap_8 FILLER_80_871 ();
 sg13g2_decap_8 FILLER_80_878 ();
 sg13g2_decap_8 FILLER_80_885 ();
 sg13g2_decap_8 FILLER_80_892 ();
 sg13g2_decap_8 FILLER_80_899 ();
 sg13g2_decap_8 FILLER_80_906 ();
 sg13g2_decap_8 FILLER_80_913 ();
 sg13g2_decap_8 FILLER_80_920 ();
 sg13g2_decap_8 FILLER_80_927 ();
 sg13g2_decap_8 FILLER_80_934 ();
 sg13g2_decap_8 FILLER_80_941 ();
 sg13g2_decap_8 FILLER_80_948 ();
 sg13g2_decap_8 FILLER_80_955 ();
 sg13g2_decap_8 FILLER_80_962 ();
 sg13g2_decap_8 FILLER_80_969 ();
 sg13g2_decap_8 FILLER_80_976 ();
 sg13g2_decap_8 FILLER_80_983 ();
 sg13g2_decap_8 FILLER_80_990 ();
 sg13g2_decap_8 FILLER_80_997 ();
 sg13g2_decap_8 FILLER_80_1004 ();
 sg13g2_decap_8 FILLER_80_1011 ();
 sg13g2_decap_8 FILLER_80_1018 ();
 sg13g2_decap_8 FILLER_80_1025 ();
 sg13g2_decap_8 FILLER_80_1032 ();
 sg13g2_decap_8 FILLER_80_1039 ();
 sg13g2_decap_8 FILLER_80_1046 ();
 sg13g2_decap_8 FILLER_80_1053 ();
 sg13g2_decap_8 FILLER_80_1060 ();
 sg13g2_decap_8 FILLER_80_1067 ();
 sg13g2_decap_8 FILLER_80_1074 ();
 sg13g2_decap_8 FILLER_80_1081 ();
 sg13g2_decap_8 FILLER_80_1088 ();
 sg13g2_decap_8 FILLER_80_1095 ();
 sg13g2_decap_8 FILLER_80_1102 ();
 sg13g2_decap_8 FILLER_80_1109 ();
 sg13g2_decap_8 FILLER_80_1116 ();
 sg13g2_decap_8 FILLER_80_1123 ();
 sg13g2_decap_8 FILLER_80_1130 ();
 sg13g2_decap_8 FILLER_80_1137 ();
 sg13g2_decap_8 FILLER_80_1144 ();
 sg13g2_decap_8 FILLER_80_1151 ();
 sg13g2_decap_8 FILLER_80_1158 ();
 sg13g2_decap_8 FILLER_80_1165 ();
 sg13g2_decap_8 FILLER_80_1172 ();
 sg13g2_decap_8 FILLER_80_1179 ();
 sg13g2_decap_8 FILLER_80_1186 ();
 sg13g2_decap_8 FILLER_80_1193 ();
 sg13g2_decap_8 FILLER_80_1200 ();
 sg13g2_decap_8 FILLER_80_1207 ();
 sg13g2_decap_8 FILLER_80_1214 ();
 sg13g2_decap_8 FILLER_80_1221 ();
 sg13g2_decap_8 FILLER_80_1228 ();
 sg13g2_decap_8 FILLER_80_1235 ();
 sg13g2_decap_8 FILLER_80_1242 ();
 sg13g2_decap_8 FILLER_80_1249 ();
 sg13g2_decap_8 FILLER_80_1256 ();
 sg13g2_decap_8 FILLER_80_1263 ();
 sg13g2_decap_8 FILLER_80_1270 ();
 sg13g2_decap_8 FILLER_80_1277 ();
 sg13g2_decap_8 FILLER_80_1284 ();
 sg13g2_decap_8 FILLER_80_1291 ();
 sg13g2_decap_8 FILLER_80_1298 ();
 sg13g2_decap_8 FILLER_80_1305 ();
 sg13g2_decap_8 FILLER_80_1312 ();
 sg13g2_decap_8 FILLER_80_1319 ();
 sg13g2_decap_8 FILLER_80_1326 ();
 sg13g2_decap_8 FILLER_80_1333 ();
 sg13g2_decap_8 FILLER_80_1340 ();
 sg13g2_decap_8 FILLER_80_1347 ();
 sg13g2_decap_8 FILLER_80_1354 ();
 sg13g2_decap_8 FILLER_80_1361 ();
 sg13g2_decap_8 FILLER_80_1368 ();
 sg13g2_decap_8 FILLER_80_1375 ();
 sg13g2_decap_8 FILLER_80_1382 ();
 sg13g2_decap_8 FILLER_80_1389 ();
 sg13g2_decap_8 FILLER_80_1396 ();
 sg13g2_decap_8 FILLER_80_1403 ();
 sg13g2_decap_8 FILLER_80_1410 ();
 sg13g2_decap_8 FILLER_80_1417 ();
 sg13g2_decap_8 FILLER_80_1424 ();
 sg13g2_decap_8 FILLER_80_1431 ();
 sg13g2_decap_8 FILLER_80_1438 ();
 sg13g2_decap_8 FILLER_80_1445 ();
 sg13g2_decap_8 FILLER_80_1452 ();
 sg13g2_decap_8 FILLER_80_1459 ();
 sg13g2_decap_8 FILLER_80_1466 ();
 sg13g2_decap_8 FILLER_80_1473 ();
 sg13g2_decap_8 FILLER_80_1480 ();
 sg13g2_decap_8 FILLER_80_1487 ();
 sg13g2_decap_8 FILLER_80_1494 ();
 sg13g2_decap_8 FILLER_80_1501 ();
 sg13g2_decap_8 FILLER_80_1508 ();
 sg13g2_decap_8 FILLER_80_1515 ();
 sg13g2_decap_8 FILLER_80_1522 ();
 sg13g2_decap_8 FILLER_80_1529 ();
 sg13g2_decap_8 FILLER_80_1536 ();
 sg13g2_decap_8 FILLER_80_1543 ();
 sg13g2_decap_8 FILLER_80_1550 ();
 sg13g2_decap_8 FILLER_80_1557 ();
 sg13g2_decap_8 FILLER_80_1564 ();
 sg13g2_decap_8 FILLER_80_1571 ();
 sg13g2_decap_8 FILLER_80_1578 ();
 sg13g2_decap_8 FILLER_80_1585 ();
 sg13g2_decap_8 FILLER_80_1592 ();
 sg13g2_decap_8 FILLER_80_1599 ();
 sg13g2_decap_8 FILLER_80_1606 ();
 sg13g2_decap_8 FILLER_80_1613 ();
 sg13g2_decap_8 FILLER_80_1620 ();
 sg13g2_decap_8 FILLER_80_1627 ();
 sg13g2_decap_8 FILLER_80_1634 ();
 sg13g2_decap_8 FILLER_80_1641 ();
 sg13g2_decap_8 FILLER_80_1648 ();
 sg13g2_decap_8 FILLER_80_1655 ();
 sg13g2_decap_8 FILLER_80_1662 ();
 sg13g2_decap_8 FILLER_80_1669 ();
 sg13g2_decap_8 FILLER_80_1676 ();
 sg13g2_decap_8 FILLER_80_1683 ();
 sg13g2_decap_8 FILLER_80_1690 ();
 sg13g2_decap_8 FILLER_80_1697 ();
 sg13g2_decap_8 FILLER_80_1704 ();
 sg13g2_decap_8 FILLER_80_1711 ();
 sg13g2_decap_8 FILLER_80_1718 ();
 sg13g2_decap_8 FILLER_80_1725 ();
 sg13g2_decap_8 FILLER_80_1732 ();
 sg13g2_decap_8 FILLER_80_1739 ();
 sg13g2_decap_8 FILLER_80_1746 ();
 sg13g2_decap_8 FILLER_80_1753 ();
 sg13g2_decap_8 FILLER_80_1760 ();
 sg13g2_fill_1 FILLER_80_1767 ();
 assign uio_oe[0] = net4;
 assign uio_oe[1] = net5;
 assign uio_oe[2] = net6;
 assign uio_oe[3] = net7;
 assign uio_oe[4] = net8;
 assign uio_oe[5] = net9;
 assign uio_oe[6] = net10;
 assign uio_oe[7] = net11;
 assign uio_out[0] = net12;
 assign uio_out[1] = net13;
 assign uio_out[2] = net14;
 assign uio_out[3] = net15;
 assign uio_out[4] = net16;
 assign uio_out[5] = net17;
 assign uio_out[6] = net18;
 assign uio_out[7] = net19;
endmodule

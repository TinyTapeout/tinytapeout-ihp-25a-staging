module tt_um_snn_with_delays_paolaunisa (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire MISO;
 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire _07353_;
 wire _07354_;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire _07421_;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire _07435_;
 wire _07436_;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire _07495_;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire _07515_;
 wire _07516_;
 wire _07517_;
 wire _07518_;
 wire _07519_;
 wire _07520_;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire _07524_;
 wire _07525_;
 wire _07526_;
 wire _07527_;
 wire _07528_;
 wire _07529_;
 wire _07530_;
 wire _07531_;
 wire _07532_;
 wire _07533_;
 wire _07534_;
 wire _07535_;
 wire _07536_;
 wire _07537_;
 wire _07538_;
 wire _07539_;
 wire _07540_;
 wire _07541_;
 wire _07542_;
 wire _07543_;
 wire _07544_;
 wire _07545_;
 wire _07546_;
 wire _07547_;
 wire _07548_;
 wire _07549_;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire _07557_;
 wire _07558_;
 wire _07559_;
 wire _07560_;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire _07565_;
 wire _07566_;
 wire _07567_;
 wire _07568_;
 wire _07569_;
 wire _07570_;
 wire _07571_;
 wire _07572_;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire _07576_;
 wire _07577_;
 wire _07578_;
 wire _07579_;
 wire _07580_;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire _07585_;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire _07589_;
 wire _07590_;
 wire _07591_;
 wire _07592_;
 wire _07593_;
 wire _07594_;
 wire _07595_;
 wire _07596_;
 wire _07597_;
 wire _07598_;
 wire _07599_;
 wire _07600_;
 wire _07601_;
 wire _07602_;
 wire _07603_;
 wire _07604_;
 wire _07605_;
 wire _07606_;
 wire _07607_;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire _07611_;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07615_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire _07620_;
 wire _07621_;
 wire _07622_;
 wire _07623_;
 wire _07624_;
 wire _07625_;
 wire _07626_;
 wire _07627_;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire _07631_;
 wire _07632_;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07636_;
 wire _07637_;
 wire _07638_;
 wire _07639_;
 wire _07640_;
 wire _07641_;
 wire _07642_;
 wire _07643_;
 wire _07644_;
 wire _07645_;
 wire _07646_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07656_;
 wire _07657_;
 wire _07658_;
 wire _07659_;
 wire _07660_;
 wire _07661_;
 wire _07662_;
 wire _07663_;
 wire _07664_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire _07672_;
 wire _07673_;
 wire _07674_;
 wire _07675_;
 wire _07676_;
 wire _07677_;
 wire _07678_;
 wire _07679_;
 wire _07680_;
 wire _07681_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07686_;
 wire _07687_;
 wire _07688_;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire _07693_;
 wire _07694_;
 wire _07695_;
 wire _07696_;
 wire _07697_;
 wire _07698_;
 wire _07699_;
 wire _07700_;
 wire _07701_;
 wire _07702_;
 wire _07703_;
 wire _07704_;
 wire _07705_;
 wire _07706_;
 wire _07707_;
 wire _07708_;
 wire _07709_;
 wire _07710_;
 wire _07711_;
 wire _07712_;
 wire _07713_;
 wire _07714_;
 wire _07715_;
 wire _07716_;
 wire _07717_;
 wire _07718_;
 wire _07719_;
 wire _07720_;
 wire _07721_;
 wire _07722_;
 wire _07723_;
 wire _07724_;
 wire _07725_;
 wire _07726_;
 wire _07727_;
 wire _07728_;
 wire _07729_;
 wire _07730_;
 wire _07731_;
 wire _07732_;
 wire _07733_;
 wire _07734_;
 wire _07735_;
 wire _07736_;
 wire _07737_;
 wire _07738_;
 wire _07739_;
 wire _07740_;
 wire _07741_;
 wire _07742_;
 wire _07743_;
 wire _07744_;
 wire _07745_;
 wire _07746_;
 wire _07747_;
 wire _07748_;
 wire _07749_;
 wire _07750_;
 wire _07751_;
 wire _07752_;
 wire _07753_;
 wire _07754_;
 wire _07755_;
 wire _07756_;
 wire _07757_;
 wire _07758_;
 wire _07759_;
 wire _07760_;
 wire _07761_;
 wire _07762_;
 wire _07763_;
 wire _07764_;
 wire _07765_;
 wire _07766_;
 wire _07767_;
 wire _07768_;
 wire _07769_;
 wire _07770_;
 wire _07771_;
 wire _07772_;
 wire _07773_;
 wire _07774_;
 wire _07775_;
 wire _07776_;
 wire _07777_;
 wire _07778_;
 wire _07779_;
 wire _07780_;
 wire _07781_;
 wire _07782_;
 wire _07783_;
 wire _07784_;
 wire _07785_;
 wire _07786_;
 wire _07787_;
 wire _07788_;
 wire _07789_;
 wire _07790_;
 wire _07791_;
 wire _07792_;
 wire _07793_;
 wire _07794_;
 wire _07795_;
 wire _07796_;
 wire _07797_;
 wire _07798_;
 wire _07799_;
 wire _07800_;
 wire _07801_;
 wire _07802_;
 wire _07803_;
 wire _07804_;
 wire _07805_;
 wire _07806_;
 wire _07807_;
 wire _07808_;
 wire _07809_;
 wire _07810_;
 wire _07811_;
 wire _07812_;
 wire _07813_;
 wire _07814_;
 wire _07815_;
 wire _07816_;
 wire _07817_;
 wire _07818_;
 wire _07819_;
 wire _07820_;
 wire _07821_;
 wire _07822_;
 wire _07823_;
 wire _07824_;
 wire _07825_;
 wire _07826_;
 wire _07827_;
 wire _07828_;
 wire _07829_;
 wire _07830_;
 wire _07831_;
 wire _07832_;
 wire _07833_;
 wire _07834_;
 wire _07835_;
 wire _07836_;
 wire _07837_;
 wire _07838_;
 wire _07839_;
 wire _07840_;
 wire _07841_;
 wire _07842_;
 wire _07843_;
 wire _07844_;
 wire _07845_;
 wire _07846_;
 wire _07847_;
 wire _07848_;
 wire _07849_;
 wire _07850_;
 wire _07851_;
 wire _07852_;
 wire _07853_;
 wire _07854_;
 wire _07855_;
 wire _07856_;
 wire _07857_;
 wire _07858_;
 wire _07859_;
 wire _07860_;
 wire _07861_;
 wire _07862_;
 wire _07863_;
 wire _07864_;
 wire _07865_;
 wire _07866_;
 wire _07867_;
 wire _07868_;
 wire _07869_;
 wire _07870_;
 wire _07871_;
 wire _07872_;
 wire _07873_;
 wire _07874_;
 wire _07875_;
 wire _07876_;
 wire _07877_;
 wire _07878_;
 wire _07879_;
 wire _07880_;
 wire _07881_;
 wire _07882_;
 wire _07883_;
 wire _07884_;
 wire _07885_;
 wire _07886_;
 wire _07887_;
 wire _07888_;
 wire _07889_;
 wire _07890_;
 wire _07891_;
 wire _07892_;
 wire _07893_;
 wire _07894_;
 wire _07895_;
 wire _07896_;
 wire _07897_;
 wire _07898_;
 wire _07899_;
 wire _07900_;
 wire _07901_;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire _07905_;
 wire _07906_;
 wire _07907_;
 wire _07908_;
 wire _07909_;
 wire _07910_;
 wire _07911_;
 wire _07912_;
 wire _07913_;
 wire _07914_;
 wire _07915_;
 wire _07916_;
 wire _07917_;
 wire _07918_;
 wire _07919_;
 wire _07920_;
 wire _07921_;
 wire _07922_;
 wire _07923_;
 wire _07924_;
 wire _07925_;
 wire _07926_;
 wire _07927_;
 wire _07928_;
 wire _07929_;
 wire _07930_;
 wire _07931_;
 wire _07932_;
 wire _07933_;
 wire _07934_;
 wire _07935_;
 wire _07936_;
 wire _07937_;
 wire _07938_;
 wire _07939_;
 wire _07940_;
 wire _07941_;
 wire _07942_;
 wire _07943_;
 wire _07944_;
 wire _07945_;
 wire _07946_;
 wire _07947_;
 wire _07948_;
 wire _07949_;
 wire _07950_;
 wire _07951_;
 wire _07952_;
 wire _07953_;
 wire _07954_;
 wire _07955_;
 wire _07956_;
 wire _07957_;
 wire _07958_;
 wire _07959_;
 wire _07960_;
 wire _07961_;
 wire _07962_;
 wire _07963_;
 wire _07964_;
 wire _07965_;
 wire _07966_;
 wire _07967_;
 wire _07968_;
 wire _07969_;
 wire _07970_;
 wire _07971_;
 wire _07972_;
 wire _07973_;
 wire _07974_;
 wire _07975_;
 wire _07976_;
 wire _07977_;
 wire _07978_;
 wire _07979_;
 wire _07980_;
 wire _07981_;
 wire _07982_;
 wire _07983_;
 wire _07984_;
 wire _07985_;
 wire _07986_;
 wire _07987_;
 wire _07988_;
 wire _07989_;
 wire _07990_;
 wire _07991_;
 wire _07992_;
 wire _07993_;
 wire _07994_;
 wire _07995_;
 wire _07996_;
 wire _07997_;
 wire _07998_;
 wire _07999_;
 wire _08000_;
 wire _08001_;
 wire _08002_;
 wire _08003_;
 wire _08004_;
 wire _08005_;
 wire _08006_;
 wire _08007_;
 wire _08008_;
 wire _08009_;
 wire _08010_;
 wire _08011_;
 wire _08012_;
 wire _08013_;
 wire _08014_;
 wire _08015_;
 wire _08016_;
 wire _08017_;
 wire _08018_;
 wire _08019_;
 wire _08020_;
 wire _08021_;
 wire _08022_;
 wire _08023_;
 wire _08024_;
 wire _08025_;
 wire _08026_;
 wire _08027_;
 wire _08028_;
 wire _08029_;
 wire _08030_;
 wire _08031_;
 wire _08032_;
 wire _08033_;
 wire _08034_;
 wire _08035_;
 wire _08036_;
 wire _08037_;
 wire _08038_;
 wire _08039_;
 wire _08040_;
 wire _08041_;
 wire _08042_;
 wire _08043_;
 wire _08044_;
 wire _08045_;
 wire _08046_;
 wire _08047_;
 wire _08048_;
 wire _08049_;
 wire _08050_;
 wire _08051_;
 wire _08052_;
 wire _08053_;
 wire _08054_;
 wire _08055_;
 wire _08056_;
 wire _08057_;
 wire _08058_;
 wire _08059_;
 wire _08060_;
 wire _08061_;
 wire _08062_;
 wire _08063_;
 wire _08064_;
 wire _08065_;
 wire _08066_;
 wire _08067_;
 wire _08068_;
 wire _08069_;
 wire _08070_;
 wire _08071_;
 wire _08072_;
 wire _08073_;
 wire _08074_;
 wire _08075_;
 wire _08076_;
 wire _08077_;
 wire _08078_;
 wire _08079_;
 wire _08080_;
 wire _08081_;
 wire _08082_;
 wire _08083_;
 wire _08084_;
 wire _08085_;
 wire _08086_;
 wire _08087_;
 wire _08088_;
 wire _08089_;
 wire _08090_;
 wire _08091_;
 wire _08092_;
 wire _08093_;
 wire _08094_;
 wire _08095_;
 wire _08096_;
 wire _08097_;
 wire _08098_;
 wire _08099_;
 wire _08100_;
 wire _08101_;
 wire _08102_;
 wire _08103_;
 wire _08104_;
 wire _08105_;
 wire _08106_;
 wire _08107_;
 wire _08108_;
 wire _08109_;
 wire _08110_;
 wire _08111_;
 wire _08112_;
 wire _08113_;
 wire _08114_;
 wire _08115_;
 wire _08116_;
 wire _08117_;
 wire _08118_;
 wire _08119_;
 wire _08120_;
 wire _08121_;
 wire _08122_;
 wire _08123_;
 wire _08124_;
 wire _08125_;
 wire _08126_;
 wire _08127_;
 wire _08128_;
 wire _08129_;
 wire _08130_;
 wire _08131_;
 wire _08132_;
 wire _08133_;
 wire _08134_;
 wire _08135_;
 wire _08136_;
 wire _08137_;
 wire _08138_;
 wire _08139_;
 wire _08140_;
 wire _08141_;
 wire _08142_;
 wire _08143_;
 wire _08144_;
 wire _08145_;
 wire _08146_;
 wire _08147_;
 wire _08148_;
 wire _08149_;
 wire _08150_;
 wire _08151_;
 wire _08152_;
 wire _08153_;
 wire _08154_;
 wire _08155_;
 wire _08156_;
 wire _08157_;
 wire _08158_;
 wire _08159_;
 wire _08160_;
 wire _08161_;
 wire _08162_;
 wire _08163_;
 wire _08164_;
 wire _08165_;
 wire _08166_;
 wire _08167_;
 wire _08168_;
 wire _08169_;
 wire _08170_;
 wire _08171_;
 wire _08172_;
 wire _08173_;
 wire _08174_;
 wire _08175_;
 wire _08176_;
 wire _08177_;
 wire _08178_;
 wire _08179_;
 wire _08180_;
 wire _08181_;
 wire _08182_;
 wire _08183_;
 wire _08184_;
 wire _08185_;
 wire _08186_;
 wire _08187_;
 wire _08188_;
 wire _08189_;
 wire _08190_;
 wire _08191_;
 wire _08192_;
 wire _08193_;
 wire _08194_;
 wire _08195_;
 wire _08196_;
 wire _08197_;
 wire _08198_;
 wire _08199_;
 wire _08200_;
 wire _08201_;
 wire _08202_;
 wire _08203_;
 wire _08204_;
 wire _08205_;
 wire _08206_;
 wire _08207_;
 wire _08208_;
 wire _08209_;
 wire _08210_;
 wire _08211_;
 wire _08212_;
 wire _08213_;
 wire _08214_;
 wire _08215_;
 wire _08216_;
 wire _08217_;
 wire _08218_;
 wire _08219_;
 wire _08220_;
 wire _08221_;
 wire _08222_;
 wire _08223_;
 wire _08224_;
 wire _08225_;
 wire _08226_;
 wire _08227_;
 wire _08228_;
 wire _08229_;
 wire _08230_;
 wire _08231_;
 wire _08232_;
 wire _08233_;
 wire _08234_;
 wire _08235_;
 wire _08236_;
 wire _08237_;
 wire _08238_;
 wire _08239_;
 wire _08240_;
 wire _08241_;
 wire _08242_;
 wire _08243_;
 wire _08244_;
 wire _08245_;
 wire _08246_;
 wire _08247_;
 wire _08248_;
 wire _08249_;
 wire _08250_;
 wire _08251_;
 wire _08252_;
 wire _08253_;
 wire _08254_;
 wire _08255_;
 wire _08256_;
 wire _08257_;
 wire _08258_;
 wire _08259_;
 wire _08260_;
 wire _08261_;
 wire _08262_;
 wire _08263_;
 wire _08264_;
 wire _08265_;
 wire _08266_;
 wire _08267_;
 wire _08268_;
 wire _08269_;
 wire _08270_;
 wire _08271_;
 wire _08272_;
 wire _08273_;
 wire _08274_;
 wire _08275_;
 wire _08276_;
 wire _08277_;
 wire _08278_;
 wire _08279_;
 wire _08280_;
 wire _08281_;
 wire _08282_;
 wire _08283_;
 wire _08284_;
 wire _08285_;
 wire _08286_;
 wire _08287_;
 wire _08288_;
 wire _08289_;
 wire _08290_;
 wire _08291_;
 wire _08292_;
 wire _08293_;
 wire _08294_;
 wire _08295_;
 wire _08296_;
 wire _08297_;
 wire _08298_;
 wire _08299_;
 wire _08300_;
 wire _08301_;
 wire _08302_;
 wire _08303_;
 wire _08304_;
 wire _08305_;
 wire _08306_;
 wire _08307_;
 wire _08308_;
 wire _08309_;
 wire _08310_;
 wire _08311_;
 wire _08312_;
 wire _08313_;
 wire _08314_;
 wire _08315_;
 wire _08316_;
 wire _08317_;
 wire _08318_;
 wire _08319_;
 wire _08320_;
 wire _08321_;
 wire _08322_;
 wire _08323_;
 wire _08324_;
 wire _08325_;
 wire _08326_;
 wire _08327_;
 wire _08328_;
 wire _08329_;
 wire _08330_;
 wire _08331_;
 wire _08332_;
 wire _08333_;
 wire _08334_;
 wire _08335_;
 wire _08336_;
 wire _08337_;
 wire _08338_;
 wire _08339_;
 wire _08340_;
 wire _08341_;
 wire _08342_;
 wire _08343_;
 wire _08344_;
 wire _08345_;
 wire _08346_;
 wire _08347_;
 wire _08348_;
 wire _08349_;
 wire _08350_;
 wire _08351_;
 wire _08352_;
 wire _08353_;
 wire _08354_;
 wire _08355_;
 wire _08356_;
 wire _08357_;
 wire _08358_;
 wire _08359_;
 wire _08360_;
 wire _08361_;
 wire _08362_;
 wire _08363_;
 wire _08364_;
 wire _08365_;
 wire _08366_;
 wire _08367_;
 wire _08368_;
 wire _08369_;
 wire _08370_;
 wire _08371_;
 wire _08372_;
 wire _08373_;
 wire _08374_;
 wire _08375_;
 wire _08376_;
 wire _08377_;
 wire _08378_;
 wire _08379_;
 wire _08380_;
 wire _08381_;
 wire _08382_;
 wire _08383_;
 wire _08384_;
 wire _08385_;
 wire _08386_;
 wire _08387_;
 wire _08388_;
 wire _08389_;
 wire _08390_;
 wire _08391_;
 wire _08392_;
 wire _08393_;
 wire _08394_;
 wire _08395_;
 wire _08396_;
 wire _08397_;
 wire _08398_;
 wire _08399_;
 wire _08400_;
 wire _08401_;
 wire _08402_;
 wire _08403_;
 wire _08404_;
 wire _08405_;
 wire _08406_;
 wire _08407_;
 wire _08408_;
 wire _08409_;
 wire _08410_;
 wire _08411_;
 wire _08412_;
 wire _08413_;
 wire _08414_;
 wire _08415_;
 wire _08416_;
 wire _08417_;
 wire _08418_;
 wire _08419_;
 wire _08420_;
 wire _08421_;
 wire _08422_;
 wire _08423_;
 wire _08424_;
 wire _08425_;
 wire _08426_;
 wire _08427_;
 wire _08428_;
 wire _08429_;
 wire _08430_;
 wire _08431_;
 wire _08432_;
 wire _08433_;
 wire _08434_;
 wire _08435_;
 wire _08436_;
 wire _08437_;
 wire _08438_;
 wire _08439_;
 wire _08440_;
 wire _08441_;
 wire _08442_;
 wire _08443_;
 wire _08444_;
 wire _08445_;
 wire _08446_;
 wire _08447_;
 wire _08448_;
 wire _08449_;
 wire _08450_;
 wire _08451_;
 wire _08452_;
 wire _08453_;
 wire _08454_;
 wire _08455_;
 wire _08456_;
 wire _08457_;
 wire _08458_;
 wire _08459_;
 wire _08460_;
 wire _08461_;
 wire _08462_;
 wire _08463_;
 wire _08464_;
 wire _08465_;
 wire _08466_;
 wire _08467_;
 wire _08468_;
 wire _08469_;
 wire _08470_;
 wire _08471_;
 wire _08472_;
 wire _08473_;
 wire _08474_;
 wire _08475_;
 wire _08476_;
 wire _08477_;
 wire _08478_;
 wire _08479_;
 wire _08480_;
 wire _08481_;
 wire _08482_;
 wire _08483_;
 wire _08484_;
 wire _08485_;
 wire _08486_;
 wire _08487_;
 wire _08488_;
 wire _08489_;
 wire _08490_;
 wire _08491_;
 wire _08492_;
 wire _08493_;
 wire _08494_;
 wire _08495_;
 wire _08496_;
 wire _08497_;
 wire _08498_;
 wire _08499_;
 wire _08500_;
 wire _08501_;
 wire _08502_;
 wire _08503_;
 wire _08504_;
 wire _08505_;
 wire _08506_;
 wire _08507_;
 wire _08508_;
 wire _08509_;
 wire _08510_;
 wire _08511_;
 wire _08512_;
 wire _08513_;
 wire _08514_;
 wire _08515_;
 wire _08516_;
 wire _08517_;
 wire _08518_;
 wire _08519_;
 wire _08520_;
 wire _08521_;
 wire _08522_;
 wire _08523_;
 wire _08524_;
 wire _08525_;
 wire _08526_;
 wire _08527_;
 wire _08528_;
 wire _08529_;
 wire _08530_;
 wire _08531_;
 wire _08532_;
 wire _08533_;
 wire _08534_;
 wire _08535_;
 wire _08536_;
 wire _08537_;
 wire _08538_;
 wire _08539_;
 wire _08540_;
 wire _08541_;
 wire _08542_;
 wire _08543_;
 wire _08544_;
 wire _08545_;
 wire _08546_;
 wire _08547_;
 wire _08548_;
 wire _08549_;
 wire _08550_;
 wire _08551_;
 wire _08552_;
 wire _08553_;
 wire _08554_;
 wire _08555_;
 wire _08556_;
 wire _08557_;
 wire _08558_;
 wire _08559_;
 wire _08560_;
 wire _08561_;
 wire _08562_;
 wire _08563_;
 wire _08564_;
 wire _08565_;
 wire _08566_;
 wire _08567_;
 wire _08568_;
 wire _08569_;
 wire _08570_;
 wire _08571_;
 wire _08572_;
 wire _08573_;
 wire _08574_;
 wire _08575_;
 wire _08576_;
 wire _08577_;
 wire _08578_;
 wire _08579_;
 wire _08580_;
 wire _08581_;
 wire _08582_;
 wire _08583_;
 wire _08584_;
 wire _08585_;
 wire _08586_;
 wire _08587_;
 wire _08588_;
 wire _08589_;
 wire _08590_;
 wire _08591_;
 wire _08592_;
 wire _08593_;
 wire _08594_;
 wire _08595_;
 wire _08596_;
 wire _08597_;
 wire _08598_;
 wire _08599_;
 wire _08600_;
 wire _08601_;
 wire _08602_;
 wire _08603_;
 wire _08604_;
 wire _08605_;
 wire _08606_;
 wire _08607_;
 wire _08608_;
 wire _08609_;
 wire _08610_;
 wire _08611_;
 wire _08612_;
 wire _08613_;
 wire _08614_;
 wire _08615_;
 wire _08616_;
 wire _08617_;
 wire _08618_;
 wire _08619_;
 wire _08620_;
 wire _08621_;
 wire _08622_;
 wire _08623_;
 wire _08624_;
 wire _08625_;
 wire _08626_;
 wire _08627_;
 wire _08628_;
 wire _08629_;
 wire _08630_;
 wire _08631_;
 wire _08632_;
 wire _08633_;
 wire _08634_;
 wire _08635_;
 wire _08636_;
 wire _08637_;
 wire _08638_;
 wire _08639_;
 wire _08640_;
 wire _08641_;
 wire _08642_;
 wire _08643_;
 wire _08644_;
 wire _08645_;
 wire _08646_;
 wire _08647_;
 wire _08648_;
 wire _08649_;
 wire _08650_;
 wire _08651_;
 wire _08652_;
 wire _08653_;
 wire _08654_;
 wire _08655_;
 wire _08656_;
 wire _08657_;
 wire _08658_;
 wire _08659_;
 wire _08660_;
 wire _08661_;
 wire _08662_;
 wire _08663_;
 wire _08664_;
 wire _08665_;
 wire _08666_;
 wire _08667_;
 wire _08668_;
 wire _08669_;
 wire _08670_;
 wire _08671_;
 wire _08672_;
 wire _08673_;
 wire _08674_;
 wire _08675_;
 wire _08676_;
 wire _08677_;
 wire _08678_;
 wire _08679_;
 wire _08680_;
 wire _08681_;
 wire _08682_;
 wire _08683_;
 wire _08684_;
 wire _08685_;
 wire _08686_;
 wire _08687_;
 wire _08688_;
 wire _08689_;
 wire _08690_;
 wire _08691_;
 wire _08692_;
 wire _08693_;
 wire _08694_;
 wire _08695_;
 wire _08696_;
 wire _08697_;
 wire _08698_;
 wire _08699_;
 wire _08700_;
 wire _08701_;
 wire _08702_;
 wire _08703_;
 wire _08704_;
 wire _08705_;
 wire _08706_;
 wire _08707_;
 wire _08708_;
 wire _08709_;
 wire _08710_;
 wire _08711_;
 wire _08712_;
 wire _08713_;
 wire _08714_;
 wire _08715_;
 wire _08716_;
 wire _08717_;
 wire _08718_;
 wire _08719_;
 wire _08720_;
 wire _08721_;
 wire _08722_;
 wire _08723_;
 wire _08724_;
 wire _08725_;
 wire _08726_;
 wire _08727_;
 wire _08728_;
 wire _08729_;
 wire _08730_;
 wire _08731_;
 wire _08732_;
 wire _08733_;
 wire _08734_;
 wire _08735_;
 wire _08736_;
 wire _08737_;
 wire _08738_;
 wire _08739_;
 wire _08740_;
 wire _08741_;
 wire _08742_;
 wire _08743_;
 wire _08744_;
 wire _08745_;
 wire _08746_;
 wire _08747_;
 wire _08748_;
 wire _08749_;
 wire _08750_;
 wire _08751_;
 wire _08752_;
 wire _08753_;
 wire _08754_;
 wire _08755_;
 wire _08756_;
 wire _08757_;
 wire _08758_;
 wire _08759_;
 wire _08760_;
 wire _08761_;
 wire _08762_;
 wire _08763_;
 wire _08764_;
 wire _08765_;
 wire _08766_;
 wire _08767_;
 wire _08768_;
 wire _08769_;
 wire _08770_;
 wire _08771_;
 wire _08772_;
 wire _08773_;
 wire _08774_;
 wire _08775_;
 wire _08776_;
 wire _08777_;
 wire _08778_;
 wire _08779_;
 wire _08780_;
 wire _08781_;
 wire _08782_;
 wire _08783_;
 wire _08784_;
 wire _08785_;
 wire _08786_;
 wire _08787_;
 wire _08788_;
 wire _08789_;
 wire _08790_;
 wire _08791_;
 wire _08792_;
 wire _08793_;
 wire _08794_;
 wire _08795_;
 wire _08796_;
 wire _08797_;
 wire _08798_;
 wire _08799_;
 wire _08800_;
 wire _08801_;
 wire _08802_;
 wire _08803_;
 wire _08804_;
 wire _08805_;
 wire _08806_;
 wire _08807_;
 wire _08808_;
 wire _08809_;
 wire _08810_;
 wire _08811_;
 wire _08812_;
 wire _08813_;
 wire _08814_;
 wire _08815_;
 wire _08816_;
 wire _08817_;
 wire _08818_;
 wire _08819_;
 wire _08820_;
 wire _08821_;
 wire _08822_;
 wire _08823_;
 wire _08824_;
 wire _08825_;
 wire _08826_;
 wire _08827_;
 wire _08828_;
 wire _08829_;
 wire _08830_;
 wire _08831_;
 wire _08832_;
 wire _08833_;
 wire _08834_;
 wire _08835_;
 wire _08836_;
 wire _08837_;
 wire _08838_;
 wire _08839_;
 wire _08840_;
 wire _08841_;
 wire _08842_;
 wire _08843_;
 wire _08844_;
 wire _08845_;
 wire _08846_;
 wire _08847_;
 wire _08848_;
 wire _08849_;
 wire _08850_;
 wire _08851_;
 wire _08852_;
 wire _08853_;
 wire _08854_;
 wire _08855_;
 wire _08856_;
 wire _08857_;
 wire _08858_;
 wire _08859_;
 wire _08860_;
 wire _08861_;
 wire _08862_;
 wire _08863_;
 wire _08864_;
 wire _08865_;
 wire _08866_;
 wire _08867_;
 wire _08868_;
 wire _08869_;
 wire _08870_;
 wire _08871_;
 wire _08872_;
 wire _08873_;
 wire _08874_;
 wire _08875_;
 wire _08876_;
 wire _08877_;
 wire _08878_;
 wire _08879_;
 wire _08880_;
 wire _08881_;
 wire _08882_;
 wire _08883_;
 wire _08884_;
 wire _08885_;
 wire _08886_;
 wire _08887_;
 wire _08888_;
 wire _08889_;
 wire _08890_;
 wire _08891_;
 wire _08892_;
 wire _08893_;
 wire _08894_;
 wire _08895_;
 wire _08896_;
 wire _08897_;
 wire _08898_;
 wire _08899_;
 wire _08900_;
 wire _08901_;
 wire _08902_;
 wire _08903_;
 wire _08904_;
 wire _08905_;
 wire _08906_;
 wire _08907_;
 wire _08908_;
 wire _08909_;
 wire _08910_;
 wire _08911_;
 wire _08912_;
 wire _08913_;
 wire _08914_;
 wire _08915_;
 wire _08916_;
 wire _08917_;
 wire _08918_;
 wire _08919_;
 wire _08920_;
 wire _08921_;
 wire _08922_;
 wire _08923_;
 wire _08924_;
 wire _08925_;
 wire _08926_;
 wire _08927_;
 wire _08928_;
 wire _08929_;
 wire _08930_;
 wire _08931_;
 wire _08932_;
 wire _08933_;
 wire _08934_;
 wire _08935_;
 wire _08936_;
 wire _08937_;
 wire _08938_;
 wire _08939_;
 wire _08940_;
 wire _08941_;
 wire _08942_;
 wire _08943_;
 wire _08944_;
 wire _08945_;
 wire _08946_;
 wire _08947_;
 wire _08948_;
 wire _08949_;
 wire _08950_;
 wire _08951_;
 wire _08952_;
 wire _08953_;
 wire _08954_;
 wire _08955_;
 wire _08956_;
 wire _08957_;
 wire _08958_;
 wire _08959_;
 wire _08960_;
 wire _08961_;
 wire _08962_;
 wire _08963_;
 wire _08964_;
 wire _08965_;
 wire _08966_;
 wire _08967_;
 wire _08968_;
 wire _08969_;
 wire _08970_;
 wire _08971_;
 wire _08972_;
 wire _08973_;
 wire _08974_;
 wire _08975_;
 wire _08976_;
 wire _08977_;
 wire _08978_;
 wire _08979_;
 wire _08980_;
 wire _08981_;
 wire _08982_;
 wire _08983_;
 wire _08984_;
 wire _08985_;
 wire _08986_;
 wire _08987_;
 wire _08988_;
 wire _08989_;
 wire _08990_;
 wire _08991_;
 wire _08992_;
 wire _08993_;
 wire _08994_;
 wire _08995_;
 wire _08996_;
 wire _08997_;
 wire _08998_;
 wire _08999_;
 wire _09000_;
 wire _09001_;
 wire _09002_;
 wire _09003_;
 wire _09004_;
 wire _09005_;
 wire _09006_;
 wire _09007_;
 wire _09008_;
 wire _09009_;
 wire _09010_;
 wire _09011_;
 wire _09012_;
 wire _09013_;
 wire _09014_;
 wire _09015_;
 wire _09016_;
 wire _09017_;
 wire _09018_;
 wire _09019_;
 wire _09020_;
 wire _09021_;
 wire _09022_;
 wire _09023_;
 wire _09024_;
 wire _09025_;
 wire _09026_;
 wire _09027_;
 wire _09028_;
 wire _09029_;
 wire _09030_;
 wire _09031_;
 wire _09032_;
 wire _09033_;
 wire _09034_;
 wire _09035_;
 wire _09036_;
 wire _09037_;
 wire _09038_;
 wire _09039_;
 wire _09040_;
 wire _09041_;
 wire _09042_;
 wire _09043_;
 wire _09044_;
 wire _09045_;
 wire _09046_;
 wire _09047_;
 wire _09048_;
 wire _09049_;
 wire _09050_;
 wire _09051_;
 wire _09052_;
 wire _09053_;
 wire _09054_;
 wire _09055_;
 wire _09056_;
 wire _09057_;
 wire _09058_;
 wire _09059_;
 wire _09060_;
 wire _09061_;
 wire _09062_;
 wire _09063_;
 wire _09064_;
 wire _09065_;
 wire _09066_;
 wire _09067_;
 wire _09068_;
 wire _09069_;
 wire _09070_;
 wire _09071_;
 wire _09072_;
 wire _09073_;
 wire _09074_;
 wire _09075_;
 wire _09076_;
 wire _09077_;
 wire _09078_;
 wire _09079_;
 wire _09080_;
 wire _09081_;
 wire _09082_;
 wire _09083_;
 wire _09084_;
 wire _09085_;
 wire _09086_;
 wire _09087_;
 wire _09088_;
 wire _09089_;
 wire _09090_;
 wire _09091_;
 wire _09092_;
 wire _09093_;
 wire _09094_;
 wire _09095_;
 wire _09096_;
 wire _09097_;
 wire _09098_;
 wire _09099_;
 wire _09100_;
 wire _09101_;
 wire _09102_;
 wire _09103_;
 wire _09104_;
 wire _09105_;
 wire _09106_;
 wire _09107_;
 wire _09108_;
 wire _09109_;
 wire _09110_;
 wire _09111_;
 wire _09112_;
 wire _09113_;
 wire _09114_;
 wire _09115_;
 wire _09116_;
 wire _09117_;
 wire _09118_;
 wire _09119_;
 wire _09120_;
 wire _09121_;
 wire _09122_;
 wire _09123_;
 wire _09124_;
 wire _09125_;
 wire _09126_;
 wire _09127_;
 wire _09128_;
 wire _09129_;
 wire _09130_;
 wire _09131_;
 wire _09132_;
 wire _09133_;
 wire _09134_;
 wire _09135_;
 wire _09136_;
 wire _09137_;
 wire _09138_;
 wire _09139_;
 wire _09140_;
 wire _09141_;
 wire _09142_;
 wire _09143_;
 wire _09144_;
 wire _09145_;
 wire _09146_;
 wire _09147_;
 wire _09148_;
 wire _09149_;
 wire _09150_;
 wire _09151_;
 wire _09152_;
 wire _09153_;
 wire _09154_;
 wire _09155_;
 wire _09156_;
 wire _09157_;
 wire _09158_;
 wire _09159_;
 wire _09160_;
 wire _09161_;
 wire _09162_;
 wire _09163_;
 wire _09164_;
 wire _09165_;
 wire _09166_;
 wire _09167_;
 wire _09168_;
 wire _09169_;
 wire _09170_;
 wire _09171_;
 wire _09172_;
 wire _09173_;
 wire _09174_;
 wire _09175_;
 wire _09176_;
 wire _09177_;
 wire _09178_;
 wire _09179_;
 wire _09180_;
 wire _09181_;
 wire _09182_;
 wire _09183_;
 wire _09184_;
 wire _09185_;
 wire _09186_;
 wire _09187_;
 wire _09188_;
 wire _09189_;
 wire _09190_;
 wire _09191_;
 wire _09192_;
 wire _09193_;
 wire _09194_;
 wire _09195_;
 wire _09196_;
 wire _09197_;
 wire _09198_;
 wire _09199_;
 wire _09200_;
 wire _09201_;
 wire _09202_;
 wire _09203_;
 wire _09204_;
 wire _09205_;
 wire _09206_;
 wire _09207_;
 wire _09208_;
 wire _09209_;
 wire _09210_;
 wire _09211_;
 wire _09212_;
 wire _09213_;
 wire _09214_;
 wire _09215_;
 wire _09216_;
 wire _09217_;
 wire _09218_;
 wire _09219_;
 wire _09220_;
 wire _09221_;
 wire _09222_;
 wire _09223_;
 wire _09224_;
 wire _09225_;
 wire _09226_;
 wire _09227_;
 wire _09228_;
 wire _09229_;
 wire _09230_;
 wire _09231_;
 wire _09232_;
 wire _09233_;
 wire _09234_;
 wire _09235_;
 wire _09236_;
 wire _09237_;
 wire _09238_;
 wire _09239_;
 wire _09240_;
 wire _09241_;
 wire _09242_;
 wire _09243_;
 wire _09244_;
 wire _09245_;
 wire _09246_;
 wire _09247_;
 wire _09248_;
 wire _09249_;
 wire _09250_;
 wire _09251_;
 wire _09252_;
 wire _09253_;
 wire _09254_;
 wire _09255_;
 wire _09256_;
 wire _09257_;
 wire _09258_;
 wire _09259_;
 wire _09260_;
 wire _09261_;
 wire _09262_;
 wire _09263_;
 wire _09264_;
 wire _09265_;
 wire _09266_;
 wire _09267_;
 wire _09268_;
 wire _09269_;
 wire _09270_;
 wire _09271_;
 wire _09272_;
 wire _09273_;
 wire _09274_;
 wire _09275_;
 wire _09276_;
 wire _09277_;
 wire _09278_;
 wire _09279_;
 wire _09280_;
 wire _09281_;
 wire _09282_;
 wire _09283_;
 wire _09284_;
 wire _09285_;
 wire _09286_;
 wire _09287_;
 wire _09288_;
 wire _09289_;
 wire _09290_;
 wire _09291_;
 wire _09292_;
 wire _09293_;
 wire _09294_;
 wire _09295_;
 wire _09296_;
 wire _09297_;
 wire _09298_;
 wire _09299_;
 wire _09300_;
 wire _09301_;
 wire _09302_;
 wire _09303_;
 wire _09304_;
 wire _09305_;
 wire _09306_;
 wire _09307_;
 wire _09308_;
 wire _09309_;
 wire _09310_;
 wire _09311_;
 wire _09312_;
 wire _09313_;
 wire _09314_;
 wire _09315_;
 wire _09316_;
 wire _09317_;
 wire _09318_;
 wire _09319_;
 wire _09320_;
 wire _09321_;
 wire _09322_;
 wire _09323_;
 wire _09324_;
 wire _09325_;
 wire _09326_;
 wire _09327_;
 wire _09328_;
 wire _09329_;
 wire _09330_;
 wire _09331_;
 wire _09332_;
 wire _09333_;
 wire _09334_;
 wire _09335_;
 wire _09336_;
 wire _09337_;
 wire _09338_;
 wire _09339_;
 wire _09340_;
 wire _09341_;
 wire _09342_;
 wire _09343_;
 wire _09344_;
 wire _09345_;
 wire _09346_;
 wire _09347_;
 wire _09348_;
 wire _09349_;
 wire _09350_;
 wire _09351_;
 wire _09352_;
 wire _09353_;
 wire _09354_;
 wire _09355_;
 wire _09356_;
 wire _09357_;
 wire _09358_;
 wire _09359_;
 wire _09360_;
 wire _09361_;
 wire _09362_;
 wire _09363_;
 wire _09364_;
 wire _09365_;
 wire _09366_;
 wire _09367_;
 wire _09368_;
 wire _09369_;
 wire _09370_;
 wire _09371_;
 wire _09372_;
 wire _09373_;
 wire _09374_;
 wire _09375_;
 wire _09376_;
 wire _09377_;
 wire _09378_;
 wire _09379_;
 wire _09380_;
 wire _09381_;
 wire _09382_;
 wire _09383_;
 wire _09384_;
 wire _09385_;
 wire _09386_;
 wire _09387_;
 wire _09388_;
 wire _09389_;
 wire _09390_;
 wire _09391_;
 wire _09392_;
 wire _09393_;
 wire _09394_;
 wire _09395_;
 wire _09396_;
 wire _09397_;
 wire _09398_;
 wire _09399_;
 wire _09400_;
 wire _09401_;
 wire _09402_;
 wire _09403_;
 wire _09404_;
 wire _09405_;
 wire _09406_;
 wire _09407_;
 wire _09408_;
 wire _09409_;
 wire _09410_;
 wire _09411_;
 wire _09412_;
 wire _09413_;
 wire _09414_;
 wire _09415_;
 wire _09416_;
 wire _09417_;
 wire _09418_;
 wire _09419_;
 wire _09420_;
 wire _09421_;
 wire _09422_;
 wire _09423_;
 wire _09424_;
 wire _09425_;
 wire _09426_;
 wire _09427_;
 wire _09428_;
 wire _09429_;
 wire _09430_;
 wire _09431_;
 wire _09432_;
 wire _09433_;
 wire _09434_;
 wire _09435_;
 wire _09436_;
 wire _09437_;
 wire _09438_;
 wire _09439_;
 wire _09440_;
 wire _09441_;
 wire _09442_;
 wire _09443_;
 wire _09444_;
 wire _09445_;
 wire _09446_;
 wire _09447_;
 wire _09448_;
 wire _09449_;
 wire _09450_;
 wire _09451_;
 wire _09452_;
 wire _09453_;
 wire _09454_;
 wire _09455_;
 wire _09456_;
 wire _09457_;
 wire _09458_;
 wire _09459_;
 wire _09460_;
 wire _09461_;
 wire _09462_;
 wire _09463_;
 wire _09464_;
 wire _09465_;
 wire _09466_;
 wire _09467_;
 wire _09468_;
 wire _09469_;
 wire _09470_;
 wire _09471_;
 wire _09472_;
 wire _09473_;
 wire _09474_;
 wire _09475_;
 wire _09476_;
 wire _09477_;
 wire _09478_;
 wire _09479_;
 wire _09480_;
 wire _09481_;
 wire _09482_;
 wire _09483_;
 wire _09484_;
 wire _09485_;
 wire _09486_;
 wire _09487_;
 wire _09488_;
 wire _09489_;
 wire _09490_;
 wire _09491_;
 wire _09492_;
 wire _09493_;
 wire _09494_;
 wire _09495_;
 wire _09496_;
 wire _09497_;
 wire _09498_;
 wire _09499_;
 wire _09500_;
 wire _09501_;
 wire _09502_;
 wire _09503_;
 wire _09504_;
 wire _09505_;
 wire _09506_;
 wire _09507_;
 wire _09508_;
 wire _09509_;
 wire _09510_;
 wire _09511_;
 wire _09512_;
 wire _09513_;
 wire _09514_;
 wire _09515_;
 wire _09516_;
 wire _09517_;
 wire _09518_;
 wire _09519_;
 wire _09520_;
 wire _09521_;
 wire _09522_;
 wire _09523_;
 wire _09524_;
 wire _09525_;
 wire _09526_;
 wire _09527_;
 wire _09528_;
 wire _09529_;
 wire _09530_;
 wire _09531_;
 wire _09532_;
 wire _09533_;
 wire _09534_;
 wire _09535_;
 wire _09536_;
 wire _09537_;
 wire _09538_;
 wire _09539_;
 wire _09540_;
 wire _09541_;
 wire _09542_;
 wire _09543_;
 wire _09544_;
 wire _09545_;
 wire _09546_;
 wire _09547_;
 wire _09548_;
 wire _09549_;
 wire _09550_;
 wire _09551_;
 wire _09552_;
 wire _09553_;
 wire _09554_;
 wire _09555_;
 wire _09556_;
 wire _09557_;
 wire _09558_;
 wire _09559_;
 wire _09560_;
 wire _09561_;
 wire _09562_;
 wire _09563_;
 wire _09564_;
 wire _09565_;
 wire _09566_;
 wire _09567_;
 wire _09568_;
 wire _09569_;
 wire _09570_;
 wire _09571_;
 wire _09572_;
 wire _09573_;
 wire _09574_;
 wire _09575_;
 wire _09576_;
 wire _09577_;
 wire _09578_;
 wire _09579_;
 wire _09580_;
 wire _09581_;
 wire _09582_;
 wire _09583_;
 wire _09584_;
 wire _09585_;
 wire _09586_;
 wire _09587_;
 wire _09588_;
 wire _09589_;
 wire _09590_;
 wire _09591_;
 wire _09592_;
 wire _09593_;
 wire _09594_;
 wire _09595_;
 wire _09596_;
 wire _09597_;
 wire _09598_;
 wire _09599_;
 wire _09600_;
 wire _09601_;
 wire _09602_;
 wire _09603_;
 wire _09604_;
 wire _09605_;
 wire _09606_;
 wire _09607_;
 wire _09608_;
 wire _09609_;
 wire _09610_;
 wire _09611_;
 wire _09612_;
 wire _09613_;
 wire _09614_;
 wire _09615_;
 wire _09616_;
 wire _09617_;
 wire _09618_;
 wire _09619_;
 wire _09620_;
 wire _09621_;
 wire _09622_;
 wire _09623_;
 wire _09624_;
 wire _09625_;
 wire _09626_;
 wire _09627_;
 wire _09628_;
 wire _09629_;
 wire _09630_;
 wire _09631_;
 wire _09632_;
 wire _09633_;
 wire _09634_;
 wire _09635_;
 wire _09636_;
 wire _09637_;
 wire _09638_;
 wire _09639_;
 wire _09640_;
 wire _09641_;
 wire _09642_;
 wire _09643_;
 wire _09644_;
 wire _09645_;
 wire _09646_;
 wire _09647_;
 wire _09648_;
 wire _09649_;
 wire _09650_;
 wire _09651_;
 wire _09652_;
 wire _09653_;
 wire _09654_;
 wire _09655_;
 wire _09656_;
 wire _09657_;
 wire _09658_;
 wire _09659_;
 wire _09660_;
 wire _09661_;
 wire _09662_;
 wire _09663_;
 wire _09664_;
 wire _09665_;
 wire _09666_;
 wire _09667_;
 wire _09668_;
 wire _09669_;
 wire _09670_;
 wire _09671_;
 wire _09672_;
 wire _09673_;
 wire _09674_;
 wire _09675_;
 wire _09676_;
 wire _09677_;
 wire _09678_;
 wire _09679_;
 wire _09680_;
 wire _09681_;
 wire _09682_;
 wire _09683_;
 wire _09684_;
 wire _09685_;
 wire _09686_;
 wire _09687_;
 wire _09688_;
 wire _09689_;
 wire _09690_;
 wire _09691_;
 wire _09692_;
 wire _09693_;
 wire _09694_;
 wire _09695_;
 wire _09696_;
 wire _09697_;
 wire _09698_;
 wire _09699_;
 wire _09700_;
 wire _09701_;
 wire _09702_;
 wire _09703_;
 wire _09704_;
 wire _09705_;
 wire _09706_;
 wire _09707_;
 wire _09708_;
 wire _09709_;
 wire _09710_;
 wire _09711_;
 wire _09712_;
 wire _09713_;
 wire _09714_;
 wire _09715_;
 wire _09716_;
 wire _09717_;
 wire _09718_;
 wire _09719_;
 wire _09720_;
 wire _09721_;
 wire _09722_;
 wire _09723_;
 wire _09724_;
 wire _09725_;
 wire _09726_;
 wire _09727_;
 wire _09728_;
 wire _09729_;
 wire _09730_;
 wire _09731_;
 wire _09732_;
 wire _09733_;
 wire _09734_;
 wire _09735_;
 wire _09736_;
 wire _09737_;
 wire _09738_;
 wire _09739_;
 wire _09740_;
 wire _09741_;
 wire _09742_;
 wire _09743_;
 wire _09744_;
 wire _09745_;
 wire _09746_;
 wire _09747_;
 wire _09748_;
 wire _09749_;
 wire _09750_;
 wire _09751_;
 wire _09752_;
 wire _09753_;
 wire _09754_;
 wire _09755_;
 wire _09756_;
 wire _09757_;
 wire _09758_;
 wire _09759_;
 wire _09760_;
 wire _09761_;
 wire _09762_;
 wire _09763_;
 wire _09764_;
 wire _09765_;
 wire _09766_;
 wire _09767_;
 wire _09768_;
 wire _09769_;
 wire _09770_;
 wire _09771_;
 wire _09772_;
 wire _09773_;
 wire _09774_;
 wire _09775_;
 wire _09776_;
 wire _09777_;
 wire _09778_;
 wire _09779_;
 wire _09780_;
 wire _09781_;
 wire _09782_;
 wire _09783_;
 wire _09784_;
 wire _09785_;
 wire _09786_;
 wire _09787_;
 wire _09788_;
 wire _09789_;
 wire _09790_;
 wire _09791_;
 wire _09792_;
 wire _09793_;
 wire _09794_;
 wire _09795_;
 wire _09796_;
 wire _09797_;
 wire _09798_;
 wire _09799_;
 wire _09800_;
 wire _09801_;
 wire _09802_;
 wire _09803_;
 wire _09804_;
 wire _09805_;
 wire _09806_;
 wire _09807_;
 wire _09808_;
 wire _09809_;
 wire _09810_;
 wire _09811_;
 wire _09812_;
 wire _09813_;
 wire _09814_;
 wire _09815_;
 wire _09816_;
 wire _09817_;
 wire _09818_;
 wire _09819_;
 wire _09820_;
 wire _09821_;
 wire _09822_;
 wire _09823_;
 wire _09824_;
 wire _09825_;
 wire _09826_;
 wire _09827_;
 wire _09828_;
 wire _09829_;
 wire _09830_;
 wire _09831_;
 wire _09832_;
 wire _09833_;
 wire _09834_;
 wire _09835_;
 wire _09836_;
 wire _09837_;
 wire _09838_;
 wire _09839_;
 wire _09840_;
 wire _09841_;
 wire _09842_;
 wire _09843_;
 wire _09844_;
 wire _09845_;
 wire _09846_;
 wire _09847_;
 wire _09848_;
 wire _09849_;
 wire _09850_;
 wire _09851_;
 wire _09852_;
 wire _09853_;
 wire _09854_;
 wire _09855_;
 wire _09856_;
 wire _09857_;
 wire _09858_;
 wire _09859_;
 wire _09860_;
 wire _09861_;
 wire _09862_;
 wire _09863_;
 wire _09864_;
 wire _09865_;
 wire _09866_;
 wire _09867_;
 wire _09868_;
 wire _09869_;
 wire _09870_;
 wire _09871_;
 wire _09872_;
 wire _09873_;
 wire _09874_;
 wire _09875_;
 wire _09876_;
 wire _09877_;
 wire _09878_;
 wire _09879_;
 wire _09880_;
 wire _09881_;
 wire _09882_;
 wire _09883_;
 wire _09884_;
 wire _09885_;
 wire _09886_;
 wire _09887_;
 wire _09888_;
 wire _09889_;
 wire _09890_;
 wire _09891_;
 wire _09892_;
 wire _09893_;
 wire _09894_;
 wire _09895_;
 wire _09896_;
 wire _09897_;
 wire _09898_;
 wire _09899_;
 wire _09900_;
 wire _09901_;
 wire _09902_;
 wire _09903_;
 wire _09904_;
 wire _09905_;
 wire _09906_;
 wire _09907_;
 wire _09908_;
 wire _09909_;
 wire _09910_;
 wire _09911_;
 wire _09912_;
 wire _09913_;
 wire _09914_;
 wire _09915_;
 wire _09916_;
 wire _09917_;
 wire _09918_;
 wire _09919_;
 wire _09920_;
 wire _09921_;
 wire _09922_;
 wire _09923_;
 wire _09924_;
 wire _09925_;
 wire _09926_;
 wire _09927_;
 wire _09928_;
 wire _09929_;
 wire _09930_;
 wire _09931_;
 wire _09932_;
 wire _09933_;
 wire _09934_;
 wire _09935_;
 wire _09936_;
 wire _09937_;
 wire _09938_;
 wire _09939_;
 wire _09940_;
 wire _09941_;
 wire _09942_;
 wire _09943_;
 wire _09944_;
 wire _09945_;
 wire _09946_;
 wire _09947_;
 wire _09948_;
 wire _09949_;
 wire _09950_;
 wire _09951_;
 wire _09952_;
 wire _09953_;
 wire _09954_;
 wire _09955_;
 wire _09956_;
 wire _09957_;
 wire _09958_;
 wire _09959_;
 wire _09960_;
 wire _09961_;
 wire _09962_;
 wire _09963_;
 wire _09964_;
 wire _09965_;
 wire _09966_;
 wire _09967_;
 wire _09968_;
 wire _09969_;
 wire _09970_;
 wire _09971_;
 wire _09972_;
 wire _09973_;
 wire _09974_;
 wire _09975_;
 wire _09976_;
 wire _09977_;
 wire _09978_;
 wire _09979_;
 wire _09980_;
 wire _09981_;
 wire _09982_;
 wire _09983_;
 wire _09984_;
 wire _09985_;
 wire _09986_;
 wire _09987_;
 wire _09988_;
 wire _09989_;
 wire _09990_;
 wire _09991_;
 wire _09992_;
 wire _09993_;
 wire _09994_;
 wire _09995_;
 wire _09996_;
 wire _09997_;
 wire _09998_;
 wire _09999_;
 wire _10000_;
 wire _10001_;
 wire _10002_;
 wire _10003_;
 wire _10004_;
 wire _10005_;
 wire _10006_;
 wire _10007_;
 wire _10008_;
 wire _10009_;
 wire _10010_;
 wire _10011_;
 wire _10012_;
 wire _10013_;
 wire _10014_;
 wire _10015_;
 wire _10016_;
 wire _10017_;
 wire _10018_;
 wire _10019_;
 wire _10020_;
 wire _10021_;
 wire _10022_;
 wire _10023_;
 wire _10024_;
 wire _10025_;
 wire _10026_;
 wire _10027_;
 wire _10028_;
 wire _10029_;
 wire _10030_;
 wire _10031_;
 wire _10032_;
 wire _10033_;
 wire _10034_;
 wire _10035_;
 wire _10036_;
 wire _10037_;
 wire _10038_;
 wire _10039_;
 wire _10040_;
 wire _10041_;
 wire _10042_;
 wire _10043_;
 wire _10044_;
 wire _10045_;
 wire _10046_;
 wire _10047_;
 wire _10048_;
 wire _10049_;
 wire _10050_;
 wire _10051_;
 wire _10052_;
 wire _10053_;
 wire _10054_;
 wire _10055_;
 wire _10056_;
 wire _10057_;
 wire _10058_;
 wire _10059_;
 wire _10060_;
 wire _10061_;
 wire _10062_;
 wire _10063_;
 wire _10064_;
 wire _10065_;
 wire _10066_;
 wire _10067_;
 wire _10068_;
 wire _10069_;
 wire _10070_;
 wire _10071_;
 wire _10072_;
 wire _10073_;
 wire _10074_;
 wire _10075_;
 wire _10076_;
 wire _10077_;
 wire _10078_;
 wire _10079_;
 wire _10080_;
 wire _10081_;
 wire _10082_;
 wire _10083_;
 wire _10084_;
 wire _10085_;
 wire _10086_;
 wire _10087_;
 wire _10088_;
 wire _10089_;
 wire _10090_;
 wire _10091_;
 wire _10092_;
 wire _10093_;
 wire _10094_;
 wire _10095_;
 wire _10096_;
 wire _10097_;
 wire _10098_;
 wire _10099_;
 wire _10100_;
 wire _10101_;
 wire _10102_;
 wire _10103_;
 wire _10104_;
 wire _10105_;
 wire _10106_;
 wire _10107_;
 wire _10108_;
 wire _10109_;
 wire _10110_;
 wire _10111_;
 wire _10112_;
 wire _10113_;
 wire _10114_;
 wire _10115_;
 wire _10116_;
 wire _10117_;
 wire _10118_;
 wire _10119_;
 wire _10120_;
 wire _10121_;
 wire _10122_;
 wire _10123_;
 wire _10124_;
 wire _10125_;
 wire _10126_;
 wire _10127_;
 wire _10128_;
 wire _10129_;
 wire _10130_;
 wire _10131_;
 wire _10132_;
 wire _10133_;
 wire _10134_;
 wire _10135_;
 wire _10136_;
 wire _10137_;
 wire _10138_;
 wire _10139_;
 wire _10140_;
 wire _10141_;
 wire _10142_;
 wire _10143_;
 wire _10144_;
 wire _10145_;
 wire _10146_;
 wire _10147_;
 wire _10148_;
 wire _10149_;
 wire _10150_;
 wire _10151_;
 wire _10152_;
 wire _10153_;
 wire _10154_;
 wire _10155_;
 wire _10156_;
 wire _10157_;
 wire _10158_;
 wire _10159_;
 wire _10160_;
 wire _10161_;
 wire _10162_;
 wire _10163_;
 wire _10164_;
 wire _10165_;
 wire _10166_;
 wire _10167_;
 wire _10168_;
 wire _10169_;
 wire _10170_;
 wire _10171_;
 wire _10172_;
 wire _10173_;
 wire _10174_;
 wire _10175_;
 wire _10176_;
 wire _10177_;
 wire _10178_;
 wire _10179_;
 wire _10180_;
 wire _10181_;
 wire _10182_;
 wire _10183_;
 wire _10184_;
 wire _10185_;
 wire _10186_;
 wire _10187_;
 wire _10188_;
 wire _10189_;
 wire _10190_;
 wire _10191_;
 wire _10192_;
 wire _10193_;
 wire _10194_;
 wire _10195_;
 wire _10196_;
 wire _10197_;
 wire _10198_;
 wire _10199_;
 wire _10200_;
 wire _10201_;
 wire _10202_;
 wire _10203_;
 wire _10204_;
 wire _10205_;
 wire _10206_;
 wire _10207_;
 wire _10208_;
 wire _10209_;
 wire _10210_;
 wire _10211_;
 wire _10212_;
 wire _10213_;
 wire _10214_;
 wire _10215_;
 wire _10216_;
 wire _10217_;
 wire _10218_;
 wire _10219_;
 wire _10220_;
 wire _10221_;
 wire _10222_;
 wire _10223_;
 wire _10224_;
 wire _10225_;
 wire _10226_;
 wire _10227_;
 wire _10228_;
 wire _10229_;
 wire _10230_;
 wire _10231_;
 wire _10232_;
 wire _10233_;
 wire _10234_;
 wire _10235_;
 wire _10236_;
 wire _10237_;
 wire _10238_;
 wire _10239_;
 wire _10240_;
 wire _10241_;
 wire _10242_;
 wire _10243_;
 wire _10244_;
 wire _10245_;
 wire _10246_;
 wire _10247_;
 wire _10248_;
 wire _10249_;
 wire _10250_;
 wire _10251_;
 wire _10252_;
 wire _10253_;
 wire _10254_;
 wire _10255_;
 wire _10256_;
 wire _10257_;
 wire _10258_;
 wire _10259_;
 wire _10260_;
 wire _10261_;
 wire _10262_;
 wire _10263_;
 wire _10264_;
 wire _10265_;
 wire _10266_;
 wire _10267_;
 wire _10268_;
 wire _10269_;
 wire _10270_;
 wire _10271_;
 wire _10272_;
 wire _10273_;
 wire _10274_;
 wire _10275_;
 wire _10276_;
 wire _10277_;
 wire _10278_;
 wire _10279_;
 wire _10280_;
 wire _10281_;
 wire _10282_;
 wire _10283_;
 wire _10284_;
 wire _10285_;
 wire _10286_;
 wire _10287_;
 wire _10288_;
 wire _10289_;
 wire _10290_;
 wire _10291_;
 wire _10292_;
 wire _10293_;
 wire _10294_;
 wire _10295_;
 wire _10296_;
 wire _10297_;
 wire _10298_;
 wire _10299_;
 wire _10300_;
 wire _10301_;
 wire _10302_;
 wire _10303_;
 wire _10304_;
 wire _10305_;
 wire _10306_;
 wire _10307_;
 wire _10308_;
 wire _10309_;
 wire _10310_;
 wire _10311_;
 wire _10312_;
 wire _10313_;
 wire _10314_;
 wire _10315_;
 wire _10316_;
 wire _10317_;
 wire _10318_;
 wire _10319_;
 wire _10320_;
 wire _10321_;
 wire _10322_;
 wire _10323_;
 wire _10324_;
 wire _10325_;
 wire _10326_;
 wire _10327_;
 wire _10328_;
 wire _10329_;
 wire _10330_;
 wire _10331_;
 wire _10332_;
 wire _10333_;
 wire _10334_;
 wire _10335_;
 wire _10336_;
 wire _10337_;
 wire _10338_;
 wire _10339_;
 wire _10340_;
 wire _10341_;
 wire _10342_;
 wire _10343_;
 wire _10344_;
 wire _10345_;
 wire _10346_;
 wire _10347_;
 wire _10348_;
 wire _10349_;
 wire _10350_;
 wire _10351_;
 wire _10352_;
 wire _10353_;
 wire _10354_;
 wire _10355_;
 wire _10356_;
 wire _10357_;
 wire _10358_;
 wire _10359_;
 wire _10360_;
 wire _10361_;
 wire _10362_;
 wire _10363_;
 wire _10364_;
 wire _10365_;
 wire _10366_;
 wire net27;
 wire net28;
 wire _10369_;
 wire _10370_;
 wire output_ready;
 wire spi_instruction_done;
 wire \spiking_network_top_uut.SNN_en_sync ;
 wire \spiking_network_top_uut.SPI_reset_synchr ;
 wire \spiking_network_top_uut.all_data_out[0] ;
 wire \spiking_network_top_uut.all_data_out[100] ;
 wire \spiking_network_top_uut.all_data_out[101] ;
 wire \spiking_network_top_uut.all_data_out[102] ;
 wire \spiking_network_top_uut.all_data_out[103] ;
 wire \spiking_network_top_uut.all_data_out[104] ;
 wire \spiking_network_top_uut.all_data_out[105] ;
 wire \spiking_network_top_uut.all_data_out[106] ;
 wire \spiking_network_top_uut.all_data_out[107] ;
 wire \spiking_network_top_uut.all_data_out[108] ;
 wire \spiking_network_top_uut.all_data_out[109] ;
 wire \spiking_network_top_uut.all_data_out[10] ;
 wire \spiking_network_top_uut.all_data_out[110] ;
 wire \spiking_network_top_uut.all_data_out[111] ;
 wire \spiking_network_top_uut.all_data_out[112] ;
 wire \spiking_network_top_uut.all_data_out[113] ;
 wire \spiking_network_top_uut.all_data_out[114] ;
 wire \spiking_network_top_uut.all_data_out[115] ;
 wire \spiking_network_top_uut.all_data_out[116] ;
 wire \spiking_network_top_uut.all_data_out[117] ;
 wire \spiking_network_top_uut.all_data_out[118] ;
 wire \spiking_network_top_uut.all_data_out[119] ;
 wire \spiking_network_top_uut.all_data_out[11] ;
 wire \spiking_network_top_uut.all_data_out[120] ;
 wire \spiking_network_top_uut.all_data_out[121] ;
 wire \spiking_network_top_uut.all_data_out[122] ;
 wire \spiking_network_top_uut.all_data_out[123] ;
 wire \spiking_network_top_uut.all_data_out[124] ;
 wire \spiking_network_top_uut.all_data_out[125] ;
 wire \spiking_network_top_uut.all_data_out[126] ;
 wire \spiking_network_top_uut.all_data_out[127] ;
 wire \spiking_network_top_uut.all_data_out[128] ;
 wire \spiking_network_top_uut.all_data_out[129] ;
 wire \spiking_network_top_uut.all_data_out[12] ;
 wire \spiking_network_top_uut.all_data_out[130] ;
 wire \spiking_network_top_uut.all_data_out[131] ;
 wire \spiking_network_top_uut.all_data_out[132] ;
 wire \spiking_network_top_uut.all_data_out[133] ;
 wire \spiking_network_top_uut.all_data_out[134] ;
 wire \spiking_network_top_uut.all_data_out[135] ;
 wire \spiking_network_top_uut.all_data_out[136] ;
 wire \spiking_network_top_uut.all_data_out[137] ;
 wire \spiking_network_top_uut.all_data_out[138] ;
 wire \spiking_network_top_uut.all_data_out[139] ;
 wire \spiking_network_top_uut.all_data_out[13] ;
 wire \spiking_network_top_uut.all_data_out[140] ;
 wire \spiking_network_top_uut.all_data_out[141] ;
 wire \spiking_network_top_uut.all_data_out[142] ;
 wire \spiking_network_top_uut.all_data_out[143] ;
 wire \spiking_network_top_uut.all_data_out[144] ;
 wire \spiking_network_top_uut.all_data_out[145] ;
 wire \spiking_network_top_uut.all_data_out[146] ;
 wire \spiking_network_top_uut.all_data_out[147] ;
 wire \spiking_network_top_uut.all_data_out[148] ;
 wire \spiking_network_top_uut.all_data_out[149] ;
 wire \spiking_network_top_uut.all_data_out[14] ;
 wire \spiking_network_top_uut.all_data_out[150] ;
 wire \spiking_network_top_uut.all_data_out[151] ;
 wire \spiking_network_top_uut.all_data_out[152] ;
 wire \spiking_network_top_uut.all_data_out[153] ;
 wire \spiking_network_top_uut.all_data_out[154] ;
 wire \spiking_network_top_uut.all_data_out[155] ;
 wire \spiking_network_top_uut.all_data_out[156] ;
 wire \spiking_network_top_uut.all_data_out[157] ;
 wire \spiking_network_top_uut.all_data_out[158] ;
 wire \spiking_network_top_uut.all_data_out[159] ;
 wire \spiking_network_top_uut.all_data_out[15] ;
 wire \spiking_network_top_uut.all_data_out[160] ;
 wire \spiking_network_top_uut.all_data_out[161] ;
 wire \spiking_network_top_uut.all_data_out[162] ;
 wire \spiking_network_top_uut.all_data_out[163] ;
 wire \spiking_network_top_uut.all_data_out[164] ;
 wire \spiking_network_top_uut.all_data_out[165] ;
 wire \spiking_network_top_uut.all_data_out[166] ;
 wire \spiking_network_top_uut.all_data_out[167] ;
 wire \spiking_network_top_uut.all_data_out[168] ;
 wire \spiking_network_top_uut.all_data_out[169] ;
 wire \spiking_network_top_uut.all_data_out[16] ;
 wire \spiking_network_top_uut.all_data_out[170] ;
 wire \spiking_network_top_uut.all_data_out[171] ;
 wire \spiking_network_top_uut.all_data_out[172] ;
 wire \spiking_network_top_uut.all_data_out[173] ;
 wire \spiking_network_top_uut.all_data_out[174] ;
 wire \spiking_network_top_uut.all_data_out[175] ;
 wire \spiking_network_top_uut.all_data_out[176] ;
 wire \spiking_network_top_uut.all_data_out[177] ;
 wire \spiking_network_top_uut.all_data_out[178] ;
 wire \spiking_network_top_uut.all_data_out[179] ;
 wire \spiking_network_top_uut.all_data_out[17] ;
 wire \spiking_network_top_uut.all_data_out[180] ;
 wire \spiking_network_top_uut.all_data_out[181] ;
 wire \spiking_network_top_uut.all_data_out[182] ;
 wire \spiking_network_top_uut.all_data_out[183] ;
 wire \spiking_network_top_uut.all_data_out[184] ;
 wire \spiking_network_top_uut.all_data_out[185] ;
 wire \spiking_network_top_uut.all_data_out[186] ;
 wire \spiking_network_top_uut.all_data_out[187] ;
 wire \spiking_network_top_uut.all_data_out[188] ;
 wire \spiking_network_top_uut.all_data_out[189] ;
 wire \spiking_network_top_uut.all_data_out[18] ;
 wire \spiking_network_top_uut.all_data_out[190] ;
 wire \spiking_network_top_uut.all_data_out[191] ;
 wire \spiking_network_top_uut.all_data_out[192] ;
 wire \spiking_network_top_uut.all_data_out[193] ;
 wire \spiking_network_top_uut.all_data_out[194] ;
 wire \spiking_network_top_uut.all_data_out[195] ;
 wire \spiking_network_top_uut.all_data_out[196] ;
 wire \spiking_network_top_uut.all_data_out[197] ;
 wire \spiking_network_top_uut.all_data_out[198] ;
 wire \spiking_network_top_uut.all_data_out[199] ;
 wire \spiking_network_top_uut.all_data_out[19] ;
 wire \spiking_network_top_uut.all_data_out[1] ;
 wire \spiking_network_top_uut.all_data_out[200] ;
 wire \spiking_network_top_uut.all_data_out[201] ;
 wire \spiking_network_top_uut.all_data_out[202] ;
 wire \spiking_network_top_uut.all_data_out[203] ;
 wire \spiking_network_top_uut.all_data_out[204] ;
 wire \spiking_network_top_uut.all_data_out[205] ;
 wire \spiking_network_top_uut.all_data_out[206] ;
 wire \spiking_network_top_uut.all_data_out[207] ;
 wire \spiking_network_top_uut.all_data_out[208] ;
 wire \spiking_network_top_uut.all_data_out[209] ;
 wire \spiking_network_top_uut.all_data_out[20] ;
 wire \spiking_network_top_uut.all_data_out[210] ;
 wire \spiking_network_top_uut.all_data_out[211] ;
 wire \spiking_network_top_uut.all_data_out[212] ;
 wire \spiking_network_top_uut.all_data_out[213] ;
 wire \spiking_network_top_uut.all_data_out[214] ;
 wire \spiking_network_top_uut.all_data_out[215] ;
 wire \spiking_network_top_uut.all_data_out[216] ;
 wire \spiking_network_top_uut.all_data_out[217] ;
 wire \spiking_network_top_uut.all_data_out[218] ;
 wire \spiking_network_top_uut.all_data_out[219] ;
 wire \spiking_network_top_uut.all_data_out[21] ;
 wire \spiking_network_top_uut.all_data_out[220] ;
 wire \spiking_network_top_uut.all_data_out[221] ;
 wire \spiking_network_top_uut.all_data_out[222] ;
 wire \spiking_network_top_uut.all_data_out[223] ;
 wire \spiking_network_top_uut.all_data_out[224] ;
 wire \spiking_network_top_uut.all_data_out[225] ;
 wire \spiking_network_top_uut.all_data_out[226] ;
 wire \spiking_network_top_uut.all_data_out[227] ;
 wire \spiking_network_top_uut.all_data_out[228] ;
 wire \spiking_network_top_uut.all_data_out[229] ;
 wire \spiking_network_top_uut.all_data_out[22] ;
 wire \spiking_network_top_uut.all_data_out[230] ;
 wire \spiking_network_top_uut.all_data_out[231] ;
 wire \spiking_network_top_uut.all_data_out[232] ;
 wire \spiking_network_top_uut.all_data_out[233] ;
 wire \spiking_network_top_uut.all_data_out[234] ;
 wire \spiking_network_top_uut.all_data_out[235] ;
 wire \spiking_network_top_uut.all_data_out[236] ;
 wire \spiking_network_top_uut.all_data_out[237] ;
 wire \spiking_network_top_uut.all_data_out[238] ;
 wire \spiking_network_top_uut.all_data_out[239] ;
 wire \spiking_network_top_uut.all_data_out[23] ;
 wire \spiking_network_top_uut.all_data_out[240] ;
 wire \spiking_network_top_uut.all_data_out[241] ;
 wire \spiking_network_top_uut.all_data_out[242] ;
 wire \spiking_network_top_uut.all_data_out[243] ;
 wire \spiking_network_top_uut.all_data_out[244] ;
 wire \spiking_network_top_uut.all_data_out[245] ;
 wire \spiking_network_top_uut.all_data_out[246] ;
 wire \spiking_network_top_uut.all_data_out[247] ;
 wire \spiking_network_top_uut.all_data_out[248] ;
 wire \spiking_network_top_uut.all_data_out[249] ;
 wire \spiking_network_top_uut.all_data_out[24] ;
 wire \spiking_network_top_uut.all_data_out[250] ;
 wire \spiking_network_top_uut.all_data_out[251] ;
 wire \spiking_network_top_uut.all_data_out[252] ;
 wire \spiking_network_top_uut.all_data_out[253] ;
 wire \spiking_network_top_uut.all_data_out[254] ;
 wire \spiking_network_top_uut.all_data_out[255] ;
 wire \spiking_network_top_uut.all_data_out[256] ;
 wire \spiking_network_top_uut.all_data_out[257] ;
 wire \spiking_network_top_uut.all_data_out[258] ;
 wire \spiking_network_top_uut.all_data_out[259] ;
 wire \spiking_network_top_uut.all_data_out[25] ;
 wire \spiking_network_top_uut.all_data_out[260] ;
 wire \spiking_network_top_uut.all_data_out[261] ;
 wire \spiking_network_top_uut.all_data_out[262] ;
 wire \spiking_network_top_uut.all_data_out[263] ;
 wire \spiking_network_top_uut.all_data_out[264] ;
 wire \spiking_network_top_uut.all_data_out[265] ;
 wire \spiking_network_top_uut.all_data_out[266] ;
 wire \spiking_network_top_uut.all_data_out[267] ;
 wire \spiking_network_top_uut.all_data_out[268] ;
 wire \spiking_network_top_uut.all_data_out[269] ;
 wire \spiking_network_top_uut.all_data_out[26] ;
 wire \spiking_network_top_uut.all_data_out[270] ;
 wire \spiking_network_top_uut.all_data_out[271] ;
 wire \spiking_network_top_uut.all_data_out[272] ;
 wire \spiking_network_top_uut.all_data_out[273] ;
 wire \spiking_network_top_uut.all_data_out[274] ;
 wire \spiking_network_top_uut.all_data_out[275] ;
 wire \spiking_network_top_uut.all_data_out[276] ;
 wire \spiking_network_top_uut.all_data_out[277] ;
 wire \spiking_network_top_uut.all_data_out[278] ;
 wire \spiking_network_top_uut.all_data_out[279] ;
 wire \spiking_network_top_uut.all_data_out[27] ;
 wire \spiking_network_top_uut.all_data_out[280] ;
 wire \spiking_network_top_uut.all_data_out[281] ;
 wire \spiking_network_top_uut.all_data_out[282] ;
 wire \spiking_network_top_uut.all_data_out[283] ;
 wire \spiking_network_top_uut.all_data_out[284] ;
 wire \spiking_network_top_uut.all_data_out[285] ;
 wire \spiking_network_top_uut.all_data_out[286] ;
 wire \spiking_network_top_uut.all_data_out[287] ;
 wire \spiking_network_top_uut.all_data_out[288] ;
 wire \spiking_network_top_uut.all_data_out[289] ;
 wire \spiking_network_top_uut.all_data_out[28] ;
 wire \spiking_network_top_uut.all_data_out[290] ;
 wire \spiking_network_top_uut.all_data_out[291] ;
 wire \spiking_network_top_uut.all_data_out[292] ;
 wire \spiking_network_top_uut.all_data_out[293] ;
 wire \spiking_network_top_uut.all_data_out[294] ;
 wire \spiking_network_top_uut.all_data_out[295] ;
 wire \spiking_network_top_uut.all_data_out[296] ;
 wire \spiking_network_top_uut.all_data_out[297] ;
 wire \spiking_network_top_uut.all_data_out[298] ;
 wire \spiking_network_top_uut.all_data_out[299] ;
 wire \spiking_network_top_uut.all_data_out[29] ;
 wire \spiking_network_top_uut.all_data_out[2] ;
 wire \spiking_network_top_uut.all_data_out[300] ;
 wire \spiking_network_top_uut.all_data_out[301] ;
 wire \spiking_network_top_uut.all_data_out[302] ;
 wire \spiking_network_top_uut.all_data_out[303] ;
 wire \spiking_network_top_uut.all_data_out[304] ;
 wire \spiking_network_top_uut.all_data_out[305] ;
 wire \spiking_network_top_uut.all_data_out[306] ;
 wire \spiking_network_top_uut.all_data_out[307] ;
 wire \spiking_network_top_uut.all_data_out[308] ;
 wire \spiking_network_top_uut.all_data_out[309] ;
 wire \spiking_network_top_uut.all_data_out[30] ;
 wire \spiking_network_top_uut.all_data_out[310] ;
 wire \spiking_network_top_uut.all_data_out[311] ;
 wire \spiking_network_top_uut.all_data_out[312] ;
 wire \spiking_network_top_uut.all_data_out[313] ;
 wire \spiking_network_top_uut.all_data_out[314] ;
 wire \spiking_network_top_uut.all_data_out[315] ;
 wire \spiking_network_top_uut.all_data_out[316] ;
 wire \spiking_network_top_uut.all_data_out[317] ;
 wire \spiking_network_top_uut.all_data_out[318] ;
 wire \spiking_network_top_uut.all_data_out[319] ;
 wire \spiking_network_top_uut.all_data_out[31] ;
 wire \spiking_network_top_uut.all_data_out[320] ;
 wire \spiking_network_top_uut.all_data_out[321] ;
 wire \spiking_network_top_uut.all_data_out[322] ;
 wire \spiking_network_top_uut.all_data_out[323] ;
 wire \spiking_network_top_uut.all_data_out[324] ;
 wire \spiking_network_top_uut.all_data_out[325] ;
 wire \spiking_network_top_uut.all_data_out[326] ;
 wire \spiking_network_top_uut.all_data_out[327] ;
 wire \spiking_network_top_uut.all_data_out[328] ;
 wire \spiking_network_top_uut.all_data_out[329] ;
 wire \spiking_network_top_uut.all_data_out[32] ;
 wire \spiking_network_top_uut.all_data_out[330] ;
 wire \spiking_network_top_uut.all_data_out[331] ;
 wire \spiking_network_top_uut.all_data_out[332] ;
 wire \spiking_network_top_uut.all_data_out[333] ;
 wire \spiking_network_top_uut.all_data_out[334] ;
 wire \spiking_network_top_uut.all_data_out[335] ;
 wire \spiking_network_top_uut.all_data_out[336] ;
 wire \spiking_network_top_uut.all_data_out[337] ;
 wire \spiking_network_top_uut.all_data_out[338] ;
 wire \spiking_network_top_uut.all_data_out[339] ;
 wire \spiking_network_top_uut.all_data_out[33] ;
 wire \spiking_network_top_uut.all_data_out[340] ;
 wire \spiking_network_top_uut.all_data_out[341] ;
 wire \spiking_network_top_uut.all_data_out[342] ;
 wire \spiking_network_top_uut.all_data_out[343] ;
 wire \spiking_network_top_uut.all_data_out[344] ;
 wire \spiking_network_top_uut.all_data_out[345] ;
 wire \spiking_network_top_uut.all_data_out[346] ;
 wire \spiking_network_top_uut.all_data_out[347] ;
 wire \spiking_network_top_uut.all_data_out[348] ;
 wire \spiking_network_top_uut.all_data_out[349] ;
 wire \spiking_network_top_uut.all_data_out[34] ;
 wire \spiking_network_top_uut.all_data_out[350] ;
 wire \spiking_network_top_uut.all_data_out[351] ;
 wire \spiking_network_top_uut.all_data_out[352] ;
 wire \spiking_network_top_uut.all_data_out[353] ;
 wire \spiking_network_top_uut.all_data_out[354] ;
 wire \spiking_network_top_uut.all_data_out[355] ;
 wire \spiking_network_top_uut.all_data_out[356] ;
 wire \spiking_network_top_uut.all_data_out[357] ;
 wire \spiking_network_top_uut.all_data_out[358] ;
 wire \spiking_network_top_uut.all_data_out[359] ;
 wire \spiking_network_top_uut.all_data_out[35] ;
 wire \spiking_network_top_uut.all_data_out[360] ;
 wire \spiking_network_top_uut.all_data_out[361] ;
 wire \spiking_network_top_uut.all_data_out[362] ;
 wire \spiking_network_top_uut.all_data_out[363] ;
 wire \spiking_network_top_uut.all_data_out[364] ;
 wire \spiking_network_top_uut.all_data_out[365] ;
 wire \spiking_network_top_uut.all_data_out[366] ;
 wire \spiking_network_top_uut.all_data_out[367] ;
 wire \spiking_network_top_uut.all_data_out[368] ;
 wire \spiking_network_top_uut.all_data_out[369] ;
 wire \spiking_network_top_uut.all_data_out[36] ;
 wire \spiking_network_top_uut.all_data_out[370] ;
 wire \spiking_network_top_uut.all_data_out[371] ;
 wire \spiking_network_top_uut.all_data_out[372] ;
 wire \spiking_network_top_uut.all_data_out[373] ;
 wire \spiking_network_top_uut.all_data_out[374] ;
 wire \spiking_network_top_uut.all_data_out[375] ;
 wire \spiking_network_top_uut.all_data_out[376] ;
 wire \spiking_network_top_uut.all_data_out[377] ;
 wire \spiking_network_top_uut.all_data_out[378] ;
 wire \spiking_network_top_uut.all_data_out[379] ;
 wire \spiking_network_top_uut.all_data_out[37] ;
 wire \spiking_network_top_uut.all_data_out[380] ;
 wire \spiking_network_top_uut.all_data_out[381] ;
 wire \spiking_network_top_uut.all_data_out[382] ;
 wire \spiking_network_top_uut.all_data_out[383] ;
 wire \spiking_network_top_uut.all_data_out[384] ;
 wire \spiking_network_top_uut.all_data_out[385] ;
 wire \spiking_network_top_uut.all_data_out[386] ;
 wire \spiking_network_top_uut.all_data_out[387] ;
 wire \spiking_network_top_uut.all_data_out[388] ;
 wire \spiking_network_top_uut.all_data_out[389] ;
 wire \spiking_network_top_uut.all_data_out[38] ;
 wire \spiking_network_top_uut.all_data_out[390] ;
 wire \spiking_network_top_uut.all_data_out[391] ;
 wire \spiking_network_top_uut.all_data_out[392] ;
 wire \spiking_network_top_uut.all_data_out[393] ;
 wire \spiking_network_top_uut.all_data_out[394] ;
 wire \spiking_network_top_uut.all_data_out[395] ;
 wire \spiking_network_top_uut.all_data_out[396] ;
 wire \spiking_network_top_uut.all_data_out[397] ;
 wire \spiking_network_top_uut.all_data_out[398] ;
 wire \spiking_network_top_uut.all_data_out[399] ;
 wire \spiking_network_top_uut.all_data_out[39] ;
 wire \spiking_network_top_uut.all_data_out[3] ;
 wire \spiking_network_top_uut.all_data_out[400] ;
 wire \spiking_network_top_uut.all_data_out[401] ;
 wire \spiking_network_top_uut.all_data_out[402] ;
 wire \spiking_network_top_uut.all_data_out[403] ;
 wire \spiking_network_top_uut.all_data_out[404] ;
 wire \spiking_network_top_uut.all_data_out[405] ;
 wire \spiking_network_top_uut.all_data_out[406] ;
 wire \spiking_network_top_uut.all_data_out[407] ;
 wire \spiking_network_top_uut.all_data_out[408] ;
 wire \spiking_network_top_uut.all_data_out[409] ;
 wire \spiking_network_top_uut.all_data_out[40] ;
 wire \spiking_network_top_uut.all_data_out[410] ;
 wire \spiking_network_top_uut.all_data_out[411] ;
 wire \spiking_network_top_uut.all_data_out[412] ;
 wire \spiking_network_top_uut.all_data_out[413] ;
 wire \spiking_network_top_uut.all_data_out[414] ;
 wire \spiking_network_top_uut.all_data_out[415] ;
 wire \spiking_network_top_uut.all_data_out[416] ;
 wire \spiking_network_top_uut.all_data_out[417] ;
 wire \spiking_network_top_uut.all_data_out[418] ;
 wire \spiking_network_top_uut.all_data_out[419] ;
 wire \spiking_network_top_uut.all_data_out[41] ;
 wire \spiking_network_top_uut.all_data_out[420] ;
 wire \spiking_network_top_uut.all_data_out[421] ;
 wire \spiking_network_top_uut.all_data_out[422] ;
 wire \spiking_network_top_uut.all_data_out[423] ;
 wire \spiking_network_top_uut.all_data_out[424] ;
 wire \spiking_network_top_uut.all_data_out[425] ;
 wire \spiking_network_top_uut.all_data_out[426] ;
 wire \spiking_network_top_uut.all_data_out[427] ;
 wire \spiking_network_top_uut.all_data_out[428] ;
 wire \spiking_network_top_uut.all_data_out[429] ;
 wire \spiking_network_top_uut.all_data_out[42] ;
 wire \spiking_network_top_uut.all_data_out[430] ;
 wire \spiking_network_top_uut.all_data_out[431] ;
 wire \spiking_network_top_uut.all_data_out[432] ;
 wire \spiking_network_top_uut.all_data_out[433] ;
 wire \spiking_network_top_uut.all_data_out[434] ;
 wire \spiking_network_top_uut.all_data_out[435] ;
 wire \spiking_network_top_uut.all_data_out[436] ;
 wire \spiking_network_top_uut.all_data_out[437] ;
 wire \spiking_network_top_uut.all_data_out[438] ;
 wire \spiking_network_top_uut.all_data_out[439] ;
 wire \spiking_network_top_uut.all_data_out[43] ;
 wire \spiking_network_top_uut.all_data_out[440] ;
 wire \spiking_network_top_uut.all_data_out[441] ;
 wire \spiking_network_top_uut.all_data_out[442] ;
 wire \spiking_network_top_uut.all_data_out[443] ;
 wire \spiking_network_top_uut.all_data_out[444] ;
 wire \spiking_network_top_uut.all_data_out[445] ;
 wire \spiking_network_top_uut.all_data_out[446] ;
 wire \spiking_network_top_uut.all_data_out[447] ;
 wire \spiking_network_top_uut.all_data_out[448] ;
 wire \spiking_network_top_uut.all_data_out[449] ;
 wire \spiking_network_top_uut.all_data_out[44] ;
 wire \spiking_network_top_uut.all_data_out[450] ;
 wire \spiking_network_top_uut.all_data_out[451] ;
 wire \spiking_network_top_uut.all_data_out[452] ;
 wire \spiking_network_top_uut.all_data_out[453] ;
 wire \spiking_network_top_uut.all_data_out[454] ;
 wire \spiking_network_top_uut.all_data_out[455] ;
 wire \spiking_network_top_uut.all_data_out[456] ;
 wire \spiking_network_top_uut.all_data_out[457] ;
 wire \spiking_network_top_uut.all_data_out[458] ;
 wire \spiking_network_top_uut.all_data_out[459] ;
 wire \spiking_network_top_uut.all_data_out[45] ;
 wire \spiking_network_top_uut.all_data_out[460] ;
 wire \spiking_network_top_uut.all_data_out[461] ;
 wire \spiking_network_top_uut.all_data_out[462] ;
 wire \spiking_network_top_uut.all_data_out[463] ;
 wire \spiking_network_top_uut.all_data_out[464] ;
 wire \spiking_network_top_uut.all_data_out[465] ;
 wire \spiking_network_top_uut.all_data_out[466] ;
 wire \spiking_network_top_uut.all_data_out[467] ;
 wire \spiking_network_top_uut.all_data_out[468] ;
 wire \spiking_network_top_uut.all_data_out[469] ;
 wire \spiking_network_top_uut.all_data_out[46] ;
 wire \spiking_network_top_uut.all_data_out[470] ;
 wire \spiking_network_top_uut.all_data_out[471] ;
 wire \spiking_network_top_uut.all_data_out[472] ;
 wire \spiking_network_top_uut.all_data_out[473] ;
 wire \spiking_network_top_uut.all_data_out[474] ;
 wire \spiking_network_top_uut.all_data_out[475] ;
 wire \spiking_network_top_uut.all_data_out[476] ;
 wire \spiking_network_top_uut.all_data_out[477] ;
 wire \spiking_network_top_uut.all_data_out[478] ;
 wire \spiking_network_top_uut.all_data_out[479] ;
 wire \spiking_network_top_uut.all_data_out[47] ;
 wire \spiking_network_top_uut.all_data_out[480] ;
 wire \spiking_network_top_uut.all_data_out[481] ;
 wire \spiking_network_top_uut.all_data_out[482] ;
 wire \spiking_network_top_uut.all_data_out[483] ;
 wire \spiking_network_top_uut.all_data_out[484] ;
 wire \spiking_network_top_uut.all_data_out[485] ;
 wire \spiking_network_top_uut.all_data_out[486] ;
 wire \spiking_network_top_uut.all_data_out[487] ;
 wire \spiking_network_top_uut.all_data_out[488] ;
 wire \spiking_network_top_uut.all_data_out[489] ;
 wire \spiking_network_top_uut.all_data_out[48] ;
 wire \spiking_network_top_uut.all_data_out[490] ;
 wire \spiking_network_top_uut.all_data_out[491] ;
 wire \spiking_network_top_uut.all_data_out[492] ;
 wire \spiking_network_top_uut.all_data_out[493] ;
 wire \spiking_network_top_uut.all_data_out[494] ;
 wire \spiking_network_top_uut.all_data_out[495] ;
 wire \spiking_network_top_uut.all_data_out[496] ;
 wire \spiking_network_top_uut.all_data_out[497] ;
 wire \spiking_network_top_uut.all_data_out[498] ;
 wire \spiking_network_top_uut.all_data_out[499] ;
 wire \spiking_network_top_uut.all_data_out[49] ;
 wire \spiking_network_top_uut.all_data_out[4] ;
 wire \spiking_network_top_uut.all_data_out[500] ;
 wire \spiking_network_top_uut.all_data_out[501] ;
 wire \spiking_network_top_uut.all_data_out[502] ;
 wire \spiking_network_top_uut.all_data_out[503] ;
 wire \spiking_network_top_uut.all_data_out[504] ;
 wire \spiking_network_top_uut.all_data_out[505] ;
 wire \spiking_network_top_uut.all_data_out[506] ;
 wire \spiking_network_top_uut.all_data_out[507] ;
 wire \spiking_network_top_uut.all_data_out[508] ;
 wire \spiking_network_top_uut.all_data_out[509] ;
 wire \spiking_network_top_uut.all_data_out[50] ;
 wire \spiking_network_top_uut.all_data_out[510] ;
 wire \spiking_network_top_uut.all_data_out[511] ;
 wire \spiking_network_top_uut.all_data_out[512] ;
 wire \spiking_network_top_uut.all_data_out[513] ;
 wire \spiking_network_top_uut.all_data_out[514] ;
 wire \spiking_network_top_uut.all_data_out[515] ;
 wire \spiking_network_top_uut.all_data_out[516] ;
 wire \spiking_network_top_uut.all_data_out[517] ;
 wire \spiking_network_top_uut.all_data_out[518] ;
 wire \spiking_network_top_uut.all_data_out[519] ;
 wire \spiking_network_top_uut.all_data_out[51] ;
 wire \spiking_network_top_uut.all_data_out[520] ;
 wire \spiking_network_top_uut.all_data_out[521] ;
 wire \spiking_network_top_uut.all_data_out[522] ;
 wire \spiking_network_top_uut.all_data_out[523] ;
 wire \spiking_network_top_uut.all_data_out[524] ;
 wire \spiking_network_top_uut.all_data_out[525] ;
 wire \spiking_network_top_uut.all_data_out[526] ;
 wire \spiking_network_top_uut.all_data_out[527] ;
 wire \spiking_network_top_uut.all_data_out[528] ;
 wire \spiking_network_top_uut.all_data_out[529] ;
 wire \spiking_network_top_uut.all_data_out[52] ;
 wire \spiking_network_top_uut.all_data_out[530] ;
 wire \spiking_network_top_uut.all_data_out[531] ;
 wire \spiking_network_top_uut.all_data_out[532] ;
 wire \spiking_network_top_uut.all_data_out[533] ;
 wire \spiking_network_top_uut.all_data_out[534] ;
 wire \spiking_network_top_uut.all_data_out[535] ;
 wire \spiking_network_top_uut.all_data_out[536] ;
 wire \spiking_network_top_uut.all_data_out[537] ;
 wire \spiking_network_top_uut.all_data_out[538] ;
 wire \spiking_network_top_uut.all_data_out[539] ;
 wire \spiking_network_top_uut.all_data_out[53] ;
 wire \spiking_network_top_uut.all_data_out[540] ;
 wire \spiking_network_top_uut.all_data_out[541] ;
 wire \spiking_network_top_uut.all_data_out[542] ;
 wire \spiking_network_top_uut.all_data_out[543] ;
 wire \spiking_network_top_uut.all_data_out[544] ;
 wire \spiking_network_top_uut.all_data_out[545] ;
 wire \spiking_network_top_uut.all_data_out[546] ;
 wire \spiking_network_top_uut.all_data_out[547] ;
 wire \spiking_network_top_uut.all_data_out[548] ;
 wire \spiking_network_top_uut.all_data_out[549] ;
 wire \spiking_network_top_uut.all_data_out[54] ;
 wire \spiking_network_top_uut.all_data_out[550] ;
 wire \spiking_network_top_uut.all_data_out[551] ;
 wire \spiking_network_top_uut.all_data_out[552] ;
 wire \spiking_network_top_uut.all_data_out[553] ;
 wire \spiking_network_top_uut.all_data_out[554] ;
 wire \spiking_network_top_uut.all_data_out[555] ;
 wire \spiking_network_top_uut.all_data_out[556] ;
 wire \spiking_network_top_uut.all_data_out[557] ;
 wire \spiking_network_top_uut.all_data_out[558] ;
 wire \spiking_network_top_uut.all_data_out[559] ;
 wire \spiking_network_top_uut.all_data_out[55] ;
 wire \spiking_network_top_uut.all_data_out[560] ;
 wire \spiking_network_top_uut.all_data_out[561] ;
 wire \spiking_network_top_uut.all_data_out[562] ;
 wire \spiking_network_top_uut.all_data_out[563] ;
 wire \spiking_network_top_uut.all_data_out[564] ;
 wire \spiking_network_top_uut.all_data_out[565] ;
 wire \spiking_network_top_uut.all_data_out[566] ;
 wire \spiking_network_top_uut.all_data_out[567] ;
 wire \spiking_network_top_uut.all_data_out[568] ;
 wire \spiking_network_top_uut.all_data_out[569] ;
 wire \spiking_network_top_uut.all_data_out[56] ;
 wire \spiking_network_top_uut.all_data_out[570] ;
 wire \spiking_network_top_uut.all_data_out[571] ;
 wire \spiking_network_top_uut.all_data_out[572] ;
 wire \spiking_network_top_uut.all_data_out[573] ;
 wire \spiking_network_top_uut.all_data_out[574] ;
 wire \spiking_network_top_uut.all_data_out[575] ;
 wire \spiking_network_top_uut.all_data_out[576] ;
 wire \spiking_network_top_uut.all_data_out[577] ;
 wire \spiking_network_top_uut.all_data_out[578] ;
 wire \spiking_network_top_uut.all_data_out[579] ;
 wire \spiking_network_top_uut.all_data_out[57] ;
 wire \spiking_network_top_uut.all_data_out[580] ;
 wire \spiking_network_top_uut.all_data_out[581] ;
 wire \spiking_network_top_uut.all_data_out[582] ;
 wire \spiking_network_top_uut.all_data_out[583] ;
 wire \spiking_network_top_uut.all_data_out[584] ;
 wire \spiking_network_top_uut.all_data_out[585] ;
 wire \spiking_network_top_uut.all_data_out[586] ;
 wire \spiking_network_top_uut.all_data_out[587] ;
 wire \spiking_network_top_uut.all_data_out[588] ;
 wire \spiking_network_top_uut.all_data_out[589] ;
 wire \spiking_network_top_uut.all_data_out[58] ;
 wire \spiking_network_top_uut.all_data_out[590] ;
 wire \spiking_network_top_uut.all_data_out[591] ;
 wire \spiking_network_top_uut.all_data_out[592] ;
 wire \spiking_network_top_uut.all_data_out[593] ;
 wire \spiking_network_top_uut.all_data_out[594] ;
 wire \spiking_network_top_uut.all_data_out[595] ;
 wire \spiking_network_top_uut.all_data_out[596] ;
 wire \spiking_network_top_uut.all_data_out[597] ;
 wire \spiking_network_top_uut.all_data_out[598] ;
 wire \spiking_network_top_uut.all_data_out[599] ;
 wire \spiking_network_top_uut.all_data_out[59] ;
 wire \spiking_network_top_uut.all_data_out[5] ;
 wire \spiking_network_top_uut.all_data_out[600] ;
 wire \spiking_network_top_uut.all_data_out[601] ;
 wire \spiking_network_top_uut.all_data_out[602] ;
 wire \spiking_network_top_uut.all_data_out[603] ;
 wire \spiking_network_top_uut.all_data_out[604] ;
 wire \spiking_network_top_uut.all_data_out[605] ;
 wire \spiking_network_top_uut.all_data_out[606] ;
 wire \spiking_network_top_uut.all_data_out[607] ;
 wire \spiking_network_top_uut.all_data_out[608] ;
 wire \spiking_network_top_uut.all_data_out[609] ;
 wire \spiking_network_top_uut.all_data_out[60] ;
 wire \spiking_network_top_uut.all_data_out[610] ;
 wire \spiking_network_top_uut.all_data_out[611] ;
 wire \spiking_network_top_uut.all_data_out[612] ;
 wire \spiking_network_top_uut.all_data_out[613] ;
 wire \spiking_network_top_uut.all_data_out[614] ;
 wire \spiking_network_top_uut.all_data_out[615] ;
 wire \spiking_network_top_uut.all_data_out[616] ;
 wire \spiking_network_top_uut.all_data_out[617] ;
 wire \spiking_network_top_uut.all_data_out[618] ;
 wire \spiking_network_top_uut.all_data_out[619] ;
 wire \spiking_network_top_uut.all_data_out[61] ;
 wire \spiking_network_top_uut.all_data_out[620] ;
 wire \spiking_network_top_uut.all_data_out[621] ;
 wire \spiking_network_top_uut.all_data_out[622] ;
 wire \spiking_network_top_uut.all_data_out[623] ;
 wire \spiking_network_top_uut.all_data_out[624] ;
 wire \spiking_network_top_uut.all_data_out[625] ;
 wire \spiking_network_top_uut.all_data_out[626] ;
 wire \spiking_network_top_uut.all_data_out[627] ;
 wire \spiking_network_top_uut.all_data_out[628] ;
 wire \spiking_network_top_uut.all_data_out[629] ;
 wire \spiking_network_top_uut.all_data_out[62] ;
 wire \spiking_network_top_uut.all_data_out[630] ;
 wire \spiking_network_top_uut.all_data_out[631] ;
 wire \spiking_network_top_uut.all_data_out[632] ;
 wire \spiking_network_top_uut.all_data_out[633] ;
 wire \spiking_network_top_uut.all_data_out[634] ;
 wire \spiking_network_top_uut.all_data_out[635] ;
 wire \spiking_network_top_uut.all_data_out[636] ;
 wire \spiking_network_top_uut.all_data_out[637] ;
 wire \spiking_network_top_uut.all_data_out[638] ;
 wire \spiking_network_top_uut.all_data_out[639] ;
 wire \spiking_network_top_uut.all_data_out[63] ;
 wire \spiking_network_top_uut.all_data_out[640] ;
 wire \spiking_network_top_uut.all_data_out[641] ;
 wire \spiking_network_top_uut.all_data_out[642] ;
 wire \spiking_network_top_uut.all_data_out[643] ;
 wire \spiking_network_top_uut.all_data_out[644] ;
 wire \spiking_network_top_uut.all_data_out[645] ;
 wire \spiking_network_top_uut.all_data_out[646] ;
 wire \spiking_network_top_uut.all_data_out[647] ;
 wire \spiking_network_top_uut.all_data_out[648] ;
 wire \spiking_network_top_uut.all_data_out[649] ;
 wire \spiking_network_top_uut.all_data_out[64] ;
 wire \spiking_network_top_uut.all_data_out[650] ;
 wire \spiking_network_top_uut.all_data_out[651] ;
 wire \spiking_network_top_uut.all_data_out[652] ;
 wire \spiking_network_top_uut.all_data_out[653] ;
 wire \spiking_network_top_uut.all_data_out[654] ;
 wire \spiking_network_top_uut.all_data_out[655] ;
 wire \spiking_network_top_uut.all_data_out[656] ;
 wire \spiking_network_top_uut.all_data_out[657] ;
 wire \spiking_network_top_uut.all_data_out[658] ;
 wire \spiking_network_top_uut.all_data_out[659] ;
 wire \spiking_network_top_uut.all_data_out[65] ;
 wire \spiking_network_top_uut.all_data_out[660] ;
 wire \spiking_network_top_uut.all_data_out[661] ;
 wire \spiking_network_top_uut.all_data_out[662] ;
 wire \spiking_network_top_uut.all_data_out[663] ;
 wire \spiking_network_top_uut.all_data_out[664] ;
 wire \spiking_network_top_uut.all_data_out[665] ;
 wire \spiking_network_top_uut.all_data_out[666] ;
 wire \spiking_network_top_uut.all_data_out[667] ;
 wire \spiking_network_top_uut.all_data_out[668] ;
 wire \spiking_network_top_uut.all_data_out[669] ;
 wire \spiking_network_top_uut.all_data_out[66] ;
 wire \spiking_network_top_uut.all_data_out[670] ;
 wire \spiking_network_top_uut.all_data_out[671] ;
 wire \spiking_network_top_uut.all_data_out[672] ;
 wire \spiking_network_top_uut.all_data_out[673] ;
 wire \spiking_network_top_uut.all_data_out[674] ;
 wire \spiking_network_top_uut.all_data_out[675] ;
 wire \spiking_network_top_uut.all_data_out[676] ;
 wire \spiking_network_top_uut.all_data_out[677] ;
 wire \spiking_network_top_uut.all_data_out[678] ;
 wire \spiking_network_top_uut.all_data_out[679] ;
 wire \spiking_network_top_uut.all_data_out[67] ;
 wire \spiking_network_top_uut.all_data_out[680] ;
 wire \spiking_network_top_uut.all_data_out[681] ;
 wire \spiking_network_top_uut.all_data_out[682] ;
 wire \spiking_network_top_uut.all_data_out[683] ;
 wire \spiking_network_top_uut.all_data_out[684] ;
 wire \spiking_network_top_uut.all_data_out[685] ;
 wire \spiking_network_top_uut.all_data_out[686] ;
 wire \spiking_network_top_uut.all_data_out[687] ;
 wire \spiking_network_top_uut.all_data_out[688] ;
 wire \spiking_network_top_uut.all_data_out[689] ;
 wire \spiking_network_top_uut.all_data_out[68] ;
 wire \spiking_network_top_uut.all_data_out[690] ;
 wire \spiking_network_top_uut.all_data_out[691] ;
 wire \spiking_network_top_uut.all_data_out[692] ;
 wire \spiking_network_top_uut.all_data_out[693] ;
 wire \spiking_network_top_uut.all_data_out[694] ;
 wire \spiking_network_top_uut.all_data_out[695] ;
 wire \spiking_network_top_uut.all_data_out[696] ;
 wire \spiking_network_top_uut.all_data_out[697] ;
 wire \spiking_network_top_uut.all_data_out[698] ;
 wire \spiking_network_top_uut.all_data_out[699] ;
 wire \spiking_network_top_uut.all_data_out[69] ;
 wire \spiking_network_top_uut.all_data_out[6] ;
 wire \spiking_network_top_uut.all_data_out[700] ;
 wire \spiking_network_top_uut.all_data_out[701] ;
 wire \spiking_network_top_uut.all_data_out[702] ;
 wire \spiking_network_top_uut.all_data_out[703] ;
 wire \spiking_network_top_uut.all_data_out[704] ;
 wire \spiking_network_top_uut.all_data_out[705] ;
 wire \spiking_network_top_uut.all_data_out[706] ;
 wire \spiking_network_top_uut.all_data_out[707] ;
 wire \spiking_network_top_uut.all_data_out[708] ;
 wire \spiking_network_top_uut.all_data_out[709] ;
 wire \spiking_network_top_uut.all_data_out[70] ;
 wire \spiking_network_top_uut.all_data_out[710] ;
 wire \spiking_network_top_uut.all_data_out[711] ;
 wire \spiking_network_top_uut.all_data_out[712] ;
 wire \spiking_network_top_uut.all_data_out[713] ;
 wire \spiking_network_top_uut.all_data_out[714] ;
 wire \spiking_network_top_uut.all_data_out[715] ;
 wire \spiking_network_top_uut.all_data_out[716] ;
 wire \spiking_network_top_uut.all_data_out[717] ;
 wire \spiking_network_top_uut.all_data_out[718] ;
 wire \spiking_network_top_uut.all_data_out[719] ;
 wire \spiking_network_top_uut.all_data_out[71] ;
 wire \spiking_network_top_uut.all_data_out[720] ;
 wire \spiking_network_top_uut.all_data_out[721] ;
 wire \spiking_network_top_uut.all_data_out[722] ;
 wire \spiking_network_top_uut.all_data_out[723] ;
 wire \spiking_network_top_uut.all_data_out[724] ;
 wire \spiking_network_top_uut.all_data_out[725] ;
 wire \spiking_network_top_uut.all_data_out[726] ;
 wire \spiking_network_top_uut.all_data_out[727] ;
 wire \spiking_network_top_uut.all_data_out[728] ;
 wire \spiking_network_top_uut.all_data_out[729] ;
 wire \spiking_network_top_uut.all_data_out[72] ;
 wire \spiking_network_top_uut.all_data_out[730] ;
 wire \spiking_network_top_uut.all_data_out[731] ;
 wire \spiking_network_top_uut.all_data_out[732] ;
 wire \spiking_network_top_uut.all_data_out[733] ;
 wire \spiking_network_top_uut.all_data_out[734] ;
 wire \spiking_network_top_uut.all_data_out[735] ;
 wire \spiking_network_top_uut.all_data_out[736] ;
 wire \spiking_network_top_uut.all_data_out[737] ;
 wire \spiking_network_top_uut.all_data_out[738] ;
 wire \spiking_network_top_uut.all_data_out[739] ;
 wire \spiking_network_top_uut.all_data_out[73] ;
 wire \spiking_network_top_uut.all_data_out[740] ;
 wire \spiking_network_top_uut.all_data_out[741] ;
 wire \spiking_network_top_uut.all_data_out[742] ;
 wire \spiking_network_top_uut.all_data_out[743] ;
 wire \spiking_network_top_uut.all_data_out[744] ;
 wire \spiking_network_top_uut.all_data_out[745] ;
 wire \spiking_network_top_uut.all_data_out[746] ;
 wire \spiking_network_top_uut.all_data_out[747] ;
 wire \spiking_network_top_uut.all_data_out[748] ;
 wire \spiking_network_top_uut.all_data_out[749] ;
 wire \spiking_network_top_uut.all_data_out[74] ;
 wire \spiking_network_top_uut.all_data_out[750] ;
 wire \spiking_network_top_uut.all_data_out[751] ;
 wire \spiking_network_top_uut.all_data_out[752] ;
 wire \spiking_network_top_uut.all_data_out[753] ;
 wire \spiking_network_top_uut.all_data_out[754] ;
 wire \spiking_network_top_uut.all_data_out[755] ;
 wire \spiking_network_top_uut.all_data_out[756] ;
 wire \spiking_network_top_uut.all_data_out[757] ;
 wire \spiking_network_top_uut.all_data_out[758] ;
 wire \spiking_network_top_uut.all_data_out[759] ;
 wire \spiking_network_top_uut.all_data_out[75] ;
 wire \spiking_network_top_uut.all_data_out[760] ;
 wire \spiking_network_top_uut.all_data_out[761] ;
 wire \spiking_network_top_uut.all_data_out[762] ;
 wire \spiking_network_top_uut.all_data_out[763] ;
 wire \spiking_network_top_uut.all_data_out[764] ;
 wire \spiking_network_top_uut.all_data_out[765] ;
 wire \spiking_network_top_uut.all_data_out[766] ;
 wire \spiking_network_top_uut.all_data_out[767] ;
 wire \spiking_network_top_uut.all_data_out[768] ;
 wire \spiking_network_top_uut.all_data_out[769] ;
 wire \spiking_network_top_uut.all_data_out[76] ;
 wire \spiking_network_top_uut.all_data_out[770] ;
 wire \spiking_network_top_uut.all_data_out[771] ;
 wire \spiking_network_top_uut.all_data_out[772] ;
 wire \spiking_network_top_uut.all_data_out[773] ;
 wire \spiking_network_top_uut.all_data_out[774] ;
 wire \spiking_network_top_uut.all_data_out[775] ;
 wire \spiking_network_top_uut.all_data_out[776] ;
 wire \spiking_network_top_uut.all_data_out[777] ;
 wire \spiking_network_top_uut.all_data_out[778] ;
 wire \spiking_network_top_uut.all_data_out[779] ;
 wire \spiking_network_top_uut.all_data_out[77] ;
 wire \spiking_network_top_uut.all_data_out[780] ;
 wire \spiking_network_top_uut.all_data_out[781] ;
 wire \spiking_network_top_uut.all_data_out[782] ;
 wire \spiking_network_top_uut.all_data_out[783] ;
 wire \spiking_network_top_uut.all_data_out[784] ;
 wire \spiking_network_top_uut.all_data_out[785] ;
 wire \spiking_network_top_uut.all_data_out[786] ;
 wire \spiking_network_top_uut.all_data_out[787] ;
 wire \spiking_network_top_uut.all_data_out[788] ;
 wire \spiking_network_top_uut.all_data_out[789] ;
 wire \spiking_network_top_uut.all_data_out[78] ;
 wire \spiking_network_top_uut.all_data_out[790] ;
 wire \spiking_network_top_uut.all_data_out[791] ;
 wire \spiking_network_top_uut.all_data_out[792] ;
 wire \spiking_network_top_uut.all_data_out[793] ;
 wire \spiking_network_top_uut.all_data_out[794] ;
 wire \spiking_network_top_uut.all_data_out[795] ;
 wire \spiking_network_top_uut.all_data_out[796] ;
 wire \spiking_network_top_uut.all_data_out[797] ;
 wire \spiking_network_top_uut.all_data_out[798] ;
 wire \spiking_network_top_uut.all_data_out[799] ;
 wire \spiking_network_top_uut.all_data_out[79] ;
 wire \spiking_network_top_uut.all_data_out[7] ;
 wire \spiking_network_top_uut.all_data_out[800] ;
 wire \spiking_network_top_uut.all_data_out[801] ;
 wire \spiking_network_top_uut.all_data_out[802] ;
 wire \spiking_network_top_uut.all_data_out[803] ;
 wire \spiking_network_top_uut.all_data_out[804] ;
 wire \spiking_network_top_uut.all_data_out[805] ;
 wire \spiking_network_top_uut.all_data_out[806] ;
 wire \spiking_network_top_uut.all_data_out[807] ;
 wire \spiking_network_top_uut.all_data_out[808] ;
 wire \spiking_network_top_uut.all_data_out[809] ;
 wire \spiking_network_top_uut.all_data_out[80] ;
 wire \spiking_network_top_uut.all_data_out[810] ;
 wire \spiking_network_top_uut.all_data_out[811] ;
 wire \spiking_network_top_uut.all_data_out[812] ;
 wire \spiking_network_top_uut.all_data_out[813] ;
 wire \spiking_network_top_uut.all_data_out[814] ;
 wire \spiking_network_top_uut.all_data_out[815] ;
 wire \spiking_network_top_uut.all_data_out[816] ;
 wire \spiking_network_top_uut.all_data_out[817] ;
 wire \spiking_network_top_uut.all_data_out[818] ;
 wire \spiking_network_top_uut.all_data_out[819] ;
 wire \spiking_network_top_uut.all_data_out[81] ;
 wire \spiking_network_top_uut.all_data_out[820] ;
 wire \spiking_network_top_uut.all_data_out[821] ;
 wire \spiking_network_top_uut.all_data_out[822] ;
 wire \spiking_network_top_uut.all_data_out[823] ;
 wire \spiking_network_top_uut.all_data_out[824] ;
 wire \spiking_network_top_uut.all_data_out[825] ;
 wire \spiking_network_top_uut.all_data_out[826] ;
 wire \spiking_network_top_uut.all_data_out[827] ;
 wire \spiking_network_top_uut.all_data_out[828] ;
 wire \spiking_network_top_uut.all_data_out[829] ;
 wire \spiking_network_top_uut.all_data_out[82] ;
 wire \spiking_network_top_uut.all_data_out[830] ;
 wire \spiking_network_top_uut.all_data_out[831] ;
 wire \spiking_network_top_uut.all_data_out[832] ;
 wire \spiking_network_top_uut.all_data_out[833] ;
 wire \spiking_network_top_uut.all_data_out[834] ;
 wire \spiking_network_top_uut.all_data_out[835] ;
 wire \spiking_network_top_uut.all_data_out[836] ;
 wire \spiking_network_top_uut.all_data_out[837] ;
 wire \spiking_network_top_uut.all_data_out[838] ;
 wire \spiking_network_top_uut.all_data_out[839] ;
 wire \spiking_network_top_uut.all_data_out[83] ;
 wire \spiking_network_top_uut.all_data_out[840] ;
 wire \spiking_network_top_uut.all_data_out[841] ;
 wire \spiking_network_top_uut.all_data_out[842] ;
 wire \spiking_network_top_uut.all_data_out[843] ;
 wire \spiking_network_top_uut.all_data_out[844] ;
 wire \spiking_network_top_uut.all_data_out[845] ;
 wire \spiking_network_top_uut.all_data_out[846] ;
 wire \spiking_network_top_uut.all_data_out[847] ;
 wire \spiking_network_top_uut.all_data_out[848] ;
 wire \spiking_network_top_uut.all_data_out[849] ;
 wire \spiking_network_top_uut.all_data_out[84] ;
 wire \spiking_network_top_uut.all_data_out[850] ;
 wire \spiking_network_top_uut.all_data_out[851] ;
 wire \spiking_network_top_uut.all_data_out[852] ;
 wire \spiking_network_top_uut.all_data_out[853] ;
 wire \spiking_network_top_uut.all_data_out[854] ;
 wire \spiking_network_top_uut.all_data_out[855] ;
 wire \spiking_network_top_uut.all_data_out[856] ;
 wire \spiking_network_top_uut.all_data_out[857] ;
 wire \spiking_network_top_uut.all_data_out[858] ;
 wire \spiking_network_top_uut.all_data_out[859] ;
 wire \spiking_network_top_uut.all_data_out[85] ;
 wire \spiking_network_top_uut.all_data_out[860] ;
 wire \spiking_network_top_uut.all_data_out[861] ;
 wire \spiking_network_top_uut.all_data_out[862] ;
 wire \spiking_network_top_uut.all_data_out[863] ;
 wire \spiking_network_top_uut.all_data_out[864] ;
 wire \spiking_network_top_uut.all_data_out[865] ;
 wire \spiking_network_top_uut.all_data_out[866] ;
 wire \spiking_network_top_uut.all_data_out[867] ;
 wire \spiking_network_top_uut.all_data_out[868] ;
 wire \spiking_network_top_uut.all_data_out[869] ;
 wire \spiking_network_top_uut.all_data_out[86] ;
 wire \spiking_network_top_uut.all_data_out[870] ;
 wire \spiking_network_top_uut.all_data_out[871] ;
 wire \spiking_network_top_uut.all_data_out[872] ;
 wire \spiking_network_top_uut.all_data_out[873] ;
 wire \spiking_network_top_uut.all_data_out[874] ;
 wire \spiking_network_top_uut.all_data_out[875] ;
 wire \spiking_network_top_uut.all_data_out[876] ;
 wire \spiking_network_top_uut.all_data_out[877] ;
 wire \spiking_network_top_uut.all_data_out[878] ;
 wire \spiking_network_top_uut.all_data_out[879] ;
 wire \spiking_network_top_uut.all_data_out[87] ;
 wire \spiking_network_top_uut.all_data_out[880] ;
 wire \spiking_network_top_uut.all_data_out[881] ;
 wire \spiking_network_top_uut.all_data_out[882] ;
 wire \spiking_network_top_uut.all_data_out[883] ;
 wire \spiking_network_top_uut.all_data_out[884] ;
 wire \spiking_network_top_uut.all_data_out[885] ;
 wire \spiking_network_top_uut.all_data_out[886] ;
 wire \spiking_network_top_uut.all_data_out[887] ;
 wire \spiking_network_top_uut.all_data_out[888] ;
 wire \spiking_network_top_uut.all_data_out[889] ;
 wire \spiking_network_top_uut.all_data_out[88] ;
 wire \spiking_network_top_uut.all_data_out[890] ;
 wire \spiking_network_top_uut.all_data_out[891] ;
 wire \spiking_network_top_uut.all_data_out[892] ;
 wire \spiking_network_top_uut.all_data_out[893] ;
 wire \spiking_network_top_uut.all_data_out[894] ;
 wire \spiking_network_top_uut.all_data_out[895] ;
 wire \spiking_network_top_uut.all_data_out[896] ;
 wire \spiking_network_top_uut.all_data_out[897] ;
 wire \spiking_network_top_uut.all_data_out[898] ;
 wire \spiking_network_top_uut.all_data_out[899] ;
 wire \spiking_network_top_uut.all_data_out[89] ;
 wire \spiking_network_top_uut.all_data_out[8] ;
 wire \spiking_network_top_uut.all_data_out[900] ;
 wire \spiking_network_top_uut.all_data_out[901] ;
 wire \spiking_network_top_uut.all_data_out[902] ;
 wire \spiking_network_top_uut.all_data_out[903] ;
 wire \spiking_network_top_uut.all_data_out[90] ;
 wire \spiking_network_top_uut.all_data_out[91] ;
 wire \spiking_network_top_uut.all_data_out[92] ;
 wire \spiking_network_top_uut.all_data_out[93] ;
 wire \spiking_network_top_uut.all_data_out[94] ;
 wire \spiking_network_top_uut.all_data_out[95] ;
 wire \spiking_network_top_uut.all_data_out[96] ;
 wire \spiking_network_top_uut.all_data_out[97] ;
 wire \spiking_network_top_uut.all_data_out[98] ;
 wire \spiking_network_top_uut.all_data_out[99] ;
 wire \spiking_network_top_uut.all_data_out[9] ;
 wire \spiking_network_top_uut.clk_div_inst.clk_out ;
 wire \spiking_network_top_uut.clk_div_inst.counter[0] ;
 wire \spiking_network_top_uut.clk_div_inst.counter[1] ;
 wire \spiking_network_top_uut.clk_div_inst.counter[2] ;
 wire \spiking_network_top_uut.clk_div_inst.counter[3] ;
 wire \spiking_network_top_uut.clk_div_inst.counter[4] ;
 wire \spiking_network_top_uut.clk_div_inst.counter[5] ;
 wire \spiking_network_top_uut.clk_div_inst.counter[6] ;
 wire \spiking_network_top_uut.clk_div_inst.counter[7] ;
 wire \spiking_network_top_uut.clk_div_inst.enable ;
 wire \spiking_network_top_uut.clk_div_ready_reg_out ;
 wire \spiking_network_top_uut.clk_div_sync.sync_ff1 ;
 wire \spiking_network_top_uut.data_valid_out ;
 wire \spiking_network_top_uut.debug_config_ready_reg_out ;
 wire \spiking_network_top_uut.debug_config_ready_sync ;
 wire \spiking_network_top_uut.debug_config_sync.sync_ff1 ;
 wire \spiking_network_top_uut.debug_inst.debug_config[0] ;
 wire \spiking_network_top_uut.debug_inst.debug_config[1] ;
 wire \spiking_network_top_uut.debug_inst.debug_config[2] ;
 wire \spiking_network_top_uut.debug_inst.debug_config[3] ;
 wire \spiking_network_top_uut.debug_inst.debug_config[4] ;
 wire \spiking_network_top_uut.debug_inst.debug_config[5] ;
 wire \spiking_network_top_uut.debug_inst.debug_config[6] ;
 wire \spiking_network_top_uut.debug_inst.debug_config[7] ;
 wire \spiking_network_top_uut.input_ready_sync ;
 wire \spiking_network_top_uut.input_ready_sync_inst.sync_ff1 ;
 wire \spiking_network_top_uut.output_data_ready ;
 wire \spiking_network_top_uut.snn_en_sync_inst.sync_ff1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.enable_LYR_2 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.enable_LYR_3 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[0] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[0] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[1] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[2] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[3] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[4] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.spike_out ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.din ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[0] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[1] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[2] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[3] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[4] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[5] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[6] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[7] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.din ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[0] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[1] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[2] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[3] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[4] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[5] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[6] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[7] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.din ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[0] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[1] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[2] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[3] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[4] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[5] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[6] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[7] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.din ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[0] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[1] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[2] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[3] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[4] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[5] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[6] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[7] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.din ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[0] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[1] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[2] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[3] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[4] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[5] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[6] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[7] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.din ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[0] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[1] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[2] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[3] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[4] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[5] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[6] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[7] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.din ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[0] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[1] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[2] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[3] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[4] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[5] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[6] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[7] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.din ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[0] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[1] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[2] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[3] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[4] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[5] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[6] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[7] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[0] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[0] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[1] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[2] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[3] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[4] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.spike_out ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[0] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[0] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[1] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[2] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[3] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[4] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.spike_out ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[0] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[0] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[1] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[2] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[3] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[4] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.spike_out ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[0] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[0] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[1] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[2] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[3] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[4] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.spike_out ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[0] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[0] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[1] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[2] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[3] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[4] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.spike_out ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[0] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[0] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[1] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[2] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[3] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[4] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.spike_out ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[0] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[0] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[1] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[2] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[3] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[4] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.spike_out ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[0] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[0] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[1] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[2] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[3] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[4] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.spike_out ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[0] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[1] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[2] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[3] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[4] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[5] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[6] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[7] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[0] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[1] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[2] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[3] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[4] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[5] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[6] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[7] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[0] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[1] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[2] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[3] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[4] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[5] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[6] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[7] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[0] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[1] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[2] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[3] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[4] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[5] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[6] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[7] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[0] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[1] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[2] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[3] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[4] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[5] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[6] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[7] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[0] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[1] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[2] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[3] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[4] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[5] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[6] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[7] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[0] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[1] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[2] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[3] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[4] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[5] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[6] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[7] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[0] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[1] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[2] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[3] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[4] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[5] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[6] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[7] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[0] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[0] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[1] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[2] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[3] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[4] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.spike_out ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[0] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[0] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[1] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[2] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[3] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[4] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.spike_out ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[0] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[0] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[1] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[2] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[3] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[4] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.spike_out ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[0] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[0] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[1] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[2] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[3] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[4] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.spike_out ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[0] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[0] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[1] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[2] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[3] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[4] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.spike_out ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[0] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[0] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[1] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[2] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[3] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[4] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.spike_out ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[0] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[0] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[1] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[2] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[3] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[4] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.spike_out ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[0] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[0] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[1] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[2] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[3] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[4] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.spike_out ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[0] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[1] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[2] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[3] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[4] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[5] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[6] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[7] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[0] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[1] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[2] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[3] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[4] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[5] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[6] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[7] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[0] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[1] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[2] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[3] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[4] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[5] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[6] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[7] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[0] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[1] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[2] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[3] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[4] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[5] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[6] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[7] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[0] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[1] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[2] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[3] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[4] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[5] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[6] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[7] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[0] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[1] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[2] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[3] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[4] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[5] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[6] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[7] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[0] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[1] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[2] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[3] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[4] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[5] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[6] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[7] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[0] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[1] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[2] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[3] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[4] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[5] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[6] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[7] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[0] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[0] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[1] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[2] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[3] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[4] ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.spike_out ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[1].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[1].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[1].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[1].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[1].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[1].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[1].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[1].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[1].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[1].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[1].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[1].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[1].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[1].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[1].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_dout ;
 wire \spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[1].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_reg1 ;
 wire \spiking_network_top_uut.spi_inst.LSB_Address_reg[0] ;
 wire \spiking_network_top_uut.spi_inst.LSB_Address_reg[1] ;
 wire \spiking_network_top_uut.spi_inst.LSB_Address_reg[2] ;
 wire \spiking_network_top_uut.spi_inst.LSB_Address_reg[3] ;
 wire \spiking_network_top_uut.spi_inst.LSB_Address_reg[4] ;
 wire \spiking_network_top_uut.spi_inst.LSB_Address_reg[5] ;
 wire \spiking_network_top_uut.spi_inst.LSB_Address_reg[6] ;
 wire \spiking_network_top_uut.spi_inst.SPI_address_LSB_reg_en ;
 wire \spiking_network_top_uut.spi_inst.SPI_instruction_reg[0] ;
 wire \spiking_network_top_uut.spi_inst.SPI_instruction_reg[1] ;
 wire \spiking_network_top_uut.spi_inst.SPI_instruction_reg[2] ;
 wire \spiking_network_top_uut.spi_inst.SPI_instruction_reg[3] ;
 wire \spiking_network_top_uut.spi_inst.SPI_instruction_reg[4] ;
 wire \spiking_network_top_uut.spi_inst.SPI_instruction_reg[5] ;
 wire \spiking_network_top_uut.spi_inst.SPI_instruction_reg[6] ;
 wire \spiking_network_top_uut.spi_inst.SPI_instruction_reg[7] ;
 wire \spiking_network_top_uut.spi_inst.SPI_instruction_reg_en ;
 wire \spiking_network_top_uut.spi_inst.SPI_instruction_reg_in[0] ;
 wire \spiking_network_top_uut.spi_inst.SPI_instruction_reg_in[1] ;
 wire \spiking_network_top_uut.spi_inst.SPI_instruction_reg_in[2] ;
 wire \spiking_network_top_uut.spi_inst.SPI_instruction_reg_in[3] ;
 wire \spiking_network_top_uut.spi_inst.SPI_instruction_reg_in[4] ;
 wire \spiking_network_top_uut.spi_inst.SPI_instruction_reg_in[5] ;
 wire \spiking_network_top_uut.spi_inst.SPI_instruction_reg_in[6] ;
 wire \spiking_network_top_uut.spi_inst.SPI_instruction_reg_in[7] ;
 wire \spiking_network_top_uut.spi_inst.clk_div_ready_reg_en ;
 wire \spiking_network_top_uut.spi_inst.clk_div_ready_reg_in ;
 wire \spiking_network_top_uut.spi_inst.debug_config_ready_reg_en ;
 wire \spiking_network_top_uut.spi_inst.debug_config_ready_reg_in ;
 wire \spiking_network_top_uut.spi_inst.memory_inst.addr_reg_out[0] ;
 wire \spiking_network_top_uut.spi_inst.memory_inst.addr_reg_out[1] ;
 wire \spiking_network_top_uut.spi_inst.memory_inst.addr_reg_out[2] ;
 wire \spiking_network_top_uut.spi_inst.memory_inst.addr_reg_out[3] ;
 wire \spiking_network_top_uut.spi_inst.memory_inst.addr_reg_out[4] ;
 wire \spiking_network_top_uut.spi_inst.memory_inst.addr_reg_out[5] ;
 wire \spiking_network_top_uut.spi_inst.memory_inst.addr_reg_out[6] ;
 wire \spiking_network_top_uut.spi_inst.memory_inst.write_enable ;
 wire \spiking_network_top_uut.spi_inst.spi_control_unit_inst.current_state[0] ;
 wire \spiking_network_top_uut.spi_inst.spi_control_unit_inst.current_state[1] ;
 wire \spiking_network_top_uut.spi_inst.spi_control_unit_inst.current_state[2] ;
 wire \spiking_network_top_uut.spi_inst.spi_slave_inst.bit_cnt[0] ;
 wire \spiking_network_top_uut.spi_inst.spi_slave_inst.bit_cnt[1] ;
 wire \spiking_network_top_uut.spi_inst.spi_slave_inst.bit_cnt[2] ;
 wire \spiking_network_top_uut.spi_inst.spi_slave_inst.shift_reg[0] ;
 wire \spiking_network_top_uut.spi_inst.spi_slave_inst.shift_reg[1] ;
 wire \spiking_network_top_uut.spi_inst.spi_slave_inst.shift_reg[2] ;
 wire \spiking_network_top_uut.spi_inst.spi_slave_inst.shift_reg[3] ;
 wire \spiking_network_top_uut.spi_inst.spi_slave_inst.shift_reg[4] ;
 wire \spiking_network_top_uut.spi_inst.spi_slave_inst.shift_reg[5] ;
 wire \spiking_network_top_uut.spi_inst.spi_slave_inst.shift_reg[6] ;
 wire \spiking_network_top_uut.sys_clk_reset_synchr ;
 wire \spiking_network_top_uut.u_SPI_reset.reset_ff1 ;
 wire \spiking_network_top_uut.u_sys_clk_reset.reset_ff1 ;
 wire net17;
 wire net18;
 wire net29;
 wire net19;
 wire net20;
 wire net30;
 wire net21;
 wire clknet_leaf_0_clk;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net3616;
 wire net3617;
 wire net3618;
 wire net3619;
 wire net3620;
 wire net3621;
 wire net3622;
 wire net3623;
 wire net3624;
 wire net3625;
 wire net3626;
 wire net3627;
 wire net3628;
 wire net3629;
 wire net3630;
 wire net3631;
 wire net3632;
 wire net3633;
 wire net3634;
 wire net3635;
 wire net3636;
 wire net3637;
 wire net3638;
 wire net3639;
 wire net3640;
 wire net3641;
 wire net3642;
 wire net3643;
 wire net3644;
 wire net3645;
 wire net3646;
 wire net3647;
 wire net3648;
 wire net3649;
 wire net3650;
 wire net3651;
 wire net3652;
 wire net3653;
 wire net3654;
 wire net3655;
 wire net3656;
 wire net3657;
 wire net3658;
 wire net3659;
 wire net3660;
 wire net3661;
 wire net3662;
 wire net3663;
 wire net3664;
 wire net3665;
 wire net3666;
 wire net3667;
 wire net3668;
 wire net3669;
 wire net3670;
 wire net3671;
 wire net3672;
 wire net3673;
 wire net3674;
 wire net3675;
 wire net3676;
 wire net3677;
 wire net3678;
 wire net3679;
 wire net3680;
 wire net3681;
 wire net3682;
 wire net3683;
 wire net3684;
 wire net3685;
 wire net3686;
 wire net3687;
 wire net3688;
 wire net3689;
 wire net3690;
 wire net3691;
 wire net3692;
 wire net3693;
 wire net3694;
 wire net3695;
 wire net3696;
 wire net3697;
 wire net3698;
 wire net3699;
 wire net3700;
 wire net3701;
 wire net3702;
 wire net3703;
 wire net3704;
 wire net3705;
 wire net3706;
 wire net3707;
 wire net3708;
 wire net3709;
 wire net3710;
 wire net3711;
 wire net3712;
 wire net3713;
 wire net3714;
 wire net3715;
 wire net3716;
 wire net3717;
 wire net3718;
 wire net3719;
 wire net3720;
 wire net3721;
 wire net3722;
 wire net3723;
 wire net3724;
 wire net3725;
 wire net3726;
 wire net3727;
 wire net3728;
 wire net3729;
 wire net3730;
 wire net3731;
 wire net3732;
 wire net3733;
 wire net3734;
 wire net3735;
 wire net3736;
 wire net3737;
 wire net3738;
 wire net3739;
 wire net3740;
 wire net3741;
 wire net3742;
 wire net3743;
 wire net3744;
 wire net3745;
 wire net3746;
 wire net3747;
 wire net3748;
 wire net3749;
 wire net3750;
 wire net3751;
 wire net3752;
 wire net3753;
 wire net3754;
 wire net3755;
 wire net3756;
 wire net3757;
 wire net3758;
 wire net3759;
 wire net3760;
 wire net3761;
 wire net3762;
 wire net3763;
 wire net3764;
 wire net3765;
 wire net3766;
 wire net3767;
 wire net3768;
 wire net3769;
 wire net3770;
 wire net3771;
 wire net3772;
 wire net3773;
 wire net3774;
 wire net3775;
 wire net3776;
 wire net3777;
 wire net3778;
 wire net3779;
 wire net3780;
 wire net3781;
 wire net3782;
 wire net3783;
 wire net3784;
 wire net3785;
 wire net3786;
 wire net3787;
 wire net3788;
 wire net3789;
 wire net3790;
 wire net3791;
 wire net3792;
 wire net3793;
 wire net3794;
 wire net3795;
 wire net3796;
 wire net3797;
 wire net3798;
 wire net3799;
 wire net3800;
 wire net3801;
 wire net3802;
 wire net3803;
 wire net3804;
 wire net3805;
 wire net3806;
 wire net3807;
 wire net3808;
 wire net3809;
 wire net3810;
 wire net3811;
 wire net3812;
 wire net3813;
 wire net3814;
 wire net3815;
 wire net3816;
 wire net3817;
 wire net3818;
 wire net3819;
 wire net3820;
 wire net3821;
 wire net3822;
 wire net3823;
 wire net3824;
 wire net3825;
 wire net3826;
 wire net3827;
 wire net3828;
 wire net3829;
 wire net3830;
 wire net3831;
 wire net3832;
 wire net3833;
 wire net3834;
 wire net3835;
 wire net3836;
 wire net3837;
 wire net3838;
 wire net3839;
 wire net3840;
 wire net3841;
 wire net3842;
 wire net3843;
 wire net3844;
 wire net3845;
 wire net3846;
 wire net3847;
 wire net3848;
 wire net3849;
 wire net3850;
 wire net3851;
 wire net3852;
 wire net3853;
 wire net3854;
 wire net3855;
 wire net3856;
 wire net3857;
 wire net3858;
 wire net3859;
 wire net3860;
 wire net3861;
 wire net3862;
 wire net3863;
 wire net3864;
 wire net3865;
 wire net3866;
 wire net3867;
 wire net3868;
 wire net3869;
 wire net3870;
 wire net3871;
 wire net3872;
 wire net3873;
 wire net3874;
 wire net3875;
 wire net3876;
 wire net3877;
 wire net3878;
 wire net3879;
 wire net3880;
 wire net3881;
 wire net3882;
 wire net3883;
 wire net3884;
 wire net3885;
 wire net3886;
 wire net3887;
 wire net3888;
 wire net3889;
 wire net3890;
 wire net3891;
 wire net3892;
 wire net3893;
 wire net3894;
 wire net3895;
 wire net3896;
 wire net3897;
 wire net3898;
 wire net3899;
 wire net3900;
 wire net3901;
 wire net3902;
 wire net3903;
 wire net3904;
 wire net3905;
 wire net3906;
 wire net3907;
 wire net3908;
 wire net3909;
 wire net3910;
 wire net3911;
 wire net3912;
 wire net3913;
 wire net3914;
 wire net3915;
 wire net3916;
 wire net3917;
 wire net3918;
 wire net3919;
 wire net3920;
 wire net3921;
 wire net3922;
 wire net3923;
 wire net3924;
 wire net3925;
 wire net3926;
 wire net3927;
 wire net3928;
 wire net3929;
 wire net3930;
 wire net3931;
 wire net3932;
 wire net3933;
 wire net3934;
 wire net3935;
 wire net3936;
 wire net3937;
 wire net3938;
 wire net3939;
 wire net3940;
 wire net3941;
 wire net3942;
 wire net3943;
 wire net3944;
 wire net3945;
 wire net3946;
 wire net3947;
 wire net3948;
 wire net3949;
 wire net3950;
 wire net3951;
 wire net3952;
 wire net3953;
 wire net3954;
 wire net3955;
 wire net3956;
 wire net3957;
 wire net3958;
 wire net3959;
 wire net3960;
 wire net3961;
 wire net3962;
 wire net3963;
 wire net3964;
 wire net3965;
 wire net3966;
 wire net3967;
 wire net3968;
 wire net3969;
 wire net3970;
 wire net3971;
 wire net3972;
 wire net3973;
 wire net3974;
 wire net3975;
 wire net3976;
 wire net3977;
 wire net3978;
 wire net3979;
 wire net3980;
 wire net3981;
 wire net3982;
 wire net3983;
 wire net3984;
 wire net3985;
 wire net3986;
 wire net3987;
 wire net3988;
 wire net3989;
 wire net3990;
 wire net3991;
 wire net3992;
 wire net3993;
 wire net3994;
 wire net3995;
 wire net3996;
 wire net3997;
 wire net3998;
 wire net3999;
 wire net4000;
 wire net4001;
 wire net4002;
 wire net4003;
 wire net4004;
 wire net4005;
 wire net4006;
 wire net4007;
 wire net4008;
 wire net4009;
 wire net4010;
 wire net4011;
 wire net4012;
 wire net4013;
 wire net4014;
 wire net4015;
 wire net4016;
 wire net4017;
 wire net4018;
 wire net4019;
 wire net4020;
 wire net4021;
 wire net4022;
 wire net4023;
 wire net4024;
 wire net4025;
 wire net4026;
 wire net4027;
 wire net4028;
 wire net4029;
 wire net4030;
 wire net4031;
 wire net4032;
 wire net4033;
 wire net4034;
 wire net4035;
 wire net4036;
 wire net4037;
 wire net4038;
 wire net4039;
 wire net4040;
 wire net4041;
 wire net4042;
 wire net4043;
 wire net4044;
 wire net4045;
 wire net4046;
 wire net4047;
 wire net4048;
 wire net4049;
 wire net4050;
 wire net4051;
 wire net4052;
 wire net4053;
 wire net4054;
 wire net4055;
 wire net4056;
 wire net4057;
 wire net4058;
 wire net4059;
 wire net4060;
 wire net4061;
 wire net4062;
 wire net4063;
 wire net4064;
 wire net4065;
 wire net4066;
 wire net4067;
 wire net4068;
 wire net4069;
 wire net4070;
 wire net4071;
 wire net4072;
 wire net4073;
 wire net4074;
 wire net4075;
 wire net4076;
 wire net4077;
 wire net4078;
 wire net4079;
 wire net4080;
 wire net4081;
 wire net4082;
 wire net4083;
 wire net4084;
 wire net4085;
 wire net4086;
 wire net4087;
 wire net4088;
 wire net4089;
 wire net4090;
 wire net4091;
 wire net4092;
 wire net4093;
 wire net4094;
 wire net4095;
 wire net4096;
 wire net4097;
 wire net4098;
 wire net4099;
 wire net4100;
 wire net4101;
 wire net4102;
 wire net4103;
 wire net4104;
 wire net4105;
 wire net4106;
 wire net4107;
 wire net4108;
 wire net4109;
 wire net4110;
 wire net4111;
 wire net4112;
 wire net4113;
 wire net4114;
 wire net4115;
 wire net4116;
 wire net4117;
 wire net4118;
 wire net4119;
 wire net4120;
 wire net4121;
 wire net4122;
 wire net4123;
 wire net4124;
 wire net4125;
 wire net4126;
 wire net4127;
 wire net4128;
 wire net4129;
 wire net4130;
 wire net4131;
 wire net4132;
 wire net4133;
 wire net4134;
 wire net4135;
 wire net4136;
 wire net4137;
 wire net4138;
 wire net4139;
 wire net4140;
 wire net4141;
 wire net4142;
 wire net4143;
 wire net4144;
 wire net4145;
 wire net4146;
 wire net4147;
 wire net4148;
 wire net4149;
 wire net4150;
 wire net4151;
 wire net4152;
 wire net4153;
 wire net4154;
 wire net4155;
 wire net4156;
 wire net4157;
 wire net4158;
 wire net4159;
 wire net4160;
 wire net4161;
 wire net4162;
 wire net4163;
 wire net4164;
 wire net4165;
 wire net4166;
 wire net4167;
 wire net4168;
 wire net4169;
 wire net4170;
 wire net4171;
 wire net4172;
 wire net4173;
 wire net4174;
 wire net4175;
 wire net4176;
 wire net4177;
 wire net4178;
 wire net4179;
 wire net4180;
 wire net4181;
 wire net4182;
 wire net4183;
 wire net4184;
 wire net4185;
 wire net4186;
 wire net4187;
 wire net4188;
 wire net4189;
 wire net4190;
 wire net4191;
 wire net4192;
 wire net4193;
 wire net4194;
 wire net4195;
 wire net4196;
 wire net4197;
 wire net4198;
 wire net4199;
 wire net4200;
 wire net4201;
 wire net4202;
 wire net4203;
 wire net4204;
 wire net4205;
 wire net4206;
 wire net4207;
 wire net4208;
 wire net4209;
 wire net4210;
 wire net4211;
 wire net4212;
 wire net4213;
 wire net4214;
 wire net4215;
 wire net4216;
 wire net4217;
 wire net4218;
 wire net4219;
 wire net4220;
 wire net4221;
 wire net4222;
 wire net4223;
 wire net4224;
 wire net4225;
 wire net4226;
 wire net4227;
 wire net4228;
 wire net4229;
 wire net4230;
 wire net4231;
 wire net4232;
 wire net4233;
 wire net4234;
 wire net4235;
 wire net4236;
 wire net4237;
 wire net4238;
 wire net4239;
 wire net4240;
 wire net4241;
 wire net4242;
 wire net4243;
 wire net4244;
 wire net4245;
 wire net4246;
 wire net4247;
 wire net4248;
 wire net4249;
 wire net4250;
 wire net4251;
 wire net4252;
 wire net4253;
 wire net4254;
 wire net4255;
 wire net4256;
 wire net4257;
 wire net4258;
 wire net4259;
 wire net4260;
 wire net4261;
 wire net4262;
 wire net4263;
 wire net4264;
 wire net4265;
 wire net4266;
 wire net4267;
 wire net4268;
 wire net4269;
 wire net4270;
 wire net4271;
 wire net4272;
 wire net4273;
 wire net4274;
 wire net4275;
 wire net4276;
 wire net4277;
 wire net4278;
 wire net4279;
 wire net4280;
 wire net4281;
 wire net4282;
 wire net4283;
 wire net4284;
 wire net4285;
 wire net4286;
 wire net4287;
 wire net4288;
 wire net4289;
 wire net4290;
 wire net4291;
 wire net4292;
 wire net4293;
 wire net4294;
 wire net4295;
 wire net4296;
 wire net4297;
 wire net4298;
 wire net4299;
 wire net4300;
 wire net4301;
 wire net4302;
 wire net4303;
 wire net4304;
 wire net4305;
 wire net4306;
 wire net4307;
 wire net4308;
 wire net4309;
 wire net4310;
 wire net4311;
 wire net4312;
 wire net4313;
 wire net4314;
 wire net4315;
 wire net4316;
 wire net4317;
 wire net4318;
 wire net4319;
 wire net4320;
 wire net4321;
 wire net4322;
 wire net4323;
 wire net4324;
 wire net4325;
 wire net4326;
 wire net4327;
 wire net4328;
 wire net4329;
 wire net4330;
 wire net4331;
 wire net4332;
 wire net4333;
 wire net4334;
 wire net4335;
 wire net4336;
 wire net4337;
 wire net4338;
 wire net4339;
 wire net4340;
 wire net4341;
 wire net4342;
 wire net4343;
 wire net4344;
 wire net4345;
 wire net4346;
 wire net4347;
 wire net4348;
 wire net4349;
 wire net4350;
 wire net4351;
 wire net4352;
 wire net4353;
 wire net4354;
 wire net4355;
 wire net4356;
 wire net4357;
 wire net4358;
 wire net4359;
 wire net4360;
 wire net4361;
 wire net4362;
 wire net4363;
 wire net4364;
 wire net4365;
 wire net4366;
 wire net4367;
 wire net4368;
 wire net4369;
 wire net4370;
 wire net4371;
 wire net4372;
 wire net4373;
 wire net4374;
 wire net4375;
 wire net4376;
 wire net4377;
 wire net4378;
 wire net4379;
 wire net4380;
 wire net4381;
 wire net4382;
 wire net4383;
 wire net4384;
 wire net4385;
 wire net4386;
 wire net4387;
 wire net4388;
 wire net4389;
 wire net4390;
 wire net4391;
 wire net4392;
 wire net4393;
 wire net4394;
 wire net4395;
 wire net4396;
 wire net4397;
 wire net4398;
 wire net4399;
 wire net4400;
 wire net4401;
 wire net4402;
 wire net4403;
 wire net4404;
 wire net4405;
 wire net4406;
 wire net4407;
 wire net4408;
 wire net4409;
 wire net4410;
 wire net4411;
 wire net4412;
 wire net4413;
 wire net4414;
 wire net4415;
 wire net4416;
 wire net4417;
 wire net4418;
 wire net4419;
 wire net4420;
 wire net4421;
 wire net4422;
 wire net4423;
 wire net4424;
 wire net4425;
 wire net4426;
 wire net4427;
 wire net4428;
 wire net4429;
 wire net4430;
 wire net4431;
 wire net4432;
 wire net4433;
 wire net4434;
 wire net4435;
 wire net4436;
 wire net4437;
 wire net4438;
 wire net4439;
 wire net4440;
 wire net4441;
 wire net4442;
 wire net4443;
 wire net4444;
 wire net4445;
 wire net4446;
 wire net4447;
 wire net4448;
 wire net4449;
 wire net4450;
 wire net4451;
 wire net4452;
 wire net4453;
 wire net4454;
 wire net4455;
 wire net4456;
 wire net4457;
 wire net4458;
 wire net4459;
 wire net4460;
 wire net4461;
 wire net4462;
 wire net4463;
 wire net4464;
 wire net4465;
 wire net4466;
 wire net4467;
 wire net4468;
 wire net4469;
 wire net4470;
 wire net4471;
 wire net4472;
 wire net4473;
 wire net4474;
 wire net4475;
 wire net4476;
 wire net4477;
 wire net4478;
 wire net4479;
 wire net4480;
 wire net4481;
 wire net4482;
 wire net4483;
 wire net4484;
 wire net4485;
 wire net4486;
 wire net4487;
 wire net4488;
 wire net4489;
 wire net4490;
 wire net4491;
 wire net4492;
 wire net4493;
 wire net4494;
 wire net4495;
 wire net4496;
 wire net4497;
 wire net4498;
 wire net4499;
 wire net4500;
 wire net4501;
 wire net4502;
 wire net4503;
 wire net4504;
 wire net4505;
 wire net4506;
 wire net4507;
 wire net4508;
 wire net4509;
 wire net4510;
 wire net4511;
 wire net4512;
 wire net4513;
 wire net4514;
 wire net4515;
 wire net4516;
 wire net4517;
 wire net4518;
 wire net4519;
 wire net4520;
 wire net4521;
 wire net4522;
 wire net4523;
 wire net4524;
 wire net4525;
 wire net4526;
 wire net4527;
 wire net4528;
 wire net4529;
 wire net4530;
 wire net4531;
 wire net4532;
 wire net4533;
 wire net4534;
 wire net4535;
 wire net4536;
 wire net4537;
 wire net4538;
 wire net4539;
 wire net4540;
 wire net4541;
 wire net4542;
 wire net4543;
 wire net4544;
 wire net4545;
 wire net4546;
 wire net4547;
 wire net4548;
 wire net4549;
 wire net4550;
 wire net4551;
 wire net4552;
 wire net4553;
 wire net4554;
 wire net4555;
 wire net4556;
 wire net4557;
 wire net4558;
 wire net4559;
 wire net4560;
 wire net4561;
 wire net4562;
 wire net4563;
 wire net4564;
 wire net4565;
 wire net4566;
 wire net4567;
 wire net4568;
 wire net4569;
 wire net4570;
 wire net4571;
 wire net4572;
 wire net4573;
 wire net4574;
 wire net4575;
 wire net4576;
 wire net4577;
 wire net4578;
 wire net4579;
 wire net4580;
 wire net4581;
 wire net4582;
 wire net4583;
 wire net4584;
 wire net4585;
 wire net4586;
 wire net4587;
 wire net4588;
 wire net4589;
 wire net4590;
 wire net4591;
 wire net4592;
 wire net4593;
 wire net4594;
 wire net4595;
 wire net4596;
 wire net4597;
 wire net4598;
 wire net4599;
 wire net4600;
 wire net4601;
 wire net4602;
 wire net4603;
 wire net4604;
 wire net4605;
 wire net4606;
 wire net4607;
 wire net4608;
 wire net4609;
 wire net4610;
 wire net4611;
 wire net4612;
 wire net4613;
 wire net4614;
 wire net4615;
 wire net4616;
 wire net4617;
 wire net4618;
 wire net4619;
 wire net4620;
 wire net4621;
 wire net4622;
 wire net4623;
 wire net4624;
 wire net4625;
 wire net4626;
 wire net4627;
 wire net4628;
 wire net4629;
 wire net4630;
 wire net4631;
 wire net4632;
 wire net4633;
 wire net4634;
 wire net4635;
 wire net4636;
 wire net4637;
 wire net4638;
 wire net4639;
 wire net4640;
 wire net4641;
 wire net4642;
 wire net4643;
 wire net4644;
 wire net4645;
 wire net4646;
 wire net4647;
 wire net4648;
 wire net4649;
 wire net4650;
 wire net4651;
 wire net4652;
 wire net4653;
 wire net4654;
 wire net4655;
 wire net4656;
 wire net4657;
 wire net4658;
 wire net4659;
 wire net4660;
 wire net4661;
 wire net4662;
 wire net4663;
 wire net4664;
 wire net4665;
 wire net4666;
 wire net4667;
 wire net4668;
 wire net4669;
 wire net4670;
 wire net4671;
 wire net4672;
 wire net4673;
 wire net4674;
 wire net4675;
 wire net4676;
 wire net4677;
 wire net4678;
 wire net4679;
 wire net4680;
 wire net4681;
 wire net4682;
 wire net4683;
 wire net4684;
 wire net4685;
 wire net4686;
 wire net4687;
 wire net4688;
 wire net4689;
 wire net4690;
 wire net4691;
 wire net4692;
 wire net4693;
 wire net4694;
 wire net4695;
 wire net4696;
 wire net4697;
 wire net4698;
 wire net4699;
 wire net4700;
 wire net4701;
 wire net4702;
 wire net4703;
 wire net4704;
 wire net4705;
 wire net4706;
 wire net4707;
 wire net4708;
 wire net4709;
 wire net4710;
 wire net4711;
 wire net4712;
 wire net4713;
 wire net4714;
 wire net4715;
 wire net4716;
 wire net4717;
 wire net4718;
 wire net4719;
 wire net4720;
 wire net4721;
 wire net4722;
 wire net4723;
 wire net4724;
 wire net4725;
 wire net4726;
 wire net4727;
 wire net4728;
 wire net4729;
 wire net4730;
 wire net4731;
 wire net4732;
 wire net4733;
 wire net4734;
 wire net4735;
 wire net4736;
 wire net4737;
 wire net4738;
 wire net4739;
 wire net4740;
 wire net4741;
 wire net4742;
 wire net4743;
 wire net4744;
 wire net4745;
 wire net4746;
 wire net4747;
 wire net4748;
 wire net4749;
 wire net4750;
 wire net4751;
 wire net4752;
 wire net4753;
 wire net4754;
 wire net4755;
 wire net4756;
 wire net4757;
 wire net4758;
 wire net4759;
 wire net4760;
 wire net4761;
 wire net4762;
 wire net4763;
 wire net4764;
 wire net4765;
 wire net4766;
 wire net4767;
 wire net4768;
 wire net4769;
 wire net4770;
 wire net4771;
 wire net4772;
 wire net4773;
 wire net4774;
 wire net4775;
 wire net4776;
 wire net4777;
 wire net4778;
 wire net4779;
 wire net4780;
 wire net4781;
 wire net4782;
 wire net4783;
 wire net4784;
 wire net4785;
 wire net4786;
 wire net4787;
 wire net4788;
 wire net4789;
 wire net4790;
 wire net4791;
 wire net4792;
 wire net4793;
 wire net4794;
 wire net4795;
 wire net4796;
 wire net4797;
 wire net4798;
 wire net4799;
 wire net4800;
 wire net4801;
 wire net4802;
 wire net4803;
 wire net4804;
 wire net4805;
 wire net4806;
 wire net4807;
 wire net4808;
 wire net4809;
 wire net4810;
 wire net4811;
 wire net4812;
 wire net4813;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_72_clk;
 wire clknet_leaf_73_clk;
 wire clknet_leaf_74_clk;
 wire clknet_leaf_75_clk;
 wire clknet_0_clk;
 wire clknet_2_0_0_clk;
 wire clknet_2_1_0_clk;
 wire clknet_2_2_0_clk;
 wire clknet_2_3_0_clk;
 wire clknet_4_0__leaf_clk;
 wire clknet_4_1__leaf_clk;
 wire clknet_4_2__leaf_clk;
 wire clknet_4_3__leaf_clk;
 wire clknet_4_4__leaf_clk;
 wire clknet_4_5__leaf_clk;
 wire clknet_4_6__leaf_clk;
 wire clknet_4_7__leaf_clk;
 wire clknet_4_8__leaf_clk;
 wire clknet_4_9__leaf_clk;
 wire clknet_4_10__leaf_clk;
 wire clknet_4_11__leaf_clk;
 wire clknet_4_12__leaf_clk;
 wire clknet_4_13__leaf_clk;
 wire clknet_4_14__leaf_clk;
 wire clknet_4_15__leaf_clk;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;

 sg13g2_inv_1 _10371_ (.Y(_03389_),
    .A(net452));
 sg13g2_inv_1 _10372_ (.Y(_03390_),
    .A(\spiking_network_top_uut.all_data_out[31] ));
 sg13g2_inv_1 _10373_ (.Y(_03391_),
    .A(net474));
 sg13g2_inv_1 _10374_ (.Y(_03392_),
    .A(\spiking_network_top_uut.all_data_out[29] ));
 sg13g2_inv_1 _10375_ (.Y(_03393_),
    .A(\spiking_network_top_uut.clk_div_inst.counter[4] ));
 sg13g2_inv_1 _10376_ (.Y(_03394_),
    .A(\spiking_network_top_uut.all_data_out[28] ));
 sg13g2_inv_1 _10377_ (.Y(_03395_),
    .A(\spiking_network_top_uut.clk_div_inst.counter[3] ));
 sg13g2_inv_1 _10378_ (.Y(_03396_),
    .A(\spiking_network_top_uut.clk_div_inst.counter[2] ));
 sg13g2_inv_1 _10379_ (.Y(_03397_),
    .A(\spiking_network_top_uut.clk_div_inst.counter[1] ));
 sg13g2_inv_1 _10380_ (.Y(_03398_),
    .A(\spiking_network_top_uut.clk_div_inst.counter[0] ));
 sg13g2_inv_1 _10381_ (.Y(_03399_),
    .A(net552));
 sg13g2_inv_1 _10382_ (.Y(_03400_),
    .A(net541));
 sg13g2_inv_2 _10383_ (.Y(_03401_),
    .A(net4310));
 sg13g2_inv_8 _10384_ (.Y(_03402_),
    .A(net4640));
 sg13g2_inv_1 _10385_ (.Y(_03403_),
    .A(net455));
 sg13g2_inv_1 _10386_ (.Y(_03404_),
    .A(net494));
 sg13g2_inv_2 _10387_ (.Y(_03405_),
    .A(\spiking_network_top_uut.spi_inst.LSB_Address_reg[2] ));
 sg13g2_inv_1 _10388_ (.Y(_03406_),
    .A(net4317));
 sg13g2_inv_1 _10389_ (.Y(_03407_),
    .A(net464));
 sg13g2_inv_1 _10390_ (.Y(_03408_),
    .A(net547));
 sg13g2_inv_1 _10391_ (.Y(_03409_),
    .A(net544));
 sg13g2_inv_1 _10392_ (.Y(_03410_),
    .A(net492));
 sg13g2_inv_1 _10393_ (.Y(_03411_),
    .A(net526));
 sg13g2_inv_1 _10394_ (.Y(_03412_),
    .A(net4574));
 sg13g2_inv_1 _10395_ (.Y(_03413_),
    .A(net489));
 sg13g2_inv_1 _10396_ (.Y(_03414_),
    .A(net509));
 sg13g2_inv_1 _10397_ (.Y(_03415_),
    .A(net453));
 sg13g2_inv_1 _10398_ (.Y(_03416_),
    .A(net472));
 sg13g2_inv_1 _10399_ (.Y(_03417_),
    .A(net418));
 sg13g2_inv_8 _10400_ (.Y(_03418_),
    .A(net4529));
 sg13g2_inv_1 _10401_ (.Y(_03419_),
    .A(net454));
 sg13g2_inv_1 _10402_ (.Y(_03420_),
    .A(net497));
 sg13g2_inv_1 _10403_ (.Y(_03421_),
    .A(net534));
 sg13g2_inv_1 _10404_ (.Y(_03422_),
    .A(net530));
 sg13g2_inv_1 _10405_ (.Y(_03423_),
    .A(net532));
 sg13g2_inv_1 _10406_ (.Y(_03424_),
    .A(net538));
 sg13g2_inv_1 _10407_ (.Y(_03425_),
    .A(net507));
 sg13g2_inv_1 _10408_ (.Y(_03426_),
    .A(net521));
 sg13g2_inv_1 _10409_ (.Y(_03427_),
    .A(net451));
 sg13g2_inv_1 _10410_ (.Y(_03428_),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ));
 sg13g2_inv_1 _10411_ (.Y(_03429_),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ));
 sg13g2_inv_1 _10412_ (.Y(_03430_),
    .A(net539));
 sg13g2_inv_1 _10413_ (.Y(_03431_),
    .A(net545));
 sg13g2_inv_1 _10414_ (.Y(_03432_),
    .A(net506));
 sg13g2_inv_1 _10415_ (.Y(_03433_),
    .A(net528));
 sg13g2_inv_1 _10416_ (.Y(_03434_),
    .A(net463));
 sg13g2_inv_1 _10417_ (.Y(_03435_),
    .A(net460));
 sg13g2_inv_1 _10418_ (.Y(_03436_),
    .A(net485));
 sg13g2_inv_1 _10419_ (.Y(_03437_),
    .A(net488));
 sg13g2_inv_1 _10420_ (.Y(_03438_),
    .A(net523));
 sg13g2_inv_1 _10421_ (.Y(_03439_),
    .A(net512));
 sg13g2_inv_1 _10422_ (.Y(_03440_),
    .A(net499));
 sg13g2_inv_1 _10423_ (.Y(_03441_),
    .A(net490));
 sg13g2_inv_1 _10424_ (.Y(_03442_),
    .A(net482));
 sg13g2_inv_1 _10425_ (.Y(_03443_),
    .A(net450));
 sg13g2_inv_1 _10426_ (.Y(_03444_),
    .A(net457));
 sg13g2_inv_1 _10427_ (.Y(_03445_),
    .A(net493));
 sg13g2_inv_1 _10428_ (.Y(_03446_),
    .A(net513));
 sg13g2_inv_1 _10429_ (.Y(_03447_),
    .A(net514));
 sg13g2_inv_1 _10430_ (.Y(_03448_),
    .A(net542));
 sg13g2_inv_1 _10431_ (.Y(_03449_),
    .A(net505));
 sg13g2_inv_1 _10432_ (.Y(_03450_),
    .A(net510));
 sg13g2_inv_1 _10433_ (.Y(_03451_),
    .A(net473));
 sg13g2_inv_1 _10434_ (.Y(_03452_),
    .A(net487));
 sg13g2_inv_1 _10435_ (.Y(_03453_),
    .A(net445));
 sg13g2_inv_1 _10436_ (.Y(_03454_),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ));
 sg13g2_inv_1 _10437_ (.Y(_03455_),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ));
 sg13g2_inv_1 _10438_ (.Y(_03456_),
    .A(net535));
 sg13g2_inv_1 _10439_ (.Y(_03457_),
    .A(net546));
 sg13g2_inv_1 _10440_ (.Y(_03458_),
    .A(net500));
 sg13g2_inv_1 _10441_ (.Y(_03459_),
    .A(net529));
 sg13g2_inv_1 _10442_ (.Y(_03460_),
    .A(net511));
 sg13g2_inv_1 _10443_ (.Y(_03461_),
    .A(net516));
 sg13g2_inv_1 _10444_ (.Y(_03462_),
    .A(net471));
 sg13g2_inv_1 _10445_ (.Y(_03463_),
    .A(net508));
 sg13g2_inv_1 _10446_ (.Y(_03464_),
    .A(net504));
 sg13g2_inv_1 _10447_ (.Y(_03465_),
    .A(net467));
 sg13g2_inv_1 _10448_ (.Y(_03466_),
    .A(net477));
 sg13g2_inv_1 _10449_ (.Y(_03467_),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ));
 sg13g2_inv_1 _10450_ (.Y(_03468_),
    .A(net484));
 sg13g2_inv_1 _10451_ (.Y(_03469_),
    .A(\spiking_network_top_uut.spi_inst.spi_control_unit_inst.current_state[1] ));
 sg13g2_inv_4 _10452_ (.A(net10),
    .Y(_03470_));
 sg13g2_inv_1 _10453_ (.Y(_03471_),
    .A(\spiking_network_top_uut.spi_inst.spi_slave_inst.bit_cnt[0] ));
 sg13g2_inv_1 _10454_ (.Y(_03472_),
    .A(\spiking_network_top_uut.spi_inst.SPI_instruction_reg[3] ));
 sg13g2_inv_1 _10455_ (.Y(_03473_),
    .A(\spiking_network_top_uut.all_data_out[2] ));
 sg13g2_inv_1 _10456_ (.Y(_03474_),
    .A(_00035_));
 sg13g2_inv_1 _10457_ (.Y(_03475_),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.spike_out ));
 sg13g2_inv_1 _10458_ (.Y(_03476_),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.spike_out ));
 sg13g2_inv_4 _10459_ (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.spike_out ),
    .Y(_03477_));
 sg13g2_inv_1 _10460_ (.Y(_03478_),
    .A(_00041_));
 sg13g2_inv_1 _10461_ (.Y(_03479_),
    .A(_00045_));
 sg13g2_inv_1 _10462_ (.Y(_03480_),
    .A(_00046_));
 sg13g2_inv_1 _10463_ (.Y(_03481_),
    .A(_00053_));
 sg13g2_inv_1 _10464_ (.Y(_03482_),
    .A(_00059_));
 sg13g2_inv_1 _10465_ (.Y(_03483_),
    .A(_00071_));
 sg13g2_inv_1 _10466_ (.Y(_03484_),
    .A(_00075_));
 sg13g2_inv_1 _10467_ (.Y(_03485_),
    .A(_00076_));
 sg13g2_inv_1 _10468_ (.Y(_03486_),
    .A(_00080_));
 sg13g2_inv_1 _10469_ (.Y(_03487_),
    .A(_00081_));
 sg13g2_inv_1 _10470_ (.Y(_03488_),
    .A(_00082_));
 sg13g2_inv_1 _10471_ (.Y(_03489_),
    .A(_00087_));
 sg13g2_inv_1 _10472_ (.Y(_03490_),
    .A(_00088_));
 sg13g2_inv_1 _10473_ (.Y(_03491_),
    .A(_00092_));
 sg13g2_inv_1 _10474_ (.Y(_03492_),
    .A(_00093_));
 sg13g2_inv_1 _10475_ (.Y(_03493_),
    .A(_00094_));
 sg13g2_inv_1 _10476_ (.Y(_03494_),
    .A(_00098_));
 sg13g2_inv_1 _10477_ (.Y(_03495_),
    .A(_00099_));
 sg13g2_inv_1 _10478_ (.Y(_03496_),
    .A(_00104_));
 sg13g2_inv_1 _10479_ (.Y(_03497_),
    .A(_00105_));
 sg13g2_inv_1 _10480_ (.Y(_03498_),
    .A(_00106_));
 sg13g2_inv_1 _10481_ (.Y(_03499_),
    .A(_00111_));
 sg13g2_inv_1 _10482_ (.Y(_03500_),
    .A(_00117_));
 sg13g2_inv_1 _10483_ (.Y(_03501_),
    .A(_00118_));
 sg13g2_inv_1 _10484_ (.Y(_03502_),
    .A(_00123_));
 sg13g2_inv_1 _10485_ (.Y(_03503_),
    .A(_00124_));
 sg13g2_inv_1 _10486_ (.Y(_03504_),
    .A(_00128_));
 sg13g2_inv_1 _10487_ (.Y(_03505_),
    .A(_00129_));
 sg13g2_inv_1 _10488_ (.Y(_03506_),
    .A(_00135_));
 sg13g2_inv_1 _10489_ (.Y(_03507_),
    .A(_00136_));
 sg13g2_inv_1 _10490_ (.Y(_03508_),
    .A(\spiking_network_top_uut.spi_inst.memory_inst.addr_reg_out[3] ));
 sg13g2_inv_4 _10491_ (.A(_00144_),
    .Y(_03509_));
 sg13g2_inv_1 _10492_ (.Y(_03510_),
    .A(_00150_));
 sg13g2_inv_1 _10493_ (.Y(_03511_),
    .A(\spiking_network_top_uut.all_data_out[814] ));
 sg13g2_inv_1 _10494_ (.Y(_03512_),
    .A(_00154_));
 sg13g2_inv_1 _10495_ (.Y(_03513_),
    .A(\spiking_network_top_uut.all_data_out[774] ));
 sg13g2_inv_1 _10496_ (.Y(_03514_),
    .A(_00156_));
 sg13g2_inv_1 _10497_ (.Y(_03515_),
    .A(\spiking_network_top_uut.all_data_out[766] ));
 sg13g2_inv_1 _10498_ (.Y(_03516_),
    .A(_00157_));
 sg13g2_inv_1 _10499_ (.Y(_03517_),
    .A(_00158_));
 sg13g2_inv_4 _10500_ (.A(_00159_),
    .Y(_03518_));
 sg13g2_inv_1 _10501_ (.Y(_03519_),
    .A(_00160_));
 sg13g2_inv_1 _10502_ (.Y(_03520_),
    .A(\spiking_network_top_uut.all_data_out[734] ));
 sg13g2_inv_2 _10503_ (.Y(_03521_),
    .A(_00161_));
 sg13g2_inv_2 _10504_ (.Y(_03522_),
    .A(_00162_));
 sg13g2_inv_1 _10505_ (.Y(_03523_),
    .A(\spiking_network_top_uut.all_data_out[718] ));
 sg13g2_inv_2 _10506_ (.Y(_03524_),
    .A(_00163_));
 sg13g2_inv_2 _10507_ (.Y(_03525_),
    .A(_00166_));
 sg13g2_inv_2 _10508_ (.Y(_03526_),
    .A(_00167_));
 sg13g2_inv_1 _10509_ (.Y(_03527_),
    .A(_00170_));
 sg13g2_inv_1 _10510_ (.Y(_03528_),
    .A(\spiking_network_top_uut.all_data_out[646] ));
 sg13g2_inv_1 _10511_ (.Y(_03529_),
    .A(_00173_));
 sg13g2_inv_1 _10512_ (.Y(_03530_),
    .A(\spiking_network_top_uut.all_data_out[630] ));
 sg13g2_inv_1 _10513_ (.Y(_03531_),
    .A(\spiking_network_top_uut.all_data_out[614] ));
 sg13g2_inv_1 _10514_ (.Y(_03532_),
    .A(_00177_));
 sg13g2_inv_2 _10515_ (.Y(_03533_),
    .A(_00179_));
 sg13g2_inv_4 _10516_ (.A(_00181_),
    .Y(_03534_));
 sg13g2_inv_1 _10517_ (.Y(_03535_),
    .A(_00182_));
 sg13g2_inv_2 _10518_ (.Y(_03536_),
    .A(_00184_));
 sg13g2_inv_2 _10519_ (.Y(_03537_),
    .A(_00190_));
 sg13g2_inv_1 _10520_ (.Y(_03538_),
    .A(\spiking_network_top_uut.all_data_out[486] ));
 sg13g2_inv_1 _10521_ (.Y(_03539_),
    .A(\spiking_network_top_uut.all_data_out[438] ));
 sg13g2_inv_1 _10522_ (.Y(_03540_),
    .A(\spiking_network_top_uut.all_data_out[430] ));
 sg13g2_inv_2 _10523_ (.Y(_03541_),
    .A(_00202_));
 sg13g2_inv_1 _10524_ (.Y(_03542_),
    .A(\spiking_network_top_uut.all_data_out[398] ));
 sg13g2_inv_4 _10525_ (.A(_00204_),
    .Y(_03543_));
 sg13g2_inv_4 _10526_ (.A(_00205_),
    .Y(_03544_));
 sg13g2_inv_1 _10527_ (.Y(_03545_),
    .A(\spiking_network_top_uut.all_data_out[374] ));
 sg13g2_inv_4 _10528_ (.A(_00207_),
    .Y(_03546_));
 sg13g2_inv_1 _10529_ (.Y(_03547_),
    .A(_00210_));
 sg13g2_inv_4 _10530_ (.A(_00215_),
    .Y(_03548_));
 sg13g2_inv_4 _10531_ (.A(_00216_),
    .Y(_03549_));
 sg13g2_inv_4 _10532_ (.A(_00222_),
    .Y(_03550_));
 sg13g2_inv_4 _10533_ (.A(_00225_),
    .Y(_03551_));
 sg13g2_inv_1 _10534_ (.Y(_03552_),
    .A(_00227_));
 sg13g2_inv_2 _10535_ (.Y(_03553_),
    .A(_00228_));
 sg13g2_inv_1 _10536_ (.Y(_03554_),
    .A(_00230_));
 sg13g2_inv_1 _10537_ (.Y(_03555_),
    .A(_00231_));
 sg13g2_inv_1 _10538_ (.Y(_03556_),
    .A(_00232_));
 sg13g2_inv_1 _10539_ (.Y(_03557_),
    .A(_00234_));
 sg13g2_inv_1 _10540_ (.Y(_03558_),
    .A(_00236_));
 sg13g2_inv_1 _10541_ (.Y(_03559_),
    .A(_00237_));
 sg13g2_inv_2 _10542_ (.Y(_03560_),
    .A(_00238_));
 sg13g2_inv_1 _10543_ (.Y(_03561_),
    .A(_00239_));
 sg13g2_inv_1 _10544_ (.Y(_03562_),
    .A(_00246_));
 sg13g2_inv_1 _10545_ (.Y(_03563_),
    .A(_00247_));
 sg13g2_inv_1 _10546_ (.Y(_03564_),
    .A(_00248_));
 sg13g2_inv_2 _10547_ (.Y(_03565_),
    .A(_00252_));
 sg13g2_inv_1 _10548_ (.Y(_03566_),
    .A(_00253_));
 sg13g2_inv_2 _10549_ (.Y(_03567_),
    .A(_00266_));
 sg13g2_inv_2 _10550_ (.Y(_03568_),
    .A(_00267_));
 sg13g2_inv_2 _10551_ (.Y(_03569_),
    .A(_00268_));
 sg13g2_inv_1 _10552_ (.Y(_03570_),
    .A(_00272_));
 sg13g2_inv_4 _10553_ (.A(_00274_),
    .Y(_03571_));
 sg13g2_inv_1 _10554_ (.Y(_03572_),
    .A(_00276_));
 sg13g2_inv_4 _10555_ (.A(_00277_),
    .Y(_03573_));
 sg13g2_inv_4 _10556_ (.A(_00280_),
    .Y(_03574_));
 sg13g2_inv_1 _10557_ (.Y(_03575_),
    .A(\spiking_network_top_uut.all_data_out[4] ));
 sg13g2_inv_2 _10558_ (.Y(_03576_),
    .A(_00281_));
 sg13g2_inv_1 _10559_ (.Y(_03577_),
    .A(\spiking_network_top_uut.all_data_out[882] ));
 sg13g2_inv_4 _10560_ (.A(_00282_),
    .Y(_03578_));
 sg13g2_inv_1 _10561_ (.Y(_03579_),
    .A(_00285_));
 sg13g2_inv_4 _10562_ (.A(_00286_),
    .Y(_03580_));
 sg13g2_inv_1 _10563_ (.Y(_03581_),
    .A(\spiking_network_top_uut.all_data_out[842] ));
 sg13g2_inv_4 _10564_ (.A(_00287_),
    .Y(_03582_));
 sg13g2_inv_1 _10565_ (.Y(_03583_),
    .A(\spiking_network_top_uut.all_data_out[818] ));
 sg13g2_inv_2 _10566_ (.Y(_03584_),
    .A(_00290_));
 sg13g2_inv_1 _10567_ (.Y(_03585_),
    .A(\spiking_network_top_uut.all_data_out[802] ));
 sg13g2_inv_1 _10568_ (.Y(_03586_),
    .A(_00292_));
 sg13g2_inv_2 _10569_ (.Y(_03587_),
    .A(_00294_));
 sg13g2_inv_4 _10570_ (.A(_00295_),
    .Y(_03588_));
 sg13g2_inv_2 _10571_ (.Y(_03589_),
    .A(_00296_));
 sg13g2_inv_2 _10572_ (.Y(_03590_),
    .A(_00297_));
 sg13g2_inv_1 _10573_ (.Y(_03591_),
    .A(_00301_));
 sg13g2_inv_2 _10574_ (.Y(_03592_),
    .A(_00302_));
 sg13g2_inv_1 _10575_ (.Y(_03593_),
    .A(_00304_));
 sg13g2_inv_1 _10576_ (.Y(_03594_),
    .A(_00305_));
 sg13g2_inv_2 _10577_ (.Y(_03595_),
    .A(_00306_));
 sg13g2_inv_1 _10578_ (.Y(_03596_),
    .A(\spiking_network_top_uut.all_data_out[682] ));
 sg13g2_inv_4 _10579_ (.A(_00307_),
    .Y(_03597_));
 sg13g2_inv_2 _10580_ (.Y(_03598_),
    .A(_00308_));
 sg13g2_inv_2 _10581_ (.Y(_03599_),
    .A(_00310_));
 sg13g2_inv_1 _10582_ (.Y(_03600_),
    .A(\spiking_network_top_uut.all_data_out[650] ));
 sg13g2_inv_1 _10583_ (.Y(_03601_),
    .A(_00311_));
 sg13g2_inv_2 _10584_ (.Y(_03602_),
    .A(_00312_));
 sg13g2_inv_1 _10585_ (.Y(_03603_),
    .A(\spiking_network_top_uut.all_data_out[634] ));
 sg13g2_inv_1 _10586_ (.Y(_03604_),
    .A(_00313_));
 sg13g2_inv_2 _10587_ (.Y(_03605_),
    .A(_00316_));
 sg13g2_inv_1 _10588_ (.Y(_03606_),
    .A(_00317_));
 sg13g2_inv_2 _10589_ (.Y(_03607_),
    .A(_00318_));
 sg13g2_inv_1 _10590_ (.Y(_03608_),
    .A(_00320_));
 sg13g2_inv_4 _10591_ (.A(_00321_),
    .Y(_03609_));
 sg13g2_inv_4 _10592_ (.A(_00323_),
    .Y(_03610_));
 sg13g2_inv_4 _10593_ (.A(_00324_),
    .Y(_03611_));
 sg13g2_inv_1 _10594_ (.Y(_03612_),
    .A(\spiking_network_top_uut.all_data_out[538] ));
 sg13g2_inv_4 _10595_ (.A(_00325_),
    .Y(_03613_));
 sg13g2_inv_2 _10596_ (.Y(_03614_),
    .A(_00326_));
 sg13g2_inv_2 _10597_ (.Y(_03615_),
    .A(_00327_));
 sg13g2_inv_2 _10598_ (.Y(_03616_),
    .A(_00330_));
 sg13g2_inv_1 _10599_ (.Y(_03617_),
    .A(\spiking_network_top_uut.all_data_out[490] ));
 sg13g2_inv_4 _10600_ (.A(_00331_),
    .Y(_03618_));
 sg13g2_inv_4 _10601_ (.A(_00332_),
    .Y(_03619_));
 sg13g2_inv_2 _10602_ (.Y(_03620_),
    .A(_00333_));
 sg13g2_inv_1 _10603_ (.Y(_03621_),
    .A(\spiking_network_top_uut.all_data_out[466] ));
 sg13g2_inv_4 _10604_ (.A(_00335_),
    .Y(_03622_));
 sg13g2_inv_1 _10605_ (.Y(_03623_),
    .A(\spiking_network_top_uut.all_data_out[450] ));
 sg13g2_inv_4 _10606_ (.A(_00337_),
    .Y(_03624_));
 sg13g2_inv_4 _10607_ (.A(_00339_),
    .Y(_03625_));
 sg13g2_inv_4 _10608_ (.A(_00341_),
    .Y(_03626_));
 sg13g2_inv_2 _10609_ (.Y(_03627_),
    .A(_00342_));
 sg13g2_inv_4 _10610_ (.A(_00344_),
    .Y(_03628_));
 sg13g2_inv_4 _10611_ (.A(_00345_),
    .Y(_03629_));
 sg13g2_inv_1 _10612_ (.Y(_03630_),
    .A(_00346_));
 sg13g2_inv_4 _10613_ (.A(_00348_),
    .Y(_03631_));
 sg13g2_inv_1 _10614_ (.Y(_03632_),
    .A(_00350_));
 sg13g2_inv_4 _10615_ (.A(_00353_),
    .Y(_03633_));
 sg13g2_inv_2 _10616_ (.Y(_03634_),
    .A(_00360_));
 sg13g2_inv_1 _10617_ (.Y(_03635_),
    .A(_00370_));
 sg13g2_inv_1 _10618_ (.Y(_03636_),
    .A(_00371_));
 sg13g2_inv_1 _10619_ (.Y(_03637_),
    .A(_00372_));
 sg13g2_inv_1 _10620_ (.Y(_03638_),
    .A(_00374_));
 sg13g2_inv_1 _10621_ (.Y(_03639_),
    .A(_00375_));
 sg13g2_inv_4 _10622_ (.A(_00376_),
    .Y(_03640_));
 sg13g2_inv_2 _10623_ (.Y(_03641_),
    .A(_00378_));
 sg13g2_inv_1 _10624_ (.Y(_03642_),
    .A(_00379_));
 sg13g2_inv_1 _10625_ (.Y(_03643_),
    .A(_00380_));
 sg13g2_inv_1 _10626_ (.Y(_03644_),
    .A(_00381_));
 sg13g2_inv_1 _10627_ (.Y(_03645_),
    .A(_00383_));
 sg13g2_inv_1 _10628_ (.Y(_03646_),
    .A(_00387_));
 sg13g2_inv_2 _10629_ (.Y(_03647_),
    .A(_00396_));
 sg13g2_inv_4 _10630_ (.A(_00405_),
    .Y(_03648_));
 sg13g2_inv_4 _10631_ (.A(_00407_),
    .Y(_03649_));
 sg13g2_inv_4 _10632_ (.A(_00414_),
    .Y(_03650_));
 sg13g2_inv_2 _10633_ (.Y(_03651_),
    .A(_00416_));
 sg13g2_inv_4 _10634_ (.A(_00417_),
    .Y(_03652_));
 sg13g2_inv_4 _10635_ (.A(_00418_),
    .Y(_03653_));
 sg13g2_inv_4 _10636_ (.A(_00420_),
    .Y(_03654_));
 sg13g2_inv_1 _10637_ (.Y(_03655_),
    .A(_00140_));
 sg13g2_inv_1 _10638_ (.Y(_03656_),
    .A(net4422));
 sg13g2_inv_1 _10639_ (.Y(_03657_),
    .A(net4402));
 sg13g2_inv_2 _10640_ (.Y(_03658_),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[5] ));
 sg13g2_inv_2 _10641_ (.Y(_03659_),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[5] ));
 sg13g2_inv_2 _10642_ (.Y(_03660_),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[5] ));
 sg13g2_inv_2 _10643_ (.Y(_03661_),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[5] ));
 sg13g2_inv_1 _10644_ (.Y(_03662_),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[5] ));
 sg13g2_inv_2 _10645_ (.Y(_03663_),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[5] ));
 sg13g2_inv_4 _10646_ (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[5] ),
    .Y(_03664_));
 sg13g2_inv_2 _10647_ (.Y(_03665_),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[5] ));
 sg13g2_inv_2 _10648_ (.Y(_03666_),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[5] ));
 sg13g2_inv_2 _10649_ (.Y(_03667_),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[5] ));
 sg13g2_inv_1 _10650_ (.Y(_03668_),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[5] ));
 sg13g2_inv_1 _10651_ (.Y(_03669_),
    .A(net65));
 sg13g2_inv_1 _10652_ (.Y(_03670_),
    .A(net107));
 sg13g2_inv_1 _10653_ (.Y(_03671_),
    .A(net142));
 sg13g2_inv_1 _10654_ (.Y(_03672_),
    .A(net86));
 sg13g2_inv_1 _10655_ (.Y(_03673_),
    .A(net120));
 sg13g2_inv_1 _10656_ (.Y(_03674_),
    .A(net113));
 sg13g2_inv_1 _10657_ (.Y(_03675_),
    .A(net251));
 sg13g2_inv_1 _10658_ (.Y(_03676_),
    .A(net108));
 sg13g2_inv_1 _10659_ (.Y(_03677_),
    .A(net148));
 sg13g2_inv_1 _10660_ (.Y(_03678_),
    .A(net115));
 sg13g2_inv_1 _10661_ (.Y(_03679_),
    .A(net58));
 sg13g2_inv_1 _10662_ (.Y(_03680_),
    .A(net76));
 sg13g2_inv_1 _10663_ (.Y(_03681_),
    .A(net53));
 sg13g2_inv_1 _10664_ (.Y(_03682_),
    .A(net94));
 sg13g2_inv_1 _10665_ (.Y(_03683_),
    .A(net136));
 sg13g2_inv_1 _10666_ (.Y(_03684_),
    .A(net38));
 sg13g2_inv_1 _10667_ (.Y(_03685_),
    .A(net78));
 sg13g2_inv_1 _10668_ (.Y(_03686_),
    .A(net122));
 sg13g2_inv_1 _10669_ (.Y(_03687_),
    .A(net149));
 sg13g2_inv_1 _10670_ (.Y(_03688_),
    .A(net97));
 sg13g2_inv_1 _10671_ (.Y(_03689_),
    .A(net114));
 sg13g2_inv_1 _10672_ (.Y(_03690_),
    .A(net171));
 sg13g2_inv_1 _10673_ (.Y(_03691_),
    .A(net87));
 sg13g2_inv_1 _10674_ (.Y(_03692_),
    .A(net106));
 sg13g2_inv_1 _10675_ (.Y(_03693_),
    .A(net159));
 sg13g2_inv_1 _10676_ (.Y(_00421_),
    .A(net4705));
 sg13g2_and2_2 _10677_ (.A(\spiking_network_top_uut.spi_inst.spi_slave_inst.bit_cnt[0] ),
    .B(\spiking_network_top_uut.spi_inst.spi_slave_inst.bit_cnt[1] ),
    .X(_03694_));
 sg13g2_and3_2 _10678_ (.X(_00026_),
    .A(_03470_),
    .B(\spiking_network_top_uut.spi_inst.spi_slave_inst.bit_cnt[2] ),
    .C(_03694_));
 sg13g2_nand3_1 _10679_ (.B(\spiking_network_top_uut.spi_inst.spi_control_unit_inst.current_state[0] ),
    .C(\spiking_network_top_uut.spi_inst.spi_control_unit_inst.current_state[2] ),
    .A(_03469_),
    .Y(_03695_));
 sg13g2_or4_1 _10680_ (.A(\spiking_network_top_uut.spi_inst.SPI_instruction_reg[5] ),
    .B(\spiking_network_top_uut.spi_inst.SPI_instruction_reg[4] ),
    .C(\spiking_network_top_uut.spi_inst.SPI_instruction_reg[7] ),
    .D(\spiking_network_top_uut.spi_inst.SPI_instruction_reg[6] ),
    .X(_03696_));
 sg13g2_nand2b_1 _10681_ (.Y(_03697_),
    .B(\spiking_network_top_uut.spi_inst.SPI_instruction_reg[0] ),
    .A_N(\spiking_network_top_uut.spi_inst.SPI_instruction_reg[1] ));
 sg13g2_or4_2 _10682_ (.A(\spiking_network_top_uut.spi_inst.SPI_instruction_reg[2] ),
    .B(_03472_),
    .C(_03696_),
    .D(_03697_),
    .X(_03698_));
 sg13g2_inv_1 _10683_ (.Y(_03699_),
    .A(_03698_));
 sg13g2_nor2_2 _10684_ (.A(_03695_),
    .B(_03698_),
    .Y(_02057_));
 sg13g2_nor3_2 _10685_ (.A(\spiking_network_top_uut.spi_inst.SPI_instruction_reg[3] ),
    .B(_03696_),
    .C(_03697_),
    .Y(_03700_));
 sg13g2_nand2_2 _10686_ (.Y(_03701_),
    .A(\spiking_network_top_uut.spi_inst.SPI_instruction_reg[2] ),
    .B(_03700_));
 sg13g2_nor2_2 _10687_ (.A(_03695_),
    .B(_03701_),
    .Y(_02058_));
 sg13g2_nor2_2 _10688_ (.A(\spiking_network_top_uut.spi_inst.memory_inst.addr_reg_out[5] ),
    .B(\spiking_network_top_uut.spi_inst.memory_inst.addr_reg_out[4] ),
    .Y(_03702_));
 sg13g2_nand2b_1 _10689_ (.Y(_03703_),
    .B(_03702_),
    .A_N(\spiking_network_top_uut.spi_inst.memory_inst.addr_reg_out[6] ));
 sg13g2_nor2_2 _10690_ (.A(\spiking_network_top_uut.spi_inst.memory_inst.addr_reg_out[2] ),
    .B(\spiking_network_top_uut.spi_inst.memory_inst.addr_reg_out[3] ),
    .Y(_03704_));
 sg13g2_nand3_1 _10691_ (.B(net4262),
    .C(_03704_),
    .A(net4265),
    .Y(_03705_));
 sg13g2_nor2_2 _10692_ (.A(net3782),
    .B(_03705_),
    .Y(_03706_));
 sg13g2_nor2b_2 _10693_ (.A(\spiking_network_top_uut.spi_inst.memory_inst.addr_reg_out[3] ),
    .B_N(\spiking_network_top_uut.spi_inst.memory_inst.addr_reg_out[2] ),
    .Y(_03707_));
 sg13g2_nand3_1 _10694_ (.B(net4262),
    .C(_03707_),
    .A(net4264),
    .Y(_03708_));
 sg13g2_nor2_1 _10695_ (.A(net3781),
    .B(net3779),
    .Y(_03709_));
 sg13g2_nand3_1 _10696_ (.B(\spiking_network_top_uut.spi_inst.memory_inst.addr_reg_out[2] ),
    .C(\spiking_network_top_uut.spi_inst.memory_inst.addr_reg_out[3] ),
    .A(net4264),
    .Y(_03710_));
 sg13g2_nor2_2 _10697_ (.A(net4263),
    .B(_03710_),
    .Y(_03711_));
 sg13g2_or2_2 _10698_ (.X(_03712_),
    .B(_03710_),
    .A(net4262));
 sg13g2_nor2_2 _10699_ (.A(net3781),
    .B(_03712_),
    .Y(_03713_));
 sg13g2_nand3b_1 _10700_ (.B(_03707_),
    .C(net4264),
    .Y(_03714_),
    .A_N(net4262));
 sg13g2_nor2_1 _10701_ (.A(net3782),
    .B(net3778),
    .Y(_03715_));
 sg13g2_nand2_2 _10702_ (.Y(_03716_),
    .A(\spiking_network_top_uut.spi_inst.memory_inst.addr_reg_out[5] ),
    .B(\spiking_network_top_uut.spi_inst.memory_inst.addr_reg_out[4] ));
 sg13g2_inv_1 _10703_ (.Y(_03717_),
    .A(_03716_));
 sg13g2_nor2_2 _10704_ (.A(\spiking_network_top_uut.spi_inst.memory_inst.addr_reg_out[6] ),
    .B(_03716_),
    .Y(_03718_));
 sg13g2_or2_1 _10705_ (.X(_03719_),
    .B(_03716_),
    .A(\spiking_network_top_uut.spi_inst.memory_inst.addr_reg_out[6] ));
 sg13g2_nor2_2 _10706_ (.A(net4264),
    .B(net4262),
    .Y(_03720_));
 sg13g2_and2_2 _10707_ (.A(_03704_),
    .B(_03720_),
    .X(_03721_));
 sg13g2_nand2_2 _10708_ (.Y(_03722_),
    .A(_03704_),
    .B(_03720_));
 sg13g2_nor2_2 _10709_ (.A(net3775),
    .B(_03722_),
    .Y(_03723_));
 sg13g2_nand3_1 _10710_ (.B(\spiking_network_top_uut.spi_inst.memory_inst.addr_reg_out[3] ),
    .C(_03720_),
    .A(\spiking_network_top_uut.spi_inst.memory_inst.addr_reg_out[2] ),
    .Y(_03724_));
 sg13g2_nor2_1 _10711_ (.A(net3782),
    .B(_03724_),
    .Y(_03725_));
 sg13g2_nor2b_2 _10712_ (.A(net4264),
    .B_N(net4263),
    .Y(_03726_));
 sg13g2_nand3_1 _10713_ (.B(\spiking_network_top_uut.spi_inst.memory_inst.addr_reg_out[3] ),
    .C(_03726_),
    .A(\spiking_network_top_uut.spi_inst.memory_inst.addr_reg_out[2] ),
    .Y(_03727_));
 sg13g2_nor2_1 _10714_ (.A(net3781),
    .B(net3774),
    .Y(_03728_));
 sg13g2_nand4_1 _10715_ (.B(net4262),
    .C(\spiking_network_top_uut.spi_inst.memory_inst.addr_reg_out[2] ),
    .A(net4264),
    .Y(_03729_),
    .D(\spiking_network_top_uut.spi_inst.memory_inst.addr_reg_out[3] ));
 sg13g2_nor2_1 _10716_ (.A(net3781),
    .B(net3919),
    .Y(_03730_));
 sg13g2_nand2_1 _10717_ (.Y(_03731_),
    .A(_03707_),
    .B(_03720_));
 sg13g2_nor2_1 _10718_ (.A(net3782),
    .B(net3773),
    .Y(_03732_));
 sg13g2_nand3b_1 _10719_ (.B(_03704_),
    .C(net4264),
    .Y(_03733_),
    .A_N(net4262));
 sg13g2_nor2_2 _10720_ (.A(\spiking_network_top_uut.spi_inst.memory_inst.addr_reg_out[2] ),
    .B(_03508_),
    .Y(_03734_));
 sg13g2_nand2_2 _10721_ (.Y(_03735_),
    .A(_03726_),
    .B(_03734_));
 sg13g2_nand2_2 _10722_ (.Y(_03736_),
    .A(_03707_),
    .B(_03726_));
 sg13g2_nor2_1 _10723_ (.A(net3781),
    .B(_03736_),
    .Y(_03737_));
 sg13g2_and2_2 _10724_ (.A(_03720_),
    .B(_03734_),
    .X(_03738_));
 sg13g2_nand2_2 _10725_ (.Y(_03739_),
    .A(_03720_),
    .B(_03734_));
 sg13g2_nor2_1 _10726_ (.A(net3781),
    .B(_03739_),
    .Y(_03740_));
 sg13g2_nand2_1 _10727_ (.Y(_03741_),
    .A(_03704_),
    .B(_03726_));
 sg13g2_nor2_2 _10728_ (.A(net3782),
    .B(net3771),
    .Y(_03742_));
 sg13g2_a21oi_2 _10729_ (.B1(\spiking_network_top_uut.spi_inst.memory_inst.addr_reg_out[6] ),
    .Y(_03743_),
    .A2(net3772),
    .A1(_03702_));
 sg13g2_nor3_2 _10730_ (.A(_00139_),
    .B(_03716_),
    .C(_03722_),
    .Y(_03744_));
 sg13g2_a21oi_2 _10731_ (.B1(_00139_),
    .Y(_03745_),
    .A2(_03722_),
    .A1(_03717_));
 sg13g2_nand3_1 _10732_ (.B(net4263),
    .C(_03734_),
    .A(net4265),
    .Y(_03746_));
 sg13g2_nor2_2 _10733_ (.A(net3781),
    .B(net3708),
    .Y(_03747_));
 sg13g2_nor2_2 _10734_ (.A(net3781),
    .B(_03735_),
    .Y(_03748_));
 sg13g2_nand3b_1 _10735_ (.B(_03734_),
    .C(net4264),
    .Y(_03749_),
    .A_N(net4262));
 sg13g2_nor2_1 _10736_ (.A(net3782),
    .B(net3707),
    .Y(_03750_));
 sg13g2_or4_1 _10737_ (.A(net3717),
    .B(_03728_),
    .C(net3710),
    .D(net3695),
    .X(_03751_));
 sg13g2_nor3_1 _10738_ (.A(net3715),
    .B(_03725_),
    .C(net3709),
    .Y(_03752_));
 sg13g2_nor4_1 _10739_ (.A(net3716),
    .B(_03730_),
    .C(net3711),
    .D(_03750_),
    .Y(_03753_));
 sg13g2_nor4_1 _10740_ (.A(net3719),
    .B(_03709_),
    .C(net3696),
    .D(net3694),
    .Y(_03754_));
 sg13g2_nand3_1 _10741_ (.B(_03753_),
    .C(_03754_),
    .A(_03752_),
    .Y(_03755_));
 sg13g2_nor4_2 _10742_ (.A(_03743_),
    .B(_03745_),
    .C(_03751_),
    .Y(_03756_),
    .D(_03755_));
 sg13g2_or4_2 _10743_ (.A(_03743_),
    .B(_03745_),
    .C(_03751_),
    .D(_03755_),
    .X(_03757_));
 sg13g2_nor3_2 _10744_ (.A(\spiking_network_top_uut.spi_inst.memory_inst.addr_reg_out[5] ),
    .B(\spiking_network_top_uut.spi_inst.memory_inst.addr_reg_out[4] ),
    .C(_00139_),
    .Y(_03758_));
 sg13g2_nand2b_1 _10745_ (.Y(_03759_),
    .B(_03702_),
    .A_N(_00139_));
 sg13g2_nor2_2 _10746_ (.A(net3708),
    .B(net3770),
    .Y(_03760_));
 sg13g2_nor2b_2 _10747_ (.A(\spiking_network_top_uut.spi_inst.memory_inst.addr_reg_out[5] ),
    .B_N(\spiking_network_top_uut.spi_inst.memory_inst.addr_reg_out[4] ),
    .Y(_03761_));
 sg13g2_nand2b_1 _10748_ (.Y(_03762_),
    .B(_03761_),
    .A_N(\spiking_network_top_uut.spi_inst.memory_inst.addr_reg_out[6] ));
 sg13g2_nor2_2 _10749_ (.A(_03708_),
    .B(net3767),
    .Y(_03763_));
 sg13g2_nor2_2 _10750_ (.A(net3778),
    .B(net3768),
    .Y(_03764_));
 sg13g2_nor2b_2 _10751_ (.A(_00139_),
    .B_N(_03761_),
    .Y(_03765_));
 sg13g2_nand2b_2 _10752_ (.Y(_03766_),
    .B(_03761_),
    .A_N(_00139_));
 sg13g2_nor2_2 _10753_ (.A(net3772),
    .B(net3765),
    .Y(_03767_));
 sg13g2_nand2b_1 _10754_ (.Y(_03768_),
    .B(_03765_),
    .A_N(net3772));
 sg13g2_nor2_2 _10755_ (.A(net3780),
    .B(net3763),
    .Y(_03769_));
 sg13g2_nor2b_1 _10756_ (.A(\spiking_network_top_uut.spi_inst.memory_inst.addr_reg_out[4] ),
    .B_N(\spiking_network_top_uut.spi_inst.memory_inst.addr_reg_out[5] ),
    .Y(_03770_));
 sg13g2_nand2b_1 _10757_ (.Y(_03771_),
    .B(_03770_),
    .A_N(\spiking_network_top_uut.spi_inst.memory_inst.addr_reg_out[6] ));
 sg13g2_nor2_2 _10758_ (.A(_03729_),
    .B(net3760),
    .Y(_03772_));
 sg13g2_nor2b_2 _10759_ (.A(_00139_),
    .B_N(_03770_),
    .Y(_03773_));
 sg13g2_nand2b_1 _10760_ (.Y(_03774_),
    .B(_03770_),
    .A_N(_00139_));
 sg13g2_nor2_2 _10761_ (.A(net3708),
    .B(net3757),
    .Y(_03775_));
 sg13g2_nor2_2 _10762_ (.A(net3778),
    .B(net3766),
    .Y(_03776_));
 sg13g2_nor2_2 _10763_ (.A(net3780),
    .B(net3775),
    .Y(_03777_));
 sg13g2_nand2b_2 _10764_ (.Y(_03778_),
    .B(_03718_),
    .A_N(net3780));
 sg13g2_nor2_2 _10765_ (.A(net3782),
    .B(net3772),
    .Y(_03779_));
 sg13g2_nor2_2 _10766_ (.A(net3708),
    .B(_03762_),
    .Y(_03780_));
 sg13g2_nor2_2 _10767_ (.A(net3919),
    .B(net3770),
    .Y(_03781_));
 sg13g2_nor2_2 _10768_ (.A(net3772),
    .B(net3767),
    .Y(_03782_));
 sg13g2_nor2_2 _10769_ (.A(net3775),
    .B(_03749_),
    .Y(_03783_));
 sg13g2_nor2_2 _10770_ (.A(net3707),
    .B(net3768),
    .Y(_03784_));
 sg13g2_nor2_2 _10771_ (.A(net3919),
    .B(net3766),
    .Y(_03785_));
 sg13g2_nor2_2 _10772_ (.A(_03712_),
    .B(net3775),
    .Y(_03786_));
 sg13g2_nand2_2 _10773_ (.Y(_03787_),
    .A(_03711_),
    .B(_03718_));
 sg13g2_nor2_2 _10774_ (.A(net3780),
    .B(net3766),
    .Y(_03788_));
 sg13g2_nor2_2 _10775_ (.A(_03712_),
    .B(net3757),
    .Y(_03789_));
 sg13g2_nor2_2 _10776_ (.A(net3919),
    .B(net3757),
    .Y(_03790_));
 sg13g2_nand2b_2 _10777_ (.Y(_03791_),
    .B(_03773_),
    .A_N(net3919));
 sg13g2_nor2_2 _10778_ (.A(_03712_),
    .B(net3766),
    .Y(_03792_));
 sg13g2_a22oi_1 _10779_ (.Y(_03793_),
    .B1(_03792_),
    .B2(\spiking_network_top_uut.all_data_out[232] ),
    .A2(_03790_),
    .A1(\spiking_network_top_uut.all_data_out[888] ));
 sg13g2_nor2_2 _10780_ (.A(net3780),
    .B(net3768),
    .Y(_03794_));
 sg13g2_nor2_2 _10781_ (.A(net3772),
    .B(net3761),
    .Y(_03795_));
 sg13g2_nor2_2 _10782_ (.A(net3776),
    .B(net3919),
    .Y(_03796_));
 sg13g2_or2_2 _10783_ (.X(_03797_),
    .B(net3919),
    .A(net3776));
 sg13g2_nor2_2 _10784_ (.A(net3708),
    .B(net3764),
    .Y(_03798_));
 sg13g2_nor2_2 _10785_ (.A(net3778),
    .B(net3776),
    .Y(_03799_));
 sg13g2_nand2b_2 _10786_ (.Y(_03800_),
    .B(_03718_),
    .A_N(net3778));
 sg13g2_nor2_2 _10787_ (.A(net3707),
    .B(net3767),
    .Y(_03801_));
 sg13g2_nor2_2 _10788_ (.A(_03736_),
    .B(net3764),
    .Y(_03802_));
 sg13g2_nor2_2 _10789_ (.A(_03736_),
    .B(net3766),
    .Y(_03803_));
 sg13g2_nor2_2 _10790_ (.A(net3776),
    .B(_03727_),
    .Y(_03804_));
 sg13g2_nor2_2 _10791_ (.A(_03722_),
    .B(net3767),
    .Y(_03805_));
 sg13g2_nor2_2 _10792_ (.A(_03722_),
    .B(net3761),
    .Y(_03806_));
 sg13g2_nor2_2 _10793_ (.A(_03727_),
    .B(_03766_),
    .Y(_03807_));
 sg13g2_nor2_2 _10794_ (.A(_03739_),
    .B(net3770),
    .Y(_03808_));
 sg13g2_nand2_2 _10795_ (.Y(_03809_),
    .A(_03738_),
    .B(_03758_));
 sg13g2_nor2_2 _10796_ (.A(_03735_),
    .B(_03774_),
    .Y(_03810_));
 sg13g2_nor2_2 _10797_ (.A(net3774),
    .B(net3761),
    .Y(_03811_));
 sg13g2_nor2_2 _10798_ (.A(net3774),
    .B(net3767),
    .Y(_03812_));
 sg13g2_nor2_2 _10799_ (.A(_03735_),
    .B(net3764),
    .Y(_03813_));
 sg13g2_nor2_2 _10800_ (.A(net3774),
    .B(net3768),
    .Y(_03814_));
 sg13g2_nand2b_2 _10801_ (.Y(_03815_),
    .B(_03758_),
    .A_N(net3774));
 sg13g2_nor2_2 _10802_ (.A(net3771),
    .B(net3760),
    .Y(_03816_));
 sg13g2_nor2_2 _10803_ (.A(_03736_),
    .B(net3769),
    .Y(_03817_));
 sg13g2_nand3_1 _10804_ (.B(_03726_),
    .C(_03758_),
    .A(_03707_),
    .Y(_03818_));
 sg13g2_nor2_2 _10805_ (.A(net3773),
    .B(net3761),
    .Y(_03819_));
 sg13g2_nor2_2 _10806_ (.A(net3773),
    .B(net3766),
    .Y(_03820_));
 sg13g2_nor2_2 _10807_ (.A(_03736_),
    .B(net3762),
    .Y(_03821_));
 sg13g2_nor2_2 _10808_ (.A(net3777),
    .B(_03739_),
    .Y(_03822_));
 sg13g2_nand2_2 _10809_ (.Y(_03823_),
    .A(_03718_),
    .B(_03738_));
 sg13g2_nor2_2 _10810_ (.A(net3777),
    .B(_03731_),
    .Y(_03824_));
 sg13g2_or2_2 _10811_ (.X(_03825_),
    .B(net3773),
    .A(net3777));
 sg13g2_nor2_2 _10812_ (.A(_03739_),
    .B(net3757),
    .Y(_03826_));
 sg13g2_nand2_2 _10813_ (.Y(_03827_),
    .A(_03738_),
    .B(_03773_));
 sg13g2_nor2_2 _10814_ (.A(_03724_),
    .B(net3767),
    .Y(_03828_));
 sg13g2_nor2_2 _10815_ (.A(net3773),
    .B(net3763),
    .Y(_03829_));
 sg13g2_nor2_2 _10816_ (.A(_03739_),
    .B(net3766),
    .Y(_03830_));
 sg13g2_nor2_2 _10817_ (.A(_03739_),
    .B(net3760),
    .Y(_03831_));
 sg13g2_nor2_2 _10818_ (.A(net3774),
    .B(net3757),
    .Y(_03832_));
 sg13g2_nor2_2 _10819_ (.A(net3777),
    .B(_03724_),
    .Y(_03833_));
 sg13g2_nor2_2 _10820_ (.A(_03739_),
    .B(net3763),
    .Y(_03834_));
 sg13g2_nor2_2 _10821_ (.A(_03741_),
    .B(net3765),
    .Y(_03835_));
 sg13g2_nor2_2 _10822_ (.A(_03735_),
    .B(net3768),
    .Y(_03836_));
 sg13g2_nand3_1 _10823_ (.B(_03734_),
    .C(_03758_),
    .A(_03726_),
    .Y(_03837_));
 sg13g2_nor2_2 _10824_ (.A(net3771),
    .B(net3759),
    .Y(_03838_));
 sg13g2_nor2_2 _10825_ (.A(net3773),
    .B(net3757),
    .Y(_03839_));
 sg13g2_nor2_2 _10826_ (.A(net3771),
    .B(net3768),
    .Y(_03840_));
 sg13g2_nand3_1 _10827_ (.B(_03726_),
    .C(_03758_),
    .A(_03704_),
    .Y(_03841_));
 sg13g2_nor2_2 _10828_ (.A(_03724_),
    .B(net3770),
    .Y(_03842_));
 sg13g2_nor2_2 _10829_ (.A(net3775),
    .B(_03736_),
    .Y(_03843_));
 sg13g2_nor2_2 _10830_ (.A(_03724_),
    .B(net3760),
    .Y(_03844_));
 sg13g2_nor2_2 _10831_ (.A(_03724_),
    .B(net3764),
    .Y(_03845_));
 sg13g2_nor2_2 _10832_ (.A(_03735_),
    .B(net3760),
    .Y(_03846_));
 sg13g2_nor2_2 _10833_ (.A(net3776),
    .B(net3771),
    .Y(_03847_));
 sg13g2_nor2_2 _10834_ (.A(_03736_),
    .B(net3759),
    .Y(_03848_));
 sg13g2_nor2_2 _10835_ (.A(net3775),
    .B(_03735_),
    .Y(_03849_));
 sg13g2_nand3_1 _10836_ (.B(_03726_),
    .C(_03734_),
    .A(_03718_),
    .Y(_03850_));
 sg13g2_nor2_2 _10837_ (.A(_03714_),
    .B(net3759),
    .Y(_03851_));
 sg13g2_nor2_2 _10838_ (.A(net3776),
    .B(net3772),
    .Y(_03852_));
 sg13g2_nor2_2 _10839_ (.A(_03712_),
    .B(net3765),
    .Y(_03853_));
 sg13g2_nand2_1 _10840_ (.Y(_03854_),
    .A(_03711_),
    .B(_03765_));
 sg13g2_nor2_2 _10841_ (.A(net3707),
    .B(net3761),
    .Y(_03855_));
 sg13g2_nor2_2 _10842_ (.A(_03712_),
    .B(net3768),
    .Y(_03856_));
 sg13g2_nand2_2 _10843_ (.Y(_03857_),
    .A(_03711_),
    .B(_03758_));
 sg13g2_a22oi_1 _10844_ (.Y(_03858_),
    .B1(_03856_),
    .B2(\spiking_network_top_uut.all_data_out[616] ),
    .A2(_03855_),
    .A1(\spiking_network_top_uut.all_data_out[328] ));
 sg13g2_nor2_2 _10845_ (.A(net3707),
    .B(net3765),
    .Y(_03859_));
 sg13g2_nand2b_2 _10846_ (.Y(_03860_),
    .B(_03765_),
    .A_N(net3707));
 sg13g2_nor2_2 _10847_ (.A(net3919),
    .B(net3763),
    .Y(_03861_));
 sg13g2_nor2_2 _10848_ (.A(net3779),
    .B(net3763),
    .Y(_03862_));
 sg13g2_nor2_2 _10849_ (.A(net3779),
    .B(net3777),
    .Y(_03863_));
 sg13g2_nor2_2 _10850_ (.A(net3772),
    .B(net3768),
    .Y(_03864_));
 sg13g2_nand2b_2 _10851_ (.Y(_03865_),
    .B(_03758_),
    .A_N(_03733_));
 sg13g2_nor2_2 _10852_ (.A(net3778),
    .B(net3762),
    .Y(_03866_));
 sg13g2_nor2_2 _10853_ (.A(net3779),
    .B(net3762),
    .Y(_03867_));
 sg13g2_nor2_2 _10854_ (.A(net3779),
    .B(net3757),
    .Y(_03868_));
 sg13g2_nor2_2 _10855_ (.A(_03712_),
    .B(net3761),
    .Y(_03869_));
 sg13g2_nor2_2 _10856_ (.A(_03746_),
    .B(net3760),
    .Y(_03870_));
 sg13g2_or2_2 _10857_ (.X(_03871_),
    .B(net3762),
    .A(net3708));
 sg13g2_nor2_2 _10858_ (.A(net3776),
    .B(net3708),
    .Y(_03872_));
 sg13g2_or2_2 _10859_ (.X(_03873_),
    .B(net3708),
    .A(net3776));
 sg13g2_nor2_2 _10860_ (.A(net3707),
    .B(net3758),
    .Y(_03874_));
 sg13g2_nand2b_2 _10861_ (.Y(_03875_),
    .B(_03773_),
    .A_N(net3707));
 sg13g2_nor2_2 _10862_ (.A(net3780),
    .B(net3760),
    .Y(_03876_));
 sg13g2_nor2_2 _10863_ (.A(net3771),
    .B(net3767),
    .Y(_03877_));
 sg13g2_nor2_2 _10864_ (.A(_03724_),
    .B(net3758),
    .Y(_03878_));
 sg13g2_nor2_2 _10865_ (.A(_03735_),
    .B(net3766),
    .Y(_03879_));
 sg13g2_nor2_2 _10866_ (.A(net3773),
    .B(net3769),
    .Y(_03880_));
 sg13g2_a21oi_2 _10867_ (.B1(net10),
    .Y(_03881_),
    .A2(_03694_),
    .A1(\spiking_network_top_uut.spi_inst.spi_slave_inst.bit_cnt[2] ));
 sg13g2_nor2_2 _10868_ (.A(_03733_),
    .B(net3759),
    .Y(_03882_));
 sg13g2_nor2_2 _10869_ (.A(net3778),
    .B(net3765),
    .Y(_03883_));
 sg13g2_nor2_2 _10870_ (.A(net3780),
    .B(net3758),
    .Y(_03884_));
 sg13g2_nor2_2 _10871_ (.A(_03722_),
    .B(net3769),
    .Y(_03885_));
 sg13g2_nand2_2 _10872_ (.Y(_03886_),
    .A(_03721_),
    .B(_03758_));
 sg13g2_nor2_2 _10873_ (.A(_03722_),
    .B(net3758),
    .Y(_03887_));
 sg13g2_nand2_2 _10874_ (.Y(_03888_),
    .A(_03721_),
    .B(_03773_));
 sg13g2_nor2_2 _10875_ (.A(net3779),
    .B(net3770),
    .Y(_03889_));
 sg13g2_nor2_2 _10876_ (.A(_03722_),
    .B(net3764),
    .Y(_03890_));
 sg13g2_nand2_2 _10877_ (.Y(_03891_),
    .A(_03721_),
    .B(_03765_));
 sg13g2_a22oi_1 _10878_ (.Y(_03892_),
    .B1(_03828_),
    .B2(\spiking_network_top_uut.all_data_out[224] ),
    .A2(_03822_),
    .A1(\spiking_network_top_uut.all_data_out[448] ));
 sg13g2_a22oi_1 _10879_ (.Y(_03893_),
    .B1(_03866_),
    .B2(\spiking_network_top_uut.all_data_out[296] ),
    .A2(net3694),
    .A1(\spiking_network_top_uut.all_data_out[80] ));
 sg13g2_a22oi_1 _10880_ (.Y(_03894_),
    .B1(_03868_),
    .B2(\spiking_network_top_uut.all_data_out[824] ),
    .A2(_03788_),
    .A1(\spiking_network_top_uut.all_data_out[152] ));
 sg13g2_a22oi_1 _10881_ (.Y(_03895_),
    .B1(_03889_),
    .B2(\spiking_network_top_uut.all_data_out[568] ),
    .A2(_03779_),
    .A1(net4286));
 sg13g2_a22oi_1 _10882_ (.Y(_03896_),
    .B1(_03884_),
    .B2(\spiking_network_top_uut.all_data_out[792] ),
    .A2(_03883_),
    .A1(\spiking_network_top_uut.all_data_out[680] ));
 sg13g2_a22oi_1 _10883_ (.Y(_03897_),
    .B1(_03874_),
    .B2(\spiking_network_top_uut.all_data_out[840] ),
    .A2(net3712),
    .A1(\spiking_network_top_uut.all_data_out[120] ));
 sg13g2_a22oi_1 _10884_ (.Y(_03898_),
    .B1(_03844_),
    .B2(\spiking_network_top_uut.all_data_out[352] ),
    .A2(net3717),
    .A1(\spiking_network_top_uut.all_data_out[104] ));
 sg13g2_a22oi_1 _10885_ (.Y(_03899_),
    .B1(net3718),
    .B2(\spiking_network_top_uut.all_data_out[56] ),
    .A2(net3719),
    .A1(\spiking_network_top_uut.all_data_out[24] ));
 sg13g2_nand4_1 _10886_ (.B(_03892_),
    .C(_03898_),
    .A(_03858_),
    .Y(_03900_),
    .D(_03899_));
 sg13g2_a22oi_1 _10887_ (.Y(_03901_),
    .B1(_03880_),
    .B2(\spiking_network_top_uut.all_data_out[544] ),
    .A2(_03863_),
    .A1(\spiking_network_top_uut.all_data_out[440] ));
 sg13g2_a22oi_1 _10888_ (.Y(_03902_),
    .B1(_03846_),
    .B2(\spiking_network_top_uut.all_data_out[336] ),
    .A2(_03764_),
    .A1(\spiking_network_top_uut.all_data_out[552] ));
 sg13g2_nand4_1 _10889_ (.B(_03894_),
    .C(_03901_),
    .A(_03893_),
    .Y(_03903_),
    .D(_03902_));
 sg13g2_a22oi_1 _10890_ (.Y(_03904_),
    .B1(_03867_),
    .B2(\spiking_network_top_uut.all_data_out[312] ),
    .A2(_03776_),
    .A1(\spiking_network_top_uut.all_data_out[168] ));
 sg13g2_a22oi_1 _10891_ (.Y(_03905_),
    .B1(_03851_),
    .B2(\spiking_network_top_uut.all_data_out[808] ),
    .A2(_03816_),
    .A1(\spiking_network_top_uut.all_data_out[272] ));
 sg13g2_a22oi_1 _10892_ (.Y(_03906_),
    .B1(_03842_),
    .B2(\spiking_network_top_uut.all_data_out[608] ),
    .A2(_03821_),
    .A1(\spiking_network_top_uut.all_data_out[304] ));
 sg13g2_a22oi_1 _10893_ (.Y(_03907_),
    .B1(_03848_),
    .B2(\spiking_network_top_uut.all_data_out[816] ),
    .A2(_03829_),
    .A1(\spiking_network_top_uut.all_data_out[672] ));
 sg13g2_nand4_1 _10894_ (.B(_03905_),
    .C(_03906_),
    .A(_03904_),
    .Y(_03908_),
    .D(_03907_));
 sg13g2_a22oi_1 _10895_ (.Y(_03909_),
    .B1(_03882_),
    .B2(\spiking_network_top_uut.all_data_out[776] ),
    .A2(_03767_),
    .A1(\spiking_network_top_uut.all_data_out[648] ));
 sg13g2_a22oi_1 _10896_ (.Y(_03910_),
    .B1(_03864_),
    .B2(\spiking_network_top_uut.all_data_out[520] ),
    .A2(_03859_),
    .A1(\spiking_network_top_uut.all_data_out[712] ));
 sg13g2_a22oi_1 _10897_ (.Y(_03911_),
    .B1(_03852_),
    .B2(\spiking_network_top_uut.all_data_out[392] ),
    .A2(_03849_),
    .A1(\spiking_network_top_uut.all_data_out[464] ));
 sg13g2_a22oi_1 _10898_ (.Y(_03912_),
    .B1(_03847_),
    .B2(\spiking_network_top_uut.all_data_out[400] ),
    .A2(_03843_),
    .A1(\spiking_network_top_uut.all_data_out[432] ));
 sg13g2_nand4_1 _10899_ (.B(_03910_),
    .C(_03911_),
    .A(_03909_),
    .Y(_03913_),
    .D(_03912_));
 sg13g2_nor4_1 _10900_ (.A(_03900_),
    .B(_03903_),
    .C(_03908_),
    .D(_03913_),
    .Y(_03914_));
 sg13g2_a22oi_1 _10901_ (.Y(_03915_),
    .B1(_03819_),
    .B2(\spiking_network_top_uut.all_data_out[288] ),
    .A2(net3695),
    .A1(\spiking_network_top_uut.all_data_out[88] ));
 sg13g2_a22oi_1 _10902_ (.Y(_03916_),
    .B1(_03760_),
    .B2(\spiking_network_top_uut.all_data_out[600] ),
    .A2(net3693),
    .A1(\spiking_network_top_uut.all_data_out[72] ));
 sg13g2_a22oi_1 _10903_ (.Y(_03917_),
    .B1(_03832_),
    .B2(\spiking_network_top_uut.all_data_out[880] ),
    .A2(_03830_),
    .A1(\spiking_network_top_uut.all_data_out[192] ));
 sg13g2_a22oi_1 _10904_ (.Y(_03918_),
    .B1(_03869_),
    .B2(\spiking_network_top_uut.all_data_out[360] ),
    .A2(_03782_),
    .A1(\spiking_network_top_uut.all_data_out[136] ));
 sg13g2_nand4_1 _10905_ (.B(_03916_),
    .C(_03917_),
    .A(_03915_),
    .Y(_03919_),
    .D(_03918_));
 sg13g2_a22oi_1 _10906_ (.Y(_03920_),
    .B1(_03805_),
    .B2(\spiking_network_top_uut.all_data_out[128] ),
    .A2(net3710),
    .A1(\spiking_network_top_uut.all_data_out[48] ));
 sg13g2_a22oi_1 _10907_ (.Y(_03921_),
    .B1(_03817_),
    .B2(\spiking_network_top_uut.all_data_out[560] ),
    .A2(_03744_),
    .A1(\spiking_network_top_uut.all_data_out[896] ));
 sg13g2_a22oi_1 _10908_ (.Y(_03922_),
    .B1(net3711),
    .B2(\spiking_network_top_uut.all_data_out[32] ),
    .A2(net3715),
    .A1(\spiking_network_top_uut.all_data_out[384] ));
 sg13g2_a22oi_1 _10909_ (.Y(_03923_),
    .B1(_03796_),
    .B2(\spiking_network_top_uut.all_data_out[504] ),
    .A2(_03783_),
    .A1(\spiking_network_top_uut.all_data_out[456] ));
 sg13g2_nand4_1 _10910_ (.B(_03921_),
    .C(_03922_),
    .A(_03920_),
    .Y(_03924_),
    .D(_03923_));
 sg13g2_a22oi_1 _10911_ (.Y(_03925_),
    .B1(_03885_),
    .B2(\spiking_network_top_uut.all_data_out[512] ),
    .A2(_03811_),
    .A1(\spiking_network_top_uut.all_data_out[368] ));
 sg13g2_a22oi_1 _10912_ (.Y(_03926_),
    .B1(_03831_),
    .B2(\spiking_network_top_uut.all_data_out[320] ),
    .A2(net3716),
    .A1(\spiking_network_top_uut.all_data_out[40] ));
 sg13g2_a22oi_1 _10913_ (.Y(_03927_),
    .B1(_03836_),
    .B2(\spiking_network_top_uut.all_data_out[592] ),
    .A2(_03777_),
    .A1(\spiking_network_top_uut.all_data_out[408] ));
 sg13g2_a22oi_1 _10914_ (.Y(_03928_),
    .B1(_03799_),
    .B2(\spiking_network_top_uut.all_data_out[424] ),
    .A2(net3714),
    .A1(\spiking_network_top_uut.all_data_out[96] ));
 sg13g2_nand4_1 _10915_ (.B(_03926_),
    .C(_03927_),
    .A(_03925_),
    .Y(_03929_),
    .D(_03928_));
 sg13g2_a22oi_1 _10916_ (.Y(_03930_),
    .B1(net3696),
    .B2(\spiking_network_top_uut.all_data_out[64] ),
    .A2(net3713),
    .A1(\spiking_network_top_uut.all_data_out[112] ));
 sg13g2_a22oi_1 _10917_ (.Y(_03931_),
    .B1(_03853_),
    .B2(\spiking_network_top_uut.all_data_out[744] ),
    .A2(_03824_),
    .A1(\spiking_network_top_uut.all_data_out[416] ));
 sg13g2_nand4_1 _10918_ (.B(_03896_),
    .C(_03930_),
    .A(_03895_),
    .Y(_03932_),
    .D(_03931_));
 sg13g2_nor4_2 _10919_ (.A(_03919_),
    .B(_03924_),
    .C(_03929_),
    .Y(_03933_),
    .D(_03932_));
 sg13g2_a22oi_1 _10920_ (.Y(_03934_),
    .B1(_03861_),
    .B2(\spiking_network_top_uut.all_data_out[760] ),
    .A2(_03785_),
    .A1(\spiking_network_top_uut.all_data_out[248] ));
 sg13g2_a22oi_1 _10921_ (.Y(_03935_),
    .B1(_03826_),
    .B2(\spiking_network_top_uut.all_data_out[832] ),
    .A2(_03813_),
    .A1(\spiking_network_top_uut.all_data_out[720] ));
 sg13g2_a22oi_1 _10922_ (.Y(_03936_),
    .B1(_03802_),
    .B2(\spiking_network_top_uut.all_data_out[688] ),
    .A2(_03780_),
    .A1(\spiking_network_top_uut.all_data_out[216] ));
 sg13g2_nand4_1 _10923_ (.B(_03934_),
    .C(_03935_),
    .A(_03897_),
    .Y(_03937_),
    .D(_03936_));
 sg13g2_a22oi_1 _10924_ (.Y(_03938_),
    .B1(_03807_),
    .B2(\spiking_network_top_uut.all_data_out[752] ),
    .A2(_03786_),
    .A1(\spiking_network_top_uut.all_data_out[488] ));
 sg13g2_a22oi_1 _10925_ (.Y(_03939_),
    .B1(_03803_),
    .B2(\spiking_network_top_uut.all_data_out[176] ),
    .A2(_03798_),
    .A1(\spiking_network_top_uut.all_data_out[728] ));
 sg13g2_a22oi_1 _10926_ (.Y(_03940_),
    .B1(_03810_),
    .B2(\spiking_network_top_uut.all_data_out[848] ),
    .A2(_03794_),
    .A1(\spiking_network_top_uut.all_data_out[536] ));
 sg13g2_a22oi_1 _10927_ (.Y(_03941_),
    .B1(_03833_),
    .B2(\spiking_network_top_uut.all_data_out[480] ),
    .A2(_03812_),
    .A1(\spiking_network_top_uut.all_data_out[240] ));
 sg13g2_nand4_1 _10928_ (.B(_03939_),
    .C(_03940_),
    .A(_03938_),
    .Y(_03942_),
    .D(_03941_));
 sg13g2_nor2_1 _10929_ (.A(_03937_),
    .B(_03942_),
    .Y(_03943_));
 sg13g2_a22oi_1 _10930_ (.Y(_03944_),
    .B1(_03839_),
    .B2(\spiking_network_top_uut.all_data_out[800] ),
    .A2(_03781_),
    .A1(\spiking_network_top_uut.all_data_out[632] ));
 sg13g2_a22oi_1 _10931_ (.Y(_03945_),
    .B1(_03877_),
    .B2(\spiking_network_top_uut.all_data_out[144] ),
    .A2(net3709),
    .A1(net4316));
 sg13g2_a22oi_1 _10932_ (.Y(_03946_),
    .B1(_03834_),
    .B2(\spiking_network_top_uut.all_data_out[704] ),
    .A2(_03814_),
    .A1(\spiking_network_top_uut.all_data_out[624] ));
 sg13g2_nand4_1 _10933_ (.B(_03944_),
    .C(_03945_),
    .A(_03793_),
    .Y(_03947_),
    .D(_03946_));
 sg13g2_a22oi_1 _10934_ (.Y(_03948_),
    .B1(_03862_),
    .B2(\spiking_network_top_uut.all_data_out[696] ),
    .A2(_03789_),
    .A1(\spiking_network_top_uut.all_data_out[872] ));
 sg13g2_a22oi_1 _10935_ (.Y(_03949_),
    .B1(_03890_),
    .B2(\spiking_network_top_uut.all_data_out[640] ),
    .A2(_03840_),
    .A1(\spiking_network_top_uut.all_data_out[528] ));
 sg13g2_a22oi_1 _10936_ (.Y(_03950_),
    .B1(_03876_),
    .B2(\spiking_network_top_uut.all_data_out[280] ),
    .A2(_03870_),
    .A1(\spiking_network_top_uut.all_data_out[344] ));
 sg13g2_a22oi_1 _10937_ (.Y(_03951_),
    .B1(_03872_),
    .B2(\spiking_network_top_uut.all_data_out[472] ),
    .A2(_03795_),
    .A1(\spiking_network_top_uut.all_data_out[264] ));
 sg13g2_nand4_1 _10938_ (.B(_03949_),
    .C(_03950_),
    .A(_03948_),
    .Y(_03952_),
    .D(_03951_));
 sg13g2_a22oi_1 _10939_ (.Y(_03953_),
    .B1(_03845_),
    .B2(\spiking_network_top_uut.all_data_out[736] ),
    .A2(_03838_),
    .A1(\spiking_network_top_uut.all_data_out[784] ));
 sg13g2_a22oi_1 _10940_ (.Y(_03954_),
    .B1(_03835_),
    .B2(\spiking_network_top_uut.all_data_out[656] ),
    .A2(_03763_),
    .A1(\spiking_network_top_uut.all_data_out[184] ));
 sg13g2_a22oi_1 _10941_ (.Y(_03955_),
    .B1(_03820_),
    .B2(\spiking_network_top_uut.all_data_out[160] ),
    .A2(_03769_),
    .A1(\spiking_network_top_uut.all_data_out[664] ));
 sg13g2_a22oi_1 _10942_ (.Y(_03956_),
    .B1(_03804_),
    .B2(\spiking_network_top_uut.all_data_out[496] ),
    .A2(_03784_),
    .A1(\spiking_network_top_uut.all_data_out[584] ));
 sg13g2_nand4_1 _10943_ (.B(_03954_),
    .C(_03955_),
    .A(_03953_),
    .Y(_03957_),
    .D(_03956_));
 sg13g2_a22oi_1 _10944_ (.Y(_03958_),
    .B1(_03887_),
    .B2(\spiking_network_top_uut.all_data_out[768] ),
    .A2(_03806_),
    .A1(\spiking_network_top_uut.all_data_out[256] ));
 sg13g2_a22oi_1 _10945_ (.Y(_03959_),
    .B1(_03808_),
    .B2(\spiking_network_top_uut.all_data_out[576] ),
    .A2(_03772_),
    .A1(\spiking_network_top_uut.all_data_out[376] ));
 sg13g2_a22oi_1 _10946_ (.Y(_03960_),
    .B1(_03879_),
    .B2(\spiking_network_top_uut.all_data_out[208] ),
    .A2(_03775_),
    .A1(\spiking_network_top_uut.all_data_out[856] ));
 sg13g2_a22oi_1 _10947_ (.Y(_03961_),
    .B1(_03878_),
    .B2(\spiking_network_top_uut.all_data_out[864] ),
    .A2(_03801_),
    .A1(\spiking_network_top_uut.all_data_out[200] ));
 sg13g2_nand4_1 _10948_ (.B(_03959_),
    .C(_03960_),
    .A(_03958_),
    .Y(_03962_),
    .D(_03961_));
 sg13g2_nor4_1 _10949_ (.A(_03947_),
    .B(_03952_),
    .C(_03957_),
    .D(_03962_),
    .Y(_03963_));
 sg13g2_and4_2 _10950_ (.A(_03914_),
    .B(_03933_),
    .C(_03943_),
    .D(_03963_),
    .X(_03964_));
 sg13g2_a21oi_1 _10951_ (.A1(\spiking_network_top_uut.all_data_out[0] ),
    .A2(_03756_),
    .Y(_03965_),
    .B1(_03881_));
 sg13g2_a22oi_1 _10952_ (.Y(_03966_),
    .B1(_03833_),
    .B2(\spiking_network_top_uut.all_data_out[487] ),
    .A2(_03821_),
    .A1(\spiking_network_top_uut.all_data_out[311] ));
 sg13g2_a22oi_1 _10953_ (.Y(_03967_),
    .B1(_03812_),
    .B2(\spiking_network_top_uut.all_data_out[247] ),
    .A2(_03767_),
    .A1(\spiking_network_top_uut.all_data_out[655] ));
 sg13g2_a22oi_1 _10954_ (.Y(_03968_),
    .B1(_03813_),
    .B2(\spiking_network_top_uut.all_data_out[727] ),
    .A2(_03706_),
    .A1(\spiking_network_top_uut.all_data_out[31] ));
 sg13g2_a22oi_1 _10955_ (.Y(_03969_),
    .B1(_03851_),
    .B2(\spiking_network_top_uut.all_data_out[815] ),
    .A2(_03847_),
    .A1(\spiking_network_top_uut.all_data_out[407] ));
 sg13g2_a22oi_1 _10956_ (.Y(_03970_),
    .B1(_03877_),
    .B2(\spiking_network_top_uut.all_data_out[151] ),
    .A2(_03781_),
    .A1(\spiking_network_top_uut.all_data_out[639] ));
 sg13g2_a22oi_1 _10957_ (.Y(_03971_),
    .B1(_03882_),
    .B2(\spiking_network_top_uut.all_data_out[783] ),
    .A2(_03803_),
    .A1(\spiking_network_top_uut.all_data_out[183] ));
 sg13g2_a22oi_1 _10958_ (.Y(_03972_),
    .B1(_03870_),
    .B2(\spiking_network_top_uut.all_data_out[351] ),
    .A2(_03785_),
    .A1(\spiking_network_top_uut.all_data_out[255] ));
 sg13g2_a22oi_1 _10959_ (.Y(_03973_),
    .B1(_03879_),
    .B2(\spiking_network_top_uut.all_data_out[215] ),
    .A2(_03862_),
    .A1(\spiking_network_top_uut.all_data_out[703] ));
 sg13g2_a22oi_1 _10960_ (.Y(_03974_),
    .B1(_03884_),
    .B2(\spiking_network_top_uut.all_data_out[799] ),
    .A2(_03776_),
    .A1(\spiking_network_top_uut.all_data_out[175] ));
 sg13g2_a22oi_1 _10961_ (.Y(_03975_),
    .B1(_03855_),
    .B2(\spiking_network_top_uut.all_data_out[335] ),
    .A2(_03760_),
    .A1(\spiking_network_top_uut.all_data_out[607] ));
 sg13g2_a22oi_1 _10962_ (.Y(_03976_),
    .B1(_03822_),
    .B2(\spiking_network_top_uut.all_data_out[455] ),
    .A2(net3696),
    .A1(\spiking_network_top_uut.all_data_out[71] ));
 sg13g2_a22oi_1 _10963_ (.Y(_03977_),
    .B1(_03796_),
    .B2(\spiking_network_top_uut.all_data_out[511] ),
    .A2(_03763_),
    .A1(\spiking_network_top_uut.all_data_out[191] ));
 sg13g2_a22oi_1 _10964_ (.Y(_03978_),
    .B1(_03826_),
    .B2(\spiking_network_top_uut.all_data_out[839] ),
    .A2(_03744_),
    .A1(\spiking_network_top_uut.all_data_out[903] ));
 sg13g2_a22oi_1 _10965_ (.Y(_03979_),
    .B1(_03820_),
    .B2(\spiking_network_top_uut.all_data_out[167] ),
    .A2(_03814_),
    .A1(\spiking_network_top_uut.all_data_out[631] ));
 sg13g2_a22oi_1 _10966_ (.Y(_03980_),
    .B1(_03887_),
    .B2(\spiking_network_top_uut.all_data_out[775] ),
    .A2(_03792_),
    .A1(\spiking_network_top_uut.all_data_out[239] ));
 sg13g2_nand4_1 _10967_ (.B(_03978_),
    .C(_03979_),
    .A(_03971_),
    .Y(_03981_),
    .D(_03980_));
 sg13g2_a22oi_1 _10968_ (.Y(_03982_),
    .B1(_03864_),
    .B2(\spiking_network_top_uut.all_data_out[527] ),
    .A2(_03845_),
    .A1(\spiking_network_top_uut.all_data_out[743] ));
 sg13g2_a22oi_1 _10969_ (.Y(_03983_),
    .B1(_03843_),
    .B2(\spiking_network_top_uut.all_data_out[439] ),
    .A2(net3695),
    .A1(\spiking_network_top_uut.all_data_out[95] ));
 sg13g2_a22oi_1 _10970_ (.Y(_03984_),
    .B1(_03861_),
    .B2(\spiking_network_top_uut.all_data_out[767] ),
    .A2(net3710),
    .A1(\spiking_network_top_uut.all_data_out[55] ));
 sg13g2_a22oi_1 _10971_ (.Y(_03985_),
    .B1(_03788_),
    .B2(\spiking_network_top_uut.all_data_out[159] ),
    .A2(_03777_),
    .A1(\spiking_network_top_uut.all_data_out[415] ));
 sg13g2_nand4_1 _10972_ (.B(_03983_),
    .C(_03984_),
    .A(_03982_),
    .Y(_03986_),
    .D(_03985_));
 sg13g2_a22oi_1 _10973_ (.Y(_03987_),
    .B1(_03876_),
    .B2(\spiking_network_top_uut.all_data_out[287] ),
    .A2(_03799_),
    .A1(\spiking_network_top_uut.all_data_out[431] ));
 sg13g2_a22oi_1 _10974_ (.Y(_03988_),
    .B1(_03842_),
    .B2(\spiking_network_top_uut.all_data_out[615] ),
    .A2(_03790_),
    .A1(\spiking_network_top_uut.all_data_out[895] ));
 sg13g2_a22oi_1 _10975_ (.Y(_03989_),
    .B1(_03836_),
    .B2(\spiking_network_top_uut.all_data_out[599] ),
    .A2(_03829_),
    .A1(\spiking_network_top_uut.all_data_out[679] ));
 sg13g2_a22oi_1 _10976_ (.Y(_03990_),
    .B1(_03832_),
    .B2(\spiking_network_top_uut.all_data_out[887] ),
    .A2(net3709),
    .A1(\spiking_network_top_uut.all_data_out[23] ));
 sg13g2_nand4_1 _10977_ (.B(_03988_),
    .C(_03989_),
    .A(_03987_),
    .Y(_03991_),
    .D(_03990_));
 sg13g2_a22oi_1 _10978_ (.Y(_03992_),
    .B1(_03839_),
    .B2(\spiking_network_top_uut.all_data_out[807] ),
    .A2(_03806_),
    .A1(\spiking_network_top_uut.all_data_out[263] ));
 sg13g2_a22oi_1 _10979_ (.Y(_03993_),
    .B1(_03872_),
    .B2(\spiking_network_top_uut.all_data_out[479] ),
    .A2(_03786_),
    .A1(\spiking_network_top_uut.all_data_out[495] ));
 sg13g2_a22oi_1 _10980_ (.Y(_03994_),
    .B1(_03783_),
    .B2(\spiking_network_top_uut.all_data_out[463] ),
    .A2(net3693),
    .A1(\spiking_network_top_uut.all_data_out[79] ));
 sg13g2_a22oi_1 _10981_ (.Y(_03995_),
    .B1(_03804_),
    .B2(\spiking_network_top_uut.all_data_out[503] ),
    .A2(_03784_),
    .A1(\spiking_network_top_uut.all_data_out[591] ));
 sg13g2_nand4_1 _10982_ (.B(_03993_),
    .C(_03994_),
    .A(_03992_),
    .Y(_03996_),
    .D(_03995_));
 sg13g2_or4_1 _10983_ (.A(_03981_),
    .B(_03986_),
    .C(_03991_),
    .D(_03996_),
    .X(_03997_));
 sg13g2_a22oi_1 _10984_ (.Y(_03998_),
    .B1(_03863_),
    .B2(\spiking_network_top_uut.all_data_out[447] ),
    .A2(_03828_),
    .A1(\spiking_network_top_uut.all_data_out[231] ));
 sg13g2_a22oi_1 _10985_ (.Y(_03999_),
    .B1(_03831_),
    .B2(\spiking_network_top_uut.all_data_out[327] ),
    .A2(_03764_),
    .A1(\spiking_network_top_uut.all_data_out[559] ));
 sg13g2_a22oi_1 _10986_ (.Y(_04000_),
    .B1(_03853_),
    .B2(\spiking_network_top_uut.all_data_out[751] ),
    .A2(net3716),
    .A1(\spiking_network_top_uut.all_data_out[47] ));
 sg13g2_nand4_1 _10987_ (.B(_03998_),
    .C(_03999_),
    .A(_03977_),
    .Y(_04001_),
    .D(_04000_));
 sg13g2_a22oi_1 _10988_ (.Y(_04002_),
    .B1(_03848_),
    .B2(\spiking_network_top_uut.all_data_out[823] ),
    .A2(_03810_),
    .A1(\spiking_network_top_uut.all_data_out[855] ));
 sg13g2_a22oi_1 _10989_ (.Y(_04003_),
    .B1(_03849_),
    .B2(\spiking_network_top_uut.all_data_out[471] ),
    .A2(net3717),
    .A1(\spiking_network_top_uut.all_data_out[111] ));
 sg13g2_a22oi_1 _10990_ (.Y(_04004_),
    .B1(_03852_),
    .B2(\spiking_network_top_uut.all_data_out[399] ),
    .A2(_03811_),
    .A1(\spiking_network_top_uut.all_data_out[375] ));
 sg13g2_a22oi_1 _10991_ (.Y(_04005_),
    .B1(_03878_),
    .B2(\spiking_network_top_uut.all_data_out[871] ),
    .A2(net3694),
    .A1(\spiking_network_top_uut.all_data_out[87] ));
 sg13g2_nand4_1 _10992_ (.B(_04003_),
    .C(_04004_),
    .A(_04002_),
    .Y(_04006_),
    .D(_04005_));
 sg13g2_nor4_2 _10993_ (.A(_03756_),
    .B(_03997_),
    .C(_04001_),
    .Y(_04007_),
    .D(_04006_));
 sg13g2_nand4_1 _10994_ (.B(_03972_),
    .C(_03973_),
    .A(_03970_),
    .Y(_04008_),
    .D(_03976_));
 sg13g2_a22oi_1 _10995_ (.Y(_04009_),
    .B1(_03890_),
    .B2(\spiking_network_top_uut.all_data_out[647] ),
    .A2(_03867_),
    .A1(\spiking_network_top_uut.all_data_out[319] ));
 sg13g2_a22oi_1 _10996_ (.Y(_04010_),
    .B1(_03846_),
    .B2(\spiking_network_top_uut.all_data_out[343] ),
    .A2(net3713),
    .A1(\spiking_network_top_uut.all_data_out[119] ));
 sg13g2_a22oi_1 _10997_ (.Y(_04011_),
    .B1(_03772_),
    .B2(\spiking_network_top_uut.all_data_out[383] ),
    .A2(net3718),
    .A1(\spiking_network_top_uut.all_data_out[63] ));
 sg13g2_a22oi_1 _10998_ (.Y(_04012_),
    .B1(_03844_),
    .B2(\spiking_network_top_uut.all_data_out[359] ),
    .A2(_03802_),
    .A1(\spiking_network_top_uut.all_data_out[695] ));
 sg13g2_nand4_1 _10999_ (.B(_04010_),
    .C(_04011_),
    .A(_04009_),
    .Y(_04013_),
    .D(_04012_));
 sg13g2_a22oi_1 _11000_ (.Y(_04014_),
    .B1(_03883_),
    .B2(\spiking_network_top_uut.all_data_out[687] ),
    .A2(net3711),
    .A1(\spiking_network_top_uut.all_data_out[39] ));
 sg13g2_a22oi_1 _11001_ (.Y(_04015_),
    .B1(_03856_),
    .B2(\spiking_network_top_uut.all_data_out[623] ),
    .A2(_03780_),
    .A1(\spiking_network_top_uut.all_data_out[223] ));
 sg13g2_a22oi_1 _11002_ (.Y(_04016_),
    .B1(_03789_),
    .B2(\spiking_network_top_uut.all_data_out[879] ),
    .A2(net3714),
    .A1(\spiking_network_top_uut.all_data_out[103] ));
 sg13g2_a22oi_1 _11003_ (.Y(_04017_),
    .B1(_03869_),
    .B2(\spiking_network_top_uut.all_data_out[367] ),
    .A2(_03824_),
    .A1(\spiking_network_top_uut.all_data_out[423] ));
 sg13g2_nand4_1 _11004_ (.B(_04015_),
    .C(_04016_),
    .A(_04014_),
    .Y(_04018_),
    .D(_04017_));
 sg13g2_a22oi_1 _11005_ (.Y(_04019_),
    .B1(_03808_),
    .B2(\spiking_network_top_uut.all_data_out[583] ),
    .A2(_03795_),
    .A1(\spiking_network_top_uut.all_data_out[271] ));
 sg13g2_a22oi_1 _11006_ (.Y(_04020_),
    .B1(_03889_),
    .B2(\spiking_network_top_uut.all_data_out[575] ),
    .A2(_03805_),
    .A1(\spiking_network_top_uut.all_data_out[135] ));
 sg13g2_a22oi_1 _11007_ (.Y(_04021_),
    .B1(_03840_),
    .B2(\spiking_network_top_uut.all_data_out[535] ),
    .A2(_03794_),
    .A1(\spiking_network_top_uut.all_data_out[543] ));
 sg13g2_nand4_1 _11008_ (.B(_04019_),
    .C(_04020_),
    .A(_03966_),
    .Y(_04022_),
    .D(_04021_));
 sg13g2_nor4_1 _11009_ (.A(_04008_),
    .B(_04013_),
    .C(_04018_),
    .D(_04022_),
    .Y(_04023_));
 sg13g2_a22oi_1 _11010_ (.Y(_04024_),
    .B1(_03807_),
    .B2(\spiking_network_top_uut.all_data_out[759] ),
    .A2(_03801_),
    .A1(\spiking_network_top_uut.all_data_out[207] ));
 sg13g2_a22oi_1 _11011_ (.Y(_04025_),
    .B1(_03866_),
    .B2(\spiking_network_top_uut.all_data_out[303] ),
    .A2(_03830_),
    .A1(\spiking_network_top_uut.all_data_out[199] ));
 sg13g2_a22oi_1 _11012_ (.Y(_04026_),
    .B1(_03885_),
    .B2(\spiking_network_top_uut.all_data_out[519] ),
    .A2(_03838_),
    .A1(\spiking_network_top_uut.all_data_out[791] ));
 sg13g2_nand4_1 _11013_ (.B(_04024_),
    .C(_04025_),
    .A(_03975_),
    .Y(_04027_),
    .D(_04026_));
 sg13g2_a22oi_1 _11014_ (.Y(_04028_),
    .B1(_03834_),
    .B2(\spiking_network_top_uut.all_data_out[711] ),
    .A2(_03775_),
    .A1(\spiking_network_top_uut.all_data_out[863] ));
 sg13g2_a22oi_1 _11015_ (.Y(_04029_),
    .B1(_03859_),
    .B2(\spiking_network_top_uut.all_data_out[719] ),
    .A2(net3712),
    .A1(\spiking_network_top_uut.all_data_out[127] ));
 sg13g2_a22oi_1 _11016_ (.Y(_04030_),
    .B1(_03819_),
    .B2(\spiking_network_top_uut.all_data_out[295] ),
    .A2(_03816_),
    .A1(\spiking_network_top_uut.all_data_out[279] ));
 sg13g2_nand4_1 _11017_ (.B(_04028_),
    .C(_04029_),
    .A(_03974_),
    .Y(_04031_),
    .D(_04030_));
 sg13g2_a22oi_1 _11018_ (.Y(_04032_),
    .B1(_03874_),
    .B2(\spiking_network_top_uut.all_data_out[847] ),
    .A2(_03817_),
    .A1(\spiking_network_top_uut.all_data_out[567] ));
 sg13g2_a22oi_1 _11019_ (.Y(_04033_),
    .B1(_03868_),
    .B2(\spiking_network_top_uut.all_data_out[831] ),
    .A2(net3715),
    .A1(\spiking_network_top_uut.all_data_out[391] ));
 sg13g2_a22oi_1 _11020_ (.Y(_04034_),
    .B1(_03779_),
    .B2(\spiking_network_top_uut.all_data_out[15] ),
    .A2(_03769_),
    .A1(\spiking_network_top_uut.all_data_out[671] ));
 sg13g2_a22oi_1 _11021_ (.Y(_04035_),
    .B1(_03798_),
    .B2(\spiking_network_top_uut.all_data_out[735] ),
    .A2(_03782_),
    .A1(\spiking_network_top_uut.all_data_out[143] ));
 sg13g2_nand4_1 _11022_ (.B(_04033_),
    .C(_04034_),
    .A(_04032_),
    .Y(_04036_),
    .D(_04035_));
 sg13g2_a22oi_1 _11023_ (.Y(_04037_),
    .B1(_03880_),
    .B2(\spiking_network_top_uut.all_data_out[551] ),
    .A2(_03835_),
    .A1(\spiking_network_top_uut.all_data_out[663] ));
 sg13g2_nand4_1 _11024_ (.B(_03968_),
    .C(_03969_),
    .A(_03967_),
    .Y(_04038_),
    .D(_04037_));
 sg13g2_nor4_1 _11025_ (.A(_04027_),
    .B(_04031_),
    .C(_04036_),
    .D(_04038_),
    .Y(_04039_));
 sg13g2_nand3_1 _11026_ (.B(_04023_),
    .C(_04039_),
    .A(_04007_),
    .Y(_04040_));
 sg13g2_o21ai_1 _11027_ (.B1(_04040_),
    .Y(_04041_),
    .A1(\spiking_network_top_uut.all_data_out[7] ),
    .A2(_03757_));
 sg13g2_nor2_1 _11028_ (.A(\spiking_network_top_uut.spi_inst.spi_slave_inst.bit_cnt[0] ),
    .B(_04041_),
    .Y(_04042_));
 sg13g2_nand2b_2 _11029_ (.Y(_04043_),
    .B(_03832_),
    .A_N(_00142_));
 sg13g2_nand2b_1 _11030_ (.Y(_04044_),
    .B(_03814_),
    .A_N(_00174_));
 sg13g2_nor2_2 _11031_ (.A(_00200_),
    .B(_03825_),
    .Y(_04045_));
 sg13g2_nand2b_2 _11032_ (.Y(_04046_),
    .B(_03829_),
    .A_N(_00168_));
 sg13g2_nand2b_1 _11033_ (.Y(_04047_),
    .B(_03839_),
    .A_N(_00152_));
 sg13g2_nand2b_1 _11034_ (.Y(_04048_),
    .B(_03810_),
    .A_N(_00146_));
 sg13g2_nand2b_1 _11035_ (.Y(_04049_),
    .B(_03842_),
    .A_N(_00176_));
 sg13g2_nor3_1 _11036_ (.A(_00198_),
    .B(net3775),
    .C(_03736_),
    .Y(_04050_));
 sg13g2_nand2b_2 _11037_ (.Y(_04051_),
    .B(_03844_),
    .A_N(_00208_));
 sg13g2_nand2b_1 _11038_ (.Y(_04052_),
    .B(_03811_),
    .A_N(_00206_));
 sg13g2_nand2b_1 _11039_ (.Y(_04053_),
    .B(_03826_),
    .A_N(_00148_));
 sg13g2_nand2b_1 _11040_ (.Y(_04054_),
    .B(_03799_),
    .A_N(_00199_));
 sg13g2_nand2b_2 _11041_ (.Y(_04055_),
    .B(_03775_),
    .A_N(_00145_));
 sg13g2_nand2b_1 _11042_ (.Y(_04056_),
    .B(_03794_),
    .A_N(_00185_));
 sg13g2_nand2b_2 _11043_ (.Y(_04057_),
    .B(_03789_),
    .A_N(_00143_));
 sg13g2_nand2b_2 _11044_ (.Y(_04058_),
    .B(_03868_),
    .A_N(_00149_));
 sg13g2_nor3_1 _11045_ (.A(_00169_),
    .B(net3780),
    .C(net3763),
    .Y(_04059_));
 sg13g2_nand2b_2 _11046_ (.Y(_04060_),
    .B(_03833_),
    .A_N(_00192_));
 sg13g2_nor3_1 _11047_ (.A(_00164_),
    .B(_03739_),
    .C(net3763),
    .Y(_04061_));
 sg13g2_nand2b_2 _11048_ (.Y(_04062_),
    .B(_03882_),
    .A_N(_00155_));
 sg13g2_nand2b_1 _11049_ (.Y(_04063_),
    .B(_03851_),
    .A_N(_00151_));
 sg13g2_nor3_1 _11050_ (.A(_00165_),
    .B(net3779),
    .C(net3763),
    .Y(_04064_));
 sg13g2_nand2b_1 _11051_ (.Y(_04065_),
    .B(_03863_),
    .A_N(_00197_));
 sg13g2_nand2b_2 _11052_ (.Y(_04066_),
    .B(_03884_),
    .A_N(_00153_));
 sg13g2_nor2_1 _11053_ (.A(_00209_),
    .B(_03871_),
    .Y(_04067_));
 sg13g2_nand2b_2 _11054_ (.Y(_04068_),
    .B(_03783_),
    .A_N(_00195_));
 sg13g2_nand2b_2 _11055_ (.Y(_04069_),
    .B(_03786_),
    .A_N(_00191_));
 sg13g2_nand2b_2 _11056_ (.Y(_04070_),
    .B(_03764_),
    .A_N(_00183_));
 sg13g2_nand2b_2 _11057_ (.Y(_04071_),
    .B(_03852_),
    .A_N(_00203_));
 sg13g2_o21ai_1 _11058_ (.B1(_04071_),
    .Y(_04072_),
    .A1(_00172_),
    .A2(_03891_));
 sg13g2_o21ai_1 _11059_ (.B1(_04048_),
    .Y(_04073_),
    .A1(_00194_),
    .A2(_03850_));
 sg13g2_o21ai_1 _11060_ (.B1(_04063_),
    .Y(_04074_),
    .A1(_00193_),
    .A2(_03873_));
 sg13g2_o21ai_1 _11061_ (.B1(_04057_),
    .Y(_04075_),
    .A1(_00178_),
    .A2(_03837_));
 sg13g2_o21ai_1 _11062_ (.B1(_04065_),
    .Y(_04076_),
    .A1(_00186_),
    .A2(_03841_));
 sg13g2_a22oi_1 _11063_ (.Y(_04077_),
    .B1(_03781_),
    .B2(_03529_),
    .A2(_03760_),
    .A1(_03532_));
 sg13g2_a22oi_1 _11064_ (.Y(_04078_),
    .B1(_03802_),
    .B2(_03525_),
    .A2(_03780_),
    .A1(\spiking_network_top_uut.all_data_out[222] ));
 sg13g2_o21ai_1 _11065_ (.B1(_04049_),
    .Y(_04079_),
    .A1(_00180_),
    .A2(_03809_));
 sg13g2_a22oi_1 _11066_ (.Y(_04080_),
    .B1(_03887_),
    .B2(_03514_),
    .A2(_03830_),
    .A1(\spiking_network_top_uut.all_data_out[198] ));
 sg13g2_a22oi_1 _11067_ (.Y(_04081_),
    .B1(_03779_),
    .B2(\spiking_network_top_uut.all_data_out[14] ),
    .A2(net3719),
    .A1(\spiking_network_top_uut.all_data_out[30] ));
 sg13g2_a22oi_1 _11068_ (.Y(_04082_),
    .B1(_03876_),
    .B2(\spiking_network_top_uut.all_data_out[286] ),
    .A2(net3718),
    .A1(\spiking_network_top_uut.all_data_out[62] ));
 sg13g2_a22oi_1 _11069_ (.Y(_04083_),
    .B1(_03848_),
    .B2(_03510_),
    .A2(_03838_),
    .A1(_03512_));
 sg13g2_a22oi_1 _11070_ (.Y(_04084_),
    .B1(_03807_),
    .B2(_03517_),
    .A2(_03782_),
    .A1(\spiking_network_top_uut.all_data_out[142] ));
 sg13g2_a22oi_1 _11071_ (.Y(_04085_),
    .B1(_03835_),
    .B2(_03527_),
    .A2(_03715_),
    .A1(\spiking_network_top_uut.all_data_out[46] ));
 sg13g2_a22oi_1 _11072_ (.Y(_04086_),
    .B1(_03798_),
    .B2(_03521_),
    .A2(net3715),
    .A1(_03543_));
 sg13g2_a22oi_1 _11073_ (.Y(_04087_),
    .B1(_03845_),
    .B2(_03519_),
    .A2(_03776_),
    .A1(\spiking_network_top_uut.all_data_out[174] ));
 sg13g2_nand4_1 _11074_ (.B(_04084_),
    .C(_04086_),
    .A(_04080_),
    .Y(_04088_),
    .D(_04087_));
 sg13g2_a22oi_1 _11075_ (.Y(_04089_),
    .B1(_03788_),
    .B2(\spiking_network_top_uut.all_data_out[158] ),
    .A2(net3695),
    .A1(\spiking_network_top_uut.all_data_out[94] ));
 sg13g2_a22oi_1 _11076_ (.Y(_04090_),
    .B1(net3710),
    .B2(\spiking_network_top_uut.all_data_out[54] ),
    .A2(net3714),
    .A1(\spiking_network_top_uut.all_data_out[102] ));
 sg13g2_a22oi_1 _11077_ (.Y(_04091_),
    .B1(_03820_),
    .B2(\spiking_network_top_uut.all_data_out[166] ),
    .A2(net3694),
    .A1(\spiking_network_top_uut.all_data_out[86] ));
 sg13g2_a22oi_1 _11078_ (.Y(_04092_),
    .B1(_03869_),
    .B2(_03546_),
    .A2(_03772_),
    .A1(_03544_));
 sg13g2_nand4_1 _11079_ (.B(_04090_),
    .C(_04091_),
    .A(_04089_),
    .Y(_04093_),
    .D(_04092_));
 sg13g2_a22oi_1 _11080_ (.Y(_04094_),
    .B1(_03883_),
    .B2(_03526_),
    .A2(net3717),
    .A1(\spiking_network_top_uut.all_data_out[110] ));
 sg13g2_nand4_1 _11081_ (.B(_04052_),
    .C(_04081_),
    .A(_04051_),
    .Y(_04095_),
    .D(_04094_));
 sg13g2_a221oi_1 _11082_ (.B2(\spiking_network_top_uut.all_data_out[214] ),
    .C1(_04095_),
    .B1(_03879_),
    .A1(\spiking_network_top_uut.all_data_out[230] ),
    .Y(_04096_),
    .A2(_03828_));
 sg13g2_a22oi_1 _11083_ (.Y(_04097_),
    .B1(_03821_),
    .B2(\spiking_network_top_uut.all_data_out[310] ),
    .A2(_03795_),
    .A1(\spiking_network_top_uut.all_data_out[270] ));
 sg13g2_a221oi_1 _11084_ (.B2(_03537_),
    .C1(_04079_),
    .B1(_03804_),
    .A1(\spiking_network_top_uut.all_data_out[206] ),
    .Y(_04098_),
    .A2(_03801_));
 sg13g2_nand4_1 _11085_ (.B(_04096_),
    .C(_04097_),
    .A(_04082_),
    .Y(_04099_),
    .D(_04098_));
 sg13g2_a22oi_1 _11086_ (.Y(_04100_),
    .B1(_03861_),
    .B2(_03516_),
    .A2(_03816_),
    .A1(\spiking_network_top_uut.all_data_out[278] ));
 sg13g2_a22oi_1 _11087_ (.Y(_04101_),
    .B1(_03859_),
    .B2(_03524_),
    .A2(_03744_),
    .A1(\spiking_network_top_uut.all_data_out[902] ));
 sg13g2_nand4_1 _11088_ (.B(_04068_),
    .C(_04100_),
    .A(_04060_),
    .Y(_04102_),
    .D(_04101_));
 sg13g2_a221oi_1 _11089_ (.B2(\spiking_network_top_uut.all_data_out[294] ),
    .C1(_04102_),
    .B1(_03819_),
    .A1(_03533_),
    .Y(_04103_),
    .A2(_03784_));
 sg13g2_a22oi_1 _11090_ (.Y(_04104_),
    .B1(_03813_),
    .B2(_03522_),
    .A2(net3713),
    .A1(\spiking_network_top_uut.all_data_out[118] ));
 sg13g2_a22oi_1 _11091_ (.Y(_04105_),
    .B1(_03877_),
    .B2(\spiking_network_top_uut.all_data_out[150] ),
    .A2(_03763_),
    .A1(\spiking_network_top_uut.all_data_out[190] ));
 sg13g2_a22oi_1 _11092_ (.Y(_04106_),
    .B1(net3693),
    .B2(\spiking_network_top_uut.all_data_out[78] ),
    .A2(net3696),
    .A1(\spiking_network_top_uut.all_data_out[70] ));
 sg13g2_nand3_1 _11093_ (.B(_04105_),
    .C(_04106_),
    .A(_04104_),
    .Y(_04107_));
 sg13g2_a221oi_1 _11094_ (.B2(_03518_),
    .C1(_04107_),
    .B1(_03853_),
    .A1(\spiking_network_top_uut.all_data_out[182] ),
    .Y(_04108_),
    .A2(_03803_));
 sg13g2_nand3_1 _11095_ (.B(_04103_),
    .C(_04108_),
    .A(_03757_),
    .Y(_04109_));
 sg13g2_nor4_2 _11096_ (.A(_04088_),
    .B(_04093_),
    .C(_04099_),
    .Y(_04110_),
    .D(_04109_));
 sg13g2_nor4_2 _11097_ (.A(_04059_),
    .B(_04061_),
    .C(_04064_),
    .Y(_04111_),
    .D(_04067_));
 sg13g2_nand4_1 _11098_ (.B(_04066_),
    .C(_04085_),
    .A(_04062_),
    .Y(_04112_),
    .D(_04111_));
 sg13g2_o21ai_1 _11099_ (.B1(_04043_),
    .Y(_04113_),
    .A1(_00196_),
    .A2(_03823_));
 sg13g2_o21ai_1 _11100_ (.B1(_04047_),
    .Y(_04114_),
    .A1(_00141_),
    .A2(_03791_));
 sg13g2_o21ai_1 _11101_ (.B1(_04044_),
    .Y(_04115_),
    .A1(_00189_),
    .A2(_03797_));
 sg13g2_o21ai_1 _11102_ (.B1(_04054_),
    .Y(_04116_),
    .A1(_00175_),
    .A2(_03857_));
 sg13g2_nor4_2 _11103_ (.A(_04113_),
    .B(_04114_),
    .C(_04115_),
    .Y(_04117_),
    .D(_04116_));
 sg13g2_o21ai_1 _11104_ (.B1(_04046_),
    .Y(_04118_),
    .A1(_00171_),
    .A2(_03768_));
 sg13g2_o21ai_1 _11105_ (.B1(_04056_),
    .Y(_04119_),
    .A1(_00187_),
    .A2(_03865_));
 sg13g2_nor4_1 _11106_ (.A(_04075_),
    .B(_04076_),
    .C(_04118_),
    .D(_04119_),
    .Y(_04120_));
 sg13g2_a22oi_1 _11107_ (.Y(_04121_),
    .B1(_03805_),
    .B2(\spiking_network_top_uut.all_data_out[134] ),
    .A2(_03792_),
    .A1(\spiking_network_top_uut.all_data_out[238] ));
 sg13g2_a22oi_1 _11108_ (.Y(_04122_),
    .B1(_03817_),
    .B2(_03535_),
    .A2(net3709),
    .A1(\spiking_network_top_uut.all_data_out[22] ));
 sg13g2_nand4_1 _11109_ (.B(_04070_),
    .C(_04121_),
    .A(_04069_),
    .Y(_04123_),
    .D(_04122_));
 sg13g2_a221oi_1 _11110_ (.B2(_03536_),
    .C1(_04123_),
    .B1(_03880_),
    .A1(\spiking_network_top_uut.all_data_out[262] ),
    .Y(_04124_),
    .A2(_03806_));
 sg13g2_nand3_1 _11111_ (.B(_04120_),
    .C(_04124_),
    .A(_04117_),
    .Y(_04125_));
 sg13g2_a22oi_1 _11112_ (.Y(_04126_),
    .B1(_03878_),
    .B2(_03509_),
    .A2(_03847_),
    .A1(_03541_));
 sg13g2_nand4_1 _11113_ (.B(_04078_),
    .C(_04083_),
    .A(_04077_),
    .Y(_04127_),
    .D(_04126_));
 sg13g2_a22oi_1 _11114_ (.Y(_04128_),
    .B1(_03866_),
    .B2(\spiking_network_top_uut.all_data_out[302] ),
    .A2(_03846_),
    .A1(\spiking_network_top_uut.all_data_out[342] ));
 sg13g2_a22oi_1 _11115_ (.Y(_04129_),
    .B1(_03889_),
    .B2(_03534_),
    .A2(net3712),
    .A1(\spiking_network_top_uut.all_data_out[126] ));
 sg13g2_a22oi_1 _11116_ (.Y(_04130_),
    .B1(_03867_),
    .B2(\spiking_network_top_uut.all_data_out[318] ),
    .A2(_03785_),
    .A1(\spiking_network_top_uut.all_data_out[254] ));
 sg13g2_nand3_1 _11117_ (.B(_04129_),
    .C(_04130_),
    .A(_04128_),
    .Y(_04131_));
 sg13g2_a221oi_1 _11118_ (.B2(\spiking_network_top_uut.all_data_out[334] ),
    .C1(_04131_),
    .B1(_03855_),
    .A1(_03547_),
    .Y(_04132_),
    .A2(_03831_));
 sg13g2_o21ai_1 _11119_ (.B1(_04058_),
    .Y(_04133_),
    .A1(_00201_),
    .A2(_03778_));
 sg13g2_o21ai_1 _11120_ (.B1(_04055_),
    .Y(_04134_),
    .A1(_00188_),
    .A2(_03886_));
 sg13g2_nor4_1 _11121_ (.A(_04072_),
    .B(_04074_),
    .C(_04133_),
    .D(_04134_),
    .Y(_04135_));
 sg13g2_a22oi_1 _11122_ (.Y(_04136_),
    .B1(_03812_),
    .B2(\spiking_network_top_uut.all_data_out[246] ),
    .A2(_03732_),
    .A1(\spiking_network_top_uut.all_data_out[38] ));
 sg13g2_o21ai_1 _11123_ (.B1(_04053_),
    .Y(_04137_),
    .A1(_00147_),
    .A2(_03875_));
 sg13g2_nor4_1 _11124_ (.A(_04045_),
    .B(_04050_),
    .C(_04073_),
    .D(_04137_),
    .Y(_04138_));
 sg13g2_nand4_1 _11125_ (.B(_04135_),
    .C(_04136_),
    .A(_04132_),
    .Y(_04139_),
    .D(_04138_));
 sg13g2_nor4_2 _11126_ (.A(_04112_),
    .B(_04125_),
    .C(_04127_),
    .Y(_04140_),
    .D(_04139_));
 sg13g2_o21ai_1 _11127_ (.B1(\spiking_network_top_uut.spi_inst.spi_slave_inst.bit_cnt[0] ),
    .Y(_04141_),
    .A1(\spiking_network_top_uut.all_data_out[6] ),
    .A2(_03757_));
 sg13g2_a21oi_1 _11128_ (.A1(_04110_),
    .A2(_04140_),
    .Y(_04142_),
    .B1(_04141_));
 sg13g2_nor3_1 _11129_ (.A(\spiking_network_top_uut.spi_inst.spi_slave_inst.bit_cnt[2] ),
    .B(_04042_),
    .C(_04142_),
    .Y(_04143_));
 sg13g2_a22oi_1 _11130_ (.Y(_04144_),
    .B1(_03851_),
    .B2(\spiking_network_top_uut.all_data_out[811] ),
    .A2(_03838_),
    .A1(\spiking_network_top_uut.all_data_out[787] ));
 sg13g2_a22oi_1 _11131_ (.Y(_04145_),
    .B1(_03792_),
    .B2(\spiking_network_top_uut.all_data_out[235] ),
    .A2(net3695),
    .A1(\spiking_network_top_uut.all_data_out[91] ));
 sg13g2_a22oi_1 _11132_ (.Y(_04146_),
    .B1(_03816_),
    .B2(\spiking_network_top_uut.all_data_out[275] ),
    .A2(net3713),
    .A1(\spiking_network_top_uut.all_data_out[115] ));
 sg13g2_a22oi_1 _11133_ (.Y(_04147_),
    .B1(_03849_),
    .B2(\spiking_network_top_uut.all_data_out[467] ),
    .A2(_03846_),
    .A1(\spiking_network_top_uut.all_data_out[339] ));
 sg13g2_a22oi_1 _11134_ (.Y(_04148_),
    .B1(_03867_),
    .B2(\spiking_network_top_uut.all_data_out[315] ),
    .A2(_03866_),
    .A1(\spiking_network_top_uut.all_data_out[299] ));
 sg13g2_a22oi_1 _11135_ (.Y(_04149_),
    .B1(_03821_),
    .B2(\spiking_network_top_uut.all_data_out[307] ),
    .A2(_03795_),
    .A1(\spiking_network_top_uut.all_data_out[267] ));
 sg13g2_a22oi_1 _11136_ (.Y(_04150_),
    .B1(_03813_),
    .B2(\spiking_network_top_uut.all_data_out[723] ),
    .A2(_03798_),
    .A1(\spiking_network_top_uut.all_data_out[731] ));
 sg13g2_a22oi_1 _11137_ (.Y(_04151_),
    .B1(_03853_),
    .B2(\spiking_network_top_uut.all_data_out[747] ),
    .A2(_03788_),
    .A1(\spiking_network_top_uut.all_data_out[155] ));
 sg13g2_a22oi_1 _11138_ (.Y(_04152_),
    .B1(_03887_),
    .B2(\spiking_network_top_uut.all_data_out[771] ),
    .A2(_03820_),
    .A1(\spiking_network_top_uut.all_data_out[163] ));
 sg13g2_a22oi_1 _11139_ (.Y(_04153_),
    .B1(_03811_),
    .B2(\spiking_network_top_uut.all_data_out[371] ),
    .A2(_03767_),
    .A1(\spiking_network_top_uut.all_data_out[651] ));
 sg13g2_a22oi_1 _11140_ (.Y(_04154_),
    .B1(_03834_),
    .B2(\spiking_network_top_uut.all_data_out[707] ),
    .A2(_03772_),
    .A1(\spiking_network_top_uut.all_data_out[379] ));
 sg13g2_a22oi_1 _11141_ (.Y(_04155_),
    .B1(_03862_),
    .B2(\spiking_network_top_uut.all_data_out[699] ),
    .A2(_03782_),
    .A1(\spiking_network_top_uut.all_data_out[139] ));
 sg13g2_nand4_1 _11142_ (.B(_04152_),
    .C(_04154_),
    .A(_04151_),
    .Y(_04156_),
    .D(_04155_));
 sg13g2_a22oi_1 _11143_ (.Y(_04157_),
    .B1(_03801_),
    .B2(\spiking_network_top_uut.all_data_out[203] ),
    .A2(net3709),
    .A1(net4298));
 sg13g2_a22oi_1 _11144_ (.Y(_04158_),
    .B1(_03789_),
    .B2(\spiking_network_top_uut.all_data_out[875] ),
    .A2(_03764_),
    .A1(\spiking_network_top_uut.all_data_out[555] ));
 sg13g2_a22oi_1 _11145_ (.Y(_04159_),
    .B1(_03859_),
    .B2(\spiking_network_top_uut.all_data_out[715] ),
    .A2(_03803_),
    .A1(\spiking_network_top_uut.all_data_out[179] ));
 sg13g2_a22oi_1 _11146_ (.Y(_04160_),
    .B1(_03832_),
    .B2(\spiking_network_top_uut.all_data_out[883] ),
    .A2(_03829_),
    .A1(\spiking_network_top_uut.all_data_out[675] ));
 sg13g2_nand4_1 _11147_ (.B(_04158_),
    .C(_04159_),
    .A(_04157_),
    .Y(_04161_),
    .D(_04160_));
 sg13g2_a22oi_1 _11148_ (.Y(_04162_),
    .B1(_03802_),
    .B2(\spiking_network_top_uut.all_data_out[691] ),
    .A2(net3718),
    .A1(\spiking_network_top_uut.all_data_out[59] ));
 sg13g2_a22oi_1 _11149_ (.Y(_04163_),
    .B1(_03831_),
    .B2(\spiking_network_top_uut.all_data_out[323] ),
    .A2(_03812_),
    .A1(\spiking_network_top_uut.all_data_out[243] ));
 sg13g2_a22oi_1 _11150_ (.Y(_04164_),
    .B1(_03879_),
    .B2(\spiking_network_top_uut.all_data_out[211] ),
    .A2(_03779_),
    .A1(net4275));
 sg13g2_a22oi_1 _11151_ (.Y(_04165_),
    .B1(_03830_),
    .B2(\spiking_network_top_uut.all_data_out[195] ),
    .A2(_03763_),
    .A1(\spiking_network_top_uut.all_data_out[187] ));
 sg13g2_nand4_1 _11152_ (.B(_04163_),
    .C(_04164_),
    .A(_04162_),
    .Y(_04166_),
    .D(_04165_));
 sg13g2_a22oi_1 _11153_ (.Y(_04167_),
    .B1(_03870_),
    .B2(\spiking_network_top_uut.all_data_out[347] ),
    .A2(_03835_),
    .A1(\spiking_network_top_uut.all_data_out[659] ));
 sg13g2_a22oi_1 _11154_ (.Y(_04168_),
    .B1(_03808_),
    .B2(\spiking_network_top_uut.all_data_out[579] ),
    .A2(_03769_),
    .A1(\spiking_network_top_uut.all_data_out[667] ));
 sg13g2_a22oi_1 _11155_ (.Y(_04169_),
    .B1(net3696),
    .B2(\spiking_network_top_uut.all_data_out[67] ),
    .A2(net3710),
    .A1(\spiking_network_top_uut.all_data_out[51] ));
 sg13g2_a22oi_1 _11156_ (.Y(_04170_),
    .B1(_03840_),
    .B2(\spiking_network_top_uut.all_data_out[531] ),
    .A2(_03833_),
    .A1(\spiking_network_top_uut.all_data_out[483] ));
 sg13g2_nand4_1 _11157_ (.B(_04168_),
    .C(_04169_),
    .A(_04167_),
    .Y(_04171_),
    .D(_04170_));
 sg13g2_or4_1 _11158_ (.A(_04156_),
    .B(_04161_),
    .C(_04166_),
    .D(_04171_),
    .X(_04172_));
 sg13g2_a22oi_1 _11159_ (.Y(_04173_),
    .B1(_03876_),
    .B2(\spiking_network_top_uut.all_data_out[283] ),
    .A2(_03856_),
    .A1(\spiking_network_top_uut.all_data_out[619] ));
 sg13g2_a22oi_1 _11160_ (.Y(_04174_),
    .B1(_03814_),
    .B2(\spiking_network_top_uut.all_data_out[627] ),
    .A2(_03807_),
    .A1(\spiking_network_top_uut.all_data_out[755] ));
 sg13g2_a22oi_1 _11161_ (.Y(_04175_),
    .B1(_03890_),
    .B2(\spiking_network_top_uut.all_data_out[643] ),
    .A2(_03847_),
    .A1(\spiking_network_top_uut.all_data_out[403] ));
 sg13g2_a22oi_1 _11162_ (.Y(_04176_),
    .B1(_03883_),
    .B2(\spiking_network_top_uut.all_data_out[683] ),
    .A2(_03824_),
    .A1(\spiking_network_top_uut.all_data_out[419] ));
 sg13g2_nand4_1 _11163_ (.B(_04174_),
    .C(_04175_),
    .A(_04173_),
    .Y(_04177_),
    .D(_04176_));
 sg13g2_a22oi_1 _11164_ (.Y(_04178_),
    .B1(_03861_),
    .B2(\spiking_network_top_uut.all_data_out[763] ),
    .A2(_03776_),
    .A1(\spiking_network_top_uut.all_data_out[171] ));
 sg13g2_a22oi_1 _11165_ (.Y(_04179_),
    .B1(net3693),
    .B2(\spiking_network_top_uut.all_data_out[75] ),
    .A2(net3715),
    .A1(\spiking_network_top_uut.all_data_out[387] ));
 sg13g2_a22oi_1 _11166_ (.Y(_04180_),
    .B1(_03877_),
    .B2(\spiking_network_top_uut.all_data_out[147] ),
    .A2(_03806_),
    .A1(\spiking_network_top_uut.all_data_out[259] ));
 sg13g2_a22oi_1 _11167_ (.Y(_04181_),
    .B1(_03805_),
    .B2(\spiking_network_top_uut.all_data_out[131] ),
    .A2(net3712),
    .A1(\spiking_network_top_uut.all_data_out[123] ));
 sg13g2_nand4_1 _11168_ (.B(_04179_),
    .C(_04180_),
    .A(_04178_),
    .Y(_04182_),
    .D(_04181_));
 sg13g2_nor4_1 _11169_ (.A(_03756_),
    .B(_04172_),
    .C(_04177_),
    .D(_04182_),
    .Y(_04183_));
 sg13g2_a22oi_1 _11170_ (.Y(_04184_),
    .B1(_03864_),
    .B2(\spiking_network_top_uut.all_data_out[523] ),
    .A2(_03783_),
    .A1(\spiking_network_top_uut.all_data_out[459] ));
 sg13g2_a22oi_1 _11171_ (.Y(_04185_),
    .B1(_03786_),
    .B2(\spiking_network_top_uut.all_data_out[491] ),
    .A2(_03775_),
    .A1(\spiking_network_top_uut.all_data_out[859] ));
 sg13g2_a22oi_1 _11172_ (.Y(_04186_),
    .B1(_03845_),
    .B2(\spiking_network_top_uut.all_data_out[739] ),
    .A2(_03760_),
    .A1(\spiking_network_top_uut.all_data_out[603] ));
 sg13g2_nand4_1 _11173_ (.B(_04184_),
    .C(_04185_),
    .A(_04150_),
    .Y(_04187_),
    .D(_04186_));
 sg13g2_a22oi_1 _11174_ (.Y(_04188_),
    .B1(_03889_),
    .B2(\spiking_network_top_uut.all_data_out[571] ),
    .A2(_03794_),
    .A1(\spiking_network_top_uut.all_data_out[539] ));
 sg13g2_a22oi_1 _11175_ (.Y(_04189_),
    .B1(_03880_),
    .B2(\spiking_network_top_uut.all_data_out[547] ),
    .A2(_03781_),
    .A1(\spiking_network_top_uut.all_data_out[635] ));
 sg13g2_a22oi_1 _11176_ (.Y(_04190_),
    .B1(_03790_),
    .B2(\spiking_network_top_uut.all_data_out[891] ),
    .A2(net3711),
    .A1(\spiking_network_top_uut.all_data_out[35] ));
 sg13g2_a22oi_1 _11177_ (.Y(_04191_),
    .B1(_03842_),
    .B2(\spiking_network_top_uut.all_data_out[611] ),
    .A2(net3719),
    .A1(\spiking_network_top_uut.all_data_out[27] ));
 sg13g2_nand4_1 _11178_ (.B(_04189_),
    .C(_04190_),
    .A(_04188_),
    .Y(_04192_),
    .D(_04191_));
 sg13g2_a22oi_1 _11179_ (.Y(_04193_),
    .B1(_03878_),
    .B2(\spiking_network_top_uut.all_data_out[867] ),
    .A2(_03796_),
    .A1(\spiking_network_top_uut.all_data_out[507] ));
 sg13g2_a22oi_1 _11180_ (.Y(_04194_),
    .B1(_03874_),
    .B2(\spiking_network_top_uut.all_data_out[843] ),
    .A2(_03810_),
    .A1(\spiking_network_top_uut.all_data_out[851] ));
 sg13g2_a22oi_1 _11181_ (.Y(_04195_),
    .B1(_03836_),
    .B2(\spiking_network_top_uut.all_data_out[595] ),
    .A2(_03784_),
    .A1(\spiking_network_top_uut.all_data_out[587] ));
 sg13g2_a22oi_1 _11182_ (.Y(_04196_),
    .B1(_03817_),
    .B2(\spiking_network_top_uut.all_data_out[563] ),
    .A2(_03804_),
    .A1(\spiking_network_top_uut.all_data_out[499] ));
 sg13g2_nand4_1 _11183_ (.B(_04194_),
    .C(_04195_),
    .A(_04193_),
    .Y(_04197_),
    .D(_04196_));
 sg13g2_a22oi_1 _11184_ (.Y(_04198_),
    .B1(_03855_),
    .B2(\spiking_network_top_uut.all_data_out[331] ),
    .A2(_03844_),
    .A1(\spiking_network_top_uut.all_data_out[355] ));
 sg13g2_nand4_1 _11185_ (.B(_04148_),
    .C(_04153_),
    .A(_04147_),
    .Y(_04199_),
    .D(_04198_));
 sg13g2_nor4_2 _11186_ (.A(_04187_),
    .B(_04192_),
    .C(_04197_),
    .Y(_04200_),
    .D(_04199_));
 sg13g2_a22oi_1 _11187_ (.Y(_04201_),
    .B1(net3714),
    .B2(\spiking_network_top_uut.all_data_out[99] ),
    .A2(_03713_),
    .A1(\spiking_network_top_uut.all_data_out[107] ));
 sg13g2_a22oi_1 _11188_ (.Y(_04202_),
    .B1(_03785_),
    .B2(\spiking_network_top_uut.all_data_out[251] ),
    .A2(net3694),
    .A1(\spiking_network_top_uut.all_data_out[83] ));
 sg13g2_a22oi_1 _11189_ (.Y(_04203_),
    .B1(_03869_),
    .B2(\spiking_network_top_uut.all_data_out[363] ),
    .A2(_03819_),
    .A1(\spiking_network_top_uut.all_data_out[291] ));
 sg13g2_nand4_1 _11190_ (.B(_04201_),
    .C(_04202_),
    .A(_04145_),
    .Y(_04204_),
    .D(_04203_));
 sg13g2_a22oi_1 _11191_ (.Y(_04205_),
    .B1(_03872_),
    .B2(\spiking_network_top_uut.all_data_out[475] ),
    .A2(_03780_),
    .A1(\spiking_network_top_uut.all_data_out[219] ));
 sg13g2_a22oi_1 _11192_ (.Y(_04206_),
    .B1(_03828_),
    .B2(\spiking_network_top_uut.all_data_out[227] ),
    .A2(net3716),
    .A1(\spiking_network_top_uut.all_data_out[43] ));
 sg13g2_nand4_1 _11193_ (.B(_04149_),
    .C(_04205_),
    .A(_04146_),
    .Y(_04207_),
    .D(_04206_));
 sg13g2_a22oi_1 _11194_ (.Y(_04208_),
    .B1(_03885_),
    .B2(\spiking_network_top_uut.all_data_out[515] ),
    .A2(_03884_),
    .A1(\spiking_network_top_uut.all_data_out[795] ));
 sg13g2_a22oi_1 _11195_ (.Y(_04209_),
    .B1(_03848_),
    .B2(\spiking_network_top_uut.all_data_out[819] ),
    .A2(_03744_),
    .A1(\spiking_network_top_uut.all_data_out[899] ));
 sg13g2_a22oi_1 _11196_ (.Y(_04210_),
    .B1(_03882_),
    .B2(\spiking_network_top_uut.all_data_out[779] ),
    .A2(_03843_),
    .A1(\spiking_network_top_uut.all_data_out[435] ));
 sg13g2_a22oi_1 _11197_ (.Y(_04211_),
    .B1(_03839_),
    .B2(\spiking_network_top_uut.all_data_out[803] ),
    .A2(_03777_),
    .A1(\spiking_network_top_uut.all_data_out[411] ));
 sg13g2_nand4_1 _11198_ (.B(_04209_),
    .C(_04210_),
    .A(_04208_),
    .Y(_04212_),
    .D(_04211_));
 sg13g2_a22oi_1 _11199_ (.Y(_04213_),
    .B1(_03868_),
    .B2(\spiking_network_top_uut.all_data_out[827] ),
    .A2(_03826_),
    .A1(\spiking_network_top_uut.all_data_out[835] ));
 sg13g2_a22oi_1 _11200_ (.Y(_04214_),
    .B1(_03863_),
    .B2(\spiking_network_top_uut.all_data_out[443] ),
    .A2(_03822_),
    .A1(\spiking_network_top_uut.all_data_out[451] ));
 sg13g2_a22oi_1 _11201_ (.Y(_04215_),
    .B1(_03852_),
    .B2(\spiking_network_top_uut.all_data_out[395] ),
    .A2(_03799_),
    .A1(\spiking_network_top_uut.all_data_out[427] ));
 sg13g2_nand4_1 _11202_ (.B(_04213_),
    .C(_04214_),
    .A(_04144_),
    .Y(_04216_),
    .D(_04215_));
 sg13g2_nor4_1 _11203_ (.A(_04204_),
    .B(_04207_),
    .C(_04212_),
    .D(_04216_),
    .Y(_04217_));
 sg13g2_nand3_1 _11204_ (.B(_04200_),
    .C(_04217_),
    .A(_04183_),
    .Y(_04218_));
 sg13g2_o21ai_1 _11205_ (.B1(_04218_),
    .Y(_04219_),
    .A1(\spiking_network_top_uut.all_data_out[3] ),
    .A2(_03757_));
 sg13g2_nand2b_2 _11206_ (.Y(_04220_),
    .B(_03849_),
    .A_N(_00334_));
 sg13g2_nand2b_2 _11207_ (.Y(_04221_),
    .B(_03807_),
    .A_N(_00298_));
 sg13g2_nand2b_2 _11208_ (.Y(_04222_),
    .B(_03843_),
    .A_N(_00338_));
 sg13g2_nand2b_2 _11209_ (.Y(_04223_),
    .B(_03845_),
    .A_N(_00300_));
 sg13g2_nand2b_1 _11210_ (.Y(_04224_),
    .B(_03851_),
    .A_N(_00291_));
 sg13g2_nand2b_1 _11211_ (.Y(_04225_),
    .B(_03853_),
    .A_N(_00299_));
 sg13g2_nand2b_1 _11212_ (.Y(_04226_),
    .B(_03852_),
    .A_N(_00343_));
 sg13g2_nand2b_1 _11213_ (.Y(_04227_),
    .B(_03789_),
    .A_N(_00283_));
 sg13g2_nand2b_2 _11214_ (.Y(_04228_),
    .B(_03884_),
    .A_N(_00293_));
 sg13g2_nand2b_2 _11215_ (.Y(_04229_),
    .B(_03878_),
    .A_N(_00284_));
 sg13g2_nand2b_2 _11216_ (.Y(_04230_),
    .B(_03824_),
    .A_N(_00340_));
 sg13g2_nand2b_2 _11217_ (.Y(_04231_),
    .B(_03784_),
    .A_N(_00319_));
 sg13g2_nand2b_1 _11218_ (.Y(_04232_),
    .B(_03856_),
    .A_N(_00315_));
 sg13g2_nand2b_2 _11219_ (.Y(_04233_),
    .B(_03859_),
    .A_N(_00303_));
 sg13g2_nand2b_2 _11220_ (.Y(_04234_),
    .B(_03769_),
    .A_N(_00309_));
 sg13g2_a22oi_1 _11221_ (.Y(_04235_),
    .B1(_03764_),
    .B2(_03610_),
    .A2(net3717),
    .A1(\spiking_network_top_uut.all_data_out[106] ));
 sg13g2_nand2b_1 _11222_ (.Y(_04236_),
    .B(_03869_),
    .A_N(_00347_));
 sg13g2_nand2b_2 _11223_ (.Y(_04237_),
    .B(_03868_),
    .A_N(_00289_));
 sg13g2_a22oi_1 _11224_ (.Y(_04238_),
    .B1(_03874_),
    .B2(_03582_),
    .A2(_03801_),
    .A1(\spiking_network_top_uut.all_data_out[202] ));
 sg13g2_a22oi_1 _11225_ (.Y(_04239_),
    .B1(_03836_),
    .B2(_03607_),
    .A2(_03779_),
    .A1(net4279));
 sg13g2_a22oi_1 _11226_ (.Y(_04240_),
    .B1(_03794_),
    .B2(_03613_),
    .A2(_03785_),
    .A1(\spiking_network_top_uut.all_data_out[250] ));
 sg13g2_a22oi_1 _11227_ (.Y(_04241_),
    .B1(_03812_),
    .B2(\spiking_network_top_uut.all_data_out[242] ),
    .A2(_03781_),
    .A1(_03604_));
 sg13g2_a22oi_1 _11228_ (.Y(_04242_),
    .B1(net3694),
    .B2(\spiking_network_top_uut.all_data_out[82] ),
    .A2(net3716),
    .A1(\spiking_network_top_uut.all_data_out[42] ));
 sg13g2_o21ai_1 _11229_ (.B1(_04226_),
    .Y(_04243_),
    .A1(_00314_),
    .A2(_03815_));
 sg13g2_a221oi_1 _11230_ (.B2(_03588_),
    .C1(_04243_),
    .B1(_03882_),
    .A1(_03580_),
    .Y(_04244_),
    .A2(_03810_));
 sg13g2_nand4_1 _11231_ (.B(_04236_),
    .C(_04241_),
    .A(_04223_),
    .Y(_04245_),
    .D(_04244_));
 sg13g2_o21ai_1 _11232_ (.B1(_04234_),
    .Y(_04246_),
    .A1(_00349_),
    .A2(_03871_));
 sg13g2_a221oi_1 _11233_ (.B2(_03590_),
    .C1(_04246_),
    .B1(_03861_),
    .A1(\spiking_network_top_uut.all_data_out[50] ),
    .Y(_04247_),
    .A2(_03737_));
 sg13g2_nand4_1 _11234_ (.B(_04230_),
    .C(_04242_),
    .A(_04220_),
    .Y(_04248_),
    .D(_04247_));
 sg13g2_a22oi_1 _11235_ (.Y(_04249_),
    .B1(_03883_),
    .B2(_03597_),
    .A2(_03830_),
    .A1(\spiking_network_top_uut.all_data_out[194] ));
 sg13g2_a22oi_1 _11236_ (.Y(_04250_),
    .B1(_03820_),
    .B2(\spiking_network_top_uut.all_data_out[162] ),
    .A2(_03772_),
    .A1(_03629_));
 sg13g2_a22oi_1 _11237_ (.Y(_04251_),
    .B1(_03813_),
    .B2(_03592_),
    .A2(net3718),
    .A1(\spiking_network_top_uut.all_data_out[58] ));
 sg13g2_nand4_1 _11238_ (.B(_04249_),
    .C(_04250_),
    .A(_04239_),
    .Y(_04252_),
    .D(_04251_));
 sg13g2_a22oi_1 _11239_ (.Y(_04253_),
    .B1(_03828_),
    .B2(\spiking_network_top_uut.all_data_out[226] ),
    .A2(net3693),
    .A1(\spiking_network_top_uut.all_data_out[74] ));
 sg13g2_a22oi_1 _11240_ (.Y(_04254_),
    .B1(_03855_),
    .B2(\spiking_network_top_uut.all_data_out[330] ),
    .A2(_03763_),
    .A1(\spiking_network_top_uut.all_data_out[186] ));
 sg13g2_o21ai_1 _11241_ (.B1(_04227_),
    .Y(_04255_),
    .A1(_00328_),
    .A2(_03886_));
 sg13g2_a221oi_1 _11242_ (.B2(\spiking_network_top_uut.all_data_out[298] ),
    .C1(_04255_),
    .B1(_03866_),
    .A1(_03594_),
    .Y(_04256_),
    .A2(_03862_));
 sg13g2_nand3_1 _11243_ (.B(_04254_),
    .C(_04256_),
    .A(_04253_),
    .Y(_04257_));
 sg13g2_nor4_1 _11244_ (.A(_04245_),
    .B(_04248_),
    .C(_04252_),
    .D(_04257_),
    .Y(_04258_));
 sg13g2_a22oi_1 _11245_ (.Y(_04259_),
    .B1(_03780_),
    .B2(\spiking_network_top_uut.all_data_out[218] ),
    .A2(net3715),
    .A1(_03628_));
 sg13g2_a22oi_1 _11246_ (.Y(_04260_),
    .B1(_03846_),
    .B2(\spiking_network_top_uut.all_data_out[338] ),
    .A2(_03790_),
    .A1(_03576_));
 sg13g2_a22oi_1 _11247_ (.Y(_04261_),
    .B1(_03890_),
    .B2(_03602_),
    .A2(_03833_),
    .A1(_03619_));
 sg13g2_a22oi_1 _11248_ (.Y(_04262_),
    .B1(_03838_),
    .B2(_03587_),
    .A2(_03777_),
    .A1(_03626_));
 sg13g2_nand4_1 _11249_ (.B(_04260_),
    .C(_04261_),
    .A(_04259_),
    .Y(_04263_),
    .D(_04262_));
 sg13g2_a22oi_1 _11250_ (.Y(_04264_),
    .B1(_03842_),
    .B2(_03605_),
    .A2(_03798_),
    .A1(_03591_));
 sg13g2_a22oi_1 _11251_ (.Y(_04265_),
    .B1(_03808_),
    .B2(_03608_),
    .A2(_03760_),
    .A1(_03606_));
 sg13g2_a22oi_1 _11252_ (.Y(_04266_),
    .B1(_03804_),
    .B2(_03616_),
    .A2(_03788_),
    .A1(\spiking_network_top_uut.all_data_out[154] ));
 sg13g2_a22oi_1 _11253_ (.Y(_04267_),
    .B1(_03872_),
    .B2(_03620_),
    .A2(_03831_),
    .A1(_03632_));
 sg13g2_nand4_1 _11254_ (.B(_04265_),
    .C(_04266_),
    .A(_04264_),
    .Y(_04268_),
    .D(_04267_));
 sg13g2_nor2_1 _11255_ (.A(_04263_),
    .B(_04268_),
    .Y(_04269_));
 sg13g2_a22oi_1 _11256_ (.Y(_04270_),
    .B1(_03821_),
    .B2(\spiking_network_top_uut.all_data_out[306] ),
    .A2(_03806_),
    .A1(\spiking_network_top_uut.all_data_out[258] ));
 sg13g2_o21ai_1 _11257_ (.B1(_04232_),
    .Y(_04271_),
    .A1(_00336_),
    .A2(_03823_));
 sg13g2_a221oi_1 _11258_ (.B2(\spiking_network_top_uut.all_data_out[146] ),
    .C1(_04271_),
    .B1(_03877_),
    .A1(\spiking_network_top_uut.all_data_out[266] ),
    .Y(_04272_),
    .A2(_03795_));
 sg13g2_nand4_1 _11259_ (.B(_04233_),
    .C(_04270_),
    .A(_04222_),
    .Y(_04273_),
    .D(_04272_));
 sg13g2_a22oi_1 _11260_ (.Y(_04274_),
    .B1(_03832_),
    .B2(_03578_),
    .A2(_03783_),
    .A1(_03622_));
 sg13g2_a22oi_1 _11261_ (.Y(_04275_),
    .B1(_03887_),
    .B2(_03589_),
    .A2(_03799_),
    .A1(_03625_));
 sg13g2_a22oi_1 _11262_ (.Y(_04276_),
    .B1(_03803_),
    .B2(\spiking_network_top_uut.all_data_out[178] ),
    .A2(_03786_),
    .A1(_03618_));
 sg13g2_a22oi_1 _11263_ (.Y(_04277_),
    .B1(_03880_),
    .B2(_03611_),
    .A2(_03805_),
    .A1(\spiking_network_top_uut.all_data_out[130] ));
 sg13g2_nand4_1 _11264_ (.B(_04275_),
    .C(_04276_),
    .A(_04274_),
    .Y(_04278_),
    .D(_04277_));
 sg13g2_a22oi_1 _11265_ (.Y(_04279_),
    .B1(_03848_),
    .B2(_03584_),
    .A2(net3711),
    .A1(\spiking_network_top_uut.all_data_out[34] ));
 sg13g2_a22oi_1 _11266_ (.Y(_04280_),
    .B1(_03867_),
    .B2(\spiking_network_top_uut.all_data_out[314] ),
    .A2(_03816_),
    .A1(\spiking_network_top_uut.all_data_out[274] ));
 sg13g2_a22oi_1 _11267_ (.Y(_04281_),
    .B1(_03863_),
    .B2(_03624_),
    .A2(net3696),
    .A1(\spiking_network_top_uut.all_data_out[66] ));
 sg13g2_nand4_1 _11268_ (.B(_04279_),
    .C(_04280_),
    .A(_04240_),
    .Y(_04282_),
    .D(_04281_));
 sg13g2_a22oi_1 _11269_ (.Y(_04283_),
    .B1(_03864_),
    .B2(_03615_),
    .A2(_03811_),
    .A1(_03630_));
 sg13g2_a22oi_1 _11270_ (.Y(_04284_),
    .B1(_03819_),
    .B2(\spiking_network_top_uut.all_data_out[290] ),
    .A2(_03802_),
    .A1(_03595_));
 sg13g2_a22oi_1 _11271_ (.Y(_04285_),
    .B1(_03835_),
    .B2(_03599_),
    .A2(_03776_),
    .A1(\spiking_network_top_uut.all_data_out[170] ));
 sg13g2_nand4_1 _11272_ (.B(_04283_),
    .C(_04284_),
    .A(_04238_),
    .Y(_04286_),
    .D(_04285_));
 sg13g2_or4_1 _11273_ (.A(_04273_),
    .B(_04278_),
    .C(_04282_),
    .D(_04286_),
    .X(_04287_));
 sg13g2_a22oi_1 _11274_ (.Y(_04288_),
    .B1(_03876_),
    .B2(\spiking_network_top_uut.all_data_out[282] ),
    .A2(_03844_),
    .A1(_03631_));
 sg13g2_o21ai_1 _11275_ (.B1(_04224_),
    .Y(_04289_),
    .A1(_00322_),
    .A2(_03818_));
 sg13g2_a221oi_1 _11276_ (.B2(\spiking_network_top_uut.all_data_out[234] ),
    .C1(_04289_),
    .B1(_03792_),
    .A1(_03601_),
    .Y(_04290_),
    .A2(_03767_));
 sg13g2_nand4_1 _11277_ (.B(_04228_),
    .C(_04288_),
    .A(_04225_),
    .Y(_04291_),
    .D(_04290_));
 sg13g2_a22oi_1 _11278_ (.Y(_04292_),
    .B1(_03879_),
    .B2(\spiking_network_top_uut.all_data_out[210] ),
    .A2(net3712),
    .A1(\spiking_network_top_uut.all_data_out[122] ));
 sg13g2_a22oi_1 _11279_ (.Y(_04293_),
    .B1(_03889_),
    .B2(_03609_),
    .A2(_03782_),
    .A1(\spiking_network_top_uut.all_data_out[138] ));
 sg13g2_o21ai_1 _11280_ (.B1(_04229_),
    .Y(_04294_),
    .A1(_00329_),
    .A2(_03797_));
 sg13g2_a221oi_1 _11281_ (.B2(_03627_),
    .C1(_04294_),
    .B1(_03847_),
    .A1(\spiking_network_top_uut.all_data_out[898] ),
    .Y(_04295_),
    .A2(_03744_));
 sg13g2_nand3_1 _11282_ (.B(_04293_),
    .C(_04295_),
    .A(_04292_),
    .Y(_04296_));
 sg13g2_a22oi_1 _11283_ (.Y(_04297_),
    .B1(_03834_),
    .B2(_03593_),
    .A2(net3695),
    .A1(\spiking_network_top_uut.all_data_out[90] ));
 sg13g2_nand4_1 _11284_ (.B(_04235_),
    .C(_04237_),
    .A(_04231_),
    .Y(_04298_),
    .D(_04297_));
 sg13g2_a221oi_1 _11285_ (.B2(_03598_),
    .C1(_04298_),
    .B1(_03829_),
    .A1(\spiking_network_top_uut.all_data_out[98] ),
    .Y(_04299_),
    .A2(net3714));
 sg13g2_a22oi_1 _11286_ (.Y(_04300_),
    .B1(_03839_),
    .B2(_03586_),
    .A2(net3709),
    .A1(net4305));
 sg13g2_a22oi_1 _11287_ (.Y(_04301_),
    .B1(_03775_),
    .B2(_03579_),
    .A2(net3719),
    .A1(\spiking_network_top_uut.all_data_out[26] ));
 sg13g2_o21ai_1 _11288_ (.B1(_04221_),
    .Y(_04302_),
    .A1(_00288_),
    .A2(_03827_));
 sg13g2_a221oi_1 _11289_ (.B2(_03614_),
    .C1(_04302_),
    .B1(_03840_),
    .A1(\spiking_network_top_uut.all_data_out[114] ),
    .Y(_04303_),
    .A2(net3713));
 sg13g2_nand4_1 _11290_ (.B(_04300_),
    .C(_04301_),
    .A(_04299_),
    .Y(_04304_),
    .D(_04303_));
 sg13g2_nor4_2 _11291_ (.A(_04287_),
    .B(_04291_),
    .C(_04296_),
    .Y(_04305_),
    .D(_04304_));
 sg13g2_nand4_1 _11292_ (.B(_04258_),
    .C(_04269_),
    .A(_03757_),
    .Y(_04306_),
    .D(_04305_));
 sg13g2_a21oi_1 _11293_ (.A1(_03473_),
    .A2(_03756_),
    .Y(_04307_),
    .B1(_03471_));
 sg13g2_o21ai_1 _11294_ (.B1(\spiking_network_top_uut.spi_inst.spi_slave_inst.bit_cnt[2] ),
    .Y(_04308_),
    .A1(\spiking_network_top_uut.spi_inst.spi_slave_inst.bit_cnt[0] ),
    .A2(_04219_));
 sg13g2_a21oi_1 _11295_ (.A1(_04306_),
    .A2(_04307_),
    .Y(_04309_),
    .B1(_04308_));
 sg13g2_nor3_1 _11296_ (.A(\spiking_network_top_uut.spi_inst.spi_slave_inst.bit_cnt[1] ),
    .B(_04143_),
    .C(_04309_),
    .Y(_04310_));
 sg13g2_a22oi_1 _11297_ (.Y(_04311_),
    .B1(_03805_),
    .B2(\spiking_network_top_uut.all_data_out[132] ),
    .A2(_03740_),
    .A1(\spiking_network_top_uut.all_data_out[68] ));
 sg13g2_a22oi_1 _11298_ (.Y(_04312_),
    .B1(_03863_),
    .B2(\spiking_network_top_uut.all_data_out[444] ),
    .A2(_03786_),
    .A1(\spiking_network_top_uut.all_data_out[492] ));
 sg13g2_a22oi_1 _11299_ (.Y(_04313_),
    .B1(_03877_),
    .B2(\spiking_network_top_uut.all_data_out[148] ),
    .A2(_03775_),
    .A1(\spiking_network_top_uut.all_data_out[860] ));
 sg13g2_a22oi_1 _11300_ (.Y(_04314_),
    .B1(_03853_),
    .B2(\spiking_network_top_uut.all_data_out[748] ),
    .A2(_03801_),
    .A1(\spiking_network_top_uut.all_data_out[204] ));
 sg13g2_a22oi_1 _11301_ (.Y(_04315_),
    .B1(_03799_),
    .B2(\spiking_network_top_uut.all_data_out[428] ),
    .A2(net3694),
    .A1(\spiking_network_top_uut.all_data_out[84] ));
 sg13g2_a22oi_1 _11302_ (.Y(_04316_),
    .B1(_03882_),
    .B2(\spiking_network_top_uut.all_data_out[780] ),
    .A2(_03790_),
    .A1(\spiking_network_top_uut.all_data_out[892] ));
 sg13g2_a22oi_1 _11303_ (.Y(_04317_),
    .B1(_03859_),
    .B2(\spiking_network_top_uut.all_data_out[716] ),
    .A2(_03817_),
    .A1(\spiking_network_top_uut.all_data_out[564] ));
 sg13g2_a22oi_1 _11304_ (.Y(_04318_),
    .B1(_03874_),
    .B2(\spiking_network_top_uut.all_data_out[844] ),
    .A2(_03846_),
    .A1(\spiking_network_top_uut.all_data_out[340] ));
 sg13g2_a22oi_1 _11305_ (.Y(_04319_),
    .B1(_03866_),
    .B2(\spiking_network_top_uut.all_data_out[300] ),
    .A2(_03812_),
    .A1(\spiking_network_top_uut.all_data_out[244] ));
 sg13g2_a22oi_1 _11306_ (.Y(_04320_),
    .B1(_03767_),
    .B2(\spiking_network_top_uut.all_data_out[652] ),
    .A2(net3717),
    .A1(\spiking_network_top_uut.all_data_out[108] ));
 sg13g2_a22oi_1 _11307_ (.Y(_04321_),
    .B1(_03789_),
    .B2(\spiking_network_top_uut.all_data_out[876] ),
    .A2(_03744_),
    .A1(\spiking_network_top_uut.all_data_out[900] ));
 sg13g2_a22oi_1 _11308_ (.Y(_04322_),
    .B1(_03829_),
    .B2(\spiking_network_top_uut.all_data_out[676] ),
    .A2(_03819_),
    .A1(\spiking_network_top_uut.all_data_out[292] ));
 sg13g2_a22oi_1 _11309_ (.Y(_04323_),
    .B1(_03816_),
    .B2(\spiking_network_top_uut.all_data_out[276] ),
    .A2(_03808_),
    .A1(\spiking_network_top_uut.all_data_out[580] ));
 sg13g2_a22oi_1 _11310_ (.Y(_04324_),
    .B1(_03840_),
    .B2(\spiking_network_top_uut.all_data_out[532] ),
    .A2(_03830_),
    .A1(\spiking_network_top_uut.all_data_out[196] ));
 sg13g2_nand4_1 _11311_ (.B(_04322_),
    .C(_04323_),
    .A(_04321_),
    .Y(_04325_),
    .D(_04324_));
 sg13g2_a22oi_1 _11312_ (.Y(_04326_),
    .B1(_03889_),
    .B2(\spiking_network_top_uut.all_data_out[572] ),
    .A2(_03776_),
    .A1(\spiking_network_top_uut.all_data_out[172] ));
 sg13g2_a22oi_1 _11313_ (.Y(_04327_),
    .B1(_03832_),
    .B2(\spiking_network_top_uut.all_data_out[884] ),
    .A2(_03796_),
    .A1(\spiking_network_top_uut.all_data_out[508] ));
 sg13g2_a22oi_1 _11314_ (.Y(_04328_),
    .B1(_03769_),
    .B2(\spiking_network_top_uut.all_data_out[668] ),
    .A2(_03742_),
    .A1(\spiking_network_top_uut.all_data_out[20] ));
 sg13g2_a22oi_1 _11315_ (.Y(_04329_),
    .B1(_03872_),
    .B2(\spiking_network_top_uut.all_data_out[476] ),
    .A2(_03764_),
    .A1(\spiking_network_top_uut.all_data_out[556] ));
 sg13g2_nand4_1 _11316_ (.B(_04327_),
    .C(_04328_),
    .A(_04326_),
    .Y(_04330_),
    .D(_04329_));
 sg13g2_a22oi_1 _11317_ (.Y(_04331_),
    .B1(_03870_),
    .B2(\spiking_network_top_uut.all_data_out[348] ),
    .A2(_03780_),
    .A1(\spiking_network_top_uut.all_data_out[220] ));
 sg13g2_a22oi_1 _11318_ (.Y(_04332_),
    .B1(_03828_),
    .B2(\spiking_network_top_uut.all_data_out[228] ),
    .A2(_03807_),
    .A1(\spiking_network_top_uut.all_data_out[756] ));
 sg13g2_a22oi_1 _11319_ (.Y(_04333_),
    .B1(_03868_),
    .B2(\spiking_network_top_uut.all_data_out[828] ),
    .A2(_03802_),
    .A1(\spiking_network_top_uut.all_data_out[692] ));
 sg13g2_a22oi_1 _11320_ (.Y(_04334_),
    .B1(_03890_),
    .B2(\spiking_network_top_uut.all_data_out[644] ),
    .A2(_03836_),
    .A1(\spiking_network_top_uut.all_data_out[596] ));
 sg13g2_nand4_1 _11321_ (.B(_04332_),
    .C(_04333_),
    .A(_04331_),
    .Y(_04335_),
    .D(_04334_));
 sg13g2_a22oi_1 _11322_ (.Y(_04336_),
    .B1(_03876_),
    .B2(\spiking_network_top_uut.all_data_out[284] ),
    .A2(_03798_),
    .A1(\spiking_network_top_uut.all_data_out[732] ));
 sg13g2_a22oi_1 _11323_ (.Y(_04337_),
    .B1(_03842_),
    .B2(\spiking_network_top_uut.all_data_out[612] ),
    .A2(net3710),
    .A1(\spiking_network_top_uut.all_data_out[52] ));
 sg13g2_a22oi_1 _11324_ (.Y(_04338_),
    .B1(_03824_),
    .B2(\spiking_network_top_uut.all_data_out[420] ),
    .A2(net3719),
    .A1(\spiking_network_top_uut.all_data_out[28] ));
 sg13g2_nand4_1 _11325_ (.B(_04336_),
    .C(_04337_),
    .A(_04316_),
    .Y(_04339_),
    .D(_04338_));
 sg13g2_or4_1 _11326_ (.A(_04325_),
    .B(_04330_),
    .C(_04335_),
    .D(_04339_),
    .X(_04340_));
 sg13g2_a22oi_1 _11327_ (.Y(_04341_),
    .B1(_03867_),
    .B2(\spiking_network_top_uut.all_data_out[316] ),
    .A2(_03851_),
    .A1(\spiking_network_top_uut.all_data_out[812] ));
 sg13g2_a22oi_1 _11328_ (.Y(_04342_),
    .B1(_03804_),
    .B2(\spiking_network_top_uut.all_data_out[500] ),
    .A2(_03794_),
    .A1(\spiking_network_top_uut.all_data_out[540] ));
 sg13g2_a22oi_1 _11329_ (.Y(_04343_),
    .B1(_03792_),
    .B2(\spiking_network_top_uut.all_data_out[236] ),
    .A2(_03785_),
    .A1(\spiking_network_top_uut.all_data_out[252] ));
 sg13g2_a22oi_1 _11330_ (.Y(_04344_),
    .B1(_03878_),
    .B2(\spiking_network_top_uut.all_data_out[868] ),
    .A2(_03795_),
    .A1(\spiking_network_top_uut.all_data_out[268] ));
 sg13g2_nand4_1 _11331_ (.B(_04342_),
    .C(_04343_),
    .A(_04341_),
    .Y(_04345_),
    .D(_04344_));
 sg13g2_a22oi_1 _11332_ (.Y(_04346_),
    .B1(_03856_),
    .B2(\spiking_network_top_uut.all_data_out[620] ),
    .A2(net3711),
    .A1(\spiking_network_top_uut.all_data_out[36] ));
 sg13g2_a22oi_1 _11333_ (.Y(_04347_),
    .B1(_03814_),
    .B2(\spiking_network_top_uut.all_data_out[628] ),
    .A2(_03783_),
    .A1(\spiking_network_top_uut.all_data_out[460] ));
 sg13g2_a22oi_1 _11334_ (.Y(_04348_),
    .B1(_03822_),
    .B2(\spiking_network_top_uut.all_data_out[452] ),
    .A2(_03810_),
    .A1(\spiking_network_top_uut.all_data_out[852] ));
 sg13g2_a22oi_1 _11335_ (.Y(_04349_),
    .B1(_03847_),
    .B2(\spiking_network_top_uut.all_data_out[404] ),
    .A2(_03835_),
    .A1(\spiking_network_top_uut.all_data_out[660] ));
 sg13g2_nand4_1 _11336_ (.B(_04347_),
    .C(_04348_),
    .A(_04346_),
    .Y(_04350_),
    .D(_04349_));
 sg13g2_nor4_1 _11337_ (.A(_03756_),
    .B(_04340_),
    .C(_04345_),
    .D(_04350_),
    .Y(_04351_));
 sg13g2_a22oi_1 _11338_ (.Y(_04352_),
    .B1(_03885_),
    .B2(\spiking_network_top_uut.all_data_out[516] ),
    .A2(_03813_),
    .A1(\spiking_network_top_uut.all_data_out[724] ));
 sg13g2_a22oi_1 _11339_ (.Y(_04353_),
    .B1(_03884_),
    .B2(\spiking_network_top_uut.all_data_out[796] ),
    .A2(_03862_),
    .A1(\spiking_network_top_uut.all_data_out[700] ));
 sg13g2_a22oi_1 _11340_ (.Y(_04354_),
    .B1(_03820_),
    .B2(\spiking_network_top_uut.all_data_out[164] ),
    .A2(_03788_),
    .A1(\spiking_network_top_uut.all_data_out[156] ));
 sg13g2_nand4_1 _11341_ (.B(_04352_),
    .C(_04353_),
    .A(_04311_),
    .Y(_04355_),
    .D(_04354_));
 sg13g2_a22oi_1 _11342_ (.Y(_04356_),
    .B1(_03887_),
    .B2(\spiking_network_top_uut.all_data_out[772] ),
    .A2(_03852_),
    .A1(\spiking_network_top_uut.all_data_out[396] ));
 sg13g2_a22oi_1 _11343_ (.Y(_04357_),
    .B1(_03844_),
    .B2(\spiking_network_top_uut.all_data_out[356] ),
    .A2(net3718),
    .A1(\spiking_network_top_uut.all_data_out[60] ));
 sg13g2_a22oi_1 _11344_ (.Y(_04358_),
    .B1(_03879_),
    .B2(\spiking_network_top_uut.all_data_out[212] ),
    .A2(_03861_),
    .A1(\spiking_network_top_uut.all_data_out[764] ));
 sg13g2_nand4_1 _11345_ (.B(_04356_),
    .C(_04357_),
    .A(_04312_),
    .Y(_04359_),
    .D(_04358_));
 sg13g2_a22oi_1 _11346_ (.Y(_04360_),
    .B1(_03763_),
    .B2(\spiking_network_top_uut.all_data_out[188] ),
    .A2(net3714),
    .A1(\spiking_network_top_uut.all_data_out[100] ));
 sg13g2_a22oi_1 _11347_ (.Y(_04361_),
    .B1(_03760_),
    .B2(\spiking_network_top_uut.all_data_out[604] ),
    .A2(_03747_),
    .A1(\spiking_network_top_uut.all_data_out[92] ));
 sg13g2_a22oi_1 _11348_ (.Y(_04362_),
    .B1(_03831_),
    .B2(\spiking_network_top_uut.all_data_out[324] ),
    .A2(_03777_),
    .A1(\spiking_network_top_uut.all_data_out[412] ));
 sg13g2_nand4_1 _11349_ (.B(_04360_),
    .C(_04361_),
    .A(_04313_),
    .Y(_04363_),
    .D(_04362_));
 sg13g2_a22oi_1 _11350_ (.Y(_04364_),
    .B1(_03848_),
    .B2(\spiking_network_top_uut.all_data_out[820] ),
    .A2(net3712),
    .A1(\spiking_network_top_uut.all_data_out[124] ));
 sg13g2_nand4_1 _11351_ (.B(_04319_),
    .C(_04320_),
    .A(_04315_),
    .Y(_04365_),
    .D(_04364_));
 sg13g2_nor4_1 _11352_ (.A(_04355_),
    .B(_04359_),
    .C(_04363_),
    .D(_04365_),
    .Y(_04366_));
 sg13g2_a22oi_1 _11353_ (.Y(_04367_),
    .B1(_03869_),
    .B2(\spiking_network_top_uut.all_data_out[364] ),
    .A2(_03779_),
    .A1(net4272));
 sg13g2_a22oi_1 _11354_ (.Y(_04368_),
    .B1(_03855_),
    .B2(\spiking_network_top_uut.all_data_out[332] ),
    .A2(_03781_),
    .A1(\spiking_network_top_uut.all_data_out[636] ));
 sg13g2_nand4_1 _11355_ (.B(_04317_),
    .C(_04367_),
    .A(_04314_),
    .Y(_04369_),
    .D(_04368_));
 sg13g2_a22oi_1 _11356_ (.Y(_04370_),
    .B1(_03849_),
    .B2(\spiking_network_top_uut.all_data_out[468] ),
    .A2(_03834_),
    .A1(\spiking_network_top_uut.all_data_out[708] ));
 sg13g2_a22oi_1 _11357_ (.Y(_04371_),
    .B1(_03864_),
    .B2(\spiking_network_top_uut.all_data_out[524] ),
    .A2(net3693),
    .A1(\spiking_network_top_uut.all_data_out[76] ));
 sg13g2_a22oi_1 _11358_ (.Y(_04372_),
    .B1(_03843_),
    .B2(\spiking_network_top_uut.all_data_out[436] ),
    .A2(net3716),
    .A1(\spiking_network_top_uut.all_data_out[44] ));
 sg13g2_nand4_1 _11359_ (.B(_04370_),
    .C(_04371_),
    .A(_04318_),
    .Y(_04373_),
    .D(_04372_));
 sg13g2_a22oi_1 _11360_ (.Y(_04374_),
    .B1(_03880_),
    .B2(\spiking_network_top_uut.all_data_out[548] ),
    .A2(_03784_),
    .A1(\spiking_network_top_uut.all_data_out[588] ));
 sg13g2_a22oi_1 _11361_ (.Y(_04375_),
    .B1(_03838_),
    .B2(\spiking_network_top_uut.all_data_out[788] ),
    .A2(_03723_),
    .A1(\spiking_network_top_uut.all_data_out[388] ));
 sg13g2_a22oi_1 _11362_ (.Y(_04376_),
    .B1(_03826_),
    .B2(\spiking_network_top_uut.all_data_out[836] ),
    .A2(net3713),
    .A1(\spiking_network_top_uut.all_data_out[116] ));
 sg13g2_a22oi_1 _11363_ (.Y(_04377_),
    .B1(_03845_),
    .B2(\spiking_network_top_uut.all_data_out[740] ),
    .A2(_03772_),
    .A1(\spiking_network_top_uut.all_data_out[380] ));
 sg13g2_nand4_1 _11364_ (.B(_04375_),
    .C(_04376_),
    .A(_04374_),
    .Y(_04378_),
    .D(_04377_));
 sg13g2_a22oi_1 _11365_ (.Y(_04379_),
    .B1(_03833_),
    .B2(\spiking_network_top_uut.all_data_out[484] ),
    .A2(_03821_),
    .A1(\spiking_network_top_uut.all_data_out[308] ));
 sg13g2_a22oi_1 _11366_ (.Y(_04380_),
    .B1(_03883_),
    .B2(\spiking_network_top_uut.all_data_out[684] ),
    .A2(_03839_),
    .A1(\spiking_network_top_uut.all_data_out[804] ));
 sg13g2_a22oi_1 _11367_ (.Y(_04381_),
    .B1(_03803_),
    .B2(\spiking_network_top_uut.all_data_out[180] ),
    .A2(_03782_),
    .A1(\spiking_network_top_uut.all_data_out[140] ));
 sg13g2_a22oi_1 _11368_ (.Y(_04382_),
    .B1(_03811_),
    .B2(\spiking_network_top_uut.all_data_out[372] ),
    .A2(_03806_),
    .A1(\spiking_network_top_uut.all_data_out[260] ));
 sg13g2_nand4_1 _11369_ (.B(_04380_),
    .C(_04381_),
    .A(_04379_),
    .Y(_04383_),
    .D(_04382_));
 sg13g2_nor4_2 _11370_ (.A(_04369_),
    .B(_04373_),
    .C(_04378_),
    .Y(_04384_),
    .D(_04383_));
 sg13g2_nand3_1 _11371_ (.B(_04366_),
    .C(_04384_),
    .A(_04351_),
    .Y(_04385_));
 sg13g2_a21oi_1 _11372_ (.A1(_03575_),
    .A2(_03756_),
    .Y(_04386_),
    .B1(_03471_));
 sg13g2_nand2b_2 _11373_ (.Y(_04387_),
    .B(_03878_),
    .A_N(_00214_));
 sg13g2_nand2_1 _11374_ (.Y(_04388_),
    .A(\spiking_network_top_uut.all_data_out[69] ),
    .B(net3696));
 sg13g2_nand2b_1 _11375_ (.Y(_04389_),
    .B(_03848_),
    .A_N(_00220_));
 sg13g2_nor3_2 _11376_ (.A(_00254_),
    .B(net3773),
    .C(net3769),
    .Y(_04390_));
 sg13g2_nor2_1 _11377_ (.A(_00256_),
    .B(_03841_),
    .Y(_04391_));
 sg13g2_nand2b_1 _11378_ (.Y(_04392_),
    .B(_03833_),
    .A_N(_00262_));
 sg13g2_nor3_2 _11379_ (.A(_00260_),
    .B(net3775),
    .C(net3774),
    .Y(_04393_));
 sg13g2_nand2_1 _11380_ (.Y(_04394_),
    .A(\spiking_network_top_uut.all_data_out[293] ),
    .B(_03819_));
 sg13g2_nor3_1 _11381_ (.A(_00240_),
    .B(net3771),
    .C(net3765),
    .Y(_04395_));
 sg13g2_nor3_1 _11382_ (.A(_00212_),
    .B(net3774),
    .C(net3757),
    .Y(_04396_));
 sg13g2_nand2b_2 _11383_ (.Y(_04397_),
    .B(_03784_),
    .A_N(_00249_));
 sg13g2_nand2b_2 _11384_ (.Y(_04398_),
    .B(_03862_),
    .A_N(_00235_));
 sg13g2_nand2b_1 _11385_ (.Y(_04399_),
    .B(_03868_),
    .A_N(_00219_));
 sg13g2_o21ai_1 _11386_ (.B1(_04399_),
    .Y(_04400_),
    .A1(_00211_),
    .A2(_03791_));
 sg13g2_nand2_2 _11387_ (.Y(_04401_),
    .A(\spiking_network_top_uut.all_data_out[173] ),
    .B(_03776_));
 sg13g2_nand2b_1 _11388_ (.Y(_04402_),
    .B(_03794_),
    .A_N(_00255_));
 sg13g2_o21ai_1 _11389_ (.B1(_04402_),
    .Y(_04403_),
    .A1(_00269_),
    .A2(_03800_));
 sg13g2_nand2b_1 _11390_ (.Y(_04404_),
    .B(_03783_),
    .A_N(_00265_));
 sg13g2_nand2b_2 _11391_ (.Y(_04405_),
    .B(_03844_),
    .A_N(_00278_));
 sg13g2_nor3_1 _11392_ (.A(_00224_),
    .B(net3771),
    .C(net3759),
    .Y(_04406_));
 sg13g2_nand2b_1 _11393_ (.Y(_04407_),
    .B(_03852_),
    .A_N(_00273_));
 sg13g2_nand2b_2 _11394_ (.Y(_04408_),
    .B(_03884_),
    .A_N(_00223_));
 sg13g2_nor3_2 _11395_ (.A(_00275_),
    .B(_03729_),
    .C(net3760),
    .Y(_04409_));
 sg13g2_nand2_2 _11396_ (.Y(_04410_),
    .A(\spiking_network_top_uut.all_data_out[205] ),
    .B(_03801_));
 sg13g2_nor2_1 _11397_ (.A(_00229_),
    .B(_03854_),
    .Y(_04411_));
 sg13g2_nand2b_1 _11398_ (.Y(_04412_),
    .B(_03781_),
    .A_N(_00243_));
 sg13g2_nor3_1 _11399_ (.A(_00251_),
    .B(net3779),
    .C(net3770),
    .Y(_04413_));
 sg13g2_nand2b_1 _11400_ (.Y(_04414_),
    .B(_03777_),
    .A_N(_00271_));
 sg13g2_nor2_2 _11401_ (.A(_00263_),
    .B(_03873_),
    .Y(_04415_));
 sg13g2_nand2_1 _11402_ (.Y(_04416_),
    .A(\spiking_network_top_uut.all_data_out[61] ),
    .B(net3718));
 sg13g2_nor3_2 _11403_ (.A(_00221_),
    .B(net3778),
    .C(net3759),
    .Y(_04417_));
 sg13g2_nor2_1 _11404_ (.A(_00226_),
    .B(_03888_),
    .Y(_04418_));
 sg13g2_nand2b_2 _11405_ (.Y(_04419_),
    .B(_03789_),
    .A_N(_00213_));
 sg13g2_a22oi_1 _11406_ (.Y(_04420_),
    .B1(net3709),
    .B2(\spiking_network_top_uut.all_data_out[21] ),
    .A2(net3719),
    .A1(\spiking_network_top_uut.all_data_out[29] ));
 sg13g2_a22oi_1 _11407_ (.Y(_04421_),
    .B1(_03803_),
    .B2(\spiking_network_top_uut.all_data_out[181] ),
    .A2(net3712),
    .A1(\spiking_network_top_uut.all_data_out[125] ));
 sg13g2_o21ai_1 _11408_ (.B1(_04404_),
    .Y(_04422_),
    .A1(_00244_),
    .A2(_03815_));
 sg13g2_a221oi_1 _11409_ (.B2(_03558_),
    .C1(_04422_),
    .B1(_03802_),
    .A1(\spiking_network_top_uut.all_data_out[189] ),
    .Y(_04423_),
    .A2(_03763_));
 sg13g2_nand3_1 _11410_ (.B(_04421_),
    .C(_04423_),
    .A(_04420_),
    .Y(_04424_));
 sg13g2_a221oi_1 _11411_ (.B2(\spiking_network_top_uut.all_data_out[85] ),
    .C1(_04413_),
    .B1(net3694),
    .A1(\spiking_network_top_uut.all_data_out[45] ),
    .Y(_04425_),
    .A2(net3716));
 sg13g2_nand2_1 _11412_ (.Y(_04426_),
    .A(_04419_),
    .B(_04425_));
 sg13g2_a21oi_1 _11413_ (.A1(\spiking_network_top_uut.all_data_out[277] ),
    .A2(_03816_),
    .Y(_04427_),
    .B1(_04403_));
 sg13g2_a221oi_1 _11414_ (.B2(\spiking_network_top_uut.all_data_out[149] ),
    .C1(_04391_),
    .B1(_03877_),
    .A1(_03553_),
    .Y(_04428_),
    .A2(_03807_));
 sg13g2_o21ai_1 _11415_ (.B1(_04428_),
    .Y(_04429_),
    .A1(_00241_),
    .A2(_03768_));
 sg13g2_a21oi_1 _11416_ (.A1(\spiking_network_top_uut.all_data_out[157] ),
    .A2(_03788_),
    .Y(_04430_),
    .B1(_04429_));
 sg13g2_nand2_1 _11417_ (.Y(_04431_),
    .A(_04427_),
    .B(_04430_));
 sg13g2_a22oi_1 _11418_ (.Y(_04432_),
    .B1(_03836_),
    .B2(_03564_),
    .A2(_03810_),
    .A1(_03549_));
 sg13g2_o21ai_1 _11419_ (.B1(_04432_),
    .Y(_04433_),
    .A1(_00279_),
    .A2(_03871_));
 sg13g2_a221oi_1 _11420_ (.B2(_03573_),
    .C1(_04433_),
    .B1(_03869_),
    .A1(\spiking_network_top_uut.all_data_out[269] ),
    .Y(_04434_),
    .A2(_03795_));
 sg13g2_a22oi_1 _11421_ (.Y(_04435_),
    .B1(_03846_),
    .B2(\spiking_network_top_uut.all_data_out[341] ),
    .A2(net3710),
    .A1(\spiking_network_top_uut.all_data_out[53] ));
 sg13g2_o21ai_1 _11422_ (.B1(_04435_),
    .Y(_04436_),
    .A1(_00245_),
    .A2(_03857_));
 sg13g2_a221oi_1 _11423_ (.B2(\spiking_network_top_uut.all_data_out[317] ),
    .C1(_04436_),
    .B1(_03867_),
    .A1(\spiking_network_top_uut.all_data_out[245] ),
    .Y(_04437_),
    .A2(_03812_));
 sg13g2_a221oi_1 _11424_ (.B2(\spiking_network_top_uut.all_data_out[221] ),
    .C1(_04396_),
    .B1(_03780_),
    .A1(_03563_),
    .Y(_04438_),
    .A2(_03760_));
 sg13g2_a221oi_1 _11425_ (.B2(_03556_),
    .C1(_04415_),
    .B1(_03813_),
    .A1(\spiking_network_top_uut.all_data_out[117] ),
    .Y(_04439_),
    .A2(net3713));
 sg13g2_nand4_1 _11426_ (.B(_04437_),
    .C(_04438_),
    .A(_04434_),
    .Y(_04440_),
    .D(_04439_));
 sg13g2_nor4_2 _11427_ (.A(_04424_),
    .B(_04426_),
    .C(_04431_),
    .Y(_04441_),
    .D(_04440_));
 sg13g2_a221oi_1 _11428_ (.B2(\spiking_network_top_uut.all_data_out[197] ),
    .C1(_04418_),
    .B1(_03830_),
    .A1(\spiking_network_top_uut.all_data_out[261] ),
    .Y(_04442_),
    .A2(_03806_));
 sg13g2_o21ai_1 _11429_ (.B1(_04392_),
    .Y(_04443_),
    .A1(_00270_),
    .A2(_03825_));
 sg13g2_a221oi_1 _11430_ (.B2(_03567_),
    .C1(_04443_),
    .B1(_03822_),
    .A1(\spiking_network_top_uut.all_data_out[133] ),
    .Y(_04444_),
    .A2(_03805_));
 sg13g2_nand3_1 _11431_ (.B(_04442_),
    .C(_04444_),
    .A(_04405_),
    .Y(_04445_));
 sg13g2_a22oi_1 _11432_ (.Y(_04446_),
    .B1(_03847_),
    .B2(_03570_),
    .A2(_03779_),
    .A1(\spiking_network_top_uut.all_data_out[13] ));
 sg13g2_nand4_1 _11433_ (.B(_04398_),
    .C(_04414_),
    .A(_04397_),
    .Y(_04447_),
    .D(_04446_));
 sg13g2_a22oi_1 _11434_ (.Y(_04448_),
    .B1(_03845_),
    .B2(_03554_),
    .A2(_03842_),
    .A1(_03562_));
 sg13g2_o21ai_1 _11435_ (.B1(_04448_),
    .Y(_04449_),
    .A1(_00218_),
    .A2(_03827_));
 sg13g2_a221oi_1 _11436_ (.B2(_03557_),
    .C1(_04449_),
    .B1(_03834_),
    .A1(\spiking_network_top_uut.all_data_out[901] ),
    .Y(_04450_),
    .A2(_03744_));
 sg13g2_o21ai_1 _11437_ (.B1(_04388_),
    .Y(_04451_),
    .A1(_00250_),
    .A2(_03809_));
 sg13g2_a221oi_1 _11438_ (.B2(\spiking_network_top_uut.all_data_out[165] ),
    .C1(_04451_),
    .B1(_03820_),
    .A1(\spiking_network_top_uut.all_data_out[37] ),
    .Y(_04452_),
    .A2(net3711));
 sg13g2_a221oi_1 _11439_ (.B2(\spiking_network_top_uut.all_data_out[229] ),
    .C1(_04390_),
    .B1(_03828_),
    .A1(\spiking_network_top_uut.all_data_out[101] ),
    .Y(_04453_),
    .A2(net3714));
 sg13g2_nand3_1 _11440_ (.B(_04452_),
    .C(_04453_),
    .A(_04450_),
    .Y(_04454_));
 sg13g2_nor3_2 _11441_ (.A(_04445_),
    .B(_04447_),
    .C(_04454_),
    .Y(_04455_));
 sg13g2_o21ai_1 _11442_ (.B1(_04389_),
    .Y(_04456_),
    .A1(_00233_),
    .A2(_03860_));
 sg13g2_nor3_2 _11443_ (.A(_04395_),
    .B(_04411_),
    .C(_04456_),
    .Y(_04457_));
 sg13g2_a22oi_1 _11444_ (.Y(_04458_),
    .B1(_03843_),
    .B2(_03569_),
    .A2(_03798_),
    .A1(_03555_));
 sg13g2_o21ai_1 _11445_ (.B1(_04408_),
    .Y(_04459_),
    .A1(_00259_),
    .A2(_03797_));
 sg13g2_a221oi_1 _11446_ (.B2(_03559_),
    .C1(_04459_),
    .B1(_03883_),
    .A1(_03568_),
    .Y(_04460_),
    .A2(_03863_));
 sg13g2_and4_1 _11447_ (.A(_04412_),
    .B(_04457_),
    .C(_04458_),
    .D(_04460_),
    .X(_04461_));
 sg13g2_a22oi_1 _11448_ (.Y(_04462_),
    .B1(_03811_),
    .B2(_03572_),
    .A2(_03782_),
    .A1(\spiking_network_top_uut.all_data_out[141] ));
 sg13g2_o21ai_1 _11449_ (.B1(_04462_),
    .Y(_04463_),
    .A1(_00261_),
    .A2(_03787_));
 sg13g2_o21ai_1 _11450_ (.B1(_04407_),
    .Y(_04464_),
    .A1(_00264_),
    .A2(_03850_));
 sg13g2_o21ai_1 _11451_ (.B1(_04416_),
    .Y(_04465_),
    .A1(_00217_),
    .A2(_03875_));
 sg13g2_nor4_2 _11452_ (.A(_04406_),
    .B(_04463_),
    .C(_04464_),
    .Y(_04466_),
    .D(_04465_));
 sg13g2_nand4_1 _11453_ (.B(_04455_),
    .C(_04461_),
    .A(_04441_),
    .Y(_04467_),
    .D(_04466_));
 sg13g2_a221oi_1 _11454_ (.B2(\spiking_network_top_uut.all_data_out[285] ),
    .C1(_04393_),
    .B1(_03876_),
    .A1(\spiking_network_top_uut.all_data_out[109] ),
    .Y(_04468_),
    .A2(net3717));
 sg13g2_a22oi_1 _11455_ (.Y(_04469_),
    .B1(_03817_),
    .B2(_03565_),
    .A2(net3695),
    .A1(\spiking_network_top_uut.all_data_out[93] ));
 sg13g2_a22oi_1 _11456_ (.Y(_04470_),
    .B1(_03792_),
    .B2(\spiking_network_top_uut.all_data_out[237] ),
    .A2(net3693),
    .A1(\spiking_network_top_uut.all_data_out[77] ));
 sg13g2_nand4_1 _11457_ (.B(_04468_),
    .C(_04469_),
    .A(_04410_),
    .Y(_04471_),
    .D(_04470_));
 sg13g2_o21ai_1 _11458_ (.B1(_04394_),
    .Y(_04472_),
    .A1(_00258_),
    .A2(_03886_));
 sg13g2_a221oi_1 _11459_ (.B2(_03560_),
    .C1(_04472_),
    .B1(_03829_),
    .A1(_03571_),
    .Y(_04473_),
    .A2(net3715));
 sg13g2_o21ai_1 _11460_ (.B1(_04387_),
    .Y(_04474_),
    .A1(_00242_),
    .A2(_03891_));
 sg13g2_a221oi_1 _11461_ (.B2(_03550_),
    .C1(_04474_),
    .B1(_03839_),
    .A1(_03574_),
    .Y(_04475_),
    .A2(_03831_));
 sg13g2_a221oi_1 _11462_ (.B2(_03552_),
    .C1(_04409_),
    .B1(_03861_),
    .A1(_03548_),
    .Y(_04476_),
    .A2(_03775_));
 sg13g2_nand4_1 _11463_ (.B(_04473_),
    .C(_04475_),
    .A(_03757_),
    .Y(_04477_),
    .D(_04476_));
 sg13g2_a221oi_1 _11464_ (.B2(\spiking_network_top_uut.all_data_out[213] ),
    .C1(_04400_),
    .B1(_03879_),
    .A1(_03561_),
    .Y(_04478_),
    .A2(_03769_));
 sg13g2_o21ai_1 _11465_ (.B1(_04401_),
    .Y(_04479_),
    .A1(_00257_),
    .A2(_03865_));
 sg13g2_a221oi_1 _11466_ (.B2(\spiking_network_top_uut.all_data_out[333] ),
    .C1(_04479_),
    .B1(_03855_),
    .A1(_03566_),
    .Y(_04480_),
    .A2(_03764_));
 sg13g2_a221oi_1 _11467_ (.B2(\spiking_network_top_uut.all_data_out[309] ),
    .C1(_04417_),
    .B1(_03821_),
    .A1(\spiking_network_top_uut.all_data_out[253] ),
    .Y(_04481_),
    .A2(_03785_));
 sg13g2_a22oi_1 _11468_ (.Y(_04482_),
    .B1(_03882_),
    .B2(_03551_),
    .A2(_03866_),
    .A1(\spiking_network_top_uut.all_data_out[301] ));
 sg13g2_nand4_1 _11469_ (.B(_04480_),
    .C(_04481_),
    .A(_04478_),
    .Y(_04483_),
    .D(_04482_));
 sg13g2_nor4_2 _11470_ (.A(_04467_),
    .B(_04471_),
    .C(_04477_),
    .Y(_04484_),
    .D(_04483_));
 sg13g2_o21ai_1 _11471_ (.B1(_03471_),
    .Y(_04485_),
    .A1(\spiking_network_top_uut.all_data_out[5] ),
    .A2(_03757_));
 sg13g2_a21oi_1 _11472_ (.A1(_04385_),
    .A2(_04386_),
    .Y(_04486_),
    .B1(\spiking_network_top_uut.spi_inst.spi_slave_inst.bit_cnt[2] ));
 sg13g2_o21ai_1 _11473_ (.B1(_04486_),
    .Y(_04487_),
    .A1(_04484_),
    .A2(_04485_));
 sg13g2_nand2b_2 _11474_ (.Y(_04488_),
    .B(_03885_),
    .A_N(_00398_));
 sg13g2_nand2b_1 _11475_ (.Y(_04489_),
    .B(_03852_),
    .A_N(_00413_));
 sg13g2_nand2b_1 _11476_ (.Y(_04490_),
    .B(_03887_),
    .A_N(_00366_));
 sg13g2_nand2b_2 _11477_ (.Y(_04491_),
    .B(_03784_),
    .A_N(_00389_));
 sg13g2_nand2b_1 _11478_ (.Y(_04492_),
    .B(_03868_),
    .A_N(_00359_));
 sg13g2_nand2b_2 _11479_ (.Y(_04493_),
    .B(_03884_),
    .A_N(_00363_));
 sg13g2_nand2b_1 _11480_ (.Y(_04494_),
    .B(_03882_),
    .A_N(_00365_));
 sg13g2_nand2b_2 _11481_ (.Y(_04495_),
    .B(_03889_),
    .A_N(_00391_));
 sg13g2_nand2b_1 _11482_ (.Y(_04496_),
    .B(_03883_),
    .A_N(_00377_));
 sg13g2_nand2b_1 _11483_ (.Y(_04497_),
    .B(_03870_),
    .A_N(_00419_));
 sg13g2_nand2b_2 _11484_ (.Y(_04498_),
    .B(_03764_),
    .A_N(_00393_));
 sg13g2_nand2b_2 _11485_ (.Y(_04499_),
    .B(_03796_),
    .A_N(_00399_));
 sg13g2_nand2b_2 _11486_ (.Y(_04500_),
    .B(_03842_),
    .A_N(_00386_));
 sg13g2_nand2b_1 _11487_ (.Y(_04501_),
    .B(_03810_),
    .A_N(_00356_));
 sg13g2_nand2b_2 _11488_ (.Y(_04502_),
    .B(_03843_),
    .A_N(_00408_));
 sg13g2_nor3_1 _11489_ (.A(_00368_),
    .B(_03727_),
    .C(net3765),
    .Y(_04503_));
 sg13g2_nand2b_2 _11490_ (.Y(_04504_),
    .B(_03839_),
    .A_N(_00362_));
 sg13g2_nand2b_1 _11491_ (.Y(_04505_),
    .B(_03832_),
    .A_N(_00352_));
 sg13g2_nand2b_2 _11492_ (.Y(_04506_),
    .B(_03880_),
    .A_N(_00394_));
 sg13g2_nand2b_1 _11493_ (.Y(_04507_),
    .B(_03847_),
    .A_N(_00412_));
 sg13g2_nand2b_2 _11494_ (.Y(_04508_),
    .B(_03878_),
    .A_N(_00354_));
 sg13g2_nand2b_1 _11495_ (.Y(_04509_),
    .B(_03822_),
    .A_N(_00406_));
 sg13g2_nand2b_2 _11496_ (.Y(_04510_),
    .B(_03808_),
    .A_N(_00390_));
 sg13g2_nand2b_2 _11497_ (.Y(_04511_),
    .B(_03833_),
    .A_N(_00402_));
 sg13g2_nand2b_1 _11498_ (.Y(_04512_),
    .B(_03838_),
    .A_N(_00364_));
 sg13g2_nand2b_2 _11499_ (.Y(_04513_),
    .B(_03849_),
    .A_N(_00404_));
 sg13g2_nand2b_2 _11500_ (.Y(_04514_),
    .B(_03804_),
    .A_N(_00400_));
 sg13g2_nor3_2 _11501_ (.A(_00367_),
    .B(_03729_),
    .C(net3765),
    .Y(_04515_));
 sg13g2_nand2b_1 _11502_ (.Y(_04516_),
    .B(_03851_),
    .A_N(_00361_));
 sg13g2_nand2b_1 _11503_ (.Y(_04517_),
    .B(_03794_),
    .A_N(_00395_));
 sg13g2_nand2b_1 _11504_ (.Y(_04518_),
    .B(_03772_),
    .A_N(_00415_));
 sg13g2_nand2b_1 _11505_ (.Y(_04519_),
    .B(_03872_),
    .A_N(_00403_));
 sg13g2_nand2b_1 _11506_ (.Y(_04520_),
    .B(_03775_),
    .A_N(_00355_));
 sg13g2_a22oi_1 _11507_ (.Y(_04521_),
    .B1(_03831_),
    .B2(_03654_),
    .A2(_03812_),
    .A1(\spiking_network_top_uut.all_data_out[241] ));
 sg13g2_nand2_1 _11508_ (.Y(_04522_),
    .A(_03471_),
    .B(\spiking_network_top_uut.spi_inst.spi_slave_inst.bit_cnt[2] ));
 sg13g2_o21ai_1 _11509_ (.B1(_04491_),
    .Y(_04523_),
    .A1(_00384_),
    .A2(_03815_));
 sg13g2_a221oi_1 _11510_ (.B2(\spiking_network_top_uut.all_data_out[153] ),
    .C1(_04523_),
    .B1(_03788_),
    .A1(\spiking_network_top_uut.all_data_out[89] ),
    .Y(_04524_),
    .A2(net3695));
 sg13g2_a22oi_1 _11511_ (.Y(_04525_),
    .B1(_03877_),
    .B2(\spiking_network_top_uut.all_data_out[145] ),
    .A2(_03803_),
    .A1(\spiking_network_top_uut.all_data_out[177] ));
 sg13g2_a22oi_1 _11512_ (.Y(_04526_),
    .B1(_03783_),
    .B2(_03648_),
    .A2(net3712),
    .A1(\spiking_network_top_uut.all_data_out[121] ));
 sg13g2_a22oi_1 _11513_ (.Y(_04527_),
    .B1(_03862_),
    .B2(_03639_),
    .A2(_03855_),
    .A1(\spiking_network_top_uut.all_data_out[329] ));
 sg13g2_o21ai_1 _11514_ (.B1(_04489_),
    .Y(_04528_),
    .A1(_00411_),
    .A2(_03778_));
 sg13g2_o21ai_1 _11515_ (.B1(_04516_),
    .Y(_04529_),
    .A1(_00397_),
    .A2(_03865_));
 sg13g2_o21ai_1 _11516_ (.B1(_04517_),
    .Y(_04530_),
    .A1(_00392_),
    .A2(_03818_));
 sg13g2_o21ai_1 _11517_ (.B1(_04496_),
    .Y(_04531_),
    .A1(_00369_),
    .A2(_03854_));
 sg13g2_a22oi_1 _11518_ (.Y(_04532_),
    .B1(_03779_),
    .B2(net4282),
    .A2(_03776_),
    .A1(\spiking_network_top_uut.all_data_out[169] ));
 sg13g2_o21ai_1 _11519_ (.B1(_04512_),
    .Y(_04533_),
    .A1(_00409_),
    .A2(_03800_));
 sg13g2_o21ai_1 _11520_ (.B1(_04501_),
    .Y(_04534_),
    .A1(_00357_),
    .A2(_03875_));
 sg13g2_a22oi_1 _11521_ (.Y(_04535_),
    .B1(_03835_),
    .B2(_03643_),
    .A2(_03813_),
    .A1(_03637_));
 sg13g2_a22oi_1 _11522_ (.Y(_04536_),
    .B1(_03834_),
    .B2(_03638_),
    .A2(_03820_),
    .A1(\spiking_network_top_uut.all_data_out[161] ));
 sg13g2_a22oi_1 _11523_ (.Y(_04537_),
    .B1(_03748_),
    .B2(\spiking_network_top_uut.all_data_out[81] ),
    .A2(net3713),
    .A1(\spiking_network_top_uut.all_data_out[113] ));
 sg13g2_o21ai_1 _11524_ (.B1(_04510_),
    .Y(_04538_),
    .A1(_00373_),
    .A2(_03860_));
 sg13g2_a221oi_1 _11525_ (.B2(_03635_),
    .C1(_04538_),
    .B1(_03845_),
    .A1(_03636_),
    .Y(_04539_),
    .A2(_03798_));
 sg13g2_nand4_1 _11526_ (.B(_04498_),
    .C(_04537_),
    .A(_04495_),
    .Y(_04540_),
    .D(_04539_));
 sg13g2_a22oi_1 _11527_ (.Y(_04541_),
    .B1(_03869_),
    .B2(_03652_),
    .A2(net3718),
    .A1(\spiking_network_top_uut.all_data_out[57] ));
 sg13g2_o21ai_1 _11528_ (.B1(_04490_),
    .Y(_04542_),
    .A1(_00382_),
    .A2(_03891_));
 sg13g2_a221oi_1 _11529_ (.B2(\spiking_network_top_uut.all_data_out[201] ),
    .C1(_04542_),
    .B1(_03801_),
    .A1(\spiking_network_top_uut.all_data_out[49] ),
    .Y(_04543_),
    .A2(net3710));
 sg13g2_nand4_1 _11530_ (.B(_04514_),
    .C(_04541_),
    .A(_04499_),
    .Y(_04544_),
    .D(_04543_));
 sg13g2_a22oi_1 _11531_ (.Y(_04545_),
    .B1(_03805_),
    .B2(\spiking_network_top_uut.all_data_out[129] ),
    .A2(_03802_),
    .A1(_03640_));
 sg13g2_a22oi_1 _11532_ (.Y(_04546_),
    .B1(_03866_),
    .B2(\spiking_network_top_uut.all_data_out[297] ),
    .A2(_03821_),
    .A1(\spiking_network_top_uut.all_data_out[305] ));
 sg13g2_a22oi_1 _11533_ (.Y(_04547_),
    .B1(_03876_),
    .B2(\spiking_network_top_uut.all_data_out[281] ),
    .A2(_03867_),
    .A1(\spiking_network_top_uut.all_data_out[313] ));
 sg13g2_nand4_1 _11534_ (.B(_04545_),
    .C(_04546_),
    .A(_04526_),
    .Y(_04548_),
    .D(_04547_));
 sg13g2_nand3_1 _11535_ (.B(_04525_),
    .C(_04536_),
    .A(_04524_),
    .Y(_04549_));
 sg13g2_nor4_1 _11536_ (.A(_04540_),
    .B(_04544_),
    .C(_04548_),
    .D(_04549_),
    .Y(_04550_));
 sg13g2_a22oi_1 _11537_ (.Y(_04551_),
    .B1(_03780_),
    .B2(\spiking_network_top_uut.all_data_out[217] ),
    .A2(net3716),
    .A1(\spiking_network_top_uut.all_data_out[41] ));
 sg13g2_a22oi_1 _11538_ (.Y(_04552_),
    .B1(_03848_),
    .B2(_03634_),
    .A2(_03744_),
    .A1(\spiking_network_top_uut.all_data_out[897] ));
 sg13g2_nand4_1 _11539_ (.B(_04493_),
    .C(_04551_),
    .A(_04488_),
    .Y(_04553_),
    .D(_04552_));
 sg13g2_a22oi_1 _11540_ (.Y(_04554_),
    .B1(_03844_),
    .B2(_03653_),
    .A2(net3709),
    .A1(\spiking_network_top_uut.all_data_out[17] ));
 sg13g2_a22oi_1 _11541_ (.Y(_04555_),
    .B1(net3711),
    .B2(\spiking_network_top_uut.all_data_out[33] ),
    .A2(net3719),
    .A1(\spiking_network_top_uut.all_data_out[25] ));
 sg13g2_a22oi_1 _11542_ (.Y(_04556_),
    .B1(_03879_),
    .B2(\spiking_network_top_uut.all_data_out[209] ),
    .A2(_03785_),
    .A1(\spiking_network_top_uut.all_data_out[249] ));
 sg13g2_nand4_1 _11543_ (.B(_04554_),
    .C(_04555_),
    .A(_04527_),
    .Y(_04557_),
    .D(_04556_));
 sg13g2_o21ai_1 _11544_ (.B1(_04507_),
    .Y(_04558_),
    .A1(_00410_),
    .A2(_03825_));
 sg13g2_o21ai_1 _11545_ (.B1(_04492_),
    .Y(_04559_),
    .A1(_00358_),
    .A2(_03827_));
 sg13g2_nor3_1 _11546_ (.A(_04529_),
    .B(_04558_),
    .C(_04559_),
    .Y(_04560_));
 sg13g2_o21ai_1 _11547_ (.B1(_04504_),
    .Y(_04561_),
    .A1(_00401_),
    .A2(_03787_));
 sg13g2_o21ai_1 _11548_ (.B1(_04520_),
    .Y(_04562_),
    .A1(_00351_),
    .A2(_03791_));
 sg13g2_o21ai_1 _11549_ (.B1(_04494_),
    .Y(_04563_),
    .A1(_00385_),
    .A2(_03857_));
 sg13g2_nor4_2 _11550_ (.A(_04533_),
    .B(_04561_),
    .C(_04562_),
    .Y(_04564_),
    .D(_04563_));
 sg13g2_nand4_1 _11551_ (.B(_04506_),
    .C(_04560_),
    .A(_04500_),
    .Y(_04565_),
    .D(_04564_));
 sg13g2_nor4_2 _11552_ (.A(_04528_),
    .B(_04553_),
    .C(_04557_),
    .Y(_04566_),
    .D(_04565_));
 sg13g2_a22oi_1 _11553_ (.Y(_04567_),
    .B1(_03781_),
    .B2(_03645_),
    .A2(_03760_),
    .A1(_03646_));
 sg13g2_a221oi_1 _11554_ (.B2(_03633_),
    .C1(_04534_),
    .B1(_03789_),
    .A1(\spiking_network_top_uut.all_data_out[105] ),
    .Y(_04568_),
    .A2(net3717));
 sg13g2_nand4_1 _11555_ (.B(_04511_),
    .C(_04567_),
    .A(_04505_),
    .Y(_04569_),
    .D(_04568_));
 sg13g2_a22oi_1 _11556_ (.Y(_04570_),
    .B1(_03863_),
    .B2(_03649_),
    .A2(_03816_),
    .A1(\spiking_network_top_uut.all_data_out[273] ));
 sg13g2_o21ai_1 _11557_ (.B1(_04508_),
    .Y(_04571_),
    .A1(_00388_),
    .A2(_03837_));
 sg13g2_a221oi_1 _11558_ (.B2(\spiking_network_top_uut.all_data_out[265] ),
    .C1(_04571_),
    .B1(_03795_),
    .A1(_03644_),
    .Y(_04572_),
    .A2(_03767_));
 sg13g2_nand4_1 _11559_ (.B(_04509_),
    .C(_04570_),
    .A(_04502_),
    .Y(_04573_),
    .D(_04572_));
 sg13g2_a22oi_1 _11560_ (.Y(_04574_),
    .B1(_03830_),
    .B2(\spiking_network_top_uut.all_data_out[193] ),
    .A2(_03763_),
    .A1(\spiking_network_top_uut.all_data_out[185] ));
 sg13g2_a22oi_1 _11561_ (.Y(_04575_),
    .B1(_03846_),
    .B2(\spiking_network_top_uut.all_data_out[337] ),
    .A2(_03828_),
    .A1(\spiking_network_top_uut.all_data_out[225] ));
 sg13g2_a22oi_1 _11562_ (.Y(_04576_),
    .B1(_03811_),
    .B2(_03651_),
    .A2(net3696),
    .A1(\spiking_network_top_uut.all_data_out[65] ));
 sg13g2_nand4_1 _11563_ (.B(_04574_),
    .C(_04575_),
    .A(_04521_),
    .Y(_04577_),
    .D(_04576_));
 sg13g2_nor4_2 _11564_ (.A(_04503_),
    .B(_04515_),
    .C(_04530_),
    .Y(_04578_),
    .D(_04531_));
 sg13g2_a22oi_1 _11565_ (.Y(_04579_),
    .B1(_03819_),
    .B2(\spiking_network_top_uut.all_data_out[289] ),
    .A2(_03769_),
    .A1(_03642_));
 sg13g2_nand4_1 _11566_ (.B(_04519_),
    .C(_04535_),
    .A(_04513_),
    .Y(_04580_),
    .D(_04579_));
 sg13g2_a221oi_1 _11567_ (.B2(_03641_),
    .C1(_04580_),
    .B1(_03829_),
    .A1(\spiking_network_top_uut.all_data_out[137] ),
    .Y(_04581_),
    .A2(_03782_));
 sg13g2_a22oi_1 _11568_ (.Y(_04582_),
    .B1(_03840_),
    .B2(_03647_),
    .A2(net3693),
    .A1(\spiking_network_top_uut.all_data_out[73] ));
 sg13g2_a22oi_1 _11569_ (.Y(_04583_),
    .B1(net3714),
    .B2(\spiking_network_top_uut.all_data_out[97] ),
    .A2(net3715),
    .A1(_03650_));
 sg13g2_nand4_1 _11570_ (.B(_04518_),
    .C(_04582_),
    .A(_04497_),
    .Y(_04584_),
    .D(_04583_));
 sg13g2_a221oi_1 _11571_ (.B2(\spiking_network_top_uut.all_data_out[257] ),
    .C1(_04584_),
    .B1(_03806_),
    .A1(\spiking_network_top_uut.all_data_out[233] ),
    .Y(_04585_),
    .A2(_03792_));
 sg13g2_nand4_1 _11572_ (.B(_04578_),
    .C(_04581_),
    .A(_04532_),
    .Y(_04586_),
    .D(_04585_));
 sg13g2_nor4_1 _11573_ (.A(_04569_),
    .B(_04573_),
    .C(_04577_),
    .D(_04586_),
    .Y(_04587_));
 sg13g2_a21oi_2 _11574_ (.B1(_04522_),
    .Y(_04588_),
    .A2(_03756_),
    .A1(net4267));
 sg13g2_nand4_1 _11575_ (.B(_04566_),
    .C(_04587_),
    .A(_04550_),
    .Y(_04589_),
    .D(_04588_));
 sg13g2_nand3_1 _11576_ (.B(_04487_),
    .C(_04589_),
    .A(\spiking_network_top_uut.spi_inst.spi_slave_inst.bit_cnt[1] ),
    .Y(_04590_));
 sg13g2_nor2_1 _11577_ (.A(net10),
    .B(_04310_),
    .Y(_04591_));
 sg13g2_a22oi_1 _11578_ (.Y(_00022_),
    .B1(_04590_),
    .B2(_04591_),
    .A2(_03965_),
    .A1(_03964_));
 sg13g2_nor2_1 _11579_ (.A(net10),
    .B(\spiking_network_top_uut.spi_inst.spi_slave_inst.bit_cnt[0] ),
    .Y(_00023_));
 sg13g2_nor2_1 _11580_ (.A(\spiking_network_top_uut.spi_inst.spi_slave_inst.bit_cnt[0] ),
    .B(\spiking_network_top_uut.spi_inst.spi_slave_inst.bit_cnt[1] ),
    .Y(_04592_));
 sg13g2_nor3_1 _11581_ (.A(net10),
    .B(_03694_),
    .C(_04592_),
    .Y(_00024_));
 sg13g2_o21ai_1 _11582_ (.B1(_03470_),
    .Y(_04593_),
    .A1(_03655_),
    .A2(_03694_));
 sg13g2_a21oi_1 _11583_ (.A1(_03655_),
    .A2(_03694_),
    .Y(_00025_),
    .B1(_04593_));
 sg13g2_nand2_1 _11584_ (.Y(_04594_),
    .A(\spiking_network_top_uut.spi_inst.spi_control_unit_inst.current_state[1] ),
    .B(\spiking_network_top_uut.spi_inst.spi_control_unit_inst.current_state[0] ));
 sg13g2_nand3_1 _11585_ (.B(\spiking_network_top_uut.spi_inst.spi_control_unit_inst.current_state[0] ),
    .C(_00028_),
    .A(\spiking_network_top_uut.spi_inst.spi_control_unit_inst.current_state[1] ),
    .Y(_04595_));
 sg13g2_nor2_1 _11586_ (.A(_00029_),
    .B(_04595_),
    .Y(_00020_));
 sg13g2_o21ai_1 _11587_ (.B1(_03695_),
    .Y(_04596_),
    .A1(\spiking_network_top_uut.spi_inst.spi_control_unit_inst.current_state[2] ),
    .A2(_04594_));
 sg13g2_nor2b_1 _11588_ (.A(net4444),
    .B_N(net4465),
    .Y(_04597_));
 sg13g2_nor4_2 _11589_ (.A(net4365),
    .B(net4384),
    .C(net4322),
    .Y(_04598_),
    .D(net4342));
 sg13g2_nand4_1 _11590_ (.B(_04596_),
    .C(_04597_),
    .A(_00020_),
    .Y(_04599_),
    .D(_04598_));
 sg13g2_nor3_1 _11591_ (.A(net4422),
    .B(_03657_),
    .C(_04599_),
    .Y(_04600_));
 sg13g2_or2_1 _11592_ (.X(_10369_),
    .B(_04600_),
    .A(_02057_));
 sg13g2_nor3_1 _11593_ (.A(_03656_),
    .B(net4402),
    .C(_04599_),
    .Y(_04601_));
 sg13g2_or2_1 _11594_ (.X(_10370_),
    .B(_04601_),
    .A(_02058_));
 sg13g2_nor2_1 _11595_ (.A(\spiking_network_top_uut.debug_inst.debug_config[4] ),
    .B(\spiking_network_top_uut.debug_inst.debug_config[5] ),
    .Y(_04602_));
 sg13g2_nand3b_1 _11596_ (.B(_04602_),
    .C(\spiking_network_top_uut.debug_inst.debug_config[7] ),
    .Y(_04603_),
    .A_N(\spiking_network_top_uut.debug_inst.debug_config[6] ));
 sg13g2_nor2_1 _11597_ (.A(\spiking_network_top_uut.debug_inst.debug_config[2] ),
    .B(\spiking_network_top_uut.debug_inst.debug_config[3] ),
    .Y(_04604_));
 sg13g2_nor2b_1 _11598_ (.A(net4602),
    .B_N(net4600),
    .Y(_04605_));
 sg13g2_nand2_2 _11599_ (.Y(_04606_),
    .A(_04604_),
    .B(_04605_));
 sg13g2_nor2_2 _11600_ (.A(net3756),
    .B(_04606_),
    .Y(_04607_));
 sg13g2_nor2_1 _11601_ (.A(\spiking_network_top_uut.debug_inst.debug_config[4] ),
    .B(\spiking_network_top_uut.debug_inst.debug_config[7] ),
    .Y(_04608_));
 sg13g2_nand3b_1 _11602_ (.B(\spiking_network_top_uut.debug_inst.debug_config[6] ),
    .C(_04602_),
    .Y(_04609_),
    .A_N(\spiking_network_top_uut.debug_inst.debug_config[7] ));
 sg13g2_nor2_2 _11603_ (.A(_04606_),
    .B(_04609_),
    .Y(_04610_));
 sg13g2_nand2_1 _11604_ (.Y(_04611_),
    .A(net4602),
    .B(net4600));
 sg13g2_nand4_1 _11605_ (.B(net4601),
    .C(\spiking_network_top_uut.debug_inst.debug_config[2] ),
    .A(\spiking_network_top_uut.debug_inst.debug_config[0] ),
    .Y(_04612_),
    .D(\spiking_network_top_uut.debug_inst.debug_config[3] ));
 sg13g2_nor2_1 _11606_ (.A(net3756),
    .B(_04612_),
    .Y(_04613_));
 sg13g2_nor2b_2 _11607_ (.A(\spiking_network_top_uut.debug_inst.debug_config[3] ),
    .B_N(\spiking_network_top_uut.debug_inst.debug_config[2] ),
    .Y(_04614_));
 sg13g2_nand2b_1 _11608_ (.Y(_04615_),
    .B(\spiking_network_top_uut.debug_inst.debug_config[2] ),
    .A_N(\spiking_network_top_uut.debug_inst.debug_config[3] ));
 sg13g2_nand2_2 _11609_ (.Y(_04616_),
    .A(_04605_),
    .B(_04614_));
 sg13g2_nor2_2 _11610_ (.A(_04603_),
    .B(_04616_),
    .Y(_04617_));
 sg13g2_nand2_2 _11611_ (.Y(_04618_),
    .A(net4602),
    .B(_04604_));
 sg13g2_nor4_2 _11612_ (.A(\spiking_network_top_uut.debug_inst.debug_config[2] ),
    .B(\spiking_network_top_uut.debug_inst.debug_config[3] ),
    .C(net3756),
    .Y(_04619_),
    .D(_04611_));
 sg13g2_nand3b_1 _11613_ (.B(_04608_),
    .C(\spiking_network_top_uut.debug_inst.debug_config[5] ),
    .Y(_04620_),
    .A_N(\spiking_network_top_uut.debug_inst.debug_config[6] ));
 sg13g2_nor2_2 _11614_ (.A(_04606_),
    .B(_04620_),
    .Y(_04621_));
 sg13g2_nor3_1 _11615_ (.A(\spiking_network_top_uut.debug_inst.debug_config[0] ),
    .B(net4600),
    .C(\spiking_network_top_uut.debug_inst.debug_config[2] ),
    .Y(_04622_));
 sg13g2_nand2_1 _11616_ (.Y(_04623_),
    .A(\spiking_network_top_uut.debug_inst.debug_config[3] ),
    .B(_04622_));
 sg13g2_nor2_2 _11617_ (.A(_04609_),
    .B(_04623_),
    .Y(_04624_));
 sg13g2_nand2_1 _11618_ (.Y(_04625_),
    .A(net4602),
    .B(_04614_));
 sg13g2_nor2_2 _11619_ (.A(_04612_),
    .B(_04620_),
    .Y(_04626_));
 sg13g2_nor2_2 _11620_ (.A(_04609_),
    .B(_04616_),
    .Y(_04627_));
 sg13g2_nor2_2 _11621_ (.A(net3756),
    .B(_04623_),
    .Y(_04628_));
 sg13g2_nor4_2 _11622_ (.A(net4602),
    .B(net4600),
    .C(_04609_),
    .Y(_04629_),
    .D(_04615_));
 sg13g2_nor3_2 _11623_ (.A(net4601),
    .B(net3756),
    .C(_04618_),
    .Y(_04630_));
 sg13g2_nor4_2 _11624_ (.A(net4602),
    .B(net4600),
    .C(net3756),
    .Y(_04631_),
    .D(_04615_));
 sg13g2_nor3_2 _11625_ (.A(net4601),
    .B(_04618_),
    .C(_04620_),
    .Y(_04632_));
 sg13g2_nor3_2 _11626_ (.A(net4600),
    .B(_04609_),
    .C(_04625_),
    .Y(_04633_));
 sg13g2_nand3_1 _11627_ (.B(net4600),
    .C(_04614_),
    .A(net4602),
    .Y(_04634_));
 sg13g2_nor2_2 _11628_ (.A(_04609_),
    .B(_04634_),
    .Y(_04635_));
 sg13g2_or2_1 _11629_ (.X(_04636_),
    .B(_04631_),
    .A(_04619_));
 sg13g2_nor3_2 _11630_ (.A(net4600),
    .B(net3756),
    .C(_04625_),
    .Y(_04637_));
 sg13g2_nor4_1 _11631_ (.A(_04617_),
    .B(_04621_),
    .C(_04624_),
    .D(_04637_),
    .Y(_04638_));
 sg13g2_nor4_1 _11632_ (.A(_04607_),
    .B(_04627_),
    .C(_04628_),
    .D(_04629_),
    .Y(_04639_));
 sg13g2_nor2_2 _11633_ (.A(net3756),
    .B(_04634_),
    .Y(_04640_));
 sg13g2_nor4_1 _11634_ (.A(_04626_),
    .B(_04632_),
    .C(_04635_),
    .D(_04640_),
    .Y(_04641_));
 sg13g2_nor3_2 _11635_ (.A(net4601),
    .B(_04609_),
    .C(_04618_),
    .Y(_04642_));
 sg13g2_nor4_2 _11636_ (.A(\spiking_network_top_uut.debug_inst.debug_config[2] ),
    .B(\spiking_network_top_uut.debug_inst.debug_config[3] ),
    .C(_04609_),
    .Y(_04643_),
    .D(_04611_));
 sg13g2_nor4_1 _11637_ (.A(_04610_),
    .B(_04630_),
    .C(_04642_),
    .D(_04643_),
    .Y(_04644_));
 sg13g2_nand4_1 _11638_ (.B(_04639_),
    .C(_04641_),
    .A(_04638_),
    .Y(_04645_),
    .D(_04644_));
 sg13g2_nor4_2 _11639_ (.A(net3706),
    .B(_04633_),
    .C(_04636_),
    .Y(_04646_),
    .D(_04645_));
 sg13g2_a22oi_1 _11640_ (.Y(_04647_),
    .B1(_04621_),
    .B2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[0] ),
    .A2(net3706),
    .A1(net4599));
 sg13g2_a22oi_1 _11641_ (.Y(_04648_),
    .B1(_04635_),
    .B2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[0] ),
    .A2(_04626_),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.spike_out ));
 sg13g2_a22oi_1 _11642_ (.Y(_04649_),
    .B1(_04632_),
    .B2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[0] ),
    .A2(_04619_),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[0] ));
 sg13g2_a22oi_1 _11643_ (.Y(_04650_),
    .B1(_04642_),
    .B2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[0] ),
    .A2(_04629_),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[0] ));
 sg13g2_nand4_1 _11644_ (.B(_04648_),
    .C(_04649_),
    .A(_04647_),
    .Y(_04651_),
    .D(_04650_));
 sg13g2_a22oi_1 _11645_ (.Y(_04652_),
    .B1(_04637_),
    .B2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[0] ),
    .A2(_04607_),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[0] ));
 sg13g2_a22oi_1 _11646_ (.Y(_04653_),
    .B1(_04643_),
    .B2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[0] ),
    .A2(_04640_),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[0] ));
 sg13g2_nand2_1 _11647_ (.Y(_04654_),
    .A(_04652_),
    .B(_04653_));
 sg13g2_a22oi_1 _11648_ (.Y(_04655_),
    .B1(_04628_),
    .B2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[0] ),
    .A2(_04624_),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[0] ));
 sg13g2_a22oi_1 _11649_ (.Y(_04656_),
    .B1(_04633_),
    .B2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[0] ),
    .A2(_04617_),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[0] ));
 sg13g2_a22oi_1 _11650_ (.Y(_04657_),
    .B1(_04627_),
    .B2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[0] ),
    .A2(_04610_),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[0] ));
 sg13g2_a22oi_1 _11651_ (.Y(_04658_),
    .B1(_04631_),
    .B2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[0] ),
    .A2(_04630_),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[0] ));
 sg13g2_nand4_1 _11652_ (.B(_04656_),
    .C(_04657_),
    .A(_04655_),
    .Y(_04659_),
    .D(_04658_));
 sg13g2_nor4_1 _11653_ (.A(net3667),
    .B(_04651_),
    .C(_04654_),
    .D(_04659_),
    .Y(_04660_));
 sg13g2_a21oi_2 _11654_ (.B1(_04660_),
    .Y(uo_out[0]),
    .A2(net3667),
    .A1(_03477_));
 sg13g2_a22oi_1 _11655_ (.Y(_04661_),
    .B1(_04621_),
    .B2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ),
    .A2(_04619_),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ));
 sg13g2_a22oi_1 _11656_ (.Y(_04662_),
    .B1(_04626_),
    .B2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.spike_out ),
    .A2(net3706),
    .A1(net4598));
 sg13g2_a22oi_1 _11657_ (.Y(_04663_),
    .B1(_04637_),
    .B2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ),
    .A2(_04628_),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ));
 sg13g2_a22oi_1 _11658_ (.Y(_04664_),
    .B1(_04635_),
    .B2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ),
    .A2(_04610_),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ));
 sg13g2_a22oi_1 _11659_ (.Y(_04665_),
    .B1(_04643_),
    .B2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ),
    .A2(_04632_),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ));
 sg13g2_nand4_1 _11660_ (.B(_04663_),
    .C(_04664_),
    .A(_04662_),
    .Y(_04666_),
    .D(_04665_));
 sg13g2_a22oi_1 _11661_ (.Y(_04667_),
    .B1(_04642_),
    .B2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ),
    .A2(_04617_),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ));
 sg13g2_a22oi_1 _11662_ (.Y(_04668_),
    .B1(_04640_),
    .B2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ),
    .A2(_04633_),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ));
 sg13g2_nand2_1 _11663_ (.Y(_04669_),
    .A(_04667_),
    .B(_04668_));
 sg13g2_a22oi_1 _11664_ (.Y(_04670_),
    .B1(_04629_),
    .B2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ),
    .A2(_04627_),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ));
 sg13g2_a22oi_1 _11665_ (.Y(_04671_),
    .B1(_04624_),
    .B2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ),
    .A2(_04607_),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ));
 sg13g2_a22oi_1 _11666_ (.Y(_04672_),
    .B1(_04631_),
    .B2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ),
    .A2(_04630_),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ));
 sg13g2_nand4_1 _11667_ (.B(_04670_),
    .C(_04671_),
    .A(_04661_),
    .Y(_04673_),
    .D(_04672_));
 sg13g2_nor4_1 _11668_ (.A(net3667),
    .B(_04666_),
    .C(_04669_),
    .D(_04673_),
    .Y(_04674_));
 sg13g2_a21oi_2 _11669_ (.B1(_04674_),
    .Y(uo_out[1]),
    .A2(net3667),
    .A1(_03476_));
 sg13g2_a22oi_1 _11670_ (.Y(_04675_),
    .B1(_04643_),
    .B2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ),
    .A2(net3706),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.spike_out ));
 sg13g2_a22oi_1 _11671_ (.Y(_04676_),
    .B1(_04637_),
    .B2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ),
    .A2(_04628_),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ));
 sg13g2_a22oi_1 _11672_ (.Y(_04677_),
    .B1(_04629_),
    .B2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ),
    .A2(_04619_),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ));
 sg13g2_a22oi_1 _11673_ (.Y(_04678_),
    .B1(_04633_),
    .B2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ),
    .A2(_04631_),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ));
 sg13g2_nand3_1 _11674_ (.B(_04677_),
    .C(_04678_),
    .A(_04676_),
    .Y(_04679_));
 sg13g2_a221oi_1 _11675_ (.B2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ),
    .C1(_04679_),
    .B1(_04627_),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ),
    .Y(_04680_),
    .A2(_04607_));
 sg13g2_nand2_1 _11676_ (.Y(_04681_),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ),
    .B(_04635_));
 sg13g2_a22oi_1 _11677_ (.Y(_04682_),
    .B1(_04640_),
    .B2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ),
    .A2(_04624_),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ));
 sg13g2_a22oi_1 _11678_ (.Y(_04683_),
    .B1(_04632_),
    .B2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ),
    .A2(_04617_),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ));
 sg13g2_a22oi_1 _11679_ (.Y(_04684_),
    .B1(_04630_),
    .B2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ),
    .A2(_04621_),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ));
 sg13g2_nand3_1 _11680_ (.B(_04683_),
    .C(_04684_),
    .A(_04675_),
    .Y(_04685_));
 sg13g2_a221oi_1 _11681_ (.B2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ),
    .C1(_04685_),
    .B1(_04642_),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ),
    .Y(_04686_),
    .A2(_04610_));
 sg13g2_nand4_1 _11682_ (.B(_04681_),
    .C(_04682_),
    .A(_04680_),
    .Y(_04687_),
    .D(_04686_));
 sg13g2_a21o_2 _11683_ (.A2(net3667),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.spike_out ),
    .B1(_04687_),
    .X(uo_out[2]));
 sg13g2_nand2_1 _11684_ (.Y(_04688_),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ),
    .B(_04635_));
 sg13g2_a22oi_1 _11685_ (.Y(_04689_),
    .B1(_04642_),
    .B2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ),
    .A2(_04637_),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ));
 sg13g2_a22oi_1 _11686_ (.Y(_04690_),
    .B1(_04628_),
    .B2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ),
    .A2(_04624_),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ));
 sg13g2_a22oi_1 _11687_ (.Y(_04691_),
    .B1(_04630_),
    .B2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ),
    .A2(_04607_),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ));
 sg13g2_a22oi_1 _11688_ (.Y(_04692_),
    .B1(_04633_),
    .B2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ),
    .A2(_04629_),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ));
 sg13g2_nand4_1 _11689_ (.B(_04690_),
    .C(_04691_),
    .A(_04689_),
    .Y(_04693_),
    .D(_04692_));
 sg13g2_a22oi_1 _11690_ (.Y(_04694_),
    .B1(_04632_),
    .B2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ),
    .A2(net3706),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.spike_out ));
 sg13g2_nand2_1 _11691_ (.Y(_04695_),
    .A(_04688_),
    .B(_04694_));
 sg13g2_a22oi_1 _11692_ (.Y(_04696_),
    .B1(_04631_),
    .B2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ),
    .A2(_04627_),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ));
 sg13g2_a22oi_1 _11693_ (.Y(_04697_),
    .B1(_04621_),
    .B2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ),
    .A2(_04617_),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ));
 sg13g2_a22oi_1 _11694_ (.Y(_04698_),
    .B1(_04619_),
    .B2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ),
    .A2(_04610_),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ));
 sg13g2_a22oi_1 _11695_ (.Y(_04699_),
    .B1(_04643_),
    .B2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ),
    .A2(_04640_),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ));
 sg13g2_nand4_1 _11696_ (.B(_04697_),
    .C(_04698_),
    .A(_04696_),
    .Y(_04700_),
    .D(_04699_));
 sg13g2_nor4_1 _11697_ (.A(net3667),
    .B(_04693_),
    .C(_04695_),
    .D(_04700_),
    .Y(_04701_));
 sg13g2_a21oi_2 _11698_ (.B1(_04701_),
    .Y(uo_out[3]),
    .A2(net3667),
    .A1(_03475_));
 sg13g2_a22oi_1 _11699_ (.Y(_04702_),
    .B1(_04632_),
    .B2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ),
    .A2(_04628_),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ));
 sg13g2_a22oi_1 _11700_ (.Y(_04703_),
    .B1(_04624_),
    .B2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ),
    .A2(_04617_),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ));
 sg13g2_a22oi_1 _11701_ (.Y(_04704_),
    .B1(_04619_),
    .B2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ),
    .A2(net3706),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.spike_out ));
 sg13g2_a22oi_1 _11702_ (.Y(_04705_),
    .B1(_04630_),
    .B2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ),
    .A2(_04610_),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ));
 sg13g2_a22oi_1 _11703_ (.Y(_04706_),
    .B1(_04643_),
    .B2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ),
    .A2(_04627_),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ));
 sg13g2_nand3_1 _11704_ (.B(_04705_),
    .C(_04706_),
    .A(_04703_),
    .Y(_04707_));
 sg13g2_a221oi_1 _11705_ (.B2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ),
    .C1(_04707_),
    .B1(_04637_),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ),
    .Y(_04708_),
    .A2(_04631_));
 sg13g2_nand2_1 _11706_ (.Y(_04709_),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ),
    .B(_04635_));
 sg13g2_a22oi_1 _11707_ (.Y(_04710_),
    .B1(_04640_),
    .B2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ),
    .A2(_04621_),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ));
 sg13g2_a22oi_1 _11708_ (.Y(_04711_),
    .B1(_04642_),
    .B2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ),
    .A2(_04607_),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ));
 sg13g2_nand3_1 _11709_ (.B(_04704_),
    .C(_04711_),
    .A(_04702_),
    .Y(_04712_));
 sg13g2_a221oi_1 _11710_ (.B2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ),
    .C1(_04712_),
    .B1(_04633_),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ),
    .Y(_04713_),
    .A2(_04629_));
 sg13g2_nand4_1 _11711_ (.B(_04709_),
    .C(_04710_),
    .A(_04708_),
    .Y(_04714_),
    .D(_04713_));
 sg13g2_a21o_2 _11712_ (.A2(net3667),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.spike_out ),
    .B1(_04714_),
    .X(uo_out[4]));
 sg13g2_a22oi_1 _11713_ (.Y(_04715_),
    .B1(_04646_),
    .B2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.spike_out ),
    .A2(_04613_),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.spike_out ));
 sg13g2_inv_4 _11714_ (.A(_04715_),
    .Y(uo_out[5]));
 sg13g2_a22oi_1 _11715_ (.Y(_04716_),
    .B1(_04646_),
    .B2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.spike_out ),
    .A2(net3706),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.spike_out ));
 sg13g2_inv_4 _11716_ (.A(_04716_),
    .Y(uo_out[6]));
 sg13g2_a22oi_1 _11717_ (.Y(_04717_),
    .B1(_04646_),
    .B2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.spike_out ),
    .A2(net3706),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.spike_out ));
 sg13g2_inv_4 _11718_ (.A(_04717_),
    .Y(uo_out[7]));
 sg13g2_nor2b_1 _11719_ (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ),
    .B_N(net4287),
    .Y(_04718_));
 sg13g2_xnor2_1 _11720_ (.Y(_04719_),
    .A(net4293),
    .B(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ));
 sg13g2_nor2_1 _11721_ (.A(net4299),
    .B(_03430_),
    .Y(_04720_));
 sg13g2_xnor2_1 _11722_ (.Y(_04721_),
    .A(net4299),
    .B(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ));
 sg13g2_nor2_1 _11723_ (.A(net4306),
    .B(_03431_),
    .Y(_04722_));
 sg13g2_xnor2_1 _11724_ (.Y(_04723_),
    .A(net4306),
    .B(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ));
 sg13g2_nand2_1 _11725_ (.Y(_04724_),
    .A(net4311),
    .B(_03432_));
 sg13g2_a21oi_2 _11726_ (.B1(_04722_),
    .Y(_04725_),
    .A2(_04724_),
    .A1(_04723_));
 sg13g2_nor2b_1 _11727_ (.A(_04725_),
    .B_N(_04721_),
    .Y(_04726_));
 sg13g2_o21ai_1 _11728_ (.B1(_04719_),
    .Y(_04727_),
    .A1(_04720_),
    .A2(_04726_));
 sg13g2_o21ai_1 _11729_ (.B1(_04727_),
    .Y(_04728_),
    .A1(net4293),
    .A2(_03429_));
 sg13g2_o21ai_1 _11730_ (.B1(_04728_),
    .Y(_04729_),
    .A1(net4287),
    .A2(_03428_));
 sg13g2_nand2b_1 _11731_ (.Y(_04730_),
    .B(_04729_),
    .A_N(_04718_));
 sg13g2_and2_1 _11732_ (.A(net4574),
    .B(net3634),
    .X(_00017_));
 sg13g2_nor2b_1 _11733_ (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ),
    .B_N(net4287),
    .Y(_04731_));
 sg13g2_xnor2_1 _11734_ (.Y(_04732_),
    .A(net4293),
    .B(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ));
 sg13g2_nor2_1 _11735_ (.A(net4299),
    .B(_03410_),
    .Y(_04733_));
 sg13g2_xnor2_1 _11736_ (.Y(_04734_),
    .A(net4299),
    .B(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ));
 sg13g2_nor2_1 _11737_ (.A(net4306),
    .B(_03408_),
    .Y(_04735_));
 sg13g2_xnor2_1 _11738_ (.Y(_04736_),
    .A(net4306),
    .B(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ));
 sg13g2_nand2_1 _11739_ (.Y(_04737_),
    .A(net4311),
    .B(_03407_));
 sg13g2_a21oi_1 _11740_ (.A1(_04736_),
    .A2(_04737_),
    .Y(_04738_),
    .B1(_04735_));
 sg13g2_nor2b_1 _11741_ (.A(_04738_),
    .B_N(_04734_),
    .Y(_04739_));
 sg13g2_o21ai_1 _11742_ (.B1(_04732_),
    .Y(_04740_),
    .A1(_04733_),
    .A2(_04739_));
 sg13g2_o21ai_1 _11743_ (.B1(_04740_),
    .Y(_04741_),
    .A1(net4293),
    .A2(_03409_));
 sg13g2_o21ai_1 _11744_ (.B1(_04741_),
    .Y(_04742_),
    .A1(net4287),
    .A2(_03411_));
 sg13g2_nand2b_1 _11745_ (.Y(_04743_),
    .B(_04742_),
    .A_N(_04731_));
 sg13g2_and2_1 _11746_ (.A(net4574),
    .B(net3631),
    .X(_00018_));
 sg13g2_nand2b_1 _11747_ (.Y(_04744_),
    .B(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ),
    .A_N(net4289));
 sg13g2_nor2b_1 _11748_ (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ),
    .B_N(net4289),
    .Y(_04745_));
 sg13g2_xnor2_1 _11749_ (.Y(_04746_),
    .A(net4295),
    .B(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ));
 sg13g2_nor2_1 _11750_ (.A(net4303),
    .B(_03437_),
    .Y(_04747_));
 sg13g2_xnor2_1 _11751_ (.Y(_04748_),
    .A(net4303),
    .B(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ));
 sg13g2_nor2_1 _11752_ (.A(net4309),
    .B(_03438_),
    .Y(_04749_));
 sg13g2_xnor2_1 _11753_ (.Y(_04750_),
    .A(net4309),
    .B(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ));
 sg13g2_nand2b_1 _11754_ (.Y(_04751_),
    .B(net4315),
    .A_N(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[0] ));
 sg13g2_a21oi_1 _11755_ (.A1(_04750_),
    .A2(_04751_),
    .Y(_04752_),
    .B1(_04749_));
 sg13g2_nor2b_1 _11756_ (.A(_04752_),
    .B_N(_04748_),
    .Y(_04753_));
 sg13g2_o21ai_1 _11757_ (.B1(_04746_),
    .Y(_04754_),
    .A1(_04747_),
    .A2(_04753_));
 sg13g2_o21ai_1 _11758_ (.B1(_04754_),
    .Y(_04755_),
    .A1(net4295),
    .A2(_03436_));
 sg13g2_a21o_1 _11759_ (.A2(_04755_),
    .A1(_04744_),
    .B1(_04745_),
    .X(_04756_));
 sg13g2_inv_1 _11760_ (.Y(_04757_),
    .A(net3661));
 sg13g2_nor2_2 _11761_ (.A(net3930),
    .B(_04757_),
    .Y(_00009_));
 sg13g2_nor2_1 _11762_ (.A(net4288),
    .B(_03439_),
    .Y(_04758_));
 sg13g2_nand2_1 _11763_ (.Y(_04759_),
    .A(net4288),
    .B(_03439_));
 sg13g2_nand2b_1 _11764_ (.Y(_04760_),
    .B(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ),
    .A_N(net4294));
 sg13g2_xnor2_1 _11765_ (.Y(_04761_),
    .A(net4294),
    .B(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ));
 sg13g2_nor2_1 _11766_ (.A(net4300),
    .B(_03441_),
    .Y(_04762_));
 sg13g2_xnor2_1 _11767_ (.Y(_04763_),
    .A(net4299),
    .B(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ));
 sg13g2_nor2b_1 _11768_ (.A(net4308),
    .B_N(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ),
    .Y(_04764_));
 sg13g2_xnor2_1 _11769_ (.Y(_04765_),
    .A(net4308),
    .B(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ));
 sg13g2_nand2b_1 _11770_ (.Y(_04766_),
    .B(net4312),
    .A_N(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[0] ));
 sg13g2_a21oi_2 _11771_ (.B1(_04764_),
    .Y(_04767_),
    .A2(_04766_),
    .A1(_04765_));
 sg13g2_nor2b_1 _11772_ (.A(_04767_),
    .B_N(_04763_),
    .Y(_04768_));
 sg13g2_o21ai_1 _11773_ (.B1(_04761_),
    .Y(_04769_),
    .A1(_04762_),
    .A2(_04768_));
 sg13g2_and2_1 _11774_ (.A(_04760_),
    .B(_04769_),
    .X(_04770_));
 sg13g2_o21ai_1 _11775_ (.B1(_04759_),
    .Y(_04771_),
    .A1(_04758_),
    .A2(_04770_));
 sg13g2_inv_2 _11776_ (.Y(_04772_),
    .A(net3666));
 sg13g2_nor2_2 _11777_ (.A(net3920),
    .B(_04772_),
    .Y(_00010_));
 sg13g2_nor2_1 _11778_ (.A(net4289),
    .B(_03442_),
    .Y(_04773_));
 sg13g2_nand2_1 _11779_ (.Y(_04774_),
    .A(net4289),
    .B(_03442_));
 sg13g2_nand2b_1 _11780_ (.Y(_04775_),
    .B(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ),
    .A_N(net4295));
 sg13g2_xnor2_1 _11781_ (.Y(_04776_),
    .A(net4295),
    .B(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ));
 sg13g2_nor2_1 _11782_ (.A(net4300),
    .B(_03443_),
    .Y(_04777_));
 sg13g2_xnor2_1 _11783_ (.Y(_04778_),
    .A(net4299),
    .B(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ));
 sg13g2_nor2b_1 _11784_ (.A(net4309),
    .B_N(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ),
    .Y(_04779_));
 sg13g2_nand2_1 _11785_ (.Y(_04780_),
    .A(net4311),
    .B(_03444_));
 sg13g2_xnor2_1 _11786_ (.Y(_04781_),
    .A(net4309),
    .B(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ));
 sg13g2_a21oi_1 _11787_ (.A1(_04780_),
    .A2(_04781_),
    .Y(_04782_),
    .B1(_04779_));
 sg13g2_nor2b_1 _11788_ (.A(_04782_),
    .B_N(_04778_),
    .Y(_04783_));
 sg13g2_o21ai_1 _11789_ (.B1(_04776_),
    .Y(_04784_),
    .A1(_04777_),
    .A2(_04783_));
 sg13g2_and2_1 _11790_ (.A(_04775_),
    .B(_04784_),
    .X(_04785_));
 sg13g2_o21ai_1 _11791_ (.B1(_04774_),
    .Y(_04786_),
    .A1(_04773_),
    .A2(_04785_));
 sg13g2_inv_1 _11792_ (.Y(_04787_),
    .A(net3658));
 sg13g2_nor2_2 _11793_ (.A(net3929),
    .B(_04787_),
    .Y(_00011_));
 sg13g2_nand2b_1 _11794_ (.Y(_04788_),
    .B(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ),
    .A_N(net4287));
 sg13g2_nor2b_1 _11795_ (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ),
    .B_N(net4287),
    .Y(_04789_));
 sg13g2_xnor2_1 _11796_ (.Y(_04790_),
    .A(net4293),
    .B(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ));
 sg13g2_nor2_1 _11797_ (.A(net4299),
    .B(_03447_),
    .Y(_04791_));
 sg13g2_xnor2_1 _11798_ (.Y(_04792_),
    .A(net4299),
    .B(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ));
 sg13g2_nor2_1 _11799_ (.A(net4306),
    .B(_03448_),
    .Y(_04793_));
 sg13g2_xnor2_1 _11800_ (.Y(_04794_),
    .A(net4306),
    .B(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ));
 sg13g2_nand2b_1 _11801_ (.Y(_04795_),
    .B(net4311),
    .A_N(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[0] ));
 sg13g2_a21oi_2 _11802_ (.B1(_04793_),
    .Y(_04796_),
    .A2(_04795_),
    .A1(_04794_));
 sg13g2_nor2b_1 _11803_ (.A(_04796_),
    .B_N(_04792_),
    .Y(_04797_));
 sg13g2_o21ai_1 _11804_ (.B1(_04790_),
    .Y(_04798_),
    .A1(_04791_),
    .A2(_04797_));
 sg13g2_o21ai_1 _11805_ (.B1(_04798_),
    .Y(_04799_),
    .A1(net4293),
    .A2(_03446_));
 sg13g2_a21o_1 _11806_ (.A2(_04799_),
    .A1(_04788_),
    .B1(_04789_),
    .X(_04800_));
 sg13g2_and2_1 _11807_ (.A(net4531),
    .B(net3655),
    .X(_00012_));
 sg13g2_nand2b_1 _11808_ (.Y(_04801_),
    .B(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ),
    .A_N(net4288));
 sg13g2_nor2b_1 _11809_ (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ),
    .B_N(net4291),
    .Y(_04802_));
 sg13g2_xnor2_1 _11810_ (.Y(_04803_),
    .A(net4297),
    .B(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ));
 sg13g2_nor2_1 _11811_ (.A(net4301),
    .B(_03415_),
    .Y(_04804_));
 sg13g2_xnor2_1 _11812_ (.Y(_04805_),
    .A(net4301),
    .B(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ));
 sg13g2_nor2_1 _11813_ (.A(net4307),
    .B(_03416_),
    .Y(_04806_));
 sg13g2_xnor2_1 _11814_ (.Y(_04807_),
    .A(net4307),
    .B(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ));
 sg13g2_nand2_1 _11815_ (.Y(_04808_),
    .A(net4313),
    .B(_03417_));
 sg13g2_a21oi_1 _11816_ (.A1(_04807_),
    .A2(_04808_),
    .Y(_04809_),
    .B1(_04806_));
 sg13g2_nor2b_1 _11817_ (.A(_04809_),
    .B_N(_04805_),
    .Y(_04810_));
 sg13g2_o21ai_1 _11818_ (.B1(_04803_),
    .Y(_04811_),
    .A1(_04804_),
    .A2(_04810_));
 sg13g2_o21ai_1 _11819_ (.B1(_04811_),
    .Y(_04812_),
    .A1(net4294),
    .A2(_03414_));
 sg13g2_a21o_1 _11820_ (.A2(_04812_),
    .A1(_04801_),
    .B1(_04802_),
    .X(_04813_));
 sg13g2_and2_2 _11821_ (.A(net4531),
    .B(_04813_),
    .X(_00013_));
 sg13g2_nor2_1 _11822_ (.A(net4290),
    .B(_03419_),
    .Y(_04814_));
 sg13g2_nand2_1 _11823_ (.Y(_04815_),
    .A(net4290),
    .B(_03419_));
 sg13g2_nand2b_1 _11824_ (.Y(_04816_),
    .B(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ),
    .A_N(net4296));
 sg13g2_xnor2_1 _11825_ (.Y(_04817_),
    .A(net4296),
    .B(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ));
 sg13g2_nor2b_1 _11826_ (.A(net4302),
    .B_N(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ),
    .Y(_04818_));
 sg13g2_nor2_1 _11827_ (.A(net4308),
    .B(_03420_),
    .Y(_04819_));
 sg13g2_xnor2_1 _11828_ (.Y(_04820_),
    .A(net4308),
    .B(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ));
 sg13g2_nand2b_1 _11829_ (.Y(_04821_),
    .B(net4314),
    .A_N(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[0] ));
 sg13g2_a21oi_1 _11830_ (.A1(_04820_),
    .A2(_04821_),
    .Y(_04822_),
    .B1(_04819_));
 sg13g2_xor2_1 _11831_ (.B(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ),
    .A(net4302),
    .X(_04823_));
 sg13g2_nor2_1 _11832_ (.A(_04822_),
    .B(_04823_),
    .Y(_04824_));
 sg13g2_o21ai_1 _11833_ (.B1(_04817_),
    .Y(_04825_),
    .A1(_04818_),
    .A2(_04824_));
 sg13g2_and2_1 _11834_ (.A(_04816_),
    .B(_04825_),
    .X(_04826_));
 sg13g2_o21ai_1 _11835_ (.B1(_04815_),
    .Y(_04827_),
    .A1(_04814_),
    .A2(_04826_));
 sg13g2_inv_1 _11836_ (.Y(_04828_),
    .A(net3650));
 sg13g2_nor2_2 _11837_ (.A(net3927),
    .B(_04828_),
    .Y(_00014_));
 sg13g2_nor2b_1 _11838_ (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ),
    .B_N(net4287),
    .Y(_04829_));
 sg13g2_xnor2_1 _11839_ (.Y(_04830_),
    .A(net4294),
    .B(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ));
 sg13g2_nor2b_1 _11840_ (.A(net4300),
    .B_N(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ),
    .Y(_04831_));
 sg13g2_xnor2_1 _11841_ (.Y(_04832_),
    .A(net4300),
    .B(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ));
 sg13g2_nor2_1 _11842_ (.A(net4306),
    .B(_03423_),
    .Y(_04833_));
 sg13g2_xnor2_1 _11843_ (.Y(_04834_),
    .A(net4306),
    .B(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ));
 sg13g2_nand2b_1 _11844_ (.Y(_04835_),
    .B(net4312),
    .A_N(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[0] ));
 sg13g2_a21oi_1 _11845_ (.A1(_04834_),
    .A2(_04835_),
    .Y(_04836_),
    .B1(_04833_));
 sg13g2_nor2b_1 _11846_ (.A(_04836_),
    .B_N(_04832_),
    .Y(_04837_));
 sg13g2_o21ai_1 _11847_ (.B1(_04830_),
    .Y(_04838_),
    .A1(_04831_),
    .A2(_04837_));
 sg13g2_o21ai_1 _11848_ (.B1(_04838_),
    .Y(_04839_),
    .A1(net4293),
    .A2(_03422_));
 sg13g2_o21ai_1 _11849_ (.B1(_04839_),
    .Y(_04840_),
    .A1(net4287),
    .A2(_03421_));
 sg13g2_nand2b_1 _11850_ (.Y(_04841_),
    .B(_04840_),
    .A_N(_04829_));
 sg13g2_and2_2 _11851_ (.A(net4530),
    .B(net3628),
    .X(_00015_));
 sg13g2_nor2b_1 _11852_ (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ),
    .B_N(net4292),
    .Y(_04842_));
 sg13g2_xnor2_1 _11853_ (.Y(_04843_),
    .A(net4298),
    .B(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ));
 sg13g2_nor2_1 _11854_ (.A(net4304),
    .B(_03426_),
    .Y(_04844_));
 sg13g2_xnor2_1 _11855_ (.Y(_04845_),
    .A(net4304),
    .B(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ));
 sg13g2_nor2b_1 _11856_ (.A(net4310),
    .B_N(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ),
    .Y(_04846_));
 sg13g2_nand2_1 _11857_ (.Y(_04847_),
    .A(\spiking_network_top_uut.all_data_out[16] ),
    .B(_03427_));
 sg13g2_xnor2_1 _11858_ (.Y(_04848_),
    .A(net4310),
    .B(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ));
 sg13g2_a21oi_1 _11859_ (.A1(_04847_),
    .A2(_04848_),
    .Y(_04849_),
    .B1(_04846_));
 sg13g2_nor2b_1 _11860_ (.A(_04849_),
    .B_N(_04845_),
    .Y(_04850_));
 sg13g2_o21ai_1 _11861_ (.B1(_04843_),
    .Y(_04851_),
    .A1(_04844_),
    .A2(_04850_));
 sg13g2_o21ai_1 _11862_ (.B1(_04851_),
    .Y(_04852_),
    .A1(net4298),
    .A2(_03425_));
 sg13g2_o21ai_1 _11863_ (.B1(_04852_),
    .Y(_04853_),
    .A1(net4292),
    .A2(_03424_));
 sg13g2_nand2b_1 _11864_ (.Y(_04854_),
    .B(_04853_),
    .A_N(_04842_));
 sg13g2_and2_1 _11865_ (.A(net4533),
    .B(net3625),
    .X(_00016_));
 sg13g2_nor2b_1 _11866_ (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ),
    .B_N(net4292),
    .Y(_04855_));
 sg13g2_xnor2_1 _11867_ (.Y(_04856_),
    .A(net4298),
    .B(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ));
 sg13g2_nor2b_1 _11868_ (.A(net4305),
    .B_N(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ),
    .Y(_04857_));
 sg13g2_nor2b_1 _11869_ (.A(net4310),
    .B_N(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ),
    .Y(_04858_));
 sg13g2_nand2b_1 _11870_ (.Y(_04859_),
    .B(net4316),
    .A_N(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[0] ));
 sg13g2_xnor2_1 _11871_ (.Y(_04860_),
    .A(net4310),
    .B(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ));
 sg13g2_a21oi_1 _11872_ (.A1(_04859_),
    .A2(_04860_),
    .Y(_04861_),
    .B1(_04858_));
 sg13g2_xnor2_1 _11873_ (.Y(_04862_),
    .A(net4305),
    .B(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ));
 sg13g2_nor2b_1 _11874_ (.A(_04861_),
    .B_N(_04862_),
    .Y(_04863_));
 sg13g2_o21ai_1 _11875_ (.B1(_04856_),
    .Y(_04864_),
    .A1(_04857_),
    .A2(_04863_));
 sg13g2_o21ai_1 _11876_ (.B1(_04864_),
    .Y(_04865_),
    .A1(net4298),
    .A2(_03400_));
 sg13g2_o21ai_1 _11877_ (.B1(_04865_),
    .Y(_04866_),
    .A1(net4292),
    .A2(_03399_));
 sg13g2_nand2b_1 _11878_ (.Y(_04867_),
    .B(_04866_),
    .A_N(_04855_));
 sg13g2_and2_2 _11879_ (.A(net4606),
    .B(net3647),
    .X(_00001_));
 sg13g2_nor2b_1 _11880_ (.A(net4289),
    .B_N(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ),
    .Y(_04868_));
 sg13g2_nand2b_1 _11881_ (.Y(_04869_),
    .B(net4289),
    .A_N(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ));
 sg13g2_nand2b_1 _11882_ (.Y(_04870_),
    .B(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ),
    .A_N(net4296));
 sg13g2_xnor2_1 _11883_ (.Y(_04871_),
    .A(net4296),
    .B(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ));
 sg13g2_nor2_1 _11884_ (.A(net4303),
    .B(_03404_),
    .Y(_04872_));
 sg13g2_xor2_1 _11885_ (.B(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ),
    .A(net4303),
    .X(_04873_));
 sg13g2_nand2_1 _11886_ (.Y(_04874_),
    .A(_03401_),
    .B(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ));
 sg13g2_nor2b_1 _11887_ (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[0] ),
    .B_N(net4315),
    .Y(_04875_));
 sg13g2_xor2_1 _11888_ (.B(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ),
    .A(net4309),
    .X(_04876_));
 sg13g2_or2_1 _11889_ (.X(_04877_),
    .B(_04876_),
    .A(_04875_));
 sg13g2_a21oi_1 _11890_ (.A1(_04874_),
    .A2(_04877_),
    .Y(_04878_),
    .B1(_04873_));
 sg13g2_o21ai_1 _11891_ (.B1(_04871_),
    .Y(_04879_),
    .A1(_04872_),
    .A2(_04878_));
 sg13g2_and2_1 _11892_ (.A(_04870_),
    .B(_04879_),
    .X(_04880_));
 sg13g2_o21ai_1 _11893_ (.B1(_04869_),
    .Y(_04881_),
    .A1(_04868_),
    .A2(_04880_));
 sg13g2_and2_2 _11894_ (.A(net4605),
    .B(net3664),
    .X(_00002_));
 sg13g2_nor2b_1 _11895_ (.A(net477),
    .B_N(net4289),
    .Y(_04882_));
 sg13g2_xnor2_1 _11896_ (.Y(_04883_),
    .A(net4295),
    .B(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ));
 sg13g2_nor2b_1 _11897_ (.A(net4303),
    .B_N(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ),
    .Y(_04884_));
 sg13g2_xor2_1 _11898_ (.B(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ),
    .A(net4309),
    .X(_04885_));
 sg13g2_nor2b_1 _11899_ (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[0] ),
    .B_N(net4315),
    .Y(_04886_));
 sg13g2_nor2_1 _11900_ (.A(_04885_),
    .B(_04886_),
    .Y(_04887_));
 sg13g2_a21oi_1 _11901_ (.A1(_03401_),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ),
    .Y(_04888_),
    .B1(_04887_));
 sg13g2_xnor2_1 _11902_ (.Y(_04889_),
    .A(net4303),
    .B(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ));
 sg13g2_nor2b_1 _11903_ (.A(_04888_),
    .B_N(_04889_),
    .Y(_04890_));
 sg13g2_o21ai_1 _11904_ (.B1(_04883_),
    .Y(_04891_),
    .A1(_04884_),
    .A2(_04890_));
 sg13g2_o21ai_1 _11905_ (.B1(_04891_),
    .Y(_04892_),
    .A1(net4295),
    .A2(_03467_));
 sg13g2_o21ai_1 _11906_ (.B1(_04892_),
    .Y(_04893_),
    .A1(net4289),
    .A2(_03466_));
 sg13g2_nand2b_1 _11907_ (.Y(_04894_),
    .B(_04893_),
    .A_N(_04882_));
 sg13g2_and2_2 _11908_ (.A(net4606),
    .B(net3622),
    .X(_00003_));
 sg13g2_nor2b_1 _11909_ (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ),
    .B_N(net4288),
    .Y(_04895_));
 sg13g2_xnor2_1 _11910_ (.Y(_04896_),
    .A(net4294),
    .B(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ));
 sg13g2_nor2_1 _11911_ (.A(net4301),
    .B(_03451_),
    .Y(_04897_));
 sg13g2_xnor2_1 _11912_ (.Y(_04898_),
    .A(net4301),
    .B(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ));
 sg13g2_nor2_1 _11913_ (.A(net4307),
    .B(_03452_),
    .Y(_04899_));
 sg13g2_xnor2_1 _11914_ (.Y(_04900_),
    .A(net4307),
    .B(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ));
 sg13g2_nand2_1 _11915_ (.Y(_04901_),
    .A(net4313),
    .B(_03453_));
 sg13g2_a21oi_1 _11916_ (.A1(_04900_),
    .A2(_04901_),
    .Y(_04902_),
    .B1(_04899_));
 sg13g2_nor2b_1 _11917_ (.A(_04902_),
    .B_N(_04898_),
    .Y(_04903_));
 sg13g2_o21ai_1 _11918_ (.B1(_04896_),
    .Y(_04904_),
    .A1(_04897_),
    .A2(_04903_));
 sg13g2_o21ai_1 _11919_ (.B1(_04904_),
    .Y(_04905_),
    .A1(net4294),
    .A2(_03450_));
 sg13g2_o21ai_1 _11920_ (.B1(_04905_),
    .Y(_04906_),
    .A1(net4288),
    .A2(_03449_));
 sg13g2_nand2b_1 _11921_ (.Y(_04907_),
    .B(_04906_),
    .A_N(_04895_));
 sg13g2_and2_1 _11922_ (.A(net4604),
    .B(net3619),
    .X(_00004_));
 sg13g2_nor2_1 _11923_ (.A(net4292),
    .B(_03454_),
    .Y(_04908_));
 sg13g2_nand2_1 _11924_ (.Y(_04909_),
    .A(net4292),
    .B(_03454_));
 sg13g2_nand2b_1 _11925_ (.Y(_04910_),
    .B(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ),
    .A_N(net4298));
 sg13g2_xnor2_1 _11926_ (.Y(_04911_),
    .A(net4298),
    .B(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ));
 sg13g2_nor2_1 _11927_ (.A(net4305),
    .B(_03456_),
    .Y(_04912_));
 sg13g2_xnor2_1 _11928_ (.Y(_04913_),
    .A(net4305),
    .B(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ));
 sg13g2_nor2_1 _11929_ (.A(net4310),
    .B(_03457_),
    .Y(_04914_));
 sg13g2_xnor2_1 _11930_ (.Y(_04915_),
    .A(net4310),
    .B(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ));
 sg13g2_nand2_1 _11931_ (.Y(_04916_),
    .A(net4316),
    .B(_03458_));
 sg13g2_a21oi_1 _11932_ (.A1(_04915_),
    .A2(_04916_),
    .Y(_04917_),
    .B1(_04914_));
 sg13g2_nor2b_1 _11933_ (.A(_04917_),
    .B_N(_04913_),
    .Y(_04918_));
 sg13g2_o21ai_1 _11934_ (.B1(_04911_),
    .Y(_04919_),
    .A1(_04912_),
    .A2(_04918_));
 sg13g2_and2_1 _11935_ (.A(_04910_),
    .B(_04919_),
    .X(_04920_));
 sg13g2_o21ai_1 _11936_ (.B1(_04909_),
    .Y(_04921_),
    .A1(_04908_),
    .A2(_04920_));
 sg13g2_inv_1 _11937_ (.Y(_04922_),
    .A(net3645));
 sg13g2_nor2_1 _11938_ (.A(net3958),
    .B(_04922_),
    .Y(_00005_));
 sg13g2_nor2_1 _11939_ (.A(net4291),
    .B(_03459_),
    .Y(_04923_));
 sg13g2_nand2_1 _11940_ (.Y(_04924_),
    .A(net4291),
    .B(_03459_));
 sg13g2_nand2b_1 _11941_ (.Y(_04925_),
    .B(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ),
    .A_N(net4297));
 sg13g2_xnor2_1 _11942_ (.Y(_04926_),
    .A(net4297),
    .B(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ));
 sg13g2_nor2_1 _11943_ (.A(net4301),
    .B(_03460_),
    .Y(_04927_));
 sg13g2_xnor2_1 _11944_ (.Y(_04928_),
    .A(net4301),
    .B(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ));
 sg13g2_nor2_1 _11945_ (.A(net4307),
    .B(_03461_),
    .Y(_04929_));
 sg13g2_xnor2_1 _11946_ (.Y(_04930_),
    .A(net4307),
    .B(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ));
 sg13g2_nand2b_1 _11947_ (.Y(_04931_),
    .B(net4313),
    .A_N(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[0] ));
 sg13g2_a21oi_1 _11948_ (.A1(_04930_),
    .A2(_04931_),
    .Y(_04932_),
    .B1(_04929_));
 sg13g2_nor2b_1 _11949_ (.A(_04932_),
    .B_N(_04928_),
    .Y(_04933_));
 sg13g2_o21ai_1 _11950_ (.B1(_04926_),
    .Y(_04934_),
    .A1(_04927_),
    .A2(_04933_));
 sg13g2_and2_1 _11951_ (.A(_04925_),
    .B(_04934_),
    .X(_04935_));
 sg13g2_o21ai_1 _11952_ (.B1(_04924_),
    .Y(_04936_),
    .A1(_04923_),
    .A2(_04935_));
 sg13g2_inv_1 _11953_ (.Y(_04937_),
    .A(net3642));
 sg13g2_nor2_2 _11954_ (.A(net3947),
    .B(_04937_),
    .Y(_00006_));
 sg13g2_nor2_1 _11955_ (.A(net4288),
    .B(_03462_),
    .Y(_04938_));
 sg13g2_nand2_1 _11956_ (.Y(_04939_),
    .A(net4288),
    .B(_03462_));
 sg13g2_nand2b_1 _11957_ (.Y(_04940_),
    .B(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ),
    .A_N(net4294));
 sg13g2_xnor2_1 _11958_ (.Y(_04941_),
    .A(net4293),
    .B(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ));
 sg13g2_nor2b_1 _11959_ (.A(net4301),
    .B_N(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ),
    .Y(_04942_));
 sg13g2_nor2_1 _11960_ (.A(net4307),
    .B(_03464_),
    .Y(_04943_));
 sg13g2_xnor2_1 _11961_ (.Y(_04944_),
    .A(net4307),
    .B(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ));
 sg13g2_nand2_1 _11962_ (.Y(_04945_),
    .A(net4313),
    .B(_03465_));
 sg13g2_a21oi_1 _11963_ (.A1(_04944_),
    .A2(_04945_),
    .Y(_04946_),
    .B1(_04943_));
 sg13g2_xor2_1 _11964_ (.B(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ),
    .A(net4301),
    .X(_04947_));
 sg13g2_nor2_1 _11965_ (.A(_04946_),
    .B(_04947_),
    .Y(_04948_));
 sg13g2_o21ai_1 _11966_ (.B1(_04941_),
    .Y(_04949_),
    .A1(_04942_),
    .A2(_04948_));
 sg13g2_and2_1 _11967_ (.A(_04940_),
    .B(_04949_),
    .X(_04950_));
 sg13g2_o21ai_1 _11968_ (.B1(_04939_),
    .Y(_04951_),
    .A1(_04938_),
    .A2(_04950_));
 sg13g2_inv_1 _11969_ (.Y(_04952_),
    .A(net3639));
 sg13g2_nor2_2 _11970_ (.A(net3948),
    .B(_04952_),
    .Y(_00007_));
 sg13g2_nor2_1 _11971_ (.A(net4290),
    .B(_03433_),
    .Y(_04953_));
 sg13g2_nand2_1 _11972_ (.Y(_04954_),
    .A(net4290),
    .B(_03433_));
 sg13g2_nand2b_1 _11973_ (.Y(_04955_),
    .B(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ),
    .A_N(net4295));
 sg13g2_xnor2_1 _11974_ (.Y(_04956_),
    .A(net4295),
    .B(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ));
 sg13g2_nor2_1 _11975_ (.A(net4303),
    .B(_03434_),
    .Y(_04957_));
 sg13g2_xnor2_1 _11976_ (.Y(_04958_),
    .A(net4303),
    .B(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ));
 sg13g2_xnor2_1 _11977_ (.Y(_04959_),
    .A(net4309),
    .B(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ));
 sg13g2_nor2b_1 _11978_ (.A(net447),
    .B_N(net4315),
    .Y(_04960_));
 sg13g2_nor2b_1 _11979_ (.A(_04960_),
    .B_N(_04959_),
    .Y(_04961_));
 sg13g2_a21oi_1 _11980_ (.A1(_03401_),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ),
    .Y(_04962_),
    .B1(_04961_));
 sg13g2_nor2b_1 _11981_ (.A(_04962_),
    .B_N(_04958_),
    .Y(_04963_));
 sg13g2_o21ai_1 _11982_ (.B1(_04956_),
    .Y(_04964_),
    .A1(_04957_),
    .A2(_04963_));
 sg13g2_and2_1 _11983_ (.A(_04955_),
    .B(_04964_),
    .X(_04965_));
 sg13g2_o21ai_1 _11984_ (.B1(_04954_),
    .Y(_04966_),
    .A1(_04953_),
    .A2(_04965_));
 sg13g2_inv_2 _11985_ (.Y(_04967_),
    .A(net3636));
 sg13g2_nor2_2 _11986_ (.A(net3952),
    .B(_04967_),
    .Y(_00008_));
 sg13g2_nand2b_1 _11987_ (.Y(_04968_),
    .B(_00028_),
    .A_N(\spiking_network_top_uut.spi_inst.spi_control_unit_inst.current_state[0] ));
 sg13g2_nor3_2 _11988_ (.A(_03469_),
    .B(_00029_),
    .C(_04968_),
    .Y(_00019_));
 sg13g2_nor2_2 _11989_ (.A(_03699_),
    .B(_03700_),
    .Y(_04969_));
 sg13g2_nor2_1 _11990_ (.A(\spiking_network_top_uut.spi_inst.spi_control_unit_inst.current_state[1] ),
    .B(\spiking_network_top_uut.spi_inst.spi_control_unit_inst.current_state[0] ),
    .Y(_04970_));
 sg13g2_and2_1 _11991_ (.A(\spiking_network_top_uut.spi_inst.spi_control_unit_inst.current_state[2] ),
    .B(_04970_),
    .X(_04971_));
 sg13g2_nand2_1 _11992_ (.Y(_04972_),
    .A(\spiking_network_top_uut.spi_inst.spi_control_unit_inst.current_state[2] ),
    .B(_04970_));
 sg13g2_nor3_2 _11993_ (.A(_00029_),
    .B(_04969_),
    .C(_04972_),
    .Y(_00021_));
 sg13g2_or2_1 _11994_ (.X(output_ready),
    .B(\spiking_network_top_uut.output_data_ready ),
    .A(\spiking_network_top_uut.data_valid_out ));
 sg13g2_a22oi_1 _11995_ (.Y(_04973_),
    .B1(_03881_),
    .B2(net11),
    .A2(net3722),
    .A1(\spiking_network_top_uut.spi_inst.spi_slave_inst.shift_reg[0] ));
 sg13g2_inv_1 _11996_ (.Y(_00425_),
    .A(_04973_));
 sg13g2_a22oi_1 _11997_ (.Y(_04974_),
    .B1(_03881_),
    .B2(\spiking_network_top_uut.spi_inst.spi_slave_inst.shift_reg[0] ),
    .A2(net3720),
    .A1(\spiking_network_top_uut.spi_inst.spi_slave_inst.shift_reg[1] ));
 sg13g2_inv_1 _11998_ (.Y(_00426_),
    .A(_04974_));
 sg13g2_a22oi_1 _11999_ (.Y(_04975_),
    .B1(_03881_),
    .B2(\spiking_network_top_uut.spi_inst.spi_slave_inst.shift_reg[1] ),
    .A2(net3720),
    .A1(\spiking_network_top_uut.spi_inst.spi_slave_inst.shift_reg[2] ));
 sg13g2_inv_1 _12000_ (.Y(_00427_),
    .A(_04975_));
 sg13g2_a22oi_1 _12001_ (.Y(_04976_),
    .B1(_03881_),
    .B2(\spiking_network_top_uut.spi_inst.spi_slave_inst.shift_reg[2] ),
    .A2(net3721),
    .A1(\spiking_network_top_uut.spi_inst.spi_slave_inst.shift_reg[3] ));
 sg13g2_inv_1 _12002_ (.Y(_00428_),
    .A(_04976_));
 sg13g2_a22oi_1 _12003_ (.Y(_04977_),
    .B1(_03881_),
    .B2(\spiking_network_top_uut.spi_inst.spi_slave_inst.shift_reg[3] ),
    .A2(net3721),
    .A1(\spiking_network_top_uut.spi_inst.spi_slave_inst.shift_reg[4] ));
 sg13g2_inv_1 _12004_ (.Y(_00429_),
    .A(_04977_));
 sg13g2_a22oi_1 _12005_ (.Y(_04978_),
    .B1(_03881_),
    .B2(\spiking_network_top_uut.spi_inst.spi_slave_inst.shift_reg[4] ),
    .A2(net3721),
    .A1(\spiking_network_top_uut.spi_inst.spi_slave_inst.shift_reg[5] ));
 sg13g2_inv_1 _12006_ (.Y(_00430_),
    .A(_04978_));
 sg13g2_a22oi_1 _12007_ (.Y(_04979_),
    .B1(_03881_),
    .B2(\spiking_network_top_uut.spi_inst.spi_slave_inst.shift_reg[5] ),
    .A2(net3720),
    .A1(\spiking_network_top_uut.spi_inst.spi_slave_inst.shift_reg[6] ));
 sg13g2_inv_1 _12008_ (.Y(_00431_),
    .A(_04979_));
 sg13g2_mux4_1 _12009_ (.S0(\spiking_network_top_uut.all_data_out[860] ),
    .A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[0] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[1] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[2] ),
    .A3(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[3] ),
    .S1(\spiking_network_top_uut.all_data_out[861] ),
    .X(_04980_));
 sg13g2_mux2_1 _12010_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[6] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[7] ),
    .S(\spiking_network_top_uut.all_data_out[860] ),
    .X(_04981_));
 sg13g2_nor2b_1 _12011_ (.A(\spiking_network_top_uut.all_data_out[860] ),
    .B_N(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[4] ),
    .Y(_04982_));
 sg13g2_a21oi_1 _12012_ (.A1(\spiking_network_top_uut.all_data_out[860] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[5] ),
    .Y(_04983_),
    .B1(_04982_));
 sg13g2_o21ai_1 _12013_ (.B1(\spiking_network_top_uut.all_data_out[862] ),
    .Y(_04984_),
    .A1(\spiking_network_top_uut.all_data_out[861] ),
    .A2(_04983_));
 sg13g2_a21oi_1 _12014_ (.A1(\spiking_network_top_uut.all_data_out[861] ),
    .A2(_04981_),
    .Y(_04985_),
    .B1(_04984_));
 sg13g2_o21ai_1 _12015_ (.B1(net4584),
    .Y(_04986_),
    .A1(\spiking_network_top_uut.all_data_out[862] ),
    .A2(_04980_));
 sg13g2_nand2_1 _12016_ (.Y(_04987_),
    .A(net3945),
    .B(net131));
 sg13g2_o21ai_1 _12017_ (.B1(_04987_),
    .Y(_00432_),
    .A1(_04985_),
    .A2(_04986_));
 sg13g2_mux2_1 _12018_ (.A0(net313),
    .A1(net131),
    .S(net4585),
    .X(_00433_));
 sg13g2_mux2_1 _12019_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[2] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[3] ),
    .S(\spiking_network_top_uut.all_data_out[856] ),
    .X(_04988_));
 sg13g2_nor2b_1 _12020_ (.A(\spiking_network_top_uut.all_data_out[856] ),
    .B_N(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[0] ),
    .Y(_04989_));
 sg13g2_a21oi_1 _12021_ (.A1(\spiking_network_top_uut.all_data_out[856] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[1] ),
    .Y(_04990_),
    .B1(_04989_));
 sg13g2_a21oi_1 _12022_ (.A1(\spiking_network_top_uut.all_data_out[857] ),
    .A2(_04988_),
    .Y(_04991_),
    .B1(\spiking_network_top_uut.all_data_out[858] ));
 sg13g2_o21ai_1 _12023_ (.B1(_04991_),
    .Y(_04992_),
    .A1(\spiking_network_top_uut.all_data_out[857] ),
    .A2(_04990_));
 sg13g2_mux2_1 _12024_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[6] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[7] ),
    .S(\spiking_network_top_uut.all_data_out[856] ),
    .X(_04993_));
 sg13g2_nor2b_1 _12025_ (.A(\spiking_network_top_uut.all_data_out[856] ),
    .B_N(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[4] ),
    .Y(_04994_));
 sg13g2_a21oi_1 _12026_ (.A1(\spiking_network_top_uut.all_data_out[856] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[5] ),
    .Y(_04995_),
    .B1(_04994_));
 sg13g2_o21ai_1 _12027_ (.B1(\spiking_network_top_uut.all_data_out[858] ),
    .Y(_04996_),
    .A1(\spiking_network_top_uut.all_data_out[857] ),
    .A2(_04995_));
 sg13g2_a21oi_2 _12028_ (.B1(_04996_),
    .Y(_04997_),
    .A2(_04993_),
    .A1(\spiking_network_top_uut.all_data_out[857] ));
 sg13g2_nand2_1 _12029_ (.Y(_04998_),
    .A(net4588),
    .B(_04992_));
 sg13g2_nand2_1 _12030_ (.Y(_04999_),
    .A(net3945),
    .B(net186));
 sg13g2_o21ai_1 _12031_ (.B1(_04999_),
    .Y(_00434_),
    .A1(_04997_),
    .A2(_04998_));
 sg13g2_mux2_1 _12032_ (.A0(net230),
    .A1(net186),
    .S(net4589),
    .X(_00435_));
 sg13g2_a21oi_1 _12033_ (.A1(\spiking_network_top_uut.all_data_out[852] ),
    .A2(_03668_),
    .Y(_05000_),
    .B1(\spiking_network_top_uut.all_data_out[853] ));
 sg13g2_o21ai_1 _12034_ (.B1(_05000_),
    .Y(_05001_),
    .A1(\spiking_network_top_uut.all_data_out[852] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[4] ));
 sg13g2_mux2_1 _12035_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[6] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[7] ),
    .S(\spiking_network_top_uut.all_data_out[852] ),
    .X(_05002_));
 sg13g2_nand2_1 _12036_ (.Y(_05003_),
    .A(\spiking_network_top_uut.all_data_out[853] ),
    .B(_05002_));
 sg13g2_nand3_1 _12037_ (.B(_05001_),
    .C(_05003_),
    .A(\spiking_network_top_uut.all_data_out[854] ),
    .Y(_05004_));
 sg13g2_mux2_1 _12038_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[2] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[3] ),
    .S(\spiking_network_top_uut.all_data_out[852] ),
    .X(_05005_));
 sg13g2_nor2b_1 _12039_ (.A(\spiking_network_top_uut.all_data_out[852] ),
    .B_N(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[0] ),
    .Y(_05006_));
 sg13g2_a21oi_1 _12040_ (.A1(\spiking_network_top_uut.all_data_out[852] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[1] ),
    .Y(_05007_),
    .B1(_05006_));
 sg13g2_a21oi_1 _12041_ (.A1(\spiking_network_top_uut.all_data_out[853] ),
    .A2(_05005_),
    .Y(_05008_),
    .B1(\spiking_network_top_uut.all_data_out[854] ));
 sg13g2_o21ai_1 _12042_ (.B1(_05008_),
    .Y(_05009_),
    .A1(\spiking_network_top_uut.all_data_out[853] ),
    .A2(_05007_));
 sg13g2_nand3_1 _12043_ (.B(_05004_),
    .C(_05009_),
    .A(net4582),
    .Y(_05010_));
 sg13g2_o21ai_1 _12044_ (.B1(_05010_),
    .Y(_00436_),
    .A1(net4581),
    .A2(_03669_));
 sg13g2_nor2_1 _12045_ (.A(net4581),
    .B(net84),
    .Y(_05011_));
 sg13g2_a21oi_1 _12046_ (.A1(net4581),
    .A2(_03669_),
    .Y(_00437_),
    .B1(_05011_));
 sg13g2_mux2_1 _12047_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[2] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[3] ),
    .S(\spiking_network_top_uut.all_data_out[848] ),
    .X(_05012_));
 sg13g2_nor2b_1 _12048_ (.A(\spiking_network_top_uut.all_data_out[848] ),
    .B_N(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[0] ),
    .Y(_05013_));
 sg13g2_a21oi_1 _12049_ (.A1(\spiking_network_top_uut.all_data_out[848] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[1] ),
    .Y(_05014_),
    .B1(_05013_));
 sg13g2_a21oi_1 _12050_ (.A1(\spiking_network_top_uut.all_data_out[849] ),
    .A2(_05012_),
    .Y(_05015_),
    .B1(\spiking_network_top_uut.all_data_out[850] ));
 sg13g2_o21ai_1 _12051_ (.B1(_05015_),
    .Y(_05016_),
    .A1(\spiking_network_top_uut.all_data_out[849] ),
    .A2(_05014_));
 sg13g2_mux2_1 _12052_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[6] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[7] ),
    .S(\spiking_network_top_uut.all_data_out[848] ),
    .X(_05017_));
 sg13g2_nor2b_1 _12053_ (.A(\spiking_network_top_uut.all_data_out[848] ),
    .B_N(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[4] ),
    .Y(_05018_));
 sg13g2_a21oi_1 _12054_ (.A1(\spiking_network_top_uut.all_data_out[848] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[5] ),
    .Y(_05019_),
    .B1(_05018_));
 sg13g2_o21ai_1 _12055_ (.B1(\spiking_network_top_uut.all_data_out[850] ),
    .Y(_05020_),
    .A1(\spiking_network_top_uut.all_data_out[849] ),
    .A2(_05019_));
 sg13g2_a21oi_1 _12056_ (.A1(\spiking_network_top_uut.all_data_out[849] ),
    .A2(_05017_),
    .Y(_05021_),
    .B1(_05020_));
 sg13g2_nand2_1 _12057_ (.Y(_05022_),
    .A(net4586),
    .B(_05016_));
 sg13g2_nand2_1 _12058_ (.Y(_05023_),
    .A(net3945),
    .B(net91));
 sg13g2_o21ai_1 _12059_ (.B1(_05023_),
    .Y(_00438_),
    .A1(_05021_),
    .A2(_05022_));
 sg13g2_mux2_1 _12060_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_dout ),
    .A1(net91),
    .S(net4586),
    .X(_00439_));
 sg13g2_mux4_1 _12061_ (.S0(\spiking_network_top_uut.all_data_out[844] ),
    .A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[0] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[1] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[2] ),
    .A3(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[3] ),
    .S1(\spiking_network_top_uut.all_data_out[845] ),
    .X(_05024_));
 sg13g2_mux2_1 _12062_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[6] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[7] ),
    .S(\spiking_network_top_uut.all_data_out[844] ),
    .X(_05025_));
 sg13g2_nor2b_1 _12063_ (.A(\spiking_network_top_uut.all_data_out[844] ),
    .B_N(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[4] ),
    .Y(_05026_));
 sg13g2_a21oi_1 _12064_ (.A1(\spiking_network_top_uut.all_data_out[844] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[5] ),
    .Y(_05027_),
    .B1(_05026_));
 sg13g2_o21ai_1 _12065_ (.B1(\spiking_network_top_uut.all_data_out[846] ),
    .Y(_05028_),
    .A1(\spiking_network_top_uut.all_data_out[845] ),
    .A2(_05027_));
 sg13g2_a21oi_1 _12066_ (.A1(\spiking_network_top_uut.all_data_out[845] ),
    .A2(_05025_),
    .Y(_05029_),
    .B1(_05028_));
 sg13g2_o21ai_1 _12067_ (.B1(net4573),
    .Y(_05030_),
    .A1(\spiking_network_top_uut.all_data_out[846] ),
    .A2(_05024_));
 sg13g2_nand2_1 _12068_ (.Y(_05031_),
    .A(net3946),
    .B(net70));
 sg13g2_o21ai_1 _12069_ (.B1(_05031_),
    .Y(_00440_),
    .A1(_05029_),
    .A2(_05030_));
 sg13g2_mux2_1 _12070_ (.A0(net222),
    .A1(net70),
    .S(net4577),
    .X(_00441_));
 sg13g2_nand2b_1 _12071_ (.Y(_05032_),
    .B(\spiking_network_top_uut.all_data_out[840] ),
    .A_N(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[5] ));
 sg13g2_nor2_1 _12072_ (.A(\spiking_network_top_uut.all_data_out[840] ),
    .B(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[4] ),
    .Y(_05033_));
 sg13g2_nor2_1 _12073_ (.A(\spiking_network_top_uut.all_data_out[841] ),
    .B(_05033_),
    .Y(_05034_));
 sg13g2_mux2_1 _12074_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[6] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[7] ),
    .S(\spiking_network_top_uut.all_data_out[840] ),
    .X(_05035_));
 sg13g2_a221oi_1 _12075_ (.B2(\spiking_network_top_uut.all_data_out[841] ),
    .C1(_03581_),
    .B1(_05035_),
    .A1(_05032_),
    .Y(_05036_),
    .A2(_05034_));
 sg13g2_mux4_1 _12076_ (.S0(\spiking_network_top_uut.all_data_out[840] ),
    .A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[0] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[1] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[2] ),
    .A3(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[3] ),
    .S1(\spiking_network_top_uut.all_data_out[841] ),
    .X(_05037_));
 sg13g2_o21ai_1 _12077_ (.B1(net4579),
    .Y(_05038_),
    .A1(\spiking_network_top_uut.all_data_out[842] ),
    .A2(_05037_));
 sg13g2_nand2_1 _12078_ (.Y(_05039_),
    .A(net3944),
    .B(net178));
 sg13g2_o21ai_1 _12079_ (.B1(_05039_),
    .Y(_00442_),
    .A1(_05036_),
    .A2(_05038_));
 sg13g2_mux2_1 _12080_ (.A0(net356),
    .A1(net178),
    .S(net4578),
    .X(_00443_));
 sg13g2_mux2_1 _12081_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[2] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[3] ),
    .S(\spiking_network_top_uut.all_data_out[836] ),
    .X(_05040_));
 sg13g2_nor2b_1 _12082_ (.A(\spiking_network_top_uut.all_data_out[836] ),
    .B_N(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[0] ),
    .Y(_05041_));
 sg13g2_a21oi_1 _12083_ (.A1(\spiking_network_top_uut.all_data_out[836] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[1] ),
    .Y(_05042_),
    .B1(_05041_));
 sg13g2_a21oi_1 _12084_ (.A1(\spiking_network_top_uut.all_data_out[837] ),
    .A2(_05040_),
    .Y(_05043_),
    .B1(\spiking_network_top_uut.all_data_out[838] ));
 sg13g2_o21ai_1 _12085_ (.B1(_05043_),
    .Y(_05044_),
    .A1(\spiking_network_top_uut.all_data_out[837] ),
    .A2(_05042_));
 sg13g2_mux2_1 _12086_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[6] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[7] ),
    .S(\spiking_network_top_uut.all_data_out[836] ),
    .X(_05045_));
 sg13g2_nor2b_1 _12087_ (.A(\spiking_network_top_uut.all_data_out[836] ),
    .B_N(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[4] ),
    .Y(_05046_));
 sg13g2_a21oi_1 _12088_ (.A1(\spiking_network_top_uut.all_data_out[836] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[5] ),
    .Y(_05047_),
    .B1(_05046_));
 sg13g2_o21ai_1 _12089_ (.B1(\spiking_network_top_uut.all_data_out[838] ),
    .Y(_05048_),
    .A1(\spiking_network_top_uut.all_data_out[837] ),
    .A2(_05047_));
 sg13g2_a21oi_1 _12090_ (.A1(\spiking_network_top_uut.all_data_out[837] ),
    .A2(_05045_),
    .Y(_05049_),
    .B1(_05048_));
 sg13g2_nand2_1 _12091_ (.Y(_05050_),
    .A(net4576),
    .B(_05044_));
 sg13g2_nand2_1 _12092_ (.Y(_05051_),
    .A(net3944),
    .B(net104));
 sg13g2_o21ai_1 _12093_ (.B1(_05051_),
    .Y(_00444_),
    .A1(_05049_),
    .A2(_05050_));
 sg13g2_mux2_1 _12094_ (.A0(net248),
    .A1(net104),
    .S(net4575),
    .X(_00445_));
 sg13g2_mux4_1 _12095_ (.S0(\spiking_network_top_uut.all_data_out[832] ),
    .A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[0] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[1] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[2] ),
    .A3(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[3] ),
    .S1(\spiking_network_top_uut.all_data_out[833] ),
    .X(_05052_));
 sg13g2_mux2_1 _12096_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[6] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[7] ),
    .S(\spiking_network_top_uut.all_data_out[832] ),
    .X(_05053_));
 sg13g2_nor2b_1 _12097_ (.A(\spiking_network_top_uut.all_data_out[832] ),
    .B_N(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[4] ),
    .Y(_05054_));
 sg13g2_a21oi_1 _12098_ (.A1(\spiking_network_top_uut.all_data_out[832] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[5] ),
    .Y(_05055_),
    .B1(_05054_));
 sg13g2_o21ai_1 _12099_ (.B1(\spiking_network_top_uut.all_data_out[834] ),
    .Y(_05056_),
    .A1(\spiking_network_top_uut.all_data_out[833] ),
    .A2(_05055_));
 sg13g2_a21oi_1 _12100_ (.A1(\spiking_network_top_uut.all_data_out[833] ),
    .A2(_05053_),
    .Y(_05057_),
    .B1(_05056_));
 sg13g2_o21ai_1 _12101_ (.B1(net4580),
    .Y(_05058_),
    .A1(\spiking_network_top_uut.all_data_out[834] ),
    .A2(_05052_));
 sg13g2_nand2_1 _12102_ (.Y(_05059_),
    .A(net3944),
    .B(net405));
 sg13g2_o21ai_1 _12103_ (.B1(_05059_),
    .Y(_00446_),
    .A1(_05057_),
    .A2(_05058_));
 sg13g2_nor3_2 _12104_ (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[2] ),
    .B(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[0] ),
    .C(net554),
    .Y(_05060_));
 sg13g2_nor2b_2 _12105_ (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[3] ),
    .B_N(_05060_),
    .Y(_05061_));
 sg13g2_nor2b_2 _12106_ (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[4] ),
    .B_N(_05061_),
    .Y(_05062_));
 sg13g2_nand2b_2 _12107_ (.Y(_05063_),
    .B(_05061_),
    .A_N(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[4] ));
 sg13g2_o21ai_1 _12108_ (.B1(net4574),
    .Y(_05064_),
    .A1(net3633),
    .A2(_05063_));
 sg13g2_nor2b_1 _12109_ (.A(net3632),
    .B_N(_00036_),
    .Y(_05065_));
 sg13g2_a21oi_1 _12110_ (.A1(net4283),
    .A2(net3632),
    .Y(_05066_),
    .B1(_05065_));
 sg13g2_nand2_1 _12111_ (.Y(_05067_),
    .A(net377),
    .B(_05064_));
 sg13g2_o21ai_1 _12112_ (.B1(_05067_),
    .Y(_00447_),
    .A1(_05064_),
    .A2(_05066_));
 sg13g2_xor2_1 _12113_ (.B(net351),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[0] ),
    .X(_05068_));
 sg13g2_nor2_1 _12114_ (.A(net3632),
    .B(_05068_),
    .Y(_05069_));
 sg13g2_a21oi_1 _12115_ (.A1(net4280),
    .A2(net3632),
    .Y(_05070_),
    .B1(_05069_));
 sg13g2_nand2_1 _12116_ (.Y(_05071_),
    .A(net351),
    .B(_05064_));
 sg13g2_o21ai_1 _12117_ (.B1(_05071_),
    .Y(_00448_),
    .A1(_05064_),
    .A2(_05070_));
 sg13g2_o21ai_1 _12118_ (.B1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[2] ),
    .Y(_05072_),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[0] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[1] ));
 sg13g2_nor2b_1 _12119_ (.A(_05060_),
    .B_N(_05072_),
    .Y(_05073_));
 sg13g2_nor2_1 _12120_ (.A(net3632),
    .B(_05073_),
    .Y(_05074_));
 sg13g2_a21oi_1 _12121_ (.A1(net4276),
    .A2(net3632),
    .Y(_05075_),
    .B1(_05074_));
 sg13g2_nand2_1 _12122_ (.Y(_05076_),
    .A(net212),
    .B(_05064_));
 sg13g2_o21ai_1 _12123_ (.B1(_05076_),
    .Y(_00449_),
    .A1(_05064_),
    .A2(_05075_));
 sg13g2_nand2_1 _12124_ (.Y(_05077_),
    .A(net4273),
    .B(net3632));
 sg13g2_xnor2_1 _12125_ (.Y(_05078_),
    .A(net434),
    .B(_05060_));
 sg13g2_o21ai_1 _12126_ (.B1(_05077_),
    .Y(_05079_),
    .A1(net3632),
    .A2(_05078_));
 sg13g2_mux2_1 _12127_ (.A0(_05079_),
    .A1(net434),
    .S(_05064_),
    .X(_00450_));
 sg13g2_nand2_1 _12128_ (.Y(_05080_),
    .A(net3942),
    .B(net275));
 sg13g2_nand2b_1 _12129_ (.Y(_05081_),
    .B(net275),
    .A_N(_05061_));
 sg13g2_a21oi_1 _12130_ (.A1(_05063_),
    .A2(_05081_),
    .Y(_05082_),
    .B1(net3633));
 sg13g2_a21oi_1 _12131_ (.A1(net4269),
    .A2(net3633),
    .Y(_05083_),
    .B1(_05082_));
 sg13g2_o21ai_1 _12132_ (.B1(_05080_),
    .Y(_00451_),
    .A1(_05064_),
    .A2(_05083_));
 sg13g2_mux2_1 _12133_ (.A0(net425),
    .A1(net405),
    .S(net4576),
    .X(_00452_));
 sg13g2_mux2_1 _12134_ (.A0(net3900),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[6] ),
    .S(net4551),
    .X(_00453_));
 sg13g2_nand2_2 _12135_ (.Y(_05084_),
    .A(net4268),
    .B(_00031_));
 sg13g2_nor2_1 _12136_ (.A(net4266),
    .B(_05084_),
    .Y(_05085_));
 sg13g2_nand3b_1 _12137_ (.B(net4268),
    .C(_00031_),
    .Y(_05086_),
    .A_N(net4267));
 sg13g2_nand2_1 _12138_ (.Y(_05087_),
    .A(net4266),
    .B(_00031_));
 sg13g2_or3_1 _12139_ (.A(net4266),
    .B(net4268),
    .C(_00031_),
    .X(_05088_));
 sg13g2_and2_1 _12140_ (.A(net3913),
    .B(net3909),
    .X(_05089_));
 sg13g2_nand2_2 _12141_ (.Y(_05090_),
    .A(net3913),
    .B(net3909));
 sg13g2_a21oi_1 _12142_ (.A1(net3913),
    .A2(net3909),
    .Y(_05091_),
    .B1(_00030_));
 sg13g2_nor2_2 _12143_ (.A(net3743),
    .B(_05091_),
    .Y(_05092_));
 sg13g2_nor2_1 _12144_ (.A(_00030_),
    .B(_05092_),
    .Y(_05093_));
 sg13g2_nand2b_1 _12145_ (.Y(_05094_),
    .B(_05092_),
    .A_N(_00030_));
 sg13g2_nor2_1 _12146_ (.A(_03429_),
    .B(_05093_),
    .Y(_05095_));
 sg13g2_a21o_1 _12147_ (.A2(net3743),
    .A1(_00032_),
    .B1(_05092_),
    .X(_05096_));
 sg13g2_nor2_1 _12148_ (.A(net4268),
    .B(net3915),
    .Y(_05097_));
 sg13g2_nand3b_1 _12149_ (.B(_00031_),
    .C(net4266),
    .Y(_05098_),
    .A_N(net4268));
 sg13g2_o21ai_1 _12150_ (.B1(net3916),
    .Y(_05099_),
    .A1(_00032_),
    .A2(net3903));
 sg13g2_a21oi_1 _12151_ (.A1(_05091_),
    .A2(net3903),
    .Y(_05100_),
    .B1(_05099_));
 sg13g2_a21oi_1 _12152_ (.A1(_00033_),
    .A2(net3743),
    .Y(_05101_),
    .B1(_05100_));
 sg13g2_or2_1 _12153_ (.X(_05102_),
    .B(_05101_),
    .A(_03431_));
 sg13g2_o21ai_1 _12154_ (.B1(net3913),
    .Y(_05103_),
    .A1(_00030_),
    .A2(net3909));
 sg13g2_and3_2 _12155_ (.X(_05104_),
    .A(net4267),
    .B(net4268),
    .C(_00031_));
 sg13g2_nand3_1 _12156_ (.B(net4268),
    .C(_00031_),
    .A(net4266),
    .Y(_05105_));
 sg13g2_a221oi_1 _12157_ (.B2(_00032_),
    .C1(net3743),
    .B1(net3901),
    .A1(_00033_),
    .Y(_05106_),
    .A2(net3738));
 sg13g2_a22oi_1 _12158_ (.Y(_05107_),
    .B1(_05103_),
    .B2(_05106_),
    .A2(net3743),
    .A1(_03474_));
 sg13g2_nor2b_1 _12159_ (.A(_05107_),
    .B_N(_00034_),
    .Y(_05108_));
 sg13g2_xnor2_1 _12160_ (.Y(_05109_),
    .A(_03431_),
    .B(_05101_));
 sg13g2_o21ai_1 _12161_ (.B1(_05102_),
    .Y(_05110_),
    .A1(_05108_),
    .A2(_05109_));
 sg13g2_xor2_1 _12162_ (.B(_05096_),
    .A(_00033_),
    .X(_05111_));
 sg13g2_nor2b_1 _12163_ (.A(_05111_),
    .B_N(_05110_),
    .Y(_05112_));
 sg13g2_a21o_1 _12164_ (.A2(_05096_),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ),
    .B1(_05112_),
    .X(_05113_));
 sg13g2_xnor2_1 _12165_ (.Y(_05114_),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ),
    .B(_05093_));
 sg13g2_a21oi_1 _12166_ (.A1(_05113_),
    .A2(_05114_),
    .Y(_05115_),
    .B1(_05095_));
 sg13g2_a22oi_1 _12167_ (.Y(_05116_),
    .B1(_05094_),
    .B2(_05115_),
    .A2(_05092_),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ));
 sg13g2_a21oi_2 _12168_ (.B1(_05116_),
    .Y(_05117_),
    .A2(_00030_),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ));
 sg13g2_nor2_1 _12169_ (.A(_05062_),
    .B(_05117_),
    .Y(_05118_));
 sg13g2_mux2_1 _12170_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.spike_out ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[839] ),
    .X(_05119_));
 sg13g2_nand2_1 _12171_ (.Y(_05120_),
    .A(\spiking_network_top_uut.all_data_out[291] ),
    .B(_05119_));
 sg13g2_mux2_1 _12172_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.spike_out ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[835] ),
    .X(_05121_));
 sg13g2_nand2_1 _12173_ (.Y(_05122_),
    .A(\spiking_network_top_uut.all_data_out[289] ),
    .B(_05121_));
 sg13g2_nor2_1 _12174_ (.A(_05120_),
    .B(_05122_),
    .Y(_05123_));
 sg13g2_nand4_1 _12175_ (.B(\spiking_network_top_uut.all_data_out[288] ),
    .C(_05119_),
    .A(\spiking_network_top_uut.all_data_out[290] ),
    .Y(_05124_),
    .D(_05121_));
 sg13g2_inv_1 _12176_ (.Y(_05125_),
    .A(_05124_));
 sg13g2_xor2_1 _12177_ (.B(_05122_),
    .A(_05120_),
    .X(_05126_));
 sg13g2_a21oi_2 _12178_ (.B1(_05123_),
    .Y(_05127_),
    .A2(_05126_),
    .A1(_05124_));
 sg13g2_mux2_1 _12179_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.spike_out ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[847] ),
    .X(_05128_));
 sg13g2_nand2_1 _12180_ (.Y(_05129_),
    .A(\spiking_network_top_uut.all_data_out[295] ),
    .B(_05128_));
 sg13g2_mux2_1 _12181_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.spike_out ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[843] ),
    .X(_05130_));
 sg13g2_nand2_1 _12182_ (.Y(_05131_),
    .A(\spiking_network_top_uut.all_data_out[293] ),
    .B(_05130_));
 sg13g2_nor2_1 _12183_ (.A(_05129_),
    .B(_05131_),
    .Y(_05132_));
 sg13g2_nand2_1 _12184_ (.Y(_05133_),
    .A(\spiking_network_top_uut.all_data_out[294] ),
    .B(_05128_));
 sg13g2_nand2_1 _12185_ (.Y(_05134_),
    .A(\spiking_network_top_uut.all_data_out[292] ),
    .B(_05130_));
 sg13g2_or2_2 _12186_ (.X(_05135_),
    .B(_05134_),
    .A(_05133_));
 sg13g2_xor2_1 _12187_ (.B(_05131_),
    .A(_05129_),
    .X(_05136_));
 sg13g2_a21oi_2 _12188_ (.B1(_05132_),
    .Y(_05137_),
    .A2(_05136_),
    .A1(_05135_));
 sg13g2_mux2_2 _12189_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.spike_out ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[855] ),
    .X(_05138_));
 sg13g2_mux2_2 _12190_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.spike_out ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[851] ),
    .X(_05139_));
 sg13g2_a22oi_1 _12191_ (.Y(_05140_),
    .B1(_05139_),
    .B2(\spiking_network_top_uut.all_data_out[297] ),
    .A2(_05138_),
    .A1(\spiking_network_top_uut.all_data_out[299] ));
 sg13g2_and4_1 _12192_ (.A(\spiking_network_top_uut.all_data_out[298] ),
    .B(\spiking_network_top_uut.all_data_out[296] ),
    .C(_05138_),
    .D(_05139_),
    .X(_05141_));
 sg13g2_nand4_1 _12193_ (.B(\spiking_network_top_uut.all_data_out[296] ),
    .C(_05138_),
    .A(\spiking_network_top_uut.all_data_out[298] ),
    .Y(_05142_),
    .D(_05139_));
 sg13g2_and4_1 _12194_ (.A(\spiking_network_top_uut.all_data_out[299] ),
    .B(\spiking_network_top_uut.all_data_out[297] ),
    .C(_05138_),
    .D(_05139_),
    .X(_05143_));
 sg13g2_nand4_1 _12195_ (.B(\spiking_network_top_uut.all_data_out[297] ),
    .C(_05138_),
    .A(\spiking_network_top_uut.all_data_out[299] ),
    .Y(_05144_),
    .D(_05139_));
 sg13g2_nand3b_1 _12196_ (.B(_05141_),
    .C(_05144_),
    .Y(_05145_),
    .A_N(_05140_));
 sg13g2_a21oi_2 _12197_ (.B1(_05140_),
    .Y(_05146_),
    .A2(_05144_),
    .A1(_05141_));
 sg13g2_mux2_2 _12198_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.spike_out ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[859] ),
    .X(_05147_));
 sg13g2_mux2_2 _12199_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.spike_out ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[863] ),
    .X(_05148_));
 sg13g2_and4_1 _12200_ (.A(\spiking_network_top_uut.all_data_out[301] ),
    .B(\spiking_network_top_uut.all_data_out[303] ),
    .C(_05147_),
    .D(_05148_),
    .X(_05149_));
 sg13g2_nand4_1 _12201_ (.B(\spiking_network_top_uut.all_data_out[303] ),
    .C(_05147_),
    .A(\spiking_network_top_uut.all_data_out[301] ),
    .Y(_05150_),
    .D(_05148_));
 sg13g2_and4_1 _12202_ (.A(\spiking_network_top_uut.all_data_out[300] ),
    .B(\spiking_network_top_uut.all_data_out[302] ),
    .C(_05147_),
    .D(_05148_),
    .X(_05151_));
 sg13g2_a22oi_1 _12203_ (.Y(_05152_),
    .B1(_05148_),
    .B2(\spiking_network_top_uut.all_data_out[303] ),
    .A2(_05147_),
    .A1(\spiking_network_top_uut.all_data_out[301] ));
 sg13g2_or3_2 _12204_ (.A(_05149_),
    .B(_05151_),
    .C(_05152_),
    .X(_05153_));
 sg13g2_o21ai_1 _12205_ (.B1(_05150_),
    .Y(_05154_),
    .A1(_05151_),
    .A2(_05152_));
 sg13g2_nand3b_1 _12206_ (.B(_05146_),
    .C(_05154_),
    .Y(_05155_),
    .A_N(_05137_));
 sg13g2_inv_1 _12207_ (.Y(_05156_),
    .A(_05155_));
 sg13g2_or2_1 _12208_ (.X(_05157_),
    .B(_05155_),
    .A(_05127_));
 sg13g2_nor2_1 _12209_ (.A(_05146_),
    .B(_05154_),
    .Y(_05158_));
 sg13g2_and2_1 _12210_ (.A(_05137_),
    .B(_05158_),
    .X(_05159_));
 sg13g2_nand2_1 _12211_ (.Y(_05160_),
    .A(_05127_),
    .B(_05159_));
 sg13g2_and2_1 _12212_ (.A(_05157_),
    .B(_05160_),
    .X(_05161_));
 sg13g2_xnor2_1 _12213_ (.Y(_05162_),
    .A(_05094_),
    .B(_05115_));
 sg13g2_nand2_1 _12214_ (.Y(_05163_),
    .A(_05161_),
    .B(_05162_));
 sg13g2_nand2_1 _12215_ (.Y(_05164_),
    .A(_05157_),
    .B(_05163_));
 sg13g2_xor2_1 _12216_ (.B(_05161_),
    .A(_05117_),
    .X(_05165_));
 sg13g2_nand2_1 _12217_ (.Y(_05166_),
    .A(_05164_),
    .B(_05165_));
 sg13g2_xnor2_1 _12218_ (.Y(_05167_),
    .A(_05161_),
    .B(_05162_));
 sg13g2_o21ai_1 _12219_ (.B1(_05151_),
    .Y(_05168_),
    .A1(_05149_),
    .A2(_05152_));
 sg13g2_o21ai_1 _12220_ (.B1(_05142_),
    .Y(_05169_),
    .A1(_05140_),
    .A2(_05143_));
 sg13g2_o21ai_1 _12221_ (.B1(_05141_),
    .Y(_05170_),
    .A1(_05140_),
    .A2(_05143_));
 sg13g2_nand3b_1 _12222_ (.B(_05142_),
    .C(_05144_),
    .Y(_05171_),
    .A_N(_05140_));
 sg13g2_a22oi_1 _12223_ (.Y(_05172_),
    .B1(_05170_),
    .B2(_05171_),
    .A2(_05168_),
    .A1(_05153_));
 sg13g2_xor2_1 _12224_ (.B(_05136_),
    .A(_05135_),
    .X(_05173_));
 sg13g2_xnor2_1 _12225_ (.Y(_05174_),
    .A(_05135_),
    .B(_05136_));
 sg13g2_and4_1 _12226_ (.A(_05153_),
    .B(_05168_),
    .C(_05170_),
    .D(_05171_),
    .X(_05175_));
 sg13g2_nand4_1 _12227_ (.B(_05168_),
    .C(_05170_),
    .A(_05153_),
    .Y(_05176_),
    .D(_05171_));
 sg13g2_and4_1 _12228_ (.A(_05145_),
    .B(_05153_),
    .C(_05168_),
    .D(_05169_),
    .X(_05177_));
 sg13g2_a22oi_1 _12229_ (.Y(_05178_),
    .B1(_05169_),
    .B2(_05145_),
    .A2(_05168_),
    .A1(_05153_));
 sg13g2_nor3_2 _12230_ (.A(_05172_),
    .B(_05173_),
    .C(_05175_),
    .Y(_05179_));
 sg13g2_a21oi_2 _12231_ (.B1(_05172_),
    .Y(_05180_),
    .A2(_05176_),
    .A1(_05174_));
 sg13g2_xor2_1 _12232_ (.B(_05154_),
    .A(_05146_),
    .X(_05181_));
 sg13g2_xnor2_1 _12233_ (.Y(_05182_),
    .A(_05137_),
    .B(_05181_));
 sg13g2_nand2b_1 _12234_ (.Y(_05183_),
    .B(_05182_),
    .A_N(_05180_));
 sg13g2_xnor2_1 _12235_ (.Y(_05184_),
    .A(_05180_),
    .B(_05182_));
 sg13g2_nand2b_1 _12236_ (.Y(_05185_),
    .B(_05184_),
    .A_N(_05127_));
 sg13g2_nand2_2 _12237_ (.Y(_05186_),
    .A(_05183_),
    .B(_05185_));
 sg13g2_nor2_1 _12238_ (.A(_05156_),
    .B(_05159_),
    .Y(_05187_));
 sg13g2_xnor2_1 _12239_ (.Y(_05188_),
    .A(_05127_),
    .B(_05187_));
 sg13g2_and2_1 _12240_ (.A(_05186_),
    .B(_05188_),
    .X(_05189_));
 sg13g2_xor2_1 _12241_ (.B(_05188_),
    .A(_05186_),
    .X(_05190_));
 sg13g2_xnor2_1 _12242_ (.Y(_05191_),
    .A(_05113_),
    .B(_05114_));
 sg13g2_inv_1 _12243_ (.Y(_05192_),
    .A(_05191_));
 sg13g2_a21oi_1 _12244_ (.A1(_05190_),
    .A2(_05192_),
    .Y(_05193_),
    .B1(_05189_));
 sg13g2_nor2_1 _12245_ (.A(_05167_),
    .B(_05193_),
    .Y(_05194_));
 sg13g2_xnor2_1 _12246_ (.Y(_05195_),
    .A(_05190_),
    .B(_05191_));
 sg13g2_a22oi_1 _12247_ (.Y(_05196_),
    .B1(_05148_),
    .B2(\spiking_network_top_uut.all_data_out[302] ),
    .A2(_05147_),
    .A1(\spiking_network_top_uut.all_data_out[300] ));
 sg13g2_nor2_2 _12248_ (.A(_05151_),
    .B(_05196_),
    .Y(_05197_));
 sg13g2_a22oi_1 _12249_ (.Y(_05198_),
    .B1(_05139_),
    .B2(\spiking_network_top_uut.all_data_out[296] ),
    .A2(_05138_),
    .A1(\spiking_network_top_uut.all_data_out[298] ));
 sg13g2_nor2_1 _12250_ (.A(_05141_),
    .B(_05198_),
    .Y(_05199_));
 sg13g2_and2_1 _12251_ (.A(_05197_),
    .B(_05199_),
    .X(_05200_));
 sg13g2_xor2_1 _12252_ (.B(_05134_),
    .A(_05133_),
    .X(_05201_));
 sg13g2_xor2_1 _12253_ (.B(_05199_),
    .A(_05197_),
    .X(_05202_));
 sg13g2_a21oi_2 _12254_ (.B1(_05200_),
    .Y(_05203_),
    .A2(_05202_),
    .A1(_05201_));
 sg13g2_nor3_2 _12255_ (.A(_05174_),
    .B(_05177_),
    .C(_05178_),
    .Y(_05204_));
 sg13g2_nor3_1 _12256_ (.A(_05179_),
    .B(_05203_),
    .C(_05204_),
    .Y(_05205_));
 sg13g2_or3_1 _12257_ (.A(_05179_),
    .B(_05203_),
    .C(_05204_),
    .X(_05206_));
 sg13g2_xnor2_1 _12258_ (.Y(_05207_),
    .A(_05124_),
    .B(_05126_));
 sg13g2_o21ai_1 _12259_ (.B1(_05203_),
    .Y(_05208_),
    .A1(_05179_),
    .A2(_05204_));
 sg13g2_nand3_1 _12260_ (.B(_05207_),
    .C(_05208_),
    .A(_05206_),
    .Y(_05209_));
 sg13g2_a21o_2 _12261_ (.A2(_05208_),
    .A1(_05207_),
    .B1(_05205_),
    .X(_05210_));
 sg13g2_xnor2_1 _12262_ (.Y(_05211_),
    .A(_05127_),
    .B(_05184_));
 sg13g2_nand2_1 _12263_ (.Y(_05212_),
    .A(_05210_),
    .B(_05211_));
 sg13g2_xnor2_1 _12264_ (.Y(_05213_),
    .A(_05210_),
    .B(_05211_));
 sg13g2_xor2_1 _12265_ (.B(_05111_),
    .A(_05110_),
    .X(_05214_));
 sg13g2_o21ai_1 _12266_ (.B1(_05212_),
    .Y(_05215_),
    .A1(_05213_),
    .A2(_05214_));
 sg13g2_nand2_1 _12267_ (.Y(_05216_),
    .A(_05195_),
    .B(_05215_));
 sg13g2_xor2_1 _12268_ (.B(_05214_),
    .A(_05213_),
    .X(_05217_));
 sg13g2_a22oi_1 _12269_ (.Y(_05218_),
    .B1(_05121_),
    .B2(\spiking_network_top_uut.all_data_out[288] ),
    .A2(_05119_),
    .A1(\spiking_network_top_uut.all_data_out[290] ));
 sg13g2_xnor2_1 _12270_ (.Y(_05219_),
    .A(_05201_),
    .B(_05202_));
 sg13g2_nor3_2 _12271_ (.A(_05125_),
    .B(_05218_),
    .C(_05219_),
    .Y(_05220_));
 sg13g2_a21o_2 _12272_ (.A2(_05208_),
    .A1(_05206_),
    .B1(_05207_),
    .X(_05221_));
 sg13g2_nand3_1 _12273_ (.B(_05220_),
    .C(_05221_),
    .A(_05209_),
    .Y(_05222_));
 sg13g2_a21oi_1 _12274_ (.A1(_05209_),
    .A2(_05221_),
    .Y(_05223_),
    .B1(_05220_));
 sg13g2_a21o_1 _12275_ (.A2(_05221_),
    .A1(_05209_),
    .B1(_05220_),
    .X(_05224_));
 sg13g2_xnor2_1 _12276_ (.Y(_05225_),
    .A(_05108_),
    .B(_05109_));
 sg13g2_inv_1 _12277_ (.Y(_05226_),
    .A(_05225_));
 sg13g2_and3_1 _12278_ (.X(_05227_),
    .A(_05222_),
    .B(_05224_),
    .C(_05226_));
 sg13g2_o21ai_1 _12279_ (.B1(_05222_),
    .Y(_05228_),
    .A1(_05223_),
    .A2(_05225_));
 sg13g2_and2_1 _12280_ (.A(_05217_),
    .B(_05228_),
    .X(_05229_));
 sg13g2_a21oi_1 _12281_ (.A1(_05222_),
    .A2(_05224_),
    .Y(_05230_),
    .B1(_05226_));
 sg13g2_nor2_1 _12282_ (.A(_05227_),
    .B(_05230_),
    .Y(_05231_));
 sg13g2_xnor2_1 _12283_ (.Y(_05232_),
    .A(_00034_),
    .B(_05107_));
 sg13g2_o21ai_1 _12284_ (.B1(_05219_),
    .Y(_05233_),
    .A1(_05125_),
    .A2(_05218_));
 sg13g2_nand2b_2 _12285_ (.Y(_05234_),
    .B(_05233_),
    .A_N(_05220_));
 sg13g2_nor2_1 _12286_ (.A(_05232_),
    .B(_05234_),
    .Y(_05235_));
 sg13g2_nor4_2 _12287_ (.A(_05227_),
    .B(_05230_),
    .C(_05232_),
    .Y(_05236_),
    .D(_05234_));
 sg13g2_xor2_1 _12288_ (.B(_05228_),
    .A(_05217_),
    .X(_05237_));
 sg13g2_a21oi_1 _12289_ (.A1(_05236_),
    .A2(_05237_),
    .Y(_05238_),
    .B1(_05229_));
 sg13g2_xnor2_1 _12290_ (.Y(_05239_),
    .A(_05195_),
    .B(_05215_));
 sg13g2_o21ai_1 _12291_ (.B1(_05216_),
    .Y(_05240_),
    .A1(_05238_),
    .A2(_05239_));
 sg13g2_nand2_1 _12292_ (.Y(_05241_),
    .A(_05167_),
    .B(_05193_));
 sg13g2_nand2b_1 _12293_ (.Y(_05242_),
    .B(_05241_),
    .A_N(_05194_));
 sg13g2_a21oi_1 _12294_ (.A1(_05240_),
    .A2(_05241_),
    .Y(_05243_),
    .B1(_05194_));
 sg13g2_xnor2_1 _12295_ (.Y(_05244_),
    .A(_05164_),
    .B(_05165_));
 sg13g2_o21ai_1 _12296_ (.B1(_05166_),
    .Y(_05245_),
    .A1(_05243_),
    .A2(_05244_));
 sg13g2_mux2_1 _12297_ (.A0(_05160_),
    .A1(_05157_),
    .S(_05117_),
    .X(_05246_));
 sg13g2_xnor2_1 _12298_ (.Y(_05247_),
    .A(_05245_),
    .B(_05246_));
 sg13g2_a21oi_2 _12299_ (.B1(_05118_),
    .Y(_05248_),
    .A2(_05247_),
    .A1(_05062_));
 sg13g2_xnor2_1 _12300_ (.Y(_05249_),
    .A(_05243_),
    .B(_05244_));
 sg13g2_a21oi_1 _12301_ (.A1(_05062_),
    .A2(_05249_),
    .Y(_05250_),
    .B1(_05118_));
 sg13g2_xnor2_1 _12302_ (.Y(_05251_),
    .A(_05240_),
    .B(_05242_));
 sg13g2_mux2_1 _12303_ (.A0(_05162_),
    .A1(_05251_),
    .S(_05062_),
    .X(_05252_));
 sg13g2_nand2_1 _12304_ (.Y(_05253_),
    .A(_05250_),
    .B(_05252_));
 sg13g2_a21oi_2 _12305_ (.B1(net3634),
    .Y(_05254_),
    .A2(_05253_),
    .A1(_05248_));
 sg13g2_nor2_1 _12306_ (.A(_05250_),
    .B(_05252_),
    .Y(_05255_));
 sg13g2_nor2_2 _12307_ (.A(_05248_),
    .B(_05255_),
    .Y(_05256_));
 sg13g2_nor2_1 _12308_ (.A(_05063_),
    .B(_05234_),
    .Y(_05257_));
 sg13g2_xnor2_1 _12309_ (.Y(_05258_),
    .A(_05232_),
    .B(_05257_));
 sg13g2_o21ai_1 _12310_ (.B1(_05254_),
    .Y(_05259_),
    .A1(_05256_),
    .A2(_05258_));
 sg13g2_xor2_1 _12311_ (.B(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[0] ),
    .A(net4311),
    .X(_05260_));
 sg13g2_a21oi_1 _12312_ (.A1(net3634),
    .A2(_05260_),
    .Y(_05261_),
    .B1(net3943));
 sg13g2_a22oi_1 _12313_ (.Y(_00454_),
    .B1(_05259_),
    .B2(_05261_),
    .A2(_03432_),
    .A1(net3943));
 sg13g2_nor2_1 _12314_ (.A(_05063_),
    .B(_05236_),
    .Y(_05262_));
 sg13g2_o21ai_1 _12315_ (.B1(_05262_),
    .Y(_05263_),
    .A1(_05231_),
    .A2(_05235_));
 sg13g2_o21ai_1 _12316_ (.B1(_05263_),
    .Y(_05264_),
    .A1(_05062_),
    .A2(_05225_));
 sg13g2_o21ai_1 _12317_ (.B1(_05254_),
    .Y(_05265_),
    .A1(_05256_),
    .A2(_05264_));
 sg13g2_xor2_1 _12318_ (.B(_04724_),
    .A(_04723_),
    .X(_05266_));
 sg13g2_a21oi_1 _12319_ (.A1(net3634),
    .A2(_05266_),
    .Y(_05267_),
    .B1(net3943));
 sg13g2_a22oi_1 _12320_ (.Y(_00455_),
    .B1(_05265_),
    .B2(_05267_),
    .A2(_03431_),
    .A1(net3943));
 sg13g2_and2_1 _12321_ (.A(_05063_),
    .B(_05214_),
    .X(_05268_));
 sg13g2_xnor2_1 _12322_ (.Y(_05269_),
    .A(_05236_),
    .B(_05237_));
 sg13g2_a21oi_1 _12323_ (.A1(_05062_),
    .A2(_05269_),
    .Y(_05270_),
    .B1(_05268_));
 sg13g2_o21ai_1 _12324_ (.B1(_05254_),
    .Y(_05271_),
    .A1(_05256_),
    .A2(_05270_));
 sg13g2_xnor2_1 _12325_ (.Y(_05272_),
    .A(_04721_),
    .B(_04725_));
 sg13g2_a21oi_1 _12326_ (.A1(net3634),
    .A2(_05272_),
    .Y(_05273_),
    .B1(net3941));
 sg13g2_a22oi_1 _12327_ (.Y(_00456_),
    .B1(_05271_),
    .B2(_05273_),
    .A2(_03430_),
    .A1(net3941));
 sg13g2_xor2_1 _12328_ (.B(_05239_),
    .A(_05238_),
    .X(_05274_));
 sg13g2_nand2_1 _12329_ (.Y(_05275_),
    .A(_05062_),
    .B(_05274_));
 sg13g2_o21ai_1 _12330_ (.B1(_05275_),
    .Y(_05276_),
    .A1(_05062_),
    .A2(_05191_));
 sg13g2_o21ai_1 _12331_ (.B1(_05254_),
    .Y(_05277_),
    .A1(_05256_),
    .A2(_05276_));
 sg13g2_or3_1 _12332_ (.A(_04719_),
    .B(_04720_),
    .C(_04726_),
    .X(_05278_));
 sg13g2_and2_1 _12333_ (.A(_04727_),
    .B(_05278_),
    .X(_05279_));
 sg13g2_a21oi_1 _12334_ (.A1(net3634),
    .A2(_05279_),
    .Y(_05280_),
    .B1(net3941));
 sg13g2_a22oi_1 _12335_ (.Y(_00457_),
    .B1(_05277_),
    .B2(_05280_),
    .A2(_03429_),
    .A1(net3941));
 sg13g2_nand2b_1 _12336_ (.Y(_05281_),
    .B(_05248_),
    .A_N(net3634));
 sg13g2_a21oi_1 _12337_ (.A1(_04718_),
    .A2(_04728_),
    .Y(_05282_),
    .B1(net3941));
 sg13g2_a22oi_1 _12338_ (.Y(_00458_),
    .B1(_05281_),
    .B2(_05282_),
    .A2(_03428_),
    .A1(net3941));
 sg13g2_mux2_1 _12339_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[2] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[3] ),
    .S(\spiking_network_top_uut.all_data_out[892] ),
    .X(_05283_));
 sg13g2_nor2b_1 _12340_ (.A(\spiking_network_top_uut.all_data_out[892] ),
    .B_N(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[0] ),
    .Y(_05284_));
 sg13g2_a21oi_1 _12341_ (.A1(\spiking_network_top_uut.all_data_out[892] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[1] ),
    .Y(_05285_),
    .B1(_05284_));
 sg13g2_a21oi_1 _12342_ (.A1(\spiking_network_top_uut.all_data_out[893] ),
    .A2(_05283_),
    .Y(_05286_),
    .B1(\spiking_network_top_uut.all_data_out[894] ));
 sg13g2_o21ai_1 _12343_ (.B1(_05286_),
    .Y(_05287_),
    .A1(\spiking_network_top_uut.all_data_out[893] ),
    .A2(_05285_));
 sg13g2_mux2_1 _12344_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[6] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[7] ),
    .S(\spiking_network_top_uut.all_data_out[892] ),
    .X(_05288_));
 sg13g2_nor2b_1 _12345_ (.A(\spiking_network_top_uut.all_data_out[892] ),
    .B_N(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[4] ),
    .Y(_05289_));
 sg13g2_a21oi_1 _12346_ (.A1(\spiking_network_top_uut.all_data_out[892] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[5] ),
    .Y(_05290_),
    .B1(_05289_));
 sg13g2_o21ai_1 _12347_ (.B1(\spiking_network_top_uut.all_data_out[894] ),
    .Y(_05291_),
    .A1(\spiking_network_top_uut.all_data_out[893] ),
    .A2(_05290_));
 sg13g2_a21oi_1 _12348_ (.A1(\spiking_network_top_uut.all_data_out[893] ),
    .A2(_05288_),
    .Y(_05292_),
    .B1(_05291_));
 sg13g2_nand2_1 _12349_ (.Y(_05293_),
    .A(net4585),
    .B(_05287_));
 sg13g2_nand2_1 _12350_ (.Y(_05294_),
    .A(net3945),
    .B(net60));
 sg13g2_o21ai_1 _12351_ (.B1(_05294_),
    .Y(_00459_),
    .A1(_05292_),
    .A2(_05293_));
 sg13g2_mux2_1 _12352_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[0] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.spike_out ),
    .S(net4589),
    .X(_00460_));
 sg13g2_mux2_1 _12353_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[1] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[0] ),
    .S(net4588),
    .X(_00461_));
 sg13g2_mux2_1 _12354_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[2] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[1] ),
    .S(net4589),
    .X(_00462_));
 sg13g2_mux2_1 _12355_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[3] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[2] ),
    .S(net4588),
    .X(_00463_));
 sg13g2_mux2_1 _12356_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[4] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[3] ),
    .S(net4588),
    .X(_00464_));
 sg13g2_mux2_1 _12357_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[5] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[4] ),
    .S(net4588),
    .X(_00465_));
 sg13g2_mux2_1 _12358_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[6] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[5] ),
    .S(net4588),
    .X(_00466_));
 sg13g2_mux2_1 _12359_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[7] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[6] ),
    .S(net4588),
    .X(_00467_));
 sg13g2_mux2_1 _12360_ (.A0(net237),
    .A1(net60),
    .S(net4585),
    .X(_00468_));
 sg13g2_mux2_1 _12361_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[2] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[3] ),
    .S(\spiking_network_top_uut.all_data_out[888] ),
    .X(_05295_));
 sg13g2_nor2b_1 _12362_ (.A(\spiking_network_top_uut.all_data_out[888] ),
    .B_N(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[0] ),
    .Y(_05296_));
 sg13g2_a21oi_1 _12363_ (.A1(\spiking_network_top_uut.all_data_out[888] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[1] ),
    .Y(_05297_),
    .B1(_05296_));
 sg13g2_a21oi_1 _12364_ (.A1(\spiking_network_top_uut.all_data_out[889] ),
    .A2(_05295_),
    .Y(_05298_),
    .B1(\spiking_network_top_uut.all_data_out[890] ));
 sg13g2_o21ai_1 _12365_ (.B1(_05298_),
    .Y(_05299_),
    .A1(\spiking_network_top_uut.all_data_out[889] ),
    .A2(_05297_));
 sg13g2_mux2_1 _12366_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[6] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[7] ),
    .S(\spiking_network_top_uut.all_data_out[888] ),
    .X(_05300_));
 sg13g2_nor2b_1 _12367_ (.A(\spiking_network_top_uut.all_data_out[888] ),
    .B_N(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[4] ),
    .Y(_05301_));
 sg13g2_a21oi_1 _12368_ (.A1(\spiking_network_top_uut.all_data_out[888] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[5] ),
    .Y(_05302_),
    .B1(_05301_));
 sg13g2_o21ai_1 _12369_ (.B1(\spiking_network_top_uut.all_data_out[890] ),
    .Y(_05303_),
    .A1(\spiking_network_top_uut.all_data_out[889] ),
    .A2(_05302_));
 sg13g2_a21oi_2 _12370_ (.B1(_05303_),
    .Y(_05304_),
    .A2(_05300_),
    .A1(\spiking_network_top_uut.all_data_out[889] ));
 sg13g2_nand2_1 _12371_ (.Y(_05305_),
    .A(net4588),
    .B(_05299_));
 sg13g2_nand2_1 _12372_ (.Y(_05306_),
    .A(net3944),
    .B(net204));
 sg13g2_o21ai_1 _12373_ (.B1(_05306_),
    .Y(_00469_),
    .A1(_05304_),
    .A2(_05305_));
 sg13g2_mux2_1 _12374_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[0] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.spike_out ),
    .S(net4582),
    .X(_00470_));
 sg13g2_mux2_1 _12375_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[1] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[0] ),
    .S(net4582),
    .X(_00471_));
 sg13g2_mux2_1 _12376_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[2] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[1] ),
    .S(net4582),
    .X(_00472_));
 sg13g2_mux2_1 _12377_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[3] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[2] ),
    .S(net4582),
    .X(_00473_));
 sg13g2_mux2_1 _12378_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[4] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[3] ),
    .S(net4582),
    .X(_00474_));
 sg13g2_nand2_1 _12379_ (.Y(_05307_),
    .A(net4581),
    .B(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[4] ));
 sg13g2_o21ai_1 _12380_ (.B1(_05307_),
    .Y(_00475_),
    .A1(net4581),
    .A2(_03668_));
 sg13g2_nor2_1 _12381_ (.A(net4581),
    .B(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[6] ),
    .Y(_05308_));
 sg13g2_a21oi_1 _12382_ (.A1(net4581),
    .A2(_03668_),
    .Y(_00476_),
    .B1(_05308_));
 sg13g2_mux2_1 _12383_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[7] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[6] ),
    .S(net4581),
    .X(_00477_));
 sg13g2_mux2_1 _12384_ (.A0(net299),
    .A1(net204),
    .S(net4589),
    .X(_00478_));
 sg13g2_mux4_1 _12385_ (.S0(\spiking_network_top_uut.all_data_out[884] ),
    .A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[0] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[1] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[2] ),
    .A3(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[3] ),
    .S1(\spiking_network_top_uut.all_data_out[885] ),
    .X(_05309_));
 sg13g2_mux2_1 _12386_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[6] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[7] ),
    .S(\spiking_network_top_uut.all_data_out[884] ),
    .X(_05310_));
 sg13g2_nor2b_1 _12387_ (.A(\spiking_network_top_uut.all_data_out[884] ),
    .B_N(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[4] ),
    .Y(_05311_));
 sg13g2_a21oi_1 _12388_ (.A1(\spiking_network_top_uut.all_data_out[884] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[5] ),
    .Y(_05312_),
    .B1(_05311_));
 sg13g2_o21ai_1 _12389_ (.B1(\spiking_network_top_uut.all_data_out[886] ),
    .Y(_05313_),
    .A1(\spiking_network_top_uut.all_data_out[885] ),
    .A2(_05312_));
 sg13g2_a21oi_1 _12390_ (.A1(\spiking_network_top_uut.all_data_out[885] ),
    .A2(_05310_),
    .Y(_05314_),
    .B1(_05313_));
 sg13g2_o21ai_1 _12391_ (.B1(net4583),
    .Y(_05315_),
    .A1(\spiking_network_top_uut.all_data_out[886] ),
    .A2(_05309_));
 sg13g2_nand2_1 _12392_ (.Y(_05316_),
    .A(net3945),
    .B(net137));
 sg13g2_o21ai_1 _12393_ (.B1(_05316_),
    .Y(_00479_),
    .A1(_05314_),
    .A2(_05315_));
 sg13g2_mux2_1 _12394_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[0] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.spike_out ),
    .S(net4586),
    .X(_00480_));
 sg13g2_mux2_1 _12395_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[1] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[0] ),
    .S(net4587),
    .X(_00481_));
 sg13g2_mux2_1 _12396_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[2] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[1] ),
    .S(net4587),
    .X(_00482_));
 sg13g2_mux2_1 _12397_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[3] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[2] ),
    .S(net4586),
    .X(_00483_));
 sg13g2_mux2_1 _12398_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[4] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[3] ),
    .S(net4586),
    .X(_00484_));
 sg13g2_mux2_1 _12399_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[5] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[4] ),
    .S(net4586),
    .X(_00485_));
 sg13g2_mux2_1 _12400_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[6] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[5] ),
    .S(net4590),
    .X(_00486_));
 sg13g2_mux2_1 _12401_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[7] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[6] ),
    .S(net4590),
    .X(_00487_));
 sg13g2_mux2_1 _12402_ (.A0(net289),
    .A1(net137),
    .S(net4582),
    .X(_00488_));
 sg13g2_nand2b_1 _12403_ (.Y(_05317_),
    .B(\spiking_network_top_uut.all_data_out[880] ),
    .A_N(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[5] ));
 sg13g2_nor2_1 _12404_ (.A(\spiking_network_top_uut.all_data_out[880] ),
    .B(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[4] ),
    .Y(_05318_));
 sg13g2_nor2_1 _12405_ (.A(\spiking_network_top_uut.all_data_out[881] ),
    .B(_05318_),
    .Y(_05319_));
 sg13g2_mux2_1 _12406_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[6] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[7] ),
    .S(\spiking_network_top_uut.all_data_out[880] ),
    .X(_05320_));
 sg13g2_a221oi_1 _12407_ (.B2(\spiking_network_top_uut.all_data_out[881] ),
    .C1(_03577_),
    .B1(_05320_),
    .A1(_05317_),
    .Y(_05321_),
    .A2(_05319_));
 sg13g2_mux4_1 _12408_ (.S0(\spiking_network_top_uut.all_data_out[880] ),
    .A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[0] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[1] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[2] ),
    .A3(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[3] ),
    .S1(\spiking_network_top_uut.all_data_out[881] ),
    .X(_05322_));
 sg13g2_o21ai_1 _12409_ (.B1(net4586),
    .Y(_05323_),
    .A1(\spiking_network_top_uut.all_data_out[882] ),
    .A2(_05322_));
 sg13g2_nand2_1 _12410_ (.Y(_05324_),
    .A(net3944),
    .B(net83));
 sg13g2_o21ai_1 _12411_ (.B1(_05324_),
    .Y(_00489_),
    .A1(_05321_),
    .A2(_05323_));
 sg13g2_mux2_1 _12412_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[0] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.spike_out ),
    .S(net4573),
    .X(_00490_));
 sg13g2_mux2_1 _12413_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[1] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[0] ),
    .S(net4573),
    .X(_00491_));
 sg13g2_mux2_1 _12414_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[2] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[1] ),
    .S(net4574),
    .X(_00492_));
 sg13g2_mux2_1 _12415_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[3] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[2] ),
    .S(net4573),
    .X(_00493_));
 sg13g2_mux2_1 _12416_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[4] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[3] ),
    .S(net4573),
    .X(_00494_));
 sg13g2_mux2_1 _12417_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[5] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[4] ),
    .S(net4573),
    .X(_00495_));
 sg13g2_mux2_1 _12418_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[6] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[5] ),
    .S(net4573),
    .X(_00496_));
 sg13g2_mux2_1 _12419_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[7] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[6] ),
    .S(net4577),
    .X(_00497_));
 sg13g2_mux2_1 _12420_ (.A0(net147),
    .A1(net83),
    .S(net4586),
    .X(_00498_));
 sg13g2_mux2_1 _12421_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[2] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[3] ),
    .S(\spiking_network_top_uut.all_data_out[876] ),
    .X(_05325_));
 sg13g2_nor2b_1 _12422_ (.A(\spiking_network_top_uut.all_data_out[876] ),
    .B_N(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[0] ),
    .Y(_05326_));
 sg13g2_a21oi_1 _12423_ (.A1(\spiking_network_top_uut.all_data_out[876] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[1] ),
    .Y(_05327_),
    .B1(_05326_));
 sg13g2_a21oi_1 _12424_ (.A1(\spiking_network_top_uut.all_data_out[877] ),
    .A2(_05325_),
    .Y(_05328_),
    .B1(\spiking_network_top_uut.all_data_out[878] ));
 sg13g2_o21ai_1 _12425_ (.B1(_05328_),
    .Y(_05329_),
    .A1(\spiking_network_top_uut.all_data_out[877] ),
    .A2(_05327_));
 sg13g2_mux2_1 _12426_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[6] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[7] ),
    .S(\spiking_network_top_uut.all_data_out[876] ),
    .X(_05330_));
 sg13g2_nor2b_1 _12427_ (.A(\spiking_network_top_uut.all_data_out[876] ),
    .B_N(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[4] ),
    .Y(_05331_));
 sg13g2_a21oi_1 _12428_ (.A1(\spiking_network_top_uut.all_data_out[876] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[5] ),
    .Y(_05332_),
    .B1(_05331_));
 sg13g2_o21ai_1 _12429_ (.B1(\spiking_network_top_uut.all_data_out[878] ),
    .Y(_05333_),
    .A1(\spiking_network_top_uut.all_data_out[877] ),
    .A2(_05332_));
 sg13g2_a21oi_1 _12430_ (.A1(\spiking_network_top_uut.all_data_out[877] ),
    .A2(_05330_),
    .Y(_05334_),
    .B1(_05333_));
 sg13g2_nand2_1 _12431_ (.Y(_05335_),
    .A(net4573),
    .B(_05329_));
 sg13g2_nand2_1 _12432_ (.Y(_05336_),
    .A(net3946),
    .B(net54));
 sg13g2_o21ai_1 _12433_ (.B1(_05336_),
    .Y(_00499_),
    .A1(_05334_),
    .A2(_05335_));
 sg13g2_mux2_1 _12434_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[0] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.spike_out ),
    .S(net4578),
    .X(_00500_));
 sg13g2_mux2_1 _12435_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[1] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[0] ),
    .S(net4578),
    .X(_00501_));
 sg13g2_mux2_1 _12436_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[2] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[1] ),
    .S(net4578),
    .X(_00502_));
 sg13g2_mux2_1 _12437_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[3] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[2] ),
    .S(net4578),
    .X(_00503_));
 sg13g2_mux2_1 _12438_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[4] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[3] ),
    .S(net4579),
    .X(_00504_));
 sg13g2_mux2_1 _12439_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[5] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[4] ),
    .S(net4579),
    .X(_00505_));
 sg13g2_mux2_1 _12440_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[6] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[5] ),
    .S(net4579),
    .X(_00506_));
 sg13g2_mux2_1 _12441_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[7] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[6] ),
    .S(net4579),
    .X(_00507_));
 sg13g2_mux2_1 _12442_ (.A0(net203),
    .A1(net54),
    .S(net4577),
    .X(_00508_));
 sg13g2_mux4_1 _12443_ (.S0(\spiking_network_top_uut.all_data_out[872] ),
    .A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[0] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[1] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[2] ),
    .A3(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[3] ),
    .S1(\spiking_network_top_uut.all_data_out[873] ),
    .X(_05337_));
 sg13g2_mux2_1 _12444_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[6] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[7] ),
    .S(\spiking_network_top_uut.all_data_out[872] ),
    .X(_05338_));
 sg13g2_nor2b_1 _12445_ (.A(\spiking_network_top_uut.all_data_out[872] ),
    .B_N(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[4] ),
    .Y(_05339_));
 sg13g2_a21oi_1 _12446_ (.A1(\spiking_network_top_uut.all_data_out[872] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[5] ),
    .Y(_05340_),
    .B1(_05339_));
 sg13g2_o21ai_1 _12447_ (.B1(\spiking_network_top_uut.all_data_out[874] ),
    .Y(_05341_),
    .A1(\spiking_network_top_uut.all_data_out[873] ),
    .A2(_05340_));
 sg13g2_a21oi_1 _12448_ (.A1(\spiking_network_top_uut.all_data_out[873] ),
    .A2(_05338_),
    .Y(_05342_),
    .B1(_05341_));
 sg13g2_o21ai_1 _12449_ (.B1(net4579),
    .Y(_05343_),
    .A1(\spiking_network_top_uut.all_data_out[874] ),
    .A2(_05337_));
 sg13g2_nand2_1 _12450_ (.Y(_05344_),
    .A(net3944),
    .B(net143));
 sg13g2_o21ai_1 _12451_ (.B1(_05344_),
    .Y(_00509_),
    .A1(_05342_),
    .A2(_05343_));
 sg13g2_mux2_1 _12452_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[0] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.spike_out ),
    .S(net4575),
    .X(_00510_));
 sg13g2_mux2_1 _12453_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[1] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[0] ),
    .S(net4575),
    .X(_00511_));
 sg13g2_mux2_1 _12454_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[2] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[1] ),
    .S(net4575),
    .X(_00512_));
 sg13g2_mux2_1 _12455_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[3] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[2] ),
    .S(net4575),
    .X(_00513_));
 sg13g2_mux2_1 _12456_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[4] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[3] ),
    .S(net4575),
    .X(_00514_));
 sg13g2_mux2_1 _12457_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[5] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[4] ),
    .S(net4575),
    .X(_00515_));
 sg13g2_mux2_1 _12458_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[6] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[5] ),
    .S(net4575),
    .X(_00516_));
 sg13g2_mux2_1 _12459_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[7] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[6] ),
    .S(net4578),
    .X(_00517_));
 sg13g2_mux2_1 _12460_ (.A0(net302),
    .A1(net143),
    .S(net4578),
    .X(_00518_));
 sg13g2_mux4_1 _12461_ (.S0(\spiking_network_top_uut.all_data_out[868] ),
    .A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[0] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[1] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[2] ),
    .A3(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[3] ),
    .S1(\spiking_network_top_uut.all_data_out[869] ),
    .X(_05345_));
 sg13g2_mux2_1 _12462_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[6] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[7] ),
    .S(\spiking_network_top_uut.all_data_out[868] ),
    .X(_05346_));
 sg13g2_nor2b_1 _12463_ (.A(\spiking_network_top_uut.all_data_out[868] ),
    .B_N(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[4] ),
    .Y(_05347_));
 sg13g2_a21oi_1 _12464_ (.A1(\spiking_network_top_uut.all_data_out[868] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[5] ),
    .Y(_05348_),
    .B1(_05347_));
 sg13g2_o21ai_1 _12465_ (.B1(\spiking_network_top_uut.all_data_out[870] ),
    .Y(_05349_),
    .A1(\spiking_network_top_uut.all_data_out[869] ),
    .A2(_05348_));
 sg13g2_a21oi_1 _12466_ (.A1(\spiking_network_top_uut.all_data_out[869] ),
    .A2(_05346_),
    .Y(_05350_),
    .B1(_05349_));
 sg13g2_o21ai_1 _12467_ (.B1(net4578),
    .Y(_05351_),
    .A1(\spiking_network_top_uut.all_data_out[870] ),
    .A2(_05345_));
 sg13g2_nand2_1 _12468_ (.Y(_05352_),
    .A(net3944),
    .B(net127));
 sg13g2_o21ai_1 _12469_ (.B1(_05352_),
    .Y(_00519_),
    .A1(_05350_),
    .A2(_05351_));
 sg13g2_mux2_1 _12470_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[0] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.spike_out ),
    .S(net4576),
    .X(_00520_));
 sg13g2_mux2_1 _12471_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[1] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[0] ),
    .S(net4580),
    .X(_00521_));
 sg13g2_mux2_1 _12472_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[2] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[1] ),
    .S(net4580),
    .X(_00522_));
 sg13g2_mux2_1 _12473_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[3] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[2] ),
    .S(net4580),
    .X(_00523_));
 sg13g2_mux2_1 _12474_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[4] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[3] ),
    .S(net4580),
    .X(_00524_));
 sg13g2_mux2_1 _12475_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[5] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[4] ),
    .S(net4580),
    .X(_00525_));
 sg13g2_mux2_1 _12476_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[6] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[5] ),
    .S(net4580),
    .X(_00526_));
 sg13g2_mux2_1 _12477_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[7] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[6] ),
    .S(net4583),
    .X(_00527_));
 sg13g2_mux2_1 _12478_ (.A0(net325),
    .A1(net127),
    .S(net4577),
    .X(_00528_));
 sg13g2_mux4_1 _12479_ (.S0(\spiking_network_top_uut.all_data_out[864] ),
    .A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[0] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[1] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[2] ),
    .A3(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[3] ),
    .S1(\spiking_network_top_uut.all_data_out[865] ),
    .X(_05353_));
 sg13g2_mux2_1 _12480_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[6] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[7] ),
    .S(\spiking_network_top_uut.all_data_out[864] ),
    .X(_05354_));
 sg13g2_nor2b_1 _12481_ (.A(\spiking_network_top_uut.all_data_out[864] ),
    .B_N(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[4] ),
    .Y(_05355_));
 sg13g2_a21oi_1 _12482_ (.A1(\spiking_network_top_uut.all_data_out[864] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[5] ),
    .Y(_05356_),
    .B1(_05355_));
 sg13g2_o21ai_1 _12483_ (.B1(\spiking_network_top_uut.all_data_out[866] ),
    .Y(_05357_),
    .A1(\spiking_network_top_uut.all_data_out[865] ),
    .A2(_05356_));
 sg13g2_a21oi_1 _12484_ (.A1(\spiking_network_top_uut.all_data_out[865] ),
    .A2(_05354_),
    .Y(_05358_),
    .B1(_05357_));
 sg13g2_o21ai_1 _12485_ (.B1(net4580),
    .Y(_05359_),
    .A1(\spiking_network_top_uut.all_data_out[866] ),
    .A2(_05353_));
 sg13g2_nand2_1 _12486_ (.Y(_05360_),
    .A(net3944),
    .B(net219));
 sg13g2_o21ai_1 _12487_ (.B1(_05360_),
    .Y(_00529_),
    .A1(_05358_),
    .A2(_05359_));
 sg13g2_nor3_2 _12488_ (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[2] ),
    .B(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[1] ),
    .C(net555),
    .Y(_05361_));
 sg13g2_nor2b_2 _12489_ (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[3] ),
    .B_N(_05361_),
    .Y(_05362_));
 sg13g2_nor2b_2 _12490_ (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[4] ),
    .B_N(_05362_),
    .Y(_05363_));
 sg13g2_nand2b_2 _12491_ (.Y(_05364_),
    .B(_05362_),
    .A_N(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[4] ));
 sg13g2_o21ai_1 _12492_ (.B1(net4574),
    .Y(_05365_),
    .A1(net3630),
    .A2(_05364_));
 sg13g2_nor2b_1 _12493_ (.A(net3629),
    .B_N(_00042_),
    .Y(_05366_));
 sg13g2_a21oi_1 _12494_ (.A1(net4283),
    .A2(net3629),
    .Y(_05367_),
    .B1(_05366_));
 sg13g2_nand2_1 _12495_ (.Y(_05368_),
    .A(net337),
    .B(_05365_));
 sg13g2_o21ai_1 _12496_ (.B1(_05368_),
    .Y(_00530_),
    .A1(_05365_),
    .A2(_05367_));
 sg13g2_xor2_1 _12497_ (.B(net337),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[1] ),
    .X(_05369_));
 sg13g2_nor2_1 _12498_ (.A(net3629),
    .B(_05369_),
    .Y(_05370_));
 sg13g2_a21oi_1 _12499_ (.A1(net4280),
    .A2(net3629),
    .Y(_05371_),
    .B1(_05370_));
 sg13g2_nand2_1 _12500_ (.Y(_05372_),
    .A(net409),
    .B(_05365_));
 sg13g2_o21ai_1 _12501_ (.B1(_05372_),
    .Y(_00531_),
    .A1(_05365_),
    .A2(_05371_));
 sg13g2_o21ai_1 _12502_ (.B1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[2] ),
    .Y(_05373_),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[1] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[0] ));
 sg13g2_nor2b_1 _12503_ (.A(net556),
    .B_N(_05373_),
    .Y(_05374_));
 sg13g2_nor2_1 _12504_ (.A(net3629),
    .B(_05374_),
    .Y(_05375_));
 sg13g2_a21oi_1 _12505_ (.A1(net4276),
    .A2(net3629),
    .Y(_05376_),
    .B1(_05375_));
 sg13g2_nand2_1 _12506_ (.Y(_05377_),
    .A(net156),
    .B(_05365_));
 sg13g2_o21ai_1 _12507_ (.B1(_05377_),
    .Y(_00532_),
    .A1(_05365_),
    .A2(_05376_));
 sg13g2_nand2_1 _12508_ (.Y(_05378_),
    .A(net4273),
    .B(net3629));
 sg13g2_xnor2_1 _12509_ (.Y(_05379_),
    .A(net427),
    .B(_05361_));
 sg13g2_o21ai_1 _12510_ (.B1(_05378_),
    .Y(_05380_),
    .A1(net3629),
    .A2(_05379_));
 sg13g2_mux2_1 _12511_ (.A0(_05380_),
    .A1(net427),
    .S(_05365_),
    .X(_00533_));
 sg13g2_nand2_1 _12512_ (.Y(_05381_),
    .A(net225),
    .B(net3942));
 sg13g2_nand2b_1 _12513_ (.Y(_05382_),
    .B(net225),
    .A_N(_05362_));
 sg13g2_a21oi_1 _12514_ (.A1(_05364_),
    .A2(_05382_),
    .Y(_05383_),
    .B1(net3630));
 sg13g2_a21oi_1 _12515_ (.A1(net4269),
    .A2(net3630),
    .Y(_05384_),
    .B1(_05383_));
 sg13g2_o21ai_1 _12516_ (.B1(_05381_),
    .Y(_00534_),
    .A1(_05365_),
    .A2(_05384_));
 sg13g2_mux2_1 _12517_ (.A0(net437),
    .A1(net219),
    .S(net4576),
    .X(_00535_));
 sg13g2_a21oi_1 _12518_ (.A1(net3913),
    .A2(net3909),
    .Y(_05385_),
    .B1(_00037_));
 sg13g2_nor2_2 _12519_ (.A(net3742),
    .B(_05385_),
    .Y(_05386_));
 sg13g2_nor2_1 _12520_ (.A(_00037_),
    .B(_05386_),
    .Y(_05387_));
 sg13g2_nand2b_1 _12521_ (.Y(_05388_),
    .B(_05386_),
    .A_N(_00037_));
 sg13g2_nor2_1 _12522_ (.A(_03409_),
    .B(_05387_),
    .Y(_05389_));
 sg13g2_a21o_1 _12523_ (.A2(net3742),
    .A1(_00038_),
    .B1(_05386_),
    .X(_05390_));
 sg13g2_o21ai_1 _12524_ (.B1(net3916),
    .Y(_05391_),
    .A1(_00038_),
    .A2(net3903));
 sg13g2_a21oi_1 _12525_ (.A1(net3903),
    .A2(_05385_),
    .Y(_05392_),
    .B1(_05391_));
 sg13g2_a21oi_1 _12526_ (.A1(_00039_),
    .A2(net3742),
    .Y(_05393_),
    .B1(_05392_));
 sg13g2_or2_1 _12527_ (.X(_05394_),
    .B(_05393_),
    .A(_03408_));
 sg13g2_o21ai_1 _12528_ (.B1(net3913),
    .Y(_05395_),
    .A1(_00037_),
    .A2(net3909));
 sg13g2_a221oi_1 _12529_ (.B2(_00038_),
    .C1(net3742),
    .B1(net3901),
    .A1(_00039_),
    .Y(_05396_),
    .A2(net3738));
 sg13g2_a22oi_1 _12530_ (.Y(_05397_),
    .B1(_05395_),
    .B2(_05396_),
    .A2(net3742),
    .A1(_03478_));
 sg13g2_nor2b_1 _12531_ (.A(_05397_),
    .B_N(_00040_),
    .Y(_05398_));
 sg13g2_xnor2_1 _12532_ (.Y(_05399_),
    .A(_03408_),
    .B(_05393_));
 sg13g2_o21ai_1 _12533_ (.B1(_05394_),
    .Y(_05400_),
    .A1(_05398_),
    .A2(_05399_));
 sg13g2_xor2_1 _12534_ (.B(_05390_),
    .A(_00039_),
    .X(_05401_));
 sg13g2_nor2b_1 _12535_ (.A(_05401_),
    .B_N(_05400_),
    .Y(_05402_));
 sg13g2_a21o_1 _12536_ (.A2(_05390_),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ),
    .B1(_05402_),
    .X(_05403_));
 sg13g2_xnor2_1 _12537_ (.Y(_05404_),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ),
    .B(_05387_));
 sg13g2_a21oi_2 _12538_ (.B1(_05389_),
    .Y(_05405_),
    .A2(_05404_),
    .A1(_05403_));
 sg13g2_a22oi_1 _12539_ (.Y(_05406_),
    .B1(_05388_),
    .B2(_05405_),
    .A2(_05386_),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ));
 sg13g2_a21oi_2 _12540_ (.B1(_05406_),
    .Y(_05407_),
    .A2(_00037_),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ));
 sg13g2_nor2_1 _12541_ (.A(_05363_),
    .B(_05407_),
    .Y(_05408_));
 sg13g2_mux2_1 _12542_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.spike_out ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[1].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[867] ),
    .X(_05409_));
 sg13g2_nand2_1 _12543_ (.Y(_05410_),
    .A(\spiking_network_top_uut.all_data_out[305] ),
    .B(_05409_));
 sg13g2_mux2_1 _12544_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.spike_out ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[1].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[871] ),
    .X(_05411_));
 sg13g2_nand2_1 _12545_ (.Y(_05412_),
    .A(\spiking_network_top_uut.all_data_out[307] ),
    .B(_05411_));
 sg13g2_nor2_1 _12546_ (.A(_05410_),
    .B(_05412_),
    .Y(_05413_));
 sg13g2_nand4_1 _12547_ (.B(\spiking_network_top_uut.all_data_out[306] ),
    .C(_05409_),
    .A(\spiking_network_top_uut.all_data_out[304] ),
    .Y(_05414_),
    .D(_05411_));
 sg13g2_inv_1 _12548_ (.Y(_05415_),
    .A(_05414_));
 sg13g2_xor2_1 _12549_ (.B(_05412_),
    .A(_05410_),
    .X(_05416_));
 sg13g2_a21oi_2 _12550_ (.B1(_05413_),
    .Y(_05417_),
    .A2(_05416_),
    .A1(_05414_));
 sg13g2_mux2_1 _12551_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.spike_out ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[1].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[879] ),
    .X(_05418_));
 sg13g2_nand2_1 _12552_ (.Y(_05419_),
    .A(\spiking_network_top_uut.all_data_out[311] ),
    .B(_05418_));
 sg13g2_mux2_1 _12553_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.spike_out ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[1].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[875] ),
    .X(_05420_));
 sg13g2_nand2_1 _12554_ (.Y(_05421_),
    .A(\spiking_network_top_uut.all_data_out[309] ),
    .B(_05420_));
 sg13g2_nor2_1 _12555_ (.A(_05419_),
    .B(_05421_),
    .Y(_05422_));
 sg13g2_nand2_1 _12556_ (.Y(_05423_),
    .A(\spiking_network_top_uut.all_data_out[310] ),
    .B(_05418_));
 sg13g2_nand2_1 _12557_ (.Y(_05424_),
    .A(\spiking_network_top_uut.all_data_out[308] ),
    .B(_05420_));
 sg13g2_or2_1 _12558_ (.X(_05425_),
    .B(_05424_),
    .A(_05423_));
 sg13g2_xor2_1 _12559_ (.B(_05421_),
    .A(_05419_),
    .X(_05426_));
 sg13g2_a21oi_2 _12560_ (.B1(_05422_),
    .Y(_05427_),
    .A2(_05426_),
    .A1(_05425_));
 sg13g2_mux2_2 _12561_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.spike_out ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[1].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[883] ),
    .X(_05428_));
 sg13g2_mux2_2 _12562_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.spike_out ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[1].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[887] ),
    .X(_05429_));
 sg13g2_a22oi_1 _12563_ (.Y(_05430_),
    .B1(_05429_),
    .B2(\spiking_network_top_uut.all_data_out[315] ),
    .A2(_05428_),
    .A1(\spiking_network_top_uut.all_data_out[313] ));
 sg13g2_and4_2 _12564_ (.A(\spiking_network_top_uut.all_data_out[312] ),
    .B(\spiking_network_top_uut.all_data_out[314] ),
    .C(_05428_),
    .D(_05429_),
    .X(_05431_));
 sg13g2_nand4_1 _12565_ (.B(\spiking_network_top_uut.all_data_out[314] ),
    .C(_05428_),
    .A(\spiking_network_top_uut.all_data_out[312] ),
    .Y(_05432_),
    .D(_05429_));
 sg13g2_and4_1 _12566_ (.A(\spiking_network_top_uut.all_data_out[313] ),
    .B(\spiking_network_top_uut.all_data_out[315] ),
    .C(_05428_),
    .D(_05429_),
    .X(_05433_));
 sg13g2_nand4_1 _12567_ (.B(\spiking_network_top_uut.all_data_out[315] ),
    .C(_05428_),
    .A(\spiking_network_top_uut.all_data_out[313] ),
    .Y(_05434_),
    .D(_05429_));
 sg13g2_nand3b_1 _12568_ (.B(_05431_),
    .C(_05434_),
    .Y(_05435_),
    .A_N(_05430_));
 sg13g2_a21oi_2 _12569_ (.B1(_05430_),
    .Y(_05436_),
    .A2(_05434_),
    .A1(_05431_));
 sg13g2_mux2_1 _12570_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.spike_out ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[1].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[895] ),
    .X(_05437_));
 sg13g2_mux2_2 _12571_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.spike_out ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[1].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[891] ),
    .X(_05438_));
 sg13g2_and4_1 _12572_ (.A(\spiking_network_top_uut.all_data_out[319] ),
    .B(\spiking_network_top_uut.all_data_out[317] ),
    .C(_05437_),
    .D(_05438_),
    .X(_05439_));
 sg13g2_nand4_1 _12573_ (.B(\spiking_network_top_uut.all_data_out[317] ),
    .C(_05437_),
    .A(\spiking_network_top_uut.all_data_out[319] ),
    .Y(_05440_),
    .D(_05438_));
 sg13g2_and4_1 _12574_ (.A(\spiking_network_top_uut.all_data_out[318] ),
    .B(\spiking_network_top_uut.all_data_out[316] ),
    .C(_05437_),
    .D(_05438_),
    .X(_05441_));
 sg13g2_a22oi_1 _12575_ (.Y(_05442_),
    .B1(_05438_),
    .B2(\spiking_network_top_uut.all_data_out[317] ),
    .A2(_05437_),
    .A1(\spiking_network_top_uut.all_data_out[319] ));
 sg13g2_or3_2 _12576_ (.A(_05439_),
    .B(_05441_),
    .C(_05442_),
    .X(_05443_));
 sg13g2_o21ai_1 _12577_ (.B1(_05440_),
    .Y(_05444_),
    .A1(_05441_),
    .A2(_05442_));
 sg13g2_nand3b_1 _12578_ (.B(_05436_),
    .C(_05444_),
    .Y(_05445_),
    .A_N(_05427_));
 sg13g2_inv_1 _12579_ (.Y(_05446_),
    .A(_05445_));
 sg13g2_or2_1 _12580_ (.X(_05447_),
    .B(_05445_),
    .A(_05417_));
 sg13g2_nor2_1 _12581_ (.A(_05436_),
    .B(_05444_),
    .Y(_05448_));
 sg13g2_and2_1 _12582_ (.A(_05427_),
    .B(_05448_),
    .X(_05449_));
 sg13g2_nand2_2 _12583_ (.Y(_05450_),
    .A(_05417_),
    .B(_05449_));
 sg13g2_and2_1 _12584_ (.A(_05447_),
    .B(_05450_),
    .X(_05451_));
 sg13g2_xnor2_1 _12585_ (.Y(_05452_),
    .A(_05388_),
    .B(_05405_));
 sg13g2_nand2_1 _12586_ (.Y(_05453_),
    .A(_05451_),
    .B(_05452_));
 sg13g2_nand2_1 _12587_ (.Y(_05454_),
    .A(_05447_),
    .B(_05453_));
 sg13g2_xor2_1 _12588_ (.B(_05451_),
    .A(_05407_),
    .X(_05455_));
 sg13g2_nand2_1 _12589_ (.Y(_05456_),
    .A(_05454_),
    .B(_05455_));
 sg13g2_xnor2_1 _12590_ (.Y(_05457_),
    .A(_05451_),
    .B(_05452_));
 sg13g2_o21ai_1 _12591_ (.B1(_05441_),
    .Y(_05458_),
    .A1(_05439_),
    .A2(_05442_));
 sg13g2_o21ai_1 _12592_ (.B1(_05432_),
    .Y(_05459_),
    .A1(_05430_),
    .A2(_05433_));
 sg13g2_o21ai_1 _12593_ (.B1(_05431_),
    .Y(_05460_),
    .A1(_05430_),
    .A2(_05433_));
 sg13g2_nand3b_1 _12594_ (.B(_05432_),
    .C(_05434_),
    .Y(_05461_),
    .A_N(_05430_));
 sg13g2_a22oi_1 _12595_ (.Y(_05462_),
    .B1(_05460_),
    .B2(_05461_),
    .A2(_05458_),
    .A1(_05443_));
 sg13g2_xor2_1 _12596_ (.B(_05426_),
    .A(_05425_),
    .X(_05463_));
 sg13g2_xnor2_1 _12597_ (.Y(_05464_),
    .A(_05425_),
    .B(_05426_));
 sg13g2_and4_1 _12598_ (.A(_05443_),
    .B(_05458_),
    .C(_05460_),
    .D(_05461_),
    .X(_05465_));
 sg13g2_nand4_1 _12599_ (.B(_05458_),
    .C(_05460_),
    .A(_05443_),
    .Y(_05466_),
    .D(_05461_));
 sg13g2_and4_1 _12600_ (.A(_05435_),
    .B(_05443_),
    .C(_05458_),
    .D(_05459_),
    .X(_05467_));
 sg13g2_a22oi_1 _12601_ (.Y(_05468_),
    .B1(_05459_),
    .B2(_05435_),
    .A2(_05458_),
    .A1(_05443_));
 sg13g2_nor3_2 _12602_ (.A(_05462_),
    .B(_05463_),
    .C(_05465_),
    .Y(_05469_));
 sg13g2_a21oi_2 _12603_ (.B1(_05462_),
    .Y(_05470_),
    .A2(_05466_),
    .A1(_05464_));
 sg13g2_xor2_1 _12604_ (.B(_05444_),
    .A(_05436_),
    .X(_05471_));
 sg13g2_xnor2_1 _12605_ (.Y(_05472_),
    .A(_05427_),
    .B(_05471_));
 sg13g2_nand2b_1 _12606_ (.Y(_05473_),
    .B(_05472_),
    .A_N(_05470_));
 sg13g2_xnor2_1 _12607_ (.Y(_05474_),
    .A(_05470_),
    .B(_05472_));
 sg13g2_nand2b_1 _12608_ (.Y(_05475_),
    .B(_05474_),
    .A_N(_05417_));
 sg13g2_nand2_2 _12609_ (.Y(_05476_),
    .A(_05473_),
    .B(_05475_));
 sg13g2_nor2_1 _12610_ (.A(_05446_),
    .B(_05449_),
    .Y(_05477_));
 sg13g2_xnor2_1 _12611_ (.Y(_05478_),
    .A(_05417_),
    .B(_05477_));
 sg13g2_and2_1 _12612_ (.A(_05476_),
    .B(_05478_),
    .X(_05479_));
 sg13g2_xor2_1 _12613_ (.B(_05478_),
    .A(_05476_),
    .X(_05480_));
 sg13g2_xnor2_1 _12614_ (.Y(_05481_),
    .A(_05403_),
    .B(_05404_));
 sg13g2_inv_1 _12615_ (.Y(_05482_),
    .A(_05481_));
 sg13g2_a21oi_1 _12616_ (.A1(_05480_),
    .A2(_05482_),
    .Y(_05483_),
    .B1(_05479_));
 sg13g2_nor2_1 _12617_ (.A(_05457_),
    .B(_05483_),
    .Y(_05484_));
 sg13g2_xnor2_1 _12618_ (.Y(_05485_),
    .A(_05480_),
    .B(_05481_));
 sg13g2_a22oi_1 _12619_ (.Y(_05486_),
    .B1(_05438_),
    .B2(\spiking_network_top_uut.all_data_out[316] ),
    .A2(_05437_),
    .A1(\spiking_network_top_uut.all_data_out[318] ));
 sg13g2_nor2_2 _12620_ (.A(_05441_),
    .B(_05486_),
    .Y(_05487_));
 sg13g2_a22oi_1 _12621_ (.Y(_05488_),
    .B1(_05429_),
    .B2(\spiking_network_top_uut.all_data_out[314] ),
    .A2(_05428_),
    .A1(\spiking_network_top_uut.all_data_out[312] ));
 sg13g2_nor2_1 _12622_ (.A(_05431_),
    .B(_05488_),
    .Y(_05489_));
 sg13g2_and2_1 _12623_ (.A(_05487_),
    .B(_05489_),
    .X(_05490_));
 sg13g2_xor2_1 _12624_ (.B(_05424_),
    .A(_05423_),
    .X(_05491_));
 sg13g2_xor2_1 _12625_ (.B(_05489_),
    .A(_05487_),
    .X(_05492_));
 sg13g2_a21oi_1 _12626_ (.A1(_05491_),
    .A2(_05492_),
    .Y(_05493_),
    .B1(_05490_));
 sg13g2_nor3_2 _12627_ (.A(_05464_),
    .B(_05467_),
    .C(_05468_),
    .Y(_05494_));
 sg13g2_nor3_1 _12628_ (.A(_05469_),
    .B(_05493_),
    .C(_05494_),
    .Y(_05495_));
 sg13g2_or3_1 _12629_ (.A(_05469_),
    .B(_05493_),
    .C(_05494_),
    .X(_05496_));
 sg13g2_xnor2_1 _12630_ (.Y(_05497_),
    .A(_05414_),
    .B(_05416_));
 sg13g2_o21ai_1 _12631_ (.B1(_05493_),
    .Y(_05498_),
    .A1(_05469_),
    .A2(_05494_));
 sg13g2_nand3_1 _12632_ (.B(_05497_),
    .C(_05498_),
    .A(_05496_),
    .Y(_05499_));
 sg13g2_a21o_2 _12633_ (.A2(_05498_),
    .A1(_05497_),
    .B1(_05495_),
    .X(_05500_));
 sg13g2_xnor2_1 _12634_ (.Y(_05501_),
    .A(_05417_),
    .B(_05474_));
 sg13g2_nand2_1 _12635_ (.Y(_05502_),
    .A(_05500_),
    .B(_05501_));
 sg13g2_xnor2_1 _12636_ (.Y(_05503_),
    .A(_05500_),
    .B(_05501_));
 sg13g2_xor2_1 _12637_ (.B(_05401_),
    .A(_05400_),
    .X(_05504_));
 sg13g2_o21ai_1 _12638_ (.B1(_05502_),
    .Y(_05505_),
    .A1(_05503_),
    .A2(_05504_));
 sg13g2_nand2_1 _12639_ (.Y(_05506_),
    .A(_05485_),
    .B(_05505_));
 sg13g2_xor2_1 _12640_ (.B(_05504_),
    .A(_05503_),
    .X(_05507_));
 sg13g2_a22oi_1 _12641_ (.Y(_05508_),
    .B1(_05411_),
    .B2(\spiking_network_top_uut.all_data_out[306] ),
    .A2(_05409_),
    .A1(\spiking_network_top_uut.all_data_out[304] ));
 sg13g2_xnor2_1 _12642_ (.Y(_05509_),
    .A(_05491_),
    .B(_05492_));
 sg13g2_nor3_2 _12643_ (.A(_05415_),
    .B(_05508_),
    .C(_05509_),
    .Y(_05510_));
 sg13g2_a21o_2 _12644_ (.A2(_05498_),
    .A1(_05496_),
    .B1(_05497_),
    .X(_05511_));
 sg13g2_nand3_1 _12645_ (.B(_05510_),
    .C(_05511_),
    .A(_05499_),
    .Y(_05512_));
 sg13g2_a21oi_1 _12646_ (.A1(_05499_),
    .A2(_05511_),
    .Y(_05513_),
    .B1(_05510_));
 sg13g2_a21o_1 _12647_ (.A2(_05511_),
    .A1(_05499_),
    .B1(_05510_),
    .X(_05514_));
 sg13g2_xnor2_1 _12648_ (.Y(_05515_),
    .A(_05398_),
    .B(_05399_));
 sg13g2_inv_1 _12649_ (.Y(_05516_),
    .A(_05515_));
 sg13g2_and3_1 _12650_ (.X(_05517_),
    .A(_05512_),
    .B(_05514_),
    .C(_05516_));
 sg13g2_o21ai_1 _12651_ (.B1(_05512_),
    .Y(_05518_),
    .A1(_05513_),
    .A2(_05515_));
 sg13g2_and2_1 _12652_ (.A(_05507_),
    .B(_05518_),
    .X(_05519_));
 sg13g2_a21oi_1 _12653_ (.A1(_05512_),
    .A2(_05514_),
    .Y(_05520_),
    .B1(_05516_));
 sg13g2_nor2_1 _12654_ (.A(_05517_),
    .B(_05520_),
    .Y(_05521_));
 sg13g2_xnor2_1 _12655_ (.Y(_05522_),
    .A(_00040_),
    .B(_05397_));
 sg13g2_o21ai_1 _12656_ (.B1(_05509_),
    .Y(_05523_),
    .A1(_05415_),
    .A2(_05508_));
 sg13g2_nand2b_2 _12657_ (.Y(_05524_),
    .B(_05523_),
    .A_N(_05510_));
 sg13g2_nor2_1 _12658_ (.A(_05522_),
    .B(_05524_),
    .Y(_05525_));
 sg13g2_nor4_2 _12659_ (.A(_05517_),
    .B(_05520_),
    .C(_05522_),
    .Y(_05526_),
    .D(_05524_));
 sg13g2_xor2_1 _12660_ (.B(_05518_),
    .A(_05507_),
    .X(_05527_));
 sg13g2_a21oi_1 _12661_ (.A1(_05526_),
    .A2(_05527_),
    .Y(_05528_),
    .B1(_05519_));
 sg13g2_xnor2_1 _12662_ (.Y(_05529_),
    .A(_05485_),
    .B(_05505_));
 sg13g2_o21ai_1 _12663_ (.B1(_05506_),
    .Y(_05530_),
    .A1(_05528_),
    .A2(_05529_));
 sg13g2_nand2_1 _12664_ (.Y(_05531_),
    .A(_05457_),
    .B(_05483_));
 sg13g2_nand2b_1 _12665_ (.Y(_05532_),
    .B(_05531_),
    .A_N(_05484_));
 sg13g2_a21oi_1 _12666_ (.A1(_05530_),
    .A2(_05531_),
    .Y(_05533_),
    .B1(_05484_));
 sg13g2_xnor2_1 _12667_ (.Y(_05534_),
    .A(_05454_),
    .B(_05455_));
 sg13g2_o21ai_1 _12668_ (.B1(_05456_),
    .Y(_05535_),
    .A1(_05533_),
    .A2(_05534_));
 sg13g2_mux2_1 _12669_ (.A0(_05450_),
    .A1(_05447_),
    .S(_05407_),
    .X(_05536_));
 sg13g2_xnor2_1 _12670_ (.Y(_05537_),
    .A(_05535_),
    .B(_05536_));
 sg13g2_a21oi_2 _12671_ (.B1(_05408_),
    .Y(_05538_),
    .A2(_05537_),
    .A1(_05363_));
 sg13g2_xnor2_1 _12672_ (.Y(_05539_),
    .A(_05533_),
    .B(_05534_));
 sg13g2_a21oi_1 _12673_ (.A1(_05363_),
    .A2(_05539_),
    .Y(_05540_),
    .B1(_05408_));
 sg13g2_nand2_1 _12674_ (.Y(_05541_),
    .A(_05364_),
    .B(_05452_));
 sg13g2_xor2_1 _12675_ (.B(_05532_),
    .A(_05530_),
    .X(_05542_));
 sg13g2_o21ai_1 _12676_ (.B1(_05541_),
    .Y(_05543_),
    .A1(_05364_),
    .A2(_05542_));
 sg13g2_nand2_1 _12677_ (.Y(_05544_),
    .A(_05540_),
    .B(_05543_));
 sg13g2_a21oi_2 _12678_ (.B1(net3631),
    .Y(_05545_),
    .A2(_05544_),
    .A1(_05538_));
 sg13g2_nor2_1 _12679_ (.A(_05540_),
    .B(_05543_),
    .Y(_05546_));
 sg13g2_nor2_2 _12680_ (.A(_05538_),
    .B(_05546_),
    .Y(_05547_));
 sg13g2_nor2_1 _12681_ (.A(_05364_),
    .B(_05524_),
    .Y(_05548_));
 sg13g2_xnor2_1 _12682_ (.Y(_05549_),
    .A(_05522_),
    .B(_05548_));
 sg13g2_o21ai_1 _12683_ (.B1(_05545_),
    .Y(_05550_),
    .A1(_05547_),
    .A2(_05549_));
 sg13g2_xor2_1 _12684_ (.B(net464),
    .A(net4311),
    .X(_05551_));
 sg13g2_a21oi_1 _12685_ (.A1(net3631),
    .A2(_05551_),
    .Y(_05552_),
    .B1(net3941));
 sg13g2_a22oi_1 _12686_ (.Y(_00536_),
    .B1(_05550_),
    .B2(_05552_),
    .A2(net3941),
    .A1(_03407_));
 sg13g2_nor2_1 _12687_ (.A(_05364_),
    .B(_05526_),
    .Y(_05553_));
 sg13g2_o21ai_1 _12688_ (.B1(_05553_),
    .Y(_05554_),
    .A1(_05521_),
    .A2(_05525_));
 sg13g2_o21ai_1 _12689_ (.B1(_05554_),
    .Y(_05555_),
    .A1(_05363_),
    .A2(_05515_));
 sg13g2_o21ai_1 _12690_ (.B1(_05545_),
    .Y(_05556_),
    .A1(_05547_),
    .A2(_05555_));
 sg13g2_xor2_1 _12691_ (.B(_04737_),
    .A(_04736_),
    .X(_05557_));
 sg13g2_a21oi_1 _12692_ (.A1(net3631),
    .A2(_05557_),
    .Y(_05558_),
    .B1(net3940));
 sg13g2_a22oi_1 _12693_ (.Y(_00537_),
    .B1(_05556_),
    .B2(_05558_),
    .A2(net3940),
    .A1(_03408_));
 sg13g2_and2_1 _12694_ (.A(_05364_),
    .B(_05504_),
    .X(_05559_));
 sg13g2_xnor2_1 _12695_ (.Y(_05560_),
    .A(_05526_),
    .B(_05527_));
 sg13g2_a21oi_1 _12696_ (.A1(_05363_),
    .A2(_05560_),
    .Y(_05561_),
    .B1(_05559_));
 sg13g2_o21ai_1 _12697_ (.B1(_05545_),
    .Y(_05562_),
    .A1(_05547_),
    .A2(_05561_));
 sg13g2_xnor2_1 _12698_ (.Y(_05563_),
    .A(_04734_),
    .B(_04738_));
 sg13g2_a21oi_1 _12699_ (.A1(net3631),
    .A2(_05563_),
    .Y(_05564_),
    .B1(net3940));
 sg13g2_a22oi_1 _12700_ (.Y(_00538_),
    .B1(_05562_),
    .B2(_05564_),
    .A2(net3940),
    .A1(_03410_));
 sg13g2_xor2_1 _12701_ (.B(_05529_),
    .A(_05528_),
    .X(_05565_));
 sg13g2_mux2_1 _12702_ (.A0(_05482_),
    .A1(_05565_),
    .S(_05363_),
    .X(_05566_));
 sg13g2_o21ai_1 _12703_ (.B1(_05545_),
    .Y(_05567_),
    .A1(_05547_),
    .A2(_05566_));
 sg13g2_or3_1 _12704_ (.A(_04732_),
    .B(_04733_),
    .C(_04739_),
    .X(_05568_));
 sg13g2_and2_1 _12705_ (.A(_04740_),
    .B(_05568_),
    .X(_05569_));
 sg13g2_a21oi_1 _12706_ (.A1(net3631),
    .A2(_05569_),
    .Y(_05570_),
    .B1(net3940));
 sg13g2_a22oi_1 _12707_ (.Y(_00539_),
    .B1(_05567_),
    .B2(_05570_),
    .A2(net3940),
    .A1(_03409_));
 sg13g2_nand2b_1 _12708_ (.Y(_05571_),
    .B(_05538_),
    .A_N(net3631));
 sg13g2_a21oi_1 _12709_ (.A1(_04731_),
    .A2(_04741_),
    .Y(_05572_),
    .B1(net3940));
 sg13g2_a22oi_1 _12710_ (.Y(_00540_),
    .B1(_05571_),
    .B2(_05572_),
    .A2(net3940),
    .A1(_03411_));
 sg13g2_mux4_1 _12711_ (.S0(\spiking_network_top_uut.all_data_out[604] ),
    .A0(net3846),
    .A1(net3845),
    .A2(net3844),
    .A3(net3843),
    .S1(\spiking_network_top_uut.all_data_out[605] ),
    .X(_05573_));
 sg13g2_mux2_1 _12712_ (.A0(net3841),
    .A1(net3900),
    .S(\spiking_network_top_uut.all_data_out[604] ),
    .X(_05574_));
 sg13g2_nor2b_1 _12713_ (.A(\spiking_network_top_uut.all_data_out[604] ),
    .B_N(net3842),
    .Y(_05575_));
 sg13g2_a21oi_1 _12714_ (.A1(\spiking_network_top_uut.all_data_out[604] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[5] ),
    .Y(_05576_),
    .B1(_05575_));
 sg13g2_o21ai_1 _12715_ (.B1(\spiking_network_top_uut.all_data_out[606] ),
    .Y(_05577_),
    .A1(\spiking_network_top_uut.all_data_out[605] ),
    .A2(_05576_));
 sg13g2_a21oi_1 _12716_ (.A1(\spiking_network_top_uut.all_data_out[605] ),
    .A2(_05574_),
    .Y(_05578_),
    .B1(_05577_));
 sg13g2_o21ai_1 _12717_ (.B1(net4551),
    .Y(_05579_),
    .A1(\spiking_network_top_uut.all_data_out[606] ),
    .A2(_05573_));
 sg13g2_nand2_1 _12718_ (.Y(_05580_),
    .A(net3934),
    .B(net181));
 sg13g2_o21ai_1 _12719_ (.B1(_05580_),
    .Y(_00541_),
    .A1(_05578_),
    .A2(_05579_));
 sg13g2_mux2_1 _12720_ (.A0(net314),
    .A1(net181),
    .S(net4553),
    .X(_00542_));
 sg13g2_mux4_1 _12721_ (.S0(\spiking_network_top_uut.all_data_out[600] ),
    .A0(net3898),
    .A1(net3897),
    .A2(net3896),
    .A3(net3895),
    .S1(\spiking_network_top_uut.all_data_out[601] ),
    .X(_05581_));
 sg13g2_mux2_1 _12722_ (.A0(net3893),
    .A1(net3892),
    .S(\spiking_network_top_uut.all_data_out[600] ),
    .X(_05582_));
 sg13g2_nor2b_1 _12723_ (.A(\spiking_network_top_uut.all_data_out[600] ),
    .B_N(net3894),
    .Y(_05583_));
 sg13g2_a21oi_1 _12724_ (.A1(\spiking_network_top_uut.all_data_out[600] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[5] ),
    .Y(_05584_),
    .B1(_05583_));
 sg13g2_o21ai_1 _12725_ (.B1(\spiking_network_top_uut.all_data_out[602] ),
    .Y(_05585_),
    .A1(\spiking_network_top_uut.all_data_out[601] ),
    .A2(_05584_));
 sg13g2_a21oi_1 _12726_ (.A1(\spiking_network_top_uut.all_data_out[601] ),
    .A2(_05582_),
    .Y(_05586_),
    .B1(_05585_));
 sg13g2_o21ai_1 _12727_ (.B1(net4545),
    .Y(_05587_),
    .A1(\spiking_network_top_uut.all_data_out[602] ),
    .A2(_05581_));
 sg13g2_nand2_1 _12728_ (.Y(_05588_),
    .A(net3933),
    .B(net57));
 sg13g2_o21ai_1 _12729_ (.B1(_05588_),
    .Y(_00543_),
    .A1(_05586_),
    .A2(_05587_));
 sg13g2_mux2_1 _12730_ (.A0(net257),
    .A1(net57),
    .S(net4544),
    .X(_00544_));
 sg13g2_a21oi_1 _12731_ (.A1(\spiking_network_top_uut.all_data_out[596] ),
    .A2(_03665_),
    .Y(_05589_),
    .B1(\spiking_network_top_uut.all_data_out[597] ));
 sg13g2_o21ai_1 _12732_ (.B1(_05589_),
    .Y(_05590_),
    .A1(\spiking_network_top_uut.all_data_out[596] ),
    .A2(net3887));
 sg13g2_mux2_1 _12733_ (.A0(net3886),
    .A1(net3885),
    .S(\spiking_network_top_uut.all_data_out[596] ),
    .X(_05591_));
 sg13g2_nand2_1 _12734_ (.Y(_05592_),
    .A(\spiking_network_top_uut.all_data_out[597] ),
    .B(_05591_));
 sg13g2_nand3_1 _12735_ (.B(_05590_),
    .C(_05592_),
    .A(\spiking_network_top_uut.all_data_out[598] ),
    .Y(_05593_));
 sg13g2_mux2_1 _12736_ (.A0(net3889),
    .A1(net3888),
    .S(\spiking_network_top_uut.all_data_out[596] ),
    .X(_05594_));
 sg13g2_nor2b_1 _12737_ (.A(\spiking_network_top_uut.all_data_out[596] ),
    .B_N(net3891),
    .Y(_05595_));
 sg13g2_a21oi_1 _12738_ (.A1(\spiking_network_top_uut.all_data_out[596] ),
    .A2(net3890),
    .Y(_05596_),
    .B1(_05595_));
 sg13g2_a21oi_1 _12739_ (.A1(\spiking_network_top_uut.all_data_out[597] ),
    .A2(_05594_),
    .Y(_05597_),
    .B1(\spiking_network_top_uut.all_data_out[598] ));
 sg13g2_o21ai_1 _12740_ (.B1(_05597_),
    .Y(_05598_),
    .A1(\spiking_network_top_uut.all_data_out[597] ),
    .A2(_05596_));
 sg13g2_nand3_1 _12741_ (.B(_05593_),
    .C(_05598_),
    .A(net4558),
    .Y(_05599_));
 sg13g2_o21ai_1 _12742_ (.B1(_05599_),
    .Y(_00545_),
    .A1(net4558),
    .A2(_03670_));
 sg13g2_nor2_1 _12743_ (.A(net4558),
    .B(net179),
    .Y(_05600_));
 sg13g2_a21oi_1 _12744_ (.A1(net4558),
    .A2(_03670_),
    .Y(_00546_),
    .B1(_05600_));
 sg13g2_mux4_1 _12745_ (.S0(\spiking_network_top_uut.all_data_out[592] ),
    .A0(net3884),
    .A1(net3883),
    .A2(net3882),
    .A3(net3881),
    .S1(\spiking_network_top_uut.all_data_out[593] ),
    .X(_05601_));
 sg13g2_mux2_1 _12746_ (.A0(net3878),
    .A1(net3877),
    .S(\spiking_network_top_uut.all_data_out[592] ),
    .X(_05602_));
 sg13g2_nor2b_1 _12747_ (.A(\spiking_network_top_uut.all_data_out[592] ),
    .B_N(net3880),
    .Y(_05603_));
 sg13g2_a21oi_1 _12748_ (.A1(\spiking_network_top_uut.all_data_out[592] ),
    .A2(net3879),
    .Y(_05604_),
    .B1(_05603_));
 sg13g2_o21ai_1 _12749_ (.B1(\spiking_network_top_uut.all_data_out[594] ),
    .Y(_05605_),
    .A1(\spiking_network_top_uut.all_data_out[593] ),
    .A2(_05604_));
 sg13g2_a21oi_1 _12750_ (.A1(\spiking_network_top_uut.all_data_out[593] ),
    .A2(_05602_),
    .Y(_05606_),
    .B1(_05605_));
 sg13g2_o21ai_1 _12751_ (.B1(net4557),
    .Y(_05607_),
    .A1(\spiking_network_top_uut.all_data_out[594] ),
    .A2(_05601_));
 sg13g2_nand2_1 _12752_ (.Y(_05608_),
    .A(net3938),
    .B(net187));
 sg13g2_o21ai_1 _12753_ (.B1(_05608_),
    .Y(_00547_),
    .A1(_05606_),
    .A2(_05607_));
 sg13g2_mux2_1 _12754_ (.A0(net279),
    .A1(net187),
    .S(net4557),
    .X(_00548_));
 sg13g2_mux2_1 _12755_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[2] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[3] ),
    .S(\spiking_network_top_uut.all_data_out[588] ),
    .X(_05609_));
 sg13g2_nor2b_1 _12756_ (.A(\spiking_network_top_uut.all_data_out[588] ),
    .B_N(net3876),
    .Y(_05610_));
 sg13g2_a21oi_1 _12757_ (.A1(\spiking_network_top_uut.all_data_out[588] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[1] ),
    .Y(_05611_),
    .B1(_05610_));
 sg13g2_a21oi_1 _12758_ (.A1(\spiking_network_top_uut.all_data_out[589] ),
    .A2(_05609_),
    .Y(_05612_),
    .B1(\spiking_network_top_uut.all_data_out[590] ));
 sg13g2_o21ai_1 _12759_ (.B1(_05612_),
    .Y(_05613_),
    .A1(\spiking_network_top_uut.all_data_out[589] ),
    .A2(_05611_));
 sg13g2_mux2_1 _12760_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[6] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[7] ),
    .S(\spiking_network_top_uut.all_data_out[588] ),
    .X(_05614_));
 sg13g2_nor2b_1 _12761_ (.A(\spiking_network_top_uut.all_data_out[588] ),
    .B_N(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[4] ),
    .Y(_05615_));
 sg13g2_a21oi_1 _12762_ (.A1(\spiking_network_top_uut.all_data_out[588] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[5] ),
    .Y(_05616_),
    .B1(_05615_));
 sg13g2_o21ai_1 _12763_ (.B1(\spiking_network_top_uut.all_data_out[590] ),
    .Y(_05617_),
    .A1(\spiking_network_top_uut.all_data_out[589] ),
    .A2(_05616_));
 sg13g2_a21oi_1 _12764_ (.A1(\spiking_network_top_uut.all_data_out[589] ),
    .A2(_05614_),
    .Y(_05618_),
    .B1(_05617_));
 sg13g2_nand2_1 _12765_ (.Y(_05619_),
    .A(net4569),
    .B(_05613_));
 sg13g2_nand2_1 _12766_ (.Y(_05620_),
    .A(net3939),
    .B(net155));
 sg13g2_o21ai_1 _12767_ (.B1(_05620_),
    .Y(_00549_),
    .A1(_05618_),
    .A2(_05619_));
 sg13g2_mux2_1 _12768_ (.A0(net319),
    .A1(net155),
    .S(net4569),
    .X(_00550_));
 sg13g2_mux4_1 _12769_ (.S0(\spiking_network_top_uut.all_data_out[584] ),
    .A0(net3868),
    .A1(net3867),
    .A2(net3866),
    .A3(net3865),
    .S1(\spiking_network_top_uut.all_data_out[585] ),
    .X(_05621_));
 sg13g2_mux2_1 _12770_ (.A0(net3862),
    .A1(net3861),
    .S(\spiking_network_top_uut.all_data_out[584] ),
    .X(_05622_));
 sg13g2_nor2b_1 _12771_ (.A(\spiking_network_top_uut.all_data_out[584] ),
    .B_N(net3864),
    .Y(_05623_));
 sg13g2_a21oi_1 _12772_ (.A1(\spiking_network_top_uut.all_data_out[584] ),
    .A2(net3863),
    .Y(_05624_),
    .B1(_05623_));
 sg13g2_o21ai_1 _12773_ (.B1(\spiking_network_top_uut.all_data_out[586] ),
    .Y(_05625_),
    .A1(\spiking_network_top_uut.all_data_out[585] ),
    .A2(_05624_));
 sg13g2_a21oi_1 _12774_ (.A1(\spiking_network_top_uut.all_data_out[585] ),
    .A2(_05622_),
    .Y(_05626_),
    .B1(_05625_));
 sg13g2_o21ai_1 _12775_ (.B1(net4563),
    .Y(_05627_),
    .A1(\spiking_network_top_uut.all_data_out[586] ),
    .A2(_05621_));
 sg13g2_nand2_1 _12776_ (.Y(_05628_),
    .A(net3936),
    .B(net164));
 sg13g2_o21ai_1 _12777_ (.B1(_05628_),
    .Y(_00551_),
    .A1(_05626_),
    .A2(_05627_));
 sg13g2_mux2_1 _12778_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_dout ),
    .A1(net164),
    .S(net4563),
    .X(_00552_));
 sg13g2_mux4_1 _12779_ (.S0(\spiking_network_top_uut.all_data_out[580] ),
    .A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[0] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[1] ),
    .A2(net3858),
    .A3(net3857),
    .S1(\spiking_network_top_uut.all_data_out[581] ),
    .X(_05629_));
 sg13g2_mux2_1 _12780_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[6] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[7] ),
    .S(\spiking_network_top_uut.all_data_out[580] ),
    .X(_05630_));
 sg13g2_nor2b_1 _12781_ (.A(\spiking_network_top_uut.all_data_out[580] ),
    .B_N(net3856),
    .Y(_05631_));
 sg13g2_a21oi_1 _12782_ (.A1(\spiking_network_top_uut.all_data_out[580] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[5] ),
    .Y(_05632_),
    .B1(_05631_));
 sg13g2_o21ai_1 _12783_ (.B1(\spiking_network_top_uut.all_data_out[582] ),
    .Y(_05633_),
    .A1(\spiking_network_top_uut.all_data_out[581] ),
    .A2(_05632_));
 sg13g2_a21oi_1 _12784_ (.A1(\spiking_network_top_uut.all_data_out[581] ),
    .A2(_05630_),
    .Y(_05634_),
    .B1(_05633_));
 sg13g2_o21ai_1 _12785_ (.B1(net4540),
    .Y(_05635_),
    .A1(\spiking_network_top_uut.all_data_out[582] ),
    .A2(_05629_));
 sg13g2_nand2_1 _12786_ (.Y(_05636_),
    .A(net3932),
    .B(net75));
 sg13g2_o21ai_1 _12787_ (.B1(_05636_),
    .Y(_00553_),
    .A1(_05634_),
    .A2(_05635_));
 sg13g2_mux2_1 _12788_ (.A0(net226),
    .A1(net75),
    .S(net4541),
    .X(_00554_));
 sg13g2_mux4_1 _12789_ (.S0(\spiking_network_top_uut.all_data_out[576] ),
    .A0(net3853),
    .A1(net3852),
    .A2(net3851),
    .A3(net3850),
    .S1(\spiking_network_top_uut.all_data_out[577] ),
    .X(_05637_));
 sg13g2_mux2_1 _12790_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[6] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[7] ),
    .S(\spiking_network_top_uut.all_data_out[576] ),
    .X(_05638_));
 sg13g2_nor2b_1 _12791_ (.A(\spiking_network_top_uut.all_data_out[576] ),
    .B_N(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[4] ),
    .Y(_05639_));
 sg13g2_a21oi_1 _12792_ (.A1(\spiking_network_top_uut.all_data_out[576] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[5] ),
    .Y(_05640_),
    .B1(_05639_));
 sg13g2_o21ai_1 _12793_ (.B1(\spiking_network_top_uut.all_data_out[578] ),
    .Y(_05641_),
    .A1(\spiking_network_top_uut.all_data_out[577] ),
    .A2(_05640_));
 sg13g2_a21oi_1 _12794_ (.A1(\spiking_network_top_uut.all_data_out[577] ),
    .A2(_05638_),
    .Y(_05642_),
    .B1(_05641_));
 sg13g2_o21ai_1 _12795_ (.B1(net4543),
    .Y(_05643_),
    .A1(\spiking_network_top_uut.all_data_out[578] ),
    .A2(_05637_));
 sg13g2_nand2_1 _12796_ (.Y(_05644_),
    .A(net3933),
    .B(net93));
 sg13g2_o21ai_1 _12797_ (.B1(_05644_),
    .Y(_00555_),
    .A1(_05642_),
    .A2(_05643_));
 sg13g2_nor3_2 _12798_ (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[2] ),
    .B(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[1] ),
    .C(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[0] ),
    .Y(_05645_));
 sg13g2_nor2b_2 _12799_ (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[3] ),
    .B_N(_05645_),
    .Y(_05646_));
 sg13g2_nor2b_2 _12800_ (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[4] ),
    .B_N(_05646_),
    .Y(_05647_));
 sg13g2_nand2b_2 _12801_ (.Y(_05648_),
    .B(_05646_),
    .A_N(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[4] ));
 sg13g2_o21ai_1 _12802_ (.B1(net4529),
    .Y(_05649_),
    .A1(net3660),
    .A2(_05648_));
 sg13g2_nor2b_1 _12803_ (.A(net3659),
    .B_N(_00048_),
    .Y(_05650_));
 sg13g2_a21oi_1 _12804_ (.A1(net4283),
    .A2(net3659),
    .Y(_05651_),
    .B1(_05650_));
 sg13g2_nand2_1 _12805_ (.Y(_05652_),
    .A(net375),
    .B(_05649_));
 sg13g2_o21ai_1 _12806_ (.B1(_05652_),
    .Y(_00556_),
    .A1(_05649_),
    .A2(_05651_));
 sg13g2_xor2_1 _12807_ (.B(net375),
    .A(net392),
    .X(_05653_));
 sg13g2_nor2_1 _12808_ (.A(net3659),
    .B(_05653_),
    .Y(_05654_));
 sg13g2_a21oi_1 _12809_ (.A1(net4280),
    .A2(net3659),
    .Y(_05655_),
    .B1(_05654_));
 sg13g2_nand2_1 _12810_ (.Y(_05656_),
    .A(net392),
    .B(_05649_));
 sg13g2_o21ai_1 _12811_ (.B1(_05656_),
    .Y(_00557_),
    .A1(_05649_),
    .A2(_05655_));
 sg13g2_o21ai_1 _12812_ (.B1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[2] ),
    .Y(_05657_),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[1] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[0] ));
 sg13g2_nor2b_1 _12813_ (.A(_05645_),
    .B_N(_05657_),
    .Y(_05658_));
 sg13g2_nor2_1 _12814_ (.A(net3659),
    .B(_05658_),
    .Y(_05659_));
 sg13g2_a21oi_1 _12815_ (.A1(net4276),
    .A2(net3659),
    .Y(_05660_),
    .B1(_05659_));
 sg13g2_nand2_1 _12816_ (.Y(_05661_),
    .A(net153),
    .B(_05649_));
 sg13g2_o21ai_1 _12817_ (.B1(_05661_),
    .Y(_00558_),
    .A1(_05649_),
    .A2(_05660_));
 sg13g2_nand2_1 _12818_ (.Y(_05662_),
    .A(net4273),
    .B(net3659));
 sg13g2_xnor2_1 _12819_ (.Y(_05663_),
    .A(net417),
    .B(_05645_));
 sg13g2_o21ai_1 _12820_ (.B1(_05662_),
    .Y(_05664_),
    .A1(net3659),
    .A2(_05663_));
 sg13g2_mux2_1 _12821_ (.A0(_05664_),
    .A1(net417),
    .S(_05649_),
    .X(_00559_));
 sg13g2_nand2_1 _12822_ (.Y(_05665_),
    .A(net3922),
    .B(net293));
 sg13g2_nand2b_1 _12823_ (.Y(_05666_),
    .B(net293),
    .A_N(_05646_));
 sg13g2_a21oi_1 _12824_ (.A1(_05648_),
    .A2(_05666_),
    .Y(_05667_),
    .B1(net3660));
 sg13g2_a21oi_1 _12825_ (.A1(net4269),
    .A2(net3660),
    .Y(_05668_),
    .B1(_05667_));
 sg13g2_o21ai_1 _12826_ (.B1(_05665_),
    .Y(_00560_),
    .A1(_05649_),
    .A2(_05668_));
 sg13g2_mux2_1 _12827_ (.A0(net273),
    .A1(net93),
    .S(net4543),
    .X(_00561_));
 sg13g2_mux2_1 _12828_ (.A0(net3899),
    .A1(net3783),
    .S(net4637),
    .X(_00562_));
 sg13g2_a21oi_1 _12829_ (.A1(net3915),
    .A2(net3911),
    .Y(_05669_),
    .B1(_00043_));
 sg13g2_nor2_2 _12830_ (.A(net3755),
    .B(_05669_),
    .Y(_05670_));
 sg13g2_nand2b_1 _12831_ (.Y(_05671_),
    .B(_05670_),
    .A_N(_00043_));
 sg13g2_o21ai_1 _12832_ (.B1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ),
    .Y(_05672_),
    .A1(_00043_),
    .A2(_05670_));
 sg13g2_a21o_1 _12833_ (.A2(net3755),
    .A1(_00044_),
    .B1(_05670_),
    .X(_05673_));
 sg13g2_nor2_1 _12834_ (.A(_03479_),
    .B(net3918),
    .Y(_05674_));
 sg13g2_o21ai_1 _12835_ (.B1(net3918),
    .Y(_05675_),
    .A1(_00044_),
    .A2(net3907));
 sg13g2_a21oi_1 _12836_ (.A1(net3907),
    .A2(_05669_),
    .Y(_05676_),
    .B1(_05675_));
 sg13g2_o21ai_1 _12837_ (.B1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ),
    .Y(_05677_),
    .A1(_05674_),
    .A2(_05676_));
 sg13g2_or2_1 _12838_ (.X(_05678_),
    .B(net3918),
    .A(_00047_));
 sg13g2_o21ai_1 _12839_ (.B1(net3915),
    .Y(_05679_),
    .A1(_00043_),
    .A2(net3911));
 sg13g2_or2_1 _12840_ (.X(_05680_),
    .B(net3907),
    .A(_03479_));
 sg13g2_nand2_1 _12841_ (.Y(_05681_),
    .A(_00044_),
    .B(net3902));
 sg13g2_nand4_1 _12842_ (.B(_05679_),
    .C(_05680_),
    .A(net3918),
    .Y(_05682_),
    .D(_05681_));
 sg13g2_and2_1 _12843_ (.A(_05678_),
    .B(_05682_),
    .X(_05683_));
 sg13g2_a21oi_1 _12844_ (.A1(_05678_),
    .A2(_05682_),
    .Y(_05684_),
    .B1(_03480_));
 sg13g2_nor3_1 _12845_ (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ),
    .B(_05674_),
    .C(_05676_),
    .Y(_05685_));
 sg13g2_or3_1 _12846_ (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ),
    .B(_05674_),
    .C(_05676_),
    .X(_05686_));
 sg13g2_nand2_1 _12847_ (.Y(_05687_),
    .A(_05677_),
    .B(_05686_));
 sg13g2_o21ai_1 _12848_ (.B1(_05677_),
    .Y(_05688_),
    .A1(_05684_),
    .A2(_05685_));
 sg13g2_xnor2_1 _12849_ (.Y(_05689_),
    .A(_03479_),
    .B(_05673_));
 sg13g2_nor2b_1 _12850_ (.A(_05689_),
    .B_N(_05688_),
    .Y(_05690_));
 sg13g2_a21o_1 _12851_ (.A2(_05673_),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ),
    .B1(_05690_),
    .X(_05691_));
 sg13g2_or3_1 _12852_ (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ),
    .B(_00043_),
    .C(_05670_),
    .X(_05692_));
 sg13g2_and2_1 _12853_ (.A(_05672_),
    .B(_05692_),
    .X(_05693_));
 sg13g2_nand2_1 _12854_ (.Y(_05694_),
    .A(_05691_),
    .B(_05693_));
 sg13g2_and2_1 _12855_ (.A(_05672_),
    .B(_05694_),
    .X(_05695_));
 sg13g2_a22oi_1 _12856_ (.Y(_05696_),
    .B1(_05671_),
    .B2(_05695_),
    .A2(_05670_),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ));
 sg13g2_a21oi_2 _12857_ (.B1(_05696_),
    .Y(_05697_),
    .A2(_00043_),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ));
 sg13g2_mux2_1 _12858_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.spike_out ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[579] ),
    .X(_05698_));
 sg13g2_nand2_1 _12859_ (.Y(_05699_),
    .A(\spiking_network_top_uut.all_data_out[161] ),
    .B(_05698_));
 sg13g2_mux2_2 _12860_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.spike_out ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[583] ),
    .X(_05700_));
 sg13g2_nand2_1 _12861_ (.Y(_05701_),
    .A(\spiking_network_top_uut.all_data_out[163] ),
    .B(_05700_));
 sg13g2_nor2_1 _12862_ (.A(_05699_),
    .B(_05701_),
    .Y(_05702_));
 sg13g2_nand4_1 _12863_ (.B(\spiking_network_top_uut.all_data_out[162] ),
    .C(_05698_),
    .A(\spiking_network_top_uut.all_data_out[160] ),
    .Y(_05703_),
    .D(_05700_));
 sg13g2_inv_1 _12864_ (.Y(_05704_),
    .A(_05703_));
 sg13g2_xor2_1 _12865_ (.B(_05701_),
    .A(_05699_),
    .X(_05705_));
 sg13g2_a21oi_2 _12866_ (.B1(_05702_),
    .Y(_05706_),
    .A2(_05705_),
    .A1(_05703_));
 sg13g2_mux2_2 _12867_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.spike_out ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[587] ),
    .X(_05707_));
 sg13g2_nand2_1 _12868_ (.Y(_05708_),
    .A(\spiking_network_top_uut.all_data_out[165] ),
    .B(_05707_));
 sg13g2_mux2_2 _12869_ (.A0(net4596),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[591] ),
    .X(_05709_));
 sg13g2_nand2_1 _12870_ (.Y(_05710_),
    .A(\spiking_network_top_uut.all_data_out[167] ),
    .B(_05709_));
 sg13g2_nor2_1 _12871_ (.A(_05708_),
    .B(_05710_),
    .Y(_05711_));
 sg13g2_nand2_1 _12872_ (.Y(_05712_),
    .A(\spiking_network_top_uut.all_data_out[164] ),
    .B(_05707_));
 sg13g2_nand2_1 _12873_ (.Y(_05713_),
    .A(\spiking_network_top_uut.all_data_out[166] ),
    .B(_05709_));
 sg13g2_or2_1 _12874_ (.X(_05714_),
    .B(_05713_),
    .A(_05712_));
 sg13g2_xor2_1 _12875_ (.B(_05710_),
    .A(_05708_),
    .X(_05715_));
 sg13g2_a21oi_2 _12876_ (.B1(_05711_),
    .Y(_05716_),
    .A2(_05715_),
    .A1(_05714_));
 sg13g2_mux2_2 _12877_ (.A0(net4595),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[595] ),
    .X(_05717_));
 sg13g2_mux2_2 _12878_ (.A0(net4594),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[599] ),
    .X(_05718_));
 sg13g2_a22oi_1 _12879_ (.Y(_05719_),
    .B1(_05718_),
    .B2(\spiking_network_top_uut.all_data_out[171] ),
    .A2(_05717_),
    .A1(\spiking_network_top_uut.all_data_out[169] ));
 sg13g2_and4_1 _12880_ (.A(\spiking_network_top_uut.all_data_out[169] ),
    .B(\spiking_network_top_uut.all_data_out[171] ),
    .C(_05717_),
    .D(_05718_),
    .X(_05720_));
 sg13g2_nand4_1 _12881_ (.B(\spiking_network_top_uut.all_data_out[171] ),
    .C(_05717_),
    .A(\spiking_network_top_uut.all_data_out[169] ),
    .Y(_05721_),
    .D(_05718_));
 sg13g2_and4_2 _12882_ (.A(\spiking_network_top_uut.all_data_out[168] ),
    .B(\spiking_network_top_uut.all_data_out[170] ),
    .C(_05717_),
    .D(_05718_),
    .X(_05722_));
 sg13g2_nand4_1 _12883_ (.B(\spiking_network_top_uut.all_data_out[170] ),
    .C(_05717_),
    .A(\spiking_network_top_uut.all_data_out[168] ),
    .Y(_05723_),
    .D(_05718_));
 sg13g2_nand3b_1 _12884_ (.B(_05721_),
    .C(_05722_),
    .Y(_05724_),
    .A_N(_05719_));
 sg13g2_a21oi_2 _12885_ (.B1(_05719_),
    .Y(_05725_),
    .A2(_05722_),
    .A1(_05721_));
 sg13g2_mux2_2 _12886_ (.A0(net4593),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[603] ),
    .X(_05726_));
 sg13g2_mux2_2 _12887_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.spike_out ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[607] ),
    .X(_05727_));
 sg13g2_and4_1 _12888_ (.A(\spiking_network_top_uut.all_data_out[173] ),
    .B(\spiking_network_top_uut.all_data_out[175] ),
    .C(_05726_),
    .D(_05727_),
    .X(_05728_));
 sg13g2_nand4_1 _12889_ (.B(\spiking_network_top_uut.all_data_out[175] ),
    .C(_05726_),
    .A(\spiking_network_top_uut.all_data_out[173] ),
    .Y(_05729_),
    .D(_05727_));
 sg13g2_and4_1 _12890_ (.A(\spiking_network_top_uut.all_data_out[172] ),
    .B(\spiking_network_top_uut.all_data_out[174] ),
    .C(_05726_),
    .D(_05727_),
    .X(_05730_));
 sg13g2_a22oi_1 _12891_ (.Y(_05731_),
    .B1(_05727_),
    .B2(\spiking_network_top_uut.all_data_out[175] ),
    .A2(_05726_),
    .A1(\spiking_network_top_uut.all_data_out[173] ));
 sg13g2_or3_2 _12892_ (.A(_05728_),
    .B(_05730_),
    .C(_05731_),
    .X(_05732_));
 sg13g2_o21ai_1 _12893_ (.B1(_05729_),
    .Y(_05733_),
    .A1(_05730_),
    .A2(_05731_));
 sg13g2_nand3b_1 _12894_ (.B(_05725_),
    .C(_05733_),
    .Y(_05734_),
    .A_N(_05716_));
 sg13g2_inv_1 _12895_ (.Y(_05735_),
    .A(_05734_));
 sg13g2_or2_1 _12896_ (.X(_05736_),
    .B(_05734_),
    .A(_05706_));
 sg13g2_inv_2 _12897_ (.Y(_05737_),
    .A(_05736_));
 sg13g2_xnor2_1 _12898_ (.Y(_05738_),
    .A(_05671_),
    .B(_05695_));
 sg13g2_nor2_1 _12899_ (.A(_05725_),
    .B(_05733_),
    .Y(_05739_));
 sg13g2_and2_1 _12900_ (.A(_05716_),
    .B(_05739_),
    .X(_05740_));
 sg13g2_a21oi_2 _12901_ (.B1(_05737_),
    .Y(_05741_),
    .A2(_05740_),
    .A1(_05706_));
 sg13g2_xnor2_1 _12902_ (.Y(_05742_),
    .A(_05738_),
    .B(_05741_));
 sg13g2_o21ai_1 _12903_ (.B1(_05730_),
    .Y(_05743_),
    .A1(_05728_),
    .A2(_05731_));
 sg13g2_o21ai_1 _12904_ (.B1(_05723_),
    .Y(_05744_),
    .A1(_05719_),
    .A2(_05720_));
 sg13g2_o21ai_1 _12905_ (.B1(_05722_),
    .Y(_05745_),
    .A1(_05719_),
    .A2(_05720_));
 sg13g2_nand3b_1 _12906_ (.B(_05721_),
    .C(_05723_),
    .Y(_05746_),
    .A_N(_05719_));
 sg13g2_a22oi_1 _12907_ (.Y(_05747_),
    .B1(_05745_),
    .B2(_05746_),
    .A2(_05743_),
    .A1(_05732_));
 sg13g2_xor2_1 _12908_ (.B(_05715_),
    .A(_05714_),
    .X(_05748_));
 sg13g2_xnor2_1 _12909_ (.Y(_05749_),
    .A(_05714_),
    .B(_05715_));
 sg13g2_and4_1 _12910_ (.A(_05732_),
    .B(_05743_),
    .C(_05745_),
    .D(_05746_),
    .X(_05750_));
 sg13g2_nand4_1 _12911_ (.B(_05743_),
    .C(_05745_),
    .A(_05732_),
    .Y(_05751_),
    .D(_05746_));
 sg13g2_and4_1 _12912_ (.A(_05724_),
    .B(_05732_),
    .C(_05743_),
    .D(_05744_),
    .X(_05752_));
 sg13g2_a22oi_1 _12913_ (.Y(_05753_),
    .B1(_05744_),
    .B2(_05724_),
    .A2(_05743_),
    .A1(_05732_));
 sg13g2_nor3_1 _12914_ (.A(_05747_),
    .B(_05748_),
    .C(_05750_),
    .Y(_05754_));
 sg13g2_o21ai_1 _12915_ (.B1(_05749_),
    .Y(_05755_),
    .A1(_05752_),
    .A2(_05753_));
 sg13g2_a21oi_2 _12916_ (.B1(_05747_),
    .Y(_05756_),
    .A2(_05751_),
    .A1(_05749_));
 sg13g2_xor2_1 _12917_ (.B(_05733_),
    .A(_05725_),
    .X(_05757_));
 sg13g2_xnor2_1 _12918_ (.Y(_05758_),
    .A(_05716_),
    .B(_05757_));
 sg13g2_nand2b_1 _12919_ (.Y(_05759_),
    .B(_05758_),
    .A_N(_05756_));
 sg13g2_xnor2_1 _12920_ (.Y(_05760_),
    .A(_05756_),
    .B(_05758_));
 sg13g2_nand2b_1 _12921_ (.Y(_05761_),
    .B(_05760_),
    .A_N(_05706_));
 sg13g2_nand2_1 _12922_ (.Y(_05762_),
    .A(_05759_),
    .B(_05761_));
 sg13g2_nor2_1 _12923_ (.A(_05735_),
    .B(_05740_),
    .Y(_05763_));
 sg13g2_xnor2_1 _12924_ (.Y(_05764_),
    .A(_05706_),
    .B(_05763_));
 sg13g2_and2_1 _12925_ (.A(_05762_),
    .B(_05764_),
    .X(_05765_));
 sg13g2_xor2_1 _12926_ (.B(_05764_),
    .A(_05762_),
    .X(_05766_));
 sg13g2_xnor2_1 _12927_ (.Y(_05767_),
    .A(_05691_),
    .B(_05693_));
 sg13g2_inv_1 _12928_ (.Y(_05768_),
    .A(_05767_));
 sg13g2_a21oi_1 _12929_ (.A1(_05766_),
    .A2(_05768_),
    .Y(_05769_),
    .B1(_05765_));
 sg13g2_nor2_1 _12930_ (.A(_05742_),
    .B(_05769_),
    .Y(_05770_));
 sg13g2_xnor2_1 _12931_ (.Y(_05771_),
    .A(_05766_),
    .B(_05768_));
 sg13g2_a22oi_1 _12932_ (.Y(_05772_),
    .B1(_05727_),
    .B2(\spiking_network_top_uut.all_data_out[174] ),
    .A2(_05726_),
    .A1(\spiking_network_top_uut.all_data_out[172] ));
 sg13g2_nor2_1 _12933_ (.A(_05730_),
    .B(_05772_),
    .Y(_05773_));
 sg13g2_a22oi_1 _12934_ (.Y(_05774_),
    .B1(_05718_),
    .B2(\spiking_network_top_uut.all_data_out[170] ),
    .A2(_05717_),
    .A1(\spiking_network_top_uut.all_data_out[168] ));
 sg13g2_nor2_1 _12935_ (.A(_05722_),
    .B(_05774_),
    .Y(_05775_));
 sg13g2_and2_1 _12936_ (.A(_05773_),
    .B(_05775_),
    .X(_05776_));
 sg13g2_xor2_1 _12937_ (.B(_05713_),
    .A(_05712_),
    .X(_05777_));
 sg13g2_xor2_1 _12938_ (.B(_05775_),
    .A(_05773_),
    .X(_05778_));
 sg13g2_a21oi_1 _12939_ (.A1(_05777_),
    .A2(_05778_),
    .Y(_05779_),
    .B1(_05776_));
 sg13g2_a21o_1 _12940_ (.A2(_05778_),
    .A1(_05777_),
    .B1(_05776_),
    .X(_05780_));
 sg13g2_nor3_1 _12941_ (.A(_05749_),
    .B(_05752_),
    .C(_05753_),
    .Y(_05781_));
 sg13g2_o21ai_1 _12942_ (.B1(_05748_),
    .Y(_05782_),
    .A1(_05747_),
    .A2(_05750_));
 sg13g2_nor3_2 _12943_ (.A(_05754_),
    .B(_05779_),
    .C(_05781_),
    .Y(_05783_));
 sg13g2_nand3_1 _12944_ (.B(_05780_),
    .C(_05782_),
    .A(_05755_),
    .Y(_05784_));
 sg13g2_xnor2_1 _12945_ (.Y(_05785_),
    .A(_05704_),
    .B(_05705_));
 sg13g2_xnor2_1 _12946_ (.Y(_05786_),
    .A(_05703_),
    .B(_05705_));
 sg13g2_a21oi_2 _12947_ (.B1(_05780_),
    .Y(_05787_),
    .A2(_05782_),
    .A1(_05755_));
 sg13g2_o21ai_1 _12948_ (.B1(_05779_),
    .Y(_05788_),
    .A1(_05754_),
    .A2(_05781_));
 sg13g2_nor3_1 _12949_ (.A(_05783_),
    .B(_05785_),
    .C(_05787_),
    .Y(_05789_));
 sg13g2_nand3_1 _12950_ (.B(_05786_),
    .C(_05788_),
    .A(_05784_),
    .Y(_05790_));
 sg13g2_o21ai_1 _12951_ (.B1(_05784_),
    .Y(_05791_),
    .A1(_05785_),
    .A2(_05787_));
 sg13g2_xnor2_1 _12952_ (.Y(_05792_),
    .A(_05706_),
    .B(_05760_));
 sg13g2_nand2_1 _12953_ (.Y(_05793_),
    .A(_05791_),
    .B(_05792_));
 sg13g2_xnor2_1 _12954_ (.Y(_05794_),
    .A(_05791_),
    .B(_05792_));
 sg13g2_xor2_1 _12955_ (.B(_05689_),
    .A(_05688_),
    .X(_05795_));
 sg13g2_o21ai_1 _12956_ (.B1(_05793_),
    .Y(_05796_),
    .A1(_05794_),
    .A2(_05795_));
 sg13g2_nand2b_1 _12957_ (.Y(_05797_),
    .B(_05796_),
    .A_N(_05771_));
 sg13g2_xor2_1 _12958_ (.B(_05795_),
    .A(_05794_),
    .X(_05798_));
 sg13g2_a22oi_1 _12959_ (.Y(_05799_),
    .B1(_05700_),
    .B2(\spiking_network_top_uut.all_data_out[162] ),
    .A2(_05698_),
    .A1(\spiking_network_top_uut.all_data_out[160] ));
 sg13g2_xnor2_1 _12960_ (.Y(_05800_),
    .A(_05777_),
    .B(_05778_));
 sg13g2_nor3_2 _12961_ (.A(_05704_),
    .B(_05799_),
    .C(_05800_),
    .Y(_05801_));
 sg13g2_a21oi_1 _12962_ (.A1(_05784_),
    .A2(_05788_),
    .Y(_05802_),
    .B1(_05786_));
 sg13g2_o21ai_1 _12963_ (.B1(_05785_),
    .Y(_05803_),
    .A1(_05783_),
    .A2(_05787_));
 sg13g2_nand3_1 _12964_ (.B(_05801_),
    .C(_05803_),
    .A(_05790_),
    .Y(_05804_));
 sg13g2_a21oi_2 _12965_ (.B1(_05801_),
    .Y(_05805_),
    .A2(_05803_),
    .A1(_05790_));
 sg13g2_nor3_1 _12966_ (.A(_05789_),
    .B(_05801_),
    .C(_05802_),
    .Y(_05806_));
 sg13g2_o21ai_1 _12967_ (.B1(_05801_),
    .Y(_05807_),
    .A1(_05789_),
    .A2(_05802_));
 sg13g2_nand2b_2 _12968_ (.Y(_05808_),
    .B(_05807_),
    .A_N(_05806_));
 sg13g2_xnor2_1 _12969_ (.Y(_05809_),
    .A(_05684_),
    .B(_05687_));
 sg13g2_o21ai_1 _12970_ (.B1(_05804_),
    .Y(_05810_),
    .A1(_05805_),
    .A2(_05809_));
 sg13g2_nand2_1 _12971_ (.Y(_05811_),
    .A(_05798_),
    .B(_05810_));
 sg13g2_xnor2_1 _12972_ (.Y(_05812_),
    .A(_05808_),
    .B(_05809_));
 sg13g2_xnor2_1 _12973_ (.Y(_05813_),
    .A(_00046_),
    .B(_05683_));
 sg13g2_o21ai_1 _12974_ (.B1(_05800_),
    .Y(_05814_),
    .A1(_05704_),
    .A2(_05799_));
 sg13g2_nand2b_2 _12975_ (.Y(_05815_),
    .B(_05814_),
    .A_N(_05801_));
 sg13g2_nor2_2 _12976_ (.A(_05813_),
    .B(_05815_),
    .Y(_05816_));
 sg13g2_xor2_1 _12977_ (.B(_05810_),
    .A(_05798_),
    .X(_05817_));
 sg13g2_nand3_1 _12978_ (.B(_05816_),
    .C(_05817_),
    .A(_05812_),
    .Y(_05818_));
 sg13g2_xor2_1 _12979_ (.B(_05796_),
    .A(_05771_),
    .X(_05819_));
 sg13g2_a21o_1 _12980_ (.A2(_05818_),
    .A1(_05811_),
    .B1(_05819_),
    .X(_05820_));
 sg13g2_xnor2_1 _12981_ (.Y(_05821_),
    .A(_05742_),
    .B(_05769_));
 sg13g2_a21oi_1 _12982_ (.A1(_05797_),
    .A2(_05820_),
    .Y(_05822_),
    .B1(_05821_));
 sg13g2_a21oi_1 _12983_ (.A1(_05738_),
    .A2(_05741_),
    .Y(_05823_),
    .B1(_05737_));
 sg13g2_xor2_1 _12984_ (.B(_05741_),
    .A(_05697_),
    .X(_05824_));
 sg13g2_nor2b_1 _12985_ (.A(_05823_),
    .B_N(_05824_),
    .Y(_05825_));
 sg13g2_xnor2_1 _12986_ (.Y(_05826_),
    .A(_05823_),
    .B(_05824_));
 sg13g2_o21ai_1 _12987_ (.B1(_05826_),
    .Y(_05827_),
    .A1(_05770_),
    .A2(_05822_));
 sg13g2_or3_1 _12988_ (.A(_05697_),
    .B(_05737_),
    .C(_05741_),
    .X(_05828_));
 sg13g2_nand3b_1 _12989_ (.B(_05827_),
    .C(_05828_),
    .Y(_05829_),
    .A_N(_05825_));
 sg13g2_nor2_1 _12990_ (.A(_05647_),
    .B(_05697_),
    .Y(_05830_));
 sg13g2_a21oi_1 _12991_ (.A1(_05697_),
    .A2(_05737_),
    .Y(_05831_),
    .B1(_05648_));
 sg13g2_a21oi_2 _12992_ (.B1(_05830_),
    .Y(_05832_),
    .A2(_05831_),
    .A1(_05829_));
 sg13g2_or3_1 _12993_ (.A(_05770_),
    .B(_05822_),
    .C(_05826_),
    .X(_05833_));
 sg13g2_a21oi_1 _12994_ (.A1(_05827_),
    .A2(_05833_),
    .Y(_05834_),
    .B1(_05648_));
 sg13g2_nand3_1 _12995_ (.B(_05820_),
    .C(_05821_),
    .A(_05797_),
    .Y(_05835_));
 sg13g2_nor2_1 _12996_ (.A(_05648_),
    .B(_05822_),
    .Y(_05836_));
 sg13g2_a22oi_1 _12997_ (.Y(_05837_),
    .B1(_05835_),
    .B2(_05836_),
    .A2(_05738_),
    .A1(_05648_));
 sg13g2_or3_1 _12998_ (.A(_05830_),
    .B(_05834_),
    .C(_05837_),
    .X(_05838_));
 sg13g2_a21oi_2 _12999_ (.B1(net3661),
    .Y(_05839_),
    .A2(_05838_),
    .A1(_05832_));
 sg13g2_o21ai_1 _13000_ (.B1(_05837_),
    .Y(_05840_),
    .A1(_05830_),
    .A2(_05834_));
 sg13g2_nor2b_2 _13001_ (.A(_05832_),
    .B_N(_05840_),
    .Y(_05841_));
 sg13g2_nor2_1 _13002_ (.A(_05648_),
    .B(_05815_),
    .Y(_05842_));
 sg13g2_xnor2_1 _13003_ (.Y(_05843_),
    .A(_05813_),
    .B(_05842_));
 sg13g2_nor2_1 _13004_ (.A(_05841_),
    .B(_05843_),
    .Y(_05844_));
 sg13g2_nand2_1 _13005_ (.Y(_05845_),
    .A(net4533),
    .B(_05839_));
 sg13g2_xor2_1 _13006_ (.B(net491),
    .A(net4316),
    .X(_05846_));
 sg13g2_a22oi_1 _13007_ (.Y(_05847_),
    .B1(_00009_),
    .B2(_05846_),
    .A2(net491),
    .A1(net3930));
 sg13g2_o21ai_1 _13008_ (.B1(_05847_),
    .Y(_00563_),
    .A1(_05844_),
    .A2(_05845_));
 sg13g2_a21oi_1 _13009_ (.A1(_05812_),
    .A2(_05816_),
    .Y(_05848_),
    .B1(_05648_));
 sg13g2_o21ai_1 _13010_ (.B1(_05848_),
    .Y(_05849_),
    .A1(_05812_),
    .A2(_05816_));
 sg13g2_o21ai_1 _13011_ (.B1(_05849_),
    .Y(_05850_),
    .A1(_05647_),
    .A2(_05809_));
 sg13g2_o21ai_1 _13012_ (.B1(_05839_),
    .Y(_05851_),
    .A1(_05841_),
    .A2(_05850_));
 sg13g2_xor2_1 _13013_ (.B(_04751_),
    .A(_04750_),
    .X(_05852_));
 sg13g2_a21oi_1 _13014_ (.A1(net3661),
    .A2(_05852_),
    .Y(_05853_),
    .B1(net3930));
 sg13g2_a22oi_1 _13015_ (.Y(_00564_),
    .B1(_05851_),
    .B2(_05853_),
    .A2(_03438_),
    .A1(net3930));
 sg13g2_a21o_1 _13016_ (.A2(_05816_),
    .A1(_05812_),
    .B1(_05817_),
    .X(_05854_));
 sg13g2_nand3_1 _13017_ (.B(_05818_),
    .C(_05854_),
    .A(_05647_),
    .Y(_05855_));
 sg13g2_o21ai_1 _13018_ (.B1(_05855_),
    .Y(_05856_),
    .A1(_05647_),
    .A2(_05795_));
 sg13g2_o21ai_1 _13019_ (.B1(_05839_),
    .Y(_05857_),
    .A1(_05841_),
    .A2(_05856_));
 sg13g2_xnor2_1 _13020_ (.Y(_05858_),
    .A(_04748_),
    .B(_04752_));
 sg13g2_a21oi_1 _13021_ (.A1(net3661),
    .A2(_05858_),
    .Y(_05859_),
    .B1(net3930));
 sg13g2_a22oi_1 _13022_ (.Y(_00565_),
    .B1(_05857_),
    .B2(_05859_),
    .A2(_03437_),
    .A1(net3930));
 sg13g2_nand3_1 _13023_ (.B(_05818_),
    .C(_05819_),
    .A(_05811_),
    .Y(_05860_));
 sg13g2_nand3_1 _13024_ (.B(_05820_),
    .C(_05860_),
    .A(_05647_),
    .Y(_05861_));
 sg13g2_o21ai_1 _13025_ (.B1(_05861_),
    .Y(_05862_),
    .A1(_05647_),
    .A2(_05767_));
 sg13g2_o21ai_1 _13026_ (.B1(_05839_),
    .Y(_05863_),
    .A1(_05841_),
    .A2(_05862_));
 sg13g2_or3_1 _13027_ (.A(_04746_),
    .B(_04747_),
    .C(_04753_),
    .X(_05864_));
 sg13g2_and2_1 _13028_ (.A(_04754_),
    .B(_05864_),
    .X(_05865_));
 sg13g2_a21oi_1 _13029_ (.A1(net3661),
    .A2(_05865_),
    .Y(_05866_),
    .B1(net3930));
 sg13g2_a22oi_1 _13030_ (.Y(_00566_),
    .B1(_05863_),
    .B2(_05866_),
    .A2(_03436_),
    .A1(net3930));
 sg13g2_nor2_1 _13031_ (.A(net4533),
    .B(net449),
    .Y(_05867_));
 sg13g2_a22oi_1 _13032_ (.Y(_05868_),
    .B1(_04757_),
    .B2(_05832_),
    .A2(_04755_),
    .A1(_04745_));
 sg13g2_a21oi_1 _13033_ (.A1(net4533),
    .A2(_05868_),
    .Y(_00567_),
    .B1(_05867_));
 sg13g2_mux4_1 _13034_ (.S0(\spiking_network_top_uut.all_data_out[636] ),
    .A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[0] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[1] ),
    .A2(net3844),
    .A3(net3843),
    .S1(\spiking_network_top_uut.all_data_out[637] ),
    .X(_05869_));
 sg13g2_mux2_1 _13035_ (.A0(net3841),
    .A1(net3900),
    .S(\spiking_network_top_uut.all_data_out[636] ),
    .X(_05870_));
 sg13g2_nor2b_1 _13036_ (.A(\spiking_network_top_uut.all_data_out[636] ),
    .B_N(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[4] ),
    .Y(_05871_));
 sg13g2_a21oi_1 _13037_ (.A1(\spiking_network_top_uut.all_data_out[636] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[5] ),
    .Y(_05872_),
    .B1(_05871_));
 sg13g2_o21ai_1 _13038_ (.B1(\spiking_network_top_uut.all_data_out[638] ),
    .Y(_05873_),
    .A1(\spiking_network_top_uut.all_data_out[637] ),
    .A2(_05872_));
 sg13g2_a21oi_1 _13039_ (.A1(\spiking_network_top_uut.all_data_out[637] ),
    .A2(_05870_),
    .Y(_05874_),
    .B1(_05873_));
 sg13g2_o21ai_1 _13040_ (.B1(net4552),
    .Y(_05875_),
    .A1(\spiking_network_top_uut.all_data_out[638] ),
    .A2(_05869_));
 sg13g2_nand2_1 _13041_ (.Y(_05876_),
    .A(net3934),
    .B(net476));
 sg13g2_o21ai_1 _13042_ (.B1(_05876_),
    .Y(_00568_),
    .A1(_05874_),
    .A2(_05875_));
 sg13g2_mux2_1 _13043_ (.A0(net480),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_reg1 ),
    .S(net4543),
    .X(_00569_));
 sg13g2_nand2_1 _13044_ (.Y(_05877_),
    .A(\spiking_network_top_uut.all_data_out[632] ),
    .B(_03666_));
 sg13g2_nor2_1 _13045_ (.A(\spiking_network_top_uut.all_data_out[632] ),
    .B(net3894),
    .Y(_05878_));
 sg13g2_nor2_1 _13046_ (.A(\spiking_network_top_uut.all_data_out[633] ),
    .B(_05878_),
    .Y(_05879_));
 sg13g2_mux2_1 _13047_ (.A0(net3893),
    .A1(net3892),
    .S(\spiking_network_top_uut.all_data_out[632] ),
    .X(_05880_));
 sg13g2_a221oi_1 _13048_ (.B2(\spiking_network_top_uut.all_data_out[633] ),
    .C1(_03603_),
    .B1(_05880_),
    .A1(_05877_),
    .Y(_05881_),
    .A2(_05879_));
 sg13g2_mux4_1 _13049_ (.S0(\spiking_network_top_uut.all_data_out[632] ),
    .A0(net3898),
    .A1(net3897),
    .A2(net3896),
    .A3(net3895),
    .S1(\spiking_network_top_uut.all_data_out[633] ),
    .X(_05882_));
 sg13g2_o21ai_1 _13050_ (.B1(net4545),
    .Y(_05883_),
    .A1(\spiking_network_top_uut.all_data_out[634] ),
    .A2(_05882_));
 sg13g2_nand2_1 _13051_ (.Y(_05884_),
    .A(net3933),
    .B(net176));
 sg13g2_o21ai_1 _13052_ (.B1(_05884_),
    .Y(_00570_),
    .A1(_05881_),
    .A2(_05883_));
 sg13g2_mux2_1 _13053_ (.A0(net285),
    .A1(net176),
    .S(net4543),
    .X(_00571_));
 sg13g2_nand2_1 _13054_ (.Y(_05885_),
    .A(\spiking_network_top_uut.all_data_out[628] ),
    .B(_03665_));
 sg13g2_nor2_1 _13055_ (.A(\spiking_network_top_uut.all_data_out[628] ),
    .B(net3887),
    .Y(_05886_));
 sg13g2_nor2_1 _13056_ (.A(\spiking_network_top_uut.all_data_out[629] ),
    .B(_05886_),
    .Y(_05887_));
 sg13g2_mux2_1 _13057_ (.A0(net3886),
    .A1(net3885),
    .S(\spiking_network_top_uut.all_data_out[628] ),
    .X(_05888_));
 sg13g2_a221oi_1 _13058_ (.B2(\spiking_network_top_uut.all_data_out[629] ),
    .C1(_03530_),
    .B1(_05888_),
    .A1(_05885_),
    .Y(_05889_),
    .A2(_05887_));
 sg13g2_mux4_1 _13059_ (.S0(\spiking_network_top_uut.all_data_out[628] ),
    .A0(net3891),
    .A1(net3890),
    .A2(net3889),
    .A3(net3888),
    .S1(\spiking_network_top_uut.all_data_out[629] ),
    .X(_05890_));
 sg13g2_o21ai_1 _13060_ (.B1(net4558),
    .Y(_05891_),
    .A1(\spiking_network_top_uut.all_data_out[630] ),
    .A2(_05890_));
 sg13g2_nand2_1 _13061_ (.Y(_05892_),
    .A(net3935),
    .B(net254));
 sg13g2_o21ai_1 _13062_ (.B1(_05892_),
    .Y(_00572_),
    .A1(_05889_),
    .A2(_05891_));
 sg13g2_mux2_1 _13063_ (.A0(net411),
    .A1(net254),
    .S(net4554),
    .X(_00573_));
 sg13g2_mux2_1 _13064_ (.A0(net3882),
    .A1(net3881),
    .S(\spiking_network_top_uut.all_data_out[624] ),
    .X(_05893_));
 sg13g2_nor2b_1 _13065_ (.A(\spiking_network_top_uut.all_data_out[624] ),
    .B_N(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[0] ),
    .Y(_05894_));
 sg13g2_a21oi_1 _13066_ (.A1(\spiking_network_top_uut.all_data_out[624] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[1] ),
    .Y(_05895_),
    .B1(_05894_));
 sg13g2_a21oi_1 _13067_ (.A1(\spiking_network_top_uut.all_data_out[625] ),
    .A2(_05893_),
    .Y(_05896_),
    .B1(\spiking_network_top_uut.all_data_out[626] ));
 sg13g2_o21ai_1 _13068_ (.B1(_05896_),
    .Y(_05897_),
    .A1(\spiking_network_top_uut.all_data_out[625] ),
    .A2(_05895_));
 sg13g2_mux2_1 _13069_ (.A0(net3878),
    .A1(net3877),
    .S(\spiking_network_top_uut.all_data_out[624] ),
    .X(_05898_));
 sg13g2_nor2b_1 _13070_ (.A(\spiking_network_top_uut.all_data_out[624] ),
    .B_N(net3880),
    .Y(_05899_));
 sg13g2_a21oi_1 _13071_ (.A1(\spiking_network_top_uut.all_data_out[624] ),
    .A2(net3879),
    .Y(_05900_),
    .B1(_05899_));
 sg13g2_o21ai_1 _13072_ (.B1(\spiking_network_top_uut.all_data_out[626] ),
    .Y(_05901_),
    .A1(\spiking_network_top_uut.all_data_out[625] ),
    .A2(_05900_));
 sg13g2_a21oi_1 _13073_ (.A1(\spiking_network_top_uut.all_data_out[625] ),
    .A2(_05898_),
    .Y(_05902_),
    .B1(_05901_));
 sg13g2_nand2_1 _13074_ (.Y(_05903_),
    .A(net4555),
    .B(_05897_));
 sg13g2_nand2_1 _13075_ (.Y(_05904_),
    .A(net3938),
    .B(net128));
 sg13g2_o21ai_1 _13076_ (.B1(_05904_),
    .Y(_00574_),
    .A1(_05902_),
    .A2(_05903_));
 sg13g2_mux2_1 _13077_ (.A0(net524),
    .A1(net128),
    .S(net4555),
    .X(_00575_));
 sg13g2_mux4_1 _13078_ (.S0(\spiking_network_top_uut.all_data_out[620] ),
    .A0(net3876),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[1] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[2] ),
    .A3(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[3] ),
    .S1(\spiking_network_top_uut.all_data_out[621] ),
    .X(_05905_));
 sg13g2_mux2_1 _13079_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[6] ),
    .A1(net3869),
    .S(\spiking_network_top_uut.all_data_out[620] ),
    .X(_05906_));
 sg13g2_nor2b_1 _13080_ (.A(\spiking_network_top_uut.all_data_out[620] ),
    .B_N(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[4] ),
    .Y(_05907_));
 sg13g2_a21oi_1 _13081_ (.A1(\spiking_network_top_uut.all_data_out[620] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[5] ),
    .Y(_05908_),
    .B1(_05907_));
 sg13g2_o21ai_1 _13082_ (.B1(\spiking_network_top_uut.all_data_out[622] ),
    .Y(_05909_),
    .A1(\spiking_network_top_uut.all_data_out[621] ),
    .A2(_05908_));
 sg13g2_a21oi_1 _13083_ (.A1(\spiking_network_top_uut.all_data_out[621] ),
    .A2(_05906_),
    .Y(_05910_),
    .B1(_05909_));
 sg13g2_o21ai_1 _13084_ (.B1(net4569),
    .Y(_05911_),
    .A1(\spiking_network_top_uut.all_data_out[622] ),
    .A2(_05905_));
 sg13g2_nand2_1 _13085_ (.Y(_05912_),
    .A(net3939),
    .B(net168));
 sg13g2_o21ai_1 _13086_ (.B1(_05912_),
    .Y(_00576_),
    .A1(_05910_),
    .A2(_05911_));
 sg13g2_mux2_1 _13087_ (.A0(net300),
    .A1(net168),
    .S(net4569),
    .X(_00577_));
 sg13g2_mux4_1 _13088_ (.S0(\spiking_network_top_uut.all_data_out[616] ),
    .A0(net3868),
    .A1(net3867),
    .A2(net3866),
    .A3(net3865),
    .S1(\spiking_network_top_uut.all_data_out[617] ),
    .X(_05913_));
 sg13g2_mux2_1 _13089_ (.A0(net3862),
    .A1(net3861),
    .S(\spiking_network_top_uut.all_data_out[616] ),
    .X(_05914_));
 sg13g2_nor2b_1 _13090_ (.A(\spiking_network_top_uut.all_data_out[616] ),
    .B_N(net3864),
    .Y(_05915_));
 sg13g2_a21oi_1 _13091_ (.A1(\spiking_network_top_uut.all_data_out[616] ),
    .A2(net3863),
    .Y(_05916_),
    .B1(_05915_));
 sg13g2_o21ai_1 _13092_ (.B1(\spiking_network_top_uut.all_data_out[618] ),
    .Y(_05917_),
    .A1(\spiking_network_top_uut.all_data_out[617] ),
    .A2(_05916_));
 sg13g2_a21oi_1 _13093_ (.A1(\spiking_network_top_uut.all_data_out[617] ),
    .A2(_05914_),
    .Y(_05918_),
    .B1(_05917_));
 sg13g2_o21ai_1 _13094_ (.B1(net4562),
    .Y(_05919_),
    .A1(\spiking_network_top_uut.all_data_out[618] ),
    .A2(_05913_));
 sg13g2_nand2_1 _13095_ (.Y(_05920_),
    .A(net3936),
    .B(net64));
 sg13g2_o21ai_1 _13096_ (.B1(_05920_),
    .Y(_00578_),
    .A1(_05918_),
    .A2(_05919_));
 sg13g2_mux2_1 _13097_ (.A0(net268),
    .A1(net64),
    .S(net4562),
    .X(_00579_));
 sg13g2_nand2_1 _13098_ (.Y(_05921_),
    .A(\spiking_network_top_uut.all_data_out[612] ),
    .B(_03664_));
 sg13g2_nor2_1 _13099_ (.A(\spiking_network_top_uut.all_data_out[612] ),
    .B(net3856),
    .Y(_05922_));
 sg13g2_nor2_1 _13100_ (.A(\spiking_network_top_uut.all_data_out[613] ),
    .B(_05922_),
    .Y(_05923_));
 sg13g2_mux2_1 _13101_ (.A0(net3855),
    .A1(net3854),
    .S(\spiking_network_top_uut.all_data_out[612] ),
    .X(_05924_));
 sg13g2_a221oi_1 _13102_ (.B2(\spiking_network_top_uut.all_data_out[613] ),
    .C1(_03531_),
    .B1(_05924_),
    .A1(_05921_),
    .Y(_05925_),
    .A2(_05923_));
 sg13g2_mux4_1 _13103_ (.S0(\spiking_network_top_uut.all_data_out[612] ),
    .A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[0] ),
    .A1(net3859),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[2] ),
    .A3(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[3] ),
    .S1(\spiking_network_top_uut.all_data_out[613] ),
    .X(_05926_));
 sg13g2_o21ai_1 _13104_ (.B1(net4540),
    .Y(_05927_),
    .A1(\spiking_network_top_uut.all_data_out[614] ),
    .A2(_05926_));
 sg13g2_nand2_1 _13105_ (.Y(_05928_),
    .A(net3932),
    .B(net61));
 sg13g2_o21ai_1 _13106_ (.B1(_05928_),
    .Y(_00580_),
    .A1(_05925_),
    .A2(_05927_));
 sg13g2_mux2_1 _13107_ (.A0(net124),
    .A1(net61),
    .S(net4541),
    .X(_00581_));
 sg13g2_mux4_1 _13108_ (.S0(\spiking_network_top_uut.all_data_out[608] ),
    .A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[0] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[1] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[2] ),
    .A3(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[3] ),
    .S1(\spiking_network_top_uut.all_data_out[609] ),
    .X(_05929_));
 sg13g2_mux2_1 _13109_ (.A0(net3848),
    .A1(net3847),
    .S(\spiking_network_top_uut.all_data_out[608] ),
    .X(_05930_));
 sg13g2_nor2b_1 _13110_ (.A(\spiking_network_top_uut.all_data_out[608] ),
    .B_N(net3849),
    .Y(_05931_));
 sg13g2_a21oi_1 _13111_ (.A1(\spiking_network_top_uut.all_data_out[608] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[5] ),
    .Y(_05932_),
    .B1(_05931_));
 sg13g2_o21ai_1 _13112_ (.B1(\spiking_network_top_uut.all_data_out[610] ),
    .Y(_05933_),
    .A1(\spiking_network_top_uut.all_data_out[609] ),
    .A2(_05932_));
 sg13g2_a21oi_1 _13113_ (.A1(\spiking_network_top_uut.all_data_out[609] ),
    .A2(_05930_),
    .Y(_05934_),
    .B1(_05933_));
 sg13g2_o21ai_1 _13114_ (.B1(net4544),
    .Y(_05935_),
    .A1(\spiking_network_top_uut.all_data_out[610] ),
    .A2(_05929_));
 sg13g2_nand2_1 _13115_ (.Y(_05936_),
    .A(net3933),
    .B(net150));
 sg13g2_o21ai_1 _13116_ (.B1(_05936_),
    .Y(_00582_),
    .A1(_05934_),
    .A2(_05935_));
 sg13g2_nor3_2 _13117_ (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[2] ),
    .B(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[0] ),
    .C(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[1] ),
    .Y(_05937_));
 sg13g2_nor2b_2 _13118_ (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[3] ),
    .B_N(_05937_),
    .Y(_05938_));
 sg13g2_nor2b_2 _13119_ (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[4] ),
    .B_N(_05938_),
    .Y(_05939_));
 sg13g2_nand2b_2 _13120_ (.Y(_05940_),
    .B(_05938_),
    .A_N(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[4] ));
 sg13g2_o21ai_1 _13121_ (.B1(net4529),
    .Y(_05941_),
    .A1(net3666),
    .A2(_05940_));
 sg13g2_nor2b_1 _13122_ (.A(net3665),
    .B_N(net331),
    .Y(_05942_));
 sg13g2_a21oi_1 _13123_ (.A1(net4283),
    .A2(net3665),
    .Y(_05943_),
    .B1(_05942_));
 sg13g2_nand2_1 _13124_ (.Y(_05944_),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[0] ),
    .B(_05941_));
 sg13g2_o21ai_1 _13125_ (.B1(_05944_),
    .Y(_00583_),
    .A1(_05941_),
    .A2(_05943_));
 sg13g2_xor2_1 _13126_ (.B(net370),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[0] ),
    .X(_05945_));
 sg13g2_nor2_1 _13127_ (.A(net3665),
    .B(_05945_),
    .Y(_05946_));
 sg13g2_a21oi_1 _13128_ (.A1(net4280),
    .A2(net3665),
    .Y(_05947_),
    .B1(_05946_));
 sg13g2_nand2_1 _13129_ (.Y(_05948_),
    .A(net370),
    .B(_05941_));
 sg13g2_o21ai_1 _13130_ (.B1(_05948_),
    .Y(_00584_),
    .A1(_05941_),
    .A2(_05947_));
 sg13g2_nand2_1 _13131_ (.Y(_05949_),
    .A(net4276),
    .B(net3665));
 sg13g2_o21ai_1 _13132_ (.B1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[2] ),
    .Y(_05950_),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[0] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[1] ));
 sg13g2_nor2b_1 _13133_ (.A(_05937_),
    .B_N(_05950_),
    .Y(_05951_));
 sg13g2_o21ai_1 _13134_ (.B1(_05949_),
    .Y(_05952_),
    .A1(net3665),
    .A2(_05951_));
 sg13g2_mux2_1 _13135_ (.A0(_05952_),
    .A1(net401),
    .S(_05941_),
    .X(_00585_));
 sg13g2_nand2_1 _13136_ (.Y(_05953_),
    .A(net4273),
    .B(net3665));
 sg13g2_xnor2_1 _13137_ (.Y(_05954_),
    .A(net438),
    .B(_05937_));
 sg13g2_o21ai_1 _13138_ (.B1(_05953_),
    .Y(_05955_),
    .A1(net3665),
    .A2(_05954_));
 sg13g2_mux2_1 _13139_ (.A0(_05955_),
    .A1(net438),
    .S(_05941_),
    .X(_00586_));
 sg13g2_nand2_1 _13140_ (.Y(_05956_),
    .A(net3922),
    .B(net298));
 sg13g2_nor2_1 _13141_ (.A(net4269),
    .B(_04772_),
    .Y(_05957_));
 sg13g2_nor2b_1 _13142_ (.A(_05938_),
    .B_N(net298),
    .Y(_05958_));
 sg13g2_o21ai_1 _13143_ (.B1(net4529),
    .Y(_05959_),
    .A1(net3666),
    .A2(_05958_));
 sg13g2_o21ai_1 _13144_ (.B1(_05956_),
    .Y(_00587_),
    .A1(_05957_),
    .A2(_05959_));
 sg13g2_mux2_1 _13145_ (.A0(net335),
    .A1(net150),
    .S(net4538),
    .X(_00588_));
 sg13g2_nor2_1 _13146_ (.A(_00049_),
    .B(net3740),
    .Y(_05960_));
 sg13g2_nor2_2 _13147_ (.A(net3743),
    .B(_05960_),
    .Y(_05961_));
 sg13g2_nor2_1 _13148_ (.A(_00049_),
    .B(_05961_),
    .Y(_05962_));
 sg13g2_nand2b_1 _13149_ (.Y(_05963_),
    .B(_05961_),
    .A_N(_00049_));
 sg13g2_o21ai_1 _13150_ (.B1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ),
    .Y(_05964_),
    .A1(_00049_),
    .A2(_05961_));
 sg13g2_inv_1 _13151_ (.Y(_05965_),
    .A(_05964_));
 sg13g2_a21o_1 _13152_ (.A2(net3746),
    .A1(_00050_),
    .B1(_05961_),
    .X(_05966_));
 sg13g2_and2_1 _13153_ (.A(_00051_),
    .B(net3746),
    .X(_05967_));
 sg13g2_o21ai_1 _13154_ (.B1(net3917),
    .Y(_05968_),
    .A1(_00050_),
    .A2(net3905));
 sg13g2_a21oi_1 _13155_ (.A1(net3905),
    .A2(_05960_),
    .Y(_05969_),
    .B1(_05968_));
 sg13g2_o21ai_1 _13156_ (.B1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ),
    .Y(_05970_),
    .A1(_05967_),
    .A2(_05969_));
 sg13g2_o21ai_1 _13157_ (.B1(net3914),
    .Y(_05971_),
    .A1(_00049_),
    .A2(net3912));
 sg13g2_a221oi_1 _13158_ (.B2(_00050_),
    .C1(net3746),
    .B1(net3901),
    .A1(_00051_),
    .Y(_05972_),
    .A2(net3739));
 sg13g2_a22oi_1 _13159_ (.Y(_05973_),
    .B1(_05971_),
    .B2(_05972_),
    .A2(net3746),
    .A1(_03481_));
 sg13g2_nor2b_1 _13160_ (.A(_05973_),
    .B_N(_00052_),
    .Y(_05974_));
 sg13g2_nor3_1 _13161_ (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ),
    .B(_05967_),
    .C(_05969_),
    .Y(_05975_));
 sg13g2_or3_1 _13162_ (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ),
    .B(_05967_),
    .C(_05969_),
    .X(_05976_));
 sg13g2_nand2_1 _13163_ (.Y(_05977_),
    .A(_05970_),
    .B(_05976_));
 sg13g2_o21ai_1 _13164_ (.B1(_05970_),
    .Y(_05978_),
    .A1(_05974_),
    .A2(_05975_));
 sg13g2_xor2_1 _13165_ (.B(_05966_),
    .A(_00051_),
    .X(_05979_));
 sg13g2_nor2b_1 _13166_ (.A(_05979_),
    .B_N(_05978_),
    .Y(_05980_));
 sg13g2_a21o_1 _13167_ (.A2(_05966_),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ),
    .B1(_05980_),
    .X(_05981_));
 sg13g2_xnor2_1 _13168_ (.Y(_05982_),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ),
    .B(_05962_));
 sg13g2_a21oi_1 _13169_ (.A1(_05981_),
    .A2(_05982_),
    .Y(_05983_),
    .B1(_05965_));
 sg13g2_a22oi_1 _13170_ (.Y(_05984_),
    .B1(_05963_),
    .B2(_05983_),
    .A2(_05961_),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ));
 sg13g2_a21oi_2 _13171_ (.B1(_05984_),
    .Y(_05985_),
    .A2(_00049_),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ));
 sg13g2_mux2_1 _13172_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.spike_out ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[611] ),
    .X(_05986_));
 sg13g2_nand2_1 _13173_ (.Y(_05987_),
    .A(\spiking_network_top_uut.all_data_out[177] ),
    .B(_05986_));
 sg13g2_mux2_2 _13174_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.spike_out ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[615] ),
    .X(_05988_));
 sg13g2_nand2_1 _13175_ (.Y(_05989_),
    .A(\spiking_network_top_uut.all_data_out[179] ),
    .B(_05988_));
 sg13g2_nor2_1 _13176_ (.A(_05987_),
    .B(_05989_),
    .Y(_05990_));
 sg13g2_nand4_1 _13177_ (.B(\spiking_network_top_uut.all_data_out[178] ),
    .C(_05986_),
    .A(\spiking_network_top_uut.all_data_out[176] ),
    .Y(_05991_),
    .D(_05988_));
 sg13g2_inv_1 _13178_ (.Y(_05992_),
    .A(_05991_));
 sg13g2_xor2_1 _13179_ (.B(_05989_),
    .A(_05987_),
    .X(_05993_));
 sg13g2_a21oi_2 _13180_ (.B1(_05990_),
    .Y(_05994_),
    .A2(_05993_),
    .A1(_05991_));
 sg13g2_mux2_2 _13181_ (.A0(net4597),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[619] ),
    .X(_05995_));
 sg13g2_nand2_1 _13182_ (.Y(_05996_),
    .A(\spiking_network_top_uut.all_data_out[181] ),
    .B(_05995_));
 sg13g2_mux2_2 _13183_ (.A0(net4596),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[623] ),
    .X(_05997_));
 sg13g2_nand2_1 _13184_ (.Y(_05998_),
    .A(\spiking_network_top_uut.all_data_out[183] ),
    .B(_05997_));
 sg13g2_nor2_1 _13185_ (.A(_05996_),
    .B(_05998_),
    .Y(_05999_));
 sg13g2_nand2_1 _13186_ (.Y(_06000_),
    .A(\spiking_network_top_uut.all_data_out[180] ),
    .B(_05995_));
 sg13g2_nand2_1 _13187_ (.Y(_06001_),
    .A(\spiking_network_top_uut.all_data_out[182] ),
    .B(_05997_));
 sg13g2_or2_1 _13188_ (.X(_06002_),
    .B(_06001_),
    .A(_06000_));
 sg13g2_xor2_1 _13189_ (.B(_05998_),
    .A(_05996_),
    .X(_06003_));
 sg13g2_a21oi_2 _13190_ (.B1(_05999_),
    .Y(_06004_),
    .A2(_06003_),
    .A1(_06002_));
 sg13g2_mux2_2 _13191_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.spike_out ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[627] ),
    .X(_06005_));
 sg13g2_mux2_2 _13192_ (.A0(net4594),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[631] ),
    .X(_06006_));
 sg13g2_a22oi_1 _13193_ (.Y(_06007_),
    .B1(_06006_),
    .B2(\spiking_network_top_uut.all_data_out[187] ),
    .A2(_06005_),
    .A1(\spiking_network_top_uut.all_data_out[185] ));
 sg13g2_and4_1 _13194_ (.A(\spiking_network_top_uut.all_data_out[185] ),
    .B(\spiking_network_top_uut.all_data_out[187] ),
    .C(_06005_),
    .D(_06006_),
    .X(_06008_));
 sg13g2_nand4_1 _13195_ (.B(\spiking_network_top_uut.all_data_out[187] ),
    .C(_06005_),
    .A(\spiking_network_top_uut.all_data_out[185] ),
    .Y(_06009_),
    .D(_06006_));
 sg13g2_and4_2 _13196_ (.A(\spiking_network_top_uut.all_data_out[184] ),
    .B(\spiking_network_top_uut.all_data_out[186] ),
    .C(_06005_),
    .D(_06006_),
    .X(_06010_));
 sg13g2_nand4_1 _13197_ (.B(\spiking_network_top_uut.all_data_out[186] ),
    .C(_06005_),
    .A(\spiking_network_top_uut.all_data_out[184] ),
    .Y(_06011_),
    .D(_06006_));
 sg13g2_nand3b_1 _13198_ (.B(_06009_),
    .C(_06010_),
    .Y(_06012_),
    .A_N(_06007_));
 sg13g2_a21oi_2 _13199_ (.B1(_06007_),
    .Y(_06013_),
    .A2(_06010_),
    .A1(_06009_));
 sg13g2_mux2_1 _13200_ (.A0(net4593),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[635] ),
    .X(_06014_));
 sg13g2_mux2_2 _13201_ (.A0(net4592),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[639] ),
    .X(_06015_));
 sg13g2_and4_1 _13202_ (.A(\spiking_network_top_uut.all_data_out[189] ),
    .B(\spiking_network_top_uut.all_data_out[191] ),
    .C(_06014_),
    .D(_06015_),
    .X(_06016_));
 sg13g2_nand4_1 _13203_ (.B(\spiking_network_top_uut.all_data_out[191] ),
    .C(_06014_),
    .A(\spiking_network_top_uut.all_data_out[189] ),
    .Y(_06017_),
    .D(_06015_));
 sg13g2_and4_2 _13204_ (.A(\spiking_network_top_uut.all_data_out[188] ),
    .B(\spiking_network_top_uut.all_data_out[190] ),
    .C(_06014_),
    .D(_06015_),
    .X(_06018_));
 sg13g2_a22oi_1 _13205_ (.Y(_06019_),
    .B1(_06015_),
    .B2(\spiking_network_top_uut.all_data_out[191] ),
    .A2(_06014_),
    .A1(\spiking_network_top_uut.all_data_out[189] ));
 sg13g2_or3_2 _13206_ (.A(_06016_),
    .B(_06018_),
    .C(_06019_),
    .X(_06020_));
 sg13g2_o21ai_1 _13207_ (.B1(_06017_),
    .Y(_06021_),
    .A1(_06018_),
    .A2(_06019_));
 sg13g2_nand3b_1 _13208_ (.B(_06013_),
    .C(_06021_),
    .Y(_06022_),
    .A_N(_06004_));
 sg13g2_or2_1 _13209_ (.X(_06023_),
    .B(_06022_),
    .A(_05994_));
 sg13g2_inv_1 _13210_ (.Y(_06024_),
    .A(_06023_));
 sg13g2_nor2_1 _13211_ (.A(_06013_),
    .B(_06021_),
    .Y(_06025_));
 sg13g2_nand2_1 _13212_ (.Y(_06026_),
    .A(_06004_),
    .B(_06025_));
 sg13g2_mux2_2 _13213_ (.A0(_06022_),
    .A1(_06026_),
    .S(_05994_),
    .X(_06027_));
 sg13g2_xor2_1 _13214_ (.B(_05983_),
    .A(_05963_),
    .X(_06028_));
 sg13g2_nor2b_1 _13215_ (.A(_06028_),
    .B_N(_06027_),
    .Y(_06029_));
 sg13g2_xnor2_1 _13216_ (.Y(_06030_),
    .A(_06027_),
    .B(_06028_));
 sg13g2_o21ai_1 _13217_ (.B1(_06018_),
    .Y(_06031_),
    .A1(_06016_),
    .A2(_06019_));
 sg13g2_o21ai_1 _13218_ (.B1(_06011_),
    .Y(_06032_),
    .A1(_06007_),
    .A2(_06008_));
 sg13g2_o21ai_1 _13219_ (.B1(_06010_),
    .Y(_06033_),
    .A1(_06007_),
    .A2(_06008_));
 sg13g2_nand3b_1 _13220_ (.B(_06009_),
    .C(_06011_),
    .Y(_06034_),
    .A_N(_06007_));
 sg13g2_a22oi_1 _13221_ (.Y(_06035_),
    .B1(_06033_),
    .B2(_06034_),
    .A2(_06031_),
    .A1(_06020_));
 sg13g2_xor2_1 _13222_ (.B(_06003_),
    .A(_06002_),
    .X(_06036_));
 sg13g2_xnor2_1 _13223_ (.Y(_06037_),
    .A(_06002_),
    .B(_06003_));
 sg13g2_and4_1 _13224_ (.A(_06020_),
    .B(_06031_),
    .C(_06033_),
    .D(_06034_),
    .X(_06038_));
 sg13g2_nand4_1 _13225_ (.B(_06031_),
    .C(_06033_),
    .A(_06020_),
    .Y(_06039_),
    .D(_06034_));
 sg13g2_and4_1 _13226_ (.A(_06012_),
    .B(_06020_),
    .C(_06031_),
    .D(_06032_),
    .X(_06040_));
 sg13g2_a22oi_1 _13227_ (.Y(_06041_),
    .B1(_06032_),
    .B2(_06012_),
    .A2(_06031_),
    .A1(_06020_));
 sg13g2_nor3_2 _13228_ (.A(_06035_),
    .B(_06036_),
    .C(_06038_),
    .Y(_06042_));
 sg13g2_a21oi_2 _13229_ (.B1(_06035_),
    .Y(_06043_),
    .A2(_06039_),
    .A1(_06037_));
 sg13g2_xor2_1 _13230_ (.B(_06021_),
    .A(_06013_),
    .X(_06044_));
 sg13g2_xnor2_1 _13231_ (.Y(_06045_),
    .A(_06004_),
    .B(_06044_));
 sg13g2_nand2b_1 _13232_ (.Y(_06046_),
    .B(_06045_),
    .A_N(_06043_));
 sg13g2_xnor2_1 _13233_ (.Y(_06047_),
    .A(_06043_),
    .B(_06045_));
 sg13g2_nand2b_1 _13234_ (.Y(_06048_),
    .B(_06047_),
    .A_N(_05994_));
 sg13g2_nand2_1 _13235_ (.Y(_06049_),
    .A(_06046_),
    .B(_06048_));
 sg13g2_nand2_1 _13236_ (.Y(_06050_),
    .A(_06022_),
    .B(_06026_));
 sg13g2_xor2_1 _13237_ (.B(_06050_),
    .A(_05994_),
    .X(_06051_));
 sg13g2_and2_1 _13238_ (.A(_06049_),
    .B(_06051_),
    .X(_06052_));
 sg13g2_xor2_1 _13239_ (.B(_06051_),
    .A(_06049_),
    .X(_06053_));
 sg13g2_xnor2_1 _13240_ (.Y(_06054_),
    .A(_05981_),
    .B(_05982_));
 sg13g2_inv_1 _13241_ (.Y(_06055_),
    .A(_06054_));
 sg13g2_a21oi_1 _13242_ (.A1(_06053_),
    .A2(_06055_),
    .Y(_06056_),
    .B1(_06052_));
 sg13g2_nor2b_1 _13243_ (.A(_06056_),
    .B_N(_06030_),
    .Y(_06057_));
 sg13g2_xor2_1 _13244_ (.B(_06054_),
    .A(_06053_),
    .X(_06058_));
 sg13g2_a22oi_1 _13245_ (.Y(_06059_),
    .B1(_06015_),
    .B2(\spiking_network_top_uut.all_data_out[190] ),
    .A2(_06014_),
    .A1(\spiking_network_top_uut.all_data_out[188] ));
 sg13g2_nor2_2 _13246_ (.A(_06018_),
    .B(_06059_),
    .Y(_06060_));
 sg13g2_a22oi_1 _13247_ (.Y(_06061_),
    .B1(_06006_),
    .B2(\spiking_network_top_uut.all_data_out[186] ),
    .A2(_06005_),
    .A1(\spiking_network_top_uut.all_data_out[184] ));
 sg13g2_nor2_1 _13248_ (.A(_06010_),
    .B(_06061_),
    .Y(_06062_));
 sg13g2_and2_1 _13249_ (.A(_06060_),
    .B(_06062_),
    .X(_06063_));
 sg13g2_xor2_1 _13250_ (.B(_06001_),
    .A(_06000_),
    .X(_06064_));
 sg13g2_xor2_1 _13251_ (.B(_06062_),
    .A(_06060_),
    .X(_06065_));
 sg13g2_a21oi_2 _13252_ (.B1(_06063_),
    .Y(_06066_),
    .A2(_06065_),
    .A1(_06064_));
 sg13g2_nor3_2 _13253_ (.A(_06037_),
    .B(_06040_),
    .C(_06041_),
    .Y(_06067_));
 sg13g2_nor3_1 _13254_ (.A(_06042_),
    .B(_06066_),
    .C(_06067_),
    .Y(_06068_));
 sg13g2_or3_1 _13255_ (.A(_06042_),
    .B(_06066_),
    .C(_06067_),
    .X(_06069_));
 sg13g2_xnor2_1 _13256_ (.Y(_06070_),
    .A(_05991_),
    .B(_05993_));
 sg13g2_o21ai_1 _13257_ (.B1(_06066_),
    .Y(_06071_),
    .A1(_06042_),
    .A2(_06067_));
 sg13g2_nand3_1 _13258_ (.B(_06070_),
    .C(_06071_),
    .A(_06069_),
    .Y(_06072_));
 sg13g2_a21o_2 _13259_ (.A2(_06071_),
    .A1(_06070_),
    .B1(_06068_),
    .X(_06073_));
 sg13g2_xnor2_1 _13260_ (.Y(_06074_),
    .A(_05994_),
    .B(_06047_));
 sg13g2_nand2_1 _13261_ (.Y(_06075_),
    .A(_06073_),
    .B(_06074_));
 sg13g2_xnor2_1 _13262_ (.Y(_06076_),
    .A(_06073_),
    .B(_06074_));
 sg13g2_xor2_1 _13263_ (.B(_05979_),
    .A(_05978_),
    .X(_06077_));
 sg13g2_o21ai_1 _13264_ (.B1(_06075_),
    .Y(_06078_),
    .A1(_06076_),
    .A2(_06077_));
 sg13g2_nand2b_1 _13265_ (.Y(_06079_),
    .B(_06078_),
    .A_N(_06058_));
 sg13g2_xor2_1 _13266_ (.B(_06077_),
    .A(_06076_),
    .X(_06080_));
 sg13g2_a22oi_1 _13267_ (.Y(_06081_),
    .B1(_05988_),
    .B2(\spiking_network_top_uut.all_data_out[178] ),
    .A2(_05986_),
    .A1(\spiking_network_top_uut.all_data_out[176] ));
 sg13g2_nor2_2 _13268_ (.A(_05992_),
    .B(_06081_),
    .Y(_06082_));
 sg13g2_inv_1 _13269_ (.Y(_06083_),
    .A(_06082_));
 sg13g2_xnor2_1 _13270_ (.Y(_06084_),
    .A(_06064_),
    .B(_06065_));
 sg13g2_nor2_1 _13271_ (.A(_06083_),
    .B(_06084_),
    .Y(_06085_));
 sg13g2_a21o_2 _13272_ (.A2(_06071_),
    .A1(_06069_),
    .B1(_06070_),
    .X(_06086_));
 sg13g2_and3_1 _13273_ (.X(_06087_),
    .A(_06072_),
    .B(_06085_),
    .C(_06086_));
 sg13g2_nand3_1 _13274_ (.B(_06085_),
    .C(_06086_),
    .A(_06072_),
    .Y(_06088_));
 sg13g2_a21oi_1 _13275_ (.A1(_06072_),
    .A2(_06086_),
    .Y(_06089_),
    .B1(_06085_));
 sg13g2_xnor2_1 _13276_ (.Y(_06090_),
    .A(_05974_),
    .B(_05977_));
 sg13g2_nor3_1 _13277_ (.A(_06087_),
    .B(_06089_),
    .C(_06090_),
    .Y(_06091_));
 sg13g2_o21ai_1 _13278_ (.B1(_06088_),
    .Y(_06092_),
    .A1(_06089_),
    .A2(_06090_));
 sg13g2_nand2_1 _13279_ (.Y(_06093_),
    .A(_06080_),
    .B(_06092_));
 sg13g2_o21ai_1 _13280_ (.B1(_06090_),
    .Y(_06094_),
    .A1(_06087_),
    .A2(_06089_));
 sg13g2_nor2b_1 _13281_ (.A(_06091_),
    .B_N(_06094_),
    .Y(_06095_));
 sg13g2_xnor2_1 _13282_ (.Y(_06096_),
    .A(_00052_),
    .B(_05973_));
 sg13g2_xnor2_1 _13283_ (.Y(_06097_),
    .A(_06083_),
    .B(_06084_));
 sg13g2_nor2_1 _13284_ (.A(_06096_),
    .B(_06097_),
    .Y(_06098_));
 sg13g2_xor2_1 _13285_ (.B(_06092_),
    .A(_06080_),
    .X(_06099_));
 sg13g2_nand3_1 _13286_ (.B(_06098_),
    .C(_06099_),
    .A(_06095_),
    .Y(_06100_));
 sg13g2_xor2_1 _13287_ (.B(_06078_),
    .A(_06058_),
    .X(_06101_));
 sg13g2_a21o_1 _13288_ (.A2(_06100_),
    .A1(_06093_),
    .B1(_06101_),
    .X(_06102_));
 sg13g2_xor2_1 _13289_ (.B(_06056_),
    .A(_06030_),
    .X(_06103_));
 sg13g2_a21oi_1 _13290_ (.A1(_06079_),
    .A2(_06102_),
    .Y(_06104_),
    .B1(_06103_));
 sg13g2_nor2_1 _13291_ (.A(_06024_),
    .B(_06029_),
    .Y(_06105_));
 sg13g2_xor2_1 _13292_ (.B(_06027_),
    .A(_05985_),
    .X(_06106_));
 sg13g2_nand2b_1 _13293_ (.Y(_06107_),
    .B(_06106_),
    .A_N(_06105_));
 sg13g2_xnor2_1 _13294_ (.Y(_06108_),
    .A(_06105_),
    .B(_06106_));
 sg13g2_or3_1 _13295_ (.A(_06057_),
    .B(_06104_),
    .C(_06108_),
    .X(_06109_));
 sg13g2_o21ai_1 _13296_ (.B1(_06108_),
    .Y(_06110_),
    .A1(_06057_),
    .A2(_06104_));
 sg13g2_or2_1 _13297_ (.X(_06111_),
    .B(_05985_),
    .A(_05939_));
 sg13g2_a21o_1 _13298_ (.A2(_06110_),
    .A1(_06109_),
    .B1(_05940_),
    .X(_06112_));
 sg13g2_nand3_1 _13299_ (.B(_06102_),
    .C(_06103_),
    .A(_06079_),
    .Y(_06113_));
 sg13g2_nand3b_1 _13300_ (.B(_06113_),
    .C(_05939_),
    .Y(_06114_),
    .A_N(_06104_));
 sg13g2_o21ai_1 _13301_ (.B1(_06114_),
    .Y(_06115_),
    .A1(_05939_),
    .A2(_06028_));
 sg13g2_nand3_1 _13302_ (.B(_06112_),
    .C(_06115_),
    .A(_06111_),
    .Y(_06116_));
 sg13g2_o21ai_1 _13303_ (.B1(_05985_),
    .Y(_06117_),
    .A1(_05940_),
    .A2(_06024_));
 sg13g2_or3_1 _13304_ (.A(_05985_),
    .B(_06024_),
    .C(_06027_),
    .X(_06118_));
 sg13g2_nand3_1 _13305_ (.B(_06110_),
    .C(_06118_),
    .A(_06107_),
    .Y(_06119_));
 sg13g2_o21ai_1 _13306_ (.B1(_06117_),
    .Y(_06120_),
    .A1(_05940_),
    .A2(_06119_));
 sg13g2_a21oi_2 _13307_ (.B1(net3666),
    .Y(_06121_),
    .A2(_06120_),
    .A1(_06116_));
 sg13g2_nand2_1 _13308_ (.Y(_06122_),
    .A(net4530),
    .B(_06121_));
 sg13g2_a21oi_1 _13309_ (.A1(_06111_),
    .A2(_06112_),
    .Y(_06123_),
    .B1(_06115_));
 sg13g2_nor2_2 _13310_ (.A(_06120_),
    .B(_06123_),
    .Y(_06124_));
 sg13g2_nor2_1 _13311_ (.A(_05940_),
    .B(_06097_),
    .Y(_06125_));
 sg13g2_xnor2_1 _13312_ (.Y(_06126_),
    .A(_06096_),
    .B(_06125_));
 sg13g2_nor2_1 _13313_ (.A(_06124_),
    .B(_06126_),
    .Y(_06127_));
 sg13g2_xor2_1 _13314_ (.B(net475),
    .A(net4311),
    .X(_06128_));
 sg13g2_a22oi_1 _13315_ (.Y(_06129_),
    .B1(_00010_),
    .B2(_06128_),
    .A2(net475),
    .A1(net3927));
 sg13g2_o21ai_1 _13316_ (.B1(_06129_),
    .Y(_00589_),
    .A1(_06122_),
    .A2(_06127_));
 sg13g2_xor2_1 _13317_ (.B(_06098_),
    .A(_06095_),
    .X(_06130_));
 sg13g2_nand2_1 _13318_ (.Y(_06131_),
    .A(_05939_),
    .B(_06130_));
 sg13g2_o21ai_1 _13319_ (.B1(_06131_),
    .Y(_06132_),
    .A1(_05939_),
    .A2(_06090_));
 sg13g2_nor2_1 _13320_ (.A(_06124_),
    .B(_06132_),
    .Y(_06133_));
 sg13g2_xor2_1 _13321_ (.B(_04766_),
    .A(_04765_),
    .X(_06134_));
 sg13g2_a22oi_1 _13322_ (.Y(_06135_),
    .B1(_00010_),
    .B2(_06134_),
    .A2(net501),
    .A1(net3922));
 sg13g2_o21ai_1 _13323_ (.B1(_06135_),
    .Y(_00590_),
    .A1(_06122_),
    .A2(_06133_));
 sg13g2_a21o_1 _13324_ (.A2(_06098_),
    .A1(_06095_),
    .B1(_06099_),
    .X(_06136_));
 sg13g2_nand3_1 _13325_ (.B(_06100_),
    .C(_06136_),
    .A(_05939_),
    .Y(_06137_));
 sg13g2_o21ai_1 _13326_ (.B1(_06137_),
    .Y(_06138_),
    .A1(_05939_),
    .A2(_06077_));
 sg13g2_o21ai_1 _13327_ (.B1(_06121_),
    .Y(_06139_),
    .A1(_06124_),
    .A2(_06138_));
 sg13g2_xnor2_1 _13328_ (.Y(_06140_),
    .A(_04763_),
    .B(_04767_));
 sg13g2_a21oi_1 _13329_ (.A1(net3666),
    .A2(_06140_),
    .Y(_06141_),
    .B1(net3920));
 sg13g2_a22oi_1 _13330_ (.Y(_00591_),
    .B1(_06139_),
    .B2(_06141_),
    .A2(_03441_),
    .A1(net3920));
 sg13g2_nand3_1 _13331_ (.B(_06100_),
    .C(_06101_),
    .A(_06093_),
    .Y(_06142_));
 sg13g2_a21oi_1 _13332_ (.A1(_06102_),
    .A2(_06142_),
    .Y(_06143_),
    .B1(_05940_));
 sg13g2_a21oi_1 _13333_ (.A1(_05940_),
    .A2(_06054_),
    .Y(_06144_),
    .B1(_06143_));
 sg13g2_o21ai_1 _13334_ (.B1(_06121_),
    .Y(_06145_),
    .A1(_06124_),
    .A2(_06144_));
 sg13g2_or3_1 _13335_ (.A(_04761_),
    .B(_04762_),
    .C(_04768_),
    .X(_06146_));
 sg13g2_and2_1 _13336_ (.A(_04769_),
    .B(_06146_),
    .X(_06147_));
 sg13g2_a21oi_1 _13337_ (.A1(net3666),
    .A2(_06147_),
    .Y(_06148_),
    .B1(net3920));
 sg13g2_a22oi_1 _13338_ (.Y(_00592_),
    .B1(_06145_),
    .B2(_06148_),
    .A2(_03440_),
    .A1(net3920));
 sg13g2_o21ai_1 _13339_ (.B1(net4530),
    .Y(_06149_),
    .A1(_04759_),
    .A2(_04770_));
 sg13g2_a21oi_1 _13340_ (.A1(_04772_),
    .A2(_06120_),
    .Y(_06150_),
    .B1(_06149_));
 sg13g2_a21oi_1 _13341_ (.A1(net3920),
    .A2(_03439_),
    .Y(_00593_),
    .B1(_06150_));
 sg13g2_mux2_1 _13342_ (.A0(net3844),
    .A1(net3843),
    .S(\spiking_network_top_uut.all_data_out[668] ),
    .X(_06151_));
 sg13g2_nor2b_1 _13343_ (.A(\spiking_network_top_uut.all_data_out[668] ),
    .B_N(net3846),
    .Y(_06152_));
 sg13g2_a21oi_1 _13344_ (.A1(\spiking_network_top_uut.all_data_out[668] ),
    .A2(net3845),
    .Y(_06153_),
    .B1(_06152_));
 sg13g2_a21oi_1 _13345_ (.A1(\spiking_network_top_uut.all_data_out[669] ),
    .A2(_06151_),
    .Y(_06154_),
    .B1(\spiking_network_top_uut.all_data_out[670] ));
 sg13g2_o21ai_1 _13346_ (.B1(_06154_),
    .Y(_06155_),
    .A1(\spiking_network_top_uut.all_data_out[669] ),
    .A2(_06153_));
 sg13g2_mux2_1 _13347_ (.A0(net3841),
    .A1(net3900),
    .S(\spiking_network_top_uut.all_data_out[668] ),
    .X(_06156_));
 sg13g2_nand2_1 _13348_ (.Y(_06157_),
    .A(\spiking_network_top_uut.all_data_out[669] ),
    .B(_06156_));
 sg13g2_a21oi_1 _13349_ (.A1(\spiking_network_top_uut.all_data_out[668] ),
    .A2(_03667_),
    .Y(_06158_),
    .B1(\spiking_network_top_uut.all_data_out[669] ));
 sg13g2_o21ai_1 _13350_ (.B1(_06158_),
    .Y(_06159_),
    .A1(\spiking_network_top_uut.all_data_out[668] ),
    .A2(net3842));
 sg13g2_nand3_1 _13351_ (.B(_06157_),
    .C(_06159_),
    .A(\spiking_network_top_uut.all_data_out[670] ),
    .Y(_06160_));
 sg13g2_nand3_1 _13352_ (.B(_06155_),
    .C(_06160_),
    .A(net4553),
    .Y(_06161_));
 sg13g2_o21ai_1 _13353_ (.B1(_06161_),
    .Y(_00594_),
    .A1(net4548),
    .A2(_03671_));
 sg13g2_mux2_1 _13354_ (.A0(net253),
    .A1(net142),
    .S(net4548),
    .X(_00595_));
 sg13g2_a21oi_1 _13355_ (.A1(\spiking_network_top_uut.all_data_out[664] ),
    .A2(_03666_),
    .Y(_06162_),
    .B1(\spiking_network_top_uut.all_data_out[665] ));
 sg13g2_o21ai_1 _13356_ (.B1(_06162_),
    .Y(_06163_),
    .A1(\spiking_network_top_uut.all_data_out[664] ),
    .A2(net3894));
 sg13g2_mux2_1 _13357_ (.A0(net3893),
    .A1(net3892),
    .S(\spiking_network_top_uut.all_data_out[664] ),
    .X(_06164_));
 sg13g2_nand2_1 _13358_ (.Y(_06165_),
    .A(\spiking_network_top_uut.all_data_out[665] ),
    .B(_06164_));
 sg13g2_nand3_1 _13359_ (.B(_06163_),
    .C(_06165_),
    .A(\spiking_network_top_uut.all_data_out[666] ),
    .Y(_06166_));
 sg13g2_mux2_1 _13360_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[2] ),
    .A1(net3895),
    .S(\spiking_network_top_uut.all_data_out[664] ),
    .X(_06167_));
 sg13g2_nor2b_1 _13361_ (.A(\spiking_network_top_uut.all_data_out[664] ),
    .B_N(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[0] ),
    .Y(_06168_));
 sg13g2_a21oi_1 _13362_ (.A1(\spiking_network_top_uut.all_data_out[664] ),
    .A2(net3897),
    .Y(_06169_),
    .B1(_06168_));
 sg13g2_a21oi_1 _13363_ (.A1(\spiking_network_top_uut.all_data_out[665] ),
    .A2(_06167_),
    .Y(_06170_),
    .B1(\spiking_network_top_uut.all_data_out[666] ));
 sg13g2_o21ai_1 _13364_ (.B1(_06170_),
    .Y(_06171_),
    .A1(\spiking_network_top_uut.all_data_out[665] ),
    .A2(_06169_));
 sg13g2_nand3_1 _13365_ (.B(_06166_),
    .C(_06171_),
    .A(net4547),
    .Y(_06172_));
 sg13g2_o21ai_1 _13366_ (.B1(_06172_),
    .Y(_00596_),
    .A1(net4548),
    .A2(_03672_));
 sg13g2_nor2_1 _13367_ (.A(net4548),
    .B(net123),
    .Y(_06173_));
 sg13g2_a21oi_1 _13368_ (.A1(net4548),
    .A2(_03672_),
    .Y(_00597_),
    .B1(_06173_));
 sg13g2_mux4_1 _13369_ (.S0(\spiking_network_top_uut.all_data_out[660] ),
    .A0(net3891),
    .A1(net3890),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[2] ),
    .A3(net3888),
    .S1(\spiking_network_top_uut.all_data_out[661] ),
    .X(_06174_));
 sg13g2_mux2_1 _13370_ (.A0(net3886),
    .A1(net3885),
    .S(\spiking_network_top_uut.all_data_out[660] ),
    .X(_06175_));
 sg13g2_nor2b_1 _13371_ (.A(\spiking_network_top_uut.all_data_out[660] ),
    .B_N(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[4] ),
    .Y(_06176_));
 sg13g2_a21oi_1 _13372_ (.A1(\spiking_network_top_uut.all_data_out[660] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[5] ),
    .Y(_06177_),
    .B1(_06176_));
 sg13g2_o21ai_1 _13373_ (.B1(\spiking_network_top_uut.all_data_out[662] ),
    .Y(_06178_),
    .A1(\spiking_network_top_uut.all_data_out[661] ),
    .A2(_06177_));
 sg13g2_a21oi_1 _13374_ (.A1(\spiking_network_top_uut.all_data_out[661] ),
    .A2(_06175_),
    .Y(_06179_),
    .B1(_06178_));
 sg13g2_o21ai_1 _13375_ (.B1(net4561),
    .Y(_06180_),
    .A1(\spiking_network_top_uut.all_data_out[662] ),
    .A2(_06174_));
 sg13g2_nand2_1 _13376_ (.Y(_06181_),
    .A(net3935),
    .B(net170));
 sg13g2_o21ai_1 _13377_ (.B1(_06181_),
    .Y(_00598_),
    .A1(_06179_),
    .A2(_06180_));
 sg13g2_mux2_1 _13378_ (.A0(net466),
    .A1(net170),
    .S(net4571),
    .X(_00599_));
 sg13g2_mux4_1 _13379_ (.S0(\spiking_network_top_uut.all_data_out[656] ),
    .A0(net3884),
    .A1(net3883),
    .A2(net3882),
    .A3(net3881),
    .S1(\spiking_network_top_uut.all_data_out[657] ),
    .X(_06182_));
 sg13g2_mux2_1 _13380_ (.A0(net3878),
    .A1(net3877),
    .S(\spiking_network_top_uut.all_data_out[656] ),
    .X(_06183_));
 sg13g2_nor2b_1 _13381_ (.A(\spiking_network_top_uut.all_data_out[656] ),
    .B_N(net3880),
    .Y(_06184_));
 sg13g2_a21oi_1 _13382_ (.A1(\spiking_network_top_uut.all_data_out[656] ),
    .A2(net3879),
    .Y(_06185_),
    .B1(_06184_));
 sg13g2_o21ai_1 _13383_ (.B1(\spiking_network_top_uut.all_data_out[658] ),
    .Y(_06186_),
    .A1(\spiking_network_top_uut.all_data_out[657] ),
    .A2(_06185_));
 sg13g2_a21oi_1 _13384_ (.A1(\spiking_network_top_uut.all_data_out[657] ),
    .A2(_06183_),
    .Y(_06187_),
    .B1(_06186_));
 sg13g2_o21ai_1 _13385_ (.B1(net4555),
    .Y(_06188_),
    .A1(\spiking_network_top_uut.all_data_out[658] ),
    .A2(_06182_));
 sg13g2_nand2_1 _13386_ (.Y(_06189_),
    .A(net3938),
    .B(net199));
 sg13g2_o21ai_1 _13387_ (.B1(_06189_),
    .Y(_00600_),
    .A1(_06187_),
    .A2(_06188_));
 sg13g2_mux2_1 _13388_ (.A0(net373),
    .A1(net199),
    .S(net4556),
    .X(_00601_));
 sg13g2_mux4_1 _13389_ (.S0(\spiking_network_top_uut.all_data_out[652] ),
    .A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[0] ),
    .A1(net3875),
    .A2(net3874),
    .A3(net3873),
    .S1(\spiking_network_top_uut.all_data_out[653] ),
    .X(_06190_));
 sg13g2_mux2_1 _13390_ (.A0(net3870),
    .A1(net3869),
    .S(\spiking_network_top_uut.all_data_out[652] ),
    .X(_06191_));
 sg13g2_nor2b_1 _13391_ (.A(\spiking_network_top_uut.all_data_out[652] ),
    .B_N(net3872),
    .Y(_06192_));
 sg13g2_a21oi_1 _13392_ (.A1(\spiking_network_top_uut.all_data_out[652] ),
    .A2(net3871),
    .Y(_06193_),
    .B1(_06192_));
 sg13g2_o21ai_1 _13393_ (.B1(\spiking_network_top_uut.all_data_out[654] ),
    .Y(_06194_),
    .A1(\spiking_network_top_uut.all_data_out[653] ),
    .A2(_06193_));
 sg13g2_a21oi_1 _13394_ (.A1(\spiking_network_top_uut.all_data_out[653] ),
    .A2(_06191_),
    .Y(_06195_),
    .B1(_06194_));
 sg13g2_o21ai_1 _13395_ (.B1(net4566),
    .Y(_06196_),
    .A1(\spiking_network_top_uut.all_data_out[654] ),
    .A2(_06190_));
 sg13g2_nand2_1 _13396_ (.Y(_06197_),
    .A(net3937),
    .B(net98));
 sg13g2_o21ai_1 _13397_ (.B1(_06197_),
    .Y(_00602_),
    .A1(_06195_),
    .A2(_06196_));
 sg13g2_mux2_1 _13398_ (.A0(net284),
    .A1(net98),
    .S(net4566),
    .X(_00603_));
 sg13g2_nand2b_1 _13399_ (.Y(_06198_),
    .B(\spiking_network_top_uut.all_data_out[648] ),
    .A_N(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[5] ));
 sg13g2_nor2_1 _13400_ (.A(\spiking_network_top_uut.all_data_out[648] ),
    .B(net3864),
    .Y(_06199_));
 sg13g2_nor2_1 _13401_ (.A(\spiking_network_top_uut.all_data_out[649] ),
    .B(_06199_),
    .Y(_06200_));
 sg13g2_mux2_1 _13402_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[6] ),
    .A1(net3861),
    .S(\spiking_network_top_uut.all_data_out[648] ),
    .X(_06201_));
 sg13g2_a221oi_1 _13403_ (.B2(\spiking_network_top_uut.all_data_out[649] ),
    .C1(_03600_),
    .B1(_06201_),
    .A1(_06198_),
    .Y(_06202_),
    .A2(_06200_));
 sg13g2_mux4_1 _13404_ (.S0(\spiking_network_top_uut.all_data_out[648] ),
    .A0(net3868),
    .A1(net3867),
    .A2(net3866),
    .A3(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[3] ),
    .S1(\spiking_network_top_uut.all_data_out[649] ),
    .X(_06203_));
 sg13g2_o21ai_1 _13405_ (.B1(net4564),
    .Y(_06204_),
    .A1(\spiking_network_top_uut.all_data_out[650] ),
    .A2(_06203_));
 sg13g2_nand2_1 _13406_ (.Y(_06205_),
    .A(net3936),
    .B(net140));
 sg13g2_o21ai_1 _13407_ (.B1(_06205_),
    .Y(_00604_),
    .A1(_06202_),
    .A2(_06204_));
 sg13g2_mux2_1 _13408_ (.A0(net326),
    .A1(net140),
    .S(net4564),
    .X(_00605_));
 sg13g2_nand2_1 _13409_ (.Y(_06206_),
    .A(\spiking_network_top_uut.all_data_out[644] ),
    .B(_03664_));
 sg13g2_nor2_1 _13410_ (.A(\spiking_network_top_uut.all_data_out[644] ),
    .B(net3856),
    .Y(_06207_));
 sg13g2_nor2_1 _13411_ (.A(\spiking_network_top_uut.all_data_out[645] ),
    .B(_06207_),
    .Y(_06208_));
 sg13g2_mux2_1 _13412_ (.A0(net3855),
    .A1(net3854),
    .S(\spiking_network_top_uut.all_data_out[644] ),
    .X(_06209_));
 sg13g2_a221oi_1 _13413_ (.B2(\spiking_network_top_uut.all_data_out[645] ),
    .C1(_03528_),
    .B1(_06209_),
    .A1(_06206_),
    .Y(_06210_),
    .A2(_06208_));
 sg13g2_mux4_1 _13414_ (.S0(\spiking_network_top_uut.all_data_out[644] ),
    .A0(net3860),
    .A1(net3859),
    .A2(net3858),
    .A3(net3857),
    .S1(\spiking_network_top_uut.all_data_out[645] ),
    .X(_06211_));
 sg13g2_o21ai_1 _13415_ (.B1(net4534),
    .Y(_06212_),
    .A1(\spiking_network_top_uut.all_data_out[646] ),
    .A2(_06211_));
 sg13g2_nand2_1 _13416_ (.Y(_06213_),
    .A(net3932),
    .B(net82));
 sg13g2_o21ai_1 _13417_ (.B1(_06213_),
    .Y(_00606_),
    .A1(_06210_),
    .A2(_06212_));
 sg13g2_mux2_1 _13418_ (.A0(net231),
    .A1(net82),
    .S(net4534),
    .X(_00607_));
 sg13g2_mux2_1 _13419_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[2] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[3] ),
    .S(\spiking_network_top_uut.all_data_out[640] ),
    .X(_06214_));
 sg13g2_nor2b_1 _13420_ (.A(\spiking_network_top_uut.all_data_out[640] ),
    .B_N(net3853),
    .Y(_06215_));
 sg13g2_a21oi_1 _13421_ (.A1(\spiking_network_top_uut.all_data_out[640] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[1] ),
    .Y(_06216_),
    .B1(_06215_));
 sg13g2_a21oi_1 _13422_ (.A1(\spiking_network_top_uut.all_data_out[641] ),
    .A2(_06214_),
    .Y(_06217_),
    .B1(\spiking_network_top_uut.all_data_out[642] ));
 sg13g2_o21ai_1 _13423_ (.B1(_06217_),
    .Y(_06218_),
    .A1(\spiking_network_top_uut.all_data_out[641] ),
    .A2(_06216_));
 sg13g2_mux2_1 _13424_ (.A0(net3848),
    .A1(net3847),
    .S(\spiking_network_top_uut.all_data_out[640] ),
    .X(_06219_));
 sg13g2_nand2_1 _13425_ (.Y(_06220_),
    .A(\spiking_network_top_uut.all_data_out[641] ),
    .B(_06219_));
 sg13g2_a21oi_1 _13426_ (.A1(\spiking_network_top_uut.all_data_out[640] ),
    .A2(_03663_),
    .Y(_06221_),
    .B1(\spiking_network_top_uut.all_data_out[641] ));
 sg13g2_o21ai_1 _13427_ (.B1(_06221_),
    .Y(_06222_),
    .A1(\spiking_network_top_uut.all_data_out[640] ),
    .A2(net3849));
 sg13g2_nand3_1 _13428_ (.B(_06220_),
    .C(_06222_),
    .A(\spiking_network_top_uut.all_data_out[642] ),
    .Y(_06223_));
 sg13g2_nand3_1 _13429_ (.B(_06218_),
    .C(_06223_),
    .A(net4538),
    .Y(_06224_));
 sg13g2_o21ai_1 _13430_ (.B1(_06224_),
    .Y(_00608_),
    .A1(net4537),
    .A2(_03673_));
 sg13g2_nor3_2 _13431_ (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[2] ),
    .B(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[1] ),
    .C(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[0] ),
    .Y(_06225_));
 sg13g2_nor2b_2 _13432_ (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[3] ),
    .B_N(_06225_),
    .Y(_06226_));
 sg13g2_nor2b_2 _13433_ (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[4] ),
    .B_N(_06226_),
    .Y(_06227_));
 sg13g2_nand2b_2 _13434_ (.Y(_06228_),
    .B(_06226_),
    .A_N(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[4] ));
 sg13g2_o21ai_1 _13435_ (.B1(net4529),
    .Y(_06229_),
    .A1(net3657),
    .A2(net3705));
 sg13g2_nor2b_1 _13436_ (.A(net3656),
    .B_N(_00060_),
    .Y(_06230_));
 sg13g2_a21oi_1 _13437_ (.A1(net4283),
    .A2(net3656),
    .Y(_06231_),
    .B1(_06230_));
 sg13g2_nand2_1 _13438_ (.Y(_06232_),
    .A(net316),
    .B(_06229_));
 sg13g2_o21ai_1 _13439_ (.B1(_06232_),
    .Y(_00609_),
    .A1(_06229_),
    .A2(_06231_));
 sg13g2_xor2_1 _13440_ (.B(net316),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[1] ),
    .X(_06233_));
 sg13g2_nor2_1 _13441_ (.A(net3656),
    .B(_06233_),
    .Y(_06234_));
 sg13g2_a21oi_1 _13442_ (.A1(net4280),
    .A2(net3656),
    .Y(_06235_),
    .B1(_06234_));
 sg13g2_nand2_1 _13443_ (.Y(_06236_),
    .A(net414),
    .B(_06229_));
 sg13g2_o21ai_1 _13444_ (.B1(_06236_),
    .Y(_00610_),
    .A1(_06229_),
    .A2(_06235_));
 sg13g2_o21ai_1 _13445_ (.B1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[2] ),
    .Y(_06237_),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[1] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[0] ));
 sg13g2_nor2b_1 _13446_ (.A(_06225_),
    .B_N(_06237_),
    .Y(_06238_));
 sg13g2_nor2_1 _13447_ (.A(net3656),
    .B(_06238_),
    .Y(_06239_));
 sg13g2_a21oi_1 _13448_ (.A1(net4276),
    .A2(net3656),
    .Y(_06240_),
    .B1(_06239_));
 sg13g2_nand2_1 _13449_ (.Y(_06241_),
    .A(net160),
    .B(_06229_));
 sg13g2_o21ai_1 _13450_ (.B1(_06241_),
    .Y(_00611_),
    .A1(_06229_),
    .A2(_06240_));
 sg13g2_nand2_1 _13451_ (.Y(_06242_),
    .A(net4273),
    .B(net3656));
 sg13g2_xnor2_1 _13452_ (.Y(_06243_),
    .A(net431),
    .B(_06225_));
 sg13g2_o21ai_1 _13453_ (.B1(_06242_),
    .Y(_06244_),
    .A1(net3656),
    .A2(_06243_));
 sg13g2_mux2_1 _13454_ (.A0(_06244_),
    .A1(net431),
    .S(_06229_),
    .X(_00612_));
 sg13g2_nand2_1 _13455_ (.Y(_06245_),
    .A(net3922),
    .B(net282));
 sg13g2_nand2b_1 _13456_ (.Y(_06246_),
    .B(net282),
    .A_N(_06226_));
 sg13g2_a21oi_1 _13457_ (.A1(net3705),
    .A2(_06246_),
    .Y(_06247_),
    .B1(net3657));
 sg13g2_a21oi_1 _13458_ (.A1(net4269),
    .A2(net3657),
    .Y(_06248_),
    .B1(_06247_));
 sg13g2_o21ai_1 _13459_ (.B1(_06245_),
    .Y(_00613_),
    .A1(_06229_),
    .A2(_06248_));
 sg13g2_mux2_1 _13460_ (.A0(net306),
    .A1(net120),
    .S(net4537),
    .X(_00614_));
 sg13g2_nor2_1 _13461_ (.A(_00055_),
    .B(net3741),
    .Y(_06249_));
 sg13g2_nor2_2 _13462_ (.A(net3749),
    .B(_06249_),
    .Y(_06250_));
 sg13g2_nor2_1 _13463_ (.A(_00055_),
    .B(_06250_),
    .Y(_06251_));
 sg13g2_nand2b_1 _13464_ (.Y(_06252_),
    .B(_06250_),
    .A_N(_00055_));
 sg13g2_o21ai_1 _13465_ (.B1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ),
    .Y(_06253_),
    .A1(_00055_),
    .A2(_06250_));
 sg13g2_inv_1 _13466_ (.Y(_06254_),
    .A(_06253_));
 sg13g2_a21o_1 _13467_ (.A2(net3747),
    .A1(_00056_),
    .B1(_06250_),
    .X(_06255_));
 sg13g2_and2_1 _13468_ (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ),
    .B(_06255_),
    .X(_06256_));
 sg13g2_and2_1 _13469_ (.A(_00057_),
    .B(net3747),
    .X(_06257_));
 sg13g2_o21ai_1 _13470_ (.B1(net3917),
    .Y(_06258_),
    .A1(_00056_),
    .A2(net3905));
 sg13g2_a21oi_1 _13471_ (.A1(net3905),
    .A2(_06249_),
    .Y(_06259_),
    .B1(_06258_));
 sg13g2_o21ai_1 _13472_ (.B1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ),
    .Y(_06260_),
    .A1(_06257_),
    .A2(_06259_));
 sg13g2_o21ai_1 _13473_ (.B1(net3914),
    .Y(_06261_),
    .A1(_00055_),
    .A2(net3910));
 sg13g2_a221oi_1 _13474_ (.B2(_00056_),
    .C1(net3747),
    .B1(net3901),
    .A1(_00057_),
    .Y(_06262_),
    .A2(net3739));
 sg13g2_a22oi_1 _13475_ (.Y(_06263_),
    .B1(_06261_),
    .B2(_06262_),
    .A2(net3747),
    .A1(_03482_));
 sg13g2_nor2b_1 _13476_ (.A(_06263_),
    .B_N(_00058_),
    .Y(_06264_));
 sg13g2_or3_1 _13477_ (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ),
    .B(_06257_),
    .C(_06259_),
    .X(_06265_));
 sg13g2_nand2_1 _13478_ (.Y(_06266_),
    .A(_06260_),
    .B(_06265_));
 sg13g2_o21ai_1 _13479_ (.B1(_06260_),
    .Y(_06267_),
    .A1(_06264_),
    .A2(_06266_));
 sg13g2_xnor2_1 _13480_ (.Y(_06268_),
    .A(_00057_),
    .B(_06255_));
 sg13g2_a21o_1 _13481_ (.A2(_06268_),
    .A1(_06267_),
    .B1(_06256_),
    .X(_06269_));
 sg13g2_xnor2_1 _13482_ (.Y(_06270_),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ),
    .B(_06251_));
 sg13g2_a21oi_1 _13483_ (.A1(_06269_),
    .A2(_06270_),
    .Y(_06271_),
    .B1(_06254_));
 sg13g2_a22oi_1 _13484_ (.Y(_06272_),
    .B1(_06252_),
    .B2(_06271_),
    .A2(_06250_),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ));
 sg13g2_a21oi_2 _13485_ (.B1(_06272_),
    .Y(_06273_),
    .A2(_00055_),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ));
 sg13g2_inv_1 _13486_ (.Y(_06274_),
    .A(_06273_));
 sg13g2_mux2_1 _13487_ (.A0(net4599),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[643] ),
    .X(_06275_));
 sg13g2_nand2_1 _13488_ (.Y(_06276_),
    .A(\spiking_network_top_uut.all_data_out[193] ),
    .B(_06275_));
 sg13g2_mux2_1 _13489_ (.A0(net4598),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[647] ),
    .X(_06277_));
 sg13g2_nand2_1 _13490_ (.Y(_06278_),
    .A(\spiking_network_top_uut.all_data_out[195] ),
    .B(_06277_));
 sg13g2_nor2_1 _13491_ (.A(_06276_),
    .B(_06278_),
    .Y(_06279_));
 sg13g2_nand4_1 _13492_ (.B(\spiking_network_top_uut.all_data_out[194] ),
    .C(_06275_),
    .A(\spiking_network_top_uut.all_data_out[192] ),
    .Y(_06280_),
    .D(_06277_));
 sg13g2_inv_1 _13493_ (.Y(_06281_),
    .A(_06280_));
 sg13g2_xor2_1 _13494_ (.B(_06278_),
    .A(_06276_),
    .X(_06282_));
 sg13g2_a21oi_2 _13495_ (.B1(_06279_),
    .Y(_06283_),
    .A2(_06282_),
    .A1(_06280_));
 sg13g2_mux2_2 _13496_ (.A0(net4597),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[651] ),
    .X(_06284_));
 sg13g2_nand2_1 _13497_ (.Y(_06285_),
    .A(\spiking_network_top_uut.all_data_out[197] ),
    .B(_06284_));
 sg13g2_mux2_2 _13498_ (.A0(net4596),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[655] ),
    .X(_06286_));
 sg13g2_nand2_1 _13499_ (.Y(_06287_),
    .A(\spiking_network_top_uut.all_data_out[199] ),
    .B(_06286_));
 sg13g2_nor2_1 _13500_ (.A(_06285_),
    .B(_06287_),
    .Y(_06288_));
 sg13g2_nand2_1 _13501_ (.Y(_06289_),
    .A(\spiking_network_top_uut.all_data_out[196] ),
    .B(_06284_));
 sg13g2_nand2_1 _13502_ (.Y(_06290_),
    .A(\spiking_network_top_uut.all_data_out[198] ),
    .B(_06286_));
 sg13g2_or2_1 _13503_ (.X(_06291_),
    .B(_06290_),
    .A(_06289_));
 sg13g2_xor2_1 _13504_ (.B(_06287_),
    .A(_06285_),
    .X(_06292_));
 sg13g2_a21oi_2 _13505_ (.B1(_06288_),
    .Y(_06293_),
    .A2(_06292_),
    .A1(_06291_));
 sg13g2_mux2_2 _13506_ (.A0(net4595),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[659] ),
    .X(_06294_));
 sg13g2_mux2_2 _13507_ (.A0(net4594),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[663] ),
    .X(_06295_));
 sg13g2_a22oi_1 _13508_ (.Y(_06296_),
    .B1(_06295_),
    .B2(\spiking_network_top_uut.all_data_out[203] ),
    .A2(_06294_),
    .A1(\spiking_network_top_uut.all_data_out[201] ));
 sg13g2_and4_1 _13509_ (.A(\spiking_network_top_uut.all_data_out[201] ),
    .B(\spiking_network_top_uut.all_data_out[203] ),
    .C(_06294_),
    .D(_06295_),
    .X(_06297_));
 sg13g2_nand4_1 _13510_ (.B(\spiking_network_top_uut.all_data_out[203] ),
    .C(_06294_),
    .A(\spiking_network_top_uut.all_data_out[201] ),
    .Y(_06298_),
    .D(_06295_));
 sg13g2_and4_2 _13511_ (.A(\spiking_network_top_uut.all_data_out[200] ),
    .B(\spiking_network_top_uut.all_data_out[202] ),
    .C(_06294_),
    .D(_06295_),
    .X(_06299_));
 sg13g2_nand4_1 _13512_ (.B(\spiking_network_top_uut.all_data_out[202] ),
    .C(_06294_),
    .A(\spiking_network_top_uut.all_data_out[200] ),
    .Y(_06300_),
    .D(_06295_));
 sg13g2_nand3b_1 _13513_ (.B(_06298_),
    .C(_06299_),
    .Y(_06301_),
    .A_N(_06296_));
 sg13g2_a21oi_2 _13514_ (.B1(_06296_),
    .Y(_06302_),
    .A2(_06299_),
    .A1(_06298_));
 sg13g2_mux2_2 _13515_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.spike_out ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[667] ),
    .X(_06303_));
 sg13g2_mux2_2 _13516_ (.A0(net4592),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[671] ),
    .X(_06304_));
 sg13g2_and4_1 _13517_ (.A(\spiking_network_top_uut.all_data_out[205] ),
    .B(\spiking_network_top_uut.all_data_out[207] ),
    .C(_06303_),
    .D(_06304_),
    .X(_06305_));
 sg13g2_nand4_1 _13518_ (.B(\spiking_network_top_uut.all_data_out[207] ),
    .C(_06303_),
    .A(\spiking_network_top_uut.all_data_out[205] ),
    .Y(_06306_),
    .D(_06304_));
 sg13g2_and4_1 _13519_ (.A(\spiking_network_top_uut.all_data_out[204] ),
    .B(\spiking_network_top_uut.all_data_out[206] ),
    .C(_06303_),
    .D(_06304_),
    .X(_06307_));
 sg13g2_a22oi_1 _13520_ (.Y(_06308_),
    .B1(_06304_),
    .B2(\spiking_network_top_uut.all_data_out[207] ),
    .A2(_06303_),
    .A1(\spiking_network_top_uut.all_data_out[205] ));
 sg13g2_or3_2 _13521_ (.A(_06305_),
    .B(_06307_),
    .C(_06308_),
    .X(_06309_));
 sg13g2_o21ai_1 _13522_ (.B1(_06306_),
    .Y(_06310_),
    .A1(_06307_),
    .A2(_06308_));
 sg13g2_nand3b_1 _13523_ (.B(_06302_),
    .C(_06310_),
    .Y(_06311_),
    .A_N(_06293_));
 sg13g2_or2_1 _13524_ (.X(_06312_),
    .B(_06311_),
    .A(_06283_));
 sg13g2_inv_1 _13525_ (.Y(_06313_),
    .A(_06312_));
 sg13g2_nor2_1 _13526_ (.A(_06302_),
    .B(_06310_),
    .Y(_06314_));
 sg13g2_nand2_1 _13527_ (.Y(_06315_),
    .A(_06293_),
    .B(_06314_));
 sg13g2_mux2_2 _13528_ (.A0(_06311_),
    .A1(_06315_),
    .S(_06283_),
    .X(_06316_));
 sg13g2_xnor2_1 _13529_ (.Y(_06317_),
    .A(_06252_),
    .B(_06271_));
 sg13g2_xor2_1 _13530_ (.B(_06317_),
    .A(_06316_),
    .X(_06318_));
 sg13g2_o21ai_1 _13531_ (.B1(_06307_),
    .Y(_06319_),
    .A1(_06305_),
    .A2(_06308_));
 sg13g2_o21ai_1 _13532_ (.B1(_06300_),
    .Y(_06320_),
    .A1(_06296_),
    .A2(_06297_));
 sg13g2_o21ai_1 _13533_ (.B1(_06299_),
    .Y(_06321_),
    .A1(_06296_),
    .A2(_06297_));
 sg13g2_nand3b_1 _13534_ (.B(_06298_),
    .C(_06300_),
    .Y(_06322_),
    .A_N(_06296_));
 sg13g2_a22oi_1 _13535_ (.Y(_06323_),
    .B1(_06321_),
    .B2(_06322_),
    .A2(_06319_),
    .A1(_06309_));
 sg13g2_xor2_1 _13536_ (.B(_06292_),
    .A(_06291_),
    .X(_06324_));
 sg13g2_xnor2_1 _13537_ (.Y(_06325_),
    .A(_06291_),
    .B(_06292_));
 sg13g2_and4_1 _13538_ (.A(_06309_),
    .B(_06319_),
    .C(_06321_),
    .D(_06322_),
    .X(_06326_));
 sg13g2_nand4_1 _13539_ (.B(_06319_),
    .C(_06321_),
    .A(_06309_),
    .Y(_06327_),
    .D(_06322_));
 sg13g2_and4_1 _13540_ (.A(_06301_),
    .B(_06309_),
    .C(_06319_),
    .D(_06320_),
    .X(_06328_));
 sg13g2_a22oi_1 _13541_ (.Y(_06329_),
    .B1(_06320_),
    .B2(_06301_),
    .A2(_06319_),
    .A1(_06309_));
 sg13g2_nor3_2 _13542_ (.A(_06323_),
    .B(_06324_),
    .C(_06326_),
    .Y(_06330_));
 sg13g2_a21oi_2 _13543_ (.B1(_06323_),
    .Y(_06331_),
    .A2(_06327_),
    .A1(_06325_));
 sg13g2_xor2_1 _13544_ (.B(_06310_),
    .A(_06302_),
    .X(_06332_));
 sg13g2_xnor2_1 _13545_ (.Y(_06333_),
    .A(_06293_),
    .B(_06332_));
 sg13g2_nand2b_1 _13546_ (.Y(_06334_),
    .B(_06333_),
    .A_N(_06331_));
 sg13g2_xnor2_1 _13547_ (.Y(_06335_),
    .A(_06331_),
    .B(_06333_));
 sg13g2_nand2b_1 _13548_ (.Y(_06336_),
    .B(_06335_),
    .A_N(_06283_));
 sg13g2_nand2_1 _13549_ (.Y(_06337_),
    .A(_06334_),
    .B(_06336_));
 sg13g2_nand2_1 _13550_ (.Y(_06338_),
    .A(_06311_),
    .B(_06315_));
 sg13g2_xor2_1 _13551_ (.B(_06338_),
    .A(_06283_),
    .X(_06339_));
 sg13g2_and2_1 _13552_ (.A(_06337_),
    .B(_06339_),
    .X(_06340_));
 sg13g2_xor2_1 _13553_ (.B(_06339_),
    .A(_06337_),
    .X(_06341_));
 sg13g2_xnor2_1 _13554_ (.Y(_06342_),
    .A(_06269_),
    .B(_06270_));
 sg13g2_inv_1 _13555_ (.Y(_06343_),
    .A(_06342_));
 sg13g2_a21oi_1 _13556_ (.A1(_06341_),
    .A2(_06343_),
    .Y(_06344_),
    .B1(_06340_));
 sg13g2_nand2b_1 _13557_ (.Y(_06345_),
    .B(_06318_),
    .A_N(_06344_));
 sg13g2_xor2_1 _13558_ (.B(_06342_),
    .A(_06341_),
    .X(_06346_));
 sg13g2_a22oi_1 _13559_ (.Y(_06347_),
    .B1(_06304_),
    .B2(\spiking_network_top_uut.all_data_out[206] ),
    .A2(_06303_),
    .A1(\spiking_network_top_uut.all_data_out[204] ));
 sg13g2_nor2_2 _13560_ (.A(_06307_),
    .B(_06347_),
    .Y(_06348_));
 sg13g2_a22oi_1 _13561_ (.Y(_06349_),
    .B1(_06295_),
    .B2(\spiking_network_top_uut.all_data_out[202] ),
    .A2(_06294_),
    .A1(\spiking_network_top_uut.all_data_out[200] ));
 sg13g2_nor2_2 _13562_ (.A(_06299_),
    .B(_06349_),
    .Y(_06350_));
 sg13g2_and2_1 _13563_ (.A(_06348_),
    .B(_06350_),
    .X(_06351_));
 sg13g2_xor2_1 _13564_ (.B(_06290_),
    .A(_06289_),
    .X(_06352_));
 sg13g2_xor2_1 _13565_ (.B(_06350_),
    .A(_06348_),
    .X(_06353_));
 sg13g2_a21oi_2 _13566_ (.B1(_06351_),
    .Y(_06354_),
    .A2(_06353_),
    .A1(_06352_));
 sg13g2_nor3_2 _13567_ (.A(_06325_),
    .B(_06328_),
    .C(_06329_),
    .Y(_06355_));
 sg13g2_nor3_1 _13568_ (.A(_06330_),
    .B(_06354_),
    .C(_06355_),
    .Y(_06356_));
 sg13g2_or3_1 _13569_ (.A(_06330_),
    .B(_06354_),
    .C(_06355_),
    .X(_06357_));
 sg13g2_xnor2_1 _13570_ (.Y(_06358_),
    .A(_06280_),
    .B(_06282_));
 sg13g2_o21ai_1 _13571_ (.B1(_06354_),
    .Y(_06359_),
    .A1(_06330_),
    .A2(_06355_));
 sg13g2_nand3_1 _13572_ (.B(_06358_),
    .C(_06359_),
    .A(_06357_),
    .Y(_06360_));
 sg13g2_a21o_2 _13573_ (.A2(_06359_),
    .A1(_06358_),
    .B1(_06356_),
    .X(_06361_));
 sg13g2_xnor2_1 _13574_ (.Y(_06362_),
    .A(_06283_),
    .B(_06335_));
 sg13g2_xnor2_1 _13575_ (.Y(_06363_),
    .A(_06361_),
    .B(_06362_));
 sg13g2_xor2_1 _13576_ (.B(_06268_),
    .A(_06267_),
    .X(_06364_));
 sg13g2_nor2b_1 _13577_ (.A(_06363_),
    .B_N(_06364_),
    .Y(_06365_));
 sg13g2_a21o_1 _13578_ (.A2(_06362_),
    .A1(_06361_),
    .B1(_06365_),
    .X(_06366_));
 sg13g2_nor2b_1 _13579_ (.A(_06346_),
    .B_N(_06366_),
    .Y(_06367_));
 sg13g2_xnor2_1 _13580_ (.Y(_06368_),
    .A(_06363_),
    .B(_06364_));
 sg13g2_a22oi_1 _13581_ (.Y(_06369_),
    .B1(_06277_),
    .B2(\spiking_network_top_uut.all_data_out[194] ),
    .A2(_06275_),
    .A1(\spiking_network_top_uut.all_data_out[192] ));
 sg13g2_nor2_1 _13582_ (.A(_06281_),
    .B(_06369_),
    .Y(_06370_));
 sg13g2_inv_1 _13583_ (.Y(_06371_),
    .A(_06370_));
 sg13g2_xnor2_1 _13584_ (.Y(_06372_),
    .A(_06352_),
    .B(_06353_));
 sg13g2_nor2_1 _13585_ (.A(_06371_),
    .B(_06372_),
    .Y(_06373_));
 sg13g2_a21o_2 _13586_ (.A2(_06359_),
    .A1(_06357_),
    .B1(_06358_),
    .X(_06374_));
 sg13g2_nand3_1 _13587_ (.B(_06373_),
    .C(_06374_),
    .A(_06360_),
    .Y(_06375_));
 sg13g2_a21oi_1 _13588_ (.A1(_06360_),
    .A2(_06374_),
    .Y(_06376_),
    .B1(_06373_));
 sg13g2_a21o_1 _13589_ (.A2(_06374_),
    .A1(_06360_),
    .B1(_06373_),
    .X(_06377_));
 sg13g2_xnor2_1 _13590_ (.Y(_06378_),
    .A(_06264_),
    .B(_06266_));
 sg13g2_inv_1 _13591_ (.Y(_06379_),
    .A(_06378_));
 sg13g2_nand3_1 _13592_ (.B(_06377_),
    .C(_06379_),
    .A(_06375_),
    .Y(_06380_));
 sg13g2_o21ai_1 _13593_ (.B1(_06375_),
    .Y(_06381_),
    .A1(_06376_),
    .A2(_06378_));
 sg13g2_nand2_1 _13594_ (.Y(_06382_),
    .A(_06368_),
    .B(_06381_));
 sg13g2_a21o_1 _13595_ (.A2(_06377_),
    .A1(_06375_),
    .B1(_06379_),
    .X(_06383_));
 sg13g2_xnor2_1 _13596_ (.Y(_06384_),
    .A(_00058_),
    .B(_06263_));
 sg13g2_xnor2_1 _13597_ (.Y(_06385_),
    .A(_06371_),
    .B(_06372_));
 sg13g2_or2_1 _13598_ (.X(_06386_),
    .B(_06385_),
    .A(_06384_));
 sg13g2_inv_1 _13599_ (.Y(_06387_),
    .A(_06386_));
 sg13g2_nand3_1 _13600_ (.B(_06383_),
    .C(_06387_),
    .A(_06380_),
    .Y(_06388_));
 sg13g2_xnor2_1 _13601_ (.Y(_06389_),
    .A(_06368_),
    .B(_06381_));
 sg13g2_o21ai_1 _13602_ (.B1(_06382_),
    .Y(_06390_),
    .A1(_06388_),
    .A2(_06389_));
 sg13g2_nand2b_1 _13603_ (.Y(_06391_),
    .B(_06346_),
    .A_N(_06366_));
 sg13g2_nand2b_1 _13604_ (.Y(_06392_),
    .B(_06391_),
    .A_N(_06367_));
 sg13g2_nand2b_1 _13605_ (.Y(_06393_),
    .B(_06390_),
    .A_N(_06392_));
 sg13g2_a21oi_2 _13606_ (.B1(_06367_),
    .Y(_06394_),
    .A2(_06391_),
    .A1(_06390_));
 sg13g2_xor2_1 _13607_ (.B(_06344_),
    .A(_06318_),
    .X(_06395_));
 sg13g2_nor2_1 _13608_ (.A(_06394_),
    .B(_06395_),
    .Y(_06396_));
 sg13g2_o21ai_1 _13609_ (.B1(_06345_),
    .Y(_06397_),
    .A1(_06394_),
    .A2(_06395_));
 sg13g2_a21oi_1 _13610_ (.A1(_06316_),
    .A2(_06317_),
    .Y(_06398_),
    .B1(_06313_));
 sg13g2_nor2_1 _13611_ (.A(_06273_),
    .B(_06316_),
    .Y(_06399_));
 sg13g2_xnor2_1 _13612_ (.Y(_06400_),
    .A(_06273_),
    .B(_06316_));
 sg13g2_nor2_1 _13613_ (.A(_06398_),
    .B(_06400_),
    .Y(_06401_));
 sg13g2_xor2_1 _13614_ (.B(_06400_),
    .A(_06398_),
    .X(_06402_));
 sg13g2_xnor2_1 _13615_ (.Y(_06403_),
    .A(_06397_),
    .B(_06402_));
 sg13g2_mux2_1 _13616_ (.A0(_06274_),
    .A1(_06403_),
    .S(_06227_),
    .X(_06404_));
 sg13g2_nand2_1 _13617_ (.Y(_06405_),
    .A(_06394_),
    .B(_06395_));
 sg13g2_nor2_1 _13618_ (.A(_06228_),
    .B(_06396_),
    .Y(_06406_));
 sg13g2_a22oi_1 _13619_ (.Y(_06407_),
    .B1(_06405_),
    .B2(_06406_),
    .A2(_06317_),
    .A1(net3705));
 sg13g2_a21oi_1 _13620_ (.A1(_06227_),
    .A2(_06312_),
    .Y(_06408_),
    .B1(_06274_));
 sg13g2_a221oi_1 _13621_ (.B2(_06397_),
    .C1(_06401_),
    .B1(_06402_),
    .A1(_06312_),
    .Y(_06409_),
    .A2(_06399_));
 sg13g2_a21o_1 _13622_ (.A2(_06409_),
    .A1(_06227_),
    .B1(_06408_),
    .X(_06410_));
 sg13g2_o21ai_1 _13623_ (.B1(_06410_),
    .Y(_06411_),
    .A1(_06404_),
    .A2(_06407_));
 sg13g2_and2_1 _13624_ (.A(_04787_),
    .B(_06411_),
    .X(_06412_));
 sg13g2_a21oi_2 _13625_ (.B1(_06410_),
    .Y(_06413_),
    .A2(_06407_),
    .A1(_06404_));
 sg13g2_nor2_1 _13626_ (.A(net3705),
    .B(_06385_),
    .Y(_06414_));
 sg13g2_xnor2_1 _13627_ (.Y(_06415_),
    .A(_06384_),
    .B(_06414_));
 sg13g2_o21ai_1 _13628_ (.B1(_06412_),
    .Y(_06416_),
    .A1(_06413_),
    .A2(_06415_));
 sg13g2_xor2_1 _13629_ (.B(net457),
    .A(net4312),
    .X(_06417_));
 sg13g2_a21oi_1 _13630_ (.A1(net3658),
    .A2(_06417_),
    .Y(_06418_),
    .B1(net3929));
 sg13g2_a22oi_1 _13631_ (.Y(_00615_),
    .B1(_06416_),
    .B2(_06418_),
    .A2(_03444_),
    .A1(net3929));
 sg13g2_a21o_1 _13632_ (.A2(_06383_),
    .A1(_06380_),
    .B1(_06387_),
    .X(_06419_));
 sg13g2_and2_1 _13633_ (.A(_06227_),
    .B(_06388_),
    .X(_06420_));
 sg13g2_a221oi_1 _13634_ (.B2(_06420_),
    .C1(_06413_),
    .B1(_06419_),
    .A1(net3705),
    .Y(_06421_),
    .A2(_06379_));
 sg13g2_nand2_1 _13635_ (.Y(_06422_),
    .A(net4533),
    .B(_06412_));
 sg13g2_xor2_1 _13636_ (.B(_04781_),
    .A(_04780_),
    .X(_06423_));
 sg13g2_a22oi_1 _13637_ (.Y(_06424_),
    .B1(_00011_),
    .B2(_06423_),
    .A2(net517),
    .A1(net3929));
 sg13g2_o21ai_1 _13638_ (.B1(_06424_),
    .Y(_00616_),
    .A1(_06421_),
    .A2(_06422_));
 sg13g2_nand2_1 _13639_ (.Y(_06425_),
    .A(net3705),
    .B(_06364_));
 sg13g2_xnor2_1 _13640_ (.Y(_06426_),
    .A(_06388_),
    .B(_06389_));
 sg13g2_o21ai_1 _13641_ (.B1(_06425_),
    .Y(_06427_),
    .A1(net3705),
    .A2(_06426_));
 sg13g2_o21ai_1 _13642_ (.B1(_06412_),
    .Y(_06428_),
    .A1(_06413_),
    .A2(_06427_));
 sg13g2_xnor2_1 _13643_ (.Y(_06429_),
    .A(_04778_),
    .B(_04782_));
 sg13g2_a21oi_1 _13644_ (.A1(net3658),
    .A2(_06429_),
    .Y(_06430_),
    .B1(net3929));
 sg13g2_a22oi_1 _13645_ (.Y(_00617_),
    .B1(_06428_),
    .B2(_06430_),
    .A2(_03443_),
    .A1(net3929));
 sg13g2_nand2b_1 _13646_ (.Y(_06431_),
    .B(_06392_),
    .A_N(_06390_));
 sg13g2_and2_1 _13647_ (.A(_06227_),
    .B(_06393_),
    .X(_06432_));
 sg13g2_a221oi_1 _13648_ (.B2(_06432_),
    .C1(_06413_),
    .B1(_06431_),
    .A1(net3705),
    .Y(_06433_),
    .A2(_06343_));
 sg13g2_or3_1 _13649_ (.A(_04776_),
    .B(_04777_),
    .C(_04783_),
    .X(_06434_));
 sg13g2_and2_1 _13650_ (.A(_04784_),
    .B(_06434_),
    .X(_06435_));
 sg13g2_a22oi_1 _13651_ (.Y(_06436_),
    .B1(_00011_),
    .B2(_06435_),
    .A2(net540),
    .A1(net3929));
 sg13g2_o21ai_1 _13652_ (.B1(_06436_),
    .Y(_00618_),
    .A1(_06422_),
    .A2(_06433_));
 sg13g2_o21ai_1 _13653_ (.B1(net4531),
    .Y(_06437_),
    .A1(_04774_),
    .A2(_04785_));
 sg13g2_a21oi_1 _13654_ (.A1(_04787_),
    .A2(_06410_),
    .Y(_06438_),
    .B1(_06437_));
 sg13g2_a21oi_1 _13655_ (.A1(net3929),
    .A2(_03442_),
    .Y(_00619_),
    .B1(_06438_));
 sg13g2_mux4_1 _13656_ (.S0(\spiking_network_top_uut.all_data_out[700] ),
    .A0(net3846),
    .A1(net3845),
    .A2(net3844),
    .A3(net3843),
    .S1(\spiking_network_top_uut.all_data_out[701] ),
    .X(_06439_));
 sg13g2_mux2_1 _13657_ (.A0(net3841),
    .A1(net3900),
    .S(\spiking_network_top_uut.all_data_out[700] ),
    .X(_06440_));
 sg13g2_nor2b_1 _13658_ (.A(\spiking_network_top_uut.all_data_out[700] ),
    .B_N(net3842),
    .Y(_06441_));
 sg13g2_a21oi_1 _13659_ (.A1(\spiking_network_top_uut.all_data_out[700] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[5] ),
    .Y(_06442_),
    .B1(_06441_));
 sg13g2_o21ai_1 _13660_ (.B1(\spiking_network_top_uut.all_data_out[702] ),
    .Y(_06443_),
    .A1(\spiking_network_top_uut.all_data_out[701] ),
    .A2(_06442_));
 sg13g2_a21oi_1 _13661_ (.A1(\spiking_network_top_uut.all_data_out[701] ),
    .A2(_06440_),
    .Y(_06444_),
    .B1(_06443_));
 sg13g2_o21ai_1 _13662_ (.B1(net4550),
    .Y(_06445_),
    .A1(\spiking_network_top_uut.all_data_out[702] ),
    .A2(_06439_));
 sg13g2_nand2_1 _13663_ (.Y(_06446_),
    .A(net3934),
    .B(net349));
 sg13g2_o21ai_1 _13664_ (.B1(_06446_),
    .Y(_00620_),
    .A1(_06444_),
    .A2(_06445_));
 sg13g2_mux2_1 _13665_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_dout ),
    .A1(net349),
    .S(net4550),
    .X(_00621_));
 sg13g2_mux4_1 _13666_ (.S0(\spiking_network_top_uut.all_data_out[696] ),
    .A0(net3898),
    .A1(net3897),
    .A2(net3896),
    .A3(net3895),
    .S1(\spiking_network_top_uut.all_data_out[697] ),
    .X(_06447_));
 sg13g2_mux2_1 _13667_ (.A0(net3893),
    .A1(net3892),
    .S(\spiking_network_top_uut.all_data_out[696] ),
    .X(_06448_));
 sg13g2_nor2b_1 _13668_ (.A(\spiking_network_top_uut.all_data_out[696] ),
    .B_N(net3894),
    .Y(_06449_));
 sg13g2_a21oi_1 _13669_ (.A1(\spiking_network_top_uut.all_data_out[696] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[5] ),
    .Y(_06450_),
    .B1(_06449_));
 sg13g2_o21ai_1 _13670_ (.B1(\spiking_network_top_uut.all_data_out[698] ),
    .Y(_06451_),
    .A1(\spiking_network_top_uut.all_data_out[697] ),
    .A2(_06450_));
 sg13g2_a21oi_1 _13671_ (.A1(\spiking_network_top_uut.all_data_out[697] ),
    .A2(_06448_),
    .Y(_06452_),
    .B1(_06451_));
 sg13g2_o21ai_1 _13672_ (.B1(net4546),
    .Y(_06453_),
    .A1(\spiking_network_top_uut.all_data_out[698] ),
    .A2(_06447_));
 sg13g2_nand2_1 _13673_ (.Y(_06454_),
    .A(net3934),
    .B(net62));
 sg13g2_o21ai_1 _13674_ (.B1(_06454_),
    .Y(_00622_),
    .A1(_06452_),
    .A2(_06453_));
 sg13g2_mux2_1 _13675_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_dout ),
    .A1(net62),
    .S(net4549),
    .X(_00623_));
 sg13g2_mux4_1 _13676_ (.S0(\spiking_network_top_uut.all_data_out[692] ),
    .A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[0] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[1] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[2] ),
    .A3(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[3] ),
    .S1(\spiking_network_top_uut.all_data_out[693] ),
    .X(_06455_));
 sg13g2_mux2_1 _13677_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[6] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[7] ),
    .S(\spiking_network_top_uut.all_data_out[692] ),
    .X(_06456_));
 sg13g2_nor2b_1 _13678_ (.A(\spiking_network_top_uut.all_data_out[692] ),
    .B_N(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[4] ),
    .Y(_06457_));
 sg13g2_a21oi_1 _13679_ (.A1(\spiking_network_top_uut.all_data_out[692] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[5] ),
    .Y(_06458_),
    .B1(_06457_));
 sg13g2_o21ai_1 _13680_ (.B1(\spiking_network_top_uut.all_data_out[694] ),
    .Y(_06459_),
    .A1(\spiking_network_top_uut.all_data_out[693] ),
    .A2(_06458_));
 sg13g2_a21oi_1 _13681_ (.A1(\spiking_network_top_uut.all_data_out[693] ),
    .A2(_06456_),
    .Y(_06460_),
    .B1(_06459_));
 sg13g2_o21ai_1 _13682_ (.B1(net4561),
    .Y(_06461_),
    .A1(\spiking_network_top_uut.all_data_out[694] ),
    .A2(_06455_));
 sg13g2_nand2_1 _13683_ (.Y(_06462_),
    .A(net3935),
    .B(net81));
 sg13g2_o21ai_1 _13684_ (.B1(_06462_),
    .Y(_00624_),
    .A1(_06460_),
    .A2(_06461_));
 sg13g2_mux2_1 _13685_ (.A0(net264),
    .A1(net81),
    .S(net4561),
    .X(_00625_));
 sg13g2_mux4_1 _13686_ (.S0(\spiking_network_top_uut.all_data_out[688] ),
    .A0(net3884),
    .A1(net3883),
    .A2(net3882),
    .A3(net3881),
    .S1(\spiking_network_top_uut.all_data_out[689] ),
    .X(_06463_));
 sg13g2_mux2_1 _13687_ (.A0(net3878),
    .A1(net3877),
    .S(\spiking_network_top_uut.all_data_out[688] ),
    .X(_06464_));
 sg13g2_nor2b_1 _13688_ (.A(\spiking_network_top_uut.all_data_out[688] ),
    .B_N(net3880),
    .Y(_06465_));
 sg13g2_a21oi_1 _13689_ (.A1(\spiking_network_top_uut.all_data_out[688] ),
    .A2(net3879),
    .Y(_06466_),
    .B1(_06465_));
 sg13g2_o21ai_1 _13690_ (.B1(\spiking_network_top_uut.all_data_out[690] ),
    .Y(_06467_),
    .A1(\spiking_network_top_uut.all_data_out[689] ),
    .A2(_06466_));
 sg13g2_a21oi_1 _13691_ (.A1(\spiking_network_top_uut.all_data_out[689] ),
    .A2(_06464_),
    .Y(_06468_),
    .B1(_06467_));
 sg13g2_o21ai_1 _13692_ (.B1(net4557),
    .Y(_06469_),
    .A1(\spiking_network_top_uut.all_data_out[690] ),
    .A2(_06463_));
 sg13g2_nand2_1 _13693_ (.Y(_06470_),
    .A(net3938),
    .B(net130));
 sg13g2_o21ai_1 _13694_ (.B1(_06470_),
    .Y(_00626_),
    .A1(_06468_),
    .A2(_06469_));
 sg13g2_mux2_1 _13695_ (.A0(net261),
    .A1(net130),
    .S(net4557),
    .X(_00627_));
 sg13g2_mux4_1 _13696_ (.S0(\spiking_network_top_uut.all_data_out[684] ),
    .A0(net3876),
    .A1(net3875),
    .A2(net3874),
    .A3(net3873),
    .S1(\spiking_network_top_uut.all_data_out[685] ),
    .X(_06471_));
 sg13g2_mux2_1 _13697_ (.A0(net3870),
    .A1(net3869),
    .S(\spiking_network_top_uut.all_data_out[684] ),
    .X(_06472_));
 sg13g2_nor2b_1 _13698_ (.A(\spiking_network_top_uut.all_data_out[684] ),
    .B_N(net3872),
    .Y(_06473_));
 sg13g2_a21oi_1 _13699_ (.A1(\spiking_network_top_uut.all_data_out[684] ),
    .A2(net3871),
    .Y(_06474_),
    .B1(_06473_));
 sg13g2_o21ai_1 _13700_ (.B1(\spiking_network_top_uut.all_data_out[686] ),
    .Y(_06475_),
    .A1(\spiking_network_top_uut.all_data_out[685] ),
    .A2(_06474_));
 sg13g2_a21oi_1 _13701_ (.A1(\spiking_network_top_uut.all_data_out[685] ),
    .A2(_06472_),
    .Y(_06476_),
    .B1(_06475_));
 sg13g2_o21ai_1 _13702_ (.B1(net4566),
    .Y(_06477_),
    .A1(\spiking_network_top_uut.all_data_out[686] ),
    .A2(_06471_));
 sg13g2_nand2_1 _13703_ (.Y(_06478_),
    .A(net3937),
    .B(net36));
 sg13g2_o21ai_1 _13704_ (.B1(_06478_),
    .Y(_00628_),
    .A1(_06476_),
    .A2(_06477_));
 sg13g2_mux2_1 _13705_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_dout ),
    .A1(net36),
    .S(net4566),
    .X(_00629_));
 sg13g2_nand2b_1 _13706_ (.Y(_06479_),
    .B(\spiking_network_top_uut.all_data_out[680] ),
    .A_N(net3863));
 sg13g2_nor2_1 _13707_ (.A(\spiking_network_top_uut.all_data_out[680] ),
    .B(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[4] ),
    .Y(_06480_));
 sg13g2_nor2_1 _13708_ (.A(\spiking_network_top_uut.all_data_out[681] ),
    .B(_06480_),
    .Y(_06481_));
 sg13g2_mux2_1 _13709_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[6] ),
    .A1(net3861),
    .S(\spiking_network_top_uut.all_data_out[680] ),
    .X(_06482_));
 sg13g2_a221oi_1 _13710_ (.B2(\spiking_network_top_uut.all_data_out[681] ),
    .C1(_03596_),
    .B1(_06482_),
    .A1(_06479_),
    .Y(_06483_),
    .A2(_06481_));
 sg13g2_mux4_1 _13711_ (.S0(\spiking_network_top_uut.all_data_out[680] ),
    .A0(net3868),
    .A1(net3867),
    .A2(net3866),
    .A3(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[3] ),
    .S1(\spiking_network_top_uut.all_data_out[681] ),
    .X(_06484_));
 sg13g2_o21ai_1 _13712_ (.B1(net4563),
    .Y(_06485_),
    .A1(\spiking_network_top_uut.all_data_out[682] ),
    .A2(_06484_));
 sg13g2_nand2_1 _13713_ (.Y(_06486_),
    .A(net3936),
    .B(net224));
 sg13g2_o21ai_1 _13714_ (.B1(_06486_),
    .Y(_00630_),
    .A1(_06483_),
    .A2(_06485_));
 sg13g2_mux2_1 _13715_ (.A0(net309),
    .A1(net224),
    .S(net4564),
    .X(_00631_));
 sg13g2_a21oi_1 _13716_ (.A1(\spiking_network_top_uut.all_data_out[676] ),
    .A2(_03664_),
    .Y(_06487_),
    .B1(\spiking_network_top_uut.all_data_out[677] ));
 sg13g2_o21ai_1 _13717_ (.B1(_06487_),
    .Y(_06488_),
    .A1(\spiking_network_top_uut.all_data_out[676] ),
    .A2(net3856));
 sg13g2_mux2_1 _13718_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[6] ),
    .A1(net3854),
    .S(\spiking_network_top_uut.all_data_out[676] ),
    .X(_06489_));
 sg13g2_nand2_1 _13719_ (.Y(_06490_),
    .A(\spiking_network_top_uut.all_data_out[677] ),
    .B(_06489_));
 sg13g2_nand3_1 _13720_ (.B(_06488_),
    .C(_06490_),
    .A(\spiking_network_top_uut.all_data_out[678] ),
    .Y(_06491_));
 sg13g2_mux2_1 _13721_ (.A0(net3858),
    .A1(net3857),
    .S(\spiking_network_top_uut.all_data_out[676] ),
    .X(_06492_));
 sg13g2_nor2b_1 _13722_ (.A(\spiking_network_top_uut.all_data_out[676] ),
    .B_N(net3860),
    .Y(_06493_));
 sg13g2_a21oi_1 _13723_ (.A1(\spiking_network_top_uut.all_data_out[676] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[1] ),
    .Y(_06494_),
    .B1(_06493_));
 sg13g2_a21oi_1 _13724_ (.A1(\spiking_network_top_uut.all_data_out[677] ),
    .A2(_06492_),
    .Y(_06495_),
    .B1(\spiking_network_top_uut.all_data_out[678] ));
 sg13g2_o21ai_1 _13725_ (.B1(_06495_),
    .Y(_06496_),
    .A1(\spiking_network_top_uut.all_data_out[677] ),
    .A2(_06494_));
 sg13g2_nand3_1 _13726_ (.B(_06491_),
    .C(_06496_),
    .A(net4540),
    .Y(_06497_));
 sg13g2_o21ai_1 _13727_ (.B1(_06497_),
    .Y(_00632_),
    .A1(net4540),
    .A2(_03674_));
 sg13g2_nor2_1 _13728_ (.A(net4540),
    .B(net146),
    .Y(_06498_));
 sg13g2_a21oi_1 _13729_ (.A1(net4540),
    .A2(_03674_),
    .Y(_00633_),
    .B1(_06498_));
 sg13g2_a21oi_1 _13730_ (.A1(\spiking_network_top_uut.all_data_out[672] ),
    .A2(_03663_),
    .Y(_06499_),
    .B1(\spiking_network_top_uut.all_data_out[673] ));
 sg13g2_o21ai_1 _13731_ (.B1(_06499_),
    .Y(_06500_),
    .A1(\spiking_network_top_uut.all_data_out[672] ),
    .A2(net3849));
 sg13g2_mux2_1 _13732_ (.A0(net3848),
    .A1(net3847),
    .S(\spiking_network_top_uut.all_data_out[672] ),
    .X(_06501_));
 sg13g2_nand2_1 _13733_ (.Y(_06502_),
    .A(\spiking_network_top_uut.all_data_out[673] ),
    .B(_06501_));
 sg13g2_nand3_1 _13734_ (.B(_06500_),
    .C(_06502_),
    .A(\spiking_network_top_uut.all_data_out[674] ),
    .Y(_06503_));
 sg13g2_mux2_1 _13735_ (.A0(net3851),
    .A1(net3850),
    .S(\spiking_network_top_uut.all_data_out[672] ),
    .X(_06504_));
 sg13g2_nor2b_1 _13736_ (.A(\spiking_network_top_uut.all_data_out[672] ),
    .B_N(net3853),
    .Y(_06505_));
 sg13g2_a21oi_1 _13737_ (.A1(\spiking_network_top_uut.all_data_out[672] ),
    .A2(net3852),
    .Y(_06506_),
    .B1(_06505_));
 sg13g2_a21oi_1 _13738_ (.A1(\spiking_network_top_uut.all_data_out[673] ),
    .A2(_06504_),
    .Y(_06507_),
    .B1(\spiking_network_top_uut.all_data_out[674] ));
 sg13g2_o21ai_1 _13739_ (.B1(_06507_),
    .Y(_06508_),
    .A1(\spiking_network_top_uut.all_data_out[673] ),
    .A2(_06506_));
 sg13g2_nand3_1 _13740_ (.B(_06503_),
    .C(_06508_),
    .A(net4544),
    .Y(_06509_));
 sg13g2_o21ai_1 _13741_ (.B1(_06509_),
    .Y(_00634_),
    .A1(net4539),
    .A2(_03675_));
 sg13g2_nor3_2 _13742_ (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[2] ),
    .B(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[1] ),
    .C(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[0] ),
    .Y(_06510_));
 sg13g2_nor2b_1 _13743_ (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[3] ),
    .B_N(_06510_),
    .Y(_06511_));
 sg13g2_nor2b_2 _13744_ (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[4] ),
    .B_N(_06511_),
    .Y(_06512_));
 sg13g2_nand2b_2 _13745_ (.Y(_06513_),
    .B(_06511_),
    .A_N(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[4] ));
 sg13g2_o21ai_1 _13746_ (.B1(net4529),
    .Y(_06514_),
    .A1(net3654),
    .A2(_06513_));
 sg13g2_nor2b_1 _13747_ (.A(net3653),
    .B_N(net333),
    .Y(_06515_));
 sg13g2_a21oi_1 _13748_ (.A1(net4283),
    .A2(net3653),
    .Y(_06516_),
    .B1(_06515_));
 sg13g2_nand2_1 _13749_ (.Y(_06517_),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[0] ),
    .B(_06514_));
 sg13g2_o21ai_1 _13750_ (.B1(_06517_),
    .Y(_00635_),
    .A1(_06514_),
    .A2(_06516_));
 sg13g2_xor2_1 _13751_ (.B(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[0] ),
    .A(net343),
    .X(_06518_));
 sg13g2_nor2_1 _13752_ (.A(net3653),
    .B(_06518_),
    .Y(_06519_));
 sg13g2_a21oi_1 _13753_ (.A1(net4280),
    .A2(net3653),
    .Y(_06520_),
    .B1(_06519_));
 sg13g2_nand2_1 _13754_ (.Y(_06521_),
    .A(net343),
    .B(_06514_));
 sg13g2_o21ai_1 _13755_ (.B1(_06521_),
    .Y(_00636_),
    .A1(_06514_),
    .A2(_06520_));
 sg13g2_o21ai_1 _13756_ (.B1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[2] ),
    .Y(_06522_),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[1] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[0] ));
 sg13g2_nor2b_1 _13757_ (.A(_06510_),
    .B_N(_06522_),
    .Y(_06523_));
 sg13g2_nor2_1 _13758_ (.A(net3653),
    .B(_06523_),
    .Y(_06524_));
 sg13g2_a21oi_1 _13759_ (.A1(net4276),
    .A2(net3653),
    .Y(_06525_),
    .B1(_06524_));
 sg13g2_nand2_1 _13760_ (.Y(_06526_),
    .A(net208),
    .B(_06514_));
 sg13g2_o21ai_1 _13761_ (.B1(_06526_),
    .Y(_00637_),
    .A1(_06514_),
    .A2(_06525_));
 sg13g2_nand2_1 _13762_ (.Y(_06527_),
    .A(net4273),
    .B(net3653));
 sg13g2_xnor2_1 _13763_ (.Y(_06528_),
    .A(net406),
    .B(_06510_));
 sg13g2_o21ai_1 _13764_ (.B1(_06527_),
    .Y(_06529_),
    .A1(net3653),
    .A2(_06528_));
 sg13g2_mux2_1 _13765_ (.A0(_06529_),
    .A1(net406),
    .S(_06514_),
    .X(_00638_));
 sg13g2_nand2_1 _13766_ (.Y(_06530_),
    .A(net3922),
    .B(net367));
 sg13g2_nand2b_1 _13767_ (.Y(_06531_),
    .B(net367),
    .A_N(_06511_));
 sg13g2_a21oi_1 _13768_ (.A1(_06513_),
    .A2(_06531_),
    .Y(_06532_),
    .B1(net3654));
 sg13g2_a21oi_1 _13769_ (.A1(net4269),
    .A2(net3654),
    .Y(_06533_),
    .B1(_06532_));
 sg13g2_o21ai_1 _13770_ (.B1(_06530_),
    .Y(_00639_),
    .A1(_06514_),
    .A2(_06533_));
 sg13g2_nor2_1 _13771_ (.A(net4541),
    .B(net269),
    .Y(_06534_));
 sg13g2_a21oi_1 _13772_ (.A1(net4541),
    .A2(_03675_),
    .Y(_00640_),
    .B1(_06534_));
 sg13g2_nor2_1 _13773_ (.A(_00061_),
    .B(net3740),
    .Y(_06535_));
 sg13g2_nor2_2 _13774_ (.A(net3742),
    .B(_06535_),
    .Y(_06536_));
 sg13g2_nand2b_1 _13775_ (.Y(_06537_),
    .B(_06536_),
    .A_N(_00061_));
 sg13g2_o21ai_1 _13776_ (.B1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ),
    .Y(_06538_),
    .A1(_00061_),
    .A2(_06536_));
 sg13g2_a21o_1 _13777_ (.A2(net3742),
    .A1(_00062_),
    .B1(_06536_),
    .X(_06539_));
 sg13g2_nand2_1 _13778_ (.Y(_06540_),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ),
    .B(_06539_));
 sg13g2_nand2_1 _13779_ (.Y(_06541_),
    .A(_00063_),
    .B(net3742));
 sg13g2_o21ai_1 _13780_ (.B1(net3916),
    .Y(_06542_),
    .A1(_00062_),
    .A2(net3903));
 sg13g2_a21o_1 _13781_ (.A2(_06535_),
    .A1(net3903),
    .B1(_06542_),
    .X(_06543_));
 sg13g2_a21oi_1 _13782_ (.A1(_06541_),
    .A2(_06543_),
    .Y(_06544_),
    .B1(_03448_));
 sg13g2_nor2_1 _13783_ (.A(_00065_),
    .B(net3916),
    .Y(_06545_));
 sg13g2_o21ai_1 _13784_ (.B1(net3913),
    .Y(_06546_),
    .A1(_00061_),
    .A2(net3909));
 sg13g2_a22oi_1 _13785_ (.Y(_06547_),
    .B1(net3901),
    .B2(_00062_),
    .A2(net3738),
    .A1(_00063_));
 sg13g2_and3_1 _13786_ (.X(_06548_),
    .A(net3916),
    .B(_06546_),
    .C(_06547_));
 sg13g2_o21ai_1 _13787_ (.B1(_00064_),
    .Y(_06549_),
    .A1(_06545_),
    .A2(_06548_));
 sg13g2_inv_1 _13788_ (.Y(_06550_),
    .A(_06549_));
 sg13g2_nand3_1 _13789_ (.B(_06541_),
    .C(_06543_),
    .A(_03448_),
    .Y(_06551_));
 sg13g2_nand2b_1 _13790_ (.Y(_06552_),
    .B(_06551_),
    .A_N(_06544_));
 sg13g2_a21oi_1 _13791_ (.A1(_06549_),
    .A2(_06551_),
    .Y(_06553_),
    .B1(_06544_));
 sg13g2_xor2_1 _13792_ (.B(_06539_),
    .A(_00063_),
    .X(_06554_));
 sg13g2_o21ai_1 _13793_ (.B1(_06540_),
    .Y(_06555_),
    .A1(_06553_),
    .A2(_06554_));
 sg13g2_or3_1 _13794_ (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ),
    .B(_00061_),
    .C(_06536_),
    .X(_06556_));
 sg13g2_and2_1 _13795_ (.A(_06538_),
    .B(_06556_),
    .X(_06557_));
 sg13g2_nand2_1 _13796_ (.Y(_06558_),
    .A(_06555_),
    .B(_06557_));
 sg13g2_and2_1 _13797_ (.A(_06538_),
    .B(_06558_),
    .X(_06559_));
 sg13g2_a22oi_1 _13798_ (.Y(_06560_),
    .B1(_06537_),
    .B2(_06559_),
    .A2(_06536_),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ));
 sg13g2_a21o_1 _13799_ (.A2(_00061_),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ),
    .B1(_06560_),
    .X(_06561_));
 sg13g2_mux2_1 _13800_ (.A0(net4599),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[675] ),
    .X(_06562_));
 sg13g2_nand2_1 _13801_ (.Y(_06563_),
    .A(\spiking_network_top_uut.all_data_out[209] ),
    .B(_06562_));
 sg13g2_mux2_1 _13802_ (.A0(net4598),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[679] ),
    .X(_06564_));
 sg13g2_nand2_1 _13803_ (.Y(_06565_),
    .A(\spiking_network_top_uut.all_data_out[211] ),
    .B(_06564_));
 sg13g2_nor2_1 _13804_ (.A(_06563_),
    .B(_06565_),
    .Y(_06566_));
 sg13g2_nand4_1 _13805_ (.B(\spiking_network_top_uut.all_data_out[210] ),
    .C(_06562_),
    .A(\spiking_network_top_uut.all_data_out[208] ),
    .Y(_06567_),
    .D(_06564_));
 sg13g2_inv_1 _13806_ (.Y(_06568_),
    .A(_06567_));
 sg13g2_xor2_1 _13807_ (.B(_06565_),
    .A(_06563_),
    .X(_06569_));
 sg13g2_a21oi_2 _13808_ (.B1(_06566_),
    .Y(_06570_),
    .A2(_06569_),
    .A1(_06567_));
 sg13g2_mux2_2 _13809_ (.A0(net4597),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[683] ),
    .X(_06571_));
 sg13g2_nand2_1 _13810_ (.Y(_06572_),
    .A(\spiking_network_top_uut.all_data_out[213] ),
    .B(_06571_));
 sg13g2_mux2_2 _13811_ (.A0(net4596),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[687] ),
    .X(_06573_));
 sg13g2_nand2_2 _13812_ (.Y(_06574_),
    .A(\spiking_network_top_uut.all_data_out[215] ),
    .B(_06573_));
 sg13g2_nor2_1 _13813_ (.A(_06572_),
    .B(_06574_),
    .Y(_06575_));
 sg13g2_nand2_1 _13814_ (.Y(_06576_),
    .A(\spiking_network_top_uut.all_data_out[212] ),
    .B(_06571_));
 sg13g2_nand2_2 _13815_ (.Y(_06577_),
    .A(\spiking_network_top_uut.all_data_out[214] ),
    .B(_06573_));
 sg13g2_or2_1 _13816_ (.X(_06578_),
    .B(_06577_),
    .A(_06576_));
 sg13g2_xor2_1 _13817_ (.B(_06574_),
    .A(_06572_),
    .X(_06579_));
 sg13g2_a21oi_2 _13818_ (.B1(_06575_),
    .Y(_06580_),
    .A2(_06579_),
    .A1(_06578_));
 sg13g2_mux2_2 _13819_ (.A0(net4595),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[691] ),
    .X(_06581_));
 sg13g2_mux2_2 _13820_ (.A0(net4594),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[695] ),
    .X(_06582_));
 sg13g2_a22oi_1 _13821_ (.Y(_06583_),
    .B1(_06582_),
    .B2(\spiking_network_top_uut.all_data_out[219] ),
    .A2(_06581_),
    .A1(\spiking_network_top_uut.all_data_out[217] ));
 sg13g2_and4_1 _13822_ (.A(\spiking_network_top_uut.all_data_out[217] ),
    .B(\spiking_network_top_uut.all_data_out[219] ),
    .C(_06581_),
    .D(_06582_),
    .X(_06584_));
 sg13g2_nand4_1 _13823_ (.B(\spiking_network_top_uut.all_data_out[219] ),
    .C(_06581_),
    .A(\spiking_network_top_uut.all_data_out[217] ),
    .Y(_06585_),
    .D(_06582_));
 sg13g2_and4_2 _13824_ (.A(\spiking_network_top_uut.all_data_out[216] ),
    .B(\spiking_network_top_uut.all_data_out[218] ),
    .C(_06581_),
    .D(_06582_),
    .X(_06586_));
 sg13g2_nand4_1 _13825_ (.B(\spiking_network_top_uut.all_data_out[218] ),
    .C(_06581_),
    .A(\spiking_network_top_uut.all_data_out[216] ),
    .Y(_06587_),
    .D(_06582_));
 sg13g2_nand3b_1 _13826_ (.B(_06585_),
    .C(_06586_),
    .Y(_06588_),
    .A_N(_06583_));
 sg13g2_a21oi_2 _13827_ (.B1(_06583_),
    .Y(_06589_),
    .A2(_06586_),
    .A1(_06585_));
 sg13g2_mux2_2 _13828_ (.A0(net4593),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[699] ),
    .X(_06590_));
 sg13g2_mux2_2 _13829_ (.A0(net4592),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[703] ),
    .X(_06591_));
 sg13g2_and4_1 _13830_ (.A(\spiking_network_top_uut.all_data_out[221] ),
    .B(\spiking_network_top_uut.all_data_out[223] ),
    .C(_06590_),
    .D(_06591_),
    .X(_06592_));
 sg13g2_nand4_1 _13831_ (.B(\spiking_network_top_uut.all_data_out[223] ),
    .C(_06590_),
    .A(\spiking_network_top_uut.all_data_out[221] ),
    .Y(_06593_),
    .D(_06591_));
 sg13g2_and4_1 _13832_ (.A(\spiking_network_top_uut.all_data_out[220] ),
    .B(\spiking_network_top_uut.all_data_out[222] ),
    .C(_06590_),
    .D(_06591_),
    .X(_06594_));
 sg13g2_a22oi_1 _13833_ (.Y(_06595_),
    .B1(_06591_),
    .B2(\spiking_network_top_uut.all_data_out[223] ),
    .A2(_06590_),
    .A1(\spiking_network_top_uut.all_data_out[221] ));
 sg13g2_or3_2 _13834_ (.A(_06592_),
    .B(_06594_),
    .C(_06595_),
    .X(_06596_));
 sg13g2_o21ai_1 _13835_ (.B1(_06593_),
    .Y(_06597_),
    .A1(_06594_),
    .A2(_06595_));
 sg13g2_nand3b_1 _13836_ (.B(_06589_),
    .C(_06597_),
    .Y(_06598_),
    .A_N(_06580_));
 sg13g2_inv_1 _13837_ (.Y(_06599_),
    .A(_06598_));
 sg13g2_or2_1 _13838_ (.X(_06600_),
    .B(_06598_),
    .A(_06570_));
 sg13g2_inv_1 _13839_ (.Y(_06601_),
    .A(_06600_));
 sg13g2_a21oi_1 _13840_ (.A1(_06512_),
    .A2(_06600_),
    .Y(_06602_),
    .B1(_06561_));
 sg13g2_nor2_1 _13841_ (.A(_06589_),
    .B(_06597_),
    .Y(_06603_));
 sg13g2_and2_2 _13842_ (.A(_06580_),
    .B(_06603_),
    .X(_06604_));
 sg13g2_a21oi_2 _13843_ (.B1(_06601_),
    .Y(_06605_),
    .A2(_06604_),
    .A1(_06570_));
 sg13g2_inv_1 _13844_ (.Y(_06606_),
    .A(_06605_));
 sg13g2_and2_1 _13845_ (.A(_06561_),
    .B(_06606_),
    .X(_06607_));
 sg13g2_xnor2_1 _13846_ (.Y(_06608_),
    .A(_06537_),
    .B(_06559_));
 sg13g2_a21oi_1 _13847_ (.A1(_06605_),
    .A2(_06608_),
    .Y(_06609_),
    .B1(_06601_));
 sg13g2_xnor2_1 _13848_ (.Y(_06610_),
    .A(_06561_),
    .B(_06605_));
 sg13g2_nor2b_1 _13849_ (.A(_06609_),
    .B_N(_06610_),
    .Y(_06611_));
 sg13g2_xnor2_1 _13850_ (.Y(_06612_),
    .A(_06606_),
    .B(_06608_));
 sg13g2_o21ai_1 _13851_ (.B1(_06594_),
    .Y(_06613_),
    .A1(_06592_),
    .A2(_06595_));
 sg13g2_o21ai_1 _13852_ (.B1(_06587_),
    .Y(_06614_),
    .A1(_06583_),
    .A2(_06584_));
 sg13g2_o21ai_1 _13853_ (.B1(_06586_),
    .Y(_06615_),
    .A1(_06583_),
    .A2(_06584_));
 sg13g2_nand3b_1 _13854_ (.B(_06585_),
    .C(_06587_),
    .Y(_06616_),
    .A_N(_06583_));
 sg13g2_a22oi_1 _13855_ (.Y(_06617_),
    .B1(_06615_),
    .B2(_06616_),
    .A2(_06613_),
    .A1(_06596_));
 sg13g2_xor2_1 _13856_ (.B(_06579_),
    .A(_06578_),
    .X(_06618_));
 sg13g2_xnor2_1 _13857_ (.Y(_06619_),
    .A(_06578_),
    .B(_06579_));
 sg13g2_and4_1 _13858_ (.A(_06596_),
    .B(_06613_),
    .C(_06615_),
    .D(_06616_),
    .X(_06620_));
 sg13g2_nand4_1 _13859_ (.B(_06613_),
    .C(_06615_),
    .A(_06596_),
    .Y(_06621_),
    .D(_06616_));
 sg13g2_and4_1 _13860_ (.A(_06588_),
    .B(_06596_),
    .C(_06613_),
    .D(_06614_),
    .X(_06622_));
 sg13g2_a22oi_1 _13861_ (.Y(_06623_),
    .B1(_06614_),
    .B2(_06588_),
    .A2(_06613_),
    .A1(_06596_));
 sg13g2_nor3_2 _13862_ (.A(_06617_),
    .B(_06618_),
    .C(_06620_),
    .Y(_06624_));
 sg13g2_a21oi_2 _13863_ (.B1(_06617_),
    .Y(_06625_),
    .A2(_06621_),
    .A1(_06619_));
 sg13g2_xor2_1 _13864_ (.B(_06597_),
    .A(_06589_),
    .X(_06626_));
 sg13g2_xnor2_1 _13865_ (.Y(_06627_),
    .A(_06580_),
    .B(_06626_));
 sg13g2_nand2b_1 _13866_ (.Y(_06628_),
    .B(_06627_),
    .A_N(_06625_));
 sg13g2_xnor2_1 _13867_ (.Y(_06629_),
    .A(_06625_),
    .B(_06627_));
 sg13g2_nand2b_1 _13868_ (.Y(_06630_),
    .B(_06629_),
    .A_N(_06570_));
 sg13g2_nand2_1 _13869_ (.Y(_06631_),
    .A(_06628_),
    .B(_06630_));
 sg13g2_nor2_1 _13870_ (.A(_06599_),
    .B(_06604_),
    .Y(_06632_));
 sg13g2_xnor2_1 _13871_ (.Y(_06633_),
    .A(_06570_),
    .B(_06632_));
 sg13g2_and2_1 _13872_ (.A(_06631_),
    .B(_06633_),
    .X(_06634_));
 sg13g2_xor2_1 _13873_ (.B(_06633_),
    .A(_06631_),
    .X(_06635_));
 sg13g2_xnor2_1 _13874_ (.Y(_06636_),
    .A(_06555_),
    .B(_06557_));
 sg13g2_inv_1 _13875_ (.Y(_06637_),
    .A(_06636_));
 sg13g2_a21oi_1 _13876_ (.A1(_06635_),
    .A2(_06637_),
    .Y(_06638_),
    .B1(_06634_));
 sg13g2_nand2b_1 _13877_ (.Y(_06639_),
    .B(_06612_),
    .A_N(_06638_));
 sg13g2_xnor2_1 _13878_ (.Y(_06640_),
    .A(_06635_),
    .B(_06637_));
 sg13g2_a22oi_1 _13879_ (.Y(_06641_),
    .B1(_06591_),
    .B2(\spiking_network_top_uut.all_data_out[222] ),
    .A2(_06590_),
    .A1(\spiking_network_top_uut.all_data_out[220] ));
 sg13g2_nor2_1 _13880_ (.A(_06594_),
    .B(_06641_),
    .Y(_06642_));
 sg13g2_a22oi_1 _13881_ (.Y(_06643_),
    .B1(_06582_),
    .B2(\spiking_network_top_uut.all_data_out[218] ),
    .A2(_06581_),
    .A1(\spiking_network_top_uut.all_data_out[216] ));
 sg13g2_nor2_1 _13882_ (.A(_06586_),
    .B(_06643_),
    .Y(_06644_));
 sg13g2_and2_1 _13883_ (.A(_06642_),
    .B(_06644_),
    .X(_06645_));
 sg13g2_xor2_1 _13884_ (.B(_06577_),
    .A(_06576_),
    .X(_06646_));
 sg13g2_xor2_1 _13885_ (.B(_06644_),
    .A(_06642_),
    .X(_06647_));
 sg13g2_a21oi_2 _13886_ (.B1(_06645_),
    .Y(_06648_),
    .A2(_06647_),
    .A1(_06646_));
 sg13g2_nor3_2 _13887_ (.A(_06619_),
    .B(_06622_),
    .C(_06623_),
    .Y(_06649_));
 sg13g2_nor3_1 _13888_ (.A(_06624_),
    .B(_06648_),
    .C(_06649_),
    .Y(_06650_));
 sg13g2_or3_1 _13889_ (.A(_06624_),
    .B(_06648_),
    .C(_06649_),
    .X(_06651_));
 sg13g2_xnor2_1 _13890_ (.Y(_06652_),
    .A(_06567_),
    .B(_06569_));
 sg13g2_o21ai_1 _13891_ (.B1(_06648_),
    .Y(_06653_),
    .A1(_06624_),
    .A2(_06649_));
 sg13g2_nand3_1 _13892_ (.B(_06652_),
    .C(_06653_),
    .A(_06651_),
    .Y(_06654_));
 sg13g2_a21o_2 _13893_ (.A2(_06653_),
    .A1(_06652_),
    .B1(_06650_),
    .X(_06655_));
 sg13g2_xnor2_1 _13894_ (.Y(_06656_),
    .A(_06570_),
    .B(_06629_));
 sg13g2_nand2_1 _13895_ (.Y(_06657_),
    .A(_06655_),
    .B(_06656_));
 sg13g2_xnor2_1 _13896_ (.Y(_06658_),
    .A(_06655_),
    .B(_06656_));
 sg13g2_xnor2_1 _13897_ (.Y(_06659_),
    .A(_06553_),
    .B(_06554_));
 sg13g2_o21ai_1 _13898_ (.B1(_06657_),
    .Y(_06660_),
    .A1(_06658_),
    .A2(_06659_));
 sg13g2_nor2b_1 _13899_ (.A(_06640_),
    .B_N(_06660_),
    .Y(_06661_));
 sg13g2_xor2_1 _13900_ (.B(_06659_),
    .A(_06658_),
    .X(_06662_));
 sg13g2_a22oi_1 _13901_ (.Y(_06663_),
    .B1(_06564_),
    .B2(\spiking_network_top_uut.all_data_out[210] ),
    .A2(_06562_),
    .A1(\spiking_network_top_uut.all_data_out[208] ));
 sg13g2_xnor2_1 _13902_ (.Y(_06664_),
    .A(_06646_),
    .B(_06647_));
 sg13g2_nor3_2 _13903_ (.A(_06568_),
    .B(_06663_),
    .C(_06664_),
    .Y(_06665_));
 sg13g2_a21o_2 _13904_ (.A2(_06653_),
    .A1(_06651_),
    .B1(_06652_),
    .X(_06666_));
 sg13g2_and3_1 _13905_ (.X(_06667_),
    .A(_06654_),
    .B(_06665_),
    .C(_06666_));
 sg13g2_nand3_1 _13906_ (.B(_06665_),
    .C(_06666_),
    .A(_06654_),
    .Y(_06668_));
 sg13g2_a21oi_1 _13907_ (.A1(_06654_),
    .A2(_06666_),
    .Y(_06669_),
    .B1(_06665_));
 sg13g2_xnor2_1 _13908_ (.Y(_06670_),
    .A(_06550_),
    .B(_06552_));
 sg13g2_nor3_1 _13909_ (.A(_06667_),
    .B(_06669_),
    .C(_06670_),
    .Y(_06671_));
 sg13g2_o21ai_1 _13910_ (.B1(_06668_),
    .Y(_06672_),
    .A1(_06669_),
    .A2(_06670_));
 sg13g2_nand2_1 _13911_ (.Y(_06673_),
    .A(_06662_),
    .B(_06672_));
 sg13g2_o21ai_1 _13912_ (.B1(_06670_),
    .Y(_06674_),
    .A1(_06667_),
    .A2(_06669_));
 sg13g2_nor2b_1 _13913_ (.A(_06671_),
    .B_N(_06674_),
    .Y(_06675_));
 sg13g2_nor3_1 _13914_ (.A(_00064_),
    .B(_06545_),
    .C(_06548_),
    .Y(_06676_));
 sg13g2_nor2_1 _13915_ (.A(_06550_),
    .B(_06676_),
    .Y(_06677_));
 sg13g2_o21ai_1 _13916_ (.B1(_06664_),
    .Y(_06678_),
    .A1(_06568_),
    .A2(_06663_));
 sg13g2_nand2b_2 _13917_ (.Y(_06679_),
    .B(_06678_),
    .A_N(_06665_));
 sg13g2_nor2_1 _13918_ (.A(_06677_),
    .B(_06679_),
    .Y(_06680_));
 sg13g2_nand3b_1 _13919_ (.B(_06674_),
    .C(_06680_),
    .Y(_06681_),
    .A_N(_06671_));
 sg13g2_nor2_1 _13920_ (.A(_06662_),
    .B(_06672_),
    .Y(_06682_));
 sg13g2_xor2_1 _13921_ (.B(_06672_),
    .A(_06662_),
    .X(_06683_));
 sg13g2_o21ai_1 _13922_ (.B1(_06673_),
    .Y(_06684_),
    .A1(_06681_),
    .A2(_06682_));
 sg13g2_nand2b_1 _13923_ (.Y(_06685_),
    .B(_06640_),
    .A_N(_06660_));
 sg13g2_nand2b_1 _13924_ (.Y(_06686_),
    .B(_06685_),
    .A_N(_06661_));
 sg13g2_a21oi_1 _13925_ (.A1(_06684_),
    .A2(_06685_),
    .Y(_06687_),
    .B1(_06661_));
 sg13g2_xor2_1 _13926_ (.B(_06638_),
    .A(_06612_),
    .X(_06688_));
 sg13g2_o21ai_1 _13927_ (.B1(_06639_),
    .Y(_06689_),
    .A1(_06687_),
    .A2(_06688_));
 sg13g2_xnor2_1 _13928_ (.Y(_06690_),
    .A(_06609_),
    .B(_06610_));
 sg13g2_a221oi_1 _13929_ (.B2(_06690_),
    .C1(_06611_),
    .B1(_06689_),
    .A1(_06600_),
    .Y(_06691_),
    .A2(_06607_));
 sg13g2_nand2_1 _13930_ (.Y(_06692_),
    .A(_06513_),
    .B(_06561_));
 sg13g2_a21o_1 _13931_ (.A2(_06691_),
    .A1(_06512_),
    .B1(_06602_),
    .X(_06693_));
 sg13g2_xor2_1 _13932_ (.B(_06690_),
    .A(_06689_),
    .X(_06694_));
 sg13g2_o21ai_1 _13933_ (.B1(_06692_),
    .Y(_06695_),
    .A1(_06513_),
    .A2(_06694_));
 sg13g2_o21ai_1 _13934_ (.B1(_06512_),
    .Y(_06696_),
    .A1(_06687_),
    .A2(_06688_));
 sg13g2_a21oi_1 _13935_ (.A1(_06687_),
    .A2(_06688_),
    .Y(_06697_),
    .B1(_06696_));
 sg13g2_a21oi_1 _13936_ (.A1(_06513_),
    .A2(_06608_),
    .Y(_06698_),
    .B1(_06697_));
 sg13g2_o21ai_1 _13937_ (.B1(_06693_),
    .Y(_06699_),
    .A1(_06695_),
    .A2(_06698_));
 sg13g2_nor2b_2 _13938_ (.A(net3655),
    .B_N(_06699_),
    .Y(_06700_));
 sg13g2_a21oi_2 _13939_ (.B1(_06693_),
    .Y(_06701_),
    .A2(_06698_),
    .A1(_06695_));
 sg13g2_nor2_1 _13940_ (.A(_06513_),
    .B(_06679_),
    .Y(_06702_));
 sg13g2_xnor2_1 _13941_ (.Y(_06703_),
    .A(_06677_),
    .B(_06702_));
 sg13g2_nor2_1 _13942_ (.A(_06701_),
    .B(_06703_),
    .Y(_06704_));
 sg13g2_nand2_1 _13943_ (.Y(_06705_),
    .A(net4531),
    .B(_06700_));
 sg13g2_xor2_1 _13944_ (.B(net495),
    .A(net4311),
    .X(_06706_));
 sg13g2_a22oi_1 _13945_ (.Y(_06707_),
    .B1(_00012_),
    .B2(_06706_),
    .A2(net495),
    .A1(net3924));
 sg13g2_o21ai_1 _13946_ (.B1(_06707_),
    .Y(_00641_),
    .A1(_06704_),
    .A2(_06705_));
 sg13g2_and2_1 _13947_ (.A(_06512_),
    .B(_06681_),
    .X(_06708_));
 sg13g2_o21ai_1 _13948_ (.B1(_06708_),
    .Y(_06709_),
    .A1(_06675_),
    .A2(_06680_));
 sg13g2_o21ai_1 _13949_ (.B1(_06709_),
    .Y(_06710_),
    .A1(_06512_),
    .A2(_06670_));
 sg13g2_o21ai_1 _13950_ (.B1(_06700_),
    .Y(_06711_),
    .A1(_06701_),
    .A2(_06710_));
 sg13g2_xor2_1 _13951_ (.B(_04795_),
    .A(_04794_),
    .X(_06712_));
 sg13g2_a21oi_1 _13952_ (.A1(net3655),
    .A2(_06712_),
    .Y(_06713_),
    .B1(net3923));
 sg13g2_a22oi_1 _13953_ (.Y(_00642_),
    .B1(_06711_),
    .B2(_06713_),
    .A2(_03448_),
    .A1(net3923));
 sg13g2_xnor2_1 _13954_ (.Y(_06714_),
    .A(_06681_),
    .B(_06683_));
 sg13g2_nor2_1 _13955_ (.A(_06513_),
    .B(_06714_),
    .Y(_06715_));
 sg13g2_a21oi_1 _13956_ (.A1(_06513_),
    .A2(_06659_),
    .Y(_06716_),
    .B1(_06715_));
 sg13g2_o21ai_1 _13957_ (.B1(_06700_),
    .Y(_06717_),
    .A1(_06701_),
    .A2(_06716_));
 sg13g2_xnor2_1 _13958_ (.Y(_06718_),
    .A(_04792_),
    .B(_04796_));
 sg13g2_a21oi_1 _13959_ (.A1(net3655),
    .A2(_06718_),
    .Y(_06719_),
    .B1(net3923));
 sg13g2_a22oi_1 _13960_ (.Y(_00643_),
    .B1(_06717_),
    .B2(_06719_),
    .A2(_03447_),
    .A1(net3924));
 sg13g2_xnor2_1 _13961_ (.Y(_06720_),
    .A(_06684_),
    .B(_06686_));
 sg13g2_mux2_1 _13962_ (.A0(_06637_),
    .A1(_06720_),
    .S(_06512_),
    .X(_06721_));
 sg13g2_o21ai_1 _13963_ (.B1(_06700_),
    .Y(_06722_),
    .A1(_06701_),
    .A2(_06721_));
 sg13g2_or3_1 _13964_ (.A(_04790_),
    .B(_04791_),
    .C(_04797_),
    .X(_06723_));
 sg13g2_and2_1 _13965_ (.A(_04798_),
    .B(_06723_),
    .X(_06724_));
 sg13g2_a21oi_1 _13966_ (.A1(net3655),
    .A2(_06724_),
    .Y(_06725_),
    .B1(net3923));
 sg13g2_a22oi_1 _13967_ (.Y(_00644_),
    .B1(_06722_),
    .B2(_06725_),
    .A2(_03446_),
    .A1(net3923));
 sg13g2_nand2b_1 _13968_ (.Y(_06726_),
    .B(_06693_),
    .A_N(net3655));
 sg13g2_a21oi_1 _13969_ (.A1(_04789_),
    .A2(_04799_),
    .Y(_06727_),
    .B1(net3923));
 sg13g2_a22oi_1 _13970_ (.Y(_00645_),
    .B1(_06726_),
    .B2(_06727_),
    .A2(_03445_),
    .A1(net3923));
 sg13g2_nand2_1 _13971_ (.Y(_06728_),
    .A(\spiking_network_top_uut.all_data_out[732] ),
    .B(_03667_));
 sg13g2_nor2_1 _13972_ (.A(\spiking_network_top_uut.all_data_out[732] ),
    .B(net3842),
    .Y(_06729_));
 sg13g2_nor2_1 _13973_ (.A(\spiking_network_top_uut.all_data_out[733] ),
    .B(_06729_),
    .Y(_06730_));
 sg13g2_mux2_1 _13974_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[6] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[7] ),
    .S(\spiking_network_top_uut.all_data_out[732] ),
    .X(_06731_));
 sg13g2_a221oi_1 _13975_ (.B2(\spiking_network_top_uut.all_data_out[733] ),
    .C1(_03520_),
    .B1(_06731_),
    .A1(_06728_),
    .Y(_06732_),
    .A2(_06730_));
 sg13g2_mux4_1 _13976_ (.S0(\spiking_network_top_uut.all_data_out[732] ),
    .A0(net3846),
    .A1(net3845),
    .A2(net3844),
    .A3(net3843),
    .S1(\spiking_network_top_uut.all_data_out[733] ),
    .X(_06733_));
 sg13g2_o21ai_1 _13977_ (.B1(net4551),
    .Y(_06734_),
    .A1(\spiking_network_top_uut.all_data_out[734] ),
    .A2(_06733_));
 sg13g2_nand2_1 _13978_ (.Y(_06735_),
    .A(net3934),
    .B(net432));
 sg13g2_o21ai_1 _13979_ (.B1(_06735_),
    .Y(_00646_),
    .A1(_06732_),
    .A2(_06734_));
 sg13g2_mux2_1 _13980_ (.A0(net470),
    .A1(net432),
    .S(net4549),
    .X(_00647_));
 sg13g2_mux4_1 _13981_ (.S0(\spiking_network_top_uut.all_data_out[728] ),
    .A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[0] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[1] ),
    .A2(net3896),
    .A3(net3895),
    .S1(\spiking_network_top_uut.all_data_out[729] ),
    .X(_06736_));
 sg13g2_mux2_1 _13982_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[6] ),
    .A1(net3892),
    .S(\spiking_network_top_uut.all_data_out[728] ),
    .X(_06737_));
 sg13g2_nor2b_1 _13983_ (.A(\spiking_network_top_uut.all_data_out[728] ),
    .B_N(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[4] ),
    .Y(_06738_));
 sg13g2_a21oi_1 _13984_ (.A1(\spiking_network_top_uut.all_data_out[728] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[5] ),
    .Y(_06739_),
    .B1(_06738_));
 sg13g2_o21ai_1 _13985_ (.B1(\spiking_network_top_uut.all_data_out[730] ),
    .Y(_06740_),
    .A1(\spiking_network_top_uut.all_data_out[729] ),
    .A2(_06739_));
 sg13g2_a21oi_1 _13986_ (.A1(\spiking_network_top_uut.all_data_out[729] ),
    .A2(_06737_),
    .Y(_06741_),
    .B1(_06740_));
 sg13g2_o21ai_1 _13987_ (.B1(net4547),
    .Y(_06742_),
    .A1(\spiking_network_top_uut.all_data_out[730] ),
    .A2(_06736_));
 sg13g2_nand2_1 _13988_ (.Y(_06743_),
    .A(net3933),
    .B(net117));
 sg13g2_o21ai_1 _13989_ (.B1(_06743_),
    .Y(_00648_),
    .A1(_06741_),
    .A2(_06742_));
 sg13g2_mux2_1 _13990_ (.A0(net278),
    .A1(net117),
    .S(net4547),
    .X(_00649_));
 sg13g2_mux4_1 _13991_ (.S0(\spiking_network_top_uut.all_data_out[724] ),
    .A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[0] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[1] ),
    .A2(net3889),
    .A3(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[3] ),
    .S1(\spiking_network_top_uut.all_data_out[725] ),
    .X(_06744_));
 sg13g2_mux2_1 _13992_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[6] ),
    .A1(net3885),
    .S(\spiking_network_top_uut.all_data_out[724] ),
    .X(_06745_));
 sg13g2_nor2b_1 _13993_ (.A(\spiking_network_top_uut.all_data_out[724] ),
    .B_N(net3887),
    .Y(_06746_));
 sg13g2_a21oi_1 _13994_ (.A1(\spiking_network_top_uut.all_data_out[724] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[5] ),
    .Y(_06747_),
    .B1(_06746_));
 sg13g2_o21ai_1 _13995_ (.B1(\spiking_network_top_uut.all_data_out[726] ),
    .Y(_06748_),
    .A1(\spiking_network_top_uut.all_data_out[725] ),
    .A2(_06747_));
 sg13g2_a21oi_1 _13996_ (.A1(\spiking_network_top_uut.all_data_out[725] ),
    .A2(_06745_),
    .Y(_06749_),
    .B1(_06748_));
 sg13g2_o21ai_1 _13997_ (.B1(net4561),
    .Y(_06750_),
    .A1(\spiking_network_top_uut.all_data_out[726] ),
    .A2(_06744_));
 sg13g2_nand2_1 _13998_ (.Y(_06751_),
    .A(net3935),
    .B(net80));
 sg13g2_o21ai_1 _13999_ (.B1(_06751_),
    .Y(_00650_),
    .A1(_06749_),
    .A2(_06750_));
 sg13g2_mux2_1 _14000_ (.A0(net462),
    .A1(net80),
    .S(net4561),
    .X(_00651_));
 sg13g2_mux4_1 _14001_ (.S0(\spiking_network_top_uut.all_data_out[720] ),
    .A0(net3884),
    .A1(net3883),
    .A2(net3882),
    .A3(net3881),
    .S1(\spiking_network_top_uut.all_data_out[721] ),
    .X(_06752_));
 sg13g2_mux2_1 _14002_ (.A0(net3878),
    .A1(net3877),
    .S(\spiking_network_top_uut.all_data_out[720] ),
    .X(_06753_));
 sg13g2_nor2b_1 _14003_ (.A(\spiking_network_top_uut.all_data_out[720] ),
    .B_N(net3880),
    .Y(_06754_));
 sg13g2_a21oi_1 _14004_ (.A1(\spiking_network_top_uut.all_data_out[720] ),
    .A2(net3879),
    .Y(_06755_),
    .B1(_06754_));
 sg13g2_o21ai_1 _14005_ (.B1(\spiking_network_top_uut.all_data_out[722] ),
    .Y(_06756_),
    .A1(\spiking_network_top_uut.all_data_out[721] ),
    .A2(_06755_));
 sg13g2_a21oi_1 _14006_ (.A1(\spiking_network_top_uut.all_data_out[721] ),
    .A2(_06753_),
    .Y(_06757_),
    .B1(_06756_));
 sg13g2_o21ai_1 _14007_ (.B1(net4554),
    .Y(_06758_),
    .A1(\spiking_network_top_uut.all_data_out[722] ),
    .A2(_06752_));
 sg13g2_nand2_1 _14008_ (.Y(_06759_),
    .A(net3938),
    .B(net286));
 sg13g2_o21ai_1 _14009_ (.B1(_06759_),
    .Y(_00652_),
    .A1(_06757_),
    .A2(_06758_));
 sg13g2_mux2_1 _14010_ (.A0(net400),
    .A1(net286),
    .S(net4557),
    .X(_00653_));
 sg13g2_nand2b_1 _14011_ (.Y(_06760_),
    .B(\spiking_network_top_uut.all_data_out[716] ),
    .A_N(net3871));
 sg13g2_nor2_1 _14012_ (.A(\spiking_network_top_uut.all_data_out[716] ),
    .B(net3872),
    .Y(_06761_));
 sg13g2_nor2_1 _14013_ (.A(\spiking_network_top_uut.all_data_out[717] ),
    .B(_06761_),
    .Y(_06762_));
 sg13g2_mux2_1 _14014_ (.A0(net3870),
    .A1(net3869),
    .S(\spiking_network_top_uut.all_data_out[716] ),
    .X(_06763_));
 sg13g2_a221oi_1 _14015_ (.B2(\spiking_network_top_uut.all_data_out[717] ),
    .C1(_03523_),
    .B1(_06763_),
    .A1(_06760_),
    .Y(_06764_),
    .A2(_06762_));
 sg13g2_mux4_1 _14016_ (.S0(\spiking_network_top_uut.all_data_out[716] ),
    .A0(net3876),
    .A1(net3875),
    .A2(net3874),
    .A3(net3873),
    .S1(\spiking_network_top_uut.all_data_out[717] ),
    .X(_06765_));
 sg13g2_o21ai_1 _14017_ (.B1(net4566),
    .Y(_06766_),
    .A1(\spiking_network_top_uut.all_data_out[718] ),
    .A2(_06765_));
 sg13g2_nand2_1 _14018_ (.Y(_06767_),
    .A(net3937),
    .B(net134));
 sg13g2_o21ai_1 _14019_ (.B1(_06767_),
    .Y(_00654_),
    .A1(_06764_),
    .A2(_06766_));
 sg13g2_mux2_1 _14020_ (.A0(net263),
    .A1(net134),
    .S(net4568),
    .X(_00655_));
 sg13g2_mux4_1 _14021_ (.S0(\spiking_network_top_uut.all_data_out[712] ),
    .A0(net3868),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[1] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[2] ),
    .A3(net3865),
    .S1(\spiking_network_top_uut.all_data_out[713] ),
    .X(_06768_));
 sg13g2_mux2_1 _14022_ (.A0(net3862),
    .A1(net3861),
    .S(\spiking_network_top_uut.all_data_out[712] ),
    .X(_06769_));
 sg13g2_nor2b_1 _14023_ (.A(\spiking_network_top_uut.all_data_out[712] ),
    .B_N(net3864),
    .Y(_06770_));
 sg13g2_a21oi_1 _14024_ (.A1(\spiking_network_top_uut.all_data_out[712] ),
    .A2(net3863),
    .Y(_06771_),
    .B1(_06770_));
 sg13g2_o21ai_1 _14025_ (.B1(\spiking_network_top_uut.all_data_out[714] ),
    .Y(_06772_),
    .A1(\spiking_network_top_uut.all_data_out[713] ),
    .A2(_06771_));
 sg13g2_a21oi_1 _14026_ (.A1(\spiking_network_top_uut.all_data_out[713] ),
    .A2(_06769_),
    .Y(_06773_),
    .B1(_06772_));
 sg13g2_o21ai_1 _14027_ (.B1(net4564),
    .Y(_06774_),
    .A1(\spiking_network_top_uut.all_data_out[714] ),
    .A2(_06768_));
 sg13g2_nand2_1 _14028_ (.Y(_06775_),
    .A(net3935),
    .B(net103));
 sg13g2_o21ai_1 _14029_ (.B1(_06775_),
    .Y(_00656_),
    .A1(_06773_),
    .A2(_06774_));
 sg13g2_mux2_1 _14030_ (.A0(net423),
    .A1(net103),
    .S(net4565),
    .X(_00657_));
 sg13g2_mux4_1 _14031_ (.S0(\spiking_network_top_uut.all_data_out[708] ),
    .A0(net3860),
    .A1(net3859),
    .A2(net3858),
    .A3(net3857),
    .S1(\spiking_network_top_uut.all_data_out[709] ),
    .X(_06776_));
 sg13g2_mux2_1 _14032_ (.A0(net3855),
    .A1(net3854),
    .S(\spiking_network_top_uut.all_data_out[708] ),
    .X(_06777_));
 sg13g2_nor2b_1 _14033_ (.A(\spiking_network_top_uut.all_data_out[708] ),
    .B_N(net3856),
    .Y(_06778_));
 sg13g2_a21oi_1 _14034_ (.A1(\spiking_network_top_uut.all_data_out[708] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[5] ),
    .Y(_06779_),
    .B1(_06778_));
 sg13g2_o21ai_1 _14035_ (.B1(\spiking_network_top_uut.all_data_out[710] ),
    .Y(_06780_),
    .A1(\spiking_network_top_uut.all_data_out[709] ),
    .A2(_06779_));
 sg13g2_a21oi_1 _14036_ (.A1(\spiking_network_top_uut.all_data_out[709] ),
    .A2(_06777_),
    .Y(_06781_),
    .B1(_06780_));
 sg13g2_o21ai_1 _14037_ (.B1(net4540),
    .Y(_06782_),
    .A1(\spiking_network_top_uut.all_data_out[710] ),
    .A2(_06776_));
 sg13g2_nand2_1 _14038_ (.Y(_06783_),
    .A(net3932),
    .B(net66));
 sg13g2_o21ai_1 _14039_ (.B1(_06783_),
    .Y(_00658_),
    .A1(_06781_),
    .A2(_06782_));
 sg13g2_mux2_1 _14040_ (.A0(net158),
    .A1(net66),
    .S(net4540),
    .X(_00659_));
 sg13g2_mux4_1 _14041_ (.S0(\spiking_network_top_uut.all_data_out[704] ),
    .A0(net3853),
    .A1(net3852),
    .A2(net3851),
    .A3(net3850),
    .S1(\spiking_network_top_uut.all_data_out[705] ),
    .X(_06784_));
 sg13g2_mux2_1 _14042_ (.A0(net3848),
    .A1(net3847),
    .S(\spiking_network_top_uut.all_data_out[704] ),
    .X(_06785_));
 sg13g2_nor2b_1 _14043_ (.A(\spiking_network_top_uut.all_data_out[704] ),
    .B_N(net3849),
    .Y(_06786_));
 sg13g2_a21oi_1 _14044_ (.A1(\spiking_network_top_uut.all_data_out[704] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[5] ),
    .Y(_06787_),
    .B1(_06786_));
 sg13g2_o21ai_1 _14045_ (.B1(\spiking_network_top_uut.all_data_out[706] ),
    .Y(_06788_),
    .A1(\spiking_network_top_uut.all_data_out[705] ),
    .A2(_06787_));
 sg13g2_a21oi_2 _14046_ (.B1(_06788_),
    .Y(_06789_),
    .A2(_06785_),
    .A1(\spiking_network_top_uut.all_data_out[705] ));
 sg13g2_o21ai_1 _14047_ (.B1(net4539),
    .Y(_06790_),
    .A1(\spiking_network_top_uut.all_data_out[706] ),
    .A2(_06784_));
 sg13g2_nand2_1 _14048_ (.Y(_06791_),
    .A(net3932),
    .B(net458));
 sg13g2_o21ai_1 _14049_ (.B1(_06791_),
    .Y(_00660_),
    .A1(_06789_),
    .A2(_06790_));
 sg13g2_nor3_2 _14050_ (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[2] ),
    .B(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[1] ),
    .C(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[0] ),
    .Y(_06792_));
 sg13g2_nand2b_1 _14051_ (.Y(_06793_),
    .B(_06792_),
    .A_N(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[3] ));
 sg13g2_nor2_2 _14052_ (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[4] ),
    .B(_06793_),
    .Y(_06794_));
 sg13g2_or2_2 _14053_ (.X(_06795_),
    .B(_06793_),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[4] ));
 sg13g2_o21ai_1 _14054_ (.B1(net4531),
    .Y(_06796_),
    .A1(net3652),
    .A2(_06795_));
 sg13g2_nor2b_1 _14055_ (.A(net3651),
    .B_N(net346),
    .Y(_06797_));
 sg13g2_a21oi_1 _14056_ (.A1(net4284),
    .A2(net3651),
    .Y(_06798_),
    .B1(_06797_));
 sg13g2_nand2_1 _14057_ (.Y(_06799_),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[0] ),
    .B(_06796_));
 sg13g2_o21ai_1 _14058_ (.B1(_06799_),
    .Y(_00661_),
    .A1(_06796_),
    .A2(_06798_));
 sg13g2_xor2_1 _14059_ (.B(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[0] ),
    .A(net419),
    .X(_06800_));
 sg13g2_nor2_1 _14060_ (.A(net3651),
    .B(_06800_),
    .Y(_06801_));
 sg13g2_a21oi_1 _14061_ (.A1(net4281),
    .A2(net3651),
    .Y(_06802_),
    .B1(_06801_));
 sg13g2_nand2_1 _14062_ (.Y(_06803_),
    .A(net419),
    .B(_06796_));
 sg13g2_o21ai_1 _14063_ (.B1(_06803_),
    .Y(_00662_),
    .A1(_06796_),
    .A2(_06802_));
 sg13g2_nand2_1 _14064_ (.Y(_06804_),
    .A(net4277),
    .B(net3651));
 sg13g2_o21ai_1 _14065_ (.B1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[2] ),
    .Y(_06805_),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[1] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[0] ));
 sg13g2_nor2b_1 _14066_ (.A(_06792_),
    .B_N(_06805_),
    .Y(_06806_));
 sg13g2_o21ai_1 _14067_ (.B1(_06804_),
    .Y(_06807_),
    .A1(net3651),
    .A2(_06806_));
 sg13g2_mux2_1 _14068_ (.A0(_06807_),
    .A1(net435),
    .S(_06796_),
    .X(_00663_));
 sg13g2_nand2_1 _14069_ (.Y(_06808_),
    .A(net4274),
    .B(net3651));
 sg13g2_xnor2_1 _14070_ (.Y(_06809_),
    .A(net398),
    .B(_06792_));
 sg13g2_o21ai_1 _14071_ (.B1(_06808_),
    .Y(_06810_),
    .A1(net3651),
    .A2(_06809_));
 sg13g2_mux2_1 _14072_ (.A0(_06810_),
    .A1(net398),
    .S(_06796_),
    .X(_00664_));
 sg13g2_nand2_1 _14073_ (.Y(_06811_),
    .A(net359),
    .B(net3924));
 sg13g2_nor2b_1 _14074_ (.A(net4270),
    .B_N(net3652),
    .Y(_06812_));
 sg13g2_nand3_1 _14075_ (.B(net4531),
    .C(_06793_),
    .A(net359),
    .Y(_06813_));
 sg13g2_nor2b_1 _14076_ (.A(_00013_),
    .B_N(_06813_),
    .Y(_06814_));
 sg13g2_o21ai_1 _14077_ (.B1(_06811_),
    .Y(_00665_),
    .A1(_06812_),
    .A2(_06814_));
 sg13g2_mux2_1 _14078_ (.A0(net166),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_reg1 ),
    .S(net4541),
    .X(_00666_));
 sg13g2_nor2_1 _14079_ (.A(_00067_),
    .B(net3740),
    .Y(_06815_));
 sg13g2_nor2_2 _14080_ (.A(net3745),
    .B(_06815_),
    .Y(_06816_));
 sg13g2_nor2_1 _14081_ (.A(_00067_),
    .B(_06816_),
    .Y(_06817_));
 sg13g2_nand2b_1 _14082_ (.Y(_06818_),
    .B(_06816_),
    .A_N(_00067_));
 sg13g2_o21ai_1 _14083_ (.B1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ),
    .Y(_06819_),
    .A1(_00067_),
    .A2(_06816_));
 sg13g2_inv_1 _14084_ (.Y(_06820_),
    .A(_06819_));
 sg13g2_a21o_1 _14085_ (.A2(net3745),
    .A1(_00068_),
    .B1(_06816_),
    .X(_06821_));
 sg13g2_and2_1 _14086_ (.A(_00069_),
    .B(net3745),
    .X(_06822_));
 sg13g2_o21ai_1 _14087_ (.B1(net3916),
    .Y(_06823_),
    .A1(_00068_),
    .A2(net3904));
 sg13g2_a21oi_2 _14088_ (.B1(_06823_),
    .Y(_06824_),
    .A2(_06815_),
    .A1(net3904));
 sg13g2_o21ai_1 _14089_ (.B1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ),
    .Y(_06825_),
    .A1(_06822_),
    .A2(_06824_));
 sg13g2_o21ai_1 _14090_ (.B1(net3913),
    .Y(_06826_),
    .A1(_00067_),
    .A2(net3910));
 sg13g2_a221oi_1 _14091_ (.B2(_00068_),
    .C1(net3745),
    .B1(net3901),
    .A1(_00069_),
    .Y(_06827_),
    .A2(net3738));
 sg13g2_a22oi_1 _14092_ (.Y(_06828_),
    .B1(_06826_),
    .B2(_06827_),
    .A2(net3745),
    .A1(_03483_));
 sg13g2_nor2b_1 _14093_ (.A(_06828_),
    .B_N(_00070_),
    .Y(_06829_));
 sg13g2_nor3_1 _14094_ (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ),
    .B(_06822_),
    .C(_06824_),
    .Y(_06830_));
 sg13g2_or3_1 _14095_ (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ),
    .B(_06822_),
    .C(_06824_),
    .X(_06831_));
 sg13g2_nand2_1 _14096_ (.Y(_06832_),
    .A(_06825_),
    .B(_06831_));
 sg13g2_o21ai_1 _14097_ (.B1(_06825_),
    .Y(_06833_),
    .A1(_06829_),
    .A2(_06830_));
 sg13g2_xor2_1 _14098_ (.B(_06821_),
    .A(_00069_),
    .X(_06834_));
 sg13g2_nor2b_1 _14099_ (.A(_06834_),
    .B_N(_06833_),
    .Y(_06835_));
 sg13g2_a21o_1 _14100_ (.A2(_06821_),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ),
    .B1(_06835_),
    .X(_06836_));
 sg13g2_xnor2_1 _14101_ (.Y(_06837_),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ),
    .B(_06817_));
 sg13g2_a21oi_1 _14102_ (.A1(_06836_),
    .A2(_06837_),
    .Y(_06838_),
    .B1(_06820_));
 sg13g2_a22oi_1 _14103_ (.Y(_06839_),
    .B1(_06818_),
    .B2(_06838_),
    .A2(_06816_),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ));
 sg13g2_a21oi_2 _14104_ (.B1(_06839_),
    .Y(_06840_),
    .A2(_00067_),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ));
 sg13g2_nor2_1 _14105_ (.A(_06794_),
    .B(_06840_),
    .Y(_06841_));
 sg13g2_mux2_1 _14106_ (.A0(net4599),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[707] ),
    .X(_06842_));
 sg13g2_nand2_1 _14107_ (.Y(_06843_),
    .A(\spiking_network_top_uut.all_data_out[225] ),
    .B(_06842_));
 sg13g2_mux2_1 _14108_ (.A0(net4598),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[711] ),
    .X(_06844_));
 sg13g2_nand2_1 _14109_ (.Y(_06845_),
    .A(\spiking_network_top_uut.all_data_out[227] ),
    .B(_06844_));
 sg13g2_nor2_1 _14110_ (.A(_06843_),
    .B(_06845_),
    .Y(_06846_));
 sg13g2_nand4_1 _14111_ (.B(\spiking_network_top_uut.all_data_out[226] ),
    .C(_06842_),
    .A(\spiking_network_top_uut.all_data_out[224] ),
    .Y(_06847_),
    .D(_06844_));
 sg13g2_inv_1 _14112_ (.Y(_06848_),
    .A(_06847_));
 sg13g2_xor2_1 _14113_ (.B(_06845_),
    .A(_06843_),
    .X(_06849_));
 sg13g2_a21oi_2 _14114_ (.B1(_06846_),
    .Y(_06850_),
    .A2(_06849_),
    .A1(_06847_));
 sg13g2_mux2_2 _14115_ (.A0(net4597),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[715] ),
    .X(_06851_));
 sg13g2_nand2_1 _14116_ (.Y(_06852_),
    .A(\spiking_network_top_uut.all_data_out[229] ),
    .B(_06851_));
 sg13g2_mux2_2 _14117_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.spike_out ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[719] ),
    .X(_06853_));
 sg13g2_nand2_2 _14118_ (.Y(_06854_),
    .A(\spiking_network_top_uut.all_data_out[231] ),
    .B(_06853_));
 sg13g2_nor2_1 _14119_ (.A(_06852_),
    .B(_06854_),
    .Y(_06855_));
 sg13g2_nand2_1 _14120_ (.Y(_06856_),
    .A(\spiking_network_top_uut.all_data_out[228] ),
    .B(_06851_));
 sg13g2_nand2_2 _14121_ (.Y(_06857_),
    .A(\spiking_network_top_uut.all_data_out[230] ),
    .B(_06853_));
 sg13g2_or2_2 _14122_ (.X(_06858_),
    .B(_06857_),
    .A(_06856_));
 sg13g2_xor2_1 _14123_ (.B(_06854_),
    .A(_06852_),
    .X(_06859_));
 sg13g2_a21oi_2 _14124_ (.B1(_06855_),
    .Y(_06860_),
    .A2(_06859_),
    .A1(_06858_));
 sg13g2_mux2_2 _14125_ (.A0(net4595),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[723] ),
    .X(_06861_));
 sg13g2_mux2_2 _14126_ (.A0(net4594),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[727] ),
    .X(_06862_));
 sg13g2_a22oi_1 _14127_ (.Y(_06863_),
    .B1(_06862_),
    .B2(\spiking_network_top_uut.all_data_out[235] ),
    .A2(_06861_),
    .A1(\spiking_network_top_uut.all_data_out[233] ));
 sg13g2_and4_2 _14128_ (.A(\spiking_network_top_uut.all_data_out[232] ),
    .B(\spiking_network_top_uut.all_data_out[234] ),
    .C(_06861_),
    .D(_06862_),
    .X(_06864_));
 sg13g2_nand4_1 _14129_ (.B(\spiking_network_top_uut.all_data_out[234] ),
    .C(_06861_),
    .A(\spiking_network_top_uut.all_data_out[232] ),
    .Y(_06865_),
    .D(_06862_));
 sg13g2_and4_1 _14130_ (.A(\spiking_network_top_uut.all_data_out[233] ),
    .B(\spiking_network_top_uut.all_data_out[235] ),
    .C(_06861_),
    .D(_06862_),
    .X(_06866_));
 sg13g2_nand4_1 _14131_ (.B(\spiking_network_top_uut.all_data_out[235] ),
    .C(_06861_),
    .A(\spiking_network_top_uut.all_data_out[233] ),
    .Y(_06867_),
    .D(_06862_));
 sg13g2_nand3b_1 _14132_ (.B(_06864_),
    .C(_06867_),
    .Y(_06868_),
    .A_N(_06863_));
 sg13g2_a21oi_2 _14133_ (.B1(_06863_),
    .Y(_06869_),
    .A2(_06867_),
    .A1(_06864_));
 sg13g2_mux2_2 _14134_ (.A0(net4593),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[731] ),
    .X(_06870_));
 sg13g2_mux2_2 _14135_ (.A0(net4592),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[735] ),
    .X(_06871_));
 sg13g2_and4_1 _14136_ (.A(\spiking_network_top_uut.all_data_out[237] ),
    .B(\spiking_network_top_uut.all_data_out[239] ),
    .C(_06870_),
    .D(_06871_),
    .X(_06872_));
 sg13g2_nand4_1 _14137_ (.B(\spiking_network_top_uut.all_data_out[239] ),
    .C(_06870_),
    .A(\spiking_network_top_uut.all_data_out[237] ),
    .Y(_06873_),
    .D(_06871_));
 sg13g2_and4_2 _14138_ (.A(\spiking_network_top_uut.all_data_out[236] ),
    .B(\spiking_network_top_uut.all_data_out[238] ),
    .C(_06870_),
    .D(_06871_),
    .X(_06874_));
 sg13g2_a22oi_1 _14139_ (.Y(_06875_),
    .B1(_06871_),
    .B2(\spiking_network_top_uut.all_data_out[239] ),
    .A2(_06870_),
    .A1(\spiking_network_top_uut.all_data_out[237] ));
 sg13g2_or3_2 _14140_ (.A(_06872_),
    .B(_06874_),
    .C(_06875_),
    .X(_06876_));
 sg13g2_o21ai_1 _14141_ (.B1(_06873_),
    .Y(_06877_),
    .A1(_06874_),
    .A2(_06875_));
 sg13g2_nand3b_1 _14142_ (.B(_06869_),
    .C(_06877_),
    .Y(_06878_),
    .A_N(_06860_));
 sg13g2_inv_1 _14143_ (.Y(_06879_),
    .A(_06878_));
 sg13g2_or2_2 _14144_ (.X(_06880_),
    .B(_06878_),
    .A(_06850_));
 sg13g2_nor2_1 _14145_ (.A(_06869_),
    .B(_06877_),
    .Y(_06881_));
 sg13g2_and2_1 _14146_ (.A(_06860_),
    .B(_06881_),
    .X(_06882_));
 sg13g2_nand2_2 _14147_ (.Y(_06883_),
    .A(_06850_),
    .B(_06882_));
 sg13g2_and2_1 _14148_ (.A(_06880_),
    .B(_06883_),
    .X(_06884_));
 sg13g2_xnor2_1 _14149_ (.Y(_06885_),
    .A(_06818_),
    .B(_06838_));
 sg13g2_nand2_1 _14150_ (.Y(_06886_),
    .A(_06884_),
    .B(_06885_));
 sg13g2_nand2_1 _14151_ (.Y(_06887_),
    .A(_06880_),
    .B(_06886_));
 sg13g2_xor2_1 _14152_ (.B(_06884_),
    .A(_06840_),
    .X(_06888_));
 sg13g2_nand2_1 _14153_ (.Y(_06889_),
    .A(_06887_),
    .B(_06888_));
 sg13g2_xnor2_1 _14154_ (.Y(_06890_),
    .A(_06884_),
    .B(_06885_));
 sg13g2_o21ai_1 _14155_ (.B1(_06874_),
    .Y(_06891_),
    .A1(_06872_),
    .A2(_06875_));
 sg13g2_o21ai_1 _14156_ (.B1(_06865_),
    .Y(_06892_),
    .A1(_06863_),
    .A2(_06866_));
 sg13g2_o21ai_1 _14157_ (.B1(_06864_),
    .Y(_06893_),
    .A1(_06863_),
    .A2(_06866_));
 sg13g2_nand3b_1 _14158_ (.B(_06865_),
    .C(_06867_),
    .Y(_06894_),
    .A_N(_06863_));
 sg13g2_a22oi_1 _14159_ (.Y(_06895_),
    .B1(_06893_),
    .B2(_06894_),
    .A2(_06891_),
    .A1(_06876_));
 sg13g2_xor2_1 _14160_ (.B(_06859_),
    .A(_06858_),
    .X(_06896_));
 sg13g2_xnor2_1 _14161_ (.Y(_06897_),
    .A(_06858_),
    .B(_06859_));
 sg13g2_and4_1 _14162_ (.A(_06876_),
    .B(_06891_),
    .C(_06893_),
    .D(_06894_),
    .X(_06898_));
 sg13g2_nand4_1 _14163_ (.B(_06891_),
    .C(_06893_),
    .A(_06876_),
    .Y(_06899_),
    .D(_06894_));
 sg13g2_and4_1 _14164_ (.A(_06868_),
    .B(_06876_),
    .C(_06891_),
    .D(_06892_),
    .X(_06900_));
 sg13g2_a22oi_1 _14165_ (.Y(_06901_),
    .B1(_06892_),
    .B2(_06868_),
    .A2(_06891_),
    .A1(_06876_));
 sg13g2_nor3_2 _14166_ (.A(_06895_),
    .B(_06896_),
    .C(_06898_),
    .Y(_06902_));
 sg13g2_a21oi_2 _14167_ (.B1(_06895_),
    .Y(_06903_),
    .A2(_06899_),
    .A1(_06897_));
 sg13g2_xor2_1 _14168_ (.B(_06877_),
    .A(_06869_),
    .X(_06904_));
 sg13g2_xnor2_1 _14169_ (.Y(_06905_),
    .A(_06860_),
    .B(_06904_));
 sg13g2_nand2b_1 _14170_ (.Y(_06906_),
    .B(_06905_),
    .A_N(_06903_));
 sg13g2_xnor2_1 _14171_ (.Y(_06907_),
    .A(_06903_),
    .B(_06905_));
 sg13g2_nand2b_1 _14172_ (.Y(_06908_),
    .B(_06907_),
    .A_N(_06850_));
 sg13g2_nand2_2 _14173_ (.Y(_06909_),
    .A(_06906_),
    .B(_06908_));
 sg13g2_nor2_1 _14174_ (.A(_06879_),
    .B(_06882_),
    .Y(_06910_));
 sg13g2_xnor2_1 _14175_ (.Y(_06911_),
    .A(_06850_),
    .B(_06910_));
 sg13g2_and2_1 _14176_ (.A(_06909_),
    .B(_06911_),
    .X(_06912_));
 sg13g2_xor2_1 _14177_ (.B(_06911_),
    .A(_06909_),
    .X(_06913_));
 sg13g2_xnor2_1 _14178_ (.Y(_06914_),
    .A(_06836_),
    .B(_06837_));
 sg13g2_inv_1 _14179_ (.Y(_06915_),
    .A(_06914_));
 sg13g2_a21oi_2 _14180_ (.B1(_06912_),
    .Y(_06916_),
    .A2(_06915_),
    .A1(_06913_));
 sg13g2_nor2_1 _14181_ (.A(_06890_),
    .B(_06916_),
    .Y(_06917_));
 sg13g2_xnor2_1 _14182_ (.Y(_06918_),
    .A(_06913_),
    .B(_06914_));
 sg13g2_a22oi_1 _14183_ (.Y(_06919_),
    .B1(_06871_),
    .B2(\spiking_network_top_uut.all_data_out[238] ),
    .A2(_06870_),
    .A1(\spiking_network_top_uut.all_data_out[236] ));
 sg13g2_nor2_2 _14184_ (.A(_06874_),
    .B(_06919_),
    .Y(_06920_));
 sg13g2_a22oi_1 _14185_ (.Y(_06921_),
    .B1(_06862_),
    .B2(\spiking_network_top_uut.all_data_out[234] ),
    .A2(_06861_),
    .A1(\spiking_network_top_uut.all_data_out[232] ));
 sg13g2_nor2_1 _14186_ (.A(_06864_),
    .B(_06921_),
    .Y(_06922_));
 sg13g2_and2_1 _14187_ (.A(_06920_),
    .B(_06922_),
    .X(_06923_));
 sg13g2_xor2_1 _14188_ (.B(_06857_),
    .A(_06856_),
    .X(_06924_));
 sg13g2_xor2_1 _14189_ (.B(_06922_),
    .A(_06920_),
    .X(_06925_));
 sg13g2_a21oi_2 _14190_ (.B1(_06923_),
    .Y(_06926_),
    .A2(_06925_),
    .A1(_06924_));
 sg13g2_nor3_2 _14191_ (.A(_06897_),
    .B(_06900_),
    .C(_06901_),
    .Y(_06927_));
 sg13g2_nor3_1 _14192_ (.A(_06902_),
    .B(_06926_),
    .C(_06927_),
    .Y(_06928_));
 sg13g2_or3_1 _14193_ (.A(_06902_),
    .B(_06926_),
    .C(_06927_),
    .X(_06929_));
 sg13g2_xnor2_1 _14194_ (.Y(_06930_),
    .A(_06847_),
    .B(_06849_));
 sg13g2_o21ai_1 _14195_ (.B1(_06926_),
    .Y(_06931_),
    .A1(_06902_),
    .A2(_06927_));
 sg13g2_nand3_1 _14196_ (.B(_06930_),
    .C(_06931_),
    .A(_06929_),
    .Y(_06932_));
 sg13g2_a21o_2 _14197_ (.A2(_06931_),
    .A1(_06930_),
    .B1(_06928_),
    .X(_06933_));
 sg13g2_xnor2_1 _14198_ (.Y(_06934_),
    .A(_06850_),
    .B(_06907_));
 sg13g2_nand2_1 _14199_ (.Y(_06935_),
    .A(_06933_),
    .B(_06934_));
 sg13g2_xnor2_1 _14200_ (.Y(_06936_),
    .A(_06933_),
    .B(_06934_));
 sg13g2_xor2_1 _14201_ (.B(_06834_),
    .A(_06833_),
    .X(_06937_));
 sg13g2_o21ai_1 _14202_ (.B1(_06935_),
    .Y(_06938_),
    .A1(_06936_),
    .A2(_06937_));
 sg13g2_nand2_1 _14203_ (.Y(_06939_),
    .A(_06918_),
    .B(_06938_));
 sg13g2_xor2_1 _14204_ (.B(_06937_),
    .A(_06936_),
    .X(_06940_));
 sg13g2_a22oi_1 _14205_ (.Y(_06941_),
    .B1(_06844_),
    .B2(\spiking_network_top_uut.all_data_out[226] ),
    .A2(_06842_),
    .A1(\spiking_network_top_uut.all_data_out[224] ));
 sg13g2_xnor2_1 _14206_ (.Y(_06942_),
    .A(_06924_),
    .B(_06925_));
 sg13g2_nor3_2 _14207_ (.A(_06848_),
    .B(_06941_),
    .C(_06942_),
    .Y(_06943_));
 sg13g2_a21o_2 _14208_ (.A2(_06931_),
    .A1(_06929_),
    .B1(_06930_),
    .X(_06944_));
 sg13g2_nand3_1 _14209_ (.B(_06943_),
    .C(_06944_),
    .A(_06932_),
    .Y(_06945_));
 sg13g2_a21oi_1 _14210_ (.A1(_06932_),
    .A2(_06944_),
    .Y(_06946_),
    .B1(_06943_));
 sg13g2_a21o_1 _14211_ (.A2(_06944_),
    .A1(_06932_),
    .B1(_06943_),
    .X(_06947_));
 sg13g2_xnor2_1 _14212_ (.Y(_06948_),
    .A(_06829_),
    .B(_06832_));
 sg13g2_inv_1 _14213_ (.Y(_06949_),
    .A(_06948_));
 sg13g2_and3_1 _14214_ (.X(_06950_),
    .A(_06945_),
    .B(_06947_),
    .C(_06949_));
 sg13g2_o21ai_1 _14215_ (.B1(_06945_),
    .Y(_06951_),
    .A1(_06946_),
    .A2(_06948_));
 sg13g2_and2_1 _14216_ (.A(_06940_),
    .B(_06951_),
    .X(_06952_));
 sg13g2_a21oi_1 _14217_ (.A1(_06945_),
    .A2(_06947_),
    .Y(_06953_),
    .B1(_06949_));
 sg13g2_nor2_1 _14218_ (.A(_06950_),
    .B(_06953_),
    .Y(_06954_));
 sg13g2_xnor2_1 _14219_ (.Y(_06955_),
    .A(_00070_),
    .B(_06828_));
 sg13g2_o21ai_1 _14220_ (.B1(_06942_),
    .Y(_06956_),
    .A1(_06848_),
    .A2(_06941_));
 sg13g2_nand2b_2 _14221_ (.Y(_06957_),
    .B(_06956_),
    .A_N(_06943_));
 sg13g2_nor2_1 _14222_ (.A(_06955_),
    .B(_06957_),
    .Y(_06958_));
 sg13g2_nor4_2 _14223_ (.A(_06950_),
    .B(_06953_),
    .C(_06955_),
    .Y(_06959_),
    .D(_06957_));
 sg13g2_xor2_1 _14224_ (.B(_06951_),
    .A(_06940_),
    .X(_06960_));
 sg13g2_a21oi_2 _14225_ (.B1(_06952_),
    .Y(_06961_),
    .A2(_06960_),
    .A1(_06959_));
 sg13g2_xnor2_1 _14226_ (.Y(_06962_),
    .A(_06918_),
    .B(_06938_));
 sg13g2_o21ai_1 _14227_ (.B1(_06939_),
    .Y(_06963_),
    .A1(_06961_),
    .A2(_06962_));
 sg13g2_nand2_1 _14228_ (.Y(_06964_),
    .A(_06890_),
    .B(_06916_));
 sg13g2_xnor2_1 _14229_ (.Y(_06965_),
    .A(_06890_),
    .B(_06916_));
 sg13g2_nor2b_1 _14230_ (.A(_06965_),
    .B_N(_06963_),
    .Y(_06966_));
 sg13g2_a21oi_1 _14231_ (.A1(_06963_),
    .A2(_06964_),
    .Y(_06967_),
    .B1(_06917_));
 sg13g2_xnor2_1 _14232_ (.Y(_06968_),
    .A(_06887_),
    .B(_06888_));
 sg13g2_o21ai_1 _14233_ (.B1(_06889_),
    .Y(_06969_),
    .A1(_06967_),
    .A2(_06968_));
 sg13g2_mux2_1 _14234_ (.A0(_06883_),
    .A1(_06880_),
    .S(_06840_),
    .X(_06970_));
 sg13g2_xnor2_1 _14235_ (.Y(_06971_),
    .A(_06969_),
    .B(_06970_));
 sg13g2_a21oi_2 _14236_ (.B1(_06841_),
    .Y(_06972_),
    .A2(_06971_),
    .A1(_06794_));
 sg13g2_nand2b_1 _14237_ (.Y(_06973_),
    .B(_06965_),
    .A_N(_06963_));
 sg13g2_nor2_1 _14238_ (.A(_06795_),
    .B(_06966_),
    .Y(_06974_));
 sg13g2_a22oi_1 _14239_ (.Y(_06975_),
    .B1(_06973_),
    .B2(_06974_),
    .A2(_06885_),
    .A1(_06795_));
 sg13g2_xnor2_1 _14240_ (.Y(_06976_),
    .A(_06967_),
    .B(_06968_));
 sg13g2_nand2_1 _14241_ (.Y(_06977_),
    .A(_06794_),
    .B(_06976_));
 sg13g2_nand2b_1 _14242_ (.Y(_06978_),
    .B(_06977_),
    .A_N(_06975_));
 sg13g2_o21ai_1 _14243_ (.B1(_06977_),
    .Y(_06979_),
    .A1(_06794_),
    .A2(_06840_));
 sg13g2_a21oi_2 _14244_ (.B1(_04813_),
    .Y(_06980_),
    .A2(_06978_),
    .A1(_06972_));
 sg13g2_a21oi_2 _14245_ (.B1(_06972_),
    .Y(_06981_),
    .A2(_06979_),
    .A1(_06975_));
 sg13g2_nor2_1 _14246_ (.A(_06795_),
    .B(_06957_),
    .Y(_06982_));
 sg13g2_xnor2_1 _14247_ (.Y(_06983_),
    .A(_06955_),
    .B(_06982_));
 sg13g2_o21ai_1 _14248_ (.B1(_06980_),
    .Y(_06984_),
    .A1(_06981_),
    .A2(_06983_));
 sg13g2_xor2_1 _14249_ (.B(net418),
    .A(net4313),
    .X(_06985_));
 sg13g2_a21oi_1 _14250_ (.A1(net3652),
    .A2(_06985_),
    .Y(_06986_),
    .B1(net3926));
 sg13g2_a22oi_1 _14251_ (.Y(_00667_),
    .B1(_06984_),
    .B2(_06986_),
    .A2(net3925),
    .A1(_03417_));
 sg13g2_nor2_1 _14252_ (.A(_06795_),
    .B(_06959_),
    .Y(_06987_));
 sg13g2_o21ai_1 _14253_ (.B1(_06987_),
    .Y(_06988_),
    .A1(_06954_),
    .A2(_06958_));
 sg13g2_o21ai_1 _14254_ (.B1(_06988_),
    .Y(_06989_),
    .A1(_06794_),
    .A2(_06948_));
 sg13g2_o21ai_1 _14255_ (.B1(_06980_),
    .Y(_06990_),
    .A1(_06981_),
    .A2(_06989_));
 sg13g2_xor2_1 _14256_ (.B(_04808_),
    .A(_04807_),
    .X(_06991_));
 sg13g2_a21oi_1 _14257_ (.A1(net3652),
    .A2(_06991_),
    .Y(_06992_),
    .B1(net3925));
 sg13g2_a22oi_1 _14258_ (.Y(_00668_),
    .B1(_06990_),
    .B2(_06992_),
    .A2(net3925),
    .A1(_03416_));
 sg13g2_and2_1 _14259_ (.A(_06795_),
    .B(_06937_),
    .X(_06993_));
 sg13g2_xnor2_1 _14260_ (.Y(_06994_),
    .A(_06959_),
    .B(_06960_));
 sg13g2_a21oi_1 _14261_ (.A1(_06794_),
    .A2(_06994_),
    .Y(_06995_),
    .B1(_06993_));
 sg13g2_o21ai_1 _14262_ (.B1(_06980_),
    .Y(_06996_),
    .A1(_06981_),
    .A2(_06995_));
 sg13g2_xnor2_1 _14263_ (.Y(_06997_),
    .A(_04805_),
    .B(_04809_));
 sg13g2_a21oi_1 _14264_ (.A1(net3652),
    .A2(_06997_),
    .Y(_06998_),
    .B1(net3925));
 sg13g2_a22oi_1 _14265_ (.Y(_00669_),
    .B1(_06996_),
    .B2(_06998_),
    .A2(net3926),
    .A1(_03415_));
 sg13g2_xor2_1 _14266_ (.B(_06962_),
    .A(_06961_),
    .X(_06999_));
 sg13g2_nor2_1 _14267_ (.A(_06795_),
    .B(_06999_),
    .Y(_07000_));
 sg13g2_a21oi_1 _14268_ (.A1(_06795_),
    .A2(_06914_),
    .Y(_07001_),
    .B1(_07000_));
 sg13g2_o21ai_1 _14269_ (.B1(_06980_),
    .Y(_07002_),
    .A1(_06981_),
    .A2(_07001_));
 sg13g2_or3_1 _14270_ (.A(_04803_),
    .B(_04804_),
    .C(_04810_),
    .X(_07003_));
 sg13g2_and2_1 _14271_ (.A(_04811_),
    .B(_07003_),
    .X(_07004_));
 sg13g2_a21oi_1 _14272_ (.A1(net3652),
    .A2(_07004_),
    .Y(_07005_),
    .B1(net3925));
 sg13g2_a22oi_1 _14273_ (.Y(_00670_),
    .B1(_07002_),
    .B2(_07005_),
    .A2(net3925),
    .A1(_03414_));
 sg13g2_nand2b_1 _14274_ (.Y(_07006_),
    .B(_06972_),
    .A_N(net3652));
 sg13g2_a21oi_1 _14275_ (.A1(_04802_),
    .A2(_04812_),
    .Y(_07007_),
    .B1(net3925));
 sg13g2_a22oi_1 _14276_ (.Y(_00671_),
    .B1(_07006_),
    .B2(_07007_),
    .A2(net3925),
    .A1(_03413_));
 sg13g2_nand2_1 _14277_ (.Y(_07008_),
    .A(\spiking_network_top_uut.all_data_out[764] ),
    .B(_03667_));
 sg13g2_nor2_1 _14278_ (.A(\spiking_network_top_uut.all_data_out[764] ),
    .B(net3842),
    .Y(_07009_));
 sg13g2_nor2_1 _14279_ (.A(\spiking_network_top_uut.all_data_out[765] ),
    .B(_07009_),
    .Y(_07010_));
 sg13g2_mux2_1 _14280_ (.A0(net3841),
    .A1(net3900),
    .S(\spiking_network_top_uut.all_data_out[764] ),
    .X(_07011_));
 sg13g2_a221oi_1 _14281_ (.B2(\spiking_network_top_uut.all_data_out[765] ),
    .C1(_03515_),
    .B1(_07011_),
    .A1(_07008_),
    .Y(_07012_),
    .A2(_07010_));
 sg13g2_mux4_1 _14282_ (.S0(\spiking_network_top_uut.all_data_out[764] ),
    .A0(net3846),
    .A1(net3845),
    .A2(net3844),
    .A3(net3843),
    .S1(\spiking_network_top_uut.all_data_out[765] ),
    .X(_07013_));
 sg13g2_o21ai_1 _14283_ (.B1(net4549),
    .Y(_07014_),
    .A1(\spiking_network_top_uut.all_data_out[766] ),
    .A2(_07013_));
 sg13g2_nand2_1 _14284_ (.Y(_07015_),
    .A(net3934),
    .B(net404));
 sg13g2_o21ai_1 _14285_ (.B1(_07015_),
    .Y(_00672_),
    .A1(_07012_),
    .A2(_07014_));
 sg13g2_mux2_1 _14286_ (.A0(net479),
    .A1(net404),
    .S(net4548),
    .X(_00673_));
 sg13g2_mux2_1 _14287_ (.A0(net3896),
    .A1(net3895),
    .S(\spiking_network_top_uut.all_data_out[760] ),
    .X(_07016_));
 sg13g2_nor2b_1 _14288_ (.A(\spiking_network_top_uut.all_data_out[760] ),
    .B_N(net3898),
    .Y(_07017_));
 sg13g2_a21oi_1 _14289_ (.A1(\spiking_network_top_uut.all_data_out[760] ),
    .A2(net3897),
    .Y(_07018_),
    .B1(_07017_));
 sg13g2_a21oi_1 _14290_ (.A1(\spiking_network_top_uut.all_data_out[761] ),
    .A2(_07016_),
    .Y(_07019_),
    .B1(\spiking_network_top_uut.all_data_out[762] ));
 sg13g2_o21ai_1 _14291_ (.B1(_07019_),
    .Y(_07020_),
    .A1(\spiking_network_top_uut.all_data_out[761] ),
    .A2(_07018_));
 sg13g2_mux2_1 _14292_ (.A0(net3893),
    .A1(net3892),
    .S(\spiking_network_top_uut.all_data_out[760] ),
    .X(_07021_));
 sg13g2_nand2_1 _14293_ (.Y(_07022_),
    .A(\spiking_network_top_uut.all_data_out[761] ),
    .B(_07021_));
 sg13g2_a21oi_1 _14294_ (.A1(\spiking_network_top_uut.all_data_out[760] ),
    .A2(_03666_),
    .Y(_07023_),
    .B1(\spiking_network_top_uut.all_data_out[761] ));
 sg13g2_o21ai_1 _14295_ (.B1(_07023_),
    .Y(_07024_),
    .A1(\spiking_network_top_uut.all_data_out[760] ),
    .A2(net3894));
 sg13g2_nand3_1 _14296_ (.B(_07022_),
    .C(_07024_),
    .A(\spiking_network_top_uut.all_data_out[762] ),
    .Y(_07025_));
 sg13g2_nand3_1 _14297_ (.B(_07020_),
    .C(_07025_),
    .A(net4545),
    .Y(_07026_));
 sg13g2_o21ai_1 _14298_ (.B1(_07026_),
    .Y(_00674_),
    .A1(net4544),
    .A2(_03676_));
 sg13g2_mux2_1 _14299_ (.A0(net238),
    .A1(net108),
    .S(net4543),
    .X(_00675_));
 sg13g2_mux2_1 _14300_ (.A0(net3889),
    .A1(net3888),
    .S(\spiking_network_top_uut.all_data_out[756] ),
    .X(_07027_));
 sg13g2_nor2b_1 _14301_ (.A(\spiking_network_top_uut.all_data_out[756] ),
    .B_N(net3891),
    .Y(_07028_));
 sg13g2_a21oi_1 _14302_ (.A1(\spiking_network_top_uut.all_data_out[756] ),
    .A2(net3890),
    .Y(_07029_),
    .B1(_07028_));
 sg13g2_a21oi_1 _14303_ (.A1(\spiking_network_top_uut.all_data_out[757] ),
    .A2(_07027_),
    .Y(_07030_),
    .B1(\spiking_network_top_uut.all_data_out[758] ));
 sg13g2_o21ai_1 _14304_ (.B1(_07030_),
    .Y(_07031_),
    .A1(\spiking_network_top_uut.all_data_out[757] ),
    .A2(_07029_));
 sg13g2_mux2_1 _14305_ (.A0(net3886),
    .A1(net3885),
    .S(\spiking_network_top_uut.all_data_out[756] ),
    .X(_07032_));
 sg13g2_nand2_1 _14306_ (.Y(_07033_),
    .A(\spiking_network_top_uut.all_data_out[757] ),
    .B(_07032_));
 sg13g2_a21oi_1 _14307_ (.A1(\spiking_network_top_uut.all_data_out[756] ),
    .A2(_03665_),
    .Y(_07034_),
    .B1(\spiking_network_top_uut.all_data_out[757] ));
 sg13g2_o21ai_1 _14308_ (.B1(_07034_),
    .Y(_07035_),
    .A1(\spiking_network_top_uut.all_data_out[756] ),
    .A2(net3887));
 sg13g2_nand3_1 _14309_ (.B(_07033_),
    .C(_07035_),
    .A(\spiking_network_top_uut.all_data_out[758] ),
    .Y(_07036_));
 sg13g2_nand3_1 _14310_ (.B(_07031_),
    .C(_07036_),
    .A(net4565),
    .Y(_07037_));
 sg13g2_o21ai_1 _14311_ (.B1(_07037_),
    .Y(_00676_),
    .A1(net4561),
    .A2(_03677_));
 sg13g2_mux2_1 _14312_ (.A0(net525),
    .A1(net148),
    .S(net4566),
    .X(_00677_));
 sg13g2_mux4_1 _14313_ (.S0(\spiking_network_top_uut.all_data_out[752] ),
    .A0(net3884),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[1] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[2] ),
    .A3(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[3] ),
    .S1(\spiking_network_top_uut.all_data_out[753] ),
    .X(_07038_));
 sg13g2_mux2_1 _14314_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[6] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[7] ),
    .S(\spiking_network_top_uut.all_data_out[752] ),
    .X(_07039_));
 sg13g2_nor2b_1 _14315_ (.A(\spiking_network_top_uut.all_data_out[752] ),
    .B_N(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[4] ),
    .Y(_07040_));
 sg13g2_a21oi_1 _14316_ (.A1(\spiking_network_top_uut.all_data_out[752] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[5] ),
    .Y(_07041_),
    .B1(_07040_));
 sg13g2_o21ai_1 _14317_ (.B1(\spiking_network_top_uut.all_data_out[754] ),
    .Y(_07042_),
    .A1(\spiking_network_top_uut.all_data_out[753] ),
    .A2(_07041_));
 sg13g2_a21oi_1 _14318_ (.A1(\spiking_network_top_uut.all_data_out[753] ),
    .A2(_07039_),
    .Y(_07043_),
    .B1(_07042_));
 sg13g2_o21ai_1 _14319_ (.B1(net4554),
    .Y(_07044_),
    .A1(\spiking_network_top_uut.all_data_out[754] ),
    .A2(_07038_));
 sg13g2_nand2_1 _14320_ (.Y(_07045_),
    .A(net3938),
    .B(net192));
 sg13g2_o21ai_1 _14321_ (.B1(_07045_),
    .Y(_00678_),
    .A1(_07043_),
    .A2(_07044_));
 sg13g2_mux2_1 _14322_ (.A0(net283),
    .A1(net192),
    .S(net4555),
    .X(_00679_));
 sg13g2_mux4_1 _14323_ (.S0(\spiking_network_top_uut.all_data_out[748] ),
    .A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[0] ),
    .A1(net3875),
    .A2(net3874),
    .A3(net3873),
    .S1(\spiking_network_top_uut.all_data_out[749] ),
    .X(_07046_));
 sg13g2_mux2_1 _14324_ (.A0(net3870),
    .A1(net3869),
    .S(\spiking_network_top_uut.all_data_out[748] ),
    .X(_07047_));
 sg13g2_nor2b_1 _14325_ (.A(\spiking_network_top_uut.all_data_out[748] ),
    .B_N(net3872),
    .Y(_07048_));
 sg13g2_a21oi_1 _14326_ (.A1(\spiking_network_top_uut.all_data_out[748] ),
    .A2(net3871),
    .Y(_07049_),
    .B1(_07048_));
 sg13g2_o21ai_1 _14327_ (.B1(\spiking_network_top_uut.all_data_out[750] ),
    .Y(_07050_),
    .A1(\spiking_network_top_uut.all_data_out[749] ),
    .A2(_07049_));
 sg13g2_a21oi_1 _14328_ (.A1(\spiking_network_top_uut.all_data_out[749] ),
    .A2(_07047_),
    .Y(_07051_),
    .B1(_07050_));
 sg13g2_o21ai_1 _14329_ (.B1(net4566),
    .Y(_07052_),
    .A1(\spiking_network_top_uut.all_data_out[750] ),
    .A2(_07046_));
 sg13g2_nand2_1 _14330_ (.Y(_07053_),
    .A(net3937),
    .B(net121));
 sg13g2_o21ai_1 _14331_ (.B1(_07053_),
    .Y(_00680_),
    .A1(_07051_),
    .A2(_07052_));
 sg13g2_mux2_1 _14332_ (.A0(net280),
    .A1(net121),
    .S(net4568),
    .X(_00681_));
 sg13g2_mux4_1 _14333_ (.S0(\spiking_network_top_uut.all_data_out[744] ),
    .A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[0] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[1] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[2] ),
    .A3(net3865),
    .S1(\spiking_network_top_uut.all_data_out[745] ),
    .X(_07054_));
 sg13g2_mux2_1 _14334_ (.A0(net3862),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[7] ),
    .S(\spiking_network_top_uut.all_data_out[744] ),
    .X(_07055_));
 sg13g2_nor2b_1 _14335_ (.A(\spiking_network_top_uut.all_data_out[744] ),
    .B_N(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[4] ),
    .Y(_07056_));
 sg13g2_a21oi_1 _14336_ (.A1(\spiking_network_top_uut.all_data_out[744] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[5] ),
    .Y(_07057_),
    .B1(_07056_));
 sg13g2_o21ai_1 _14337_ (.B1(\spiking_network_top_uut.all_data_out[746] ),
    .Y(_07058_),
    .A1(\spiking_network_top_uut.all_data_out[745] ),
    .A2(_07057_));
 sg13g2_a21oi_1 _14338_ (.A1(\spiking_network_top_uut.all_data_out[745] ),
    .A2(_07055_),
    .Y(_07059_),
    .B1(_07058_));
 sg13g2_o21ai_1 _14339_ (.B1(net4564),
    .Y(_07060_),
    .A1(\spiking_network_top_uut.all_data_out[746] ),
    .A2(_07054_));
 sg13g2_nand2_1 _14340_ (.Y(_07061_),
    .A(net3935),
    .B(net383));
 sg13g2_o21ai_1 _14341_ (.B1(_07061_),
    .Y(_00682_),
    .A1(_07059_),
    .A2(_07060_));
 sg13g2_mux2_1 _14342_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_dout ),
    .A1(net383),
    .S(net4570),
    .X(_00683_));
 sg13g2_mux2_1 _14343_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[2] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[3] ),
    .S(\spiking_network_top_uut.all_data_out[740] ),
    .X(_07062_));
 sg13g2_nor2b_1 _14344_ (.A(\spiking_network_top_uut.all_data_out[740] ),
    .B_N(net3860),
    .Y(_07063_));
 sg13g2_a21oi_1 _14345_ (.A1(\spiking_network_top_uut.all_data_out[740] ),
    .A2(net3859),
    .Y(_07064_),
    .B1(_07063_));
 sg13g2_a21oi_1 _14346_ (.A1(\spiking_network_top_uut.all_data_out[741] ),
    .A2(_07062_),
    .Y(_07065_),
    .B1(\spiking_network_top_uut.all_data_out[742] ));
 sg13g2_o21ai_1 _14347_ (.B1(_07065_),
    .Y(_07066_),
    .A1(\spiking_network_top_uut.all_data_out[741] ),
    .A2(_07064_));
 sg13g2_mux2_1 _14348_ (.A0(net3855),
    .A1(net3854),
    .S(\spiking_network_top_uut.all_data_out[740] ),
    .X(_07067_));
 sg13g2_nand2_1 _14349_ (.Y(_07068_),
    .A(\spiking_network_top_uut.all_data_out[741] ),
    .B(_07067_));
 sg13g2_a21oi_1 _14350_ (.A1(\spiking_network_top_uut.all_data_out[740] ),
    .A2(_03664_),
    .Y(_07069_),
    .B1(\spiking_network_top_uut.all_data_out[741] ));
 sg13g2_o21ai_1 _14351_ (.B1(_07069_),
    .Y(_07070_),
    .A1(\spiking_network_top_uut.all_data_out[740] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[4] ));
 sg13g2_nand3_1 _14352_ (.B(_07068_),
    .C(_07070_),
    .A(\spiking_network_top_uut.all_data_out[742] ),
    .Y(_07071_));
 sg13g2_nand3_1 _14353_ (.B(_07066_),
    .C(_07071_),
    .A(net4535),
    .Y(_07072_));
 sg13g2_o21ai_1 _14354_ (.B1(_07072_),
    .Y(_00684_),
    .A1(net4535),
    .A2(_03678_));
 sg13g2_mux2_1 _14355_ (.A0(net202),
    .A1(net115),
    .S(net4535),
    .X(_00685_));
 sg13g2_mux4_1 _14356_ (.S0(\spiking_network_top_uut.all_data_out[736] ),
    .A0(net3853),
    .A1(net3852),
    .A2(net3851),
    .A3(net3850),
    .S1(\spiking_network_top_uut.all_data_out[737] ),
    .X(_07073_));
 sg13g2_mux2_1 _14357_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[6] ),
    .A1(net3847),
    .S(\spiking_network_top_uut.all_data_out[736] ),
    .X(_07074_));
 sg13g2_nor2b_1 _14358_ (.A(\spiking_network_top_uut.all_data_out[736] ),
    .B_N(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[4] ),
    .Y(_07075_));
 sg13g2_a21oi_1 _14359_ (.A1(\spiking_network_top_uut.all_data_out[736] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[5] ),
    .Y(_07076_),
    .B1(_07075_));
 sg13g2_o21ai_1 _14360_ (.B1(\spiking_network_top_uut.all_data_out[738] ),
    .Y(_07077_),
    .A1(\spiking_network_top_uut.all_data_out[737] ),
    .A2(_07076_));
 sg13g2_a21oi_1 _14361_ (.A1(\spiking_network_top_uut.all_data_out[737] ),
    .A2(_07074_),
    .Y(_07078_),
    .B1(_07077_));
 sg13g2_o21ai_1 _14362_ (.B1(net4544),
    .Y(_07079_),
    .A1(\spiking_network_top_uut.all_data_out[738] ),
    .A2(_07073_));
 sg13g2_nand2_1 _14363_ (.Y(_07080_),
    .A(net3933),
    .B(net389));
 sg13g2_o21ai_1 _14364_ (.B1(_07080_),
    .Y(_00686_),
    .A1(_07078_),
    .A2(_07079_));
 sg13g2_nor3_2 _14365_ (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[2] ),
    .B(net557),
    .C(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[0] ),
    .Y(_07081_));
 sg13g2_nor2b_2 _14366_ (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[3] ),
    .B_N(_07081_),
    .Y(_07082_));
 sg13g2_nor2b_2 _14367_ (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[4] ),
    .B_N(_07082_),
    .Y(_07083_));
 sg13g2_nand2b_2 _14368_ (.Y(_07084_),
    .B(_07082_),
    .A_N(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[4] ));
 sg13g2_o21ai_1 _14369_ (.B1(net4531),
    .Y(_07085_),
    .A1(net3648),
    .A2(_07084_));
 sg13g2_nor2b_1 _14370_ (.A(net3648),
    .B_N(_00078_),
    .Y(_07086_));
 sg13g2_a21oi_1 _14371_ (.A1(net4284),
    .A2(net3648),
    .Y(_07087_),
    .B1(_07086_));
 sg13g2_nand2_1 _14372_ (.Y(_07088_),
    .A(net353),
    .B(_07085_));
 sg13g2_o21ai_1 _14373_ (.B1(_07088_),
    .Y(_00687_),
    .A1(_07085_),
    .A2(_07087_));
 sg13g2_xor2_1 _14374_ (.B(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[0] ),
    .A(net323),
    .X(_07089_));
 sg13g2_nor2_1 _14375_ (.A(net3648),
    .B(_07089_),
    .Y(_07090_));
 sg13g2_a21oi_1 _14376_ (.A1(net4281),
    .A2(net3648),
    .Y(_07091_),
    .B1(_07090_));
 sg13g2_nand2_1 _14377_ (.Y(_07092_),
    .A(net323),
    .B(_07085_));
 sg13g2_o21ai_1 _14378_ (.B1(_07092_),
    .Y(_00688_),
    .A1(_07085_),
    .A2(_07091_));
 sg13g2_o21ai_1 _14379_ (.B1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[2] ),
    .Y(_07093_),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[1] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[0] ));
 sg13g2_nor2b_1 _14380_ (.A(_07081_),
    .B_N(_07093_),
    .Y(_07094_));
 sg13g2_nor2_1 _14381_ (.A(net3648),
    .B(_07094_),
    .Y(_07095_));
 sg13g2_a21oi_1 _14382_ (.A1(net4277),
    .A2(net3648),
    .Y(_07096_),
    .B1(_07095_));
 sg13g2_nand2_1 _14383_ (.Y(_07097_),
    .A(net183),
    .B(_07085_));
 sg13g2_o21ai_1 _14384_ (.B1(_07097_),
    .Y(_00689_),
    .A1(_07085_),
    .A2(_07096_));
 sg13g2_nand2_1 _14385_ (.Y(_07098_),
    .A(net4274),
    .B(net3648));
 sg13g2_xnor2_1 _14386_ (.Y(_07099_),
    .A(net428),
    .B(_07081_));
 sg13g2_o21ai_1 _14387_ (.B1(_07098_),
    .Y(_07100_),
    .A1(net3649),
    .A2(_07099_));
 sg13g2_mux2_1 _14388_ (.A0(_07100_),
    .A1(net428),
    .S(_07085_),
    .X(_00690_));
 sg13g2_nand2_1 _14389_ (.Y(_07101_),
    .A(net3924),
    .B(net295));
 sg13g2_nand2b_1 _14390_ (.Y(_07102_),
    .B(net295),
    .A_N(_07082_));
 sg13g2_a21oi_1 _14391_ (.A1(_07084_),
    .A2(_07102_),
    .Y(_07103_),
    .B1(net3649));
 sg13g2_a21oi_1 _14392_ (.A1(net4270),
    .A2(net3649),
    .Y(_07104_),
    .B1(_07103_));
 sg13g2_o21ai_1 _14393_ (.B1(_07101_),
    .Y(_00691_),
    .A1(_07085_),
    .A2(_07104_));
 sg13g2_mux2_1 _14394_ (.A0(net291),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_reg1 ),
    .S(net4542),
    .X(_00692_));
 sg13g2_nor2_1 _14395_ (.A(_00073_),
    .B(net3741),
    .Y(_07105_));
 sg13g2_nor3_2 _14396_ (.A(_00073_),
    .B(net3748),
    .C(_05090_),
    .Y(_07106_));
 sg13g2_nand2_1 _14397_ (.Y(_07107_),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ),
    .B(_00073_));
 sg13g2_a21oi_1 _14398_ (.A1(net3917),
    .A2(net3741),
    .Y(_07108_),
    .B1(_00073_));
 sg13g2_nor2b_1 _14399_ (.A(_07108_),
    .B_N(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ),
    .Y(_07109_));
 sg13g2_nand2_1 _14400_ (.Y(_07110_),
    .A(_00074_),
    .B(net3749));
 sg13g2_o21ai_1 _14401_ (.B1(_07110_),
    .Y(_07111_),
    .A1(net3748),
    .A2(_07105_));
 sg13g2_nor2_1 _14402_ (.A(_00074_),
    .B(net3906),
    .Y(_07112_));
 sg13g2_a221oi_1 _14403_ (.B2(_07105_),
    .C1(_07112_),
    .B1(net3906),
    .A1(_03484_),
    .Y(_07113_),
    .A2(net3748));
 sg13g2_nand2_1 _14404_ (.Y(_07114_),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ),
    .B(_07113_));
 sg13g2_nor2_1 _14405_ (.A(_00074_),
    .B(_05105_),
    .Y(_07115_));
 sg13g2_nor2_1 _14406_ (.A(_00073_),
    .B(net3910),
    .Y(_07116_));
 sg13g2_o21ai_1 _14407_ (.B1(net3917),
    .Y(_07117_),
    .A1(_00075_),
    .A2(net3906));
 sg13g2_nor3_2 _14408_ (.A(_07115_),
    .B(_07116_),
    .C(_07117_),
    .Y(_07118_));
 sg13g2_and2_1 _14409_ (.A(_00077_),
    .B(net3748),
    .X(_07119_));
 sg13g2_nor3_2 _14410_ (.A(_03485_),
    .B(_07118_),
    .C(_07119_),
    .Y(_07120_));
 sg13g2_xnor2_1 _14411_ (.Y(_07121_),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ),
    .B(_07113_));
 sg13g2_o21ai_1 _14412_ (.B1(_07114_),
    .Y(_07122_),
    .A1(_07120_),
    .A2(_07121_));
 sg13g2_xnor2_1 _14413_ (.Y(_07123_),
    .A(_03484_),
    .B(_07111_));
 sg13g2_nor2b_1 _14414_ (.A(_07123_),
    .B_N(_07122_),
    .Y(_07124_));
 sg13g2_a21o_1 _14415_ (.A2(_07111_),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ),
    .B1(_07124_),
    .X(_07125_));
 sg13g2_xnor2_1 _14416_ (.Y(_07126_),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ),
    .B(_07108_));
 sg13g2_a21oi_1 _14417_ (.A1(_07125_),
    .A2(_07126_),
    .Y(_07127_),
    .B1(_07109_));
 sg13g2_nor2b_1 _14418_ (.A(_07106_),
    .B_N(_07127_),
    .Y(_07128_));
 sg13g2_a22oi_1 _14419_ (.Y(_07129_),
    .B1(_07107_),
    .B2(_07128_),
    .A2(_07106_),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ));
 sg13g2_and2_1 _14420_ (.A(_07084_),
    .B(_07129_),
    .X(_07130_));
 sg13g2_mux2_2 _14421_ (.A0(net4599),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[739] ),
    .X(_07131_));
 sg13g2_nand2_1 _14422_ (.Y(_07132_),
    .A(\spiking_network_top_uut.all_data_out[241] ),
    .B(_07131_));
 sg13g2_mux2_1 _14423_ (.A0(net4598),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[743] ),
    .X(_07133_));
 sg13g2_nand2_1 _14424_ (.Y(_07134_),
    .A(\spiking_network_top_uut.all_data_out[243] ),
    .B(_07133_));
 sg13g2_nor2_1 _14425_ (.A(_07132_),
    .B(_07134_),
    .Y(_07135_));
 sg13g2_nand4_1 _14426_ (.B(\spiking_network_top_uut.all_data_out[242] ),
    .C(_07131_),
    .A(\spiking_network_top_uut.all_data_out[240] ),
    .Y(_07136_),
    .D(_07133_));
 sg13g2_inv_1 _14427_ (.Y(_07137_),
    .A(_07136_));
 sg13g2_xor2_1 _14428_ (.B(_07134_),
    .A(_07132_),
    .X(_07138_));
 sg13g2_a21oi_2 _14429_ (.B1(_07135_),
    .Y(_07139_),
    .A2(_07138_),
    .A1(_07136_));
 sg13g2_mux2_2 _14430_ (.A0(net4597),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[747] ),
    .X(_07140_));
 sg13g2_nand2_1 _14431_ (.Y(_07141_),
    .A(\spiking_network_top_uut.all_data_out[245] ),
    .B(_07140_));
 sg13g2_mux2_2 _14432_ (.A0(net4596),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[751] ),
    .X(_07142_));
 sg13g2_nand2_2 _14433_ (.Y(_07143_),
    .A(\spiking_network_top_uut.all_data_out[247] ),
    .B(_07142_));
 sg13g2_nor2_1 _14434_ (.A(_07141_),
    .B(_07143_),
    .Y(_07144_));
 sg13g2_nand2_1 _14435_ (.Y(_07145_),
    .A(\spiking_network_top_uut.all_data_out[244] ),
    .B(_07140_));
 sg13g2_nand2_2 _14436_ (.Y(_07146_),
    .A(\spiking_network_top_uut.all_data_out[246] ),
    .B(_07142_));
 sg13g2_or2_1 _14437_ (.X(_07147_),
    .B(_07146_),
    .A(_07145_));
 sg13g2_xor2_1 _14438_ (.B(_07143_),
    .A(_07141_),
    .X(_07148_));
 sg13g2_a21oi_2 _14439_ (.B1(_07144_),
    .Y(_07149_),
    .A2(_07148_),
    .A1(_07147_));
 sg13g2_mux2_2 _14440_ (.A0(net4595),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[755] ),
    .X(_07150_));
 sg13g2_mux2_2 _14441_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.spike_out ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[759] ),
    .X(_07151_));
 sg13g2_a22oi_1 _14442_ (.Y(_07152_),
    .B1(_07151_),
    .B2(\spiking_network_top_uut.all_data_out[251] ),
    .A2(_07150_),
    .A1(\spiking_network_top_uut.all_data_out[249] ));
 sg13g2_and4_1 _14443_ (.A(\spiking_network_top_uut.all_data_out[249] ),
    .B(\spiking_network_top_uut.all_data_out[251] ),
    .C(_07150_),
    .D(_07151_),
    .X(_07153_));
 sg13g2_nand4_1 _14444_ (.B(\spiking_network_top_uut.all_data_out[251] ),
    .C(_07150_),
    .A(\spiking_network_top_uut.all_data_out[249] ),
    .Y(_07154_),
    .D(_07151_));
 sg13g2_and4_2 _14445_ (.A(\spiking_network_top_uut.all_data_out[248] ),
    .B(\spiking_network_top_uut.all_data_out[250] ),
    .C(_07150_),
    .D(_07151_),
    .X(_07155_));
 sg13g2_a21oi_2 _14446_ (.B1(_07152_),
    .Y(_07156_),
    .A2(_07155_),
    .A1(_07154_));
 sg13g2_mux2_2 _14447_ (.A0(net4593),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[763] ),
    .X(_07157_));
 sg13g2_mux2_2 _14448_ (.A0(net4592),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[767] ),
    .X(_07158_));
 sg13g2_and4_1 _14449_ (.A(\spiking_network_top_uut.all_data_out[253] ),
    .B(\spiking_network_top_uut.all_data_out[255] ),
    .C(_07157_),
    .D(_07158_),
    .X(_07159_));
 sg13g2_nand4_1 _14450_ (.B(\spiking_network_top_uut.all_data_out[255] ),
    .C(_07157_),
    .A(\spiking_network_top_uut.all_data_out[253] ),
    .Y(_07160_),
    .D(_07158_));
 sg13g2_and4_1 _14451_ (.A(\spiking_network_top_uut.all_data_out[252] ),
    .B(\spiking_network_top_uut.all_data_out[254] ),
    .C(_07157_),
    .D(_07158_),
    .X(_07161_));
 sg13g2_a22oi_1 _14452_ (.Y(_07162_),
    .B1(_07158_),
    .B2(\spiking_network_top_uut.all_data_out[255] ),
    .A2(_07157_),
    .A1(\spiking_network_top_uut.all_data_out[253] ));
 sg13g2_or3_1 _14453_ (.A(_07159_),
    .B(_07161_),
    .C(_07162_),
    .X(_07163_));
 sg13g2_o21ai_1 _14454_ (.B1(_07160_),
    .Y(_07164_),
    .A1(_07161_),
    .A2(_07162_));
 sg13g2_nand3b_1 _14455_ (.B(_07156_),
    .C(_07164_),
    .Y(_07165_),
    .A_N(_07149_));
 sg13g2_inv_1 _14456_ (.Y(_07166_),
    .A(_07165_));
 sg13g2_or2_1 _14457_ (.X(_07167_),
    .B(_07165_),
    .A(_07139_));
 sg13g2_inv_2 _14458_ (.Y(_07168_),
    .A(_07167_));
 sg13g2_nor2_1 _14459_ (.A(_07156_),
    .B(_07164_),
    .Y(_07169_));
 sg13g2_and2_2 _14460_ (.A(_07149_),
    .B(_07169_),
    .X(_07170_));
 sg13g2_a21oi_2 _14461_ (.B1(_07168_),
    .Y(_07171_),
    .A2(_07170_),
    .A1(_07139_));
 sg13g2_xor2_1 _14462_ (.B(_07127_),
    .A(_07106_),
    .X(_07172_));
 sg13g2_a21o_1 _14463_ (.A2(_07172_),
    .A1(_07171_),
    .B1(_07168_),
    .X(_07173_));
 sg13g2_nor2b_1 _14464_ (.A(_07171_),
    .B_N(_07129_),
    .Y(_07174_));
 sg13g2_xor2_1 _14465_ (.B(_07171_),
    .A(_07129_),
    .X(_07175_));
 sg13g2_nor2b_1 _14466_ (.A(_07175_),
    .B_N(_07173_),
    .Y(_07176_));
 sg13g2_xnor2_1 _14467_ (.Y(_07177_),
    .A(_07173_),
    .B(_07175_));
 sg13g2_o21ai_1 _14468_ (.B1(_07161_),
    .Y(_07178_),
    .A1(_07159_),
    .A2(_07162_));
 sg13g2_o21ai_1 _14469_ (.B1(_07155_),
    .Y(_07179_),
    .A1(_07152_),
    .A2(_07153_));
 sg13g2_or3_1 _14470_ (.A(_07152_),
    .B(_07153_),
    .C(_07155_),
    .X(_07180_));
 sg13g2_a22oi_1 _14471_ (.Y(_07181_),
    .B1(_07179_),
    .B2(_07180_),
    .A2(_07178_),
    .A1(_07163_));
 sg13g2_xor2_1 _14472_ (.B(_07148_),
    .A(_07147_),
    .X(_07182_));
 sg13g2_xnor2_1 _14473_ (.Y(_07183_),
    .A(_07147_),
    .B(_07148_));
 sg13g2_and4_1 _14474_ (.A(_07163_),
    .B(_07178_),
    .C(_07179_),
    .D(_07180_),
    .X(_07184_));
 sg13g2_nand4_1 _14475_ (.B(_07178_),
    .C(_07179_),
    .A(_07163_),
    .Y(_07185_),
    .D(_07180_));
 sg13g2_nand3b_1 _14476_ (.B(_07183_),
    .C(_07185_),
    .Y(_07186_),
    .A_N(_07181_));
 sg13g2_a21oi_2 _14477_ (.B1(_07181_),
    .Y(_07187_),
    .A2(_07185_),
    .A1(_07183_));
 sg13g2_xor2_1 _14478_ (.B(_07164_),
    .A(_07156_),
    .X(_07188_));
 sg13g2_xnor2_1 _14479_ (.Y(_07189_),
    .A(_07149_),
    .B(_07188_));
 sg13g2_nor2b_1 _14480_ (.A(_07187_),
    .B_N(_07189_),
    .Y(_07190_));
 sg13g2_xnor2_1 _14481_ (.Y(_07191_),
    .A(_07187_),
    .B(_07189_));
 sg13g2_nor2b_1 _14482_ (.A(_07139_),
    .B_N(_07191_),
    .Y(_07192_));
 sg13g2_nor2_2 _14483_ (.A(_07190_),
    .B(_07192_),
    .Y(_07193_));
 sg13g2_nor2_1 _14484_ (.A(_07166_),
    .B(_07170_),
    .Y(_07194_));
 sg13g2_xnor2_1 _14485_ (.Y(_07195_),
    .A(_07139_),
    .B(_07194_));
 sg13g2_nor2b_1 _14486_ (.A(_07193_),
    .B_N(_07195_),
    .Y(_07196_));
 sg13g2_xnor2_1 _14487_ (.Y(_07197_),
    .A(_07193_),
    .B(_07195_));
 sg13g2_xor2_1 _14488_ (.B(_07126_),
    .A(_07125_),
    .X(_07198_));
 sg13g2_a21oi_1 _14489_ (.A1(_07197_),
    .A2(_07198_),
    .Y(_07199_),
    .B1(_07196_));
 sg13g2_xor2_1 _14490_ (.B(_07172_),
    .A(_07171_),
    .X(_07200_));
 sg13g2_nand2b_1 _14491_ (.Y(_07201_),
    .B(_07200_),
    .A_N(_07199_));
 sg13g2_xnor2_1 _14492_ (.Y(_07202_),
    .A(_07197_),
    .B(_07198_));
 sg13g2_a22oi_1 _14493_ (.Y(_07203_),
    .B1(_07158_),
    .B2(\spiking_network_top_uut.all_data_out[254] ),
    .A2(_07157_),
    .A1(\spiking_network_top_uut.all_data_out[252] ));
 sg13g2_nor2_1 _14494_ (.A(_07161_),
    .B(_07203_),
    .Y(_07204_));
 sg13g2_a22oi_1 _14495_ (.Y(_07205_),
    .B1(_07151_),
    .B2(\spiking_network_top_uut.all_data_out[250] ),
    .A2(_07150_),
    .A1(\spiking_network_top_uut.all_data_out[248] ));
 sg13g2_nor2_1 _14496_ (.A(_07155_),
    .B(_07205_),
    .Y(_07206_));
 sg13g2_and2_1 _14497_ (.A(_07204_),
    .B(_07206_),
    .X(_07207_));
 sg13g2_xor2_1 _14498_ (.B(_07146_),
    .A(_07145_),
    .X(_07208_));
 sg13g2_xor2_1 _14499_ (.B(_07206_),
    .A(_07204_),
    .X(_07209_));
 sg13g2_a21o_2 _14500_ (.A2(_07209_),
    .A1(_07208_),
    .B1(_07207_),
    .X(_07210_));
 sg13g2_o21ai_1 _14501_ (.B1(_07182_),
    .Y(_07211_),
    .A1(_07181_),
    .A2(_07184_));
 sg13g2_and3_1 _14502_ (.X(_07212_),
    .A(_07186_),
    .B(_07210_),
    .C(_07211_));
 sg13g2_nand3_1 _14503_ (.B(_07210_),
    .C(_07211_),
    .A(_07186_),
    .Y(_07213_));
 sg13g2_xnor2_1 _14504_ (.Y(_07214_),
    .A(_07137_),
    .B(_07138_));
 sg13g2_a21oi_1 _14505_ (.A1(_07186_),
    .A2(_07211_),
    .Y(_07215_),
    .B1(_07210_));
 sg13g2_or3_2 _14506_ (.A(_07212_),
    .B(_07214_),
    .C(_07215_),
    .X(_07216_));
 sg13g2_o21ai_1 _14507_ (.B1(_07213_),
    .Y(_07217_),
    .A1(_07214_),
    .A2(_07215_));
 sg13g2_xnor2_1 _14508_ (.Y(_07218_),
    .A(_07139_),
    .B(_07191_));
 sg13g2_nand2_2 _14509_ (.Y(_07219_),
    .A(_07217_),
    .B(_07218_));
 sg13g2_xnor2_1 _14510_ (.Y(_07220_),
    .A(_07217_),
    .B(_07218_));
 sg13g2_xor2_1 _14511_ (.B(_07123_),
    .A(_07122_),
    .X(_07221_));
 sg13g2_o21ai_1 _14512_ (.B1(_07219_),
    .Y(_07222_),
    .A1(_07220_),
    .A2(_07221_));
 sg13g2_nor2b_1 _14513_ (.A(_07202_),
    .B_N(_07222_),
    .Y(_07223_));
 sg13g2_xor2_1 _14514_ (.B(_07221_),
    .A(_07220_),
    .X(_07224_));
 sg13g2_a22oi_1 _14515_ (.Y(_07225_),
    .B1(_07133_),
    .B2(\spiking_network_top_uut.all_data_out[242] ),
    .A2(_07131_),
    .A1(\spiking_network_top_uut.all_data_out[240] ));
 sg13g2_nor2_2 _14516_ (.A(_07137_),
    .B(_07225_),
    .Y(_07226_));
 sg13g2_inv_1 _14517_ (.Y(_07227_),
    .A(_07226_));
 sg13g2_xnor2_1 _14518_ (.Y(_07228_),
    .A(_07208_),
    .B(_07209_));
 sg13g2_nor2_2 _14519_ (.A(_07227_),
    .B(_07228_),
    .Y(_07229_));
 sg13g2_o21ai_1 _14520_ (.B1(_07214_),
    .Y(_07230_),
    .A1(_07212_),
    .A2(_07215_));
 sg13g2_and3_1 _14521_ (.X(_07231_),
    .A(_07216_),
    .B(_07229_),
    .C(_07230_));
 sg13g2_nand3_1 _14522_ (.B(_07229_),
    .C(_07230_),
    .A(_07216_),
    .Y(_07232_));
 sg13g2_a21oi_1 _14523_ (.A1(_07216_),
    .A2(_07230_),
    .Y(_07233_),
    .B1(_07229_));
 sg13g2_xnor2_1 _14524_ (.Y(_07234_),
    .A(_07120_),
    .B(_07121_));
 sg13g2_nor3_1 _14525_ (.A(_07231_),
    .B(_07233_),
    .C(_07234_),
    .Y(_07235_));
 sg13g2_o21ai_1 _14526_ (.B1(_07232_),
    .Y(_07236_),
    .A1(_07233_),
    .A2(_07234_));
 sg13g2_nand2_1 _14527_ (.Y(_07237_),
    .A(_07224_),
    .B(_07236_));
 sg13g2_o21ai_1 _14528_ (.B1(_07234_),
    .Y(_07238_),
    .A1(_07231_),
    .A2(_07233_));
 sg13g2_nand2b_1 _14529_ (.Y(_07239_),
    .B(_07238_),
    .A_N(_07235_));
 sg13g2_xnor2_1 _14530_ (.Y(_07240_),
    .A(_07227_),
    .B(_07228_));
 sg13g2_o21ai_1 _14531_ (.B1(_03485_),
    .Y(_07241_),
    .A1(_07118_),
    .A2(_07119_));
 sg13g2_nor2b_1 _14532_ (.A(_07120_),
    .B_N(_07241_),
    .Y(_07242_));
 sg13g2_nor2_1 _14533_ (.A(_07240_),
    .B(_07242_),
    .Y(_07243_));
 sg13g2_nand3b_1 _14534_ (.B(_07238_),
    .C(_07243_),
    .Y(_07244_),
    .A_N(_07235_));
 sg13g2_nor2_1 _14535_ (.A(_07224_),
    .B(_07236_),
    .Y(_07245_));
 sg13g2_xor2_1 _14536_ (.B(_07236_),
    .A(_07224_),
    .X(_07246_));
 sg13g2_o21ai_1 _14537_ (.B1(_07237_),
    .Y(_07247_),
    .A1(_07244_),
    .A2(_07245_));
 sg13g2_nand2b_1 _14538_ (.Y(_07248_),
    .B(_07202_),
    .A_N(_07222_));
 sg13g2_nand2b_1 _14539_ (.Y(_07249_),
    .B(_07248_),
    .A_N(_07223_));
 sg13g2_a21oi_1 _14540_ (.A1(_07247_),
    .A2(_07248_),
    .Y(_07250_),
    .B1(_07223_));
 sg13g2_xor2_1 _14541_ (.B(_07200_),
    .A(_07199_),
    .X(_07251_));
 sg13g2_o21ai_1 _14542_ (.B1(_07201_),
    .Y(_07252_),
    .A1(_07250_),
    .A2(_07251_));
 sg13g2_a21oi_1 _14543_ (.A1(_07177_),
    .A2(_07252_),
    .Y(_07253_),
    .B1(_07176_));
 sg13g2_nand2_1 _14544_ (.Y(_07254_),
    .A(_07129_),
    .B(_07168_));
 sg13g2_o21ai_1 _14545_ (.B1(_07254_),
    .Y(_07255_),
    .A1(_07168_),
    .A2(_07174_));
 sg13g2_xor2_1 _14546_ (.B(_07255_),
    .A(_07253_),
    .X(_07256_));
 sg13g2_a21oi_2 _14547_ (.B1(_07130_),
    .Y(_07257_),
    .A2(_07256_),
    .A1(_07083_));
 sg13g2_xnor2_1 _14548_ (.Y(_07258_),
    .A(_07177_),
    .B(_07252_));
 sg13g2_a21o_1 _14549_ (.A2(_07258_),
    .A1(_07083_),
    .B1(_07130_),
    .X(_07259_));
 sg13g2_xnor2_1 _14550_ (.Y(_07260_),
    .A(_07250_),
    .B(_07251_));
 sg13g2_nor2_1 _14551_ (.A(_07084_),
    .B(_07260_),
    .Y(_07261_));
 sg13g2_a21oi_1 _14552_ (.A1(_07084_),
    .A2(_07172_),
    .Y(_07262_),
    .B1(_07261_));
 sg13g2_or2_1 _14553_ (.X(_07263_),
    .B(_07262_),
    .A(_07259_));
 sg13g2_a21o_1 _14554_ (.A2(_07263_),
    .A1(_07257_),
    .B1(net3650),
    .X(_07264_));
 sg13g2_or2_1 _14555_ (.X(_07265_),
    .B(_07264_),
    .A(net3926));
 sg13g2_a21o_1 _14556_ (.A2(_07262_),
    .A1(_07259_),
    .B1(_07257_),
    .X(_07266_));
 sg13g2_nor2_1 _14557_ (.A(_07084_),
    .B(_07240_),
    .Y(_07267_));
 sg13g2_xor2_1 _14558_ (.B(_07267_),
    .A(_07242_),
    .X(_07268_));
 sg13g2_and2_1 _14559_ (.A(_07266_),
    .B(_07268_),
    .X(_07269_));
 sg13g2_xor2_1 _14560_ (.B(net459),
    .A(net4314),
    .X(_07270_));
 sg13g2_a22oi_1 _14561_ (.Y(_07271_),
    .B1(_00014_),
    .B2(_07270_),
    .A2(net459),
    .A1(net3926));
 sg13g2_o21ai_1 _14562_ (.B1(_07271_),
    .Y(_00693_),
    .A1(_07265_),
    .A2(_07269_));
 sg13g2_xnor2_1 _14563_ (.Y(_07272_),
    .A(_07239_),
    .B(_07243_));
 sg13g2_nor2_1 _14564_ (.A(_07083_),
    .B(_07234_),
    .Y(_07273_));
 sg13g2_a21oi_1 _14565_ (.A1(_07083_),
    .A2(_07272_),
    .Y(_07274_),
    .B1(_07273_));
 sg13g2_a21o_1 _14566_ (.A2(_07274_),
    .A1(_07266_),
    .B1(_07264_),
    .X(_07275_));
 sg13g2_xor2_1 _14567_ (.B(_04821_),
    .A(_04820_),
    .X(_07276_));
 sg13g2_a21oi_1 _14568_ (.A1(net3650),
    .A2(_07276_),
    .Y(_07277_),
    .B1(net3927));
 sg13g2_a22oi_1 _14569_ (.Y(_00694_),
    .B1(_07275_),
    .B2(_07277_),
    .A2(_03420_),
    .A1(net3926));
 sg13g2_nand2_1 _14570_ (.Y(_07278_),
    .A(_07084_),
    .B(_07221_));
 sg13g2_xnor2_1 _14571_ (.Y(_07279_),
    .A(_07244_),
    .B(_07246_));
 sg13g2_o21ai_1 _14572_ (.B1(_07278_),
    .Y(_07280_),
    .A1(_07084_),
    .A2(_07279_));
 sg13g2_and2_1 _14573_ (.A(_07266_),
    .B(_07280_),
    .X(_07281_));
 sg13g2_xor2_1 _14574_ (.B(_04823_),
    .A(_04822_),
    .X(_07282_));
 sg13g2_a22oi_1 _14575_ (.Y(_07283_),
    .B1(_00014_),
    .B2(_07282_),
    .A2(net483),
    .A1(net3926));
 sg13g2_o21ai_1 _14576_ (.B1(_07283_),
    .Y(_00695_),
    .A1(_07265_),
    .A2(_07281_));
 sg13g2_nor2_1 _14577_ (.A(_07083_),
    .B(_07198_),
    .Y(_07284_));
 sg13g2_xor2_1 _14578_ (.B(_07249_),
    .A(_07247_),
    .X(_07285_));
 sg13g2_a21oi_1 _14579_ (.A1(_07083_),
    .A2(_07285_),
    .Y(_07286_),
    .B1(_07284_));
 sg13g2_nor2b_1 _14580_ (.A(_07286_),
    .B_N(_07266_),
    .Y(_07287_));
 sg13g2_or3_1 _14581_ (.A(_04817_),
    .B(_04818_),
    .C(_04824_),
    .X(_07288_));
 sg13g2_and2_1 _14582_ (.A(_04825_),
    .B(_07288_),
    .X(_07289_));
 sg13g2_a22oi_1 _14583_ (.Y(_07290_),
    .B1(_00014_),
    .B2(_07289_),
    .A2(net498),
    .A1(net3926));
 sg13g2_o21ai_1 _14584_ (.B1(_07290_),
    .Y(_00696_),
    .A1(_07265_),
    .A2(_07287_));
 sg13g2_o21ai_1 _14585_ (.B1(net4532),
    .Y(_07291_),
    .A1(_04815_),
    .A2(_04826_));
 sg13g2_a21oi_1 _14586_ (.A1(_04828_),
    .A2(_07257_),
    .Y(_07292_),
    .B1(_07291_));
 sg13g2_a21oi_1 _14587_ (.A1(net3927),
    .A2(_03419_),
    .Y(_00697_),
    .B1(_07292_));
 sg13g2_a21oi_1 _14588_ (.A1(\spiking_network_top_uut.all_data_out[796] ),
    .A2(_03667_),
    .Y(_07293_),
    .B1(\spiking_network_top_uut.all_data_out[797] ));
 sg13g2_o21ai_1 _14589_ (.B1(_07293_),
    .Y(_07294_),
    .A1(\spiking_network_top_uut.all_data_out[796] ),
    .A2(net3842));
 sg13g2_mux2_1 _14590_ (.A0(net3841),
    .A1(net3900),
    .S(\spiking_network_top_uut.all_data_out[796] ),
    .X(_07295_));
 sg13g2_nand2_1 _14591_ (.Y(_07296_),
    .A(\spiking_network_top_uut.all_data_out[797] ),
    .B(_07295_));
 sg13g2_nand3_1 _14592_ (.B(_07294_),
    .C(_07296_),
    .A(\spiking_network_top_uut.all_data_out[798] ),
    .Y(_07297_));
 sg13g2_mux2_1 _14593_ (.A0(net3844),
    .A1(net3843),
    .S(\spiking_network_top_uut.all_data_out[796] ),
    .X(_07298_));
 sg13g2_nor2b_1 _14594_ (.A(\spiking_network_top_uut.all_data_out[796] ),
    .B_N(net3846),
    .Y(_07299_));
 sg13g2_a21oi_1 _14595_ (.A1(\spiking_network_top_uut.all_data_out[796] ),
    .A2(net3845),
    .Y(_07300_),
    .B1(_07299_));
 sg13g2_a21oi_1 _14596_ (.A1(\spiking_network_top_uut.all_data_out[797] ),
    .A2(_07298_),
    .Y(_07301_),
    .B1(\spiking_network_top_uut.all_data_out[798] ));
 sg13g2_o21ai_1 _14597_ (.B1(_07301_),
    .Y(_07302_),
    .A1(\spiking_network_top_uut.all_data_out[797] ),
    .A2(_07300_));
 sg13g2_nand3_1 _14598_ (.B(_07297_),
    .C(_07302_),
    .A(net4552),
    .Y(_07303_));
 sg13g2_o21ai_1 _14599_ (.B1(_07303_),
    .Y(_00698_),
    .A1(net4552),
    .A2(_03679_));
 sg13g2_nor2_1 _14600_ (.A(net4552),
    .B(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_dout ),
    .Y(_07304_));
 sg13g2_a21oi_1 _14601_ (.A1(net4552),
    .A2(_03679_),
    .Y(_00699_),
    .B1(_07304_));
 sg13g2_mux4_1 _14602_ (.S0(\spiking_network_top_uut.all_data_out[792] ),
    .A0(net3898),
    .A1(net3897),
    .A2(net3896),
    .A3(net3895),
    .S1(\spiking_network_top_uut.all_data_out[793] ),
    .X(_07305_));
 sg13g2_mux2_1 _14603_ (.A0(net3893),
    .A1(net3892),
    .S(\spiking_network_top_uut.all_data_out[792] ),
    .X(_07306_));
 sg13g2_nor2b_1 _14604_ (.A(\spiking_network_top_uut.all_data_out[792] ),
    .B_N(net3894),
    .Y(_07307_));
 sg13g2_a21oi_1 _14605_ (.A1(\spiking_network_top_uut.all_data_out[792] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[5] ),
    .Y(_07308_),
    .B1(_07307_));
 sg13g2_o21ai_1 _14606_ (.B1(\spiking_network_top_uut.all_data_out[794] ),
    .Y(_07309_),
    .A1(\spiking_network_top_uut.all_data_out[793] ),
    .A2(_07308_));
 sg13g2_a21oi_1 _14607_ (.A1(\spiking_network_top_uut.all_data_out[793] ),
    .A2(_07306_),
    .Y(_07310_),
    .B1(_07309_));
 sg13g2_o21ai_1 _14608_ (.B1(net4546),
    .Y(_07311_),
    .A1(\spiking_network_top_uut.all_data_out[794] ),
    .A2(_07305_));
 sg13g2_nand2_1 _14609_ (.Y(_07312_),
    .A(net3934),
    .B(net77));
 sg13g2_o21ai_1 _14610_ (.B1(_07312_),
    .Y(_00700_),
    .A1(_07310_),
    .A2(_07311_));
 sg13g2_mux2_1 _14611_ (.A0(net175),
    .A1(net77),
    .S(net4549),
    .X(_00701_));
 sg13g2_mux4_1 _14612_ (.S0(\spiking_network_top_uut.all_data_out[788] ),
    .A0(net3891),
    .A1(net3890),
    .A2(net3889),
    .A3(net3888),
    .S1(\spiking_network_top_uut.all_data_out[789] ),
    .X(_07313_));
 sg13g2_mux2_1 _14613_ (.A0(net3886),
    .A1(net3885),
    .S(\spiking_network_top_uut.all_data_out[788] ),
    .X(_07314_));
 sg13g2_nor2b_1 _14614_ (.A(\spiking_network_top_uut.all_data_out[788] ),
    .B_N(net3887),
    .Y(_07315_));
 sg13g2_a21oi_1 _14615_ (.A1(\spiking_network_top_uut.all_data_out[788] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[5] ),
    .Y(_07316_),
    .B1(_07315_));
 sg13g2_o21ai_1 _14616_ (.B1(\spiking_network_top_uut.all_data_out[790] ),
    .Y(_07317_),
    .A1(\spiking_network_top_uut.all_data_out[789] ),
    .A2(_07316_));
 sg13g2_a21oi_1 _14617_ (.A1(\spiking_network_top_uut.all_data_out[789] ),
    .A2(_07314_),
    .Y(_07318_),
    .B1(_07317_));
 sg13g2_o21ai_1 _14618_ (.B1(net4559),
    .Y(_07319_),
    .A1(\spiking_network_top_uut.all_data_out[790] ),
    .A2(_07313_));
 sg13g2_nand2_1 _14619_ (.Y(_07320_),
    .A(net3935),
    .B(net220));
 sg13g2_o21ai_1 _14620_ (.B1(_07320_),
    .Y(_00702_),
    .A1(_07318_),
    .A2(_07319_));
 sg13g2_mux2_1 _14621_ (.A0(net360),
    .A1(net220),
    .S(net4558),
    .X(_00703_));
 sg13g2_mux4_1 _14622_ (.S0(\spiking_network_top_uut.all_data_out[784] ),
    .A0(net3884),
    .A1(net3883),
    .A2(net3882),
    .A3(net3881),
    .S1(\spiking_network_top_uut.all_data_out[785] ),
    .X(_07321_));
 sg13g2_mux2_1 _14623_ (.A0(net3878),
    .A1(net3877),
    .S(\spiking_network_top_uut.all_data_out[784] ),
    .X(_07322_));
 sg13g2_nor2b_1 _14624_ (.A(\spiking_network_top_uut.all_data_out[784] ),
    .B_N(net3880),
    .Y(_07323_));
 sg13g2_a21oi_1 _14625_ (.A1(\spiking_network_top_uut.all_data_out[784] ),
    .A2(net3879),
    .Y(_07324_),
    .B1(_07323_));
 sg13g2_o21ai_1 _14626_ (.B1(\spiking_network_top_uut.all_data_out[786] ),
    .Y(_07325_),
    .A1(\spiking_network_top_uut.all_data_out[785] ),
    .A2(_07324_));
 sg13g2_a21oi_1 _14627_ (.A1(\spiking_network_top_uut.all_data_out[785] ),
    .A2(_07322_),
    .Y(_07326_),
    .B1(_07325_));
 sg13g2_o21ai_1 _14628_ (.B1(net4554),
    .Y(_07327_),
    .A1(\spiking_network_top_uut.all_data_out[786] ),
    .A2(_07321_));
 sg13g2_nand2_1 _14629_ (.Y(_07328_),
    .A(net3938),
    .B(net85));
 sg13g2_o21ai_1 _14630_ (.B1(_07328_),
    .Y(_00704_),
    .A1(_07326_),
    .A2(_07327_));
 sg13g2_mux2_1 _14631_ (.A0(net157),
    .A1(net85),
    .S(net4554),
    .X(_00705_));
 sg13g2_mux4_1 _14632_ (.S0(\spiking_network_top_uut.all_data_out[780] ),
    .A0(net3876),
    .A1(net3875),
    .A2(net3874),
    .A3(net3873),
    .S1(\spiking_network_top_uut.all_data_out[781] ),
    .X(_07329_));
 sg13g2_mux2_1 _14633_ (.A0(net3870),
    .A1(net3869),
    .S(\spiking_network_top_uut.all_data_out[780] ),
    .X(_07330_));
 sg13g2_nor2b_1 _14634_ (.A(\spiking_network_top_uut.all_data_out[780] ),
    .B_N(net3872),
    .Y(_07331_));
 sg13g2_a21oi_1 _14635_ (.A1(\spiking_network_top_uut.all_data_out[780] ),
    .A2(net3871),
    .Y(_07332_),
    .B1(_07331_));
 sg13g2_o21ai_1 _14636_ (.B1(\spiking_network_top_uut.all_data_out[782] ),
    .Y(_07333_),
    .A1(\spiking_network_top_uut.all_data_out[781] ),
    .A2(_07332_));
 sg13g2_a21oi_1 _14637_ (.A1(\spiking_network_top_uut.all_data_out[781] ),
    .A2(_07330_),
    .Y(_07334_),
    .B1(_07333_));
 sg13g2_o21ai_1 _14638_ (.B1(net4567),
    .Y(_07335_),
    .A1(\spiking_network_top_uut.all_data_out[782] ),
    .A2(_07329_));
 sg13g2_nand2_1 _14639_ (.Y(_07336_),
    .A(net3937),
    .B(net51));
 sg13g2_o21ai_1 _14640_ (.B1(_07336_),
    .Y(_00706_),
    .A1(_07334_),
    .A2(_07335_));
 sg13g2_mux2_1 _14641_ (.A0(net260),
    .A1(net51),
    .S(net4567),
    .X(_00707_));
 sg13g2_mux4_1 _14642_ (.S0(\spiking_network_top_uut.all_data_out[776] ),
    .A0(net3868),
    .A1(net3867),
    .A2(net3866),
    .A3(net3865),
    .S1(\spiking_network_top_uut.all_data_out[777] ),
    .X(_07337_));
 sg13g2_mux2_1 _14643_ (.A0(net3862),
    .A1(net3861),
    .S(\spiking_network_top_uut.all_data_out[776] ),
    .X(_07338_));
 sg13g2_nor2b_1 _14644_ (.A(\spiking_network_top_uut.all_data_out[776] ),
    .B_N(net3864),
    .Y(_07339_));
 sg13g2_a21oi_1 _14645_ (.A1(\spiking_network_top_uut.all_data_out[776] ),
    .A2(net3863),
    .Y(_07340_),
    .B1(_07339_));
 sg13g2_o21ai_1 _14646_ (.B1(\spiking_network_top_uut.all_data_out[778] ),
    .Y(_07341_),
    .A1(\spiking_network_top_uut.all_data_out[777] ),
    .A2(_07340_));
 sg13g2_a21oi_1 _14647_ (.A1(\spiking_network_top_uut.all_data_out[777] ),
    .A2(_07338_),
    .Y(_07342_),
    .B1(_07341_));
 sg13g2_o21ai_1 _14648_ (.B1(net4563),
    .Y(_07343_),
    .A1(\spiking_network_top_uut.all_data_out[778] ),
    .A2(_07337_));
 sg13g2_nand2_1 _14649_ (.Y(_07344_),
    .A(net3936),
    .B(net270));
 sg13g2_o21ai_1 _14650_ (.B1(_07344_),
    .Y(_00708_),
    .A1(_07342_),
    .A2(_07343_));
 sg13g2_mux2_1 _14651_ (.A0(net311),
    .A1(net270),
    .S(net4562),
    .X(_00709_));
 sg13g2_nand2_1 _14652_ (.Y(_07345_),
    .A(\spiking_network_top_uut.all_data_out[772] ),
    .B(_03664_));
 sg13g2_nor2_1 _14653_ (.A(\spiking_network_top_uut.all_data_out[772] ),
    .B(net3856),
    .Y(_07346_));
 sg13g2_nor2_1 _14654_ (.A(\spiking_network_top_uut.all_data_out[773] ),
    .B(_07346_),
    .Y(_07347_));
 sg13g2_mux2_1 _14655_ (.A0(net3855),
    .A1(net3854),
    .S(\spiking_network_top_uut.all_data_out[772] ),
    .X(_07348_));
 sg13g2_a221oi_1 _14656_ (.B2(\spiking_network_top_uut.all_data_out[773] ),
    .C1(_03513_),
    .B1(_07348_),
    .A1(_07345_),
    .Y(_07349_),
    .A2(_07347_));
 sg13g2_mux4_1 _14657_ (.S0(\spiking_network_top_uut.all_data_out[772] ),
    .A0(net3860),
    .A1(net3859),
    .A2(net3858),
    .A3(net3857),
    .S1(\spiking_network_top_uut.all_data_out[773] ),
    .X(_07350_));
 sg13g2_o21ai_1 _14658_ (.B1(net4536),
    .Y(_07351_),
    .A1(\spiking_network_top_uut.all_data_out[774] ),
    .A2(_07350_));
 sg13g2_nand2_1 _14659_ (.Y(_07352_),
    .A(net3932),
    .B(net71));
 sg13g2_o21ai_1 _14660_ (.B1(_07352_),
    .Y(_00710_),
    .A1(_07349_),
    .A2(_07351_));
 sg13g2_mux2_1 _14661_ (.A0(net305),
    .A1(net71),
    .S(net4536),
    .X(_00711_));
 sg13g2_mux2_1 _14662_ (.A0(net3851),
    .A1(net3850),
    .S(\spiking_network_top_uut.all_data_out[768] ),
    .X(_07353_));
 sg13g2_nor2b_1 _14663_ (.A(\spiking_network_top_uut.all_data_out[768] ),
    .B_N(net3853),
    .Y(_07354_));
 sg13g2_a21oi_1 _14664_ (.A1(\spiking_network_top_uut.all_data_out[768] ),
    .A2(net3852),
    .Y(_07355_),
    .B1(_07354_));
 sg13g2_a21oi_1 _14665_ (.A1(\spiking_network_top_uut.all_data_out[769] ),
    .A2(_07353_),
    .Y(_07356_),
    .B1(\spiking_network_top_uut.all_data_out[770] ));
 sg13g2_o21ai_1 _14666_ (.B1(_07356_),
    .Y(_07357_),
    .A1(\spiking_network_top_uut.all_data_out[769] ),
    .A2(_07355_));
 sg13g2_mux2_1 _14667_ (.A0(net3848),
    .A1(net3847),
    .S(\spiking_network_top_uut.all_data_out[768] ),
    .X(_07358_));
 sg13g2_nand2_1 _14668_ (.Y(_07359_),
    .A(\spiking_network_top_uut.all_data_out[769] ),
    .B(_07358_));
 sg13g2_a21oi_1 _14669_ (.A1(\spiking_network_top_uut.all_data_out[768] ),
    .A2(_03663_),
    .Y(_07360_),
    .B1(\spiking_network_top_uut.all_data_out[769] ));
 sg13g2_o21ai_1 _14670_ (.B1(_07360_),
    .Y(_07361_),
    .A1(\spiking_network_top_uut.all_data_out[768] ),
    .A2(net3849));
 sg13g2_nand3_1 _14671_ (.B(_07359_),
    .C(_07361_),
    .A(\spiking_network_top_uut.all_data_out[770] ),
    .Y(_07362_));
 sg13g2_nand3_1 _14672_ (.B(_07357_),
    .C(_07362_),
    .A(net4539),
    .Y(_07363_));
 sg13g2_o21ai_1 _14673_ (.B1(_07363_),
    .Y(_00712_),
    .A1(net4534),
    .A2(_03680_));
 sg13g2_nor3_2 _14674_ (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[2] ),
    .B(net339),
    .C(net320),
    .Y(_07364_));
 sg13g2_nor2b_2 _14675_ (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[3] ),
    .B_N(_07364_),
    .Y(_07365_));
 sg13g2_nor2b_1 _14676_ (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[4] ),
    .B_N(_07365_),
    .Y(_07366_));
 sg13g2_nand2b_2 _14677_ (.Y(_07367_),
    .B(_07365_),
    .A_N(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[4] ));
 sg13g2_o21ai_1 _14678_ (.B1(net4529),
    .Y(_07368_),
    .A1(net3627),
    .A2(_07367_));
 sg13g2_nor2b_1 _14679_ (.A(net3626),
    .B_N(_00084_),
    .Y(_07369_));
 sg13g2_a21oi_1 _14680_ (.A1(net4283),
    .A2(net3626),
    .Y(_07370_),
    .B1(_07369_));
 sg13g2_nand2_1 _14681_ (.Y(_07371_),
    .A(net320),
    .B(_07368_));
 sg13g2_o21ai_1 _14682_ (.B1(_07371_),
    .Y(_00713_),
    .A1(_07368_),
    .A2(_07370_));
 sg13g2_xor2_1 _14683_ (.B(net320),
    .A(net339),
    .X(_07372_));
 sg13g2_nor2_1 _14684_ (.A(net3626),
    .B(_07372_),
    .Y(_07373_));
 sg13g2_a21oi_1 _14685_ (.A1(net4280),
    .A2(net3626),
    .Y(_07374_),
    .B1(_07373_));
 sg13g2_nand2_1 _14686_ (.Y(_07375_),
    .A(net339),
    .B(_07368_));
 sg13g2_o21ai_1 _14687_ (.B1(_07375_),
    .Y(_00714_),
    .A1(_07368_),
    .A2(_07374_));
 sg13g2_o21ai_1 _14688_ (.B1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[2] ),
    .Y(_07376_),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[1] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[0] ));
 sg13g2_nor2b_1 _14689_ (.A(_07364_),
    .B_N(_07376_),
    .Y(_07377_));
 sg13g2_nor2_1 _14690_ (.A(net3626),
    .B(_07377_),
    .Y(_07378_));
 sg13g2_a21oi_1 _14691_ (.A1(net4276),
    .A2(net3626),
    .Y(_07379_),
    .B1(_07378_));
 sg13g2_nand2_1 _14692_ (.Y(_07380_),
    .A(net213),
    .B(_07368_));
 sg13g2_o21ai_1 _14693_ (.B1(_07380_),
    .Y(_00715_),
    .A1(_07368_),
    .A2(_07379_));
 sg13g2_nand2_1 _14694_ (.Y(_07381_),
    .A(net4273),
    .B(net3626));
 sg13g2_xnor2_1 _14695_ (.Y(_07382_),
    .A(net443),
    .B(_07364_));
 sg13g2_o21ai_1 _14696_ (.B1(_07381_),
    .Y(_07383_),
    .A1(net3626),
    .A2(_07382_));
 sg13g2_mux2_1 _14697_ (.A0(_07383_),
    .A1(net443),
    .S(_07368_),
    .X(_00716_));
 sg13g2_nand2_1 _14698_ (.Y(_07384_),
    .A(net3921),
    .B(net218));
 sg13g2_nand2b_1 _14699_ (.Y(_07385_),
    .B(net218),
    .A_N(_07365_));
 sg13g2_a21oi_1 _14700_ (.A1(_07367_),
    .A2(_07385_),
    .Y(_07386_),
    .B1(net3627));
 sg13g2_a21oi_1 _14701_ (.A1(net4269),
    .A2(net3627),
    .Y(_07387_),
    .B1(_07386_));
 sg13g2_o21ai_1 _14702_ (.B1(_07384_),
    .Y(_00717_),
    .A1(_07368_),
    .A2(_07387_));
 sg13g2_mux2_1 _14703_ (.A0(net234),
    .A1(net76),
    .S(net4534),
    .X(_00718_));
 sg13g2_nor2_1 _14704_ (.A(_00079_),
    .B(net3741),
    .Y(_07388_));
 sg13g2_nor2_2 _14705_ (.A(net3746),
    .B(_07388_),
    .Y(_07389_));
 sg13g2_nor2_1 _14706_ (.A(_00079_),
    .B(_07389_),
    .Y(_07390_));
 sg13g2_nand2b_1 _14707_ (.Y(_07391_),
    .B(_07389_),
    .A_N(_00079_));
 sg13g2_o21ai_1 _14708_ (.B1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ),
    .Y(_07392_),
    .A1(_00079_),
    .A2(_07389_));
 sg13g2_inv_1 _14709_ (.Y(_07393_),
    .A(_07392_));
 sg13g2_nor2_1 _14710_ (.A(_00080_),
    .B(net3905),
    .Y(_07394_));
 sg13g2_a221oi_1 _14711_ (.B2(_07388_),
    .C1(_07394_),
    .B1(net3905),
    .A1(_03487_),
    .Y(_07395_),
    .A2(net3746));
 sg13g2_nand2_1 _14712_ (.Y(_07396_),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ),
    .B(_07395_));
 sg13g2_o21ai_1 _14713_ (.B1(net3917),
    .Y(_07397_),
    .A1(_00079_),
    .A2(net3912));
 sg13g2_a221oi_1 _14714_ (.B2(_03486_),
    .C1(_07397_),
    .B1(net3901),
    .A1(_03487_),
    .Y(_07398_),
    .A2(net3738));
 sg13g2_and2_1 _14715_ (.A(_00083_),
    .B(net3746),
    .X(_07399_));
 sg13g2_nor3_2 _14716_ (.A(_03488_),
    .B(_07398_),
    .C(_07399_),
    .Y(_07400_));
 sg13g2_xnor2_1 _14717_ (.Y(_07401_),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ),
    .B(_07395_));
 sg13g2_o21ai_1 _14718_ (.B1(_07396_),
    .Y(_07402_),
    .A1(_07400_),
    .A2(_07401_));
 sg13g2_inv_1 _14719_ (.Y(_07403_),
    .A(_07402_));
 sg13g2_a21o_1 _14720_ (.A2(net3746),
    .A1(_00080_),
    .B1(_07389_),
    .X(_07404_));
 sg13g2_xnor2_1 _14721_ (.Y(_07405_),
    .A(_03487_),
    .B(_07404_));
 sg13g2_nand2_1 _14722_ (.Y(_07406_),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ),
    .B(_07404_));
 sg13g2_o21ai_1 _14723_ (.B1(_07406_),
    .Y(_07407_),
    .A1(_07403_),
    .A2(_07405_));
 sg13g2_xnor2_1 _14724_ (.Y(_07408_),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ),
    .B(_07390_));
 sg13g2_a21oi_1 _14725_ (.A1(_07407_),
    .A2(_07408_),
    .Y(_07409_),
    .B1(_07393_));
 sg13g2_a22oi_1 _14726_ (.Y(_07410_),
    .B1(_07391_),
    .B2(_07409_),
    .A2(_07389_),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ));
 sg13g2_a21oi_2 _14727_ (.B1(_07410_),
    .Y(_07411_),
    .A2(_00079_),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ));
 sg13g2_nor2_1 _14728_ (.A(net3704),
    .B(_07411_),
    .Y(_07412_));
 sg13g2_mux2_1 _14729_ (.A0(net4599),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[771] ),
    .X(_07413_));
 sg13g2_nand2_1 _14730_ (.Y(_07414_),
    .A(\spiking_network_top_uut.all_data_out[257] ),
    .B(_07413_));
 sg13g2_mux2_1 _14731_ (.A0(net4598),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[775] ),
    .X(_07415_));
 sg13g2_nand2_1 _14732_ (.Y(_07416_),
    .A(\spiking_network_top_uut.all_data_out[259] ),
    .B(_07415_));
 sg13g2_nor2_1 _14733_ (.A(_07414_),
    .B(_07416_),
    .Y(_07417_));
 sg13g2_nand4_1 _14734_ (.B(\spiking_network_top_uut.all_data_out[258] ),
    .C(_07413_),
    .A(\spiking_network_top_uut.all_data_out[256] ),
    .Y(_07418_),
    .D(_07415_));
 sg13g2_inv_1 _14735_ (.Y(_07419_),
    .A(_07418_));
 sg13g2_xor2_1 _14736_ (.B(_07416_),
    .A(_07414_),
    .X(_07420_));
 sg13g2_a21oi_2 _14737_ (.B1(_07417_),
    .Y(_07421_),
    .A2(_07420_),
    .A1(_07418_));
 sg13g2_mux2_2 _14738_ (.A0(net4597),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[779] ),
    .X(_07422_));
 sg13g2_nand2_1 _14739_ (.Y(_07423_),
    .A(\spiking_network_top_uut.all_data_out[261] ),
    .B(_07422_));
 sg13g2_mux2_2 _14740_ (.A0(net4596),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[783] ),
    .X(_07424_));
 sg13g2_nand2_1 _14741_ (.Y(_07425_),
    .A(\spiking_network_top_uut.all_data_out[263] ),
    .B(_07424_));
 sg13g2_nor2_1 _14742_ (.A(_07423_),
    .B(_07425_),
    .Y(_07426_));
 sg13g2_nand2_1 _14743_ (.Y(_07427_),
    .A(\spiking_network_top_uut.all_data_out[260] ),
    .B(_07422_));
 sg13g2_nand2_1 _14744_ (.Y(_07428_),
    .A(\spiking_network_top_uut.all_data_out[262] ),
    .B(_07424_));
 sg13g2_or2_2 _14745_ (.X(_07429_),
    .B(_07428_),
    .A(_07427_));
 sg13g2_xor2_1 _14746_ (.B(_07425_),
    .A(_07423_),
    .X(_07430_));
 sg13g2_a21oi_2 _14747_ (.B1(_07426_),
    .Y(_07431_),
    .A2(_07430_),
    .A1(_07429_));
 sg13g2_mux2_2 _14748_ (.A0(net4595),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[787] ),
    .X(_07432_));
 sg13g2_mux2_2 _14749_ (.A0(net4594),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[791] ),
    .X(_07433_));
 sg13g2_a22oi_1 _14750_ (.Y(_07434_),
    .B1(_07433_),
    .B2(\spiking_network_top_uut.all_data_out[267] ),
    .A2(_07432_),
    .A1(\spiking_network_top_uut.all_data_out[265] ));
 sg13g2_and4_2 _14751_ (.A(\spiking_network_top_uut.all_data_out[264] ),
    .B(\spiking_network_top_uut.all_data_out[266] ),
    .C(_07432_),
    .D(_07433_),
    .X(_07435_));
 sg13g2_nand4_1 _14752_ (.B(\spiking_network_top_uut.all_data_out[266] ),
    .C(_07432_),
    .A(\spiking_network_top_uut.all_data_out[264] ),
    .Y(_07436_),
    .D(_07433_));
 sg13g2_and4_1 _14753_ (.A(\spiking_network_top_uut.all_data_out[265] ),
    .B(\spiking_network_top_uut.all_data_out[267] ),
    .C(_07432_),
    .D(_07433_),
    .X(_07437_));
 sg13g2_nand4_1 _14754_ (.B(\spiking_network_top_uut.all_data_out[267] ),
    .C(_07432_),
    .A(\spiking_network_top_uut.all_data_out[265] ),
    .Y(_07438_),
    .D(_07433_));
 sg13g2_nand3b_1 _14755_ (.B(_07435_),
    .C(_07438_),
    .Y(_07439_),
    .A_N(_07434_));
 sg13g2_a21oi_2 _14756_ (.B1(_07434_),
    .Y(_07440_),
    .A2(_07438_),
    .A1(_07435_));
 sg13g2_mux2_2 _14757_ (.A0(net4593),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[795] ),
    .X(_07441_));
 sg13g2_mux2_2 _14758_ (.A0(net4592),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[799] ),
    .X(_07442_));
 sg13g2_and4_1 _14759_ (.A(\spiking_network_top_uut.all_data_out[269] ),
    .B(\spiking_network_top_uut.all_data_out[271] ),
    .C(_07441_),
    .D(_07442_),
    .X(_07443_));
 sg13g2_nand4_1 _14760_ (.B(\spiking_network_top_uut.all_data_out[271] ),
    .C(_07441_),
    .A(\spiking_network_top_uut.all_data_out[269] ),
    .Y(_07444_),
    .D(_07442_));
 sg13g2_and4_1 _14761_ (.A(\spiking_network_top_uut.all_data_out[268] ),
    .B(\spiking_network_top_uut.all_data_out[270] ),
    .C(_07441_),
    .D(_07442_),
    .X(_07445_));
 sg13g2_a22oi_1 _14762_ (.Y(_07446_),
    .B1(_07442_),
    .B2(\spiking_network_top_uut.all_data_out[271] ),
    .A2(_07441_),
    .A1(\spiking_network_top_uut.all_data_out[269] ));
 sg13g2_or3_2 _14763_ (.A(_07443_),
    .B(_07445_),
    .C(_07446_),
    .X(_07447_));
 sg13g2_o21ai_1 _14764_ (.B1(_07444_),
    .Y(_07448_),
    .A1(_07445_),
    .A2(_07446_));
 sg13g2_nand3b_1 _14765_ (.B(_07440_),
    .C(_07448_),
    .Y(_07449_),
    .A_N(_07431_));
 sg13g2_inv_1 _14766_ (.Y(_07450_),
    .A(_07449_));
 sg13g2_or2_1 _14767_ (.X(_07451_),
    .B(_07449_),
    .A(_07421_));
 sg13g2_nor2_1 _14768_ (.A(_07440_),
    .B(_07448_),
    .Y(_07452_));
 sg13g2_and2_1 _14769_ (.A(_07431_),
    .B(_07452_),
    .X(_07453_));
 sg13g2_nand2_1 _14770_ (.Y(_07454_),
    .A(_07421_),
    .B(_07453_));
 sg13g2_and2_1 _14771_ (.A(_07451_),
    .B(_07454_),
    .X(_07455_));
 sg13g2_xnor2_1 _14772_ (.Y(_07456_),
    .A(_07391_),
    .B(_07409_));
 sg13g2_nand2_1 _14773_ (.Y(_07457_),
    .A(_07455_),
    .B(_07456_));
 sg13g2_nand2_1 _14774_ (.Y(_07458_),
    .A(_07451_),
    .B(_07457_));
 sg13g2_xor2_1 _14775_ (.B(_07455_),
    .A(_07411_),
    .X(_07459_));
 sg13g2_nand2_1 _14776_ (.Y(_07460_),
    .A(_07458_),
    .B(_07459_));
 sg13g2_xnor2_1 _14777_ (.Y(_07461_),
    .A(_07455_),
    .B(_07456_));
 sg13g2_o21ai_1 _14778_ (.B1(_07445_),
    .Y(_07462_),
    .A1(_07443_),
    .A2(_07446_));
 sg13g2_o21ai_1 _14779_ (.B1(_07436_),
    .Y(_07463_),
    .A1(_07434_),
    .A2(_07437_));
 sg13g2_o21ai_1 _14780_ (.B1(_07435_),
    .Y(_07464_),
    .A1(_07434_),
    .A2(_07437_));
 sg13g2_nand3b_1 _14781_ (.B(_07436_),
    .C(_07438_),
    .Y(_07465_),
    .A_N(_07434_));
 sg13g2_a22oi_1 _14782_ (.Y(_07466_),
    .B1(_07464_),
    .B2(_07465_),
    .A2(_07462_),
    .A1(_07447_));
 sg13g2_xor2_1 _14783_ (.B(_07430_),
    .A(_07429_),
    .X(_07467_));
 sg13g2_xnor2_1 _14784_ (.Y(_07468_),
    .A(_07429_),
    .B(_07430_));
 sg13g2_and4_1 _14785_ (.A(_07447_),
    .B(_07462_),
    .C(_07464_),
    .D(_07465_),
    .X(_07469_));
 sg13g2_nand4_1 _14786_ (.B(_07462_),
    .C(_07464_),
    .A(_07447_),
    .Y(_07470_),
    .D(_07465_));
 sg13g2_and4_1 _14787_ (.A(_07439_),
    .B(_07447_),
    .C(_07462_),
    .D(_07463_),
    .X(_07471_));
 sg13g2_a22oi_1 _14788_ (.Y(_07472_),
    .B1(_07463_),
    .B2(_07439_),
    .A2(_07462_),
    .A1(_07447_));
 sg13g2_nor3_2 _14789_ (.A(_07466_),
    .B(_07467_),
    .C(_07469_),
    .Y(_07473_));
 sg13g2_a21oi_2 _14790_ (.B1(_07466_),
    .Y(_07474_),
    .A2(_07470_),
    .A1(_07468_));
 sg13g2_xor2_1 _14791_ (.B(_07448_),
    .A(_07440_),
    .X(_07475_));
 sg13g2_xnor2_1 _14792_ (.Y(_07476_),
    .A(_07431_),
    .B(_07475_));
 sg13g2_nand2b_1 _14793_ (.Y(_07477_),
    .B(_07476_),
    .A_N(_07474_));
 sg13g2_xnor2_1 _14794_ (.Y(_07478_),
    .A(_07474_),
    .B(_07476_));
 sg13g2_nand2b_1 _14795_ (.Y(_07479_),
    .B(_07478_),
    .A_N(_07421_));
 sg13g2_nand2_1 _14796_ (.Y(_07480_),
    .A(_07477_),
    .B(_07479_));
 sg13g2_nor2_1 _14797_ (.A(_07450_),
    .B(_07453_),
    .Y(_07481_));
 sg13g2_xnor2_1 _14798_ (.Y(_07482_),
    .A(_07421_),
    .B(_07481_));
 sg13g2_and2_1 _14799_ (.A(_07480_),
    .B(_07482_),
    .X(_07483_));
 sg13g2_xor2_1 _14800_ (.B(_07482_),
    .A(_07480_),
    .X(_07484_));
 sg13g2_xnor2_1 _14801_ (.Y(_07485_),
    .A(_07407_),
    .B(_07408_));
 sg13g2_inv_1 _14802_ (.Y(_07486_),
    .A(_07485_));
 sg13g2_a21oi_1 _14803_ (.A1(_07484_),
    .A2(_07486_),
    .Y(_07487_),
    .B1(_07483_));
 sg13g2_nor2_1 _14804_ (.A(_07461_),
    .B(_07487_),
    .Y(_07488_));
 sg13g2_xnor2_1 _14805_ (.Y(_07489_),
    .A(_07484_),
    .B(_07485_));
 sg13g2_a22oi_1 _14806_ (.Y(_07490_),
    .B1(_07442_),
    .B2(\spiking_network_top_uut.all_data_out[270] ),
    .A2(_07441_),
    .A1(\spiking_network_top_uut.all_data_out[268] ));
 sg13g2_nor2_1 _14807_ (.A(_07445_),
    .B(_07490_),
    .Y(_07491_));
 sg13g2_a22oi_1 _14808_ (.Y(_07492_),
    .B1(_07433_),
    .B2(\spiking_network_top_uut.all_data_out[266] ),
    .A2(_07432_),
    .A1(\spiking_network_top_uut.all_data_out[264] ));
 sg13g2_nor2_1 _14809_ (.A(_07435_),
    .B(_07492_),
    .Y(_07493_));
 sg13g2_and2_1 _14810_ (.A(_07491_),
    .B(_07493_),
    .X(_07494_));
 sg13g2_xor2_1 _14811_ (.B(_07428_),
    .A(_07427_),
    .X(_07495_));
 sg13g2_xor2_1 _14812_ (.B(_07493_),
    .A(_07491_),
    .X(_07496_));
 sg13g2_a21oi_2 _14813_ (.B1(_07494_),
    .Y(_07497_),
    .A2(_07496_),
    .A1(_07495_));
 sg13g2_nor3_2 _14814_ (.A(_07468_),
    .B(_07471_),
    .C(_07472_),
    .Y(_07498_));
 sg13g2_nor3_1 _14815_ (.A(_07473_),
    .B(_07497_),
    .C(_07498_),
    .Y(_07499_));
 sg13g2_or3_1 _14816_ (.A(_07473_),
    .B(_07497_),
    .C(_07498_),
    .X(_07500_));
 sg13g2_xnor2_1 _14817_ (.Y(_07501_),
    .A(_07418_),
    .B(_07420_));
 sg13g2_o21ai_1 _14818_ (.B1(_07497_),
    .Y(_07502_),
    .A1(_07473_),
    .A2(_07498_));
 sg13g2_nand3_1 _14819_ (.B(_07501_),
    .C(_07502_),
    .A(_07500_),
    .Y(_07503_));
 sg13g2_a21o_2 _14820_ (.A2(_07502_),
    .A1(_07501_),
    .B1(_07499_),
    .X(_07504_));
 sg13g2_xnor2_1 _14821_ (.Y(_07505_),
    .A(_07421_),
    .B(_07478_));
 sg13g2_nand2_1 _14822_ (.Y(_07506_),
    .A(_07504_),
    .B(_07505_));
 sg13g2_xnor2_1 _14823_ (.Y(_07507_),
    .A(_07402_),
    .B(_07405_));
 sg13g2_inv_1 _14824_ (.Y(_07508_),
    .A(_07507_));
 sg13g2_xnor2_1 _14825_ (.Y(_07509_),
    .A(_07504_),
    .B(_07505_));
 sg13g2_o21ai_1 _14826_ (.B1(_07506_),
    .Y(_07510_),
    .A1(_07508_),
    .A2(_07509_));
 sg13g2_nand2_1 _14827_ (.Y(_07511_),
    .A(_07489_),
    .B(_07510_));
 sg13g2_a22oi_1 _14828_ (.Y(_07512_),
    .B1(_07415_),
    .B2(\spiking_network_top_uut.all_data_out[258] ),
    .A2(_07413_),
    .A1(\spiking_network_top_uut.all_data_out[256] ));
 sg13g2_xnor2_1 _14829_ (.Y(_07513_),
    .A(_07495_),
    .B(_07496_));
 sg13g2_nor3_2 _14830_ (.A(_07419_),
    .B(_07512_),
    .C(_07513_),
    .Y(_07514_));
 sg13g2_a21o_2 _14831_ (.A2(_07502_),
    .A1(_07500_),
    .B1(_07501_),
    .X(_07515_));
 sg13g2_nand3_1 _14832_ (.B(_07514_),
    .C(_07515_),
    .A(_07503_),
    .Y(_07516_));
 sg13g2_a21oi_1 _14833_ (.A1(_07503_),
    .A2(_07515_),
    .Y(_07517_),
    .B1(_07514_));
 sg13g2_a21o_1 _14834_ (.A2(_07515_),
    .A1(_07503_),
    .B1(_07514_),
    .X(_07518_));
 sg13g2_xnor2_1 _14835_ (.Y(_07519_),
    .A(_07400_),
    .B(_07401_));
 sg13g2_inv_1 _14836_ (.Y(_07520_),
    .A(_07519_));
 sg13g2_and3_1 _14837_ (.X(_07521_),
    .A(_07516_),
    .B(_07518_),
    .C(_07520_));
 sg13g2_o21ai_1 _14838_ (.B1(_07516_),
    .Y(_07522_),
    .A1(_07517_),
    .A2(_07519_));
 sg13g2_xnor2_1 _14839_ (.Y(_07523_),
    .A(_07508_),
    .B(_07509_));
 sg13g2_nor2b_1 _14840_ (.A(_07523_),
    .B_N(_07522_),
    .Y(_07524_));
 sg13g2_a21oi_1 _14841_ (.A1(_07516_),
    .A2(_07518_),
    .Y(_07525_),
    .B1(_07520_));
 sg13g2_o21ai_1 _14842_ (.B1(_07513_),
    .Y(_07526_),
    .A1(_07419_),
    .A2(_07512_));
 sg13g2_nand2b_1 _14843_ (.Y(_07527_),
    .B(_07526_),
    .A_N(_07514_));
 sg13g2_o21ai_1 _14844_ (.B1(_03488_),
    .Y(_07528_),
    .A1(_07398_),
    .A2(_07399_));
 sg13g2_nor2b_1 _14845_ (.A(_07400_),
    .B_N(_07528_),
    .Y(_07529_));
 sg13g2_or2_1 _14846_ (.X(_07530_),
    .B(_07529_),
    .A(_07527_));
 sg13g2_nor3_2 _14847_ (.A(_07521_),
    .B(_07525_),
    .C(_07530_),
    .Y(_07531_));
 sg13g2_nand2b_1 _14848_ (.Y(_07532_),
    .B(_07523_),
    .A_N(_07522_));
 sg13g2_nand2b_1 _14849_ (.Y(_07533_),
    .B(_07532_),
    .A_N(_07524_));
 sg13g2_a21oi_1 _14850_ (.A1(_07531_),
    .A2(_07532_),
    .Y(_07534_),
    .B1(_07524_));
 sg13g2_nor2_1 _14851_ (.A(_07489_),
    .B(_07510_),
    .Y(_07535_));
 sg13g2_xor2_1 _14852_ (.B(_07510_),
    .A(_07489_),
    .X(_07536_));
 sg13g2_nand2b_1 _14853_ (.Y(_07537_),
    .B(_07536_),
    .A_N(_07534_));
 sg13g2_o21ai_1 _14854_ (.B1(_07511_),
    .Y(_07538_),
    .A1(_07534_),
    .A2(_07535_));
 sg13g2_xor2_1 _14855_ (.B(_07487_),
    .A(_07461_),
    .X(_07539_));
 sg13g2_and2_1 _14856_ (.A(_07538_),
    .B(_07539_),
    .X(_07540_));
 sg13g2_a21oi_1 _14857_ (.A1(_07538_),
    .A2(_07539_),
    .Y(_07541_),
    .B1(_07488_));
 sg13g2_xnor2_1 _14858_ (.Y(_07542_),
    .A(_07458_),
    .B(_07459_));
 sg13g2_o21ai_1 _14859_ (.B1(_07460_),
    .Y(_07543_),
    .A1(_07541_),
    .A2(_07542_));
 sg13g2_mux2_1 _14860_ (.A0(_07454_),
    .A1(_07451_),
    .S(_07411_),
    .X(_07544_));
 sg13g2_xnor2_1 _14861_ (.Y(_07545_),
    .A(_07543_),
    .B(_07544_));
 sg13g2_a21oi_2 _14862_ (.B1(_07412_),
    .Y(_07546_),
    .A2(_07545_),
    .A1(_07366_));
 sg13g2_xnor2_1 _14863_ (.Y(_07547_),
    .A(_07541_),
    .B(_07542_));
 sg13g2_a21oi_1 _14864_ (.A1(net3704),
    .A2(_07547_),
    .Y(_07548_),
    .B1(_07412_));
 sg13g2_nor2_1 _14865_ (.A(_07538_),
    .B(_07539_),
    .Y(_07549_));
 sg13g2_nor3_1 _14866_ (.A(_07367_),
    .B(_07540_),
    .C(_07549_),
    .Y(_07550_));
 sg13g2_a21o_1 _14867_ (.A2(_07456_),
    .A1(_07367_),
    .B1(_07550_),
    .X(_07551_));
 sg13g2_nand2_1 _14868_ (.Y(_07552_),
    .A(_07548_),
    .B(_07551_));
 sg13g2_a21oi_2 _14869_ (.B1(net3628),
    .Y(_07553_),
    .A2(_07552_),
    .A1(_07546_));
 sg13g2_nand2_1 _14870_ (.Y(_07554_),
    .A(net4530),
    .B(_07553_));
 sg13g2_nor2_1 _14871_ (.A(_07548_),
    .B(_07551_),
    .Y(_07555_));
 sg13g2_nor2_2 _14872_ (.A(_07546_),
    .B(_07555_),
    .Y(_07556_));
 sg13g2_nor2_1 _14873_ (.A(_07367_),
    .B(_07527_),
    .Y(_07557_));
 sg13g2_xnor2_1 _14874_ (.Y(_07558_),
    .A(_07529_),
    .B(_07557_));
 sg13g2_nor2_1 _14875_ (.A(_07556_),
    .B(_07558_),
    .Y(_07559_));
 sg13g2_xor2_1 _14876_ (.B(net486),
    .A(net4312),
    .X(_07560_));
 sg13g2_a22oi_1 _14877_ (.Y(_07561_),
    .B1(_00015_),
    .B2(_07560_),
    .A2(net486),
    .A1(net3920));
 sg13g2_o21ai_1 _14878_ (.B1(_07561_),
    .Y(_00719_),
    .A1(_07554_),
    .A2(_07559_));
 sg13g2_o21ai_1 _14879_ (.B1(_07530_),
    .Y(_07562_),
    .A1(_07521_),
    .A2(_07525_));
 sg13g2_nand3b_1 _14880_ (.B(_07562_),
    .C(net3704),
    .Y(_07563_),
    .A_N(_07531_));
 sg13g2_o21ai_1 _14881_ (.B1(_07563_),
    .Y(_07564_),
    .A1(net3704),
    .A2(_07519_));
 sg13g2_o21ai_1 _14882_ (.B1(_07553_),
    .Y(_07565_),
    .A1(_07556_),
    .A2(_07564_));
 sg13g2_xor2_1 _14883_ (.B(_04835_),
    .A(_04834_),
    .X(_07566_));
 sg13g2_a21oi_1 _14884_ (.A1(net3628),
    .A2(_07566_),
    .Y(_07567_),
    .B1(net3921));
 sg13g2_a22oi_1 _14885_ (.Y(_00720_),
    .B1(_07565_),
    .B2(_07567_),
    .A2(_03423_),
    .A1(net3921));
 sg13g2_xnor2_1 _14886_ (.Y(_07568_),
    .A(_07531_),
    .B(_07533_));
 sg13g2_nand2_1 _14887_ (.Y(_07569_),
    .A(net3704),
    .B(_07568_));
 sg13g2_o21ai_1 _14888_ (.B1(_07569_),
    .Y(_07570_),
    .A1(net3704),
    .A2(_07508_));
 sg13g2_nor2_1 _14889_ (.A(_07556_),
    .B(_07570_),
    .Y(_07571_));
 sg13g2_xnor2_1 _14890_ (.Y(_07572_),
    .A(_04832_),
    .B(_04836_));
 sg13g2_a22oi_1 _14891_ (.Y(_07573_),
    .B1(_00015_),
    .B2(_07572_),
    .A2(net537),
    .A1(net3920));
 sg13g2_o21ai_1 _14892_ (.B1(_07573_),
    .Y(_00721_),
    .A1(_07554_),
    .A2(_07571_));
 sg13g2_nor2b_1 _14893_ (.A(_07536_),
    .B_N(_07534_),
    .Y(_07574_));
 sg13g2_nand3b_1 _14894_ (.B(net3704),
    .C(_07537_),
    .Y(_07575_),
    .A_N(_07574_));
 sg13g2_o21ai_1 _14895_ (.B1(_07575_),
    .Y(_07576_),
    .A1(net3704),
    .A2(_07485_));
 sg13g2_o21ai_1 _14896_ (.B1(_07553_),
    .Y(_07577_),
    .A1(_07556_),
    .A2(_07576_));
 sg13g2_or3_1 _14897_ (.A(_04830_),
    .B(_04831_),
    .C(_04837_),
    .X(_07578_));
 sg13g2_and2_1 _14898_ (.A(_04838_),
    .B(_07578_),
    .X(_07579_));
 sg13g2_a21oi_1 _14899_ (.A1(net3628),
    .A2(_07579_),
    .Y(_07580_),
    .B1(net3921));
 sg13g2_a22oi_1 _14900_ (.Y(_00722_),
    .B1(_07577_),
    .B2(_07580_),
    .A2(_03422_),
    .A1(net3921));
 sg13g2_nand2b_1 _14901_ (.Y(_07581_),
    .B(_07546_),
    .A_N(net3628));
 sg13g2_a21oi_1 _14902_ (.A1(_04829_),
    .A2(_04839_),
    .Y(_07582_),
    .B1(net3921));
 sg13g2_a22oi_1 _14903_ (.Y(_00723_),
    .B1(_07581_),
    .B2(_07582_),
    .A2(_03421_),
    .A1(net3921));
 sg13g2_mux4_1 _14904_ (.S0(\spiking_network_top_uut.all_data_out[828] ),
    .A0(net3846),
    .A1(net3845),
    .A2(net3844),
    .A3(net3843),
    .S1(\spiking_network_top_uut.all_data_out[829] ),
    .X(_07583_));
 sg13g2_mux2_1 _14905_ (.A0(net3841),
    .A1(net3900),
    .S(\spiking_network_top_uut.all_data_out[828] ),
    .X(_07584_));
 sg13g2_nor2b_1 _14906_ (.A(\spiking_network_top_uut.all_data_out[828] ),
    .B_N(net3842),
    .Y(_07585_));
 sg13g2_a21oi_1 _14907_ (.A1(\spiking_network_top_uut.all_data_out[828] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[5] ),
    .Y(_07586_),
    .B1(_07585_));
 sg13g2_o21ai_1 _14908_ (.B1(\spiking_network_top_uut.all_data_out[830] ),
    .Y(_07587_),
    .A1(\spiking_network_top_uut.all_data_out[829] ),
    .A2(_07586_));
 sg13g2_a21oi_1 _14909_ (.A1(\spiking_network_top_uut.all_data_out[829] ),
    .A2(_07584_),
    .Y(_07588_),
    .B1(_07587_));
 sg13g2_o21ai_1 _14910_ (.B1(net4549),
    .Y(_07589_),
    .A1(\spiking_network_top_uut.all_data_out[830] ),
    .A2(_07583_));
 sg13g2_nand2_1 _14911_ (.Y(_07590_),
    .A(net3933),
    .B(net105));
 sg13g2_o21ai_1 _14912_ (.B1(_07590_),
    .Y(_00724_),
    .A1(_07588_),
    .A2(_07589_));
 sg13g2_mux2_1 _14913_ (.A0(net3898),
    .A1(net4593),
    .S(net4547),
    .X(_00725_));
 sg13g2_mux2_1 _14914_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[1] ),
    .A1(net3898),
    .S(net4545),
    .X(_00726_));
 sg13g2_mux2_1 _14915_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[2] ),
    .A1(net3897),
    .S(net4546),
    .X(_00727_));
 sg13g2_mux2_1 _14916_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[3] ),
    .A1(net3896),
    .S(net4546),
    .X(_00728_));
 sg13g2_mux2_1 _14917_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[4] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[3] ),
    .S(net4546),
    .X(_00729_));
 sg13g2_nand2_1 _14918_ (.Y(_07591_),
    .A(net4545),
    .B(net3894));
 sg13g2_o21ai_1 _14919_ (.B1(_07591_),
    .Y(_00730_),
    .A1(net4545),
    .A2(_03666_));
 sg13g2_nor2_1 _14920_ (.A(net4545),
    .B(net3893),
    .Y(_07592_));
 sg13g2_a21oi_1 _14921_ (.A1(net4545),
    .A2(_03666_),
    .Y(_00731_),
    .B1(_07592_));
 sg13g2_mux2_1 _14922_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[7] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[6] ),
    .S(net4546),
    .X(_00732_));
 sg13g2_mux2_1 _14923_ (.A0(net267),
    .A1(net105),
    .S(net4549),
    .X(_00733_));
 sg13g2_mux2_1 _14924_ (.A0(net3896),
    .A1(net3895),
    .S(\spiking_network_top_uut.all_data_out[824] ),
    .X(_07593_));
 sg13g2_nor2b_1 _14925_ (.A(\spiking_network_top_uut.all_data_out[824] ),
    .B_N(net3898),
    .Y(_07594_));
 sg13g2_a21oi_1 _14926_ (.A1(\spiking_network_top_uut.all_data_out[824] ),
    .A2(net3897),
    .Y(_07595_),
    .B1(_07594_));
 sg13g2_a21oi_1 _14927_ (.A1(\spiking_network_top_uut.all_data_out[825] ),
    .A2(_07593_),
    .Y(_07596_),
    .B1(\spiking_network_top_uut.all_data_out[826] ));
 sg13g2_o21ai_1 _14928_ (.B1(_07596_),
    .Y(_07597_),
    .A1(\spiking_network_top_uut.all_data_out[825] ),
    .A2(_07595_));
 sg13g2_mux2_1 _14929_ (.A0(net3893),
    .A1(net3892),
    .S(\spiking_network_top_uut.all_data_out[824] ),
    .X(_07598_));
 sg13g2_nand2_1 _14930_ (.Y(_07599_),
    .A(\spiking_network_top_uut.all_data_out[825] ),
    .B(_07598_));
 sg13g2_a21oi_1 _14931_ (.A1(\spiking_network_top_uut.all_data_out[824] ),
    .A2(_03666_),
    .Y(_07600_),
    .B1(\spiking_network_top_uut.all_data_out[825] ));
 sg13g2_o21ai_1 _14932_ (.B1(_07600_),
    .Y(_07601_),
    .A1(\spiking_network_top_uut.all_data_out[824] ),
    .A2(net3894));
 sg13g2_nand3_1 _14933_ (.B(_07599_),
    .C(_07601_),
    .A(\spiking_network_top_uut.all_data_out[826] ),
    .Y(_07602_));
 sg13g2_nand3_1 _14934_ (.B(_07597_),
    .C(_07602_),
    .A(net4546),
    .Y(_07603_));
 sg13g2_o21ai_1 _14935_ (.B1(_07603_),
    .Y(_00734_),
    .A1(net4546),
    .A2(_03681_));
 sg13g2_mux2_1 _14936_ (.A0(net3891),
    .A1(net4594),
    .S(net4556),
    .X(_00735_));
 sg13g2_mux2_1 _14937_ (.A0(net3890),
    .A1(net3891),
    .S(net4558),
    .X(_00736_));
 sg13g2_mux2_1 _14938_ (.A0(net3889),
    .A1(net3890),
    .S(net4560),
    .X(_00737_));
 sg13g2_mux2_1 _14939_ (.A0(net3888),
    .A1(net3889),
    .S(net4560),
    .X(_00738_));
 sg13g2_mux2_1 _14940_ (.A0(net3887),
    .A1(net3888),
    .S(net4560),
    .X(_00739_));
 sg13g2_nand2_1 _14941_ (.Y(_07604_),
    .A(net4559),
    .B(net3887));
 sg13g2_o21ai_1 _14942_ (.B1(_07604_),
    .Y(_00740_),
    .A1(net4559),
    .A2(_03665_));
 sg13g2_nor2_1 _14943_ (.A(net4559),
    .B(net3886),
    .Y(_07605_));
 sg13g2_a21oi_1 _14944_ (.A1(net4559),
    .A2(_03665_),
    .Y(_00741_),
    .B1(_07605_));
 sg13g2_mux2_1 _14945_ (.A0(net3885),
    .A1(net3886),
    .S(net4558),
    .X(_00742_));
 sg13g2_mux2_1 _14946_ (.A0(net242),
    .A1(net53),
    .S(net4549),
    .X(_00743_));
 sg13g2_mux4_1 _14947_ (.S0(\spiking_network_top_uut.all_data_out[820] ),
    .A0(net3891),
    .A1(net3890),
    .A2(net3889),
    .A3(net3888),
    .S1(\spiking_network_top_uut.all_data_out[821] ),
    .X(_07606_));
 sg13g2_mux2_1 _14948_ (.A0(net3886),
    .A1(net3885),
    .S(\spiking_network_top_uut.all_data_out[820] ),
    .X(_07607_));
 sg13g2_nor2b_1 _14949_ (.A(\spiking_network_top_uut.all_data_out[820] ),
    .B_N(net3887),
    .Y(_07608_));
 sg13g2_a21oi_1 _14950_ (.A1(\spiking_network_top_uut.all_data_out[820] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[5] ),
    .Y(_07609_),
    .B1(_07608_));
 sg13g2_o21ai_1 _14951_ (.B1(\spiking_network_top_uut.all_data_out[822] ),
    .Y(_07610_),
    .A1(\spiking_network_top_uut.all_data_out[821] ),
    .A2(_07609_));
 sg13g2_a21oi_1 _14952_ (.A1(\spiking_network_top_uut.all_data_out[821] ),
    .A2(_07607_),
    .Y(_07611_),
    .B1(_07610_));
 sg13g2_o21ai_1 _14953_ (.B1(net4561),
    .Y(_07612_),
    .A1(\spiking_network_top_uut.all_data_out[822] ),
    .A2(_07606_));
 sg13g2_nand2_1 _14954_ (.Y(_07613_),
    .A(net3935),
    .B(net95));
 sg13g2_o21ai_1 _14955_ (.B1(_07613_),
    .Y(_00744_),
    .A1(_07611_),
    .A2(_07612_));
 sg13g2_mux2_1 _14956_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[0] ),
    .A1(net4595),
    .S(net4556),
    .X(_00745_));
 sg13g2_mux2_1 _14957_ (.A0(net3883),
    .A1(net3884),
    .S(net4554),
    .X(_00746_));
 sg13g2_mux2_1 _14958_ (.A0(net3882),
    .A1(net3883),
    .S(net4554),
    .X(_00747_));
 sg13g2_mux2_1 _14959_ (.A0(net3881),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[2] ),
    .S(net4554),
    .X(_00748_));
 sg13g2_mux2_1 _14960_ (.A0(net3880),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[3] ),
    .S(net4556),
    .X(_00749_));
 sg13g2_mux2_1 _14961_ (.A0(net3879),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[4] ),
    .S(net4555),
    .X(_00750_));
 sg13g2_mux2_1 _14962_ (.A0(net3878),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[5] ),
    .S(net4555),
    .X(_00751_));
 sg13g2_mux2_1 _14963_ (.A0(net3877),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[6] ),
    .S(net4555),
    .X(_00752_));
 sg13g2_mux2_1 _14964_ (.A0(net478),
    .A1(net95),
    .S(net4561),
    .X(_00753_));
 sg13g2_nand2b_1 _14965_ (.Y(_07614_),
    .B(\spiking_network_top_uut.all_data_out[816] ),
    .A_N(net3879));
 sg13g2_nor2_1 _14966_ (.A(\spiking_network_top_uut.all_data_out[816] ),
    .B(net3880),
    .Y(_07615_));
 sg13g2_nor2_1 _14967_ (.A(\spiking_network_top_uut.all_data_out[817] ),
    .B(_07615_),
    .Y(_07616_));
 sg13g2_mux2_1 _14968_ (.A0(net3878),
    .A1(net3877),
    .S(\spiking_network_top_uut.all_data_out[816] ),
    .X(_07617_));
 sg13g2_a221oi_1 _14969_ (.B2(\spiking_network_top_uut.all_data_out[817] ),
    .C1(_03583_),
    .B1(_07617_),
    .A1(_07614_),
    .Y(_07618_),
    .A2(_07616_));
 sg13g2_mux4_1 _14970_ (.S0(\spiking_network_top_uut.all_data_out[816] ),
    .A0(net3884),
    .A1(net3883),
    .A2(net3882),
    .A3(net3881),
    .S1(\spiking_network_top_uut.all_data_out[817] ),
    .X(_07619_));
 sg13g2_o21ai_1 _14971_ (.B1(net4557),
    .Y(_07620_),
    .A1(\spiking_network_top_uut.all_data_out[818] ),
    .A2(_07619_));
 sg13g2_nand2_1 _14972_ (.Y(_07621_),
    .A(net3938),
    .B(net215));
 sg13g2_o21ai_1 _14973_ (.B1(_07621_),
    .Y(_00754_),
    .A1(_07618_),
    .A2(_07620_));
 sg13g2_mux2_1 _14974_ (.A0(net3876),
    .A1(net4596),
    .S(net4571),
    .X(_00755_));
 sg13g2_mux2_1 _14975_ (.A0(net3875),
    .A1(net3876),
    .S(net4567),
    .X(_00756_));
 sg13g2_mux2_1 _14976_ (.A0(net3874),
    .A1(net3875),
    .S(net4567),
    .X(_00757_));
 sg13g2_mux2_1 _14977_ (.A0(net3873),
    .A1(net3874),
    .S(net4567),
    .X(_00758_));
 sg13g2_mux2_1 _14978_ (.A0(net3872),
    .A1(net3873),
    .S(net4569),
    .X(_00759_));
 sg13g2_mux2_1 _14979_ (.A0(net3871),
    .A1(net3872),
    .S(net4569),
    .X(_00760_));
 sg13g2_mux2_1 _14980_ (.A0(net3870),
    .A1(net3871),
    .S(net4569),
    .X(_00761_));
 sg13g2_mux2_1 _14981_ (.A0(net3869),
    .A1(net3870),
    .S(net4569),
    .X(_00762_));
 sg13g2_mux2_1 _14982_ (.A0(net276),
    .A1(net215),
    .S(net4557),
    .X(_00763_));
 sg13g2_nand2b_1 _14983_ (.Y(_07622_),
    .B(\spiking_network_top_uut.all_data_out[812] ),
    .A_N(net3871));
 sg13g2_nor2_1 _14984_ (.A(\spiking_network_top_uut.all_data_out[812] ),
    .B(net3872),
    .Y(_07623_));
 sg13g2_nor2_1 _14985_ (.A(\spiking_network_top_uut.all_data_out[813] ),
    .B(_07623_),
    .Y(_07624_));
 sg13g2_mux2_1 _14986_ (.A0(net3870),
    .A1(net3869),
    .S(\spiking_network_top_uut.all_data_out[812] ),
    .X(_07625_));
 sg13g2_a221oi_1 _14987_ (.B2(\spiking_network_top_uut.all_data_out[813] ),
    .C1(_03511_),
    .B1(_07625_),
    .A1(_07622_),
    .Y(_07626_),
    .A2(_07624_));
 sg13g2_mux4_1 _14988_ (.S0(\spiking_network_top_uut.all_data_out[812] ),
    .A0(net3876),
    .A1(net3875),
    .A2(net3874),
    .A3(net3873),
    .S1(\spiking_network_top_uut.all_data_out[813] ),
    .X(_07627_));
 sg13g2_o21ai_1 _14989_ (.B1(net4566),
    .Y(_07628_),
    .A1(\spiking_network_top_uut.all_data_out[814] ),
    .A2(_07627_));
 sg13g2_nand2_1 _14990_ (.Y(_07629_),
    .A(net3937),
    .B(net72));
 sg13g2_o21ai_1 _14991_ (.B1(_07629_),
    .Y(_00764_),
    .A1(_07626_),
    .A2(_07628_));
 sg13g2_mux2_1 _14992_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[0] ),
    .A1(net4597),
    .S(net4564),
    .X(_00765_));
 sg13g2_mux2_1 _14993_ (.A0(net3867),
    .A1(net3868),
    .S(net4562),
    .X(_00766_));
 sg13g2_mux2_1 _14994_ (.A0(net3866),
    .A1(net3867),
    .S(net4563),
    .X(_00767_));
 sg13g2_mux2_1 _14995_ (.A0(net3865),
    .A1(net3866),
    .S(net4564),
    .X(_00768_));
 sg13g2_mux2_1 _14996_ (.A0(net3864),
    .A1(net3865),
    .S(net4562),
    .X(_00769_));
 sg13g2_mux2_1 _14997_ (.A0(net3863),
    .A1(net3864),
    .S(net4562),
    .X(_00770_));
 sg13g2_mux2_1 _14998_ (.A0(net3862),
    .A1(net3863),
    .S(net4562),
    .X(_00771_));
 sg13g2_mux2_1 _14999_ (.A0(net3861),
    .A1(net3862),
    .S(net4562),
    .X(_00772_));
 sg13g2_mux2_1 _15000_ (.A0(net245),
    .A1(net72),
    .S(net4567),
    .X(_00773_));
 sg13g2_mux4_1 _15001_ (.S0(\spiking_network_top_uut.all_data_out[808] ),
    .A0(net3868),
    .A1(net3867),
    .A2(net3866),
    .A3(net3865),
    .S1(\spiking_network_top_uut.all_data_out[809] ),
    .X(_07630_));
 sg13g2_mux2_1 _15002_ (.A0(net3862),
    .A1(net3861),
    .S(\spiking_network_top_uut.all_data_out[808] ),
    .X(_07631_));
 sg13g2_nor2b_1 _15003_ (.A(\spiking_network_top_uut.all_data_out[808] ),
    .B_N(net3864),
    .Y(_07632_));
 sg13g2_a21oi_1 _15004_ (.A1(\spiking_network_top_uut.all_data_out[808] ),
    .A2(net3863),
    .Y(_07633_),
    .B1(_07632_));
 sg13g2_o21ai_1 _15005_ (.B1(\spiking_network_top_uut.all_data_out[810] ),
    .Y(_07634_),
    .A1(\spiking_network_top_uut.all_data_out[809] ),
    .A2(_07633_));
 sg13g2_a21oi_1 _15006_ (.A1(\spiking_network_top_uut.all_data_out[809] ),
    .A2(_07631_),
    .Y(_07635_),
    .B1(_07634_));
 sg13g2_o21ai_1 _15007_ (.B1(net4563),
    .Y(_07636_),
    .A1(\spiking_network_top_uut.all_data_out[810] ),
    .A2(_07630_));
 sg13g2_nand2_1 _15008_ (.Y(_07637_),
    .A(net3936),
    .B(net169));
 sg13g2_o21ai_1 _15009_ (.B1(_07637_),
    .Y(_00774_),
    .A1(_07635_),
    .A2(_07636_));
 sg13g2_mux2_1 _15010_ (.A0(net3860),
    .A1(net4598),
    .S(net4534),
    .X(_00775_));
 sg13g2_mux2_1 _15011_ (.A0(net3859),
    .A1(net3860),
    .S(net4537),
    .X(_00776_));
 sg13g2_mux2_1 _15012_ (.A0(net3858),
    .A1(net3859),
    .S(net4535),
    .X(_00777_));
 sg13g2_mux2_1 _15013_ (.A0(net3857),
    .A1(net3858),
    .S(net4535),
    .X(_00778_));
 sg13g2_mux2_1 _15014_ (.A0(net3856),
    .A1(net3857),
    .S(net4535),
    .X(_00779_));
 sg13g2_nand2_1 _15015_ (.Y(_07638_),
    .A(net4541),
    .B(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[4] ));
 sg13g2_o21ai_1 _15016_ (.B1(_07638_),
    .Y(_00780_),
    .A1(net4541),
    .A2(_03664_));
 sg13g2_nor2_1 _15017_ (.A(net4535),
    .B(net3855),
    .Y(_07639_));
 sg13g2_a21oi_1 _15018_ (.A1(net4535),
    .A2(_03664_),
    .Y(_00781_),
    .B1(_07639_));
 sg13g2_mux2_1 _15019_ (.A0(net3854),
    .A1(net3855),
    .S(net4536),
    .X(_00782_));
 sg13g2_mux2_1 _15020_ (.A0(net255),
    .A1(net169),
    .S(net4563),
    .X(_00783_));
 sg13g2_mux2_1 _15021_ (.A0(net3858),
    .A1(net3857),
    .S(\spiking_network_top_uut.all_data_out[804] ),
    .X(_07640_));
 sg13g2_nor2b_1 _15022_ (.A(\spiking_network_top_uut.all_data_out[804] ),
    .B_N(net3860),
    .Y(_07641_));
 sg13g2_a21oi_1 _15023_ (.A1(\spiking_network_top_uut.all_data_out[804] ),
    .A2(net3859),
    .Y(_07642_),
    .B1(_07641_));
 sg13g2_a21oi_1 _15024_ (.A1(\spiking_network_top_uut.all_data_out[805] ),
    .A2(_07640_),
    .Y(_07643_),
    .B1(\spiking_network_top_uut.all_data_out[806] ));
 sg13g2_o21ai_1 _15025_ (.B1(_07643_),
    .Y(_07644_),
    .A1(\spiking_network_top_uut.all_data_out[805] ),
    .A2(_07642_));
 sg13g2_mux2_1 _15026_ (.A0(net3855),
    .A1(net3854),
    .S(\spiking_network_top_uut.all_data_out[804] ),
    .X(_07645_));
 sg13g2_nand2_1 _15027_ (.Y(_07646_),
    .A(\spiking_network_top_uut.all_data_out[805] ),
    .B(_07645_));
 sg13g2_a21oi_1 _15028_ (.A1(\spiking_network_top_uut.all_data_out[804] ),
    .A2(_03664_),
    .Y(_07647_),
    .B1(\spiking_network_top_uut.all_data_out[805] ));
 sg13g2_o21ai_1 _15029_ (.B1(_07647_),
    .Y(_07648_),
    .A1(\spiking_network_top_uut.all_data_out[804] ),
    .A2(net3856));
 sg13g2_nand3_1 _15030_ (.B(_07646_),
    .C(_07648_),
    .A(\spiking_network_top_uut.all_data_out[806] ),
    .Y(_07649_));
 sg13g2_nand3_1 _15031_ (.B(_07644_),
    .C(_07649_),
    .A(net4534),
    .Y(_07650_));
 sg13g2_o21ai_1 _15032_ (.B1(_07650_),
    .Y(_00784_),
    .A1(net4534),
    .A2(_03682_));
 sg13g2_mux2_1 _15033_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[0] ),
    .A1(net4599),
    .S(net4544),
    .X(_00785_));
 sg13g2_mux2_1 _15034_ (.A0(net3852),
    .A1(net3853),
    .S(net4543),
    .X(_00786_));
 sg13g2_mux2_1 _15035_ (.A0(net3851),
    .A1(net3852),
    .S(net4543),
    .X(_00787_));
 sg13g2_mux2_1 _15036_ (.A0(net3850),
    .A1(net3851),
    .S(net4543),
    .X(_00788_));
 sg13g2_mux2_1 _15037_ (.A0(net3849),
    .A1(net3850),
    .S(net4538),
    .X(_00789_));
 sg13g2_nand2_1 _15038_ (.Y(_07651_),
    .A(net4538),
    .B(net3849));
 sg13g2_o21ai_1 _15039_ (.B1(_07651_),
    .Y(_00790_),
    .A1(net4538),
    .A2(_03663_));
 sg13g2_nor2_1 _15040_ (.A(net4538),
    .B(net3848),
    .Y(_07652_));
 sg13g2_a21oi_1 _15041_ (.A1(net4538),
    .A2(_03663_),
    .Y(_00791_),
    .B1(_07652_));
 sg13g2_mux2_1 _15042_ (.A0(net3847),
    .A1(net3848),
    .S(net4538),
    .X(_00792_));
 sg13g2_mux2_1 _15043_ (.A0(net207),
    .A1(net94),
    .S(net4534),
    .X(_00793_));
 sg13g2_nand2_1 _15044_ (.Y(_07653_),
    .A(\spiking_network_top_uut.all_data_out[800] ),
    .B(_03663_));
 sg13g2_nor2_1 _15045_ (.A(\spiking_network_top_uut.all_data_out[800] ),
    .B(net3849),
    .Y(_07654_));
 sg13g2_nor2_1 _15046_ (.A(\spiking_network_top_uut.all_data_out[801] ),
    .B(_07654_),
    .Y(_07655_));
 sg13g2_mux2_1 _15047_ (.A0(net3848),
    .A1(net3847),
    .S(\spiking_network_top_uut.all_data_out[800] ),
    .X(_07656_));
 sg13g2_a221oi_1 _15048_ (.B2(\spiking_network_top_uut.all_data_out[801] ),
    .C1(_03585_),
    .B1(_07656_),
    .A1(_07653_),
    .Y(_07657_),
    .A2(_07655_));
 sg13g2_mux4_1 _15049_ (.S0(\spiking_network_top_uut.all_data_out[800] ),
    .A0(net3853),
    .A1(net3852),
    .A2(net3851),
    .A3(net3850),
    .S1(\spiking_network_top_uut.all_data_out[801] ),
    .X(_07658_));
 sg13g2_o21ai_1 _15050_ (.B1(net4544),
    .Y(_07659_),
    .A1(\spiking_network_top_uut.all_data_out[802] ),
    .A2(_07658_));
 sg13g2_nand2_1 _15051_ (.Y(_07660_),
    .A(net3933),
    .B(net527));
 sg13g2_o21ai_1 _15052_ (.B1(_07660_),
    .Y(_00794_),
    .A1(_07657_),
    .A2(_07659_));
 sg13g2_nor3_2 _15053_ (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[2] ),
    .B(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[1] ),
    .C(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[0] ),
    .Y(_07661_));
 sg13g2_nor2b_2 _15054_ (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[3] ),
    .B_N(_07661_),
    .Y(_07662_));
 sg13g2_nor2b_2 _15055_ (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[4] ),
    .B_N(_07662_),
    .Y(_07663_));
 sg13g2_nand2b_2 _15056_ (.Y(_07664_),
    .B(_07662_),
    .A_N(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[4] ));
 sg13g2_o21ai_1 _15057_ (.B1(net4531),
    .Y(_07665_),
    .A1(net3623),
    .A2(_07664_));
 sg13g2_nor2b_1 _15058_ (.A(net3623),
    .B_N(_00090_),
    .Y(_07666_));
 sg13g2_a21oi_1 _15059_ (.A1(net4283),
    .A2(net3623),
    .Y(_07667_),
    .B1(_07666_));
 sg13g2_nand2_1 _15060_ (.Y(_07668_),
    .A(net365),
    .B(_07665_));
 sg13g2_o21ai_1 _15061_ (.B1(_07668_),
    .Y(_00795_),
    .A1(_07665_),
    .A2(_07667_));
 sg13g2_xor2_1 _15062_ (.B(net365),
    .A(net397),
    .X(_07669_));
 sg13g2_nor2_1 _15063_ (.A(net3623),
    .B(_07669_),
    .Y(_07670_));
 sg13g2_a21oi_1 _15064_ (.A1(net4280),
    .A2(net3623),
    .Y(_07671_),
    .B1(_07670_));
 sg13g2_nand2_1 _15065_ (.Y(_07672_),
    .A(net397),
    .B(_07665_));
 sg13g2_o21ai_1 _15066_ (.B1(_07672_),
    .Y(_00796_),
    .A1(_07665_),
    .A2(_07671_));
 sg13g2_o21ai_1 _15067_ (.B1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[2] ),
    .Y(_07673_),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[1] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[0] ));
 sg13g2_nor2b_1 _15068_ (.A(_07661_),
    .B_N(_07673_),
    .Y(_07674_));
 sg13g2_nor2_1 _15069_ (.A(net3623),
    .B(_07674_),
    .Y(_07675_));
 sg13g2_a21oi_1 _15070_ (.A1(net4276),
    .A2(net3623),
    .Y(_07676_),
    .B1(_07675_));
 sg13g2_nand2_1 _15071_ (.Y(_07677_),
    .A(net210),
    .B(_07665_));
 sg13g2_o21ai_1 _15072_ (.B1(_07677_),
    .Y(_00797_),
    .A1(_07665_),
    .A2(_07676_));
 sg13g2_nand2_1 _15073_ (.Y(_07678_),
    .A(net4273),
    .B(net3623));
 sg13g2_xnor2_1 _15074_ (.Y(_07679_),
    .A(net441),
    .B(_07661_));
 sg13g2_o21ai_1 _15075_ (.B1(_07678_),
    .Y(_07680_),
    .A1(net3624),
    .A2(_07679_));
 sg13g2_mux2_1 _15076_ (.A0(_07680_),
    .A1(net441),
    .S(_07665_),
    .X(_00798_));
 sg13g2_nand2_1 _15077_ (.Y(_07681_),
    .A(net3923),
    .B(net312));
 sg13g2_nand2b_1 _15078_ (.Y(_07682_),
    .B(net312),
    .A_N(_07662_));
 sg13g2_a21oi_1 _15079_ (.A1(_07664_),
    .A2(_07682_),
    .Y(_07683_),
    .B1(net3624));
 sg13g2_a21oi_1 _15080_ (.A1(net4270),
    .A2(net3624),
    .Y(_07684_),
    .B1(_07683_));
 sg13g2_o21ai_1 _15081_ (.B1(_07681_),
    .Y(_00799_),
    .A1(_07665_),
    .A2(_07684_));
 sg13g2_mux2_1 _15082_ (.A0(net196),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_reg1 ),
    .S(net4536),
    .X(_00800_));
 sg13g2_mux2_1 _15083_ (.A0(net3846),
    .A1(net4592),
    .S(net4549),
    .X(_00801_));
 sg13g2_mux2_1 _15084_ (.A0(net3845),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[0] ),
    .S(net4551),
    .X(_00802_));
 sg13g2_mux2_1 _15085_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[2] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[1] ),
    .S(net4550),
    .X(_00803_));
 sg13g2_mux2_1 _15086_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[3] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[2] ),
    .S(net4552),
    .X(_00804_));
 sg13g2_mux2_1 _15087_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[4] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[3] ),
    .S(net4550),
    .X(_00805_));
 sg13g2_nand2_1 _15088_ (.Y(_07685_),
    .A(net4550),
    .B(net3842));
 sg13g2_o21ai_1 _15089_ (.B1(_07685_),
    .Y(_00806_),
    .A1(net4550),
    .A2(_03667_));
 sg13g2_nor2_1 _15090_ (.A(net4550),
    .B(net3841),
    .Y(_07686_));
 sg13g2_a21oi_1 _15091_ (.A1(net4550),
    .A2(_03667_),
    .Y(_00807_),
    .B1(_07686_));
 sg13g2_a21oi_1 _15092_ (.A1(net3915),
    .A2(net3911),
    .Y(_07687_),
    .B1(_00085_));
 sg13g2_nor2_2 _15093_ (.A(net3752),
    .B(_07687_),
    .Y(_07688_));
 sg13g2_nor2_1 _15094_ (.A(_00085_),
    .B(_07688_),
    .Y(_07689_));
 sg13g2_nand2b_1 _15095_ (.Y(_07690_),
    .B(_07688_),
    .A_N(_00085_));
 sg13g2_o21ai_1 _15096_ (.B1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ),
    .Y(_07691_),
    .A1(_00085_),
    .A2(_07688_));
 sg13g2_inv_1 _15097_ (.Y(_07692_),
    .A(_07691_));
 sg13g2_a21o_1 _15098_ (.A2(net3754),
    .A1(_00086_),
    .B1(_07688_),
    .X(_07693_));
 sg13g2_nor2_1 _15099_ (.A(_00086_),
    .B(net3908),
    .Y(_07694_));
 sg13g2_a221oi_1 _15100_ (.B2(_07687_),
    .C1(_07694_),
    .B1(net3908),
    .A1(_03489_),
    .Y(_07695_),
    .A2(net3754));
 sg13g2_nand2_1 _15101_ (.Y(_07696_),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ),
    .B(_07695_));
 sg13g2_nor2_1 _15102_ (.A(_00085_),
    .B(net3911),
    .Y(_07697_));
 sg13g2_a21o_1 _15103_ (.A2(_00086_),
    .A1(net4267),
    .B1(_05084_),
    .X(_07698_));
 sg13g2_a21oi_1 _15104_ (.A1(_03489_),
    .A2(net3739),
    .Y(_07699_),
    .B1(_07697_));
 sg13g2_a22oi_1 _15105_ (.Y(_07700_),
    .B1(_07698_),
    .B2(_07699_),
    .A2(net3754),
    .A1(_00089_));
 sg13g2_a221oi_1 _15106_ (.B2(_07699_),
    .C1(_03490_),
    .B1(_07698_),
    .A1(_00089_),
    .Y(_07701_),
    .A2(net3754));
 sg13g2_xnor2_1 _15107_ (.Y(_07702_),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ),
    .B(_07695_));
 sg13g2_o21ai_1 _15108_ (.B1(_07696_),
    .Y(_07703_),
    .A1(_07701_),
    .A2(_07702_));
 sg13g2_xnor2_1 _15109_ (.Y(_07704_),
    .A(_03489_),
    .B(_07693_));
 sg13g2_nor2b_1 _15110_ (.A(_07704_),
    .B_N(_07703_),
    .Y(_07705_));
 sg13g2_a21o_1 _15111_ (.A2(_07693_),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ),
    .B1(_07705_),
    .X(_07706_));
 sg13g2_xnor2_1 _15112_ (.Y(_07707_),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ),
    .B(_07689_));
 sg13g2_a21oi_1 _15113_ (.A1(_07706_),
    .A2(_07707_),
    .Y(_07708_),
    .B1(_07692_));
 sg13g2_a22oi_1 _15114_ (.Y(_07709_),
    .B1(_07690_),
    .B2(_07708_),
    .A2(_07688_),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ));
 sg13g2_a21oi_2 _15115_ (.B1(_07709_),
    .Y(_07710_),
    .A2(_00085_),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ));
 sg13g2_nor2_1 _15116_ (.A(_07663_),
    .B(_07710_),
    .Y(_07711_));
 sg13g2_mux2_1 _15117_ (.A0(net4599),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[803] ),
    .X(_07712_));
 sg13g2_nand2_1 _15118_ (.Y(_07713_),
    .A(\spiking_network_top_uut.all_data_out[273] ),
    .B(_07712_));
 sg13g2_mux2_1 _15119_ (.A0(net4598),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[807] ),
    .X(_07714_));
 sg13g2_nand2_1 _15120_ (.Y(_07715_),
    .A(\spiking_network_top_uut.all_data_out[275] ),
    .B(_07714_));
 sg13g2_nor2_1 _15121_ (.A(_07713_),
    .B(_07715_),
    .Y(_07716_));
 sg13g2_and4_1 _15122_ (.A(\spiking_network_top_uut.all_data_out[272] ),
    .B(\spiking_network_top_uut.all_data_out[274] ),
    .C(_07712_),
    .D(_07714_),
    .X(_07717_));
 sg13g2_nand4_1 _15123_ (.B(\spiking_network_top_uut.all_data_out[274] ),
    .C(_07712_),
    .A(\spiking_network_top_uut.all_data_out[272] ),
    .Y(_07718_),
    .D(_07714_));
 sg13g2_xor2_1 _15124_ (.B(_07715_),
    .A(_07713_),
    .X(_07719_));
 sg13g2_a21oi_2 _15125_ (.B1(_07716_),
    .Y(_07720_),
    .A2(_07719_),
    .A1(_07718_));
 sg13g2_mux2_2 _15126_ (.A0(net4597),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[811] ),
    .X(_07721_));
 sg13g2_nand2_1 _15127_ (.Y(_07722_),
    .A(\spiking_network_top_uut.all_data_out[277] ),
    .B(_07721_));
 sg13g2_mux2_2 _15128_ (.A0(net4596),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[815] ),
    .X(_07723_));
 sg13g2_nand2_1 _15129_ (.Y(_07724_),
    .A(\spiking_network_top_uut.all_data_out[279] ),
    .B(_07723_));
 sg13g2_nor2_1 _15130_ (.A(_07722_),
    .B(_07724_),
    .Y(_07725_));
 sg13g2_nand2_1 _15131_ (.Y(_07726_),
    .A(\spiking_network_top_uut.all_data_out[276] ),
    .B(_07721_));
 sg13g2_nand2_1 _15132_ (.Y(_07727_),
    .A(\spiking_network_top_uut.all_data_out[278] ),
    .B(_07723_));
 sg13g2_or2_1 _15133_ (.X(_07728_),
    .B(_07727_),
    .A(_07726_));
 sg13g2_xor2_1 _15134_ (.B(_07724_),
    .A(_07722_),
    .X(_07729_));
 sg13g2_a21oi_2 _15135_ (.B1(_07725_),
    .Y(_07730_),
    .A2(_07729_),
    .A1(_07728_));
 sg13g2_mux2_2 _15136_ (.A0(net4595),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[819] ),
    .X(_07731_));
 sg13g2_mux2_2 _15137_ (.A0(net4594),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[823] ),
    .X(_07732_));
 sg13g2_a22oi_1 _15138_ (.Y(_07733_),
    .B1(_07732_),
    .B2(\spiking_network_top_uut.all_data_out[283] ),
    .A2(_07731_),
    .A1(\spiking_network_top_uut.all_data_out[281] ));
 sg13g2_and4_1 _15139_ (.A(\spiking_network_top_uut.all_data_out[280] ),
    .B(\spiking_network_top_uut.all_data_out[282] ),
    .C(_07731_),
    .D(_07732_),
    .X(_07734_));
 sg13g2_and4_1 _15140_ (.A(\spiking_network_top_uut.all_data_out[281] ),
    .B(\spiking_network_top_uut.all_data_out[283] ),
    .C(_07731_),
    .D(_07732_),
    .X(_07735_));
 sg13g2_nand4_1 _15141_ (.B(\spiking_network_top_uut.all_data_out[283] ),
    .C(_07731_),
    .A(\spiking_network_top_uut.all_data_out[281] ),
    .Y(_07736_),
    .D(_07732_));
 sg13g2_a21oi_2 _15142_ (.B1(_07733_),
    .Y(_07737_),
    .A2(_07736_),
    .A1(_07734_));
 sg13g2_mux2_2 _15143_ (.A0(net4593),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[827] ),
    .X(_07738_));
 sg13g2_mux2_2 _15144_ (.A0(net4592),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[831] ),
    .X(_07739_));
 sg13g2_and4_1 _15145_ (.A(\spiking_network_top_uut.all_data_out[285] ),
    .B(\spiking_network_top_uut.all_data_out[287] ),
    .C(_07738_),
    .D(_07739_),
    .X(_07740_));
 sg13g2_nand4_1 _15146_ (.B(\spiking_network_top_uut.all_data_out[287] ),
    .C(_07738_),
    .A(\spiking_network_top_uut.all_data_out[285] ),
    .Y(_07741_),
    .D(_07739_));
 sg13g2_and4_1 _15147_ (.A(\spiking_network_top_uut.all_data_out[284] ),
    .B(\spiking_network_top_uut.all_data_out[286] ),
    .C(_07738_),
    .D(_07739_),
    .X(_07742_));
 sg13g2_a22oi_1 _15148_ (.Y(_07743_),
    .B1(_07739_),
    .B2(\spiking_network_top_uut.all_data_out[287] ),
    .A2(_07738_),
    .A1(\spiking_network_top_uut.all_data_out[285] ));
 sg13g2_or3_1 _15149_ (.A(_07740_),
    .B(_07742_),
    .C(_07743_),
    .X(_07744_));
 sg13g2_o21ai_1 _15150_ (.B1(_07741_),
    .Y(_07745_),
    .A1(_07742_),
    .A2(_07743_));
 sg13g2_nand3b_1 _15151_ (.B(_07737_),
    .C(_07745_),
    .Y(_07746_),
    .A_N(_07730_));
 sg13g2_inv_1 _15152_ (.Y(_07747_),
    .A(_07746_));
 sg13g2_or2_1 _15153_ (.X(_07748_),
    .B(_07746_),
    .A(_07720_));
 sg13g2_nor2_1 _15154_ (.A(_07737_),
    .B(_07745_),
    .Y(_07749_));
 sg13g2_and2_1 _15155_ (.A(_07730_),
    .B(_07749_),
    .X(_07750_));
 sg13g2_nand2_1 _15156_ (.Y(_07751_),
    .A(_07720_),
    .B(_07750_));
 sg13g2_and2_1 _15157_ (.A(_07748_),
    .B(_07751_),
    .X(_07752_));
 sg13g2_xnor2_1 _15158_ (.Y(_07753_),
    .A(_07690_),
    .B(_07708_));
 sg13g2_nand2_1 _15159_ (.Y(_07754_),
    .A(_07752_),
    .B(_07753_));
 sg13g2_nand2_1 _15160_ (.Y(_07755_),
    .A(_07748_),
    .B(_07754_));
 sg13g2_xor2_1 _15161_ (.B(_07752_),
    .A(_07710_),
    .X(_07756_));
 sg13g2_nand2_1 _15162_ (.Y(_07757_),
    .A(_07755_),
    .B(_07756_));
 sg13g2_xor2_1 _15163_ (.B(_07753_),
    .A(_07752_),
    .X(_07758_));
 sg13g2_o21ai_1 _15164_ (.B1(_07742_),
    .Y(_07759_),
    .A1(_07740_),
    .A2(_07743_));
 sg13g2_o21ai_1 _15165_ (.B1(_07734_),
    .Y(_07760_),
    .A1(_07733_),
    .A2(_07735_));
 sg13g2_or3_1 _15166_ (.A(_07733_),
    .B(_07734_),
    .C(_07735_),
    .X(_07761_));
 sg13g2_a22oi_1 _15167_ (.Y(_07762_),
    .B1(_07760_),
    .B2(_07761_),
    .A2(_07759_),
    .A1(_07744_));
 sg13g2_xor2_1 _15168_ (.B(_07729_),
    .A(_07728_),
    .X(_07763_));
 sg13g2_xnor2_1 _15169_ (.Y(_07764_),
    .A(_07728_),
    .B(_07729_));
 sg13g2_and4_1 _15170_ (.A(_07744_),
    .B(_07759_),
    .C(_07760_),
    .D(_07761_),
    .X(_07765_));
 sg13g2_nand4_1 _15171_ (.B(_07759_),
    .C(_07760_),
    .A(_07744_),
    .Y(_07766_),
    .D(_07761_));
 sg13g2_nand3b_1 _15172_ (.B(_07764_),
    .C(_07766_),
    .Y(_07767_),
    .A_N(_07762_));
 sg13g2_a21oi_2 _15173_ (.B1(_07762_),
    .Y(_07768_),
    .A2(_07766_),
    .A1(_07764_));
 sg13g2_xor2_1 _15174_ (.B(_07745_),
    .A(_07737_),
    .X(_07769_));
 sg13g2_xnor2_1 _15175_ (.Y(_07770_),
    .A(_07730_),
    .B(_07769_));
 sg13g2_nand2b_1 _15176_ (.Y(_07771_),
    .B(_07770_),
    .A_N(_07768_));
 sg13g2_xnor2_1 _15177_ (.Y(_07772_),
    .A(_07768_),
    .B(_07770_));
 sg13g2_nand2b_1 _15178_ (.Y(_07773_),
    .B(_07772_),
    .A_N(_07720_));
 sg13g2_nand2_1 _15179_ (.Y(_07774_),
    .A(_07771_),
    .B(_07773_));
 sg13g2_nor2_1 _15180_ (.A(_07747_),
    .B(_07750_),
    .Y(_07775_));
 sg13g2_xnor2_1 _15181_ (.Y(_07776_),
    .A(_07720_),
    .B(_07775_));
 sg13g2_and2_1 _15182_ (.A(_07774_),
    .B(_07776_),
    .X(_07777_));
 sg13g2_xor2_1 _15183_ (.B(_07776_),
    .A(_07774_),
    .X(_07778_));
 sg13g2_xnor2_1 _15184_ (.Y(_07779_),
    .A(_07706_),
    .B(_07707_));
 sg13g2_inv_1 _15185_ (.Y(_07780_),
    .A(_07779_));
 sg13g2_a21o_1 _15186_ (.A2(_07780_),
    .A1(_07778_),
    .B1(_07777_),
    .X(_07781_));
 sg13g2_and2_1 _15187_ (.A(_07758_),
    .B(_07781_),
    .X(_07782_));
 sg13g2_a22oi_1 _15188_ (.Y(_07783_),
    .B1(_07739_),
    .B2(\spiking_network_top_uut.all_data_out[286] ),
    .A2(_07738_),
    .A1(\spiking_network_top_uut.all_data_out[284] ));
 sg13g2_nor2_1 _15189_ (.A(_07742_),
    .B(_07783_),
    .Y(_07784_));
 sg13g2_a22oi_1 _15190_ (.Y(_07785_),
    .B1(_07732_),
    .B2(\spiking_network_top_uut.all_data_out[282] ),
    .A2(_07731_),
    .A1(\spiking_network_top_uut.all_data_out[280] ));
 sg13g2_nor2_1 _15191_ (.A(_07734_),
    .B(_07785_),
    .Y(_07786_));
 sg13g2_and2_1 _15192_ (.A(_07784_),
    .B(_07786_),
    .X(_07787_));
 sg13g2_xor2_1 _15193_ (.B(_07727_),
    .A(_07726_),
    .X(_07788_));
 sg13g2_xor2_1 _15194_ (.B(_07786_),
    .A(_07784_),
    .X(_07789_));
 sg13g2_a21o_2 _15195_ (.A2(_07789_),
    .A1(_07788_),
    .B1(_07787_),
    .X(_07790_));
 sg13g2_o21ai_1 _15196_ (.B1(_07763_),
    .Y(_07791_),
    .A1(_07762_),
    .A2(_07765_));
 sg13g2_nand3_1 _15197_ (.B(_07790_),
    .C(_07791_),
    .A(_07767_),
    .Y(_07792_));
 sg13g2_xnor2_1 _15198_ (.Y(_07793_),
    .A(_07717_),
    .B(_07719_));
 sg13g2_inv_1 _15199_ (.Y(_07794_),
    .A(_07793_));
 sg13g2_a21oi_1 _15200_ (.A1(_07767_),
    .A2(_07791_),
    .Y(_07795_),
    .B1(_07790_));
 sg13g2_a21o_1 _15201_ (.A2(_07791_),
    .A1(_07767_),
    .B1(_07790_),
    .X(_07796_));
 sg13g2_nand3_1 _15202_ (.B(_07794_),
    .C(_07796_),
    .A(_07792_),
    .Y(_07797_));
 sg13g2_o21ai_1 _15203_ (.B1(_07792_),
    .Y(_07798_),
    .A1(_07793_),
    .A2(_07795_));
 sg13g2_xnor2_1 _15204_ (.Y(_07799_),
    .A(_07720_),
    .B(_07772_));
 sg13g2_nand2_1 _15205_ (.Y(_07800_),
    .A(_07798_),
    .B(_07799_));
 sg13g2_xnor2_1 _15206_ (.Y(_07801_),
    .A(_07798_),
    .B(_07799_));
 sg13g2_xor2_1 _15207_ (.B(_07704_),
    .A(_07703_),
    .X(_07802_));
 sg13g2_o21ai_1 _15208_ (.B1(_07800_),
    .Y(_07803_),
    .A1(_07801_),
    .A2(_07802_));
 sg13g2_xnor2_1 _15209_ (.Y(_07804_),
    .A(_07778_),
    .B(_07780_));
 sg13g2_nand2b_1 _15210_ (.Y(_07805_),
    .B(_07803_),
    .A_N(_07804_));
 sg13g2_a22oi_1 _15211_ (.Y(_07806_),
    .B1(_07714_),
    .B2(\spiking_network_top_uut.all_data_out[274] ),
    .A2(_07712_),
    .A1(\spiking_network_top_uut.all_data_out[272] ));
 sg13g2_xnor2_1 _15212_ (.Y(_07807_),
    .A(_07788_),
    .B(_07789_));
 sg13g2_nor3_2 _15213_ (.A(_07717_),
    .B(_07806_),
    .C(_07807_),
    .Y(_07808_));
 sg13g2_a21o_1 _15214_ (.A2(_07796_),
    .A1(_07792_),
    .B1(_07794_),
    .X(_07809_));
 sg13g2_nand3_1 _15215_ (.B(_07808_),
    .C(_07809_),
    .A(_07797_),
    .Y(_07810_));
 sg13g2_a21oi_1 _15216_ (.A1(_07797_),
    .A2(_07809_),
    .Y(_07811_),
    .B1(_07808_));
 sg13g2_a21o_1 _15217_ (.A2(_07809_),
    .A1(_07797_),
    .B1(_07808_),
    .X(_07812_));
 sg13g2_xnor2_1 _15218_ (.Y(_07813_),
    .A(_07701_),
    .B(_07702_));
 sg13g2_inv_1 _15219_ (.Y(_07814_),
    .A(_07813_));
 sg13g2_nand3_1 _15220_ (.B(_07812_),
    .C(_07814_),
    .A(_07810_),
    .Y(_07815_));
 sg13g2_o21ai_1 _15221_ (.B1(_07810_),
    .Y(_07816_),
    .A1(_07811_),
    .A2(_07813_));
 sg13g2_xor2_1 _15222_ (.B(_07802_),
    .A(_07801_),
    .X(_07817_));
 sg13g2_and2_1 _15223_ (.A(_07816_),
    .B(_07817_),
    .X(_07818_));
 sg13g2_a21o_1 _15224_ (.A2(_07812_),
    .A1(_07810_),
    .B1(_07814_),
    .X(_07819_));
 sg13g2_o21ai_1 _15225_ (.B1(_07807_),
    .Y(_07820_),
    .A1(_07717_),
    .A2(_07806_));
 sg13g2_nand2b_1 _15226_ (.Y(_07821_),
    .B(_07820_),
    .A_N(_07808_));
 sg13g2_xnor2_1 _15227_ (.Y(_07822_),
    .A(_03490_),
    .B(_07700_));
 sg13g2_nor2_1 _15228_ (.A(_07821_),
    .B(_07822_),
    .Y(_07823_));
 sg13g2_and3_1 _15229_ (.X(_07824_),
    .A(_07815_),
    .B(_07819_),
    .C(_07823_));
 sg13g2_or2_1 _15230_ (.X(_07825_),
    .B(_07817_),
    .A(_07816_));
 sg13g2_nand2b_1 _15231_ (.Y(_07826_),
    .B(_07825_),
    .A_N(_07818_));
 sg13g2_a21oi_1 _15232_ (.A1(_07824_),
    .A2(_07825_),
    .Y(_07827_),
    .B1(_07818_));
 sg13g2_xor2_1 _15233_ (.B(_07804_),
    .A(_07803_),
    .X(_07828_));
 sg13g2_o21ai_1 _15234_ (.B1(_07805_),
    .Y(_07829_),
    .A1(_07827_),
    .A2(_07828_));
 sg13g2_or2_1 _15235_ (.X(_07830_),
    .B(_07781_),
    .A(_07758_));
 sg13g2_nand2b_1 _15236_ (.Y(_07831_),
    .B(_07830_),
    .A_N(_07782_));
 sg13g2_a21oi_1 _15237_ (.A1(_07829_),
    .A2(_07830_),
    .Y(_07832_),
    .B1(_07782_));
 sg13g2_xnor2_1 _15238_ (.Y(_07833_),
    .A(_07755_),
    .B(_07756_));
 sg13g2_o21ai_1 _15239_ (.B1(_07757_),
    .Y(_07834_),
    .A1(_07832_),
    .A2(_07833_));
 sg13g2_mux2_1 _15240_ (.A0(_07751_),
    .A1(_07748_),
    .S(_07710_),
    .X(_07835_));
 sg13g2_xnor2_1 _15241_ (.Y(_07836_),
    .A(_07834_),
    .B(_07835_));
 sg13g2_a21oi_2 _15242_ (.B1(_07711_),
    .Y(_07837_),
    .A2(_07836_),
    .A1(net3703));
 sg13g2_xnor2_1 _15243_ (.Y(_07838_),
    .A(_07832_),
    .B(_07833_));
 sg13g2_a21oi_1 _15244_ (.A1(net3703),
    .A2(_07838_),
    .Y(_07839_),
    .B1(_07711_));
 sg13g2_nor2_1 _15245_ (.A(net3703),
    .B(_07753_),
    .Y(_07840_));
 sg13g2_xor2_1 _15246_ (.B(_07831_),
    .A(_07829_),
    .X(_07841_));
 sg13g2_a21oi_1 _15247_ (.A1(net3703),
    .A2(_07841_),
    .Y(_07842_),
    .B1(_07840_));
 sg13g2_nand2_1 _15248_ (.Y(_07843_),
    .A(_07839_),
    .B(_07842_));
 sg13g2_a21oi_2 _15249_ (.B1(net3625),
    .Y(_07844_),
    .A2(_07843_),
    .A1(_07837_));
 sg13g2_nor2_1 _15250_ (.A(_07839_),
    .B(_07842_),
    .Y(_07845_));
 sg13g2_nor2_2 _15251_ (.A(_07837_),
    .B(_07845_),
    .Y(_07846_));
 sg13g2_nor2_1 _15252_ (.A(_07664_),
    .B(_07821_),
    .Y(_07847_));
 sg13g2_xnor2_1 _15253_ (.Y(_07848_),
    .A(_07822_),
    .B(_07847_));
 sg13g2_o21ai_1 _15254_ (.B1(_07844_),
    .Y(_07849_),
    .A1(_07846_),
    .A2(_07848_));
 sg13g2_xor2_1 _15255_ (.B(net451),
    .A(net4316),
    .X(_07850_));
 sg13g2_a21oi_1 _15256_ (.A1(net3625),
    .A2(_07850_),
    .Y(_07851_),
    .B1(net3928));
 sg13g2_a22oi_1 _15257_ (.Y(_00808_),
    .B1(_07849_),
    .B2(_07851_),
    .A2(_03427_),
    .A1(net3928));
 sg13g2_nor2_1 _15258_ (.A(net3703),
    .B(_07813_),
    .Y(_07852_));
 sg13g2_a21oi_1 _15259_ (.A1(_07815_),
    .A2(_07819_),
    .Y(_07853_),
    .B1(_07823_));
 sg13g2_nor3_1 _15260_ (.A(_07664_),
    .B(_07824_),
    .C(_07853_),
    .Y(_07854_));
 sg13g2_nor3_1 _15261_ (.A(_07846_),
    .B(_07852_),
    .C(_07854_),
    .Y(_07855_));
 sg13g2_nand2_1 _15262_ (.Y(_07856_),
    .A(net4533),
    .B(_07844_));
 sg13g2_xor2_1 _15263_ (.B(_04848_),
    .A(_04847_),
    .X(_07857_));
 sg13g2_a22oi_1 _15264_ (.Y(_07858_),
    .B1(_00016_),
    .B2(_07857_),
    .A2(net548),
    .A1(net3931));
 sg13g2_o21ai_1 _15265_ (.B1(_07858_),
    .Y(_00809_),
    .A1(_07855_),
    .A2(_07856_));
 sg13g2_xnor2_1 _15266_ (.Y(_07859_),
    .A(_07824_),
    .B(_07826_));
 sg13g2_nand2_1 _15267_ (.Y(_07860_),
    .A(net3703),
    .B(_07859_));
 sg13g2_o21ai_1 _15268_ (.B1(_07860_),
    .Y(_07861_),
    .A1(_07663_),
    .A2(_07802_));
 sg13g2_o21ai_1 _15269_ (.B1(_07844_),
    .Y(_07862_),
    .A1(_07846_),
    .A2(_07861_));
 sg13g2_xnor2_1 _15270_ (.Y(_07863_),
    .A(_04845_),
    .B(_04849_));
 sg13g2_a21oi_1 _15271_ (.A1(net3625),
    .A2(_07863_),
    .Y(_07864_),
    .B1(net3928));
 sg13g2_a22oi_1 _15272_ (.Y(_00810_),
    .B1(_07862_),
    .B2(_07864_),
    .A2(_03426_),
    .A1(net3928));
 sg13g2_nor2_1 _15273_ (.A(net3703),
    .B(_07780_),
    .Y(_07865_));
 sg13g2_xnor2_1 _15274_ (.Y(_07866_),
    .A(_07827_),
    .B(_07828_));
 sg13g2_a21oi_1 _15275_ (.A1(net3703),
    .A2(_07866_),
    .Y(_07867_),
    .B1(_07865_));
 sg13g2_o21ai_1 _15276_ (.B1(_07844_),
    .Y(_07868_),
    .A1(_07846_),
    .A2(_07867_));
 sg13g2_or3_1 _15277_ (.A(_04843_),
    .B(_04844_),
    .C(_04850_),
    .X(_07869_));
 sg13g2_and2_1 _15278_ (.A(_04851_),
    .B(_07869_),
    .X(_07870_));
 sg13g2_a21oi_1 _15279_ (.A1(net3625),
    .A2(_07870_),
    .Y(_07871_),
    .B1(net3928));
 sg13g2_a22oi_1 _15280_ (.Y(_00811_),
    .B1(_07868_),
    .B2(_07871_),
    .A2(_03425_),
    .A1(net3928));
 sg13g2_nand2b_1 _15281_ (.Y(_07872_),
    .B(_07837_),
    .A_N(net3625));
 sg13g2_a21oi_1 _15282_ (.A1(_04842_),
    .A2(_04852_),
    .Y(_07873_),
    .B1(net3928));
 sg13g2_a22oi_1 _15283_ (.Y(_00812_),
    .B1(_07872_),
    .B2(_07873_),
    .A2(_03424_),
    .A1(net3928));
 sg13g2_mux2_1 _15284_ (.A0(net3787),
    .A1(net3786),
    .S(\spiking_network_top_uut.all_data_out[348] ),
    .X(_07874_));
 sg13g2_nor2b_1 _15285_ (.A(\spiking_network_top_uut.all_data_out[348] ),
    .B_N(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[0] ),
    .Y(_07875_));
 sg13g2_a21oi_1 _15286_ (.A1(\spiking_network_top_uut.all_data_out[348] ),
    .A2(net3788),
    .Y(_07876_),
    .B1(_07875_));
 sg13g2_a21oi_1 _15287_ (.A1(\spiking_network_top_uut.all_data_out[349] ),
    .A2(_07874_),
    .Y(_07877_),
    .B1(\spiking_network_top_uut.all_data_out[350] ));
 sg13g2_o21ai_1 _15288_ (.B1(_07877_),
    .Y(_07878_),
    .A1(\spiking_network_top_uut.all_data_out[349] ),
    .A2(_07876_));
 sg13g2_mux2_1 _15289_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[6] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[7] ),
    .S(\spiking_network_top_uut.all_data_out[348] ),
    .X(_07879_));
 sg13g2_nor2b_1 _15290_ (.A(\spiking_network_top_uut.all_data_out[348] ),
    .B_N(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[4] ),
    .Y(_07880_));
 sg13g2_a21oi_1 _15291_ (.A1(\spiking_network_top_uut.all_data_out[348] ),
    .A2(net3784),
    .Y(_07881_),
    .B1(_07880_));
 sg13g2_o21ai_1 _15292_ (.B1(\spiking_network_top_uut.all_data_out[350] ),
    .Y(_07882_),
    .A1(\spiking_network_top_uut.all_data_out[349] ),
    .A2(_07881_));
 sg13g2_a21oi_1 _15293_ (.A1(\spiking_network_top_uut.all_data_out[349] ),
    .A2(_07879_),
    .Y(_07883_),
    .B1(_07882_));
 sg13g2_nand2_1 _15294_ (.Y(_07884_),
    .A(net4637),
    .B(_07878_));
 sg13g2_nand2_1 _15295_ (.Y(_07885_),
    .A(net3962),
    .B(net99));
 sg13g2_o21ai_1 _15296_ (.B1(_07885_),
    .Y(_00813_),
    .A1(_07883_),
    .A2(_07884_));
 sg13g2_mux2_1 _15297_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_dout ),
    .A1(net99),
    .S(net4639),
    .X(_00814_));
 sg13g2_mux4_1 _15298_ (.S0(\spiking_network_top_uut.all_data_out[344] ),
    .A0(net3840),
    .A1(net3839),
    .A2(net3838),
    .A3(net3837),
    .S1(\spiking_network_top_uut.all_data_out[345] ),
    .X(_07886_));
 sg13g2_mux2_1 _15299_ (.A0(net3835),
    .A1(net3834),
    .S(\spiking_network_top_uut.all_data_out[344] ),
    .X(_07887_));
 sg13g2_nor2b_1 _15300_ (.A(\spiking_network_top_uut.all_data_out[344] ),
    .B_N(net3836),
    .Y(_07888_));
 sg13g2_a21oi_1 _15301_ (.A1(\spiking_network_top_uut.all_data_out[344] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[5] ),
    .Y(_07889_),
    .B1(_07888_));
 sg13g2_o21ai_1 _15302_ (.B1(\spiking_network_top_uut.all_data_out[346] ),
    .Y(_07890_),
    .A1(\spiking_network_top_uut.all_data_out[345] ),
    .A2(_07889_));
 sg13g2_a21oi_1 _15303_ (.A1(\spiking_network_top_uut.all_data_out[345] ),
    .A2(_07887_),
    .Y(_07891_),
    .B1(_07890_));
 sg13g2_o21ai_1 _15304_ (.B1(net4641),
    .Y(_07892_),
    .A1(\spiking_network_top_uut.all_data_out[346] ),
    .A2(_07886_));
 sg13g2_nand2_1 _15305_ (.Y(_07893_),
    .A(net3963),
    .B(net74));
 sg13g2_o21ai_1 _15306_ (.B1(_07893_),
    .Y(_00815_),
    .A1(_07891_),
    .A2(_07892_));
 sg13g2_mux2_1 _15307_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_dout ),
    .A1(net74),
    .S(net4640),
    .X(_00816_));
 sg13g2_mux4_1 _15308_ (.S0(\spiking_network_top_uut.all_data_out[340] ),
    .A0(net3833),
    .A1(net3832),
    .A2(net3831),
    .A3(net3830),
    .S1(\spiking_network_top_uut.all_data_out[341] ),
    .X(_07894_));
 sg13g2_mux2_1 _15309_ (.A0(net3828),
    .A1(net3827),
    .S(\spiking_network_top_uut.all_data_out[340] ),
    .X(_07895_));
 sg13g2_nor2b_1 _15310_ (.A(\spiking_network_top_uut.all_data_out[340] ),
    .B_N(net3829),
    .Y(_07896_));
 sg13g2_a21oi_1 _15311_ (.A1(\spiking_network_top_uut.all_data_out[340] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[5] ),
    .Y(_07897_),
    .B1(_07896_));
 sg13g2_o21ai_1 _15312_ (.B1(\spiking_network_top_uut.all_data_out[342] ),
    .Y(_07898_),
    .A1(\spiking_network_top_uut.all_data_out[341] ),
    .A2(_07897_));
 sg13g2_a21oi_1 _15313_ (.A1(\spiking_network_top_uut.all_data_out[341] ),
    .A2(_07895_),
    .Y(_07899_),
    .B1(_07898_));
 sg13g2_o21ai_1 _15314_ (.B1(net4608),
    .Y(_07900_),
    .A1(\spiking_network_top_uut.all_data_out[342] ),
    .A2(_07894_));
 sg13g2_nand2_1 _15315_ (.Y(_07901_),
    .A(net3966),
    .B(net129));
 sg13g2_o21ai_1 _15316_ (.B1(_07901_),
    .Y(_00817_),
    .A1(_07899_),
    .A2(_07900_));
 sg13g2_mux2_1 _15317_ (.A0(net200),
    .A1(net129),
    .S(net4608),
    .X(_00818_));
 sg13g2_mux4_1 _15318_ (.S0(\spiking_network_top_uut.all_data_out[336] ),
    .A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[0] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[1] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[2] ),
    .A3(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[3] ),
    .S1(\spiking_network_top_uut.all_data_out[337] ),
    .X(_07902_));
 sg13g2_mux2_1 _15319_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[6] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[7] ),
    .S(\spiking_network_top_uut.all_data_out[336] ),
    .X(_07903_));
 sg13g2_nor2b_1 _15320_ (.A(\spiking_network_top_uut.all_data_out[336] ),
    .B_N(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[4] ),
    .Y(_07904_));
 sg13g2_a21oi_1 _15321_ (.A1(\spiking_network_top_uut.all_data_out[336] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[5] ),
    .Y(_07905_),
    .B1(_07904_));
 sg13g2_o21ai_1 _15322_ (.B1(\spiking_network_top_uut.all_data_out[338] ),
    .Y(_07906_),
    .A1(\spiking_network_top_uut.all_data_out[337] ),
    .A2(_07905_));
 sg13g2_a21oi_1 _15323_ (.A1(\spiking_network_top_uut.all_data_out[337] ),
    .A2(_07903_),
    .Y(_07907_),
    .B1(_07906_));
 sg13g2_o21ai_1 _15324_ (.B1(net4615),
    .Y(_07908_),
    .A1(\spiking_network_top_uut.all_data_out[338] ),
    .A2(_07902_));
 sg13g2_nand2_1 _15325_ (.Y(_07909_),
    .A(net3965),
    .B(net118));
 sg13g2_o21ai_1 _15326_ (.B1(_07909_),
    .Y(_00819_),
    .A1(_07907_),
    .A2(_07908_));
 sg13g2_mux2_1 _15327_ (.A0(net424),
    .A1(net118),
    .S(net4615),
    .X(_00820_));
 sg13g2_mux4_1 _15328_ (.S0(\spiking_network_top_uut.all_data_out[332] ),
    .A0(net3819),
    .A1(net3818),
    .A2(net3817),
    .A3(net3816),
    .S1(\spiking_network_top_uut.all_data_out[333] ),
    .X(_07910_));
 sg13g2_mux2_1 _15329_ (.A0(net3814),
    .A1(net3813),
    .S(\spiking_network_top_uut.all_data_out[332] ),
    .X(_07911_));
 sg13g2_nor2b_1 _15330_ (.A(\spiking_network_top_uut.all_data_out[332] ),
    .B_N(net3815),
    .Y(_07912_));
 sg13g2_a21oi_1 _15331_ (.A1(\spiking_network_top_uut.all_data_out[332] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[5] ),
    .Y(_07913_),
    .B1(_07912_));
 sg13g2_o21ai_1 _15332_ (.B1(\spiking_network_top_uut.all_data_out[334] ),
    .Y(_07914_),
    .A1(\spiking_network_top_uut.all_data_out[333] ),
    .A2(_07913_));
 sg13g2_a21oi_1 _15333_ (.A1(\spiking_network_top_uut.all_data_out[333] ),
    .A2(_07911_),
    .Y(_07915_),
    .B1(_07914_));
 sg13g2_o21ai_1 _15334_ (.B1(net4626),
    .Y(_07916_),
    .A1(\spiking_network_top_uut.all_data_out[334] ),
    .A2(_07910_));
 sg13g2_nand2_1 _15335_ (.Y(_07917_),
    .A(net3960),
    .B(net68));
 sg13g2_o21ai_1 _15336_ (.B1(_07917_),
    .Y(_00821_),
    .A1(_07915_),
    .A2(_07916_));
 sg13g2_mux2_1 _15337_ (.A0(net216),
    .A1(net68),
    .S(net4626),
    .X(_00822_));
 sg13g2_mux4_1 _15338_ (.S0(\spiking_network_top_uut.all_data_out[328] ),
    .A0(net3812),
    .A1(net3811),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[2] ),
    .A3(net3809),
    .S1(\spiking_network_top_uut.all_data_out[329] ),
    .X(_07918_));
 sg13g2_mux2_1 _15339_ (.A0(net3806),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[7] ),
    .S(\spiking_network_top_uut.all_data_out[328] ),
    .X(_07919_));
 sg13g2_nor2b_1 _15340_ (.A(\spiking_network_top_uut.all_data_out[328] ),
    .B_N(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[4] ),
    .Y(_07920_));
 sg13g2_a21oi_1 _15341_ (.A1(\spiking_network_top_uut.all_data_out[328] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[5] ),
    .Y(_07921_),
    .B1(_07920_));
 sg13g2_o21ai_1 _15342_ (.B1(\spiking_network_top_uut.all_data_out[330] ),
    .Y(_07922_),
    .A1(\spiking_network_top_uut.all_data_out[329] ),
    .A2(_07921_));
 sg13g2_a21oi_1 _15343_ (.A1(\spiking_network_top_uut.all_data_out[329] ),
    .A2(_07919_),
    .Y(_07923_),
    .B1(_07922_));
 sg13g2_o21ai_1 _15344_ (.B1(net4623),
    .Y(_07924_),
    .A1(\spiking_network_top_uut.all_data_out[330] ),
    .A2(_07918_));
 sg13g2_nand2_1 _15345_ (.Y(_07925_),
    .A(net3960),
    .B(net139));
 sg13g2_o21ai_1 _15346_ (.B1(_07925_),
    .Y(_00823_),
    .A1(_07923_),
    .A2(_07924_));
 sg13g2_mux2_1 _15347_ (.A0(net247),
    .A1(net139),
    .S(net4624),
    .X(_00824_));
 sg13g2_mux4_1 _15348_ (.S0(\spiking_network_top_uut.all_data_out[324] ),
    .A0(net3804),
    .A1(net3803),
    .A2(net3802),
    .A3(net3801),
    .S1(\spiking_network_top_uut.all_data_out[325] ),
    .X(_07926_));
 sg13g2_mux2_1 _15349_ (.A0(net3798),
    .A1(net3797),
    .S(\spiking_network_top_uut.all_data_out[324] ),
    .X(_07927_));
 sg13g2_nor2b_1 _15350_ (.A(\spiking_network_top_uut.all_data_out[324] ),
    .B_N(net3800),
    .Y(_07928_));
 sg13g2_a21oi_1 _15351_ (.A1(\spiking_network_top_uut.all_data_out[324] ),
    .A2(net3799),
    .Y(_07929_),
    .B1(_07928_));
 sg13g2_o21ai_1 _15352_ (.B1(\spiking_network_top_uut.all_data_out[326] ),
    .Y(_07930_),
    .A1(\spiking_network_top_uut.all_data_out[325] ),
    .A2(_07929_));
 sg13g2_a21oi_1 _15353_ (.A1(\spiking_network_top_uut.all_data_out[325] ),
    .A2(_07927_),
    .Y(_07931_),
    .B1(_07930_));
 sg13g2_o21ai_1 _15354_ (.B1(net4631),
    .Y(_07932_),
    .A1(\spiking_network_top_uut.all_data_out[326] ),
    .A2(_07926_));
 sg13g2_nand2_1 _15355_ (.Y(_07933_),
    .A(net3961),
    .B(net288));
 sg13g2_o21ai_1 _15356_ (.B1(_07933_),
    .Y(_00825_),
    .A1(_07931_),
    .A2(_07932_));
 sg13g2_mux2_1 _15357_ (.A0(net374),
    .A1(net288),
    .S(net4633),
    .X(_00826_));
 sg13g2_mux4_1 _15358_ (.S0(\spiking_network_top_uut.all_data_out[320] ),
    .A0(net3796),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[1] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[2] ),
    .A3(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[3] ),
    .S1(\spiking_network_top_uut.all_data_out[321] ),
    .X(_07934_));
 sg13g2_mux2_1 _15359_ (.A0(net3791),
    .A1(net3790),
    .S(\spiking_network_top_uut.all_data_out[320] ),
    .X(_07935_));
 sg13g2_nor2b_1 _15360_ (.A(\spiking_network_top_uut.all_data_out[320] ),
    .B_N(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[4] ),
    .Y(_07936_));
 sg13g2_a21oi_1 _15361_ (.A1(\spiking_network_top_uut.all_data_out[320] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[5] ),
    .Y(_07937_),
    .B1(_07936_));
 sg13g2_o21ai_1 _15362_ (.B1(\spiking_network_top_uut.all_data_out[322] ),
    .Y(_07938_),
    .A1(\spiking_network_top_uut.all_data_out[321] ),
    .A2(_07937_));
 sg13g2_a21oi_1 _15363_ (.A1(\spiking_network_top_uut.all_data_out[321] ),
    .A2(_07935_),
    .Y(_07939_),
    .B1(_07938_));
 sg13g2_o21ai_1 _15364_ (.B1(net4635),
    .Y(_07940_),
    .A1(\spiking_network_top_uut.all_data_out[322] ),
    .A2(_07934_));
 sg13g2_nand2_1 _15365_ (.Y(_07941_),
    .A(net3964),
    .B(net165));
 sg13g2_o21ai_1 _15366_ (.B1(_07941_),
    .Y(_00827_),
    .A1(_07939_),
    .A2(_07940_));
 sg13g2_nor3_2 _15367_ (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[2] ),
    .B(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[1] ),
    .C(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[0] ),
    .Y(_07942_));
 sg13g2_nor2b_2 _15368_ (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[3] ),
    .B_N(_07942_),
    .Y(_07943_));
 sg13g2_nor2b_2 _15369_ (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[4] ),
    .B_N(_07943_),
    .Y(_07944_));
 sg13g2_nand2b_2 _15370_ (.Y(_07945_),
    .B(_07943_),
    .A_N(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[4] ));
 sg13g2_o21ai_1 _15371_ (.B1(net4606),
    .Y(_07946_),
    .A1(net3647),
    .A2(_07945_));
 sg13g2_nor2b_1 _15372_ (.A(net3646),
    .B_N(_00096_),
    .Y(_07947_));
 sg13g2_a21oi_1 _15373_ (.A1(net4285),
    .A2(net3646),
    .Y(_07948_),
    .B1(_07947_));
 sg13g2_nand2_1 _15374_ (.Y(_07949_),
    .A(net357),
    .B(_07946_));
 sg13g2_o21ai_1 _15375_ (.B1(_07949_),
    .Y(_00828_),
    .A1(_07946_),
    .A2(_07948_));
 sg13g2_xor2_1 _15376_ (.B(net357),
    .A(net381),
    .X(_07950_));
 sg13g2_nor2_1 _15377_ (.A(net3646),
    .B(_07950_),
    .Y(_07951_));
 sg13g2_a21oi_1 _15378_ (.A1(net4282),
    .A2(net3646),
    .Y(_07952_),
    .B1(_07951_));
 sg13g2_nand2_1 _15379_ (.Y(_07953_),
    .A(net381),
    .B(_07946_));
 sg13g2_o21ai_1 _15380_ (.B1(_07953_),
    .Y(_00829_),
    .A1(_07946_),
    .A2(_07952_));
 sg13g2_o21ai_1 _15381_ (.B1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[2] ),
    .Y(_07954_),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[1] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[0] ));
 sg13g2_nor2b_1 _15382_ (.A(_07942_),
    .B_N(_07954_),
    .Y(_07955_));
 sg13g2_nor2_1 _15383_ (.A(net3646),
    .B(_07955_),
    .Y(_07956_));
 sg13g2_a21oi_1 _15384_ (.A1(net4278),
    .A2(net3646),
    .Y(_07957_),
    .B1(_07956_));
 sg13g2_nand2_1 _15385_ (.Y(_07958_),
    .A(net173),
    .B(_07946_));
 sg13g2_o21ai_1 _15386_ (.B1(_07958_),
    .Y(_00830_),
    .A1(_07946_),
    .A2(_07957_));
 sg13g2_nand2_1 _15387_ (.Y(_07959_),
    .A(net4275),
    .B(net3647));
 sg13g2_xnor2_1 _15388_ (.Y(_07960_),
    .A(net436),
    .B(_07942_));
 sg13g2_o21ai_1 _15389_ (.B1(_07959_),
    .Y(_07961_),
    .A1(net3647),
    .A2(_07960_));
 sg13g2_mux2_1 _15390_ (.A0(_07961_),
    .A1(net436),
    .S(_07946_),
    .X(_00831_));
 sg13g2_nand2_1 _15391_ (.Y(_07962_),
    .A(net265),
    .B(net3956));
 sg13g2_nand2b_1 _15392_ (.Y(_07963_),
    .B(net265),
    .A_N(_07943_));
 sg13g2_a21oi_1 _15393_ (.A1(_07945_),
    .A2(_07963_),
    .Y(_07964_),
    .B1(net3646));
 sg13g2_a21oi_1 _15394_ (.A1(net4271),
    .A2(net3647),
    .Y(_07965_),
    .B1(_07964_));
 sg13g2_o21ai_1 _15395_ (.B1(_07962_),
    .Y(_00832_),
    .A1(_07946_),
    .A2(_07965_));
 sg13g2_mux2_1 _15396_ (.A0(net469),
    .A1(net165),
    .S(net4634),
    .X(_00833_));
 sg13g2_mux2_1 _15397_ (.A0(net4602),
    .A1(\spiking_network_top_uut.all_data_out[896] ),
    .S(\spiking_network_top_uut.debug_config_ready_sync ),
    .X(_00834_));
 sg13g2_mux2_1 _15398_ (.A0(net4601),
    .A1(\spiking_network_top_uut.all_data_out[897] ),
    .S(\spiking_network_top_uut.debug_config_ready_sync ),
    .X(_00835_));
 sg13g2_mux2_1 _15399_ (.A0(net520),
    .A1(\spiking_network_top_uut.all_data_out[898] ),
    .S(\spiking_network_top_uut.debug_config_ready_sync ),
    .X(_00836_));
 sg13g2_mux2_1 _15400_ (.A0(net515),
    .A1(\spiking_network_top_uut.all_data_out[899] ),
    .S(\spiking_network_top_uut.debug_config_ready_sync ),
    .X(_00837_));
 sg13g2_mux2_1 _15401_ (.A0(net361),
    .A1(\spiking_network_top_uut.all_data_out[900] ),
    .S(\spiking_network_top_uut.debug_config_ready_sync ),
    .X(_00838_));
 sg13g2_mux2_1 _15402_ (.A0(net294),
    .A1(\spiking_network_top_uut.all_data_out[901] ),
    .S(\spiking_network_top_uut.debug_config_ready_sync ),
    .X(_00839_));
 sg13g2_mux2_1 _15403_ (.A0(net362),
    .A1(\spiking_network_top_uut.all_data_out[902] ),
    .S(\spiking_network_top_uut.debug_config_ready_sync ),
    .X(_00840_));
 sg13g2_mux2_1 _15404_ (.A0(net355),
    .A1(\spiking_network_top_uut.all_data_out[903] ),
    .S(\spiking_network_top_uut.debug_config_ready_sync ),
    .X(_00841_));
 sg13g2_a21oi_1 _15405_ (.A1(net3915),
    .A2(net3912),
    .Y(_07966_),
    .B1(_00091_));
 sg13g2_nor2_2 _15406_ (.A(net3753),
    .B(_07966_),
    .Y(_07967_));
 sg13g2_nor2_1 _15407_ (.A(_00091_),
    .B(_07967_),
    .Y(_07968_));
 sg13g2_nand2b_1 _15408_ (.Y(_07969_),
    .B(_07967_),
    .A_N(_00091_));
 sg13g2_o21ai_1 _15409_ (.B1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ),
    .Y(_07970_),
    .A1(_00091_),
    .A2(_07967_));
 sg13g2_a21o_1 _15410_ (.A2(net3753),
    .A1(_00092_),
    .B1(_07967_),
    .X(_07971_));
 sg13g2_nor2_1 _15411_ (.A(_00092_),
    .B(net3908),
    .Y(_07972_));
 sg13g2_a221oi_1 _15412_ (.B2(_07966_),
    .C1(_07972_),
    .B1(net3908),
    .A1(_03492_),
    .Y(_07973_),
    .A2(net3753));
 sg13g2_nand2_1 _15413_ (.Y(_07974_),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ),
    .B(_07973_));
 sg13g2_o21ai_1 _15414_ (.B1(_05086_),
    .Y(_07975_),
    .A1(_00091_),
    .A2(net3912));
 sg13g2_a221oi_1 _15415_ (.B2(_03491_),
    .C1(_07975_),
    .B1(net3902),
    .A1(_03492_),
    .Y(_07976_),
    .A2(net3739));
 sg13g2_and2_1 _15416_ (.A(_00095_),
    .B(net3754),
    .X(_07977_));
 sg13g2_nor3_2 _15417_ (.A(_03493_),
    .B(_07976_),
    .C(_07977_),
    .Y(_07978_));
 sg13g2_xnor2_1 _15418_ (.Y(_07979_),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ),
    .B(_07973_));
 sg13g2_o21ai_1 _15419_ (.B1(_07974_),
    .Y(_07980_),
    .A1(_07978_),
    .A2(_07979_));
 sg13g2_xnor2_1 _15420_ (.Y(_07981_),
    .A(_03492_),
    .B(_07971_));
 sg13g2_nor2b_1 _15421_ (.A(_07981_),
    .B_N(_07980_),
    .Y(_07982_));
 sg13g2_a21o_1 _15422_ (.A2(_07971_),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ),
    .B1(_07982_),
    .X(_07983_));
 sg13g2_xnor2_1 _15423_ (.Y(_07984_),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ),
    .B(_07968_));
 sg13g2_nand2_1 _15424_ (.Y(_07985_),
    .A(_07983_),
    .B(_07984_));
 sg13g2_nand3_1 _15425_ (.B(_07970_),
    .C(_07985_),
    .A(_07969_),
    .Y(_07986_));
 sg13g2_nand2_1 _15426_ (.Y(_07987_),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ),
    .B(_07967_));
 sg13g2_a22oi_1 _15427_ (.Y(_07988_),
    .B1(_07986_),
    .B2(_07987_),
    .A2(_00091_),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ));
 sg13g2_nor2_1 _15428_ (.A(_07944_),
    .B(_07988_),
    .Y(_07989_));
 sg13g2_mux2_2 _15429_ (.A0(net4492),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[323] ),
    .X(_07990_));
 sg13g2_nand2_1 _15430_ (.Y(_07991_),
    .A(\spiking_network_top_uut.all_data_out[33] ),
    .B(_07990_));
 sg13g2_mux2_2 _15431_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.din ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[327] ),
    .X(_07992_));
 sg13g2_nand2_1 _15432_ (.Y(_07993_),
    .A(\spiking_network_top_uut.all_data_out[35] ),
    .B(_07992_));
 sg13g2_nor2_1 _15433_ (.A(_07991_),
    .B(_07993_),
    .Y(_07994_));
 sg13g2_nand4_1 _15434_ (.B(\spiking_network_top_uut.all_data_out[34] ),
    .C(_07990_),
    .A(\spiking_network_top_uut.all_data_out[32] ),
    .Y(_07995_),
    .D(_07992_));
 sg13g2_inv_1 _15435_ (.Y(_07996_),
    .A(_07995_));
 sg13g2_xor2_1 _15436_ (.B(_07993_),
    .A(_07991_),
    .X(_07997_));
 sg13g2_a21oi_2 _15437_ (.B1(_07994_),
    .Y(_07998_),
    .A2(_07997_),
    .A1(_07995_));
 sg13g2_mux2_2 _15438_ (.A0(net4489),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[335] ),
    .X(_07999_));
 sg13g2_nand2_1 _15439_ (.Y(_08000_),
    .A(\spiking_network_top_uut.all_data_out[39] ),
    .B(_07999_));
 sg13g2_mux2_2 _15440_ (.A0(net4490),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[331] ),
    .X(_08001_));
 sg13g2_nand2_1 _15441_ (.Y(_08002_),
    .A(\spiking_network_top_uut.all_data_out[37] ),
    .B(_08001_));
 sg13g2_nor2_1 _15442_ (.A(_08000_),
    .B(_08002_),
    .Y(_08003_));
 sg13g2_nand2_1 _15443_ (.Y(_08004_),
    .A(\spiking_network_top_uut.all_data_out[38] ),
    .B(_07999_));
 sg13g2_nand2_1 _15444_ (.Y(_08005_),
    .A(\spiking_network_top_uut.all_data_out[36] ),
    .B(_08001_));
 sg13g2_or2_2 _15445_ (.X(_08006_),
    .B(_08005_),
    .A(_08004_));
 sg13g2_xor2_1 _15446_ (.B(_08002_),
    .A(_08000_),
    .X(_08007_));
 sg13g2_a21oi_2 _15447_ (.B1(_08003_),
    .Y(_08008_),
    .A2(_08007_),
    .A1(_08006_));
 sg13g2_mux2_2 _15448_ (.A0(net4488),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[339] ),
    .X(_08009_));
 sg13g2_mux2_2 _15449_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.din ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[343] ),
    .X(_08010_));
 sg13g2_a22oi_1 _15450_ (.Y(_08011_),
    .B1(_08010_),
    .B2(\spiking_network_top_uut.all_data_out[43] ),
    .A2(_08009_),
    .A1(\spiking_network_top_uut.all_data_out[41] ));
 sg13g2_and4_1 _15451_ (.A(\spiking_network_top_uut.all_data_out[40] ),
    .B(\spiking_network_top_uut.all_data_out[42] ),
    .C(_08009_),
    .D(_08010_),
    .X(_08012_));
 sg13g2_nand4_1 _15452_ (.B(\spiking_network_top_uut.all_data_out[42] ),
    .C(_08009_),
    .A(\spiking_network_top_uut.all_data_out[40] ),
    .Y(_08013_),
    .D(_08010_));
 sg13g2_and4_1 _15453_ (.A(\spiking_network_top_uut.all_data_out[41] ),
    .B(\spiking_network_top_uut.all_data_out[43] ),
    .C(_08009_),
    .D(_08010_),
    .X(_08014_));
 sg13g2_nand4_1 _15454_ (.B(\spiking_network_top_uut.all_data_out[43] ),
    .C(_08009_),
    .A(\spiking_network_top_uut.all_data_out[41] ),
    .Y(_08015_),
    .D(_08010_));
 sg13g2_nand3b_1 _15455_ (.B(_08012_),
    .C(_08015_),
    .Y(_08016_),
    .A_N(_08011_));
 sg13g2_a21oi_2 _15456_ (.B1(_08011_),
    .Y(_08017_),
    .A2(_08015_),
    .A1(_08012_));
 sg13g2_mux2_1 _15457_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.din ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[351] ),
    .X(_08018_));
 sg13g2_mux2_2 _15458_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.din ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[347] ),
    .X(_08019_));
 sg13g2_and4_1 _15459_ (.A(\spiking_network_top_uut.all_data_out[47] ),
    .B(\spiking_network_top_uut.all_data_out[45] ),
    .C(_08018_),
    .D(_08019_),
    .X(_08020_));
 sg13g2_nand4_1 _15460_ (.B(\spiking_network_top_uut.all_data_out[45] ),
    .C(_08018_),
    .A(\spiking_network_top_uut.all_data_out[47] ),
    .Y(_08021_),
    .D(_08019_));
 sg13g2_and4_1 _15461_ (.A(\spiking_network_top_uut.all_data_out[46] ),
    .B(\spiking_network_top_uut.all_data_out[44] ),
    .C(_08018_),
    .D(_08019_),
    .X(_08022_));
 sg13g2_a22oi_1 _15462_ (.Y(_08023_),
    .B1(_08019_),
    .B2(\spiking_network_top_uut.all_data_out[45] ),
    .A2(_08018_),
    .A1(\spiking_network_top_uut.all_data_out[47] ));
 sg13g2_or3_2 _15463_ (.A(_08020_),
    .B(_08022_),
    .C(_08023_),
    .X(_08024_));
 sg13g2_o21ai_1 _15464_ (.B1(_08021_),
    .Y(_08025_),
    .A1(_08022_),
    .A2(_08023_));
 sg13g2_nand3b_1 _15465_ (.B(_08017_),
    .C(_08025_),
    .Y(_08026_),
    .A_N(_08008_));
 sg13g2_inv_1 _15466_ (.Y(_08027_),
    .A(_08026_));
 sg13g2_or2_2 _15467_ (.X(_08028_),
    .B(_08026_),
    .A(_07998_));
 sg13g2_a21o_1 _15468_ (.A2(_07985_),
    .A1(_07970_),
    .B1(_07969_),
    .X(_08029_));
 sg13g2_nand2_2 _15469_ (.Y(_08030_),
    .A(_07986_),
    .B(_08029_));
 sg13g2_nor2_1 _15470_ (.A(_08017_),
    .B(_08025_),
    .Y(_08031_));
 sg13g2_and2_1 _15471_ (.A(_08008_),
    .B(_08031_),
    .X(_08032_));
 sg13g2_nand2_2 _15472_ (.Y(_08033_),
    .A(_07998_),
    .B(_08032_));
 sg13g2_and2_1 _15473_ (.A(_08028_),
    .B(_08033_),
    .X(_08034_));
 sg13g2_nand2_1 _15474_ (.Y(_08035_),
    .A(_08030_),
    .B(_08034_));
 sg13g2_nand2_1 _15475_ (.Y(_08036_),
    .A(_08028_),
    .B(_08035_));
 sg13g2_xor2_1 _15476_ (.B(_08034_),
    .A(_07988_),
    .X(_08037_));
 sg13g2_nand2_1 _15477_ (.Y(_08038_),
    .A(_08036_),
    .B(_08037_));
 sg13g2_o21ai_1 _15478_ (.B1(_08022_),
    .Y(_08039_),
    .A1(_08020_),
    .A2(_08023_));
 sg13g2_o21ai_1 _15479_ (.B1(_08013_),
    .Y(_08040_),
    .A1(_08011_),
    .A2(_08014_));
 sg13g2_o21ai_1 _15480_ (.B1(_08012_),
    .Y(_08041_),
    .A1(_08011_),
    .A2(_08014_));
 sg13g2_nand3b_1 _15481_ (.B(_08013_),
    .C(_08015_),
    .Y(_08042_),
    .A_N(_08011_));
 sg13g2_a22oi_1 _15482_ (.Y(_08043_),
    .B1(_08041_),
    .B2(_08042_),
    .A2(_08039_),
    .A1(_08024_));
 sg13g2_xor2_1 _15483_ (.B(_08007_),
    .A(_08006_),
    .X(_08044_));
 sg13g2_xnor2_1 _15484_ (.Y(_08045_),
    .A(_08006_),
    .B(_08007_));
 sg13g2_and4_1 _15485_ (.A(_08024_),
    .B(_08039_),
    .C(_08041_),
    .D(_08042_),
    .X(_08046_));
 sg13g2_nand4_1 _15486_ (.B(_08039_),
    .C(_08041_),
    .A(_08024_),
    .Y(_08047_),
    .D(_08042_));
 sg13g2_and4_1 _15487_ (.A(_08016_),
    .B(_08024_),
    .C(_08039_),
    .D(_08040_),
    .X(_08048_));
 sg13g2_a22oi_1 _15488_ (.Y(_08049_),
    .B1(_08040_),
    .B2(_08016_),
    .A2(_08039_),
    .A1(_08024_));
 sg13g2_nor3_2 _15489_ (.A(_08043_),
    .B(_08044_),
    .C(_08046_),
    .Y(_08050_));
 sg13g2_a21oi_2 _15490_ (.B1(_08043_),
    .Y(_08051_),
    .A2(_08047_),
    .A1(_08045_));
 sg13g2_xor2_1 _15491_ (.B(_08025_),
    .A(_08017_),
    .X(_08052_));
 sg13g2_xnor2_1 _15492_ (.Y(_08053_),
    .A(_08008_),
    .B(_08052_));
 sg13g2_nand2b_1 _15493_ (.Y(_08054_),
    .B(_08053_),
    .A_N(_08051_));
 sg13g2_xnor2_1 _15494_ (.Y(_08055_),
    .A(_08051_),
    .B(_08053_));
 sg13g2_nand2b_1 _15495_ (.Y(_08056_),
    .B(_08055_),
    .A_N(_07998_));
 sg13g2_nand2_1 _15496_ (.Y(_08057_),
    .A(_08054_),
    .B(_08056_));
 sg13g2_nor2_1 _15497_ (.A(_08027_),
    .B(_08032_),
    .Y(_08058_));
 sg13g2_xnor2_1 _15498_ (.Y(_08059_),
    .A(_07998_),
    .B(_08058_));
 sg13g2_and2_2 _15499_ (.A(_08057_),
    .B(_08059_),
    .X(_08060_));
 sg13g2_xor2_1 _15500_ (.B(_08059_),
    .A(_08057_),
    .X(_08061_));
 sg13g2_xnor2_1 _15501_ (.Y(_08062_),
    .A(_07983_),
    .B(_07984_));
 sg13g2_inv_1 _15502_ (.Y(_08063_),
    .A(_08062_));
 sg13g2_a21oi_1 _15503_ (.A1(_08061_),
    .A2(_08063_),
    .Y(_08064_),
    .B1(_08060_));
 sg13g2_xnor2_1 _15504_ (.Y(_08065_),
    .A(_08030_),
    .B(_08034_));
 sg13g2_nor2_1 _15505_ (.A(_08064_),
    .B(_08065_),
    .Y(_08066_));
 sg13g2_a22oi_1 _15506_ (.Y(_08067_),
    .B1(_08019_),
    .B2(\spiking_network_top_uut.all_data_out[44] ),
    .A2(_08018_),
    .A1(\spiking_network_top_uut.all_data_out[46] ));
 sg13g2_nor2_1 _15507_ (.A(_08022_),
    .B(_08067_),
    .Y(_08068_));
 sg13g2_a22oi_1 _15508_ (.Y(_08069_),
    .B1(_08010_),
    .B2(\spiking_network_top_uut.all_data_out[42] ),
    .A2(_08009_),
    .A1(\spiking_network_top_uut.all_data_out[40] ));
 sg13g2_nor2_1 _15509_ (.A(_08012_),
    .B(_08069_),
    .Y(_08070_));
 sg13g2_and2_1 _15510_ (.A(_08068_),
    .B(_08070_),
    .X(_08071_));
 sg13g2_xor2_1 _15511_ (.B(_08005_),
    .A(_08004_),
    .X(_08072_));
 sg13g2_xor2_1 _15512_ (.B(_08070_),
    .A(_08068_),
    .X(_08073_));
 sg13g2_a21oi_2 _15513_ (.B1(_08071_),
    .Y(_08074_),
    .A2(_08073_),
    .A1(_08072_));
 sg13g2_nor3_1 _15514_ (.A(_08045_),
    .B(_08048_),
    .C(_08049_),
    .Y(_08075_));
 sg13g2_nor3_1 _15515_ (.A(_08050_),
    .B(_08074_),
    .C(_08075_),
    .Y(_08076_));
 sg13g2_or3_1 _15516_ (.A(_08050_),
    .B(_08074_),
    .C(_08075_),
    .X(_08077_));
 sg13g2_xnor2_1 _15517_ (.Y(_08078_),
    .A(_07995_),
    .B(_07997_));
 sg13g2_o21ai_1 _15518_ (.B1(_08074_),
    .Y(_08079_),
    .A1(_08050_),
    .A2(_08075_));
 sg13g2_nand3_1 _15519_ (.B(_08078_),
    .C(_08079_),
    .A(_08077_),
    .Y(_08080_));
 sg13g2_a21o_2 _15520_ (.A2(_08079_),
    .A1(_08078_),
    .B1(_08076_),
    .X(_08081_));
 sg13g2_xnor2_1 _15521_ (.Y(_08082_),
    .A(_07998_),
    .B(_08055_));
 sg13g2_nand2_1 _15522_ (.Y(_08083_),
    .A(_08081_),
    .B(_08082_));
 sg13g2_xnor2_1 _15523_ (.Y(_08084_),
    .A(_08081_),
    .B(_08082_));
 sg13g2_xor2_1 _15524_ (.B(_07981_),
    .A(_07980_),
    .X(_08085_));
 sg13g2_o21ai_1 _15525_ (.B1(_08083_),
    .Y(_08086_),
    .A1(_08084_),
    .A2(_08085_));
 sg13g2_xnor2_1 _15526_ (.Y(_08087_),
    .A(_08061_),
    .B(_08062_));
 sg13g2_nand2_1 _15527_ (.Y(_08088_),
    .A(_08086_),
    .B(_08087_));
 sg13g2_a22oi_1 _15528_ (.Y(_08089_),
    .B1(_07992_),
    .B2(\spiking_network_top_uut.all_data_out[34] ),
    .A2(_07990_),
    .A1(\spiking_network_top_uut.all_data_out[32] ));
 sg13g2_xnor2_1 _15529_ (.Y(_08090_),
    .A(_08072_),
    .B(_08073_));
 sg13g2_nor3_2 _15530_ (.A(_07996_),
    .B(_08089_),
    .C(_08090_),
    .Y(_08091_));
 sg13g2_a21o_2 _15531_ (.A2(_08079_),
    .A1(_08077_),
    .B1(_08078_),
    .X(_08092_));
 sg13g2_nand3_1 _15532_ (.B(_08091_),
    .C(_08092_),
    .A(_08080_),
    .Y(_08093_));
 sg13g2_a21oi_1 _15533_ (.A1(_08080_),
    .A2(_08092_),
    .Y(_08094_),
    .B1(_08091_));
 sg13g2_a21o_1 _15534_ (.A2(_08092_),
    .A1(_08080_),
    .B1(_08091_),
    .X(_08095_));
 sg13g2_xnor2_1 _15535_ (.Y(_08096_),
    .A(_07978_),
    .B(_07979_));
 sg13g2_inv_1 _15536_ (.Y(_08097_),
    .A(_08096_));
 sg13g2_and3_1 _15537_ (.X(_08098_),
    .A(_08093_),
    .B(_08095_),
    .C(_08097_));
 sg13g2_o21ai_1 _15538_ (.B1(_08093_),
    .Y(_08099_),
    .A1(_08094_),
    .A2(_08096_));
 sg13g2_xor2_1 _15539_ (.B(_08085_),
    .A(_08084_),
    .X(_08100_));
 sg13g2_and2_1 _15540_ (.A(_08099_),
    .B(_08100_),
    .X(_08101_));
 sg13g2_a21oi_1 _15541_ (.A1(_08093_),
    .A2(_08095_),
    .Y(_08102_),
    .B1(_08097_));
 sg13g2_o21ai_1 _15542_ (.B1(_03493_),
    .Y(_08103_),
    .A1(_07976_),
    .A2(_07977_));
 sg13g2_nand2b_1 _15543_ (.Y(_08104_),
    .B(_08103_),
    .A_N(_07978_));
 sg13g2_o21ai_1 _15544_ (.B1(_08090_),
    .Y(_08105_),
    .A1(_07996_),
    .A2(_08089_));
 sg13g2_nor2b_2 _15545_ (.A(_08091_),
    .B_N(_08105_),
    .Y(_08106_));
 sg13g2_nand2_1 _15546_ (.Y(_08107_),
    .A(_08104_),
    .B(_08106_));
 sg13g2_nor3_2 _15547_ (.A(_08098_),
    .B(_08102_),
    .C(_08107_),
    .Y(_08108_));
 sg13g2_or2_1 _15548_ (.X(_08109_),
    .B(_08100_),
    .A(_08099_));
 sg13g2_nand2b_1 _15549_ (.Y(_08110_),
    .B(_08109_),
    .A_N(_08101_));
 sg13g2_a21oi_2 _15550_ (.B1(_08101_),
    .Y(_08111_),
    .A2(_08109_),
    .A1(_08108_));
 sg13g2_xnor2_1 _15551_ (.Y(_08112_),
    .A(_08086_),
    .B(_08087_));
 sg13g2_o21ai_1 _15552_ (.B1(_08088_),
    .Y(_08113_),
    .A1(_08111_),
    .A2(_08112_));
 sg13g2_nand2_1 _15553_ (.Y(_08114_),
    .A(_08064_),
    .B(_08065_));
 sg13g2_nand2b_1 _15554_ (.Y(_08115_),
    .B(_08114_),
    .A_N(_08066_));
 sg13g2_a21oi_1 _15555_ (.A1(_08113_),
    .A2(_08114_),
    .Y(_08116_),
    .B1(_08066_));
 sg13g2_xnor2_1 _15556_ (.Y(_08117_),
    .A(_08036_),
    .B(_08037_));
 sg13g2_o21ai_1 _15557_ (.B1(_08038_),
    .Y(_08118_),
    .A1(_08116_),
    .A2(_08117_));
 sg13g2_mux2_1 _15558_ (.A0(_08033_),
    .A1(_08028_),
    .S(_07988_),
    .X(_08119_));
 sg13g2_xnor2_1 _15559_ (.Y(_08120_),
    .A(_08118_),
    .B(_08119_));
 sg13g2_a21oi_2 _15560_ (.B1(_07989_),
    .Y(_08121_),
    .A2(_08120_),
    .A1(_07944_));
 sg13g2_xnor2_1 _15561_ (.Y(_08122_),
    .A(_08116_),
    .B(_08117_));
 sg13g2_a21oi_1 _15562_ (.A1(_07944_),
    .A2(_08122_),
    .Y(_08123_),
    .B1(_07989_));
 sg13g2_xnor2_1 _15563_ (.Y(_08124_),
    .A(_08113_),
    .B(_08115_));
 sg13g2_mux2_1 _15564_ (.A0(_08030_),
    .A1(_08124_),
    .S(_07944_),
    .X(_08125_));
 sg13g2_nand2_1 _15565_ (.Y(_08126_),
    .A(_08123_),
    .B(_08125_));
 sg13g2_a21oi_1 _15566_ (.A1(_08121_),
    .A2(_08126_),
    .Y(_08127_),
    .B1(net3647));
 sg13g2_nand2_2 _15567_ (.Y(_08128_),
    .A(net4606),
    .B(_08127_));
 sg13g2_nor2_1 _15568_ (.A(_08123_),
    .B(_08125_),
    .Y(_08129_));
 sg13g2_nor2_2 _15569_ (.A(_08121_),
    .B(_08129_),
    .Y(_08130_));
 sg13g2_nand2_1 _15570_ (.Y(_08131_),
    .A(_07944_),
    .B(_08106_));
 sg13g2_xnor2_1 _15571_ (.Y(_08132_),
    .A(_08104_),
    .B(_08131_));
 sg13g2_nor2_1 _15572_ (.A(_08130_),
    .B(_08132_),
    .Y(_08133_));
 sg13g2_xor2_1 _15573_ (.B(net4316),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[0] ),
    .X(_08134_));
 sg13g2_a22oi_1 _15574_ (.Y(_08135_),
    .B1(_00001_),
    .B2(_08134_),
    .A2(net3957),
    .A1(net522));
 sg13g2_o21ai_1 _15575_ (.B1(_08135_),
    .Y(_00842_),
    .A1(_08128_),
    .A2(_08133_));
 sg13g2_o21ai_1 _15576_ (.B1(_08107_),
    .Y(_08136_),
    .A1(_08098_),
    .A2(_08102_));
 sg13g2_nor2_1 _15577_ (.A(_07945_),
    .B(_08108_),
    .Y(_08137_));
 sg13g2_a221oi_1 _15578_ (.B2(_08137_),
    .C1(_08130_),
    .B1(_08136_),
    .A1(_07945_),
    .Y(_08138_),
    .A2(_08097_));
 sg13g2_xor2_1 _15579_ (.B(_04860_),
    .A(_04859_),
    .X(_08139_));
 sg13g2_a22oi_1 _15580_ (.Y(_08140_),
    .B1(_00001_),
    .B2(_08139_),
    .A2(net3957),
    .A1(net550));
 sg13g2_o21ai_1 _15581_ (.B1(_08140_),
    .Y(_00843_),
    .A1(_08128_),
    .A2(_08138_));
 sg13g2_nand2_1 _15582_ (.Y(_08141_),
    .A(_07945_),
    .B(_08085_));
 sg13g2_xnor2_1 _15583_ (.Y(_08142_),
    .A(_08108_),
    .B(_08110_));
 sg13g2_nand2b_1 _15584_ (.Y(_08143_),
    .B(_07944_),
    .A_N(_08142_));
 sg13g2_a21oi_1 _15585_ (.A1(_08141_),
    .A2(_08143_),
    .Y(_08144_),
    .B1(_08130_));
 sg13g2_xnor2_1 _15586_ (.Y(_08145_),
    .A(_04861_),
    .B(_04862_));
 sg13g2_a22oi_1 _15587_ (.Y(_08146_),
    .B1(_00001_),
    .B2(_08145_),
    .A2(net3956),
    .A1(net551));
 sg13g2_o21ai_1 _15588_ (.B1(_08146_),
    .Y(_00844_),
    .A1(_08128_),
    .A2(_08144_));
 sg13g2_nor2_1 _15589_ (.A(_07944_),
    .B(_08063_),
    .Y(_08147_));
 sg13g2_xnor2_1 _15590_ (.Y(_08148_),
    .A(_08111_),
    .B(_08112_));
 sg13g2_a21oi_1 _15591_ (.A1(_07944_),
    .A2(_08148_),
    .Y(_08149_),
    .B1(_08147_));
 sg13g2_o21ai_1 _15592_ (.B1(_08127_),
    .Y(_08150_),
    .A1(_08130_),
    .A2(_08149_));
 sg13g2_or3_1 _15593_ (.A(_04856_),
    .B(_04857_),
    .C(_04863_),
    .X(_08151_));
 sg13g2_and2_1 _15594_ (.A(_04864_),
    .B(_08151_),
    .X(_08152_));
 sg13g2_a21oi_1 _15595_ (.A1(net3646),
    .A2(_08152_),
    .Y(_08153_),
    .B1(net3955));
 sg13g2_a22oi_1 _15596_ (.Y(_00845_),
    .B1(_08150_),
    .B2(_08153_),
    .A2(net3955),
    .A1(_03400_));
 sg13g2_nand2b_1 _15597_ (.Y(_08154_),
    .B(_08121_),
    .A_N(net3647));
 sg13g2_a21oi_1 _15598_ (.A1(_04855_),
    .A2(_04865_),
    .Y(_08155_),
    .B1(net3955));
 sg13g2_a22oi_1 _15599_ (.Y(_00846_),
    .B1(_08154_),
    .B2(_08155_),
    .A2(net3955),
    .A1(_03399_));
 sg13g2_mux4_1 _15600_ (.S0(\spiking_network_top_uut.all_data_out[380] ),
    .A0(net3789),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[1] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[2] ),
    .A3(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[3] ),
    .S1(\spiking_network_top_uut.all_data_out[381] ),
    .X(_08156_));
 sg13g2_mux2_1 _15601_ (.A0(net3783),
    .A1(net3899),
    .S(\spiking_network_top_uut.all_data_out[380] ),
    .X(_08157_));
 sg13g2_nor2b_1 _15602_ (.A(\spiking_network_top_uut.all_data_out[380] ),
    .B_N(net3785),
    .Y(_08158_));
 sg13g2_a21oi_1 _15603_ (.A1(\spiking_network_top_uut.all_data_out[380] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[5] ),
    .Y(_08159_),
    .B1(_08158_));
 sg13g2_o21ai_1 _15604_ (.B1(\spiking_network_top_uut.all_data_out[382] ),
    .Y(_08160_),
    .A1(\spiking_network_top_uut.all_data_out[381] ),
    .A2(_08159_));
 sg13g2_a21oi_1 _15605_ (.A1(\spiking_network_top_uut.all_data_out[381] ),
    .A2(_08157_),
    .Y(_08161_),
    .B1(_08160_));
 sg13g2_o21ai_1 _15606_ (.B1(net4637),
    .Y(_08162_),
    .A1(\spiking_network_top_uut.all_data_out[382] ),
    .A2(_08156_));
 sg13g2_nand2_1 _15607_ (.Y(_08163_),
    .A(net3962),
    .B(net249));
 sg13g2_o21ai_1 _15608_ (.B1(_08163_),
    .Y(_00847_),
    .A1(_08161_),
    .A2(_08162_));
 sg13g2_mux2_1 _15609_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_dout ),
    .A1(net249),
    .S(net4642),
    .X(_00848_));
 sg13g2_mux4_1 _15610_ (.S0(\spiking_network_top_uut.all_data_out[376] ),
    .A0(net3840),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[1] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[2] ),
    .A3(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[3] ),
    .S1(\spiking_network_top_uut.all_data_out[377] ),
    .X(_08164_));
 sg13g2_mux2_1 _15611_ (.A0(net3835),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[7] ),
    .S(\spiking_network_top_uut.all_data_out[376] ),
    .X(_08165_));
 sg13g2_nor2b_1 _15612_ (.A(\spiking_network_top_uut.all_data_out[376] ),
    .B_N(net3836),
    .Y(_08166_));
 sg13g2_a21oi_1 _15613_ (.A1(\spiking_network_top_uut.all_data_out[376] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[5] ),
    .Y(_08167_),
    .B1(_08166_));
 sg13g2_o21ai_1 _15614_ (.B1(\spiking_network_top_uut.all_data_out[378] ),
    .Y(_08168_),
    .A1(\spiking_network_top_uut.all_data_out[377] ),
    .A2(_08167_));
 sg13g2_a21oi_1 _15615_ (.A1(\spiking_network_top_uut.all_data_out[377] ),
    .A2(_08165_),
    .Y(_08169_),
    .B1(_08168_));
 sg13g2_o21ai_1 _15616_ (.B1(net4640),
    .Y(_08170_),
    .A1(\spiking_network_top_uut.all_data_out[378] ),
    .A2(_08164_));
 sg13g2_nand2_1 _15617_ (.Y(_08171_),
    .A(net3963),
    .B(net189));
 sg13g2_o21ai_1 _15618_ (.B1(_08171_),
    .Y(_00849_),
    .A1(_08169_),
    .A2(_08170_));
 sg13g2_mux2_1 _15619_ (.A0(net328),
    .A1(net189),
    .S(net4636),
    .X(_00850_));
 sg13g2_nand2_1 _15620_ (.Y(_08172_),
    .A(\spiking_network_top_uut.all_data_out[372] ),
    .B(_03661_));
 sg13g2_nor2_1 _15621_ (.A(\spiking_network_top_uut.all_data_out[372] ),
    .B(net3829),
    .Y(_08173_));
 sg13g2_nor2_1 _15622_ (.A(\spiking_network_top_uut.all_data_out[373] ),
    .B(_08173_),
    .Y(_08174_));
 sg13g2_mux2_1 _15623_ (.A0(net3828),
    .A1(net3827),
    .S(\spiking_network_top_uut.all_data_out[372] ),
    .X(_08175_));
 sg13g2_a221oi_1 _15624_ (.B2(\spiking_network_top_uut.all_data_out[373] ),
    .C1(_03545_),
    .B1(_08175_),
    .A1(_08172_),
    .Y(_08176_),
    .A2(_08174_));
 sg13g2_mux4_1 _15625_ (.S0(\spiking_network_top_uut.all_data_out[372] ),
    .A0(net3833),
    .A1(net3832),
    .A2(net3831),
    .A3(net3830),
    .S1(\spiking_network_top_uut.all_data_out[373] ),
    .X(_08177_));
 sg13g2_o21ai_1 _15626_ (.B1(net4609),
    .Y(_08178_),
    .A1(\spiking_network_top_uut.all_data_out[374] ),
    .A2(_08177_));
 sg13g2_nand2_1 _15627_ (.Y(_08179_),
    .A(net3966),
    .B(net193));
 sg13g2_o21ai_1 _15628_ (.B1(_08179_),
    .Y(_00851_),
    .A1(_08176_),
    .A2(_08178_));
 sg13g2_mux2_1 _15629_ (.A0(net125),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_reg1 ),
    .S(net4609),
    .X(_00852_));
 sg13g2_mux2_1 _15630_ (.A0(net3824),
    .A1(net3823),
    .S(\spiking_network_top_uut.all_data_out[368] ),
    .X(_08180_));
 sg13g2_nor2b_1 _15631_ (.A(\spiking_network_top_uut.all_data_out[368] ),
    .B_N(net3826),
    .Y(_08181_));
 sg13g2_a21oi_1 _15632_ (.A1(\spiking_network_top_uut.all_data_out[368] ),
    .A2(net3825),
    .Y(_08182_),
    .B1(_08181_));
 sg13g2_a21oi_1 _15633_ (.A1(\spiking_network_top_uut.all_data_out[369] ),
    .A2(_08180_),
    .Y(_08183_),
    .B1(\spiking_network_top_uut.all_data_out[370] ));
 sg13g2_o21ai_1 _15634_ (.B1(_08183_),
    .Y(_08184_),
    .A1(\spiking_network_top_uut.all_data_out[369] ),
    .A2(_08182_));
 sg13g2_mux2_1 _15635_ (.A0(net3821),
    .A1(net3820),
    .S(\spiking_network_top_uut.all_data_out[368] ),
    .X(_08185_));
 sg13g2_nand2_1 _15636_ (.Y(_08186_),
    .A(\spiking_network_top_uut.all_data_out[369] ),
    .B(_08185_));
 sg13g2_a21oi_1 _15637_ (.A1(\spiking_network_top_uut.all_data_out[368] ),
    .A2(_03660_),
    .Y(_08187_),
    .B1(\spiking_network_top_uut.all_data_out[369] ));
 sg13g2_o21ai_1 _15638_ (.B1(_08187_),
    .Y(_08188_),
    .A1(\spiking_network_top_uut.all_data_out[368] ),
    .A2(net3822));
 sg13g2_nand3_1 _15639_ (.B(_08186_),
    .C(_08188_),
    .A(\spiking_network_top_uut.all_data_out[370] ),
    .Y(_08189_));
 sg13g2_nand3_1 _15640_ (.B(_08184_),
    .C(_08189_),
    .A(net4613),
    .Y(_08190_));
 sg13g2_o21ai_1 _15641_ (.B1(_08190_),
    .Y(_00853_),
    .A1(net4614),
    .A2(_03683_));
 sg13g2_mux2_1 _15642_ (.A0(net177),
    .A1(net136),
    .S(net4614),
    .X(_00854_));
 sg13g2_a21oi_1 _15643_ (.A1(\spiking_network_top_uut.all_data_out[364] ),
    .A2(_03659_),
    .Y(_08191_),
    .B1(\spiking_network_top_uut.all_data_out[365] ));
 sg13g2_o21ai_1 _15644_ (.B1(_08191_),
    .Y(_08192_),
    .A1(\spiking_network_top_uut.all_data_out[364] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[4] ));
 sg13g2_mux2_1 _15645_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[6] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[7] ),
    .S(\spiking_network_top_uut.all_data_out[364] ),
    .X(_08193_));
 sg13g2_nand2_1 _15646_ (.Y(_08194_),
    .A(\spiking_network_top_uut.all_data_out[365] ),
    .B(_08193_));
 sg13g2_nand3_1 _15647_ (.B(_08192_),
    .C(_08194_),
    .A(\spiking_network_top_uut.all_data_out[366] ),
    .Y(_08195_));
 sg13g2_mux2_1 _15648_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[2] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[3] ),
    .S(\spiking_network_top_uut.all_data_out[364] ),
    .X(_08196_));
 sg13g2_nor2b_1 _15649_ (.A(\spiking_network_top_uut.all_data_out[364] ),
    .B_N(net3819),
    .Y(_08197_));
 sg13g2_a21oi_1 _15650_ (.A1(\spiking_network_top_uut.all_data_out[364] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[1] ),
    .Y(_08198_),
    .B1(_08197_));
 sg13g2_a21oi_1 _15651_ (.A1(\spiking_network_top_uut.all_data_out[365] ),
    .A2(_08196_),
    .Y(_08199_),
    .B1(\spiking_network_top_uut.all_data_out[366] ));
 sg13g2_o21ai_1 _15652_ (.B1(_08199_),
    .Y(_08200_),
    .A1(\spiking_network_top_uut.all_data_out[365] ),
    .A2(_08198_));
 sg13g2_nand3_1 _15653_ (.B(_08195_),
    .C(_08200_),
    .A(net4627),
    .Y(_08201_));
 sg13g2_o21ai_1 _15654_ (.B1(_08201_),
    .Y(_00855_),
    .A1(net4627),
    .A2(_03684_));
 sg13g2_nor2_1 _15655_ (.A(net4628),
    .B(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_dout ),
    .Y(_08202_));
 sg13g2_a21oi_1 _15656_ (.A1(net4628),
    .A2(_03684_),
    .Y(_00856_),
    .B1(_08202_));
 sg13g2_mux4_1 _15657_ (.S0(\spiking_network_top_uut.all_data_out[360] ),
    .A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[0] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[1] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[2] ),
    .A3(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[3] ),
    .S1(\spiking_network_top_uut.all_data_out[361] ),
    .X(_08203_));
 sg13g2_mux2_1 _15658_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[6] ),
    .A1(net3805),
    .S(\spiking_network_top_uut.all_data_out[360] ),
    .X(_08204_));
 sg13g2_nor2b_1 _15659_ (.A(\spiking_network_top_uut.all_data_out[360] ),
    .B_N(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[4] ),
    .Y(_08205_));
 sg13g2_a21oi_1 _15660_ (.A1(\spiking_network_top_uut.all_data_out[360] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[5] ),
    .Y(_08206_),
    .B1(_08205_));
 sg13g2_o21ai_1 _15661_ (.B1(\spiking_network_top_uut.all_data_out[362] ),
    .Y(_08207_),
    .A1(\spiking_network_top_uut.all_data_out[361] ),
    .A2(_08206_));
 sg13g2_a21oi_1 _15662_ (.A1(\spiking_network_top_uut.all_data_out[361] ),
    .A2(_08204_),
    .Y(_08208_),
    .B1(_08207_));
 sg13g2_o21ai_1 _15663_ (.B1(net4630),
    .Y(_08209_),
    .A1(\spiking_network_top_uut.all_data_out[362] ),
    .A2(_08203_));
 sg13g2_nand2_1 _15664_ (.Y(_08210_),
    .A(net3959),
    .B(net73));
 sg13g2_o21ai_1 _15665_ (.B1(_08210_),
    .Y(_00857_),
    .A1(_08208_),
    .A2(_08209_));
 sg13g2_mux2_1 _15666_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_dout ),
    .A1(net73),
    .S(net4630),
    .X(_00858_));
 sg13g2_mux4_1 _15667_ (.S0(\spiking_network_top_uut.all_data_out[356] ),
    .A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[0] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[1] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[2] ),
    .A3(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[3] ),
    .S1(\spiking_network_top_uut.all_data_out[357] ),
    .X(_08211_));
 sg13g2_mux2_1 _15668_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[6] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[7] ),
    .S(\spiking_network_top_uut.all_data_out[356] ),
    .X(_08212_));
 sg13g2_nor2b_1 _15669_ (.A(\spiking_network_top_uut.all_data_out[356] ),
    .B_N(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[4] ),
    .Y(_08213_));
 sg13g2_a21oi_1 _15670_ (.A1(\spiking_network_top_uut.all_data_out[356] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[5] ),
    .Y(_08214_),
    .B1(_08213_));
 sg13g2_o21ai_1 _15671_ (.B1(\spiking_network_top_uut.all_data_out[358] ),
    .Y(_08215_),
    .A1(\spiking_network_top_uut.all_data_out[357] ),
    .A2(_08214_));
 sg13g2_a21oi_1 _15672_ (.A1(\spiking_network_top_uut.all_data_out[357] ),
    .A2(_08212_),
    .Y(_08216_),
    .B1(_08215_));
 sg13g2_o21ai_1 _15673_ (.B1(net4633),
    .Y(_08217_),
    .A1(\spiking_network_top_uut.all_data_out[358] ),
    .A2(_08211_));
 sg13g2_nand2_1 _15674_ (.Y(_08218_),
    .A(net3961),
    .B(net43));
 sg13g2_o21ai_1 _15675_ (.B1(_08218_),
    .Y(_00859_),
    .A1(_08216_),
    .A2(_08217_));
 sg13g2_mux2_1 _15676_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_dout ),
    .A1(net43),
    .S(net4636),
    .X(_00860_));
 sg13g2_mux4_1 _15677_ (.S0(\spiking_network_top_uut.all_data_out[352] ),
    .A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[0] ),
    .A1(net3795),
    .A2(net3794),
    .A3(net3793),
    .S1(\spiking_network_top_uut.all_data_out[353] ),
    .X(_08219_));
 sg13g2_mux2_1 _15678_ (.A0(net3791),
    .A1(net3790),
    .S(\spiking_network_top_uut.all_data_out[352] ),
    .X(_08220_));
 sg13g2_nor2b_1 _15679_ (.A(\spiking_network_top_uut.all_data_out[352] ),
    .B_N(net3792),
    .Y(_08221_));
 sg13g2_a21oi_1 _15680_ (.A1(\spiking_network_top_uut.all_data_out[352] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[5] ),
    .Y(_08222_),
    .B1(_08221_));
 sg13g2_o21ai_1 _15681_ (.B1(\spiking_network_top_uut.all_data_out[354] ),
    .Y(_08223_),
    .A1(\spiking_network_top_uut.all_data_out[353] ),
    .A2(_08222_));
 sg13g2_a21oi_1 _15682_ (.A1(\spiking_network_top_uut.all_data_out[353] ),
    .A2(_08220_),
    .Y(_08224_),
    .B1(_08223_));
 sg13g2_o21ai_1 _15683_ (.B1(net4618),
    .Y(_08225_),
    .A1(\spiking_network_top_uut.all_data_out[354] ),
    .A2(_08219_));
 sg13g2_nand2_1 _15684_ (.Y(_08226_),
    .A(net3961),
    .B(net385));
 sg13g2_o21ai_1 _15685_ (.B1(_08226_),
    .Y(_00861_),
    .A1(_08224_),
    .A2(_08225_));
 sg13g2_nor3_2 _15686_ (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[2] ),
    .B(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[1] ),
    .C(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[0] ),
    .Y(_08227_));
 sg13g2_nor2b_2 _15687_ (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[3] ),
    .B_N(_08227_),
    .Y(_08228_));
 sg13g2_nor2b_2 _15688_ (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[4] ),
    .B_N(_08228_),
    .Y(_08229_));
 sg13g2_nand2b_2 _15689_ (.Y(_08230_),
    .B(_08228_),
    .A_N(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[4] ));
 sg13g2_o21ai_1 _15690_ (.B1(net4604),
    .Y(_08231_),
    .A1(net3663),
    .A2(net3702));
 sg13g2_nor2b_1 _15691_ (.A(net3662),
    .B_N(net379),
    .Y(_08232_));
 sg13g2_a21oi_1 _15692_ (.A1(net4284),
    .A2(net3662),
    .Y(_08233_),
    .B1(_08232_));
 sg13g2_nand2_1 _15693_ (.Y(_08234_),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[0] ),
    .B(_08231_));
 sg13g2_o21ai_1 _15694_ (.B1(_08234_),
    .Y(_00862_),
    .A1(_08231_),
    .A2(_08233_));
 sg13g2_xor2_1 _15695_ (.B(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[0] ),
    .A(net402),
    .X(_08235_));
 sg13g2_nor2_1 _15696_ (.A(net3662),
    .B(_08235_),
    .Y(_08236_));
 sg13g2_a21oi_1 _15697_ (.A1(net4281),
    .A2(net3662),
    .Y(_08237_),
    .B1(_08236_));
 sg13g2_nand2_1 _15698_ (.Y(_08238_),
    .A(net402),
    .B(_08231_));
 sg13g2_o21ai_1 _15699_ (.B1(_08238_),
    .Y(_00863_),
    .A1(_08231_),
    .A2(_08237_));
 sg13g2_o21ai_1 _15700_ (.B1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[2] ),
    .Y(_08239_),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[1] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[0] ));
 sg13g2_nor2b_1 _15701_ (.A(_08227_),
    .B_N(_08239_),
    .Y(_08240_));
 sg13g2_nor2_1 _15702_ (.A(net3662),
    .B(_08240_),
    .Y(_08241_));
 sg13g2_a21oi_1 _15703_ (.A1(net4277),
    .A2(net3662),
    .Y(_08242_),
    .B1(_08241_));
 sg13g2_nand2_1 _15704_ (.Y(_08243_),
    .A(net235),
    .B(_08231_));
 sg13g2_o21ai_1 _15705_ (.B1(_08243_),
    .Y(_00864_),
    .A1(_08231_),
    .A2(_08242_));
 sg13g2_nand2_1 _15706_ (.Y(_08244_),
    .A(net4274),
    .B(net3663));
 sg13g2_xnor2_1 _15707_ (.Y(_08245_),
    .A(net416),
    .B(_08227_));
 sg13g2_o21ai_1 _15708_ (.B1(_08244_),
    .Y(_08246_),
    .A1(net3662),
    .A2(_08245_));
 sg13g2_mux2_1 _15709_ (.A0(_08246_),
    .A1(net416),
    .S(_08231_),
    .X(_00865_));
 sg13g2_nand2_1 _15710_ (.Y(_08247_),
    .A(net3949),
    .B(net403));
 sg13g2_nand2b_1 _15711_ (.Y(_08248_),
    .B(net403),
    .A_N(_08228_));
 sg13g2_a21oi_1 _15712_ (.A1(net3702),
    .A2(_08248_),
    .Y(_08249_),
    .B1(net3663));
 sg13g2_a21oi_1 _15713_ (.A1(net4270),
    .A2(net3662),
    .Y(_08250_),
    .B1(_08249_));
 sg13g2_o21ai_1 _15714_ (.B1(_08247_),
    .Y(_00866_),
    .A1(_08231_),
    .A2(_08250_));
 sg13g2_mux2_1 _15715_ (.A0(net446),
    .A1(net385),
    .S(net4634),
    .X(_00867_));
 sg13g2_nor2_1 _15716_ (.A(_00097_),
    .B(net3741),
    .Y(_08251_));
 sg13g2_nor3_2 _15717_ (.A(_00097_),
    .B(net3749),
    .C(_05090_),
    .Y(_08252_));
 sg13g2_nand2_1 _15718_ (.Y(_08253_),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ),
    .B(_00097_));
 sg13g2_a21oi_1 _15719_ (.A1(net3918),
    .A2(net3740),
    .Y(_08254_),
    .B1(_00097_));
 sg13g2_nor2_1 _15720_ (.A(_03403_),
    .B(_08254_),
    .Y(_08255_));
 sg13g2_nand2_1 _15721_ (.Y(_08256_),
    .A(_00098_),
    .B(net3751));
 sg13g2_o21ai_1 _15722_ (.B1(_08256_),
    .Y(_08257_),
    .A1(net3751),
    .A2(_08251_));
 sg13g2_nor2_1 _15723_ (.A(_00098_),
    .B(net3907),
    .Y(_08258_));
 sg13g2_a221oi_1 _15724_ (.B2(_08251_),
    .C1(_08258_),
    .B1(net3907),
    .A1(_03495_),
    .Y(_08259_),
    .A2(net3751));
 sg13g2_nand2_1 _15725_ (.Y(_08260_),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ),
    .B(_08259_));
 sg13g2_o21ai_1 _15726_ (.B1(net3918),
    .Y(_08261_),
    .A1(_00097_),
    .A2(net3911));
 sg13g2_a221oi_1 _15727_ (.B2(_03494_),
    .C1(_08261_),
    .B1(net3902),
    .A1(_03495_),
    .Y(_08262_),
    .A2(net3739));
 sg13g2_a21oi_1 _15728_ (.A1(_00101_),
    .A2(net3752),
    .Y(_08263_),
    .B1(_08262_));
 sg13g2_and2_1 _15729_ (.A(_00100_),
    .B(_08263_),
    .X(_08264_));
 sg13g2_xnor2_1 _15730_ (.Y(_08265_),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ),
    .B(_08259_));
 sg13g2_o21ai_1 _15731_ (.B1(_08260_),
    .Y(_08266_),
    .A1(_08264_),
    .A2(_08265_));
 sg13g2_xnor2_1 _15732_ (.Y(_08267_),
    .A(_03495_),
    .B(_08257_));
 sg13g2_nor2b_1 _15733_ (.A(_08267_),
    .B_N(_08266_),
    .Y(_08268_));
 sg13g2_a21o_1 _15734_ (.A2(_08257_),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ),
    .B1(_08268_),
    .X(_08269_));
 sg13g2_xnor2_1 _15735_ (.Y(_08270_),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ),
    .B(_08254_));
 sg13g2_a21oi_1 _15736_ (.A1(_08269_),
    .A2(_08270_),
    .Y(_08271_),
    .B1(_08255_));
 sg13g2_nor2b_1 _15737_ (.A(_08252_),
    .B_N(_08271_),
    .Y(_08272_));
 sg13g2_a22oi_1 _15738_ (.Y(_08273_),
    .B1(_08253_),
    .B2(_08272_),
    .A2(_08252_),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ));
 sg13g2_and2_1 _15739_ (.A(_08230_),
    .B(_08273_),
    .X(_08274_));
 sg13g2_inv_1 _15740_ (.Y(_08275_),
    .A(_08274_));
 sg13g2_mux2_2 _15741_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.din ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[359] ),
    .X(_08276_));
 sg13g2_nand2_2 _15742_ (.Y(_08277_),
    .A(\spiking_network_top_uut.all_data_out[51] ),
    .B(_08276_));
 sg13g2_mux2_2 _15743_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.din ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[355] ),
    .X(_08278_));
 sg13g2_nand2_1 _15744_ (.Y(_08279_),
    .A(\spiking_network_top_uut.all_data_out[49] ),
    .B(_08278_));
 sg13g2_nor2_1 _15745_ (.A(_08277_),
    .B(_08279_),
    .Y(_08280_));
 sg13g2_nand2_2 _15746_ (.Y(_08281_),
    .A(\spiking_network_top_uut.all_data_out[50] ),
    .B(_08276_));
 sg13g2_nand2_1 _15747_ (.Y(_08282_),
    .A(\spiking_network_top_uut.all_data_out[48] ),
    .B(_08278_));
 sg13g2_or2_1 _15748_ (.X(_08283_),
    .B(_08282_),
    .A(_08281_));
 sg13g2_xor2_1 _15749_ (.B(_08279_),
    .A(_08277_),
    .X(_08284_));
 sg13g2_a21oi_2 _15750_ (.B1(_08280_),
    .Y(_08285_),
    .A2(_08284_),
    .A1(_08283_));
 sg13g2_mux2_2 _15751_ (.A0(net4489),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[367] ),
    .X(_08286_));
 sg13g2_nand2_1 _15752_ (.Y(_08287_),
    .A(\spiking_network_top_uut.all_data_out[55] ),
    .B(_08286_));
 sg13g2_mux2_2 _15753_ (.A0(net4490),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[363] ),
    .X(_08288_));
 sg13g2_nand2_1 _15754_ (.Y(_08289_),
    .A(\spiking_network_top_uut.all_data_out[53] ),
    .B(_08288_));
 sg13g2_nor2_1 _15755_ (.A(_08287_),
    .B(_08289_),
    .Y(_08290_));
 sg13g2_nand2_1 _15756_ (.Y(_08291_),
    .A(\spiking_network_top_uut.all_data_out[54] ),
    .B(_08286_));
 sg13g2_nand2_1 _15757_ (.Y(_08292_),
    .A(\spiking_network_top_uut.all_data_out[52] ),
    .B(_08288_));
 sg13g2_or2_1 _15758_ (.X(_08293_),
    .B(_08292_),
    .A(_08291_));
 sg13g2_xor2_1 _15759_ (.B(_08289_),
    .A(_08287_),
    .X(_08294_));
 sg13g2_a21oi_2 _15760_ (.B1(_08290_),
    .Y(_08295_),
    .A2(_08294_),
    .A1(_08293_));
 sg13g2_mux2_2 _15761_ (.A0(net4487),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[375] ),
    .X(_08296_));
 sg13g2_mux2_2 _15762_ (.A0(net4488),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[371] ),
    .X(_08297_));
 sg13g2_a22oi_1 _15763_ (.Y(_08298_),
    .B1(_08297_),
    .B2(\spiking_network_top_uut.all_data_out[57] ),
    .A2(_08296_),
    .A1(\spiking_network_top_uut.all_data_out[59] ));
 sg13g2_and4_1 _15764_ (.A(\spiking_network_top_uut.all_data_out[59] ),
    .B(\spiking_network_top_uut.all_data_out[57] ),
    .C(_08296_),
    .D(_08297_),
    .X(_08299_));
 sg13g2_nand4_1 _15765_ (.B(\spiking_network_top_uut.all_data_out[57] ),
    .C(_08296_),
    .A(\spiking_network_top_uut.all_data_out[59] ),
    .Y(_08300_),
    .D(_08297_));
 sg13g2_and4_2 _15766_ (.A(\spiking_network_top_uut.all_data_out[58] ),
    .B(\spiking_network_top_uut.all_data_out[56] ),
    .C(_08296_),
    .D(_08297_),
    .X(_08301_));
 sg13g2_a21oi_2 _15767_ (.B1(_08298_),
    .Y(_08302_),
    .A2(_08301_),
    .A1(_08300_));
 sg13g2_mux2_2 _15768_ (.A0(net4486),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[379] ),
    .X(_08303_));
 sg13g2_mux2_2 _15769_ (.A0(net4485),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[383] ),
    .X(_08304_));
 sg13g2_and4_1 _15770_ (.A(\spiking_network_top_uut.all_data_out[61] ),
    .B(\spiking_network_top_uut.all_data_out[63] ),
    .C(_08303_),
    .D(_08304_),
    .X(_08305_));
 sg13g2_nand4_1 _15771_ (.B(\spiking_network_top_uut.all_data_out[63] ),
    .C(_08303_),
    .A(\spiking_network_top_uut.all_data_out[61] ),
    .Y(_08306_),
    .D(_08304_));
 sg13g2_and4_1 _15772_ (.A(\spiking_network_top_uut.all_data_out[60] ),
    .B(\spiking_network_top_uut.all_data_out[62] ),
    .C(_08303_),
    .D(_08304_),
    .X(_08307_));
 sg13g2_a22oi_1 _15773_ (.Y(_08308_),
    .B1(_08304_),
    .B2(\spiking_network_top_uut.all_data_out[63] ),
    .A2(_08303_),
    .A1(\spiking_network_top_uut.all_data_out[61] ));
 sg13g2_or3_1 _15774_ (.A(_08305_),
    .B(_08307_),
    .C(_08308_),
    .X(_08309_));
 sg13g2_o21ai_1 _15775_ (.B1(_08306_),
    .Y(_08310_),
    .A1(_08307_),
    .A2(_08308_));
 sg13g2_nand3b_1 _15776_ (.B(_08302_),
    .C(_08310_),
    .Y(_08311_),
    .A_N(_08295_));
 sg13g2_inv_1 _15777_ (.Y(_08312_),
    .A(_08311_));
 sg13g2_or2_1 _15778_ (.X(_08313_),
    .B(_08311_),
    .A(_08285_));
 sg13g2_inv_1 _15779_ (.Y(_08314_),
    .A(_08313_));
 sg13g2_nor2_1 _15780_ (.A(_08302_),
    .B(_08310_),
    .Y(_08315_));
 sg13g2_and2_1 _15781_ (.A(_08295_),
    .B(_08315_),
    .X(_08316_));
 sg13g2_a21oi_2 _15782_ (.B1(_08314_),
    .Y(_08317_),
    .A2(_08316_),
    .A1(_08285_));
 sg13g2_xor2_1 _15783_ (.B(_08271_),
    .A(_08252_),
    .X(_08318_));
 sg13g2_a21o_1 _15784_ (.A2(_08318_),
    .A1(_08317_),
    .B1(_08314_),
    .X(_08319_));
 sg13g2_nand2b_1 _15785_ (.Y(_08320_),
    .B(_08273_),
    .A_N(_08317_));
 sg13g2_xor2_1 _15786_ (.B(_08317_),
    .A(_08273_),
    .X(_08321_));
 sg13g2_nor2b_1 _15787_ (.A(_08321_),
    .B_N(_08319_),
    .Y(_08322_));
 sg13g2_xnor2_1 _15788_ (.Y(_08323_),
    .A(_08319_),
    .B(_08321_));
 sg13g2_o21ai_1 _15789_ (.B1(_08307_),
    .Y(_08324_),
    .A1(_08305_),
    .A2(_08308_));
 sg13g2_o21ai_1 _15790_ (.B1(_08301_),
    .Y(_08325_),
    .A1(_08298_),
    .A2(_08299_));
 sg13g2_or3_1 _15791_ (.A(_08298_),
    .B(_08299_),
    .C(_08301_),
    .X(_08326_));
 sg13g2_a22oi_1 _15792_ (.Y(_08327_),
    .B1(_08325_),
    .B2(_08326_),
    .A2(_08324_),
    .A1(_08309_));
 sg13g2_xor2_1 _15793_ (.B(_08294_),
    .A(_08293_),
    .X(_08328_));
 sg13g2_xnor2_1 _15794_ (.Y(_08329_),
    .A(_08293_),
    .B(_08294_));
 sg13g2_and4_1 _15795_ (.A(_08309_),
    .B(_08324_),
    .C(_08325_),
    .D(_08326_),
    .X(_08330_));
 sg13g2_nand4_1 _15796_ (.B(_08324_),
    .C(_08325_),
    .A(_08309_),
    .Y(_08331_),
    .D(_08326_));
 sg13g2_nand3b_1 _15797_ (.B(_08329_),
    .C(_08331_),
    .Y(_08332_),
    .A_N(_08327_));
 sg13g2_a21oi_2 _15798_ (.B1(_08327_),
    .Y(_08333_),
    .A2(_08331_),
    .A1(_08329_));
 sg13g2_xor2_1 _15799_ (.B(_08310_),
    .A(_08302_),
    .X(_08334_));
 sg13g2_xnor2_1 _15800_ (.Y(_08335_),
    .A(_08295_),
    .B(_08334_));
 sg13g2_nor2b_1 _15801_ (.A(_08333_),
    .B_N(_08335_),
    .Y(_08336_));
 sg13g2_xnor2_1 _15802_ (.Y(_08337_),
    .A(_08333_),
    .B(_08335_));
 sg13g2_nor2b_1 _15803_ (.A(_08285_),
    .B_N(_08337_),
    .Y(_08338_));
 sg13g2_nor2_1 _15804_ (.A(_08336_),
    .B(_08338_),
    .Y(_08339_));
 sg13g2_nor2_1 _15805_ (.A(_08312_),
    .B(_08316_),
    .Y(_08340_));
 sg13g2_xnor2_1 _15806_ (.Y(_08341_),
    .A(_08285_),
    .B(_08340_));
 sg13g2_nor2b_1 _15807_ (.A(_08339_),
    .B_N(_08341_),
    .Y(_08342_));
 sg13g2_xnor2_1 _15808_ (.Y(_08343_),
    .A(_08339_),
    .B(_08341_));
 sg13g2_xor2_1 _15809_ (.B(_08270_),
    .A(_08269_),
    .X(_08344_));
 sg13g2_a21o_1 _15810_ (.A2(_08344_),
    .A1(_08343_),
    .B1(_08342_),
    .X(_08345_));
 sg13g2_xor2_1 _15811_ (.B(_08318_),
    .A(_08317_),
    .X(_08346_));
 sg13g2_nand2_1 _15812_ (.Y(_08347_),
    .A(_08345_),
    .B(_08346_));
 sg13g2_a22oi_1 _15813_ (.Y(_08348_),
    .B1(_08304_),
    .B2(\spiking_network_top_uut.all_data_out[62] ),
    .A2(_08303_),
    .A1(\spiking_network_top_uut.all_data_out[60] ));
 sg13g2_nor2_1 _15814_ (.A(_08307_),
    .B(_08348_),
    .Y(_08349_));
 sg13g2_a22oi_1 _15815_ (.Y(_08350_),
    .B1(_08297_),
    .B2(\spiking_network_top_uut.all_data_out[56] ),
    .A2(_08296_),
    .A1(\spiking_network_top_uut.all_data_out[58] ));
 sg13g2_nor2_2 _15816_ (.A(_08301_),
    .B(_08350_),
    .Y(_08351_));
 sg13g2_and2_1 _15817_ (.A(_08349_),
    .B(_08351_),
    .X(_08352_));
 sg13g2_xor2_1 _15818_ (.B(_08292_),
    .A(_08291_),
    .X(_08353_));
 sg13g2_xor2_1 _15819_ (.B(_08351_),
    .A(_08349_),
    .X(_08354_));
 sg13g2_a21o_1 _15820_ (.A2(_08354_),
    .A1(_08353_),
    .B1(_08352_),
    .X(_08355_));
 sg13g2_o21ai_1 _15821_ (.B1(_08328_),
    .Y(_08356_),
    .A1(_08327_),
    .A2(_08330_));
 sg13g2_nand3_1 _15822_ (.B(_08355_),
    .C(_08356_),
    .A(_08332_),
    .Y(_08357_));
 sg13g2_xor2_1 _15823_ (.B(_08284_),
    .A(_08283_),
    .X(_08358_));
 sg13g2_inv_1 _15824_ (.Y(_08359_),
    .A(_08358_));
 sg13g2_a21oi_1 _15825_ (.A1(_08332_),
    .A2(_08356_),
    .Y(_08360_),
    .B1(_08355_));
 sg13g2_a21o_1 _15826_ (.A2(_08356_),
    .A1(_08332_),
    .B1(_08355_),
    .X(_08361_));
 sg13g2_nand3_1 _15827_ (.B(_08359_),
    .C(_08361_),
    .A(_08357_),
    .Y(_08362_));
 sg13g2_o21ai_1 _15828_ (.B1(_08357_),
    .Y(_08363_),
    .A1(_08358_),
    .A2(_08360_));
 sg13g2_xnor2_1 _15829_ (.Y(_08364_),
    .A(_08285_),
    .B(_08337_));
 sg13g2_nand2_1 _15830_ (.Y(_08365_),
    .A(_08363_),
    .B(_08364_));
 sg13g2_xnor2_1 _15831_ (.Y(_08366_),
    .A(_08363_),
    .B(_08364_));
 sg13g2_xor2_1 _15832_ (.B(_08267_),
    .A(_08266_),
    .X(_08367_));
 sg13g2_o21ai_1 _15833_ (.B1(_08365_),
    .Y(_08368_),
    .A1(_08366_),
    .A2(_08367_));
 sg13g2_xnor2_1 _15834_ (.Y(_08369_),
    .A(_08343_),
    .B(_08344_));
 sg13g2_nor2b_1 _15835_ (.A(_08369_),
    .B_N(_08368_),
    .Y(_08370_));
 sg13g2_xor2_1 _15836_ (.B(_08367_),
    .A(_08366_),
    .X(_08371_));
 sg13g2_xor2_1 _15837_ (.B(_08282_),
    .A(_08281_),
    .X(_08372_));
 sg13g2_xnor2_1 _15838_ (.Y(_08373_),
    .A(_08353_),
    .B(_08354_));
 sg13g2_inv_1 _15839_ (.Y(_08374_),
    .A(_08373_));
 sg13g2_a21o_2 _15840_ (.A2(_08361_),
    .A1(_08357_),
    .B1(_08359_),
    .X(_08375_));
 sg13g2_and4_1 _15841_ (.A(_08362_),
    .B(_08372_),
    .C(_08374_),
    .D(_08375_),
    .X(_08376_));
 sg13g2_nand4_1 _15842_ (.B(_08372_),
    .C(_08374_),
    .A(_08362_),
    .Y(_08377_),
    .D(_08375_));
 sg13g2_a22oi_1 _15843_ (.Y(_08378_),
    .B1(_08375_),
    .B2(_08362_),
    .A2(_08374_),
    .A1(_08372_));
 sg13g2_xnor2_1 _15844_ (.Y(_08379_),
    .A(_08264_),
    .B(_08265_));
 sg13g2_inv_1 _15845_ (.Y(_08380_),
    .A(_08379_));
 sg13g2_nor3_1 _15846_ (.A(_08376_),
    .B(_08378_),
    .C(_08379_),
    .Y(_08381_));
 sg13g2_o21ai_1 _15847_ (.B1(_08377_),
    .Y(_08382_),
    .A1(_08378_),
    .A2(_08379_));
 sg13g2_nand2_1 _15848_ (.Y(_08383_),
    .A(_08371_),
    .B(_08382_));
 sg13g2_o21ai_1 _15849_ (.B1(_08379_),
    .Y(_08384_),
    .A1(_08376_),
    .A2(_08378_));
 sg13g2_nor2b_1 _15850_ (.A(_08381_),
    .B_N(_08384_),
    .Y(_08385_));
 sg13g2_xnor2_1 _15851_ (.Y(_08386_),
    .A(_08372_),
    .B(_08373_));
 sg13g2_xor2_1 _15852_ (.B(_08263_),
    .A(_00100_),
    .X(_08387_));
 sg13g2_nor2b_1 _15853_ (.A(_08387_),
    .B_N(_08386_),
    .Y(_08388_));
 sg13g2_nand3b_1 _15854_ (.B(_08384_),
    .C(_08388_),
    .Y(_08389_),
    .A_N(_08381_));
 sg13g2_nor2_1 _15855_ (.A(_08371_),
    .B(_08382_),
    .Y(_08390_));
 sg13g2_xor2_1 _15856_ (.B(_08382_),
    .A(_08371_),
    .X(_08391_));
 sg13g2_o21ai_1 _15857_ (.B1(_08383_),
    .Y(_08392_),
    .A1(_08389_),
    .A2(_08390_));
 sg13g2_nand2b_1 _15858_ (.Y(_08393_),
    .B(_08369_),
    .A_N(_08368_));
 sg13g2_nand2b_1 _15859_ (.Y(_08394_),
    .B(_08393_),
    .A_N(_08370_));
 sg13g2_nand2b_1 _15860_ (.Y(_08395_),
    .B(_08392_),
    .A_N(_08394_));
 sg13g2_a21oi_1 _15861_ (.A1(_08392_),
    .A2(_08393_),
    .Y(_08396_),
    .B1(_08370_));
 sg13g2_xnor2_1 _15862_ (.Y(_08397_),
    .A(_08345_),
    .B(_08346_));
 sg13g2_o21ai_1 _15863_ (.B1(_08347_),
    .Y(_08398_),
    .A1(_08396_),
    .A2(_08397_));
 sg13g2_nand2_1 _15864_ (.Y(_08399_),
    .A(_08273_),
    .B(_08314_));
 sg13g2_nand2_1 _15865_ (.Y(_08400_),
    .A(_08313_),
    .B(_08320_));
 sg13g2_a221oi_1 _15866_ (.B2(_08400_),
    .C1(_08322_),
    .B1(_08399_),
    .A1(_08323_),
    .Y(_08401_),
    .A2(_08398_));
 sg13g2_o21ai_1 _15867_ (.B1(_08229_),
    .Y(_08402_),
    .A1(_08273_),
    .A2(_08313_));
 sg13g2_nor2_1 _15868_ (.A(_08401_),
    .B(_08402_),
    .Y(_08403_));
 sg13g2_nor2_1 _15869_ (.A(_08274_),
    .B(_08403_),
    .Y(_08404_));
 sg13g2_o21ai_1 _15870_ (.B1(_08275_),
    .Y(_08405_),
    .A1(_08401_),
    .A2(_08402_));
 sg13g2_xnor2_1 _15871_ (.Y(_08406_),
    .A(_08323_),
    .B(_08398_));
 sg13g2_a21oi_1 _15872_ (.A1(_08229_),
    .A2(_08406_),
    .Y(_08407_),
    .B1(_08274_));
 sg13g2_nand2_1 _15873_ (.Y(_08408_),
    .A(net3702),
    .B(_08318_));
 sg13g2_xnor2_1 _15874_ (.Y(_08409_),
    .A(_08396_),
    .B(_08397_));
 sg13g2_o21ai_1 _15875_ (.B1(_08408_),
    .Y(_08410_),
    .A1(net3702),
    .A2(_08409_));
 sg13g2_nand2_1 _15876_ (.Y(_08411_),
    .A(_08407_),
    .B(_08410_));
 sg13g2_a21oi_2 _15877_ (.B1(net3664),
    .Y(_08412_),
    .A2(_08411_),
    .A1(_08404_));
 sg13g2_nand2_1 _15878_ (.Y(_08413_),
    .A(net4605),
    .B(_08412_));
 sg13g2_o21ai_1 _15879_ (.B1(_08405_),
    .Y(_08414_),
    .A1(_08407_),
    .A2(_08410_));
 sg13g2_nand2_1 _15880_ (.Y(_08415_),
    .A(_08229_),
    .B(_08386_));
 sg13g2_xnor2_1 _15881_ (.Y(_08416_),
    .A(_08387_),
    .B(_08415_));
 sg13g2_and2_1 _15882_ (.A(_08414_),
    .B(_08416_),
    .X(_08417_));
 sg13g2_xor2_1 _15883_ (.B(net465),
    .A(net4315),
    .X(_08418_));
 sg13g2_a22oi_1 _15884_ (.Y(_08419_),
    .B1(_00002_),
    .B2(_08418_),
    .A2(net465),
    .A1(net3953));
 sg13g2_o21ai_1 _15885_ (.B1(_08419_),
    .Y(_00868_),
    .A1(_08413_),
    .A2(_08417_));
 sg13g2_xnor2_1 _15886_ (.Y(_08420_),
    .A(_08385_),
    .B(_08388_));
 sg13g2_o21ai_1 _15887_ (.B1(_08414_),
    .Y(_08421_),
    .A1(_08230_),
    .A2(_08420_));
 sg13g2_a21oi_1 _15888_ (.A1(net3702),
    .A2(_08380_),
    .Y(_08422_),
    .B1(_08421_));
 sg13g2_xor2_1 _15889_ (.B(_04876_),
    .A(_04875_),
    .X(_08423_));
 sg13g2_a22oi_1 _15890_ (.Y(_08424_),
    .B1(_00002_),
    .B2(_08423_),
    .A2(net531),
    .A1(net3953));
 sg13g2_o21ai_1 _15891_ (.B1(_08424_),
    .Y(_00869_),
    .A1(_08413_),
    .A2(_08422_));
 sg13g2_nand2_1 _15892_ (.Y(_08425_),
    .A(net3702),
    .B(_08367_));
 sg13g2_xnor2_1 _15893_ (.Y(_08426_),
    .A(_08389_),
    .B(_08391_));
 sg13g2_o21ai_1 _15894_ (.B1(_08425_),
    .Y(_08427_),
    .A1(net3702),
    .A2(_08426_));
 sg13g2_nand2_1 _15895_ (.Y(_08428_),
    .A(_08414_),
    .B(_08427_));
 sg13g2_nand3_1 _15896_ (.B(_04874_),
    .C(_04877_),
    .A(_04873_),
    .Y(_08429_));
 sg13g2_nor2b_1 _15897_ (.A(_04878_),
    .B_N(_08429_),
    .Y(_08430_));
 sg13g2_a221oi_1 _15898_ (.B2(net3664),
    .C1(net3953),
    .B1(_08430_),
    .A1(_08412_),
    .Y(_08431_),
    .A2(_08428_));
 sg13g2_a21oi_1 _15899_ (.A1(net3953),
    .A2(_03404_),
    .Y(_00870_),
    .B1(_08431_));
 sg13g2_nand2b_1 _15900_ (.Y(_08432_),
    .B(_08394_),
    .A_N(_08392_));
 sg13g2_nor2_1 _15901_ (.A(_08229_),
    .B(_08344_),
    .Y(_08433_));
 sg13g2_a21oi_1 _15902_ (.A1(_08395_),
    .A2(_08432_),
    .Y(_08434_),
    .B1(net3702));
 sg13g2_o21ai_1 _15903_ (.B1(_08414_),
    .Y(_08435_),
    .A1(_08433_),
    .A2(_08434_));
 sg13g2_or3_1 _15904_ (.A(_04871_),
    .B(_04872_),
    .C(_04878_),
    .X(_08436_));
 sg13g2_and2_1 _15905_ (.A(_04879_),
    .B(_08436_),
    .X(_08437_));
 sg13g2_a221oi_1 _15906_ (.B2(net3664),
    .C1(net3953),
    .B1(_08437_),
    .A1(_08412_),
    .Y(_08438_),
    .A2(_08435_));
 sg13g2_a21oi_1 _15907_ (.A1(net3954),
    .A2(_03403_),
    .Y(_00871_),
    .B1(_08438_));
 sg13g2_or2_1 _15908_ (.X(_08439_),
    .B(_04880_),
    .A(_04869_));
 sg13g2_o21ai_1 _15909_ (.B1(_08439_),
    .Y(_08440_),
    .A1(net3664),
    .A2(_08405_));
 sg13g2_mux2_1 _15910_ (.A0(net461),
    .A1(_08440_),
    .S(net4604),
    .X(_00872_));
 sg13g2_mux4_1 _15911_ (.S0(\spiking_network_top_uut.all_data_out[412] ),
    .A0(net3789),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[1] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[2] ),
    .A3(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[3] ),
    .S1(\spiking_network_top_uut.all_data_out[413] ),
    .X(_08441_));
 sg13g2_mux2_1 _15912_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[6] ),
    .A1(net3899),
    .S(\spiking_network_top_uut.all_data_out[412] ),
    .X(_08442_));
 sg13g2_nor2b_1 _15913_ (.A(\spiking_network_top_uut.all_data_out[412] ),
    .B_N(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[4] ),
    .Y(_08443_));
 sg13g2_a21oi_1 _15914_ (.A1(\spiking_network_top_uut.all_data_out[412] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[5] ),
    .Y(_08444_),
    .B1(_08443_));
 sg13g2_o21ai_1 _15915_ (.B1(\spiking_network_top_uut.all_data_out[414] ),
    .Y(_08445_),
    .A1(\spiking_network_top_uut.all_data_out[413] ),
    .A2(_08444_));
 sg13g2_a21oi_1 _15916_ (.A1(\spiking_network_top_uut.all_data_out[413] ),
    .A2(_08442_),
    .Y(_08446_),
    .B1(_08445_));
 sg13g2_o21ai_1 _15917_ (.B1(net4637),
    .Y(_08447_),
    .A1(\spiking_network_top_uut.all_data_out[414] ),
    .A2(_08441_));
 sg13g2_nand2_1 _15918_ (.Y(_08448_),
    .A(net3962),
    .B(net88));
 sg13g2_o21ai_1 _15919_ (.B1(_08448_),
    .Y(_00873_),
    .A1(_08446_),
    .A2(_08447_));
 sg13g2_mux2_1 _15920_ (.A0(net256),
    .A1(net88),
    .S(net4639),
    .X(_00874_));
 sg13g2_a21oi_1 _15921_ (.A1(\spiking_network_top_uut.all_data_out[408] ),
    .A2(_03662_),
    .Y(_08449_),
    .B1(\spiking_network_top_uut.all_data_out[409] ));
 sg13g2_o21ai_1 _15922_ (.B1(_08449_),
    .Y(_08450_),
    .A1(\spiking_network_top_uut.all_data_out[408] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[4] ));
 sg13g2_mux2_1 _15923_ (.A0(net3835),
    .A1(net3834),
    .S(\spiking_network_top_uut.all_data_out[408] ),
    .X(_08451_));
 sg13g2_nand2_1 _15924_ (.Y(_08452_),
    .A(\spiking_network_top_uut.all_data_out[409] ),
    .B(_08451_));
 sg13g2_nand3_1 _15925_ (.B(_08450_),
    .C(_08452_),
    .A(\spiking_network_top_uut.all_data_out[410] ),
    .Y(_08453_));
 sg13g2_mux2_1 _15926_ (.A0(net3838),
    .A1(net3837),
    .S(\spiking_network_top_uut.all_data_out[408] ),
    .X(_08454_));
 sg13g2_nor2b_1 _15927_ (.A(\spiking_network_top_uut.all_data_out[408] ),
    .B_N(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[0] ),
    .Y(_08455_));
 sg13g2_a21oi_1 _15928_ (.A1(\spiking_network_top_uut.all_data_out[408] ),
    .A2(net3839),
    .Y(_08456_),
    .B1(_08455_));
 sg13g2_a21oi_1 _15929_ (.A1(\spiking_network_top_uut.all_data_out[409] ),
    .A2(_08454_),
    .Y(_08457_),
    .B1(\spiking_network_top_uut.all_data_out[410] ));
 sg13g2_o21ai_1 _15930_ (.B1(_08457_),
    .Y(_08458_),
    .A1(\spiking_network_top_uut.all_data_out[409] ),
    .A2(_08456_));
 sg13g2_nand3_1 _15931_ (.B(_08453_),
    .C(_08458_),
    .A(net4642),
    .Y(_08459_));
 sg13g2_o21ai_1 _15932_ (.B1(_08459_),
    .Y(_00875_),
    .A1(net4643),
    .A2(_03685_));
 sg13g2_nor2_1 _15933_ (.A(net4639),
    .B(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_dout ),
    .Y(_08460_));
 sg13g2_a21oi_1 _15934_ (.A1(net4643),
    .A2(_03685_),
    .Y(_00876_),
    .B1(_08460_));
 sg13g2_mux4_1 _15935_ (.S0(\spiking_network_top_uut.all_data_out[404] ),
    .A0(net3833),
    .A1(net3832),
    .A2(net3831),
    .A3(net3830),
    .S1(\spiking_network_top_uut.all_data_out[405] ),
    .X(_08461_));
 sg13g2_mux2_1 _15936_ (.A0(net3828),
    .A1(net3827),
    .S(\spiking_network_top_uut.all_data_out[404] ),
    .X(_08462_));
 sg13g2_nor2b_1 _15937_ (.A(\spiking_network_top_uut.all_data_out[404] ),
    .B_N(net3829),
    .Y(_08463_));
 sg13g2_a21oi_1 _15938_ (.A1(\spiking_network_top_uut.all_data_out[404] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[5] ),
    .Y(_08464_),
    .B1(_08463_));
 sg13g2_o21ai_1 _15939_ (.B1(\spiking_network_top_uut.all_data_out[406] ),
    .Y(_08465_),
    .A1(\spiking_network_top_uut.all_data_out[405] ),
    .A2(_08464_));
 sg13g2_a21oi_1 _15940_ (.A1(\spiking_network_top_uut.all_data_out[405] ),
    .A2(_08462_),
    .Y(_08466_),
    .B1(_08465_));
 sg13g2_o21ai_1 _15941_ (.B1(net4610),
    .Y(_08467_),
    .A1(\spiking_network_top_uut.all_data_out[406] ),
    .A2(_08461_));
 sg13g2_nand2_1 _15942_ (.Y(_08468_),
    .A(net3966),
    .B(net138));
 sg13g2_o21ai_1 _15943_ (.B1(_08468_),
    .Y(_00877_),
    .A1(_08466_),
    .A2(_08467_));
 sg13g2_mux2_1 _15944_ (.A0(net236),
    .A1(net138),
    .S(net4611),
    .X(_00878_));
 sg13g2_a21oi_1 _15945_ (.A1(\spiking_network_top_uut.all_data_out[400] ),
    .A2(_03660_),
    .Y(_08469_),
    .B1(\spiking_network_top_uut.all_data_out[401] ));
 sg13g2_o21ai_1 _15946_ (.B1(_08469_),
    .Y(_08470_),
    .A1(\spiking_network_top_uut.all_data_out[400] ),
    .A2(net3822));
 sg13g2_mux2_1 _15947_ (.A0(net3821),
    .A1(net3820),
    .S(\spiking_network_top_uut.all_data_out[400] ),
    .X(_08471_));
 sg13g2_nand2_1 _15948_ (.Y(_08472_),
    .A(\spiking_network_top_uut.all_data_out[401] ),
    .B(_08471_));
 sg13g2_nand3_1 _15949_ (.B(_08470_),
    .C(_08472_),
    .A(\spiking_network_top_uut.all_data_out[402] ),
    .Y(_08473_));
 sg13g2_mux2_1 _15950_ (.A0(net3824),
    .A1(net3823),
    .S(\spiking_network_top_uut.all_data_out[400] ),
    .X(_08474_));
 sg13g2_nor2b_1 _15951_ (.A(\spiking_network_top_uut.all_data_out[400] ),
    .B_N(net3826),
    .Y(_08475_));
 sg13g2_a21oi_1 _15952_ (.A1(\spiking_network_top_uut.all_data_out[400] ),
    .A2(net3825),
    .Y(_08476_),
    .B1(_08475_));
 sg13g2_a21oi_1 _15953_ (.A1(\spiking_network_top_uut.all_data_out[401] ),
    .A2(_08474_),
    .Y(_08477_),
    .B1(\spiking_network_top_uut.all_data_out[402] ));
 sg13g2_o21ai_1 _15954_ (.B1(_08477_),
    .Y(_08478_),
    .A1(\spiking_network_top_uut.all_data_out[401] ),
    .A2(_08476_));
 sg13g2_nand3_1 _15955_ (.B(_08473_),
    .C(_08478_),
    .A(net4613),
    .Y(_08479_));
 sg13g2_o21ai_1 _15956_ (.B1(_08479_),
    .Y(_00879_),
    .A1(net4611),
    .A2(_03686_));
 sg13g2_nor2_1 _15957_ (.A(net4611),
    .B(net182),
    .Y(_08480_));
 sg13g2_a21oi_1 _15958_ (.A1(net4611),
    .A2(_03686_),
    .Y(_00880_),
    .B1(_08480_));
 sg13g2_nand2_1 _15959_ (.Y(_08481_),
    .A(\spiking_network_top_uut.all_data_out[396] ),
    .B(_03659_));
 sg13g2_nor2_1 _15960_ (.A(\spiking_network_top_uut.all_data_out[396] ),
    .B(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[4] ),
    .Y(_08482_));
 sg13g2_nor2_1 _15961_ (.A(\spiking_network_top_uut.all_data_out[397] ),
    .B(_08482_),
    .Y(_08483_));
 sg13g2_mux2_1 _15962_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[6] ),
    .A1(net3813),
    .S(\spiking_network_top_uut.all_data_out[396] ),
    .X(_08484_));
 sg13g2_a221oi_1 _15963_ (.B2(\spiking_network_top_uut.all_data_out[397] ),
    .C1(_03542_),
    .B1(_08484_),
    .A1(_08481_),
    .Y(_08485_),
    .A2(_08483_));
 sg13g2_mux4_1 _15964_ (.S0(\spiking_network_top_uut.all_data_out[396] ),
    .A0(net3819),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[1] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[2] ),
    .A3(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[3] ),
    .S1(\spiking_network_top_uut.all_data_out[397] ),
    .X(_08486_));
 sg13g2_o21ai_1 _15965_ (.B1(net4629),
    .Y(_08487_),
    .A1(\spiking_network_top_uut.all_data_out[398] ),
    .A2(_08486_));
 sg13g2_nand2_1 _15966_ (.Y(_08488_),
    .A(net3960),
    .B(net69));
 sg13g2_o21ai_1 _15967_ (.B1(_08488_),
    .Y(_00881_),
    .A1(_08485_),
    .A2(_08487_));
 sg13g2_mux2_1 _15968_ (.A0(net259),
    .A1(net69),
    .S(net4627),
    .X(_00882_));
 sg13g2_mux4_1 _15969_ (.S0(\spiking_network_top_uut.all_data_out[392] ),
    .A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[0] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[1] ),
    .A2(net3810),
    .A3(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[3] ),
    .S1(\spiking_network_top_uut.all_data_out[393] ),
    .X(_08489_));
 sg13g2_mux2_1 _15970_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[6] ),
    .A1(net3805),
    .S(\spiking_network_top_uut.all_data_out[392] ),
    .X(_08490_));
 sg13g2_nor2b_1 _15971_ (.A(\spiking_network_top_uut.all_data_out[392] ),
    .B_N(net3808),
    .Y(_08491_));
 sg13g2_a21oi_1 _15972_ (.A1(\spiking_network_top_uut.all_data_out[392] ),
    .A2(net3807),
    .Y(_08492_),
    .B1(_08491_));
 sg13g2_o21ai_1 _15973_ (.B1(\spiking_network_top_uut.all_data_out[394] ),
    .Y(_08493_),
    .A1(\spiking_network_top_uut.all_data_out[393] ),
    .A2(_08492_));
 sg13g2_a21oi_1 _15974_ (.A1(\spiking_network_top_uut.all_data_out[393] ),
    .A2(_08490_),
    .Y(_08494_),
    .B1(_08493_));
 sg13g2_o21ai_1 _15975_ (.B1(net4623),
    .Y(_08495_),
    .A1(\spiking_network_top_uut.all_data_out[394] ),
    .A2(_08489_));
 sg13g2_nand2_1 _15976_ (.Y(_08496_),
    .A(net3959),
    .B(net110));
 sg13g2_o21ai_1 _15977_ (.B1(_08496_),
    .Y(_00883_),
    .A1(_08494_),
    .A2(_08495_));
 sg13g2_mux2_1 _15978_ (.A0(net239),
    .A1(net110),
    .S(net4623),
    .X(_00884_));
 sg13g2_mux4_1 _15979_ (.S0(\spiking_network_top_uut.all_data_out[388] ),
    .A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[0] ),
    .A1(net3803),
    .A2(net3802),
    .A3(net3801),
    .S1(\spiking_network_top_uut.all_data_out[389] ),
    .X(_08497_));
 sg13g2_mux2_1 _15980_ (.A0(net3798),
    .A1(net3797),
    .S(\spiking_network_top_uut.all_data_out[388] ),
    .X(_08498_));
 sg13g2_nor2b_1 _15981_ (.A(\spiking_network_top_uut.all_data_out[388] ),
    .B_N(net3800),
    .Y(_08499_));
 sg13g2_a21oi_1 _15982_ (.A1(\spiking_network_top_uut.all_data_out[388] ),
    .A2(net3799),
    .Y(_08500_),
    .B1(_08499_));
 sg13g2_o21ai_1 _15983_ (.B1(\spiking_network_top_uut.all_data_out[390] ),
    .Y(_08501_),
    .A1(\spiking_network_top_uut.all_data_out[389] ),
    .A2(_08500_));
 sg13g2_a21oi_1 _15984_ (.A1(\spiking_network_top_uut.all_data_out[389] ),
    .A2(_08498_),
    .Y(_08502_),
    .B1(_08501_));
 sg13g2_o21ai_1 _15985_ (.B1(net4631),
    .Y(_08503_),
    .A1(\spiking_network_top_uut.all_data_out[390] ),
    .A2(_08497_));
 sg13g2_nand2_1 _15986_ (.Y(_08504_),
    .A(net3961),
    .B(net132));
 sg13g2_o21ai_1 _15987_ (.B1(_08504_),
    .Y(_00885_),
    .A1(_08502_),
    .A2(_08503_));
 sg13g2_mux2_1 _15988_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_dout ),
    .A1(net132),
    .S(net4632),
    .X(_00886_));
 sg13g2_mux4_1 _15989_ (.S0(\spiking_network_top_uut.all_data_out[384] ),
    .A0(net3796),
    .A1(net3795),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[2] ),
    .A3(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[3] ),
    .S1(\spiking_network_top_uut.all_data_out[385] ),
    .X(_08505_));
 sg13g2_mux2_1 _15990_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[6] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[7] ),
    .S(\spiking_network_top_uut.all_data_out[384] ),
    .X(_08506_));
 sg13g2_nor2b_1 _15991_ (.A(\spiking_network_top_uut.all_data_out[384] ),
    .B_N(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[4] ),
    .Y(_08507_));
 sg13g2_a21oi_1 _15992_ (.A1(\spiking_network_top_uut.all_data_out[384] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[5] ),
    .Y(_08508_),
    .B1(_08507_));
 sg13g2_o21ai_1 _15993_ (.B1(\spiking_network_top_uut.all_data_out[386] ),
    .Y(_08509_),
    .A1(\spiking_network_top_uut.all_data_out[385] ),
    .A2(_08508_));
 sg13g2_a21oi_1 _15994_ (.A1(\spiking_network_top_uut.all_data_out[385] ),
    .A2(_08506_),
    .Y(_08510_),
    .B1(_08509_));
 sg13g2_o21ai_1 _15995_ (.B1(net4635),
    .Y(_08511_),
    .A1(\spiking_network_top_uut.all_data_out[386] ),
    .A2(_08505_));
 sg13g2_nand2_1 _15996_ (.Y(_08512_),
    .A(net3964),
    .B(net144));
 sg13g2_o21ai_1 _15997_ (.B1(_08512_),
    .Y(_00887_),
    .A1(_08510_),
    .A2(_08511_));
 sg13g2_nor3_2 _15998_ (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[2] ),
    .B(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[1] ),
    .C(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[0] ),
    .Y(_08513_));
 sg13g2_nor2b_2 _15999_ (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[3] ),
    .B_N(_08513_),
    .Y(_08514_));
 sg13g2_nor2b_2 _16000_ (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[4] ),
    .B_N(_08514_),
    .Y(_08515_));
 sg13g2_nand2b_2 _16001_ (.Y(_08516_),
    .B(_08514_),
    .A_N(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[4] ));
 sg13g2_o21ai_1 _16002_ (.B1(net4605),
    .Y(_08517_),
    .A1(net3620),
    .A2(_08516_));
 sg13g2_nor2b_1 _16003_ (.A(net3620),
    .B_N(_00108_),
    .Y(_08518_));
 sg13g2_a21oi_1 _16004_ (.A1(net4285),
    .A2(net3621),
    .Y(_08519_),
    .B1(_08518_));
 sg13g2_nand2_1 _16005_ (.Y(_08520_),
    .A(net303),
    .B(_08517_));
 sg13g2_o21ai_1 _16006_ (.B1(_08520_),
    .Y(_00888_),
    .A1(_08517_),
    .A2(_08519_));
 sg13g2_xor2_1 _16007_ (.B(net303),
    .A(net393),
    .X(_08521_));
 sg13g2_nor2_1 _16008_ (.A(net3620),
    .B(_08521_),
    .Y(_08522_));
 sg13g2_a21oi_1 _16009_ (.A1(net4282),
    .A2(net3620),
    .Y(_08523_),
    .B1(_08522_));
 sg13g2_nand2_1 _16010_ (.Y(_08524_),
    .A(net393),
    .B(_08517_));
 sg13g2_o21ai_1 _16011_ (.B1(_08524_),
    .Y(_00889_),
    .A1(_08517_),
    .A2(_08523_));
 sg13g2_o21ai_1 _16012_ (.B1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[2] ),
    .Y(_08525_),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[1] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[0] ));
 sg13g2_nor2b_1 _16013_ (.A(_08513_),
    .B_N(_08525_),
    .Y(_08526_));
 sg13g2_nor2_1 _16014_ (.A(net3620),
    .B(_08526_),
    .Y(_08527_));
 sg13g2_a21oi_1 _16015_ (.A1(net4278),
    .A2(net3620),
    .Y(_08528_),
    .B1(_08527_));
 sg13g2_nand2_1 _16016_ (.Y(_08529_),
    .A(net194),
    .B(_08517_));
 sg13g2_o21ai_1 _16017_ (.B1(_08529_),
    .Y(_00890_),
    .A1(_08517_),
    .A2(_08528_));
 sg13g2_nand2_1 _16018_ (.Y(_08530_),
    .A(net4275),
    .B(net3621));
 sg13g2_xnor2_1 _16019_ (.Y(_08531_),
    .A(net426),
    .B(_08513_));
 sg13g2_o21ai_1 _16020_ (.B1(_08530_),
    .Y(_08532_),
    .A1(net3621),
    .A2(_08531_));
 sg13g2_mux2_1 _16021_ (.A0(_08532_),
    .A1(net426),
    .S(_08517_),
    .X(_00891_));
 sg13g2_nand2_1 _16022_ (.Y(_08533_),
    .A(net3954),
    .B(net287));
 sg13g2_nand2b_1 _16023_ (.Y(_08534_),
    .B(net287),
    .A_N(_08514_));
 sg13g2_a21oi_1 _16024_ (.A1(_08516_),
    .A2(_08534_),
    .Y(_08535_),
    .B1(net3620));
 sg13g2_a21oi_1 _16025_ (.A1(net4271),
    .A2(net3620),
    .Y(_08536_),
    .B1(_08535_));
 sg13g2_o21ai_1 _16026_ (.B1(_08533_),
    .Y(_00892_),
    .A1(_08517_),
    .A2(_08536_));
 sg13g2_mux2_1 _16027_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_dout ),
    .A1(net144),
    .S(net4635),
    .X(_00893_));
 sg13g2_nor2_2 _16028_ (.A(_00103_),
    .B(net3740),
    .Y(_08537_));
 sg13g2_nor2_2 _16029_ (.A(net3749),
    .B(_08537_),
    .Y(_08538_));
 sg13g2_nor2_1 _16030_ (.A(_00103_),
    .B(_08538_),
    .Y(_08539_));
 sg13g2_nand2b_1 _16031_ (.Y(_08540_),
    .B(_08538_),
    .A_N(_00103_));
 sg13g2_o21ai_1 _16032_ (.B1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ),
    .Y(_08541_),
    .A1(_00103_),
    .A2(_08538_));
 sg13g2_inv_1 _16033_ (.Y(_08542_),
    .A(_08541_));
 sg13g2_a21o_1 _16034_ (.A2(net3749),
    .A1(_00104_),
    .B1(_08538_),
    .X(_08543_));
 sg13g2_nand2_1 _16035_ (.Y(_08544_),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ),
    .B(_08543_));
 sg13g2_nor2_1 _16036_ (.A(_00104_),
    .B(net3908),
    .Y(_08545_));
 sg13g2_a221oi_1 _16037_ (.B2(_08537_),
    .C1(_08545_),
    .B1(net3907),
    .A1(_03497_),
    .Y(_08546_),
    .A2(net3749));
 sg13g2_o21ai_1 _16038_ (.B1(net3918),
    .Y(_08547_),
    .A1(_00103_),
    .A2(net3910));
 sg13g2_a221oi_1 _16039_ (.B2(_03496_),
    .C1(_08547_),
    .B1(net3902),
    .A1(_03497_),
    .Y(_08548_),
    .A2(net3738));
 sg13g2_and2_1 _16040_ (.A(_00107_),
    .B(net3752),
    .X(_08549_));
 sg13g2_nor3_2 _16041_ (.A(_03498_),
    .B(_08548_),
    .C(_08549_),
    .Y(_08550_));
 sg13g2_xnor2_1 _16042_ (.Y(_08551_),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ),
    .B(_08546_));
 sg13g2_nor2_1 _16043_ (.A(_08550_),
    .B(_08551_),
    .Y(_08552_));
 sg13g2_a21oi_1 _16044_ (.A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ),
    .A2(_08546_),
    .Y(_08553_),
    .B1(_08552_));
 sg13g2_xnor2_1 _16045_ (.Y(_08554_),
    .A(_03497_),
    .B(_08543_));
 sg13g2_o21ai_1 _16046_ (.B1(_08544_),
    .Y(_08555_),
    .A1(_08553_),
    .A2(_08554_));
 sg13g2_xnor2_1 _16047_ (.Y(_08556_),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ),
    .B(_08539_));
 sg13g2_a21oi_1 _16048_ (.A1(_08555_),
    .A2(_08556_),
    .Y(_08557_),
    .B1(_08542_));
 sg13g2_a22oi_1 _16049_ (.Y(_08558_),
    .B1(_08540_),
    .B2(_08557_),
    .A2(_08538_),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ));
 sg13g2_a21oi_2 _16050_ (.B1(_08558_),
    .Y(_08559_),
    .A2(_00103_),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ));
 sg13g2_nor2_1 _16051_ (.A(_08515_),
    .B(_08559_),
    .Y(_08560_));
 sg13g2_mux2_2 _16052_ (.A0(net4492),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[387] ),
    .X(_08561_));
 sg13g2_nand2_2 _16053_ (.Y(_08562_),
    .A(\spiking_network_top_uut.all_data_out[65] ),
    .B(_08561_));
 sg13g2_mux2_2 _16054_ (.A0(net4491),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[391] ),
    .X(_08563_));
 sg13g2_nand2_1 _16055_ (.Y(_08564_),
    .A(\spiking_network_top_uut.all_data_out[67] ),
    .B(_08563_));
 sg13g2_nor2_1 _16056_ (.A(_08562_),
    .B(_08564_),
    .Y(_08565_));
 sg13g2_nand4_1 _16057_ (.B(\spiking_network_top_uut.all_data_out[66] ),
    .C(_08561_),
    .A(\spiking_network_top_uut.all_data_out[64] ),
    .Y(_08566_),
    .D(_08563_));
 sg13g2_inv_1 _16058_ (.Y(_08567_),
    .A(_08566_));
 sg13g2_xor2_1 _16059_ (.B(_08564_),
    .A(_08562_),
    .X(_08568_));
 sg13g2_a21oi_2 _16060_ (.B1(_08565_),
    .Y(_08569_),
    .A2(_08568_),
    .A1(_08566_));
 sg13g2_mux2_2 _16061_ (.A0(net4489),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[399] ),
    .X(_08570_));
 sg13g2_nand2_1 _16062_ (.Y(_08571_),
    .A(\spiking_network_top_uut.all_data_out[71] ),
    .B(_08570_));
 sg13g2_mux2_2 _16063_ (.A0(net4490),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[395] ),
    .X(_08572_));
 sg13g2_nand2_1 _16064_ (.Y(_08573_),
    .A(\spiking_network_top_uut.all_data_out[69] ),
    .B(_08572_));
 sg13g2_nor2_1 _16065_ (.A(_08571_),
    .B(_08573_),
    .Y(_08574_));
 sg13g2_nand2_1 _16066_ (.Y(_08575_),
    .A(\spiking_network_top_uut.all_data_out[70] ),
    .B(_08570_));
 sg13g2_nand2_1 _16067_ (.Y(_08576_),
    .A(\spiking_network_top_uut.all_data_out[68] ),
    .B(_08572_));
 sg13g2_or2_2 _16068_ (.X(_08577_),
    .B(_08576_),
    .A(_08575_));
 sg13g2_xor2_1 _16069_ (.B(_08573_),
    .A(_08571_),
    .X(_08578_));
 sg13g2_a21oi_2 _16070_ (.B1(_08574_),
    .Y(_08579_),
    .A2(_08578_),
    .A1(_08577_));
 sg13g2_mux2_2 _16071_ (.A0(net4487),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[407] ),
    .X(_08580_));
 sg13g2_mux2_2 _16072_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.din ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[403] ),
    .X(_08581_));
 sg13g2_a22oi_1 _16073_ (.Y(_08582_),
    .B1(_08581_),
    .B2(\spiking_network_top_uut.all_data_out[73] ),
    .A2(_08580_),
    .A1(\spiking_network_top_uut.all_data_out[75] ));
 sg13g2_and4_1 _16074_ (.A(\spiking_network_top_uut.all_data_out[74] ),
    .B(\spiking_network_top_uut.all_data_out[72] ),
    .C(_08580_),
    .D(_08581_),
    .X(_08583_));
 sg13g2_nand4_1 _16075_ (.B(\spiking_network_top_uut.all_data_out[72] ),
    .C(_08580_),
    .A(\spiking_network_top_uut.all_data_out[74] ),
    .Y(_08584_),
    .D(_08581_));
 sg13g2_and4_1 _16076_ (.A(\spiking_network_top_uut.all_data_out[75] ),
    .B(\spiking_network_top_uut.all_data_out[73] ),
    .C(_08580_),
    .D(_08581_),
    .X(_08585_));
 sg13g2_nand4_1 _16077_ (.B(\spiking_network_top_uut.all_data_out[73] ),
    .C(_08580_),
    .A(\spiking_network_top_uut.all_data_out[75] ),
    .Y(_08586_),
    .D(_08581_));
 sg13g2_nand3b_1 _16078_ (.B(_08583_),
    .C(_08586_),
    .Y(_08587_),
    .A_N(_08582_));
 sg13g2_a21oi_2 _16079_ (.B1(_08582_),
    .Y(_08588_),
    .A2(_08586_),
    .A1(_08583_));
 sg13g2_mux2_2 _16080_ (.A0(net4485),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[415] ),
    .X(_08589_));
 sg13g2_mux2_2 _16081_ (.A0(net4486),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[411] ),
    .X(_08590_));
 sg13g2_and4_1 _16082_ (.A(\spiking_network_top_uut.all_data_out[79] ),
    .B(\spiking_network_top_uut.all_data_out[77] ),
    .C(_08589_),
    .D(_08590_),
    .X(_08591_));
 sg13g2_nand4_1 _16083_ (.B(\spiking_network_top_uut.all_data_out[77] ),
    .C(_08589_),
    .A(\spiking_network_top_uut.all_data_out[79] ),
    .Y(_08592_),
    .D(_08590_));
 sg13g2_and4_1 _16084_ (.A(\spiking_network_top_uut.all_data_out[78] ),
    .B(\spiking_network_top_uut.all_data_out[76] ),
    .C(_08589_),
    .D(_08590_),
    .X(_08593_));
 sg13g2_a22oi_1 _16085_ (.Y(_08594_),
    .B1(_08590_),
    .B2(\spiking_network_top_uut.all_data_out[77] ),
    .A2(_08589_),
    .A1(\spiking_network_top_uut.all_data_out[79] ));
 sg13g2_or3_2 _16086_ (.A(_08591_),
    .B(_08593_),
    .C(_08594_),
    .X(_08595_));
 sg13g2_o21ai_1 _16087_ (.B1(_08592_),
    .Y(_08596_),
    .A1(_08593_),
    .A2(_08594_));
 sg13g2_nand3b_1 _16088_ (.B(_08588_),
    .C(_08596_),
    .Y(_08597_),
    .A_N(_08579_));
 sg13g2_inv_1 _16089_ (.Y(_08598_),
    .A(_08597_));
 sg13g2_or2_1 _16090_ (.X(_08599_),
    .B(_08597_),
    .A(_08569_));
 sg13g2_nor2_1 _16091_ (.A(_08588_),
    .B(_08596_),
    .Y(_08600_));
 sg13g2_and2_1 _16092_ (.A(_08579_),
    .B(_08600_),
    .X(_08601_));
 sg13g2_nand2_1 _16093_ (.Y(_08602_),
    .A(_08569_),
    .B(_08601_));
 sg13g2_and2_1 _16094_ (.A(_08599_),
    .B(_08602_),
    .X(_08603_));
 sg13g2_xnor2_1 _16095_ (.Y(_08604_),
    .A(_08540_),
    .B(_08557_));
 sg13g2_nand2_1 _16096_ (.Y(_08605_),
    .A(_08603_),
    .B(_08604_));
 sg13g2_nand2_1 _16097_ (.Y(_08606_),
    .A(_08599_),
    .B(_08605_));
 sg13g2_xor2_1 _16098_ (.B(_08603_),
    .A(_08559_),
    .X(_08607_));
 sg13g2_nand2_1 _16099_ (.Y(_08608_),
    .A(_08606_),
    .B(_08607_));
 sg13g2_xnor2_1 _16100_ (.Y(_08609_),
    .A(_08603_),
    .B(_08604_));
 sg13g2_o21ai_1 _16101_ (.B1(_08593_),
    .Y(_08610_),
    .A1(_08591_),
    .A2(_08594_));
 sg13g2_o21ai_1 _16102_ (.B1(_08584_),
    .Y(_08611_),
    .A1(_08582_),
    .A2(_08585_));
 sg13g2_o21ai_1 _16103_ (.B1(_08583_),
    .Y(_08612_),
    .A1(_08582_),
    .A2(_08585_));
 sg13g2_nand3b_1 _16104_ (.B(_08584_),
    .C(_08586_),
    .Y(_08613_),
    .A_N(_08582_));
 sg13g2_a22oi_1 _16105_ (.Y(_08614_),
    .B1(_08612_),
    .B2(_08613_),
    .A2(_08610_),
    .A1(_08595_));
 sg13g2_xor2_1 _16106_ (.B(_08578_),
    .A(_08577_),
    .X(_08615_));
 sg13g2_xnor2_1 _16107_ (.Y(_08616_),
    .A(_08577_),
    .B(_08578_));
 sg13g2_and4_1 _16108_ (.A(_08595_),
    .B(_08610_),
    .C(_08612_),
    .D(_08613_),
    .X(_08617_));
 sg13g2_nand4_1 _16109_ (.B(_08610_),
    .C(_08612_),
    .A(_08595_),
    .Y(_08618_),
    .D(_08613_));
 sg13g2_and4_1 _16110_ (.A(_08587_),
    .B(_08595_),
    .C(_08610_),
    .D(_08611_),
    .X(_08619_));
 sg13g2_a22oi_1 _16111_ (.Y(_08620_),
    .B1(_08611_),
    .B2(_08587_),
    .A2(_08610_),
    .A1(_08595_));
 sg13g2_nor3_2 _16112_ (.A(_08614_),
    .B(_08615_),
    .C(_08617_),
    .Y(_08621_));
 sg13g2_a21oi_2 _16113_ (.B1(_08614_),
    .Y(_08622_),
    .A2(_08618_),
    .A1(_08616_));
 sg13g2_xor2_1 _16114_ (.B(_08596_),
    .A(_08588_),
    .X(_08623_));
 sg13g2_xnor2_1 _16115_ (.Y(_08624_),
    .A(_08579_),
    .B(_08623_));
 sg13g2_nand2b_1 _16116_ (.Y(_08625_),
    .B(_08624_),
    .A_N(_08622_));
 sg13g2_xnor2_1 _16117_ (.Y(_08626_),
    .A(_08622_),
    .B(_08624_));
 sg13g2_nand2b_1 _16118_ (.Y(_08627_),
    .B(_08626_),
    .A_N(_08569_));
 sg13g2_nand2_1 _16119_ (.Y(_08628_),
    .A(_08625_),
    .B(_08627_));
 sg13g2_nor2_1 _16120_ (.A(_08598_),
    .B(_08601_),
    .Y(_08629_));
 sg13g2_xnor2_1 _16121_ (.Y(_08630_),
    .A(_08569_),
    .B(_08629_));
 sg13g2_and2_1 _16122_ (.A(_08628_),
    .B(_08630_),
    .X(_08631_));
 sg13g2_xor2_1 _16123_ (.B(_08630_),
    .A(_08628_),
    .X(_08632_));
 sg13g2_xnor2_1 _16124_ (.Y(_08633_),
    .A(_08555_),
    .B(_08556_));
 sg13g2_inv_1 _16125_ (.Y(_08634_),
    .A(_08633_));
 sg13g2_a21oi_1 _16126_ (.A1(_08632_),
    .A2(_08634_),
    .Y(_08635_),
    .B1(_08631_));
 sg13g2_nor2_1 _16127_ (.A(_08609_),
    .B(_08635_),
    .Y(_08636_));
 sg13g2_xnor2_1 _16128_ (.Y(_08637_),
    .A(_08632_),
    .B(_08633_));
 sg13g2_a22oi_1 _16129_ (.Y(_08638_),
    .B1(_08590_),
    .B2(\spiking_network_top_uut.all_data_out[76] ),
    .A2(_08589_),
    .A1(\spiking_network_top_uut.all_data_out[78] ));
 sg13g2_nor2_1 _16130_ (.A(_08593_),
    .B(_08638_),
    .Y(_08639_));
 sg13g2_a22oi_1 _16131_ (.Y(_08640_),
    .B1(_08581_),
    .B2(\spiking_network_top_uut.all_data_out[72] ),
    .A2(_08580_),
    .A1(\spiking_network_top_uut.all_data_out[74] ));
 sg13g2_nor2_1 _16132_ (.A(_08583_),
    .B(_08640_),
    .Y(_08641_));
 sg13g2_and2_1 _16133_ (.A(_08639_),
    .B(_08641_),
    .X(_08642_));
 sg13g2_xor2_1 _16134_ (.B(_08576_),
    .A(_08575_),
    .X(_08643_));
 sg13g2_xor2_1 _16135_ (.B(_08641_),
    .A(_08639_),
    .X(_08644_));
 sg13g2_a21oi_2 _16136_ (.B1(_08642_),
    .Y(_08645_),
    .A2(_08644_),
    .A1(_08643_));
 sg13g2_nor3_2 _16137_ (.A(_08616_),
    .B(_08619_),
    .C(_08620_),
    .Y(_08646_));
 sg13g2_nor3_1 _16138_ (.A(_08621_),
    .B(_08645_),
    .C(_08646_),
    .Y(_08647_));
 sg13g2_or3_1 _16139_ (.A(_08621_),
    .B(_08645_),
    .C(_08646_),
    .X(_08648_));
 sg13g2_xnor2_1 _16140_ (.Y(_08649_),
    .A(_08566_),
    .B(_08568_));
 sg13g2_o21ai_1 _16141_ (.B1(_08645_),
    .Y(_08650_),
    .A1(_08621_),
    .A2(_08646_));
 sg13g2_nand3_1 _16142_ (.B(_08649_),
    .C(_08650_),
    .A(_08648_),
    .Y(_08651_));
 sg13g2_a21o_2 _16143_ (.A2(_08650_),
    .A1(_08649_),
    .B1(_08647_),
    .X(_08652_));
 sg13g2_xnor2_1 _16144_ (.Y(_08653_),
    .A(_08569_),
    .B(_08626_));
 sg13g2_xnor2_1 _16145_ (.Y(_08654_),
    .A(_08652_),
    .B(_08653_));
 sg13g2_xor2_1 _16146_ (.B(_08554_),
    .A(_08553_),
    .X(_08655_));
 sg13g2_nor2b_1 _16147_ (.A(_08654_),
    .B_N(_08655_),
    .Y(_08656_));
 sg13g2_a21o_1 _16148_ (.A2(_08653_),
    .A1(_08652_),
    .B1(_08656_),
    .X(_08657_));
 sg13g2_nand2_1 _16149_ (.Y(_08658_),
    .A(_08637_),
    .B(_08657_));
 sg13g2_a22oi_1 _16150_ (.Y(_08659_),
    .B1(_08563_),
    .B2(\spiking_network_top_uut.all_data_out[66] ),
    .A2(_08561_),
    .A1(\spiking_network_top_uut.all_data_out[64] ));
 sg13g2_xnor2_1 _16151_ (.Y(_08660_),
    .A(_08643_),
    .B(_08644_));
 sg13g2_nor3_2 _16152_ (.A(_08567_),
    .B(_08659_),
    .C(_08660_),
    .Y(_08661_));
 sg13g2_a21o_2 _16153_ (.A2(_08650_),
    .A1(_08648_),
    .B1(_08649_),
    .X(_08662_));
 sg13g2_nand3_1 _16154_ (.B(_08661_),
    .C(_08662_),
    .A(_08651_),
    .Y(_08663_));
 sg13g2_a21oi_1 _16155_ (.A1(_08651_),
    .A2(_08662_),
    .Y(_08664_),
    .B1(_08661_));
 sg13g2_a21o_1 _16156_ (.A2(_08662_),
    .A1(_08651_),
    .B1(_08661_),
    .X(_08665_));
 sg13g2_xor2_1 _16157_ (.B(_08551_),
    .A(_08550_),
    .X(_08666_));
 sg13g2_xnor2_1 _16158_ (.Y(_08667_),
    .A(_08550_),
    .B(_08551_));
 sg13g2_and3_1 _16159_ (.X(_08668_),
    .A(_08663_),
    .B(_08665_),
    .C(_08666_));
 sg13g2_o21ai_1 _16160_ (.B1(_08663_),
    .Y(_08669_),
    .A1(_08664_),
    .A2(_08667_));
 sg13g2_xnor2_1 _16161_ (.Y(_08670_),
    .A(_08654_),
    .B(_08655_));
 sg13g2_and2_1 _16162_ (.A(_08669_),
    .B(_08670_),
    .X(_08671_));
 sg13g2_a21oi_1 _16163_ (.A1(_08663_),
    .A2(_08665_),
    .Y(_08672_),
    .B1(_08666_));
 sg13g2_o21ai_1 _16164_ (.B1(_08660_),
    .Y(_08673_),
    .A1(_08567_),
    .A2(_08659_));
 sg13g2_nand2b_2 _16165_ (.Y(_08674_),
    .B(_08673_),
    .A_N(_08661_));
 sg13g2_o21ai_1 _16166_ (.B1(_03498_),
    .Y(_08675_),
    .A1(_08548_),
    .A2(_08549_));
 sg13g2_nand2b_1 _16167_ (.Y(_08676_),
    .B(_08675_),
    .A_N(_08550_));
 sg13g2_nand2b_1 _16168_ (.Y(_08677_),
    .B(_08676_),
    .A_N(_08674_));
 sg13g2_nor3_2 _16169_ (.A(_08668_),
    .B(_08672_),
    .C(_08677_),
    .Y(_08678_));
 sg13g2_or2_1 _16170_ (.X(_08679_),
    .B(_08670_),
    .A(_08669_));
 sg13g2_nand2b_1 _16171_ (.Y(_08680_),
    .B(_08679_),
    .A_N(_08671_));
 sg13g2_a21oi_2 _16172_ (.B1(_08671_),
    .Y(_08681_),
    .A2(_08679_),
    .A1(_08678_));
 sg13g2_xnor2_1 _16173_ (.Y(_08682_),
    .A(_08637_),
    .B(_08657_));
 sg13g2_o21ai_1 _16174_ (.B1(_08658_),
    .Y(_08683_),
    .A1(_08681_),
    .A2(_08682_));
 sg13g2_xor2_1 _16175_ (.B(_08635_),
    .A(_08609_),
    .X(_08684_));
 sg13g2_a21oi_1 _16176_ (.A1(_08683_),
    .A2(_08684_),
    .Y(_08685_),
    .B1(_08636_));
 sg13g2_xnor2_1 _16177_ (.Y(_08686_),
    .A(_08606_),
    .B(_08607_));
 sg13g2_o21ai_1 _16178_ (.B1(_08608_),
    .Y(_08687_),
    .A1(_08685_),
    .A2(_08686_));
 sg13g2_mux2_1 _16179_ (.A0(_08602_),
    .A1(_08599_),
    .S(_08559_),
    .X(_08688_));
 sg13g2_xnor2_1 _16180_ (.Y(_08689_),
    .A(_08687_),
    .B(_08688_));
 sg13g2_a21oi_2 _16181_ (.B1(_08560_),
    .Y(_08690_),
    .A2(_08689_),
    .A1(_08515_));
 sg13g2_xnor2_1 _16182_ (.Y(_08691_),
    .A(_08685_),
    .B(_08686_));
 sg13g2_a21oi_1 _16183_ (.A1(_08515_),
    .A2(_08691_),
    .Y(_08692_),
    .B1(_08560_));
 sg13g2_nor2_1 _16184_ (.A(_08515_),
    .B(_08604_),
    .Y(_08693_));
 sg13g2_xnor2_1 _16185_ (.Y(_08694_),
    .A(_08683_),
    .B(_08684_));
 sg13g2_a21oi_1 _16186_ (.A1(_08515_),
    .A2(_08694_),
    .Y(_08695_),
    .B1(_08693_));
 sg13g2_nand2_1 _16187_ (.Y(_08696_),
    .A(_08692_),
    .B(_08695_));
 sg13g2_a21oi_1 _16188_ (.A1(_08690_),
    .A2(_08696_),
    .Y(_08697_),
    .B1(net3622));
 sg13g2_nor2_1 _16189_ (.A(_08692_),
    .B(_08695_),
    .Y(_08698_));
 sg13g2_nor2_2 _16190_ (.A(_08690_),
    .B(_08698_),
    .Y(_08699_));
 sg13g2_nor2_1 _16191_ (.A(_08516_),
    .B(_08674_),
    .Y(_08700_));
 sg13g2_xor2_1 _16192_ (.B(_08700_),
    .A(_08676_),
    .X(_08701_));
 sg13g2_o21ai_1 _16193_ (.B1(_08697_),
    .Y(_08702_),
    .A1(_08699_),
    .A2(_08701_));
 sg13g2_xor2_1 _16194_ (.B(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[0] ),
    .A(net4315),
    .X(_08703_));
 sg13g2_a21oi_1 _16195_ (.A1(net3622),
    .A2(_08703_),
    .Y(_08704_),
    .B1(net3952));
 sg13g2_a22oi_1 _16196_ (.Y(_00894_),
    .B1(_08702_),
    .B2(_08704_),
    .A2(_03468_),
    .A1(net3952));
 sg13g2_o21ai_1 _16197_ (.B1(_08677_),
    .Y(_08705_),
    .A1(_08668_),
    .A2(_08672_));
 sg13g2_nor2_1 _16198_ (.A(_08516_),
    .B(_08678_),
    .Y(_08706_));
 sg13g2_a221oi_1 _16199_ (.B2(_08706_),
    .C1(_08699_),
    .B1(_08705_),
    .A1(_08516_),
    .Y(_08707_),
    .A2(_08666_));
 sg13g2_nand2_1 _16200_ (.Y(_08708_),
    .A(net4605),
    .B(_08697_));
 sg13g2_xor2_1 _16201_ (.B(_04886_),
    .A(_04885_),
    .X(_08709_));
 sg13g2_a22oi_1 _16202_ (.Y(_08710_),
    .B1(_00003_),
    .B2(_08709_),
    .A2(net543),
    .A1(net3954));
 sg13g2_o21ai_1 _16203_ (.B1(_08710_),
    .Y(_00895_),
    .A1(_08707_),
    .A2(_08708_));
 sg13g2_nor2_1 _16204_ (.A(_08515_),
    .B(_08655_),
    .Y(_08711_));
 sg13g2_xor2_1 _16205_ (.B(_08680_),
    .A(_08678_),
    .X(_08712_));
 sg13g2_a21oi_1 _16206_ (.A1(_08515_),
    .A2(_08712_),
    .Y(_08713_),
    .B1(_08711_));
 sg13g2_nor2_1 _16207_ (.A(_08699_),
    .B(_08713_),
    .Y(_08714_));
 sg13g2_xnor2_1 _16208_ (.Y(_08715_),
    .A(_04888_),
    .B(_04889_));
 sg13g2_a22oi_1 _16209_ (.Y(_08716_),
    .B1(_00003_),
    .B2(_08715_),
    .A2(net503),
    .A1(net3952));
 sg13g2_o21ai_1 _16210_ (.B1(_08716_),
    .Y(_00896_),
    .A1(_08708_),
    .A2(_08714_));
 sg13g2_xor2_1 _16211_ (.B(_08682_),
    .A(_08681_),
    .X(_08717_));
 sg13g2_mux2_1 _16212_ (.A0(_08634_),
    .A1(_08717_),
    .S(_08515_),
    .X(_08718_));
 sg13g2_nor2_1 _16213_ (.A(_08699_),
    .B(_08718_),
    .Y(_08719_));
 sg13g2_or3_1 _16214_ (.A(_04883_),
    .B(_04884_),
    .C(_04890_),
    .X(_08720_));
 sg13g2_and2_1 _16215_ (.A(_04891_),
    .B(_08720_),
    .X(_08721_));
 sg13g2_a22oi_1 _16216_ (.Y(_08722_),
    .B1(_00003_),
    .B2(_08721_),
    .A2(net549),
    .A1(net3952));
 sg13g2_o21ai_1 _16217_ (.B1(_08722_),
    .Y(_00897_),
    .A1(_08708_),
    .A2(_08719_));
 sg13g2_nand2b_1 _16218_ (.Y(_08723_),
    .B(_08690_),
    .A_N(net3622));
 sg13g2_a21oi_1 _16219_ (.A1(_04882_),
    .A2(_04892_),
    .Y(_08724_),
    .B1(net3951));
 sg13g2_a22oi_1 _16220_ (.Y(_00898_),
    .B1(_08723_),
    .B2(_08724_),
    .A2(_03466_),
    .A1(net3951));
 sg13g2_mux4_1 _16221_ (.S0(\spiking_network_top_uut.all_data_out[444] ),
    .A0(net3789),
    .A1(net3788),
    .A2(net3787),
    .A3(net3786),
    .S1(\spiking_network_top_uut.all_data_out[445] ),
    .X(_08725_));
 sg13g2_mux2_1 _16222_ (.A0(net3783),
    .A1(net3899),
    .S(\spiking_network_top_uut.all_data_out[444] ),
    .X(_08726_));
 sg13g2_nor2b_1 _16223_ (.A(\spiking_network_top_uut.all_data_out[444] ),
    .B_N(net3785),
    .Y(_08727_));
 sg13g2_a21oi_1 _16224_ (.A1(\spiking_network_top_uut.all_data_out[444] ),
    .A2(net3784),
    .Y(_08728_),
    .B1(_08727_));
 sg13g2_o21ai_1 _16225_ (.B1(\spiking_network_top_uut.all_data_out[446] ),
    .Y(_08729_),
    .A1(\spiking_network_top_uut.all_data_out[445] ),
    .A2(_08728_));
 sg13g2_a21oi_1 _16226_ (.A1(\spiking_network_top_uut.all_data_out[445] ),
    .A2(_08726_),
    .Y(_08730_),
    .B1(_08729_));
 sg13g2_o21ai_1 _16227_ (.B1(net4638),
    .Y(_08731_),
    .A1(\spiking_network_top_uut.all_data_out[446] ),
    .A2(_08725_));
 sg13g2_nand2_1 _16228_ (.Y(_08732_),
    .A(net3962),
    .B(net198));
 sg13g2_o21ai_1 _16229_ (.B1(_08732_),
    .Y(_00899_),
    .A1(_08730_),
    .A2(_08731_));
 sg13g2_mux2_1 _16230_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_dout ),
    .A1(net198),
    .S(net4639),
    .X(_00900_));
 sg13g2_mux4_1 _16231_ (.S0(\spiking_network_top_uut.all_data_out[440] ),
    .A0(net3840),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[1] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[2] ),
    .A3(net3837),
    .S1(\spiking_network_top_uut.all_data_out[441] ),
    .X(_08733_));
 sg13g2_mux2_1 _16232_ (.A0(net3835),
    .A1(net3834),
    .S(\spiking_network_top_uut.all_data_out[440] ),
    .X(_08734_));
 sg13g2_nor2b_1 _16233_ (.A(\spiking_network_top_uut.all_data_out[440] ),
    .B_N(net3836),
    .Y(_08735_));
 sg13g2_a21oi_1 _16234_ (.A1(\spiking_network_top_uut.all_data_out[440] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[5] ),
    .Y(_08736_),
    .B1(_08735_));
 sg13g2_o21ai_1 _16235_ (.B1(\spiking_network_top_uut.all_data_out[442] ),
    .Y(_08737_),
    .A1(\spiking_network_top_uut.all_data_out[441] ),
    .A2(_08736_));
 sg13g2_a21oi_1 _16236_ (.A1(\spiking_network_top_uut.all_data_out[441] ),
    .A2(_08734_),
    .Y(_08738_),
    .B1(_08737_));
 sg13g2_o21ai_1 _16237_ (.B1(net4640),
    .Y(_08739_),
    .A1(\spiking_network_top_uut.all_data_out[442] ),
    .A2(_08733_));
 sg13g2_nand2_1 _16238_ (.Y(_08740_),
    .A(net3963),
    .B(net180));
 sg13g2_o21ai_1 _16239_ (.B1(_08740_),
    .Y(_00901_),
    .A1(_08738_),
    .A2(_08739_));
 sg13g2_mux2_1 _16240_ (.A0(net243),
    .A1(net180),
    .S(net4640),
    .X(_00902_));
 sg13g2_nand2_1 _16241_ (.Y(_08741_),
    .A(\spiking_network_top_uut.all_data_out[436] ),
    .B(_03661_));
 sg13g2_nor2_1 _16242_ (.A(\spiking_network_top_uut.all_data_out[436] ),
    .B(net3829),
    .Y(_08742_));
 sg13g2_nor2_1 _16243_ (.A(\spiking_network_top_uut.all_data_out[437] ),
    .B(_08742_),
    .Y(_08743_));
 sg13g2_mux2_1 _16244_ (.A0(net3828),
    .A1(net3827),
    .S(\spiking_network_top_uut.all_data_out[436] ),
    .X(_08744_));
 sg13g2_a221oi_1 _16245_ (.B2(\spiking_network_top_uut.all_data_out[437] ),
    .C1(_03539_),
    .B1(_08744_),
    .A1(_08741_),
    .Y(_08745_),
    .A2(_08743_));
 sg13g2_mux4_1 _16246_ (.S0(\spiking_network_top_uut.all_data_out[436] ),
    .A0(net3833),
    .A1(net3832),
    .A2(net3831),
    .A3(net3830),
    .S1(\spiking_network_top_uut.all_data_out[437] ),
    .X(_08746_));
 sg13g2_o21ai_1 _16247_ (.B1(net4607),
    .Y(_08747_),
    .A1(\spiking_network_top_uut.all_data_out[438] ),
    .A2(_08746_));
 sg13g2_nand2_1 _16248_ (.Y(_08748_),
    .A(net3966),
    .B(net228));
 sg13g2_o21ai_1 _16249_ (.B1(_08748_),
    .Y(_00903_),
    .A1(_08745_),
    .A2(_08747_));
 sg13g2_mux2_1 _16250_ (.A0(net162),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_reg1 ),
    .S(net4608),
    .X(_00904_));
 sg13g2_mux4_1 _16251_ (.S0(\spiking_network_top_uut.all_data_out[432] ),
    .A0(net3826),
    .A1(net3825),
    .A2(net3824),
    .A3(net3823),
    .S1(\spiking_network_top_uut.all_data_out[433] ),
    .X(_08749_));
 sg13g2_mux2_1 _16252_ (.A0(net3821),
    .A1(net3820),
    .S(\spiking_network_top_uut.all_data_out[432] ),
    .X(_08750_));
 sg13g2_nor2b_1 _16253_ (.A(\spiking_network_top_uut.all_data_out[432] ),
    .B_N(net3822),
    .Y(_08751_));
 sg13g2_a21oi_1 _16254_ (.A1(\spiking_network_top_uut.all_data_out[432] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[5] ),
    .Y(_08752_),
    .B1(_08751_));
 sg13g2_o21ai_1 _16255_ (.B1(\spiking_network_top_uut.all_data_out[434] ),
    .Y(_08753_),
    .A1(\spiking_network_top_uut.all_data_out[433] ),
    .A2(_08752_));
 sg13g2_a21oi_1 _16256_ (.A1(\spiking_network_top_uut.all_data_out[433] ),
    .A2(_08750_),
    .Y(_08754_),
    .B1(_08753_));
 sg13g2_o21ai_1 _16257_ (.B1(net4613),
    .Y(_08755_),
    .A1(\spiking_network_top_uut.all_data_out[434] ),
    .A2(_08749_));
 sg13g2_nand2_1 _16258_ (.Y(_08756_),
    .A(net3965),
    .B(net188));
 sg13g2_o21ai_1 _16259_ (.B1(_08756_),
    .Y(_00905_),
    .A1(_08754_),
    .A2(_08755_));
 sg13g2_mux2_1 _16260_ (.A0(net191),
    .A1(net188),
    .S(net4616),
    .X(_00906_));
 sg13g2_nand2_1 _16261_ (.Y(_08757_),
    .A(\spiking_network_top_uut.all_data_out[428] ),
    .B(_03659_));
 sg13g2_nor2_1 _16262_ (.A(\spiking_network_top_uut.all_data_out[428] ),
    .B(net3815),
    .Y(_08758_));
 sg13g2_nor2_1 _16263_ (.A(\spiking_network_top_uut.all_data_out[429] ),
    .B(_08758_),
    .Y(_08759_));
 sg13g2_mux2_1 _16264_ (.A0(net3814),
    .A1(net3813),
    .S(\spiking_network_top_uut.all_data_out[428] ),
    .X(_08760_));
 sg13g2_a221oi_1 _16265_ (.B2(\spiking_network_top_uut.all_data_out[429] ),
    .C1(_03540_),
    .B1(_08760_),
    .A1(_08757_),
    .Y(_08761_),
    .A2(_08759_));
 sg13g2_mux4_1 _16266_ (.S0(\spiking_network_top_uut.all_data_out[428] ),
    .A0(net3819),
    .A1(net3818),
    .A2(net3817),
    .A3(net3816),
    .S1(\spiking_network_top_uut.all_data_out[429] ),
    .X(_08762_));
 sg13g2_o21ai_1 _16267_ (.B1(net4625),
    .Y(_08763_),
    .A1(\spiking_network_top_uut.all_data_out[430] ),
    .A2(_08762_));
 sg13g2_nand2_1 _16268_ (.Y(_08764_),
    .A(net3960),
    .B(net161));
 sg13g2_o21ai_1 _16269_ (.B1(_08764_),
    .Y(_00907_),
    .A1(_08761_),
    .A2(_08763_));
 sg13g2_mux2_1 _16270_ (.A0(net223),
    .A1(net161),
    .S(net4625),
    .X(_00908_));
 sg13g2_mux2_1 _16271_ (.A0(net3810),
    .A1(net3809),
    .S(\spiking_network_top_uut.all_data_out[424] ),
    .X(_08765_));
 sg13g2_nor2b_1 _16272_ (.A(\spiking_network_top_uut.all_data_out[424] ),
    .B_N(net3812),
    .Y(_08766_));
 sg13g2_a21oi_1 _16273_ (.A1(\spiking_network_top_uut.all_data_out[424] ),
    .A2(net3811),
    .Y(_08767_),
    .B1(_08766_));
 sg13g2_a21oi_1 _16274_ (.A1(\spiking_network_top_uut.all_data_out[425] ),
    .A2(_08765_),
    .Y(_08768_),
    .B1(\spiking_network_top_uut.all_data_out[426] ));
 sg13g2_o21ai_1 _16275_ (.B1(_08768_),
    .Y(_08769_),
    .A1(\spiking_network_top_uut.all_data_out[425] ),
    .A2(_08767_));
 sg13g2_mux2_1 _16276_ (.A0(net3806),
    .A1(net3805),
    .S(\spiking_network_top_uut.all_data_out[424] ),
    .X(_08770_));
 sg13g2_nor2b_1 _16277_ (.A(\spiking_network_top_uut.all_data_out[424] ),
    .B_N(net3808),
    .Y(_08771_));
 sg13g2_a21oi_1 _16278_ (.A1(\spiking_network_top_uut.all_data_out[424] ),
    .A2(net3807),
    .Y(_08772_),
    .B1(_08771_));
 sg13g2_o21ai_1 _16279_ (.B1(\spiking_network_top_uut.all_data_out[426] ),
    .Y(_08773_),
    .A1(\spiking_network_top_uut.all_data_out[425] ),
    .A2(_08772_));
 sg13g2_a21oi_1 _16280_ (.A1(\spiking_network_top_uut.all_data_out[425] ),
    .A2(_08770_),
    .Y(_08774_),
    .B1(_08773_));
 sg13g2_nand2_1 _16281_ (.Y(_08775_),
    .A(net4621),
    .B(_08769_));
 sg13g2_nand2_1 _16282_ (.Y(_08776_),
    .A(net3959),
    .B(net89));
 sg13g2_o21ai_1 _16283_ (.B1(_08776_),
    .Y(_00909_),
    .A1(_08774_),
    .A2(_08775_));
 sg13g2_mux2_1 _16284_ (.A0(net336),
    .A1(net89),
    .S(net4624),
    .X(_00910_));
 sg13g2_mux2_1 _16285_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[2] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[3] ),
    .S(\spiking_network_top_uut.all_data_out[420] ),
    .X(_08777_));
 sg13g2_nor2b_1 _16286_ (.A(\spiking_network_top_uut.all_data_out[420] ),
    .B_N(net3804),
    .Y(_08778_));
 sg13g2_a21oi_1 _16287_ (.A1(\spiking_network_top_uut.all_data_out[420] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[1] ),
    .Y(_08779_),
    .B1(_08778_));
 sg13g2_a21oi_1 _16288_ (.A1(\spiking_network_top_uut.all_data_out[421] ),
    .A2(_08777_),
    .Y(_08780_),
    .B1(\spiking_network_top_uut.all_data_out[422] ));
 sg13g2_o21ai_1 _16289_ (.B1(_08780_),
    .Y(_08781_),
    .A1(\spiking_network_top_uut.all_data_out[421] ),
    .A2(_08779_));
 sg13g2_mux2_1 _16290_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[6] ),
    .A1(net3797),
    .S(\spiking_network_top_uut.all_data_out[420] ),
    .X(_08782_));
 sg13g2_nor2b_1 _16291_ (.A(\spiking_network_top_uut.all_data_out[420] ),
    .B_N(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[4] ),
    .Y(_08783_));
 sg13g2_a21oi_1 _16292_ (.A1(\spiking_network_top_uut.all_data_out[420] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[5] ),
    .Y(_08784_),
    .B1(_08783_));
 sg13g2_o21ai_1 _16293_ (.B1(\spiking_network_top_uut.all_data_out[422] ),
    .Y(_08785_),
    .A1(\spiking_network_top_uut.all_data_out[421] ),
    .A2(_08784_));
 sg13g2_a21oi_1 _16294_ (.A1(\spiking_network_top_uut.all_data_out[421] ),
    .A2(_08782_),
    .Y(_08786_),
    .B1(_08785_));
 sg13g2_nand2_1 _16295_ (.Y(_08787_),
    .A(net4632),
    .B(_08781_));
 sg13g2_nand2_1 _16296_ (.Y(_08788_),
    .A(net3961),
    .B(net41));
 sg13g2_o21ai_1 _16297_ (.B1(_08788_),
    .Y(_00911_),
    .A1(_08786_),
    .A2(_08787_));
 sg13g2_mux2_1 _16298_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_dout ),
    .A1(net41),
    .S(net4635),
    .X(_00912_));
 sg13g2_mux2_1 _16299_ (.A0(net3794),
    .A1(net3793),
    .S(\spiking_network_top_uut.all_data_out[416] ),
    .X(_08789_));
 sg13g2_nor2b_1 _16300_ (.A(\spiking_network_top_uut.all_data_out[416] ),
    .B_N(net3796),
    .Y(_08790_));
 sg13g2_a21oi_1 _16301_ (.A1(\spiking_network_top_uut.all_data_out[416] ),
    .A2(net3795),
    .Y(_08791_),
    .B1(_08790_));
 sg13g2_a21oi_1 _16302_ (.A1(\spiking_network_top_uut.all_data_out[417] ),
    .A2(_08789_),
    .Y(_08792_),
    .B1(\spiking_network_top_uut.all_data_out[418] ));
 sg13g2_o21ai_1 _16303_ (.B1(_08792_),
    .Y(_08793_),
    .A1(\spiking_network_top_uut.all_data_out[417] ),
    .A2(_08791_));
 sg13g2_mux2_1 _16304_ (.A0(net3791),
    .A1(net3790),
    .S(\spiking_network_top_uut.all_data_out[416] ),
    .X(_08794_));
 sg13g2_nand2_1 _16305_ (.Y(_08795_),
    .A(\spiking_network_top_uut.all_data_out[417] ),
    .B(_08794_));
 sg13g2_a21oi_1 _16306_ (.A1(\spiking_network_top_uut.all_data_out[416] ),
    .A2(_03658_),
    .Y(_08796_),
    .B1(\spiking_network_top_uut.all_data_out[417] ));
 sg13g2_o21ai_1 _16307_ (.B1(_08796_),
    .Y(_08797_),
    .A1(\spiking_network_top_uut.all_data_out[416] ),
    .A2(net3792));
 sg13g2_nand3_1 _16308_ (.B(_08795_),
    .C(_08797_),
    .A(\spiking_network_top_uut.all_data_out[418] ),
    .Y(_08798_));
 sg13g2_nand3_1 _16309_ (.B(_08793_),
    .C(_08798_),
    .A(net4617),
    .Y(_08799_));
 sg13g2_o21ai_1 _16310_ (.B1(_08799_),
    .Y(_00913_),
    .A1(net4618),
    .A2(_03687_));
 sg13g2_nor3_2 _16311_ (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[2] ),
    .B(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[1] ),
    .C(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[0] ),
    .Y(_08800_));
 sg13g2_nor2b_1 _16312_ (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[3] ),
    .B_N(_08800_),
    .Y(_08801_));
 sg13g2_nor2b_2 _16313_ (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[4] ),
    .B_N(_08801_),
    .Y(_08802_));
 sg13g2_inv_2 _16314_ (.Y(_08803_),
    .A(_08802_));
 sg13g2_o21ai_1 _16315_ (.B1(net4603),
    .Y(_08804_),
    .A1(net3617),
    .A2(_08803_));
 sg13g2_nor2b_1 _16316_ (.A(net3617),
    .B_N(net394),
    .Y(_08805_));
 sg13g2_a21oi_1 _16317_ (.A1(net4284),
    .A2(net3617),
    .Y(_08806_),
    .B1(_08805_));
 sg13g2_nand2_1 _16318_ (.Y(_08807_),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[0] ),
    .B(_08804_));
 sg13g2_o21ai_1 _16319_ (.B1(_08807_),
    .Y(_00914_),
    .A1(_08804_),
    .A2(_08806_));
 sg13g2_xor2_1 _16320_ (.B(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[0] ),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[1] ),
    .X(_08808_));
 sg13g2_nor2_1 _16321_ (.A(net3617),
    .B(_08808_),
    .Y(_08809_));
 sg13g2_a21oi_1 _16322_ (.A1(net4281),
    .A2(net3617),
    .Y(_08810_),
    .B1(_08809_));
 sg13g2_nand2_1 _16323_ (.Y(_08811_),
    .A(net412),
    .B(_08804_));
 sg13g2_o21ai_1 _16324_ (.B1(_08811_),
    .Y(_00915_),
    .A1(_08804_),
    .A2(_08810_));
 sg13g2_o21ai_1 _16325_ (.B1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[2] ),
    .Y(_08812_),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[1] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[0] ));
 sg13g2_nor2b_1 _16326_ (.A(_08800_),
    .B_N(_08812_),
    .Y(_08813_));
 sg13g2_nor2_1 _16327_ (.A(net3617),
    .B(_08813_),
    .Y(_08814_));
 sg13g2_a21oi_1 _16328_ (.A1(net4277),
    .A2(net3617),
    .Y(_08815_),
    .B1(_08814_));
 sg13g2_nand2_1 _16329_ (.Y(_08816_),
    .A(net229),
    .B(_08804_));
 sg13g2_o21ai_1 _16330_ (.B1(_08816_),
    .Y(_00916_),
    .A1(_08804_),
    .A2(_08815_));
 sg13g2_nand2_1 _16331_ (.Y(_08817_),
    .A(net4274),
    .B(net3618));
 sg13g2_xnor2_1 _16332_ (.Y(_08818_),
    .A(net422),
    .B(_08800_));
 sg13g2_o21ai_1 _16333_ (.B1(_08817_),
    .Y(_08819_),
    .A1(net3618),
    .A2(_08818_));
 sg13g2_mux2_1 _16334_ (.A0(_08819_),
    .A1(net422),
    .S(_08804_),
    .X(_00917_));
 sg13g2_nand2_1 _16335_ (.Y(_08820_),
    .A(net3949),
    .B(net258));
 sg13g2_nand2b_1 _16336_ (.Y(_08821_),
    .B(net258),
    .A_N(_08801_));
 sg13g2_a21oi_1 _16337_ (.A1(_08803_),
    .A2(_08821_),
    .Y(_08822_),
    .B1(net3618));
 sg13g2_a21oi_1 _16338_ (.A1(net4269),
    .A2(net3617),
    .Y(_08823_),
    .B1(_08822_));
 sg13g2_o21ai_1 _16339_ (.B1(_08820_),
    .Y(_00918_),
    .A1(_08804_),
    .A2(_08823_));
 sg13g2_mux2_1 _16340_ (.A0(net296),
    .A1(net149),
    .S(net4634),
    .X(_00919_));
 sg13g2_nor2_1 _16341_ (.A(_00109_),
    .B(net3740),
    .Y(_08824_));
 sg13g2_nor2_2 _16342_ (.A(net3748),
    .B(_08824_),
    .Y(_08825_));
 sg13g2_nor2_1 _16343_ (.A(_00109_),
    .B(_08825_),
    .Y(_08826_));
 sg13g2_nand2b_1 _16344_ (.Y(_08827_),
    .B(_08825_),
    .A_N(_00109_));
 sg13g2_o21ai_1 _16345_ (.B1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ),
    .Y(_08828_),
    .A1(_00109_),
    .A2(_08825_));
 sg13g2_inv_1 _16346_ (.Y(_08829_),
    .A(_08828_));
 sg13g2_a21o_1 _16347_ (.A2(net3748),
    .A1(_00110_),
    .B1(_08825_),
    .X(_08830_));
 sg13g2_nor2_1 _16348_ (.A(_00110_),
    .B(net3905),
    .Y(_08831_));
 sg13g2_a221oi_1 _16349_ (.B2(_08824_),
    .C1(_08831_),
    .B1(net3905),
    .A1(_03499_),
    .Y(_08832_),
    .A2(net3748));
 sg13g2_nand2_1 _16350_ (.Y(_08833_),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ),
    .B(_08832_));
 sg13g2_a21oi_1 _16351_ (.A1(net4266),
    .A2(_00110_),
    .Y(_08834_),
    .B1(_05084_));
 sg13g2_a21oi_1 _16352_ (.A1(_03499_),
    .A2(net3738),
    .Y(_08835_),
    .B1(_08834_));
 sg13g2_o21ai_1 _16353_ (.B1(_08835_),
    .Y(_08836_),
    .A1(_00109_),
    .A2(net3910));
 sg13g2_nand2_1 _16354_ (.Y(_08837_),
    .A(_00113_),
    .B(net3748));
 sg13g2_and3_1 _16355_ (.X(_08838_),
    .A(_00112_),
    .B(_08836_),
    .C(_08837_));
 sg13g2_xnor2_1 _16356_ (.Y(_08839_),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ),
    .B(_08832_));
 sg13g2_o21ai_1 _16357_ (.B1(_08833_),
    .Y(_08840_),
    .A1(_08838_),
    .A2(_08839_));
 sg13g2_xnor2_1 _16358_ (.Y(_08841_),
    .A(_03499_),
    .B(_08830_));
 sg13g2_nor2b_1 _16359_ (.A(_08841_),
    .B_N(_08840_),
    .Y(_08842_));
 sg13g2_a21o_1 _16360_ (.A2(_08830_),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ),
    .B1(_08842_),
    .X(_08843_));
 sg13g2_xnor2_1 _16361_ (.Y(_08844_),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ),
    .B(_08826_));
 sg13g2_a21oi_1 _16362_ (.A1(_08843_),
    .A2(_08844_),
    .Y(_08845_),
    .B1(_08829_));
 sg13g2_a22oi_1 _16363_ (.Y(_08846_),
    .B1(_08827_),
    .B2(_08845_),
    .A2(_08825_),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ));
 sg13g2_a21oi_2 _16364_ (.B1(_08846_),
    .Y(_08847_),
    .A2(_00109_),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ));
 sg13g2_nor2_1 _16365_ (.A(_08802_),
    .B(_08847_),
    .Y(_08848_));
 sg13g2_mux2_2 _16366_ (.A0(net4491),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[423] ),
    .X(_08849_));
 sg13g2_nand2_1 _16367_ (.Y(_08850_),
    .A(\spiking_network_top_uut.all_data_out[83] ),
    .B(_08849_));
 sg13g2_mux2_2 _16368_ (.A0(net4492),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[419] ),
    .X(_08851_));
 sg13g2_nand2_1 _16369_ (.Y(_08852_),
    .A(\spiking_network_top_uut.all_data_out[81] ),
    .B(_08851_));
 sg13g2_nor2_1 _16370_ (.A(_08850_),
    .B(_08852_),
    .Y(_08853_));
 sg13g2_nand4_1 _16371_ (.B(\spiking_network_top_uut.all_data_out[80] ),
    .C(_08849_),
    .A(\spiking_network_top_uut.all_data_out[82] ),
    .Y(_08854_),
    .D(_08851_));
 sg13g2_inv_1 _16372_ (.Y(_08855_),
    .A(_08854_));
 sg13g2_xor2_1 _16373_ (.B(_08852_),
    .A(_08850_),
    .X(_08856_));
 sg13g2_a21oi_2 _16374_ (.B1(_08853_),
    .Y(_08857_),
    .A2(_08856_),
    .A1(_08854_));
 sg13g2_mux2_2 _16375_ (.A0(net4490),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[427] ),
    .X(_08858_));
 sg13g2_nand2_2 _16376_ (.Y(_08859_),
    .A(\spiking_network_top_uut.all_data_out[85] ),
    .B(_08858_));
 sg13g2_mux2_2 _16377_ (.A0(net4489),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[431] ),
    .X(_08860_));
 sg13g2_nand2_1 _16378_ (.Y(_08861_),
    .A(\spiking_network_top_uut.all_data_out[87] ),
    .B(_08860_));
 sg13g2_nor2_1 _16379_ (.A(_08859_),
    .B(_08861_),
    .Y(_08862_));
 sg13g2_nand2_2 _16380_ (.Y(_08863_),
    .A(\spiking_network_top_uut.all_data_out[84] ),
    .B(_08858_));
 sg13g2_nand2_1 _16381_ (.Y(_08864_),
    .A(\spiking_network_top_uut.all_data_out[86] ),
    .B(_08860_));
 sg13g2_or2_2 _16382_ (.X(_08865_),
    .B(_08864_),
    .A(_08863_));
 sg13g2_xor2_1 _16383_ (.B(_08861_),
    .A(_08859_),
    .X(_08866_));
 sg13g2_a21oi_2 _16384_ (.B1(_08862_),
    .Y(_08867_),
    .A2(_08866_),
    .A1(_08865_));
 sg13g2_mux2_2 _16385_ (.A0(net4487),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[439] ),
    .X(_08868_));
 sg13g2_mux2_2 _16386_ (.A0(net4488),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[435] ),
    .X(_08869_));
 sg13g2_a22oi_1 _16387_ (.Y(_08870_),
    .B1(_08869_),
    .B2(\spiking_network_top_uut.all_data_out[89] ),
    .A2(_08868_),
    .A1(\spiking_network_top_uut.all_data_out[91] ));
 sg13g2_and4_1 _16388_ (.A(\spiking_network_top_uut.all_data_out[90] ),
    .B(\spiking_network_top_uut.all_data_out[88] ),
    .C(_08868_),
    .D(_08869_),
    .X(_08871_));
 sg13g2_and4_1 _16389_ (.A(\spiking_network_top_uut.all_data_out[91] ),
    .B(\spiking_network_top_uut.all_data_out[89] ),
    .C(_08868_),
    .D(_08869_),
    .X(_08872_));
 sg13g2_nand4_1 _16390_ (.B(\spiking_network_top_uut.all_data_out[89] ),
    .C(_08868_),
    .A(\spiking_network_top_uut.all_data_out[91] ),
    .Y(_08873_),
    .D(_08869_));
 sg13g2_a21oi_2 _16391_ (.B1(_08870_),
    .Y(_08874_),
    .A2(_08873_),
    .A1(_08871_));
 sg13g2_mux2_2 _16392_ (.A0(net4485),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[447] ),
    .X(_08875_));
 sg13g2_mux2_2 _16393_ (.A0(net4486),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[443] ),
    .X(_08876_));
 sg13g2_and4_1 _16394_ (.A(\spiking_network_top_uut.all_data_out[95] ),
    .B(\spiking_network_top_uut.all_data_out[93] ),
    .C(_08875_),
    .D(_08876_),
    .X(_08877_));
 sg13g2_nand4_1 _16395_ (.B(\spiking_network_top_uut.all_data_out[93] ),
    .C(_08875_),
    .A(\spiking_network_top_uut.all_data_out[95] ),
    .Y(_08878_),
    .D(_08876_));
 sg13g2_and4_1 _16396_ (.A(\spiking_network_top_uut.all_data_out[94] ),
    .B(\spiking_network_top_uut.all_data_out[92] ),
    .C(_08875_),
    .D(_08876_),
    .X(_08879_));
 sg13g2_a22oi_1 _16397_ (.Y(_08880_),
    .B1(_08876_),
    .B2(\spiking_network_top_uut.all_data_out[93] ),
    .A2(_08875_),
    .A1(\spiking_network_top_uut.all_data_out[95] ));
 sg13g2_or3_1 _16398_ (.A(_08877_),
    .B(_08879_),
    .C(_08880_),
    .X(_08881_));
 sg13g2_o21ai_1 _16399_ (.B1(_08878_),
    .Y(_08882_),
    .A1(_08879_),
    .A2(_08880_));
 sg13g2_nand3b_1 _16400_ (.B(_08874_),
    .C(_08882_),
    .Y(_08883_),
    .A_N(_08867_));
 sg13g2_inv_1 _16401_ (.Y(_08884_),
    .A(_08883_));
 sg13g2_or2_1 _16402_ (.X(_08885_),
    .B(_08883_),
    .A(_08857_));
 sg13g2_nor2_1 _16403_ (.A(_08874_),
    .B(_08882_),
    .Y(_08886_));
 sg13g2_and2_1 _16404_ (.A(_08867_),
    .B(_08886_),
    .X(_08887_));
 sg13g2_nand2_1 _16405_ (.Y(_08888_),
    .A(_08857_),
    .B(_08887_));
 sg13g2_and2_1 _16406_ (.A(_08885_),
    .B(_08888_),
    .X(_08889_));
 sg13g2_xnor2_1 _16407_ (.Y(_08890_),
    .A(_08827_),
    .B(_08845_));
 sg13g2_nand2_1 _16408_ (.Y(_08891_),
    .A(_08889_),
    .B(_08890_));
 sg13g2_nand2_1 _16409_ (.Y(_08892_),
    .A(_08885_),
    .B(_08891_));
 sg13g2_xor2_1 _16410_ (.B(_08889_),
    .A(_08847_),
    .X(_08893_));
 sg13g2_nand2_1 _16411_ (.Y(_08894_),
    .A(_08892_),
    .B(_08893_));
 sg13g2_xnor2_1 _16412_ (.Y(_08895_),
    .A(_08889_),
    .B(_08890_));
 sg13g2_o21ai_1 _16413_ (.B1(_08879_),
    .Y(_08896_),
    .A1(_08877_),
    .A2(_08880_));
 sg13g2_o21ai_1 _16414_ (.B1(_08871_),
    .Y(_08897_),
    .A1(_08870_),
    .A2(_08872_));
 sg13g2_or3_1 _16415_ (.A(_08870_),
    .B(_08871_),
    .C(_08872_),
    .X(_08898_));
 sg13g2_a22oi_1 _16416_ (.Y(_08899_),
    .B1(_08897_),
    .B2(_08898_),
    .A2(_08896_),
    .A1(_08881_));
 sg13g2_xor2_1 _16417_ (.B(_08866_),
    .A(_08865_),
    .X(_08900_));
 sg13g2_xnor2_1 _16418_ (.Y(_08901_),
    .A(_08865_),
    .B(_08866_));
 sg13g2_and4_1 _16419_ (.A(_08881_),
    .B(_08896_),
    .C(_08897_),
    .D(_08898_),
    .X(_08902_));
 sg13g2_nand4_1 _16420_ (.B(_08896_),
    .C(_08897_),
    .A(_08881_),
    .Y(_08903_),
    .D(_08898_));
 sg13g2_nand3b_1 _16421_ (.B(_08901_),
    .C(_08903_),
    .Y(_08904_),
    .A_N(_08899_));
 sg13g2_a21oi_2 _16422_ (.B1(_08899_),
    .Y(_08905_),
    .A2(_08903_),
    .A1(_08901_));
 sg13g2_xor2_1 _16423_ (.B(_08882_),
    .A(_08874_),
    .X(_08906_));
 sg13g2_xnor2_1 _16424_ (.Y(_08907_),
    .A(_08867_),
    .B(_08906_));
 sg13g2_nand2b_1 _16425_ (.Y(_08908_),
    .B(_08907_),
    .A_N(_08905_));
 sg13g2_xnor2_1 _16426_ (.Y(_08909_),
    .A(_08905_),
    .B(_08907_));
 sg13g2_nand2b_1 _16427_ (.Y(_08910_),
    .B(_08909_),
    .A_N(_08857_));
 sg13g2_nand2_1 _16428_ (.Y(_08911_),
    .A(_08908_),
    .B(_08910_));
 sg13g2_nor2_1 _16429_ (.A(_08884_),
    .B(_08887_),
    .Y(_08912_));
 sg13g2_xnor2_1 _16430_ (.Y(_08913_),
    .A(_08857_),
    .B(_08912_));
 sg13g2_and2_1 _16431_ (.A(_08911_),
    .B(_08913_),
    .X(_08914_));
 sg13g2_xor2_1 _16432_ (.B(_08913_),
    .A(_08911_),
    .X(_08915_));
 sg13g2_xnor2_1 _16433_ (.Y(_08916_),
    .A(_08843_),
    .B(_08844_));
 sg13g2_inv_1 _16434_ (.Y(_08917_),
    .A(_08916_));
 sg13g2_a21oi_1 _16435_ (.A1(_08915_),
    .A2(_08917_),
    .Y(_08918_),
    .B1(_08914_));
 sg13g2_nor2_1 _16436_ (.A(_08895_),
    .B(_08918_),
    .Y(_08919_));
 sg13g2_a22oi_1 _16437_ (.Y(_08920_),
    .B1(_08876_),
    .B2(\spiking_network_top_uut.all_data_out[92] ),
    .A2(_08875_),
    .A1(\spiking_network_top_uut.all_data_out[94] ));
 sg13g2_nor2_2 _16438_ (.A(_08879_),
    .B(_08920_),
    .Y(_08921_));
 sg13g2_a22oi_1 _16439_ (.Y(_08922_),
    .B1(_08869_),
    .B2(\spiking_network_top_uut.all_data_out[88] ),
    .A2(_08868_),
    .A1(\spiking_network_top_uut.all_data_out[90] ));
 sg13g2_nor2_1 _16440_ (.A(_08871_),
    .B(_08922_),
    .Y(_08923_));
 sg13g2_and2_1 _16441_ (.A(_08921_),
    .B(_08923_),
    .X(_08924_));
 sg13g2_xor2_1 _16442_ (.B(_08864_),
    .A(_08863_),
    .X(_08925_));
 sg13g2_xor2_1 _16443_ (.B(_08923_),
    .A(_08921_),
    .X(_08926_));
 sg13g2_a21o_1 _16444_ (.A2(_08926_),
    .A1(_08925_),
    .B1(_08924_),
    .X(_08927_));
 sg13g2_o21ai_1 _16445_ (.B1(_08900_),
    .Y(_08928_),
    .A1(_08899_),
    .A2(_08902_));
 sg13g2_nand3_1 _16446_ (.B(_08927_),
    .C(_08928_),
    .A(_08904_),
    .Y(_08929_));
 sg13g2_xnor2_1 _16447_ (.Y(_08930_),
    .A(_08855_),
    .B(_08856_));
 sg13g2_inv_1 _16448_ (.Y(_08931_),
    .A(_08930_));
 sg13g2_a21oi_1 _16449_ (.A1(_08904_),
    .A2(_08928_),
    .Y(_08932_),
    .B1(_08927_));
 sg13g2_a21o_1 _16450_ (.A2(_08928_),
    .A1(_08904_),
    .B1(_08927_),
    .X(_08933_));
 sg13g2_nand3_1 _16451_ (.B(_08931_),
    .C(_08933_),
    .A(_08929_),
    .Y(_08934_));
 sg13g2_o21ai_1 _16452_ (.B1(_08929_),
    .Y(_08935_),
    .A1(_08930_),
    .A2(_08932_));
 sg13g2_xnor2_1 _16453_ (.Y(_08936_),
    .A(_08857_),
    .B(_08909_));
 sg13g2_nand2_1 _16454_ (.Y(_08937_),
    .A(_08935_),
    .B(_08936_));
 sg13g2_xnor2_1 _16455_ (.Y(_08938_),
    .A(_08935_),
    .B(_08936_));
 sg13g2_xor2_1 _16456_ (.B(_08841_),
    .A(_08840_),
    .X(_08939_));
 sg13g2_o21ai_1 _16457_ (.B1(_08937_),
    .Y(_08940_),
    .A1(_08938_),
    .A2(_08939_));
 sg13g2_xnor2_1 _16458_ (.Y(_08941_),
    .A(_08915_),
    .B(_08916_));
 sg13g2_nand2_1 _16459_ (.Y(_08942_),
    .A(_08940_),
    .B(_08941_));
 sg13g2_xor2_1 _16460_ (.B(_08939_),
    .A(_08938_),
    .X(_08943_));
 sg13g2_a22oi_1 _16461_ (.Y(_08944_),
    .B1(_08851_),
    .B2(\spiking_network_top_uut.all_data_out[80] ),
    .A2(_08849_),
    .A1(\spiking_network_top_uut.all_data_out[82] ));
 sg13g2_xnor2_1 _16462_ (.Y(_08945_),
    .A(_08925_),
    .B(_08926_));
 sg13g2_or3_2 _16463_ (.A(_08855_),
    .B(_08944_),
    .C(_08945_),
    .X(_08946_));
 sg13g2_inv_1 _16464_ (.Y(_08947_),
    .A(_08946_));
 sg13g2_a21o_2 _16465_ (.A2(_08933_),
    .A1(_08929_),
    .B1(_08931_),
    .X(_08948_));
 sg13g2_nand3_1 _16466_ (.B(_08947_),
    .C(_08948_),
    .A(_08934_),
    .Y(_08949_));
 sg13g2_a21oi_2 _16467_ (.B1(_08947_),
    .Y(_08950_),
    .A2(_08948_),
    .A1(_08934_));
 sg13g2_a21o_2 _16468_ (.A2(_08948_),
    .A1(_08934_),
    .B1(_08947_),
    .X(_08951_));
 sg13g2_xnor2_1 _16469_ (.Y(_08952_),
    .A(_08838_),
    .B(_08839_));
 sg13g2_inv_1 _16470_ (.Y(_08953_),
    .A(_08952_));
 sg13g2_and3_1 _16471_ (.X(_08954_),
    .A(_08949_),
    .B(_08951_),
    .C(_08953_));
 sg13g2_o21ai_1 _16472_ (.B1(_08949_),
    .Y(_08955_),
    .A1(_08950_),
    .A2(_08952_));
 sg13g2_and2_1 _16473_ (.A(_08943_),
    .B(_08955_),
    .X(_08956_));
 sg13g2_a21oi_1 _16474_ (.A1(_08949_),
    .A2(_08951_),
    .Y(_08957_),
    .B1(_08953_));
 sg13g2_nor2_1 _16475_ (.A(_08954_),
    .B(_08957_),
    .Y(_08958_));
 sg13g2_o21ai_1 _16476_ (.B1(_08945_),
    .Y(_08959_),
    .A1(_08855_),
    .A2(_08944_));
 sg13g2_and2_2 _16477_ (.A(_08946_),
    .B(_08959_),
    .X(_08960_));
 sg13g2_a21oi_1 _16478_ (.A1(_08836_),
    .A2(_08837_),
    .Y(_08961_),
    .B1(_00112_));
 sg13g2_or2_1 _16479_ (.X(_08962_),
    .B(_08961_),
    .A(_08838_));
 sg13g2_nand2_1 _16480_ (.Y(_08963_),
    .A(_08960_),
    .B(_08962_));
 sg13g2_nor3_2 _16481_ (.A(_08954_),
    .B(_08957_),
    .C(_08963_),
    .Y(_08964_));
 sg13g2_xor2_1 _16482_ (.B(_08955_),
    .A(_08943_),
    .X(_08965_));
 sg13g2_a21oi_2 _16483_ (.B1(_08956_),
    .Y(_08966_),
    .A2(_08965_),
    .A1(_08964_));
 sg13g2_xnor2_1 _16484_ (.Y(_08967_),
    .A(_08940_),
    .B(_08941_));
 sg13g2_or2_1 _16485_ (.X(_08968_),
    .B(_08967_),
    .A(_08966_));
 sg13g2_o21ai_1 _16486_ (.B1(_08942_),
    .Y(_08969_),
    .A1(_08966_),
    .A2(_08967_));
 sg13g2_nand2_1 _16487_ (.Y(_08970_),
    .A(_08895_),
    .B(_08918_));
 sg13g2_nand2b_1 _16488_ (.Y(_08971_),
    .B(_08970_),
    .A_N(_08919_));
 sg13g2_a21oi_1 _16489_ (.A1(_08969_),
    .A2(_08970_),
    .Y(_08972_),
    .B1(_08919_));
 sg13g2_xnor2_1 _16490_ (.Y(_08973_),
    .A(_08892_),
    .B(_08893_));
 sg13g2_o21ai_1 _16491_ (.B1(_08894_),
    .Y(_08974_),
    .A1(_08972_),
    .A2(_08973_));
 sg13g2_mux2_1 _16492_ (.A0(_08888_),
    .A1(_08885_),
    .S(_08847_),
    .X(_08975_));
 sg13g2_xnor2_1 _16493_ (.Y(_08976_),
    .A(_08974_),
    .B(_08975_));
 sg13g2_a21oi_2 _16494_ (.B1(_08848_),
    .Y(_08977_),
    .A2(_08976_),
    .A1(_08802_));
 sg13g2_xnor2_1 _16495_ (.Y(_08978_),
    .A(_08972_),
    .B(_08973_));
 sg13g2_a21oi_1 _16496_ (.A1(_08802_),
    .A2(_08978_),
    .Y(_08979_),
    .B1(_08848_));
 sg13g2_xnor2_1 _16497_ (.Y(_08980_),
    .A(_08969_),
    .B(_08971_));
 sg13g2_mux2_1 _16498_ (.A0(_08890_),
    .A1(_08980_),
    .S(_08802_),
    .X(_08981_));
 sg13g2_nand2_1 _16499_ (.Y(_08982_),
    .A(_08979_),
    .B(_08981_));
 sg13g2_a21oi_2 _16500_ (.B1(net3619),
    .Y(_08983_),
    .A2(_08982_),
    .A1(_08977_));
 sg13g2_nor2_1 _16501_ (.A(_08979_),
    .B(_08981_),
    .Y(_08984_));
 sg13g2_nor2_2 _16502_ (.A(_08977_),
    .B(_08984_),
    .Y(_08985_));
 sg13g2_nand2_1 _16503_ (.Y(_08986_),
    .A(_08802_),
    .B(_08960_));
 sg13g2_xnor2_1 _16504_ (.Y(_08987_),
    .A(_08962_),
    .B(_08986_));
 sg13g2_o21ai_1 _16505_ (.B1(_08983_),
    .Y(_08988_),
    .A1(_08985_),
    .A2(_08987_));
 sg13g2_xor2_1 _16506_ (.B(net445),
    .A(net4313),
    .X(_08989_));
 sg13g2_a21oi_1 _16507_ (.A1(net3619),
    .A2(_08989_),
    .Y(_08990_),
    .B1(net3951));
 sg13g2_a22oi_1 _16508_ (.Y(_00920_),
    .B1(_08988_),
    .B2(_08990_),
    .A2(_03453_),
    .A1(net3950));
 sg13g2_nor2b_1 _16509_ (.A(_08958_),
    .B_N(_08963_),
    .Y(_08991_));
 sg13g2_or3_1 _16510_ (.A(_08803_),
    .B(_08964_),
    .C(_08991_),
    .X(_08992_));
 sg13g2_o21ai_1 _16511_ (.B1(_08992_),
    .Y(_08993_),
    .A1(_08802_),
    .A2(_08952_));
 sg13g2_o21ai_1 _16512_ (.B1(_08983_),
    .Y(_08994_),
    .A1(_08985_),
    .A2(_08993_));
 sg13g2_xor2_1 _16513_ (.B(_04901_),
    .A(_04900_),
    .X(_08995_));
 sg13g2_a21oi_1 _16514_ (.A1(net3619),
    .A2(_08995_),
    .Y(_08996_),
    .B1(net3951));
 sg13g2_a22oi_1 _16515_ (.Y(_00921_),
    .B1(_08994_),
    .B2(_08996_),
    .A2(_03452_),
    .A1(net3950));
 sg13g2_xnor2_1 _16516_ (.Y(_08997_),
    .A(_08964_),
    .B(_08965_));
 sg13g2_nand2b_1 _16517_ (.Y(_08998_),
    .B(_08803_),
    .A_N(_08939_));
 sg13g2_o21ai_1 _16518_ (.B1(_08998_),
    .Y(_08999_),
    .A1(_08803_),
    .A2(_08997_));
 sg13g2_o21ai_1 _16519_ (.B1(_08983_),
    .Y(_09000_),
    .A1(_08985_),
    .A2(_08999_));
 sg13g2_xnor2_1 _16520_ (.Y(_09001_),
    .A(_04898_),
    .B(_04902_));
 sg13g2_a21oi_1 _16521_ (.A1(net3619),
    .A2(_09001_),
    .Y(_09002_),
    .B1(net3950));
 sg13g2_a22oi_1 _16522_ (.Y(_00922_),
    .B1(_09000_),
    .B2(_09002_),
    .A2(_03451_),
    .A1(net3950));
 sg13g2_nand2_1 _16523_ (.Y(_09003_),
    .A(_08966_),
    .B(_08967_));
 sg13g2_a21oi_1 _16524_ (.A1(_08968_),
    .A2(_09003_),
    .Y(_09004_),
    .B1(_08803_));
 sg13g2_a21oi_1 _16525_ (.A1(_08803_),
    .A2(_08916_),
    .Y(_09005_),
    .B1(_09004_));
 sg13g2_o21ai_1 _16526_ (.B1(_08983_),
    .Y(_09006_),
    .A1(_08985_),
    .A2(_09005_));
 sg13g2_or3_1 _16527_ (.A(_04896_),
    .B(_04897_),
    .C(_04903_),
    .X(_09007_));
 sg13g2_and2_1 _16528_ (.A(_04904_),
    .B(_09007_),
    .X(_09008_));
 sg13g2_a21oi_1 _16529_ (.A1(net3619),
    .A2(_09008_),
    .Y(_09009_),
    .B1(net3950));
 sg13g2_a22oi_1 _16530_ (.Y(_00923_),
    .B1(_09006_),
    .B2(_09009_),
    .A2(_03450_),
    .A1(net3950));
 sg13g2_nand2b_1 _16531_ (.Y(_09010_),
    .B(_08977_),
    .A_N(net3619));
 sg13g2_a21oi_1 _16532_ (.A1(_04895_),
    .A2(_04905_),
    .Y(_09011_),
    .B1(net3950));
 sg13g2_a22oi_1 _16533_ (.Y(_00924_),
    .B1(_09010_),
    .B2(_09011_),
    .A2(_03449_),
    .A1(net3950));
 sg13g2_mux2_1 _16534_ (.A0(net3787),
    .A1(net3786),
    .S(\spiking_network_top_uut.all_data_out[476] ),
    .X(_09012_));
 sg13g2_nor2b_1 _16535_ (.A(\spiking_network_top_uut.all_data_out[476] ),
    .B_N(net3789),
    .Y(_09013_));
 sg13g2_a21oi_1 _16536_ (.A1(\spiking_network_top_uut.all_data_out[476] ),
    .A2(net3788),
    .Y(_09014_),
    .B1(_09013_));
 sg13g2_a21oi_1 _16537_ (.A1(\spiking_network_top_uut.all_data_out[477] ),
    .A2(_09012_),
    .Y(_09015_),
    .B1(\spiking_network_top_uut.all_data_out[478] ));
 sg13g2_o21ai_1 _16538_ (.B1(_09015_),
    .Y(_09016_),
    .A1(\spiking_network_top_uut.all_data_out[477] ),
    .A2(_09014_));
 sg13g2_mux2_1 _16539_ (.A0(net3783),
    .A1(net3899),
    .S(\spiking_network_top_uut.all_data_out[476] ),
    .X(_09017_));
 sg13g2_nor2b_1 _16540_ (.A(\spiking_network_top_uut.all_data_out[476] ),
    .B_N(net3785),
    .Y(_09018_));
 sg13g2_a21oi_1 _16541_ (.A1(\spiking_network_top_uut.all_data_out[476] ),
    .A2(net3784),
    .Y(_09019_),
    .B1(_09018_));
 sg13g2_o21ai_1 _16542_ (.B1(\spiking_network_top_uut.all_data_out[478] ),
    .Y(_09020_),
    .A1(\spiking_network_top_uut.all_data_out[477] ),
    .A2(_09019_));
 sg13g2_a21oi_1 _16543_ (.A1(\spiking_network_top_uut.all_data_out[477] ),
    .A2(_09017_),
    .Y(_09021_),
    .B1(_09020_));
 sg13g2_nand2_1 _16544_ (.Y(_09022_),
    .A(net4638),
    .B(_09016_));
 sg13g2_nand2_1 _16545_ (.Y(_09023_),
    .A(net3962),
    .B(net240));
 sg13g2_o21ai_1 _16546_ (.B1(_09023_),
    .Y(_00925_),
    .A1(_09021_),
    .A2(_09022_));
 sg13g2_mux2_1 _16547_ (.A0(net444),
    .A1(net240),
    .S(net4639),
    .X(_00926_));
 sg13g2_mux4_1 _16548_ (.S0(\spiking_network_top_uut.all_data_out[472] ),
    .A0(net3840),
    .A1(net3839),
    .A2(net3838),
    .A3(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[3] ),
    .S1(\spiking_network_top_uut.all_data_out[473] ),
    .X(_09024_));
 sg13g2_mux2_1 _16549_ (.A0(net3835),
    .A1(net3834),
    .S(\spiking_network_top_uut.all_data_out[472] ),
    .X(_09025_));
 sg13g2_nor2b_1 _16550_ (.A(\spiking_network_top_uut.all_data_out[472] ),
    .B_N(net3836),
    .Y(_09026_));
 sg13g2_a21oi_1 _16551_ (.A1(\spiking_network_top_uut.all_data_out[472] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[5] ),
    .Y(_09027_),
    .B1(_09026_));
 sg13g2_o21ai_1 _16552_ (.B1(\spiking_network_top_uut.all_data_out[474] ),
    .Y(_09028_),
    .A1(\spiking_network_top_uut.all_data_out[473] ),
    .A2(_09027_));
 sg13g2_a21oi_1 _16553_ (.A1(\spiking_network_top_uut.all_data_out[473] ),
    .A2(_09025_),
    .Y(_09029_),
    .B1(_09028_));
 sg13g2_o21ai_1 _16554_ (.B1(net4641),
    .Y(_09030_),
    .A1(\spiking_network_top_uut.all_data_out[474] ),
    .A2(_09024_));
 sg13g2_nand2_1 _16555_ (.Y(_09031_),
    .A(net3963),
    .B(net141));
 sg13g2_o21ai_1 _16556_ (.B1(_09031_),
    .Y(_00927_),
    .A1(_09029_),
    .A2(_09030_));
 sg13g2_mux2_1 _16557_ (.A0(net241),
    .A1(net141),
    .S(net4640),
    .X(_00928_));
 sg13g2_a21oi_1 _16558_ (.A1(\spiking_network_top_uut.all_data_out[468] ),
    .A2(_03661_),
    .Y(_09032_),
    .B1(\spiking_network_top_uut.all_data_out[469] ));
 sg13g2_o21ai_1 _16559_ (.B1(_09032_),
    .Y(_09033_),
    .A1(\spiking_network_top_uut.all_data_out[468] ),
    .A2(net3829));
 sg13g2_mux2_1 _16560_ (.A0(net3828),
    .A1(net3827),
    .S(\spiking_network_top_uut.all_data_out[468] ),
    .X(_09034_));
 sg13g2_nand2_1 _16561_ (.Y(_09035_),
    .A(\spiking_network_top_uut.all_data_out[469] ),
    .B(_09034_));
 sg13g2_nand3_1 _16562_ (.B(_09033_),
    .C(_09035_),
    .A(\spiking_network_top_uut.all_data_out[470] ),
    .Y(_09036_));
 sg13g2_mux2_1 _16563_ (.A0(net3831),
    .A1(net3830),
    .S(\spiking_network_top_uut.all_data_out[468] ),
    .X(_09037_));
 sg13g2_nor2b_1 _16564_ (.A(\spiking_network_top_uut.all_data_out[468] ),
    .B_N(net3833),
    .Y(_09038_));
 sg13g2_a21oi_1 _16565_ (.A1(\spiking_network_top_uut.all_data_out[468] ),
    .A2(net3832),
    .Y(_09039_),
    .B1(_09038_));
 sg13g2_a21oi_1 _16566_ (.A1(\spiking_network_top_uut.all_data_out[469] ),
    .A2(_09037_),
    .Y(_09040_),
    .B1(\spiking_network_top_uut.all_data_out[470] ));
 sg13g2_o21ai_1 _16567_ (.B1(_09040_),
    .Y(_09041_),
    .A1(\spiking_network_top_uut.all_data_out[469] ),
    .A2(_09039_));
 sg13g2_nand3_1 _16568_ (.B(_09036_),
    .C(_09041_),
    .A(net4607),
    .Y(_09042_));
 sg13g2_o21ai_1 _16569_ (.B1(_09042_),
    .Y(_00929_),
    .A1(net4608),
    .A2(_03688_));
 sg13g2_nor2_1 _16570_ (.A(net4612),
    .B(net55),
    .Y(_09043_));
 sg13g2_a21oi_1 _16571_ (.A1(net4612),
    .A2(_03688_),
    .Y(_00930_),
    .B1(_09043_));
 sg13g2_nand2_1 _16572_ (.Y(_09044_),
    .A(\spiking_network_top_uut.all_data_out[464] ),
    .B(_03660_));
 sg13g2_nor2_1 _16573_ (.A(\spiking_network_top_uut.all_data_out[464] ),
    .B(net3822),
    .Y(_09045_));
 sg13g2_nor2_1 _16574_ (.A(\spiking_network_top_uut.all_data_out[465] ),
    .B(_09045_),
    .Y(_09046_));
 sg13g2_mux2_1 _16575_ (.A0(net3821),
    .A1(net3820),
    .S(\spiking_network_top_uut.all_data_out[464] ),
    .X(_09047_));
 sg13g2_a221oi_1 _16576_ (.B2(\spiking_network_top_uut.all_data_out[465] ),
    .C1(_03621_),
    .B1(_09047_),
    .A1(_09044_),
    .Y(_09048_),
    .A2(_09046_));
 sg13g2_mux4_1 _16577_ (.S0(\spiking_network_top_uut.all_data_out[464] ),
    .A0(net3826),
    .A1(net3825),
    .A2(net3824),
    .A3(net3823),
    .S1(\spiking_network_top_uut.all_data_out[465] ),
    .X(_09049_));
 sg13g2_o21ai_1 _16578_ (.B1(net4614),
    .Y(_09050_),
    .A1(\spiking_network_top_uut.all_data_out[466] ),
    .A2(_09049_));
 sg13g2_nand2_1 _16579_ (.Y(_09051_),
    .A(net3965),
    .B(net172));
 sg13g2_o21ai_1 _16580_ (.B1(_09051_),
    .Y(_00931_),
    .A1(_09048_),
    .A2(_09050_));
 sg13g2_mux2_1 _16581_ (.A0(net290),
    .A1(net172),
    .S(net4620),
    .X(_00932_));
 sg13g2_mux4_1 _16582_ (.S0(\spiking_network_top_uut.all_data_out[460] ),
    .A0(net3819),
    .A1(net3818),
    .A2(net3817),
    .A3(net3816),
    .S1(\spiking_network_top_uut.all_data_out[461] ),
    .X(_09052_));
 sg13g2_mux2_1 _16583_ (.A0(net3814),
    .A1(net3813),
    .S(\spiking_network_top_uut.all_data_out[460] ),
    .X(_09053_));
 sg13g2_nor2b_1 _16584_ (.A(\spiking_network_top_uut.all_data_out[460] ),
    .B_N(net3815),
    .Y(_09054_));
 sg13g2_a21oi_1 _16585_ (.A1(\spiking_network_top_uut.all_data_out[460] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[5] ),
    .Y(_09055_),
    .B1(_09054_));
 sg13g2_o21ai_1 _16586_ (.B1(\spiking_network_top_uut.all_data_out[462] ),
    .Y(_09056_),
    .A1(\spiking_network_top_uut.all_data_out[461] ),
    .A2(_09055_));
 sg13g2_a21oi_1 _16587_ (.A1(\spiking_network_top_uut.all_data_out[461] ),
    .A2(_09053_),
    .Y(_09057_),
    .B1(_09056_));
 sg13g2_o21ai_1 _16588_ (.B1(net4626),
    .Y(_09058_),
    .A1(\spiking_network_top_uut.all_data_out[462] ),
    .A2(_09052_));
 sg13g2_nand2_1 _16589_ (.Y(_09059_),
    .A(net3960),
    .B(net109));
 sg13g2_o21ai_1 _16590_ (.B1(_09059_),
    .Y(_00933_),
    .A1(_09057_),
    .A2(_09058_));
 sg13g2_mux2_1 _16591_ (.A0(net185),
    .A1(net109),
    .S(net4626),
    .X(_00934_));
 sg13g2_mux2_1 _16592_ (.A0(net3810),
    .A1(net3809),
    .S(\spiking_network_top_uut.all_data_out[456] ),
    .X(_09060_));
 sg13g2_nor2b_1 _16593_ (.A(\spiking_network_top_uut.all_data_out[456] ),
    .B_N(net3812),
    .Y(_09061_));
 sg13g2_a21oi_1 _16594_ (.A1(\spiking_network_top_uut.all_data_out[456] ),
    .A2(net3811),
    .Y(_09062_),
    .B1(_09061_));
 sg13g2_a21oi_1 _16595_ (.A1(\spiking_network_top_uut.all_data_out[457] ),
    .A2(_09060_),
    .Y(_09063_),
    .B1(\spiking_network_top_uut.all_data_out[458] ));
 sg13g2_o21ai_1 _16596_ (.B1(_09063_),
    .Y(_09064_),
    .A1(\spiking_network_top_uut.all_data_out[457] ),
    .A2(_09062_));
 sg13g2_mux2_1 _16597_ (.A0(net3806),
    .A1(net3805),
    .S(\spiking_network_top_uut.all_data_out[456] ),
    .X(_09065_));
 sg13g2_nor2b_1 _16598_ (.A(\spiking_network_top_uut.all_data_out[456] ),
    .B_N(net3808),
    .Y(_09066_));
 sg13g2_a21oi_1 _16599_ (.A1(\spiking_network_top_uut.all_data_out[456] ),
    .A2(net3807),
    .Y(_09067_),
    .B1(_09066_));
 sg13g2_o21ai_1 _16600_ (.B1(\spiking_network_top_uut.all_data_out[458] ),
    .Y(_09068_),
    .A1(\spiking_network_top_uut.all_data_out[457] ),
    .A2(_09067_));
 sg13g2_a21oi_1 _16601_ (.A1(\spiking_network_top_uut.all_data_out[457] ),
    .A2(_09065_),
    .Y(_09069_),
    .B1(_09068_));
 sg13g2_nand2_1 _16602_ (.Y(_09070_),
    .A(net4622),
    .B(_09064_));
 sg13g2_nand2_1 _16603_ (.Y(_09071_),
    .A(net3959),
    .B(net96));
 sg13g2_o21ai_1 _16604_ (.B1(_09071_),
    .Y(_00935_),
    .A1(_09069_),
    .A2(_09070_));
 sg13g2_mux2_1 _16605_ (.A0(net310),
    .A1(net96),
    .S(net4621),
    .X(_00936_));
 sg13g2_mux4_1 _16606_ (.S0(\spiking_network_top_uut.all_data_out[452] ),
    .A0(net3804),
    .A1(net3803),
    .A2(net3802),
    .A3(net3801),
    .S1(\spiking_network_top_uut.all_data_out[453] ),
    .X(_09072_));
 sg13g2_mux2_1 _16607_ (.A0(net3798),
    .A1(net3797),
    .S(\spiking_network_top_uut.all_data_out[452] ),
    .X(_09073_));
 sg13g2_nor2b_1 _16608_ (.A(\spiking_network_top_uut.all_data_out[452] ),
    .B_N(net3800),
    .Y(_09074_));
 sg13g2_a21oi_1 _16609_ (.A1(\spiking_network_top_uut.all_data_out[452] ),
    .A2(net3799),
    .Y(_09075_),
    .B1(_09074_));
 sg13g2_o21ai_1 _16610_ (.B1(\spiking_network_top_uut.all_data_out[454] ),
    .Y(_09076_),
    .A1(\spiking_network_top_uut.all_data_out[453] ),
    .A2(_09075_));
 sg13g2_a21oi_1 _16611_ (.A1(\spiking_network_top_uut.all_data_out[453] ),
    .A2(_09073_),
    .Y(_09077_),
    .B1(_09076_));
 sg13g2_o21ai_1 _16612_ (.B1(net4632),
    .Y(_09078_),
    .A1(\spiking_network_top_uut.all_data_out[454] ),
    .A2(_09072_));
 sg13g2_nand2_1 _16613_ (.Y(_09079_),
    .A(net3961),
    .B(net151));
 sg13g2_o21ai_1 _16614_ (.B1(_09079_),
    .Y(_00937_),
    .A1(_09077_),
    .A2(_09078_));
 sg13g2_mux2_1 _16615_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_dout ),
    .A1(net151),
    .S(net4635),
    .X(_00938_));
 sg13g2_nand2_1 _16616_ (.Y(_09080_),
    .A(\spiking_network_top_uut.all_data_out[448] ),
    .B(_03658_));
 sg13g2_nor2_1 _16617_ (.A(\spiking_network_top_uut.all_data_out[448] ),
    .B(net3792),
    .Y(_09081_));
 sg13g2_nor2_1 _16618_ (.A(\spiking_network_top_uut.all_data_out[449] ),
    .B(_09081_),
    .Y(_09082_));
 sg13g2_mux2_1 _16619_ (.A0(net3791),
    .A1(net3790),
    .S(\spiking_network_top_uut.all_data_out[448] ),
    .X(_09083_));
 sg13g2_a221oi_1 _16620_ (.B2(\spiking_network_top_uut.all_data_out[449] ),
    .C1(_03623_),
    .B1(_09083_),
    .A1(_09080_),
    .Y(_09084_),
    .A2(_09082_));
 sg13g2_mux4_1 _16621_ (.S0(\spiking_network_top_uut.all_data_out[448] ),
    .A0(net3796),
    .A1(net3795),
    .A2(net3794),
    .A3(net3793),
    .S1(\spiking_network_top_uut.all_data_out[449] ),
    .X(_02059_));
 sg13g2_o21ai_1 _16622_ (.B1(net4617),
    .Y(_02060_),
    .A1(\spiking_network_top_uut.all_data_out[450] ),
    .A2(_02059_));
 sg13g2_nand2_1 _16623_ (.Y(_02061_),
    .A(net3965),
    .B(net217));
 sg13g2_o21ai_1 _16624_ (.B1(_02061_),
    .Y(_00939_),
    .A1(_09084_),
    .A2(_02060_));
 sg13g2_nor3_2 _16625_ (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[2] ),
    .B(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[1] ),
    .C(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[0] ),
    .Y(_02062_));
 sg13g2_nor2b_1 _16626_ (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[3] ),
    .B_N(_02062_),
    .Y(_02063_));
 sg13g2_nor2b_2 _16627_ (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[4] ),
    .B_N(_02063_),
    .Y(_02064_));
 sg13g2_nand2b_1 _16628_ (.Y(_02065_),
    .B(_02063_),
    .A_N(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[4] ));
 sg13g2_o21ai_1 _16629_ (.B1(net4606),
    .Y(_02066_),
    .A1(net3643),
    .A2(_02065_));
 sg13g2_nor2b_1 _16630_ (.A(net3643),
    .B_N(_00120_),
    .Y(_02067_));
 sg13g2_a21oi_1 _16631_ (.A1(net4286),
    .A2(net3644),
    .Y(_02068_),
    .B1(_02067_));
 sg13g2_nand2_1 _16632_ (.Y(_02069_),
    .A(net329),
    .B(_02066_));
 sg13g2_o21ai_1 _16633_ (.B1(_02069_),
    .Y(_00940_),
    .A1(_02066_),
    .A2(_02068_));
 sg13g2_xor2_1 _16634_ (.B(net329),
    .A(net342),
    .X(_02070_));
 sg13g2_nor2_1 _16635_ (.A(net3644),
    .B(_02070_),
    .Y(_02071_));
 sg13g2_a21oi_1 _16636_ (.A1(net4282),
    .A2(net3644),
    .Y(_02072_),
    .B1(_02071_));
 sg13g2_nand2_1 _16637_ (.Y(_02073_),
    .A(net342),
    .B(_02066_));
 sg13g2_o21ai_1 _16638_ (.B1(_02073_),
    .Y(_00941_),
    .A1(_02066_),
    .A2(_02072_));
 sg13g2_o21ai_1 _16639_ (.B1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[2] ),
    .Y(_02074_),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[1] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[0] ));
 sg13g2_nor2b_1 _16640_ (.A(_02062_),
    .B_N(_02074_),
    .Y(_02075_));
 sg13g2_nor2_1 _16641_ (.A(net3643),
    .B(_02075_),
    .Y(_02076_));
 sg13g2_a21oi_1 _16642_ (.A1(net4279),
    .A2(net3643),
    .Y(_02077_),
    .B1(_02076_));
 sg13g2_nand2_1 _16643_ (.Y(_02078_),
    .A(net206),
    .B(_02066_));
 sg13g2_o21ai_1 _16644_ (.B1(_02078_),
    .Y(_00942_),
    .A1(_02066_),
    .A2(_02077_));
 sg13g2_nand2_1 _16645_ (.Y(_02079_),
    .A(net4275),
    .B(net3643));
 sg13g2_xnor2_1 _16646_ (.Y(_02080_),
    .A(net421),
    .B(_02062_));
 sg13g2_o21ai_1 _16647_ (.B1(_02079_),
    .Y(_02081_),
    .A1(net3643),
    .A2(_02080_));
 sg13g2_mux2_1 _16648_ (.A0(_02081_),
    .A1(net421),
    .S(_02066_),
    .X(_00943_));
 sg13g2_nand2_1 _16649_ (.Y(_02082_),
    .A(net3958),
    .B(net348));
 sg13g2_nand2b_1 _16650_ (.Y(_02083_),
    .B(net348),
    .A_N(_02063_));
 sg13g2_a21oi_1 _16651_ (.A1(net3701),
    .A2(_02083_),
    .Y(_02084_),
    .B1(net3643));
 sg13g2_a21oi_1 _16652_ (.A1(net4272),
    .A2(net3643),
    .Y(_02085_),
    .B1(_02084_));
 sg13g2_o21ai_1 _16653_ (.B1(_02082_),
    .Y(_00944_),
    .A1(_02066_),
    .A2(_02085_));
 sg13g2_mux2_1 _16654_ (.A0(net221),
    .A1(net217),
    .S(net4619),
    .X(_00945_));
 sg13g2_a21oi_1 _16655_ (.A1(net3915),
    .A2(net3912),
    .Y(_02086_),
    .B1(_00115_));
 sg13g2_nor2_2 _16656_ (.A(net3753),
    .B(_02086_),
    .Y(_02087_));
 sg13g2_nor2_1 _16657_ (.A(_00115_),
    .B(_02087_),
    .Y(_02088_));
 sg13g2_nand2b_1 _16658_ (.Y(_02089_),
    .B(_02087_),
    .A_N(_00115_));
 sg13g2_o21ai_1 _16659_ (.B1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ),
    .Y(_02090_),
    .A1(_00115_),
    .A2(_02087_));
 sg13g2_inv_1 _16660_ (.Y(_02091_),
    .A(_02090_));
 sg13g2_a21o_1 _16661_ (.A2(net3753),
    .A1(_00116_),
    .B1(_02087_),
    .X(_02092_));
 sg13g2_nor2_1 _16662_ (.A(_00116_),
    .B(net3908),
    .Y(_02093_));
 sg13g2_a221oi_1 _16663_ (.B2(_02086_),
    .C1(_02093_),
    .B1(net3908),
    .A1(_03500_),
    .Y(_02094_),
    .A2(net3753));
 sg13g2_nand2_1 _16664_ (.Y(_02095_),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ),
    .B(_02094_));
 sg13g2_nor2_1 _16665_ (.A(_00115_),
    .B(net3911),
    .Y(_02096_));
 sg13g2_a21o_1 _16666_ (.A2(_00116_),
    .A1(net4266),
    .B1(_05084_),
    .X(_02097_));
 sg13g2_a21oi_1 _16667_ (.A1(_03500_),
    .A2(net3739),
    .Y(_02098_),
    .B1(_02096_));
 sg13g2_a22oi_1 _16668_ (.Y(_02099_),
    .B1(_02097_),
    .B2(_02098_),
    .A2(net3753),
    .A1(_00119_));
 sg13g2_a221oi_1 _16669_ (.B2(_02098_),
    .C1(_03501_),
    .B1(_02097_),
    .A1(_00119_),
    .Y(_02100_),
    .A2(net3753));
 sg13g2_xnor2_1 _16670_ (.Y(_02101_),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ),
    .B(_02094_));
 sg13g2_o21ai_1 _16671_ (.B1(_02095_),
    .Y(_02102_),
    .A1(_02100_),
    .A2(_02101_));
 sg13g2_xnor2_1 _16672_ (.Y(_02103_),
    .A(_03500_),
    .B(_02092_));
 sg13g2_nor2b_1 _16673_ (.A(_02103_),
    .B_N(_02102_),
    .Y(_02104_));
 sg13g2_a21o_1 _16674_ (.A2(_02092_),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ),
    .B1(_02104_),
    .X(_02105_));
 sg13g2_xnor2_1 _16675_ (.Y(_02106_),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ),
    .B(_02088_));
 sg13g2_a21oi_1 _16676_ (.A1(_02105_),
    .A2(_02106_),
    .Y(_02107_),
    .B1(_02091_));
 sg13g2_a22oi_1 _16677_ (.Y(_02108_),
    .B1(_02089_),
    .B2(_02107_),
    .A2(_02087_),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ));
 sg13g2_a21oi_2 _16678_ (.B1(_02108_),
    .Y(_02109_),
    .A2(_00115_),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ));
 sg13g2_nand2_1 _16679_ (.Y(_02110_),
    .A(net3701),
    .B(_02109_));
 sg13g2_mux2_2 _16680_ (.A0(net4491),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[455] ),
    .X(_02111_));
 sg13g2_nand2_1 _16681_ (.Y(_02112_),
    .A(\spiking_network_top_uut.all_data_out[99] ),
    .B(_02111_));
 sg13g2_mux2_2 _16682_ (.A0(net4492),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[451] ),
    .X(_02113_));
 sg13g2_nand2_1 _16683_ (.Y(_02114_),
    .A(\spiking_network_top_uut.all_data_out[97] ),
    .B(_02113_));
 sg13g2_nor2_1 _16684_ (.A(_02112_),
    .B(_02114_),
    .Y(_02115_));
 sg13g2_and4_2 _16685_ (.A(\spiking_network_top_uut.all_data_out[98] ),
    .B(\spiking_network_top_uut.all_data_out[96] ),
    .C(_02111_),
    .D(_02113_),
    .X(_02116_));
 sg13g2_nand4_1 _16686_ (.B(\spiking_network_top_uut.all_data_out[96] ),
    .C(_02111_),
    .A(\spiking_network_top_uut.all_data_out[98] ),
    .Y(_02117_),
    .D(_02113_));
 sg13g2_xor2_1 _16687_ (.B(_02114_),
    .A(_02112_),
    .X(_02118_));
 sg13g2_a21oi_2 _16688_ (.B1(_02115_),
    .Y(_02119_),
    .A2(_02118_),
    .A1(_02117_));
 sg13g2_mux2_2 _16689_ (.A0(net4489),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[463] ),
    .X(_02120_));
 sg13g2_nand2_2 _16690_ (.Y(_02121_),
    .A(\spiking_network_top_uut.all_data_out[103] ),
    .B(_02120_));
 sg13g2_mux2_2 _16691_ (.A0(net4490),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[459] ),
    .X(_02122_));
 sg13g2_nand2_1 _16692_ (.Y(_02123_),
    .A(\spiking_network_top_uut.all_data_out[101] ),
    .B(_02122_));
 sg13g2_nor2_1 _16693_ (.A(_02121_),
    .B(_02123_),
    .Y(_02124_));
 sg13g2_nand2_2 _16694_ (.Y(_02125_),
    .A(\spiking_network_top_uut.all_data_out[102] ),
    .B(_02120_));
 sg13g2_nand2_1 _16695_ (.Y(_02126_),
    .A(\spiking_network_top_uut.all_data_out[100] ),
    .B(_02122_));
 sg13g2_or2_2 _16696_ (.X(_02127_),
    .B(_02126_),
    .A(_02125_));
 sg13g2_xor2_1 _16697_ (.B(_02123_),
    .A(_02121_),
    .X(_02128_));
 sg13g2_a21oi_2 _16698_ (.B1(_02124_),
    .Y(_02129_),
    .A2(_02128_),
    .A1(_02127_));
 sg13g2_mux2_2 _16699_ (.A0(net4488),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[467] ),
    .X(_02130_));
 sg13g2_mux2_2 _16700_ (.A0(net4487),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[471] ),
    .X(_02131_));
 sg13g2_a22oi_1 _16701_ (.Y(_02132_),
    .B1(_02131_),
    .B2(\spiking_network_top_uut.all_data_out[107] ),
    .A2(_02130_),
    .A1(\spiking_network_top_uut.all_data_out[105] ));
 sg13g2_and4_1 _16702_ (.A(\spiking_network_top_uut.all_data_out[105] ),
    .B(\spiking_network_top_uut.all_data_out[107] ),
    .C(_02130_),
    .D(_02131_),
    .X(_02133_));
 sg13g2_nand4_1 _16703_ (.B(\spiking_network_top_uut.all_data_out[107] ),
    .C(_02130_),
    .A(\spiking_network_top_uut.all_data_out[105] ),
    .Y(_02134_),
    .D(_02131_));
 sg13g2_and4_1 _16704_ (.A(\spiking_network_top_uut.all_data_out[104] ),
    .B(\spiking_network_top_uut.all_data_out[106] ),
    .C(_02130_),
    .D(_02131_),
    .X(_02135_));
 sg13g2_nand4_1 _16705_ (.B(\spiking_network_top_uut.all_data_out[106] ),
    .C(_02130_),
    .A(\spiking_network_top_uut.all_data_out[104] ),
    .Y(_02136_),
    .D(_02131_));
 sg13g2_nand3b_1 _16706_ (.B(_02134_),
    .C(_02135_),
    .Y(_02137_),
    .A_N(_02132_));
 sg13g2_a21oi_2 _16707_ (.B1(_02132_),
    .Y(_02138_),
    .A2(_02135_),
    .A1(_02134_));
 sg13g2_mux2_2 _16708_ (.A0(net4485),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[479] ),
    .X(_02139_));
 sg13g2_mux2_2 _16709_ (.A0(net4486),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[475] ),
    .X(_02140_));
 sg13g2_and4_1 _16710_ (.A(\spiking_network_top_uut.all_data_out[111] ),
    .B(\spiking_network_top_uut.all_data_out[109] ),
    .C(_02139_),
    .D(_02140_),
    .X(_02141_));
 sg13g2_nand4_1 _16711_ (.B(\spiking_network_top_uut.all_data_out[109] ),
    .C(_02139_),
    .A(\spiking_network_top_uut.all_data_out[111] ),
    .Y(_02142_),
    .D(_02140_));
 sg13g2_and4_1 _16712_ (.A(\spiking_network_top_uut.all_data_out[110] ),
    .B(\spiking_network_top_uut.all_data_out[108] ),
    .C(_02139_),
    .D(_02140_),
    .X(_02143_));
 sg13g2_a22oi_1 _16713_ (.Y(_02144_),
    .B1(_02140_),
    .B2(\spiking_network_top_uut.all_data_out[109] ),
    .A2(_02139_),
    .A1(\spiking_network_top_uut.all_data_out[111] ));
 sg13g2_or3_2 _16714_ (.A(_02141_),
    .B(_02143_),
    .C(_02144_),
    .X(_02145_));
 sg13g2_o21ai_1 _16715_ (.B1(_02142_),
    .Y(_02146_),
    .A1(_02143_),
    .A2(_02144_));
 sg13g2_nand3b_1 _16716_ (.B(_02138_),
    .C(_02146_),
    .Y(_02147_),
    .A_N(_02129_));
 sg13g2_or2_1 _16717_ (.X(_02148_),
    .B(_02147_),
    .A(_02119_));
 sg13g2_inv_2 _16718_ (.Y(_02149_),
    .A(_02148_));
 sg13g2_nor2_1 _16719_ (.A(_02138_),
    .B(_02146_),
    .Y(_02150_));
 sg13g2_nand2_1 _16720_ (.Y(_02151_),
    .A(_02129_),
    .B(_02150_));
 sg13g2_mux2_2 _16721_ (.A0(_02147_),
    .A1(_02151_),
    .S(_02119_),
    .X(_02152_));
 sg13g2_xnor2_1 _16722_ (.Y(_02153_),
    .A(_02089_),
    .B(_02107_));
 sg13g2_xor2_1 _16723_ (.B(_02153_),
    .A(_02152_),
    .X(_02154_));
 sg13g2_o21ai_1 _16724_ (.B1(_02143_),
    .Y(_02155_),
    .A1(_02141_),
    .A2(_02144_));
 sg13g2_o21ai_1 _16725_ (.B1(_02136_),
    .Y(_02156_),
    .A1(_02132_),
    .A2(_02133_));
 sg13g2_o21ai_1 _16726_ (.B1(_02135_),
    .Y(_02157_),
    .A1(_02132_),
    .A2(_02133_));
 sg13g2_nand3b_1 _16727_ (.B(_02134_),
    .C(_02136_),
    .Y(_02158_),
    .A_N(_02132_));
 sg13g2_a22oi_1 _16728_ (.Y(_02159_),
    .B1(_02157_),
    .B2(_02158_),
    .A2(_02155_),
    .A1(_02145_));
 sg13g2_xor2_1 _16729_ (.B(_02128_),
    .A(_02127_),
    .X(_02160_));
 sg13g2_xnor2_1 _16730_ (.Y(_02161_),
    .A(_02127_),
    .B(_02128_));
 sg13g2_and4_1 _16731_ (.A(_02145_),
    .B(_02155_),
    .C(_02157_),
    .D(_02158_),
    .X(_02162_));
 sg13g2_nand4_1 _16732_ (.B(_02155_),
    .C(_02157_),
    .A(_02145_),
    .Y(_02163_),
    .D(_02158_));
 sg13g2_and4_1 _16733_ (.A(_02137_),
    .B(_02145_),
    .C(_02155_),
    .D(_02156_),
    .X(_02164_));
 sg13g2_a22oi_1 _16734_ (.Y(_02165_),
    .B1(_02156_),
    .B2(_02137_),
    .A2(_02155_),
    .A1(_02145_));
 sg13g2_nor3_1 _16735_ (.A(_02159_),
    .B(_02160_),
    .C(_02162_),
    .Y(_02166_));
 sg13g2_o21ai_1 _16736_ (.B1(_02161_),
    .Y(_02167_),
    .A1(_02164_),
    .A2(_02165_));
 sg13g2_a21oi_2 _16737_ (.B1(_02159_),
    .Y(_02168_),
    .A2(_02163_),
    .A1(_02161_));
 sg13g2_xor2_1 _16738_ (.B(_02146_),
    .A(_02138_),
    .X(_02169_));
 sg13g2_xnor2_1 _16739_ (.Y(_02170_),
    .A(_02129_),
    .B(_02169_));
 sg13g2_nand2b_1 _16740_ (.Y(_02171_),
    .B(_02170_),
    .A_N(_02168_));
 sg13g2_xnor2_1 _16741_ (.Y(_02172_),
    .A(_02168_),
    .B(_02170_));
 sg13g2_nand2b_1 _16742_ (.Y(_02173_),
    .B(_02172_),
    .A_N(_02119_));
 sg13g2_nand2_1 _16743_ (.Y(_02174_),
    .A(_02171_),
    .B(_02173_));
 sg13g2_nand2_1 _16744_ (.Y(_02175_),
    .A(_02147_),
    .B(_02151_));
 sg13g2_xor2_1 _16745_ (.B(_02175_),
    .A(_02119_),
    .X(_02176_));
 sg13g2_and2_1 _16746_ (.A(_02174_),
    .B(_02176_),
    .X(_02177_));
 sg13g2_xor2_1 _16747_ (.B(_02176_),
    .A(_02174_),
    .X(_02178_));
 sg13g2_xnor2_1 _16748_ (.Y(_02179_),
    .A(_02105_),
    .B(_02106_));
 sg13g2_inv_1 _16749_ (.Y(_02180_),
    .A(_02179_));
 sg13g2_a21o_1 _16750_ (.A2(_02180_),
    .A1(_02178_),
    .B1(_02177_),
    .X(_02181_));
 sg13g2_nand2_1 _16751_ (.Y(_02182_),
    .A(_02154_),
    .B(_02181_));
 sg13g2_a22oi_1 _16752_ (.Y(_02183_),
    .B1(_02140_),
    .B2(\spiking_network_top_uut.all_data_out[108] ),
    .A2(_02139_),
    .A1(\spiking_network_top_uut.all_data_out[110] ));
 sg13g2_nor2_1 _16753_ (.A(_02143_),
    .B(_02183_),
    .Y(_02184_));
 sg13g2_a22oi_1 _16754_ (.Y(_02185_),
    .B1(_02131_),
    .B2(\spiking_network_top_uut.all_data_out[106] ),
    .A2(_02130_),
    .A1(\spiking_network_top_uut.all_data_out[104] ));
 sg13g2_nor2_1 _16755_ (.A(_02135_),
    .B(_02185_),
    .Y(_02186_));
 sg13g2_and2_1 _16756_ (.A(_02184_),
    .B(_02186_),
    .X(_02187_));
 sg13g2_xor2_1 _16757_ (.B(_02126_),
    .A(_02125_),
    .X(_02188_));
 sg13g2_xor2_1 _16758_ (.B(_02186_),
    .A(_02184_),
    .X(_02189_));
 sg13g2_a21oi_1 _16759_ (.A1(_02188_),
    .A2(_02189_),
    .Y(_02190_),
    .B1(_02187_));
 sg13g2_a21o_1 _16760_ (.A2(_02189_),
    .A1(_02188_),
    .B1(_02187_),
    .X(_02191_));
 sg13g2_nor3_1 _16761_ (.A(_02161_),
    .B(_02164_),
    .C(_02165_),
    .Y(_02192_));
 sg13g2_o21ai_1 _16762_ (.B1(_02160_),
    .Y(_02193_),
    .A1(_02159_),
    .A2(_02162_));
 sg13g2_nor3_1 _16763_ (.A(_02166_),
    .B(_02190_),
    .C(_02192_),
    .Y(_02194_));
 sg13g2_nand3_1 _16764_ (.B(_02191_),
    .C(_02193_),
    .A(_02167_),
    .Y(_02195_));
 sg13g2_xnor2_1 _16765_ (.Y(_02196_),
    .A(_02116_),
    .B(_02118_));
 sg13g2_xnor2_1 _16766_ (.Y(_02197_),
    .A(_02117_),
    .B(_02118_));
 sg13g2_a21oi_2 _16767_ (.B1(_02191_),
    .Y(_02198_),
    .A2(_02193_),
    .A1(_02167_));
 sg13g2_o21ai_1 _16768_ (.B1(_02190_),
    .Y(_02199_),
    .A1(_02166_),
    .A2(_02192_));
 sg13g2_nor3_1 _16769_ (.A(_02194_),
    .B(_02196_),
    .C(_02198_),
    .Y(_02200_));
 sg13g2_nand3_1 _16770_ (.B(_02197_),
    .C(_02199_),
    .A(_02195_),
    .Y(_02201_));
 sg13g2_o21ai_1 _16771_ (.B1(_02195_),
    .Y(_02202_),
    .A1(_02196_),
    .A2(_02198_));
 sg13g2_xnor2_1 _16772_ (.Y(_02203_),
    .A(_02119_),
    .B(_02172_));
 sg13g2_nand2_1 _16773_ (.Y(_02204_),
    .A(_02202_),
    .B(_02203_));
 sg13g2_xnor2_1 _16774_ (.Y(_02205_),
    .A(_02202_),
    .B(_02203_));
 sg13g2_xor2_1 _16775_ (.B(_02103_),
    .A(_02102_),
    .X(_02206_));
 sg13g2_o21ai_1 _16776_ (.B1(_02204_),
    .Y(_02207_),
    .A1(_02205_),
    .A2(_02206_));
 sg13g2_xnor2_1 _16777_ (.Y(_02208_),
    .A(_02178_),
    .B(_02180_));
 sg13g2_nand2b_1 _16778_ (.Y(_02209_),
    .B(_02207_),
    .A_N(_02208_));
 sg13g2_a22oi_1 _16779_ (.Y(_02210_),
    .B1(_02113_),
    .B2(\spiking_network_top_uut.all_data_out[96] ),
    .A2(_02111_),
    .A1(\spiking_network_top_uut.all_data_out[98] ));
 sg13g2_xnor2_1 _16780_ (.Y(_02211_),
    .A(_02188_),
    .B(_02189_));
 sg13g2_nor3_2 _16781_ (.A(_02116_),
    .B(_02210_),
    .C(_02211_),
    .Y(_02212_));
 sg13g2_a21oi_1 _16782_ (.A1(_02195_),
    .A2(_02199_),
    .Y(_02213_),
    .B1(_02197_));
 sg13g2_o21ai_1 _16783_ (.B1(_02196_),
    .Y(_02214_),
    .A1(_02194_),
    .A2(_02198_));
 sg13g2_nand3_1 _16784_ (.B(_02212_),
    .C(_02214_),
    .A(_02201_),
    .Y(_02215_));
 sg13g2_a21oi_2 _16785_ (.B1(_02212_),
    .Y(_02216_),
    .A2(_02214_),
    .A1(_02201_));
 sg13g2_nor3_1 _16786_ (.A(_02200_),
    .B(_02212_),
    .C(_02213_),
    .Y(_02217_));
 sg13g2_o21ai_1 _16787_ (.B1(_02212_),
    .Y(_02218_),
    .A1(_02200_),
    .A2(_02213_));
 sg13g2_nand2b_2 _16788_ (.Y(_02219_),
    .B(_02218_),
    .A_N(_02217_));
 sg13g2_xor2_1 _16789_ (.B(_02101_),
    .A(_02100_),
    .X(_02220_));
 sg13g2_inv_1 _16790_ (.Y(_02221_),
    .A(_02220_));
 sg13g2_o21ai_1 _16791_ (.B1(_02215_),
    .Y(_02222_),
    .A1(_02216_),
    .A2(_02221_));
 sg13g2_xor2_1 _16792_ (.B(_02206_),
    .A(_02205_),
    .X(_02223_));
 sg13g2_nand2_1 _16793_ (.Y(_02224_),
    .A(_02222_),
    .B(_02223_));
 sg13g2_xnor2_1 _16794_ (.Y(_02225_),
    .A(_02219_),
    .B(_02220_));
 sg13g2_o21ai_1 _16795_ (.B1(_02211_),
    .Y(_02226_),
    .A1(_02116_),
    .A2(_02210_));
 sg13g2_nand2b_2 _16796_ (.Y(_02227_),
    .B(_02226_),
    .A_N(_02212_));
 sg13g2_xnor2_1 _16797_ (.Y(_02228_),
    .A(_03501_),
    .B(_02099_));
 sg13g2_nor2_1 _16798_ (.A(_02227_),
    .B(_02228_),
    .Y(_02229_));
 sg13g2_inv_1 _16799_ (.Y(_02230_),
    .A(_02229_));
 sg13g2_xnor2_1 _16800_ (.Y(_02231_),
    .A(_02222_),
    .B(_02223_));
 sg13g2_or3_1 _16801_ (.A(_02225_),
    .B(_02230_),
    .C(_02231_),
    .X(_02232_));
 sg13g2_xor2_1 _16802_ (.B(_02208_),
    .A(_02207_),
    .X(_02233_));
 sg13g2_a21o_1 _16803_ (.A2(_02232_),
    .A1(_02224_),
    .B1(_02233_),
    .X(_02234_));
 sg13g2_xnor2_1 _16804_ (.Y(_02235_),
    .A(_02154_),
    .B(_02181_));
 sg13g2_a21o_1 _16805_ (.A2(_02234_),
    .A1(_02209_),
    .B1(_02235_),
    .X(_02236_));
 sg13g2_a21oi_1 _16806_ (.A1(_02152_),
    .A2(_02153_),
    .Y(_02237_),
    .B1(_02149_));
 sg13g2_xnor2_1 _16807_ (.Y(_02238_),
    .A(_02109_),
    .B(_02152_));
 sg13g2_nor2_1 _16808_ (.A(_02237_),
    .B(_02238_),
    .Y(_02239_));
 sg13g2_xnor2_1 _16809_ (.Y(_02240_),
    .A(_02237_),
    .B(_02238_));
 sg13g2_nand3_1 _16810_ (.B(_02236_),
    .C(_02240_),
    .A(_02182_),
    .Y(_02241_));
 sg13g2_a21oi_1 _16811_ (.A1(_02182_),
    .A2(_02236_),
    .Y(_02242_),
    .B1(_02240_));
 sg13g2_nand3b_1 _16812_ (.B(_02064_),
    .C(_02241_),
    .Y(_02243_),
    .A_N(_02242_));
 sg13g2_and2_1 _16813_ (.A(_02110_),
    .B(_02243_),
    .X(_02244_));
 sg13g2_nand3_1 _16814_ (.B(_02234_),
    .C(_02235_),
    .A(_02209_),
    .Y(_02245_));
 sg13g2_and2_1 _16815_ (.A(_02064_),
    .B(_02236_),
    .X(_02246_));
 sg13g2_a22oi_1 _16816_ (.Y(_02247_),
    .B1(_02245_),
    .B2(_02246_),
    .A2(_02153_),
    .A1(net3701));
 sg13g2_a21o_1 _16817_ (.A2(_02243_),
    .A1(_02110_),
    .B1(_02247_),
    .X(_02248_));
 sg13g2_o21ai_1 _16818_ (.B1(_02109_),
    .Y(_02249_),
    .A1(net3701),
    .A2(_02149_));
 sg13g2_nor3_1 _16819_ (.A(_02109_),
    .B(_02149_),
    .C(_02152_),
    .Y(_02250_));
 sg13g2_or3_1 _16820_ (.A(_02239_),
    .B(_02242_),
    .C(_02250_),
    .X(_02251_));
 sg13g2_o21ai_1 _16821_ (.B1(_02249_),
    .Y(_02252_),
    .A1(net3701),
    .A2(_02251_));
 sg13g2_a21oi_2 _16822_ (.B1(net3645),
    .Y(_02253_),
    .A2(_02252_),
    .A1(_02248_));
 sg13g2_a21oi_2 _16823_ (.B1(_02252_),
    .Y(_02254_),
    .A2(_02247_),
    .A1(_02244_));
 sg13g2_nor2_1 _16824_ (.A(net3701),
    .B(_02227_),
    .Y(_02255_));
 sg13g2_xnor2_1 _16825_ (.Y(_02256_),
    .A(_02228_),
    .B(_02255_));
 sg13g2_o21ai_1 _16826_ (.B1(_02253_),
    .Y(_02257_),
    .A1(_02254_),
    .A2(_02256_));
 sg13g2_xor2_1 _16827_ (.B(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[0] ),
    .A(net4316),
    .X(_02258_));
 sg13g2_a21oi_1 _16828_ (.A1(net3645),
    .A2(_02258_),
    .Y(_02259_),
    .B1(net3957));
 sg13g2_a22oi_1 _16829_ (.Y(_00946_),
    .B1(_02257_),
    .B2(_02259_),
    .A2(_03458_),
    .A1(net3957));
 sg13g2_nand2_1 _16830_ (.Y(_02260_),
    .A(net3701),
    .B(_02220_));
 sg13g2_xnor2_1 _16831_ (.Y(_02261_),
    .A(_02225_),
    .B(_02230_));
 sg13g2_o21ai_1 _16832_ (.B1(_02260_),
    .Y(_02262_),
    .A1(net3701),
    .A2(_02261_));
 sg13g2_o21ai_1 _16833_ (.B1(_02253_),
    .Y(_02263_),
    .A1(_02254_),
    .A2(_02262_));
 sg13g2_xor2_1 _16834_ (.B(_04916_),
    .A(_04915_),
    .X(_02264_));
 sg13g2_a21oi_1 _16835_ (.A1(net3645),
    .A2(_02264_),
    .Y(_02265_),
    .B1(net3956));
 sg13g2_a22oi_1 _16836_ (.Y(_00947_),
    .B1(_02263_),
    .B2(_02265_),
    .A2(_03457_),
    .A1(net3956));
 sg13g2_o21ai_1 _16837_ (.B1(_02231_),
    .Y(_02266_),
    .A1(_02225_),
    .A2(_02230_));
 sg13g2_nand3_1 _16838_ (.B(_02232_),
    .C(_02266_),
    .A(_02064_),
    .Y(_02267_));
 sg13g2_o21ai_1 _16839_ (.B1(_02267_),
    .Y(_02268_),
    .A1(_02064_),
    .A2(_02206_));
 sg13g2_o21ai_1 _16840_ (.B1(_02253_),
    .Y(_02269_),
    .A1(_02254_),
    .A2(_02268_));
 sg13g2_xnor2_1 _16841_ (.Y(_02270_),
    .A(_04913_),
    .B(_04917_));
 sg13g2_a21oi_1 _16842_ (.A1(net3645),
    .A2(_02270_),
    .Y(_02271_),
    .B1(net3956));
 sg13g2_a22oi_1 _16843_ (.Y(_00948_),
    .B1(_02269_),
    .B2(_02271_),
    .A2(_03456_),
    .A1(net3956));
 sg13g2_nand3_1 _16844_ (.B(_02232_),
    .C(_02233_),
    .A(_02224_),
    .Y(_02272_));
 sg13g2_nand3_1 _16845_ (.B(_02234_),
    .C(_02272_),
    .A(_02064_),
    .Y(_02273_));
 sg13g2_o21ai_1 _16846_ (.B1(_02273_),
    .Y(_02274_),
    .A1(_02064_),
    .A2(_02179_));
 sg13g2_o21ai_1 _16847_ (.B1(_02253_),
    .Y(_02275_),
    .A1(_02254_),
    .A2(_02274_));
 sg13g2_or3_1 _16848_ (.A(_04911_),
    .B(_04912_),
    .C(_04918_),
    .X(_02276_));
 sg13g2_and2_1 _16849_ (.A(_04919_),
    .B(_02276_),
    .X(_02277_));
 sg13g2_a21oi_1 _16850_ (.A1(net3645),
    .A2(_02277_),
    .Y(_02278_),
    .B1(net3956));
 sg13g2_a22oi_1 _16851_ (.Y(_00949_),
    .B1(_02275_),
    .B2(_02278_),
    .A2(_03455_),
    .A1(net3956));
 sg13g2_o21ai_1 _16852_ (.B1(net4606),
    .Y(_02279_),
    .A1(_04909_),
    .A2(_04920_));
 sg13g2_a21oi_1 _16853_ (.A1(_04922_),
    .A2(_02252_),
    .Y(_02280_),
    .B1(_02279_));
 sg13g2_a21oi_1 _16854_ (.A1(net3957),
    .A2(_03454_),
    .Y(_00950_),
    .B1(_02280_));
 sg13g2_mux4_1 _16855_ (.S0(\spiking_network_top_uut.all_data_out[508] ),
    .A0(net3789),
    .A1(net3788),
    .A2(net3787),
    .A3(net3786),
    .S1(\spiking_network_top_uut.all_data_out[509] ),
    .X(_02281_));
 sg13g2_mux2_1 _16856_ (.A0(net3783),
    .A1(net3899),
    .S(\spiking_network_top_uut.all_data_out[508] ),
    .X(_02282_));
 sg13g2_nor2b_1 _16857_ (.A(\spiking_network_top_uut.all_data_out[508] ),
    .B_N(net3785),
    .Y(_02283_));
 sg13g2_a21oi_1 _16858_ (.A1(\spiking_network_top_uut.all_data_out[508] ),
    .A2(net3784),
    .Y(_02284_),
    .B1(_02283_));
 sg13g2_o21ai_1 _16859_ (.B1(\spiking_network_top_uut.all_data_out[510] ),
    .Y(_02285_),
    .A1(\spiking_network_top_uut.all_data_out[509] ),
    .A2(_02284_));
 sg13g2_a21oi_1 _16860_ (.A1(\spiking_network_top_uut.all_data_out[509] ),
    .A2(_02282_),
    .Y(_02286_),
    .B1(_02285_));
 sg13g2_o21ai_1 _16861_ (.B1(net4638),
    .Y(_02287_),
    .A1(\spiking_network_top_uut.all_data_out[510] ),
    .A2(_02281_));
 sg13g2_nand2_1 _16862_ (.Y(_02288_),
    .A(net3962),
    .B(net205));
 sg13g2_o21ai_1 _16863_ (.B1(_02288_),
    .Y(_00951_),
    .A1(_02286_),
    .A2(_02287_));
 sg13g2_mux2_1 _16864_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_dout ),
    .A1(net205),
    .S(net4644),
    .X(_00952_));
 sg13g2_mux4_1 _16865_ (.S0(\spiking_network_top_uut.all_data_out[504] ),
    .A0(net3840),
    .A1(net3839),
    .A2(net3838),
    .A3(net3837),
    .S1(\spiking_network_top_uut.all_data_out[505] ),
    .X(_02289_));
 sg13g2_mux2_1 _16866_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[6] ),
    .A1(net3834),
    .S(\spiking_network_top_uut.all_data_out[504] ),
    .X(_02290_));
 sg13g2_nor2b_1 _16867_ (.A(\spiking_network_top_uut.all_data_out[504] ),
    .B_N(net3836),
    .Y(_02291_));
 sg13g2_a21oi_1 _16868_ (.A1(\spiking_network_top_uut.all_data_out[504] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[5] ),
    .Y(_02292_),
    .B1(_02291_));
 sg13g2_o21ai_1 _16869_ (.B1(\spiking_network_top_uut.all_data_out[506] ),
    .Y(_02293_),
    .A1(\spiking_network_top_uut.all_data_out[505] ),
    .A2(_02292_));
 sg13g2_a21oi_1 _16870_ (.A1(\spiking_network_top_uut.all_data_out[505] ),
    .A2(_02290_),
    .Y(_02294_),
    .B1(_02293_));
 sg13g2_o21ai_1 _16871_ (.B1(net4642),
    .Y(_02295_),
    .A1(\spiking_network_top_uut.all_data_out[506] ),
    .A2(_02289_));
 sg13g2_nand2_1 _16872_ (.Y(_02296_),
    .A(net3963),
    .B(net227));
 sg13g2_o21ai_1 _16873_ (.B1(_02296_),
    .Y(_00953_),
    .A1(_02294_),
    .A2(_02295_));
 sg13g2_mux2_1 _16874_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_dout ),
    .A1(net227),
    .S(net4643),
    .X(_00954_));
 sg13g2_mux4_1 _16875_ (.S0(\spiking_network_top_uut.all_data_out[500] ),
    .A0(net3833),
    .A1(net3832),
    .A2(net3831),
    .A3(net3830),
    .S1(\spiking_network_top_uut.all_data_out[501] ),
    .X(_02297_));
 sg13g2_mux2_1 _16876_ (.A0(net3828),
    .A1(net3827),
    .S(\spiking_network_top_uut.all_data_out[500] ),
    .X(_02298_));
 sg13g2_nor2b_1 _16877_ (.A(\spiking_network_top_uut.all_data_out[500] ),
    .B_N(net3829),
    .Y(_02299_));
 sg13g2_a21oi_1 _16878_ (.A1(\spiking_network_top_uut.all_data_out[500] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[5] ),
    .Y(_02300_),
    .B1(_02299_));
 sg13g2_o21ai_1 _16879_ (.B1(\spiking_network_top_uut.all_data_out[502] ),
    .Y(_02301_),
    .A1(\spiking_network_top_uut.all_data_out[501] ),
    .A2(_02300_));
 sg13g2_a21oi_1 _16880_ (.A1(\spiking_network_top_uut.all_data_out[501] ),
    .A2(_02298_),
    .Y(_02302_),
    .B1(_02301_));
 sg13g2_o21ai_1 _16881_ (.B1(net4608),
    .Y(_02303_),
    .A1(\spiking_network_top_uut.all_data_out[502] ),
    .A2(_02297_));
 sg13g2_nand2_1 _16882_ (.Y(_02304_),
    .A(net3966),
    .B(net232));
 sg13g2_o21ai_1 _16883_ (.B1(_02304_),
    .Y(_00955_),
    .A1(_02302_),
    .A2(_02303_));
 sg13g2_mux2_1 _16884_ (.A0(net318),
    .A1(net232),
    .S(net4609),
    .X(_00956_));
 sg13g2_mux4_1 _16885_ (.S0(\spiking_network_top_uut.all_data_out[496] ),
    .A0(net3826),
    .A1(net3825),
    .A2(net3824),
    .A3(net3823),
    .S1(\spiking_network_top_uut.all_data_out[497] ),
    .X(_02305_));
 sg13g2_mux2_1 _16886_ (.A0(net3821),
    .A1(net3820),
    .S(\spiking_network_top_uut.all_data_out[496] ),
    .X(_02306_));
 sg13g2_nor2b_1 _16887_ (.A(\spiking_network_top_uut.all_data_out[496] ),
    .B_N(net3822),
    .Y(_02307_));
 sg13g2_a21oi_1 _16888_ (.A1(\spiking_network_top_uut.all_data_out[496] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[5] ),
    .Y(_02308_),
    .B1(_02307_));
 sg13g2_o21ai_1 _16889_ (.B1(\spiking_network_top_uut.all_data_out[498] ),
    .Y(_02309_),
    .A1(\spiking_network_top_uut.all_data_out[497] ),
    .A2(_02308_));
 sg13g2_a21oi_1 _16890_ (.A1(\spiking_network_top_uut.all_data_out[497] ),
    .A2(_02306_),
    .Y(_02310_),
    .B1(_02309_));
 sg13g2_o21ai_1 _16891_ (.B1(net4613),
    .Y(_02311_),
    .A1(\spiking_network_top_uut.all_data_out[498] ),
    .A2(_02305_));
 sg13g2_nand2_1 _16892_ (.Y(_02312_),
    .A(net3965),
    .B(net112));
 sg13g2_o21ai_1 _16893_ (.B1(_02312_),
    .Y(_00957_),
    .A1(_02310_),
    .A2(_02311_));
 sg13g2_mux2_1 _16894_ (.A0(net368),
    .A1(net112),
    .S(net4616),
    .X(_00958_));
 sg13g2_mux4_1 _16895_ (.S0(\spiking_network_top_uut.all_data_out[492] ),
    .A0(net3819),
    .A1(net3818),
    .A2(net3817),
    .A3(net3816),
    .S1(\spiking_network_top_uut.all_data_out[493] ),
    .X(_02313_));
 sg13g2_mux2_1 _16896_ (.A0(net3814),
    .A1(net3813),
    .S(\spiking_network_top_uut.all_data_out[492] ),
    .X(_02314_));
 sg13g2_nor2b_1 _16897_ (.A(\spiking_network_top_uut.all_data_out[492] ),
    .B_N(net3815),
    .Y(_02315_));
 sg13g2_a21oi_1 _16898_ (.A1(\spiking_network_top_uut.all_data_out[492] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[5] ),
    .Y(_02316_),
    .B1(_02315_));
 sg13g2_o21ai_1 _16899_ (.B1(\spiking_network_top_uut.all_data_out[494] ),
    .Y(_02317_),
    .A1(\spiking_network_top_uut.all_data_out[493] ),
    .A2(_02316_));
 sg13g2_a21oi_1 _16900_ (.A1(\spiking_network_top_uut.all_data_out[493] ),
    .A2(_02314_),
    .Y(_02318_),
    .B1(_02317_));
 sg13g2_o21ai_1 _16901_ (.B1(net4627),
    .Y(_02319_),
    .A1(\spiking_network_top_uut.all_data_out[494] ),
    .A2(_02313_));
 sg13g2_nand2_1 _16902_ (.Y(_02320_),
    .A(net3960),
    .B(net52));
 sg13g2_o21ai_1 _16903_ (.B1(_02320_),
    .Y(_00959_),
    .A1(_02318_),
    .A2(_02319_));
 sg13g2_mux2_1 _16904_ (.A0(net252),
    .A1(net52),
    .S(net4627),
    .X(_00960_));
 sg13g2_nand2b_1 _16905_ (.Y(_02321_),
    .B(\spiking_network_top_uut.all_data_out[488] ),
    .A_N(net3807));
 sg13g2_nor2_1 _16906_ (.A(\spiking_network_top_uut.all_data_out[488] ),
    .B(net3808),
    .Y(_02322_));
 sg13g2_nor2_1 _16907_ (.A(\spiking_network_top_uut.all_data_out[489] ),
    .B(_02322_),
    .Y(_02323_));
 sg13g2_mux2_1 _16908_ (.A0(net3806),
    .A1(net3805),
    .S(\spiking_network_top_uut.all_data_out[488] ),
    .X(_02324_));
 sg13g2_a221oi_1 _16909_ (.B2(\spiking_network_top_uut.all_data_out[489] ),
    .C1(_03617_),
    .B1(_02324_),
    .A1(_02321_),
    .Y(_02325_),
    .A2(_02323_));
 sg13g2_mux4_1 _16910_ (.S0(\spiking_network_top_uut.all_data_out[488] ),
    .A0(net3812),
    .A1(net3811),
    .A2(net3810),
    .A3(net3809),
    .S1(\spiking_network_top_uut.all_data_out[489] ),
    .X(_02326_));
 sg13g2_o21ai_1 _16911_ (.B1(net4621),
    .Y(_02327_),
    .A1(\spiking_network_top_uut.all_data_out[490] ),
    .A2(_02326_));
 sg13g2_nand2_1 _16912_ (.Y(_02328_),
    .A(net3959),
    .B(net135));
 sg13g2_o21ai_1 _16913_ (.B1(_02328_),
    .Y(_00961_),
    .A1(_02325_),
    .A2(_02327_));
 sg13g2_mux2_1 _16914_ (.A0(net327),
    .A1(net135),
    .S(net4621),
    .X(_00962_));
 sg13g2_nand2b_1 _16915_ (.Y(_02329_),
    .B(\spiking_network_top_uut.all_data_out[484] ),
    .A_N(net3799));
 sg13g2_nor2_1 _16916_ (.A(\spiking_network_top_uut.all_data_out[484] ),
    .B(net3800),
    .Y(_02330_));
 sg13g2_nor2_1 _16917_ (.A(\spiking_network_top_uut.all_data_out[485] ),
    .B(_02330_),
    .Y(_02331_));
 sg13g2_mux2_1 _16918_ (.A0(net3798),
    .A1(net3797),
    .S(\spiking_network_top_uut.all_data_out[484] ),
    .X(_02332_));
 sg13g2_a221oi_1 _16919_ (.B2(\spiking_network_top_uut.all_data_out[485] ),
    .C1(_03538_),
    .B1(_02332_),
    .A1(_02329_),
    .Y(_02333_),
    .A2(_02331_));
 sg13g2_mux4_1 _16920_ (.S0(\spiking_network_top_uut.all_data_out[484] ),
    .A0(net3804),
    .A1(net3803),
    .A2(net3802),
    .A3(net3801),
    .S1(\spiking_network_top_uut.all_data_out[485] ),
    .X(_02334_));
 sg13g2_o21ai_1 _16921_ (.B1(net4632),
    .Y(_02335_),
    .A1(\spiking_network_top_uut.all_data_out[486] ),
    .A2(_02334_));
 sg13g2_nand2_1 _16922_ (.Y(_02336_),
    .A(net3961),
    .B(net49));
 sg13g2_o21ai_1 _16923_ (.B1(_02336_),
    .Y(_00963_),
    .A1(_02333_),
    .A2(_02335_));
 sg13g2_mux2_1 _16924_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_dout ),
    .A1(net49),
    .S(net4632),
    .X(_00964_));
 sg13g2_mux4_1 _16925_ (.S0(\spiking_network_top_uut.all_data_out[480] ),
    .A0(net3796),
    .A1(net3795),
    .A2(net3794),
    .A3(net3793),
    .S1(\spiking_network_top_uut.all_data_out[481] ),
    .X(_02337_));
 sg13g2_mux2_1 _16926_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[6] ),
    .A1(net3790),
    .S(\spiking_network_top_uut.all_data_out[480] ),
    .X(_02338_));
 sg13g2_nor2b_1 _16927_ (.A(\spiking_network_top_uut.all_data_out[480] ),
    .B_N(net3792),
    .Y(_02339_));
 sg13g2_a21oi_1 _16928_ (.A1(\spiking_network_top_uut.all_data_out[480] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[5] ),
    .Y(_02340_),
    .B1(_02339_));
 sg13g2_o21ai_1 _16929_ (.B1(\spiking_network_top_uut.all_data_out[482] ),
    .Y(_02341_),
    .A1(\spiking_network_top_uut.all_data_out[481] ),
    .A2(_02340_));
 sg13g2_a21oi_1 _16930_ (.A1(\spiking_network_top_uut.all_data_out[481] ),
    .A2(_02338_),
    .Y(_02342_),
    .B1(_02341_));
 sg13g2_o21ai_1 _16931_ (.B1(net4635),
    .Y(_02343_),
    .A1(\spiking_network_top_uut.all_data_out[482] ),
    .A2(_02337_));
 sg13g2_nand2_1 _16932_ (.Y(_02344_),
    .A(net3964),
    .B(net133));
 sg13g2_o21ai_1 _16933_ (.B1(_02344_),
    .Y(_00965_),
    .A1(_02342_),
    .A2(_02343_));
 sg13g2_nor3_2 _16934_ (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[2] ),
    .B(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[1] ),
    .C(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[0] ),
    .Y(_02345_));
 sg13g2_nor2b_1 _16935_ (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[3] ),
    .B_N(_02345_),
    .Y(_02346_));
 sg13g2_nor2b_2 _16936_ (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[4] ),
    .B_N(_02346_),
    .Y(_02347_));
 sg13g2_nand2b_1 _16937_ (.Y(_02348_),
    .B(_02346_),
    .A_N(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[4] ));
 sg13g2_o21ai_1 _16938_ (.B1(net4604),
    .Y(_02349_),
    .A1(net3640),
    .A2(net3700));
 sg13g2_nor2b_1 _16939_ (.A(net3641),
    .B_N(net340),
    .Y(_02350_));
 sg13g2_a21oi_1 _16940_ (.A1(net4284),
    .A2(net3640),
    .Y(_02351_),
    .B1(_02350_));
 sg13g2_nand2_1 _16941_ (.Y(_02352_),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[0] ),
    .B(_02349_));
 sg13g2_o21ai_1 _16942_ (.B1(_02352_),
    .Y(_00966_),
    .A1(_02349_),
    .A2(_02351_));
 sg13g2_xor2_1 _16943_ (.B(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[0] ),
    .A(net387),
    .X(_02353_));
 sg13g2_nor2_1 _16944_ (.A(net3640),
    .B(_02353_),
    .Y(_02354_));
 sg13g2_a21oi_1 _16945_ (.A1(net4281),
    .A2(net3640),
    .Y(_02355_),
    .B1(_02354_));
 sg13g2_nand2_1 _16946_ (.Y(_02356_),
    .A(net387),
    .B(_02349_));
 sg13g2_o21ai_1 _16947_ (.B1(_02356_),
    .Y(_00967_),
    .A1(_02349_),
    .A2(_02355_));
 sg13g2_o21ai_1 _16948_ (.B1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[2] ),
    .Y(_02357_),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[1] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[0] ));
 sg13g2_nor2b_1 _16949_ (.A(_02345_),
    .B_N(_02357_),
    .Y(_02358_));
 sg13g2_nor2_1 _16950_ (.A(net3640),
    .B(_02358_),
    .Y(_02359_));
 sg13g2_a21oi_1 _16951_ (.A1(net4277),
    .A2(net3640),
    .Y(_02360_),
    .B1(_02359_));
 sg13g2_nand2_1 _16952_ (.Y(_02361_),
    .A(net190),
    .B(_02349_));
 sg13g2_o21ai_1 _16953_ (.B1(_02361_),
    .Y(_00968_),
    .A1(_02349_),
    .A2(_02360_));
 sg13g2_nand2_1 _16954_ (.Y(_02362_),
    .A(net4274),
    .B(net3640));
 sg13g2_xnor2_1 _16955_ (.Y(_02363_),
    .A(net396),
    .B(_02345_));
 sg13g2_o21ai_1 _16956_ (.B1(_02362_),
    .Y(_02364_),
    .A1(net3641),
    .A2(_02363_));
 sg13g2_mux2_1 _16957_ (.A0(_02364_),
    .A1(net396),
    .S(_02349_),
    .X(_00969_));
 sg13g2_nand2_1 _16958_ (.Y(_02365_),
    .A(net3949),
    .B(net297));
 sg13g2_nand2b_1 _16959_ (.Y(_02366_),
    .B(net297),
    .A_N(_02346_));
 sg13g2_a21oi_1 _16960_ (.A1(net3700),
    .A2(_02366_),
    .Y(_02367_),
    .B1(net3641));
 sg13g2_a21oi_1 _16961_ (.A1(net4270),
    .A2(net3640),
    .Y(_02368_),
    .B1(_02367_));
 sg13g2_o21ai_1 _16962_ (.B1(_02365_),
    .Y(_00970_),
    .A1(_02349_),
    .A2(_02368_));
 sg13g2_mux2_1 _16963_ (.A0(net277),
    .A1(net133),
    .S(net4634),
    .X(_00971_));
 sg13g2_a21oi_1 _16964_ (.A1(net3914),
    .A2(net3910),
    .Y(_02369_),
    .B1(_00121_));
 sg13g2_nor2_2 _16965_ (.A(net3745),
    .B(_02369_),
    .Y(_02370_));
 sg13g2_nor2_1 _16966_ (.A(_00121_),
    .B(_02370_),
    .Y(_02371_));
 sg13g2_nor2_1 _16967_ (.A(_00121_),
    .B(_02371_),
    .Y(_02372_));
 sg13g2_nand2b_1 _16968_ (.Y(_02373_),
    .B(_02370_),
    .A_N(_00121_));
 sg13g2_o21ai_1 _16969_ (.B1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ),
    .Y(_02374_),
    .A1(_00121_),
    .A2(_02370_));
 sg13g2_inv_1 _16970_ (.Y(_02375_),
    .A(_02374_));
 sg13g2_a21o_1 _16971_ (.A2(net3744),
    .A1(_00122_),
    .B1(_02370_),
    .X(_02376_));
 sg13g2_nor2_1 _16972_ (.A(_00122_),
    .B(net3904),
    .Y(_02377_));
 sg13g2_a221oi_1 _16973_ (.B2(_02369_),
    .C1(_02377_),
    .B1(net3904),
    .A1(_03502_),
    .Y(_02378_),
    .A2(net3744));
 sg13g2_nand2_1 _16974_ (.Y(_02379_),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ),
    .B(_02378_));
 sg13g2_and2_1 _16975_ (.A(_00125_),
    .B(net3744),
    .X(_02380_));
 sg13g2_nor2_1 _16976_ (.A(_00122_),
    .B(_05105_),
    .Y(_02381_));
 sg13g2_nor2_1 _16977_ (.A(_00121_),
    .B(net3910),
    .Y(_02382_));
 sg13g2_o21ai_1 _16978_ (.B1(net3917),
    .Y(_02383_),
    .A1(_00123_),
    .A2(net3904));
 sg13g2_nor3_1 _16979_ (.A(_02381_),
    .B(_02382_),
    .C(_02383_),
    .Y(_02384_));
 sg13g2_nor2_1 _16980_ (.A(_02380_),
    .B(_02384_),
    .Y(_02385_));
 sg13g2_nor3_1 _16981_ (.A(_03503_),
    .B(_02380_),
    .C(_02384_),
    .Y(_02386_));
 sg13g2_xnor2_1 _16982_ (.Y(_02387_),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ),
    .B(_02378_));
 sg13g2_o21ai_1 _16983_ (.B1(_02379_),
    .Y(_02388_),
    .A1(_02386_),
    .A2(_02387_));
 sg13g2_xnor2_1 _16984_ (.Y(_02389_),
    .A(_03502_),
    .B(_02376_));
 sg13g2_nor2b_1 _16985_ (.A(_02389_),
    .B_N(_02388_),
    .Y(_02390_));
 sg13g2_a21o_1 _16986_ (.A2(_02376_),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ),
    .B1(_02390_),
    .X(_02391_));
 sg13g2_xnor2_1 _16987_ (.Y(_02392_),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ),
    .B(_02371_));
 sg13g2_a21oi_1 _16988_ (.A1(_02391_),
    .A2(_02392_),
    .Y(_02393_),
    .B1(_02375_));
 sg13g2_a22oi_1 _16989_ (.Y(_02394_),
    .B1(_02373_),
    .B2(_02393_),
    .A2(_02370_),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ));
 sg13g2_a21oi_2 _16990_ (.B1(_02394_),
    .Y(_02395_),
    .A2(_00121_),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ));
 sg13g2_a21o_1 _16991_ (.A2(_00121_),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ),
    .B1(_02394_),
    .X(_02396_));
 sg13g2_mux2_2 _16992_ (.A0(net4491),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[487] ),
    .X(_02397_));
 sg13g2_nand2_1 _16993_ (.Y(_02398_),
    .A(\spiking_network_top_uut.all_data_out[115] ),
    .B(_02397_));
 sg13g2_mux2_2 _16994_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.din ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[483] ),
    .X(_02399_));
 sg13g2_nand2_1 _16995_ (.Y(_02400_),
    .A(\spiking_network_top_uut.all_data_out[113] ),
    .B(_02399_));
 sg13g2_nor2_1 _16996_ (.A(_02398_),
    .B(_02400_),
    .Y(_02401_));
 sg13g2_and4_1 _16997_ (.A(\spiking_network_top_uut.all_data_out[114] ),
    .B(\spiking_network_top_uut.all_data_out[112] ),
    .C(_02397_),
    .D(_02399_),
    .X(_02402_));
 sg13g2_nand4_1 _16998_ (.B(\spiking_network_top_uut.all_data_out[112] ),
    .C(_02397_),
    .A(\spiking_network_top_uut.all_data_out[114] ),
    .Y(_02403_),
    .D(_02399_));
 sg13g2_xor2_1 _16999_ (.B(_02400_),
    .A(_02398_),
    .X(_02404_));
 sg13g2_a21oi_2 _17000_ (.B1(_02401_),
    .Y(_02405_),
    .A2(_02404_),
    .A1(_02403_));
 sg13g2_mux2_2 _17001_ (.A0(net4489),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[495] ),
    .X(_02406_));
 sg13g2_nand2_1 _17002_ (.Y(_02407_),
    .A(\spiking_network_top_uut.all_data_out[119] ),
    .B(_02406_));
 sg13g2_mux2_2 _17003_ (.A0(net4490),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[491] ),
    .X(_02408_));
 sg13g2_nand2_1 _17004_ (.Y(_02409_),
    .A(\spiking_network_top_uut.all_data_out[117] ),
    .B(_02408_));
 sg13g2_nor2_1 _17005_ (.A(_02407_),
    .B(_02409_),
    .Y(_02410_));
 sg13g2_nand2_1 _17006_ (.Y(_02411_),
    .A(\spiking_network_top_uut.all_data_out[118] ),
    .B(_02406_));
 sg13g2_nand2_1 _17007_ (.Y(_02412_),
    .A(\spiking_network_top_uut.all_data_out[116] ),
    .B(_02408_));
 sg13g2_or2_2 _17008_ (.X(_02413_),
    .B(_02412_),
    .A(_02411_));
 sg13g2_xor2_1 _17009_ (.B(_02409_),
    .A(_02407_),
    .X(_02414_));
 sg13g2_a21oi_2 _17010_ (.B1(_02410_),
    .Y(_02415_),
    .A2(_02414_),
    .A1(_02413_));
 sg13g2_mux2_2 _17011_ (.A0(net4487),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[503] ),
    .X(_02416_));
 sg13g2_mux2_2 _17012_ (.A0(net4488),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[499] ),
    .X(_02417_));
 sg13g2_a22oi_1 _17013_ (.Y(_02418_),
    .B1(_02417_),
    .B2(\spiking_network_top_uut.all_data_out[121] ),
    .A2(_02416_),
    .A1(\spiking_network_top_uut.all_data_out[123] ));
 sg13g2_and4_1 _17014_ (.A(\spiking_network_top_uut.all_data_out[123] ),
    .B(\spiking_network_top_uut.all_data_out[121] ),
    .C(_02416_),
    .D(_02417_),
    .X(_02419_));
 sg13g2_nand4_1 _17015_ (.B(\spiking_network_top_uut.all_data_out[121] ),
    .C(_02416_),
    .A(\spiking_network_top_uut.all_data_out[123] ),
    .Y(_02420_),
    .D(_02417_));
 sg13g2_and4_2 _17016_ (.A(\spiking_network_top_uut.all_data_out[122] ),
    .B(\spiking_network_top_uut.all_data_out[120] ),
    .C(_02416_),
    .D(_02417_),
    .X(_02421_));
 sg13g2_nand4_1 _17017_ (.B(\spiking_network_top_uut.all_data_out[120] ),
    .C(_02416_),
    .A(\spiking_network_top_uut.all_data_out[122] ),
    .Y(_02422_),
    .D(_02417_));
 sg13g2_nand3b_1 _17018_ (.B(_02420_),
    .C(_02421_),
    .Y(_02423_),
    .A_N(_02418_));
 sg13g2_a21oi_2 _17019_ (.B1(_02418_),
    .Y(_02424_),
    .A2(_02421_),
    .A1(_02420_));
 sg13g2_mux2_2 _17020_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.din ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[507] ),
    .X(_02425_));
 sg13g2_mux2_2 _17021_ (.A0(net4485),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[511] ),
    .X(_02426_));
 sg13g2_and4_1 _17022_ (.A(\spiking_network_top_uut.all_data_out[125] ),
    .B(\spiking_network_top_uut.all_data_out[127] ),
    .C(_02425_),
    .D(_02426_),
    .X(_02427_));
 sg13g2_nand4_1 _17023_ (.B(\spiking_network_top_uut.all_data_out[127] ),
    .C(_02425_),
    .A(\spiking_network_top_uut.all_data_out[125] ),
    .Y(_02428_),
    .D(_02426_));
 sg13g2_and4_1 _17024_ (.A(\spiking_network_top_uut.all_data_out[124] ),
    .B(\spiking_network_top_uut.all_data_out[126] ),
    .C(_02425_),
    .D(_02426_),
    .X(_02429_));
 sg13g2_a22oi_1 _17025_ (.Y(_02430_),
    .B1(_02426_),
    .B2(\spiking_network_top_uut.all_data_out[127] ),
    .A2(_02425_),
    .A1(\spiking_network_top_uut.all_data_out[125] ));
 sg13g2_or3_2 _17026_ (.A(_02427_),
    .B(_02429_),
    .C(_02430_),
    .X(_02431_));
 sg13g2_o21ai_1 _17027_ (.B1(_02428_),
    .Y(_02432_),
    .A1(_02429_),
    .A2(_02430_));
 sg13g2_nand3b_1 _17028_ (.B(_02424_),
    .C(_02432_),
    .Y(_02433_),
    .A_N(_02415_));
 sg13g2_nor2_1 _17029_ (.A(_02405_),
    .B(_02433_),
    .Y(_02434_));
 sg13g2_or2_1 _17030_ (.X(_02435_),
    .B(_02433_),
    .A(_02405_));
 sg13g2_a21oi_1 _17031_ (.A1(_02347_),
    .A2(_02435_),
    .Y(_02436_),
    .B1(_02396_));
 sg13g2_nor2_1 _17032_ (.A(_02424_),
    .B(_02432_),
    .Y(_02437_));
 sg13g2_nand2_2 _17033_ (.Y(_02438_),
    .A(_02415_),
    .B(_02437_));
 sg13g2_mux2_2 _17034_ (.A0(_02433_),
    .A1(_02438_),
    .S(_02405_),
    .X(_02439_));
 sg13g2_xnor2_1 _17035_ (.Y(_02440_),
    .A(_02372_),
    .B(_02393_));
 sg13g2_inv_1 _17036_ (.Y(_02441_),
    .A(_02440_));
 sg13g2_xnor2_1 _17037_ (.Y(_02442_),
    .A(_02439_),
    .B(_02440_));
 sg13g2_o21ai_1 _17038_ (.B1(_02429_),
    .Y(_02443_),
    .A1(_02427_),
    .A2(_02430_));
 sg13g2_o21ai_1 _17039_ (.B1(_02422_),
    .Y(_02444_),
    .A1(_02418_),
    .A2(_02419_));
 sg13g2_o21ai_1 _17040_ (.B1(_02421_),
    .Y(_02445_),
    .A1(_02418_),
    .A2(_02419_));
 sg13g2_nand3b_1 _17041_ (.B(_02420_),
    .C(_02422_),
    .Y(_02446_),
    .A_N(_02418_));
 sg13g2_a22oi_1 _17042_ (.Y(_02447_),
    .B1(_02445_),
    .B2(_02446_),
    .A2(_02443_),
    .A1(_02431_));
 sg13g2_xor2_1 _17043_ (.B(_02414_),
    .A(_02413_),
    .X(_02448_));
 sg13g2_xnor2_1 _17044_ (.Y(_02449_),
    .A(_02413_),
    .B(_02414_));
 sg13g2_and4_1 _17045_ (.A(_02431_),
    .B(_02443_),
    .C(_02445_),
    .D(_02446_),
    .X(_02450_));
 sg13g2_nand4_1 _17046_ (.B(_02443_),
    .C(_02445_),
    .A(_02431_),
    .Y(_02451_),
    .D(_02446_));
 sg13g2_and4_1 _17047_ (.A(_02423_),
    .B(_02431_),
    .C(_02443_),
    .D(_02444_),
    .X(_02452_));
 sg13g2_a22oi_1 _17048_ (.Y(_02453_),
    .B1(_02444_),
    .B2(_02423_),
    .A2(_02443_),
    .A1(_02431_));
 sg13g2_nor3_2 _17049_ (.A(_02447_),
    .B(_02448_),
    .C(_02450_),
    .Y(_02454_));
 sg13g2_a21oi_2 _17050_ (.B1(_02447_),
    .Y(_02455_),
    .A2(_02451_),
    .A1(_02449_));
 sg13g2_xor2_1 _17051_ (.B(_02432_),
    .A(_02424_),
    .X(_02456_));
 sg13g2_xnor2_1 _17052_ (.Y(_02457_),
    .A(_02415_),
    .B(_02456_));
 sg13g2_nand2b_1 _17053_ (.Y(_02458_),
    .B(_02457_),
    .A_N(_02455_));
 sg13g2_xnor2_1 _17054_ (.Y(_02459_),
    .A(_02455_),
    .B(_02457_));
 sg13g2_nand2b_1 _17055_ (.Y(_02460_),
    .B(_02459_),
    .A_N(_02405_));
 sg13g2_nand2_2 _17056_ (.Y(_02461_),
    .A(_02458_),
    .B(_02460_));
 sg13g2_nand2_1 _17057_ (.Y(_02462_),
    .A(_02433_),
    .B(_02438_));
 sg13g2_xor2_1 _17058_ (.B(_02462_),
    .A(_02405_),
    .X(_02463_));
 sg13g2_and2_1 _17059_ (.A(_02461_),
    .B(_02463_),
    .X(_02464_));
 sg13g2_xor2_1 _17060_ (.B(_02463_),
    .A(_02461_),
    .X(_02465_));
 sg13g2_xnor2_1 _17061_ (.Y(_02466_),
    .A(_02391_),
    .B(_02392_));
 sg13g2_inv_1 _17062_ (.Y(_02467_),
    .A(_02466_));
 sg13g2_a21o_1 _17063_ (.A2(_02467_),
    .A1(_02465_),
    .B1(_02464_),
    .X(_02468_));
 sg13g2_nand2_1 _17064_ (.Y(_02469_),
    .A(_02442_),
    .B(_02468_));
 sg13g2_a22oi_1 _17065_ (.Y(_02470_),
    .B1(_02426_),
    .B2(\spiking_network_top_uut.all_data_out[126] ),
    .A2(_02425_),
    .A1(\spiking_network_top_uut.all_data_out[124] ));
 sg13g2_nor2_1 _17066_ (.A(_02429_),
    .B(_02470_),
    .Y(_02471_));
 sg13g2_a22oi_1 _17067_ (.Y(_02472_),
    .B1(_02417_),
    .B2(\spiking_network_top_uut.all_data_out[120] ),
    .A2(_02416_),
    .A1(\spiking_network_top_uut.all_data_out[122] ));
 sg13g2_nor2_1 _17068_ (.A(_02421_),
    .B(_02472_),
    .Y(_02473_));
 sg13g2_and2_1 _17069_ (.A(_02471_),
    .B(_02473_),
    .X(_02474_));
 sg13g2_xor2_1 _17070_ (.B(_02412_),
    .A(_02411_),
    .X(_02475_));
 sg13g2_xor2_1 _17071_ (.B(_02473_),
    .A(_02471_),
    .X(_02476_));
 sg13g2_a21oi_2 _17072_ (.B1(_02474_),
    .Y(_02477_),
    .A2(_02476_),
    .A1(_02475_));
 sg13g2_nor3_2 _17073_ (.A(_02449_),
    .B(_02452_),
    .C(_02453_),
    .Y(_02478_));
 sg13g2_nor3_1 _17074_ (.A(_02454_),
    .B(_02477_),
    .C(_02478_),
    .Y(_02479_));
 sg13g2_or3_1 _17075_ (.A(_02454_),
    .B(_02477_),
    .C(_02478_),
    .X(_02480_));
 sg13g2_xnor2_1 _17076_ (.Y(_02481_),
    .A(_02403_),
    .B(_02404_));
 sg13g2_o21ai_1 _17077_ (.B1(_02477_),
    .Y(_02482_),
    .A1(_02454_),
    .A2(_02478_));
 sg13g2_nand3_1 _17078_ (.B(_02481_),
    .C(_02482_),
    .A(_02480_),
    .Y(_02483_));
 sg13g2_a21o_2 _17079_ (.A2(_02482_),
    .A1(_02481_),
    .B1(_02479_),
    .X(_02484_));
 sg13g2_xnor2_1 _17080_ (.Y(_02485_),
    .A(_02405_),
    .B(_02459_));
 sg13g2_nand2_1 _17081_ (.Y(_02486_),
    .A(_02484_),
    .B(_02485_));
 sg13g2_xnor2_1 _17082_ (.Y(_02487_),
    .A(_02484_),
    .B(_02485_));
 sg13g2_xor2_1 _17083_ (.B(_02389_),
    .A(_02388_),
    .X(_02488_));
 sg13g2_o21ai_1 _17084_ (.B1(_02486_),
    .Y(_02489_),
    .A1(_02487_),
    .A2(_02488_));
 sg13g2_xnor2_1 _17085_ (.Y(_02490_),
    .A(_02465_),
    .B(_02467_));
 sg13g2_nor2b_1 _17086_ (.A(_02490_),
    .B_N(_02489_),
    .Y(_02491_));
 sg13g2_a22oi_1 _17087_ (.Y(_02492_),
    .B1(_02399_),
    .B2(\spiking_network_top_uut.all_data_out[112] ),
    .A2(_02397_),
    .A1(\spiking_network_top_uut.all_data_out[114] ));
 sg13g2_xnor2_1 _17088_ (.Y(_02493_),
    .A(_02475_),
    .B(_02476_));
 sg13g2_nor3_2 _17089_ (.A(_02402_),
    .B(_02492_),
    .C(_02493_),
    .Y(_02494_));
 sg13g2_a21o_2 _17090_ (.A2(_02482_),
    .A1(_02480_),
    .B1(_02481_),
    .X(_02495_));
 sg13g2_and3_1 _17091_ (.X(_02496_),
    .A(_02483_),
    .B(_02494_),
    .C(_02495_));
 sg13g2_nand3_1 _17092_ (.B(_02494_),
    .C(_02495_),
    .A(_02483_),
    .Y(_02497_));
 sg13g2_a21oi_1 _17093_ (.A1(_02483_),
    .A2(_02495_),
    .Y(_02498_),
    .B1(_02494_));
 sg13g2_xor2_1 _17094_ (.B(_02387_),
    .A(_02386_),
    .X(_02499_));
 sg13g2_inv_1 _17095_ (.Y(_02500_),
    .A(_02499_));
 sg13g2_nor3_1 _17096_ (.A(_02496_),
    .B(_02498_),
    .C(_02500_),
    .Y(_02501_));
 sg13g2_o21ai_1 _17097_ (.B1(_02497_),
    .Y(_02502_),
    .A1(_02498_),
    .A2(_02500_));
 sg13g2_xor2_1 _17098_ (.B(_02488_),
    .A(_02487_),
    .X(_02503_));
 sg13g2_nand2_1 _17099_ (.Y(_02504_),
    .A(_02502_),
    .B(_02503_));
 sg13g2_o21ai_1 _17100_ (.B1(_02500_),
    .Y(_02505_),
    .A1(_02496_),
    .A2(_02498_));
 sg13g2_nand2b_1 _17101_ (.Y(_02506_),
    .B(_02505_),
    .A_N(_02501_));
 sg13g2_xnor2_1 _17102_ (.Y(_02507_),
    .A(_03503_),
    .B(_02385_));
 sg13g2_o21ai_1 _17103_ (.B1(_02493_),
    .Y(_02508_),
    .A1(_02402_),
    .A2(_02492_));
 sg13g2_nand2b_2 _17104_ (.Y(_02509_),
    .B(_02508_),
    .A_N(_02494_));
 sg13g2_nor2_1 _17105_ (.A(_02507_),
    .B(_02509_),
    .Y(_02510_));
 sg13g2_nand3b_1 _17106_ (.B(_02505_),
    .C(_02510_),
    .Y(_02511_),
    .A_N(_02501_));
 sg13g2_xnor2_1 _17107_ (.Y(_02512_),
    .A(_02502_),
    .B(_02503_));
 sg13g2_or2_1 _17108_ (.X(_02513_),
    .B(_02512_),
    .A(_02511_));
 sg13g2_o21ai_1 _17109_ (.B1(_02504_),
    .Y(_02514_),
    .A1(_02511_),
    .A2(_02512_));
 sg13g2_nand2b_1 _17110_ (.Y(_02515_),
    .B(_02490_),
    .A_N(_02489_));
 sg13g2_nand2b_1 _17111_ (.Y(_02516_),
    .B(_02515_),
    .A_N(_02491_));
 sg13g2_nor2b_1 _17112_ (.A(_02516_),
    .B_N(_02514_),
    .Y(_02517_));
 sg13g2_a21oi_1 _17113_ (.A1(_02514_),
    .A2(_02515_),
    .Y(_02518_),
    .B1(_02491_));
 sg13g2_xnor2_1 _17114_ (.Y(_02519_),
    .A(_02442_),
    .B(_02468_));
 sg13g2_nor2_1 _17115_ (.A(_02518_),
    .B(_02519_),
    .Y(_02520_));
 sg13g2_o21ai_1 _17116_ (.B1(_02469_),
    .Y(_02521_),
    .A1(_02518_),
    .A2(_02519_));
 sg13g2_a21oi_1 _17117_ (.A1(_02439_),
    .A2(_02441_),
    .Y(_02522_),
    .B1(_02434_));
 sg13g2_nor2_1 _17118_ (.A(_02395_),
    .B(_02439_),
    .Y(_02523_));
 sg13g2_xnor2_1 _17119_ (.Y(_02524_),
    .A(_02395_),
    .B(_02439_));
 sg13g2_nor2_1 _17120_ (.A(_02522_),
    .B(_02524_),
    .Y(_02525_));
 sg13g2_xor2_1 _17121_ (.B(_02524_),
    .A(_02522_),
    .X(_02526_));
 sg13g2_a221oi_1 _17122_ (.B2(_02521_),
    .C1(_02525_),
    .B1(_02526_),
    .A1(_02435_),
    .Y(_02527_),
    .A2(_02523_));
 sg13g2_nand2_1 _17123_ (.Y(_02528_),
    .A(net3700),
    .B(_02396_));
 sg13g2_a21o_1 _17124_ (.A2(_02527_),
    .A1(_02347_),
    .B1(_02436_),
    .X(_02529_));
 sg13g2_xor2_1 _17125_ (.B(_02526_),
    .A(_02521_),
    .X(_02530_));
 sg13g2_o21ai_1 _17126_ (.B1(_02528_),
    .Y(_02531_),
    .A1(net3700),
    .A2(_02530_));
 sg13g2_nand2_1 _17127_ (.Y(_02532_),
    .A(_02518_),
    .B(_02519_));
 sg13g2_nor2_1 _17128_ (.A(net3700),
    .B(_02520_),
    .Y(_02533_));
 sg13g2_a22oi_1 _17129_ (.Y(_02534_),
    .B1(_02532_),
    .B2(_02533_),
    .A2(_02441_),
    .A1(net3700));
 sg13g2_or2_1 _17130_ (.X(_02535_),
    .B(_02534_),
    .A(_02531_));
 sg13g2_a21o_1 _17131_ (.A2(_02535_),
    .A1(_02529_),
    .B1(net3642),
    .X(_02536_));
 sg13g2_a21oi_2 _17132_ (.B1(_02529_),
    .Y(_02537_),
    .A2(_02534_),
    .A1(_02531_));
 sg13g2_nor2_1 _17133_ (.A(_02348_),
    .B(_02509_),
    .Y(_02538_));
 sg13g2_xnor2_1 _17134_ (.Y(_02539_),
    .A(_02507_),
    .B(_02538_));
 sg13g2_o21ai_1 _17135_ (.B1(net4603),
    .Y(_02540_),
    .A1(_02537_),
    .A2(_02539_));
 sg13g2_xor2_1 _17136_ (.B(net496),
    .A(net4313),
    .X(_02541_));
 sg13g2_a22oi_1 _17137_ (.Y(_02542_),
    .B1(_00006_),
    .B2(_02541_),
    .A2(net496),
    .A1(net3949));
 sg13g2_o21ai_1 _17138_ (.B1(_02542_),
    .Y(_00972_),
    .A1(_02536_),
    .A2(_02540_));
 sg13g2_xnor2_1 _17139_ (.Y(_02543_),
    .A(_02506_),
    .B(_02510_));
 sg13g2_nand2_1 _17140_ (.Y(_02544_),
    .A(_02348_),
    .B(_02499_));
 sg13g2_a21oi_1 _17141_ (.A1(_02347_),
    .A2(_02543_),
    .Y(_02545_),
    .B1(_02537_));
 sg13g2_a21o_1 _17142_ (.A2(_02545_),
    .A1(_02544_),
    .B1(_02536_),
    .X(_02546_));
 sg13g2_xor2_1 _17143_ (.B(_04931_),
    .A(_04930_),
    .X(_02547_));
 sg13g2_a21oi_1 _17144_ (.A1(net3642),
    .A2(_02547_),
    .Y(_02548_),
    .B1(net3947));
 sg13g2_a22oi_1 _17145_ (.Y(_00973_),
    .B1(_02546_),
    .B2(_02548_),
    .A2(_03461_),
    .A1(net3947));
 sg13g2_nor2_1 _17146_ (.A(_02347_),
    .B(_02488_),
    .Y(_02549_));
 sg13g2_nand2_1 _17147_ (.Y(_02550_),
    .A(_02347_),
    .B(_02513_));
 sg13g2_a21oi_1 _17148_ (.A1(_02511_),
    .A2(_02512_),
    .Y(_02551_),
    .B1(_02550_));
 sg13g2_nor3_1 _17149_ (.A(_02537_),
    .B(_02549_),
    .C(_02551_),
    .Y(_02552_));
 sg13g2_or2_1 _17150_ (.X(_02553_),
    .B(_02552_),
    .A(_02536_));
 sg13g2_xnor2_1 _17151_ (.Y(_02554_),
    .A(_04928_),
    .B(_04932_));
 sg13g2_a21oi_1 _17152_ (.A1(net3642),
    .A2(_02554_),
    .Y(_02555_),
    .B1(net3947));
 sg13g2_a22oi_1 _17153_ (.Y(_00974_),
    .B1(_02553_),
    .B2(_02555_),
    .A2(_03460_),
    .A1(net3947));
 sg13g2_nor2_1 _17154_ (.A(net4603),
    .B(net502),
    .Y(_02556_));
 sg13g2_nand2b_1 _17155_ (.Y(_02557_),
    .B(_02516_),
    .A_N(_02514_));
 sg13g2_nor2_1 _17156_ (.A(net3700),
    .B(_02517_),
    .Y(_02558_));
 sg13g2_a221oi_1 _17157_ (.B2(_02558_),
    .C1(_02537_),
    .B1(_02557_),
    .A1(net3700),
    .Y(_02559_),
    .A2(_02467_));
 sg13g2_or3_1 _17158_ (.A(_04926_),
    .B(_04927_),
    .C(_04933_),
    .X(_02560_));
 sg13g2_and2_1 _17159_ (.A(_04934_),
    .B(_02560_),
    .X(_02561_));
 sg13g2_a21oi_1 _17160_ (.A1(net3642),
    .A2(_02561_),
    .Y(_02562_),
    .B1(net3949));
 sg13g2_o21ai_1 _17161_ (.B1(_02562_),
    .Y(_02563_),
    .A1(_02536_),
    .A2(_02559_));
 sg13g2_nor2b_1 _17162_ (.A(_02556_),
    .B_N(_02563_),
    .Y(_00975_));
 sg13g2_o21ai_1 _17163_ (.B1(net4604),
    .Y(_02564_),
    .A1(_04924_),
    .A2(_04935_));
 sg13g2_a21oi_1 _17164_ (.A1(_04937_),
    .A2(_02529_),
    .Y(_02565_),
    .B1(_02564_));
 sg13g2_a21oi_1 _17165_ (.A1(net3949),
    .A2(_03459_),
    .Y(_00976_),
    .B1(_02565_));
 sg13g2_mux2_1 _17166_ (.A0(net3787),
    .A1(net3786),
    .S(\spiking_network_top_uut.all_data_out[540] ),
    .X(_02566_));
 sg13g2_nor2b_1 _17167_ (.A(\spiking_network_top_uut.all_data_out[540] ),
    .B_N(net3789),
    .Y(_02567_));
 sg13g2_a21oi_1 _17168_ (.A1(\spiking_network_top_uut.all_data_out[540] ),
    .A2(net3788),
    .Y(_02568_),
    .B1(_02567_));
 sg13g2_a21oi_1 _17169_ (.A1(\spiking_network_top_uut.all_data_out[541] ),
    .A2(_02566_),
    .Y(_02569_),
    .B1(\spiking_network_top_uut.all_data_out[542] ));
 sg13g2_o21ai_1 _17170_ (.B1(_02569_),
    .Y(_02570_),
    .A1(\spiking_network_top_uut.all_data_out[541] ),
    .A2(_02568_));
 sg13g2_mux2_1 _17171_ (.A0(net3783),
    .A1(net3899),
    .S(\spiking_network_top_uut.all_data_out[540] ),
    .X(_02571_));
 sg13g2_nor2b_1 _17172_ (.A(\spiking_network_top_uut.all_data_out[540] ),
    .B_N(net3785),
    .Y(_02572_));
 sg13g2_a21oi_1 _17173_ (.A1(\spiking_network_top_uut.all_data_out[540] ),
    .A2(net3784),
    .Y(_02573_),
    .B1(_02572_));
 sg13g2_o21ai_1 _17174_ (.B1(\spiking_network_top_uut.all_data_out[542] ),
    .Y(_02574_),
    .A1(\spiking_network_top_uut.all_data_out[541] ),
    .A2(_02573_));
 sg13g2_a21oi_1 _17175_ (.A1(\spiking_network_top_uut.all_data_out[541] ),
    .A2(_02571_),
    .Y(_02575_),
    .B1(_02574_));
 sg13g2_nand2_1 _17176_ (.Y(_02576_),
    .A(net4637),
    .B(_02570_));
 sg13g2_nand2_1 _17177_ (.Y(_02577_),
    .A(net3962),
    .B(net116));
 sg13g2_o21ai_1 _17178_ (.B1(_02577_),
    .Y(_00977_),
    .A1(_02575_),
    .A2(_02576_));
 sg13g2_mux2_1 _17179_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_dout ),
    .A1(net116),
    .S(net4637),
    .X(_00978_));
 sg13g2_nand2_1 _17180_ (.Y(_02578_),
    .A(\spiking_network_top_uut.all_data_out[536] ),
    .B(_03662_));
 sg13g2_nor2_1 _17181_ (.A(\spiking_network_top_uut.all_data_out[536] ),
    .B(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[4] ),
    .Y(_02579_));
 sg13g2_nor2_1 _17182_ (.A(\spiking_network_top_uut.all_data_out[537] ),
    .B(_02579_),
    .Y(_02580_));
 sg13g2_mux2_1 _17183_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[6] ),
    .A1(net3834),
    .S(\spiking_network_top_uut.all_data_out[536] ),
    .X(_02581_));
 sg13g2_a221oi_1 _17184_ (.B2(\spiking_network_top_uut.all_data_out[537] ),
    .C1(_03612_),
    .B1(_02581_),
    .A1(_02578_),
    .Y(_02582_),
    .A2(_02580_));
 sg13g2_mux4_1 _17185_ (.S0(\spiking_network_top_uut.all_data_out[536] ),
    .A0(net3840),
    .A1(net3839),
    .A2(net3838),
    .A3(net3837),
    .S1(\spiking_network_top_uut.all_data_out[537] ),
    .X(_02583_));
 sg13g2_o21ai_1 _17186_ (.B1(net4642),
    .Y(_02584_),
    .A1(\spiking_network_top_uut.all_data_out[538] ),
    .A2(_02583_));
 sg13g2_nand2_1 _17187_ (.Y(_02585_),
    .A(net3963),
    .B(net90));
 sg13g2_o21ai_1 _17188_ (.B1(_02585_),
    .Y(_00979_),
    .A1(_02582_),
    .A2(_02584_));
 sg13g2_mux2_1 _17189_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_dout ),
    .A1(net90),
    .S(net4639),
    .X(_00980_));
 sg13g2_mux4_1 _17190_ (.S0(\spiking_network_top_uut.all_data_out[532] ),
    .A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[0] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[1] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[2] ),
    .A3(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[3] ),
    .S1(\spiking_network_top_uut.all_data_out[533] ),
    .X(_02586_));
 sg13g2_mux2_1 _17191_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[6] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[7] ),
    .S(\spiking_network_top_uut.all_data_out[532] ),
    .X(_02587_));
 sg13g2_nor2b_1 _17192_ (.A(\spiking_network_top_uut.all_data_out[532] ),
    .B_N(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[4] ),
    .Y(_02588_));
 sg13g2_a21oi_1 _17193_ (.A1(\spiking_network_top_uut.all_data_out[532] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[5] ),
    .Y(_02589_),
    .B1(_02588_));
 sg13g2_o21ai_1 _17194_ (.B1(\spiking_network_top_uut.all_data_out[534] ),
    .Y(_02590_),
    .A1(\spiking_network_top_uut.all_data_out[533] ),
    .A2(_02589_));
 sg13g2_a21oi_1 _17195_ (.A1(\spiking_network_top_uut.all_data_out[533] ),
    .A2(_02587_),
    .Y(_02591_),
    .B1(_02590_));
 sg13g2_o21ai_1 _17196_ (.B1(net4610),
    .Y(_02592_),
    .A1(\spiking_network_top_uut.all_data_out[534] ),
    .A2(_02586_));
 sg13g2_nand2_1 _17197_ (.Y(_02593_),
    .A(net3966),
    .B(net307));
 sg13g2_o21ai_1 _17198_ (.B1(_02593_),
    .Y(_00981_),
    .A1(_02591_),
    .A2(_02592_));
 sg13g2_mux2_1 _17199_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_dout ),
    .A1(net307),
    .S(net4607),
    .X(_00982_));
 sg13g2_mux2_1 _17200_ (.A0(net3824),
    .A1(net3823),
    .S(\spiking_network_top_uut.all_data_out[528] ),
    .X(_02594_));
 sg13g2_nor2b_1 _17201_ (.A(\spiking_network_top_uut.all_data_out[528] ),
    .B_N(net3826),
    .Y(_02595_));
 sg13g2_a21oi_1 _17202_ (.A1(\spiking_network_top_uut.all_data_out[528] ),
    .A2(net3825),
    .Y(_02596_),
    .B1(_02595_));
 sg13g2_a21oi_1 _17203_ (.A1(\spiking_network_top_uut.all_data_out[529] ),
    .A2(_02594_),
    .Y(_02597_),
    .B1(\spiking_network_top_uut.all_data_out[530] ));
 sg13g2_o21ai_1 _17204_ (.B1(_02597_),
    .Y(_02598_),
    .A1(\spiking_network_top_uut.all_data_out[529] ),
    .A2(_02596_));
 sg13g2_mux2_1 _17205_ (.A0(net3821),
    .A1(net3820),
    .S(\spiking_network_top_uut.all_data_out[528] ),
    .X(_02599_));
 sg13g2_nand2_1 _17206_ (.Y(_02600_),
    .A(\spiking_network_top_uut.all_data_out[529] ),
    .B(_02599_));
 sg13g2_a21oi_1 _17207_ (.A1(\spiking_network_top_uut.all_data_out[528] ),
    .A2(_03660_),
    .Y(_02601_),
    .B1(\spiking_network_top_uut.all_data_out[529] ));
 sg13g2_o21ai_1 _17208_ (.B1(_02601_),
    .Y(_02602_),
    .A1(\spiking_network_top_uut.all_data_out[528] ),
    .A2(net3822));
 sg13g2_nand3_1 _17209_ (.B(_02600_),
    .C(_02602_),
    .A(\spiking_network_top_uut.all_data_out[530] ),
    .Y(_02603_));
 sg13g2_nand3_1 _17210_ (.B(_02598_),
    .C(_02603_),
    .A(net4613),
    .Y(_02604_));
 sg13g2_o21ai_1 _17211_ (.B1(_02604_),
    .Y(_00983_),
    .A1(net4611),
    .A2(_03689_));
 sg13g2_mux2_1 _17212_ (.A0(net274),
    .A1(net114),
    .S(net4611),
    .X(_00984_));
 sg13g2_mux4_1 _17213_ (.S0(\spiking_network_top_uut.all_data_out[524] ),
    .A0(net3819),
    .A1(net3818),
    .A2(net3817),
    .A3(net3816),
    .S1(\spiking_network_top_uut.all_data_out[525] ),
    .X(_02605_));
 sg13g2_mux2_1 _17214_ (.A0(net3814),
    .A1(net3813),
    .S(\spiking_network_top_uut.all_data_out[524] ),
    .X(_02606_));
 sg13g2_nor2b_1 _17215_ (.A(\spiking_network_top_uut.all_data_out[524] ),
    .B_N(net3815),
    .Y(_02607_));
 sg13g2_a21oi_1 _17216_ (.A1(\spiking_network_top_uut.all_data_out[524] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[5] ),
    .Y(_02608_),
    .B1(_02607_));
 sg13g2_o21ai_1 _17217_ (.B1(\spiking_network_top_uut.all_data_out[526] ),
    .Y(_02609_),
    .A1(\spiking_network_top_uut.all_data_out[525] ),
    .A2(_02608_));
 sg13g2_a21oi_1 _17218_ (.A1(\spiking_network_top_uut.all_data_out[525] ),
    .A2(_02606_),
    .Y(_02610_),
    .B1(_02609_));
 sg13g2_o21ai_1 _17219_ (.B1(net4627),
    .Y(_02611_),
    .A1(\spiking_network_top_uut.all_data_out[526] ),
    .A2(_02605_));
 sg13g2_nand2_1 _17220_ (.Y(_02612_),
    .A(net3960),
    .B(net45));
 sg13g2_o21ai_1 _17221_ (.B1(_02612_),
    .Y(_00985_),
    .A1(_02610_),
    .A2(_02611_));
 sg13g2_mux2_1 _17222_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_dout ),
    .A1(net45),
    .S(net4627),
    .X(_00986_));
 sg13g2_mux4_1 _17223_ (.S0(\spiking_network_top_uut.all_data_out[520] ),
    .A0(net3812),
    .A1(net3811),
    .A2(net3810),
    .A3(net3809),
    .S1(\spiking_network_top_uut.all_data_out[521] ),
    .X(_02613_));
 sg13g2_mux2_1 _17224_ (.A0(net3806),
    .A1(net3805),
    .S(\spiking_network_top_uut.all_data_out[520] ),
    .X(_02614_));
 sg13g2_nor2b_1 _17225_ (.A(\spiking_network_top_uut.all_data_out[520] ),
    .B_N(net3808),
    .Y(_02615_));
 sg13g2_a21oi_1 _17226_ (.A1(\spiking_network_top_uut.all_data_out[520] ),
    .A2(net3807),
    .Y(_02616_),
    .B1(_02615_));
 sg13g2_o21ai_1 _17227_ (.B1(\spiking_network_top_uut.all_data_out[522] ),
    .Y(_02617_),
    .A1(\spiking_network_top_uut.all_data_out[521] ),
    .A2(_02616_));
 sg13g2_a21oi_1 _17228_ (.A1(\spiking_network_top_uut.all_data_out[521] ),
    .A2(_02614_),
    .Y(_02618_),
    .B1(_02617_));
 sg13g2_o21ai_1 _17229_ (.B1(net4630),
    .Y(_02619_),
    .A1(\spiking_network_top_uut.all_data_out[522] ),
    .A2(_02613_));
 sg13g2_nand2_1 _17230_ (.Y(_02620_),
    .A(net3959),
    .B(net79));
 sg13g2_o21ai_1 _17231_ (.B1(_02620_),
    .Y(_00987_),
    .A1(_02618_),
    .A2(_02619_));
 sg13g2_mux2_1 _17232_ (.A0(net315),
    .A1(net79),
    .S(net4624),
    .X(_00988_));
 sg13g2_mux2_1 _17233_ (.A0(net3802),
    .A1(net3801),
    .S(\spiking_network_top_uut.all_data_out[516] ),
    .X(_02621_));
 sg13g2_nor2b_1 _17234_ (.A(\spiking_network_top_uut.all_data_out[516] ),
    .B_N(net3804),
    .Y(_02622_));
 sg13g2_a21oi_1 _17235_ (.A1(\spiking_network_top_uut.all_data_out[516] ),
    .A2(net3803),
    .Y(_02623_),
    .B1(_02622_));
 sg13g2_a21oi_1 _17236_ (.A1(\spiking_network_top_uut.all_data_out[517] ),
    .A2(_02621_),
    .Y(_02624_),
    .B1(\spiking_network_top_uut.all_data_out[518] ));
 sg13g2_o21ai_1 _17237_ (.B1(_02624_),
    .Y(_02625_),
    .A1(\spiking_network_top_uut.all_data_out[517] ),
    .A2(_02623_));
 sg13g2_mux2_1 _17238_ (.A0(net3798),
    .A1(net3797),
    .S(\spiking_network_top_uut.all_data_out[516] ),
    .X(_02626_));
 sg13g2_nor2b_1 _17239_ (.A(\spiking_network_top_uut.all_data_out[516] ),
    .B_N(net3800),
    .Y(_02627_));
 sg13g2_a21oi_1 _17240_ (.A1(\spiking_network_top_uut.all_data_out[516] ),
    .A2(net3799),
    .Y(_02628_),
    .B1(_02627_));
 sg13g2_o21ai_1 _17241_ (.B1(\spiking_network_top_uut.all_data_out[518] ),
    .Y(_02629_),
    .A1(\spiking_network_top_uut.all_data_out[517] ),
    .A2(_02628_));
 sg13g2_a21oi_1 _17242_ (.A1(\spiking_network_top_uut.all_data_out[517] ),
    .A2(_02626_),
    .Y(_02630_),
    .B1(_02629_));
 sg13g2_nand2_1 _17243_ (.Y(_02631_),
    .A(net4633),
    .B(_02625_));
 sg13g2_nand2_1 _17244_ (.Y(_02632_),
    .A(net3959),
    .B(net145));
 sg13g2_o21ai_1 _17245_ (.B1(_02632_),
    .Y(_00989_),
    .A1(_02630_),
    .A2(_02631_));
 sg13g2_mux2_1 _17246_ (.A0(net262),
    .A1(net145),
    .S(net4624),
    .X(_00990_));
 sg13g2_mux2_1 _17247_ (.A0(net3794),
    .A1(net3793),
    .S(\spiking_network_top_uut.all_data_out[512] ),
    .X(_02633_));
 sg13g2_nor2b_1 _17248_ (.A(\spiking_network_top_uut.all_data_out[512] ),
    .B_N(net3796),
    .Y(_02634_));
 sg13g2_a21oi_1 _17249_ (.A1(\spiking_network_top_uut.all_data_out[512] ),
    .A2(net3795),
    .Y(_02635_),
    .B1(_02634_));
 sg13g2_a21oi_1 _17250_ (.A1(\spiking_network_top_uut.all_data_out[513] ),
    .A2(_02633_),
    .Y(_02636_),
    .B1(\spiking_network_top_uut.all_data_out[514] ));
 sg13g2_o21ai_1 _17251_ (.B1(_02636_),
    .Y(_02637_),
    .A1(\spiking_network_top_uut.all_data_out[513] ),
    .A2(_02635_));
 sg13g2_mux2_1 _17252_ (.A0(net3791),
    .A1(net3790),
    .S(\spiking_network_top_uut.all_data_out[512] ),
    .X(_02638_));
 sg13g2_nand2_1 _17253_ (.Y(_02639_),
    .A(\spiking_network_top_uut.all_data_out[513] ),
    .B(_02638_));
 sg13g2_a21oi_1 _17254_ (.A1(\spiking_network_top_uut.all_data_out[512] ),
    .A2(_03658_),
    .Y(_02640_),
    .B1(\spiking_network_top_uut.all_data_out[513] ));
 sg13g2_o21ai_1 _17255_ (.B1(_02640_),
    .Y(_02641_),
    .A1(\spiking_network_top_uut.all_data_out[512] ),
    .A2(net3792));
 sg13g2_nand3_1 _17256_ (.B(_02639_),
    .C(_02641_),
    .A(\spiking_network_top_uut.all_data_out[514] ),
    .Y(_02642_));
 sg13g2_nand3_1 _17257_ (.B(_02637_),
    .C(_02642_),
    .A(net4619),
    .Y(_02643_));
 sg13g2_o21ai_1 _17258_ (.B1(_02643_),
    .Y(_00991_),
    .A1(net4619),
    .A2(_03690_));
 sg13g2_nor3_2 _17259_ (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[2] ),
    .B(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[1] ),
    .C(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[0] ),
    .Y(_02644_));
 sg13g2_nor2b_2 _17260_ (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[3] ),
    .B_N(_02644_),
    .Y(_02645_));
 sg13g2_nor2b_2 _17261_ (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[4] ),
    .B_N(_02645_),
    .Y(_02646_));
 sg13g2_nand2b_2 _17262_ (.Y(_02647_),
    .B(_02645_),
    .A_N(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[4] ));
 sg13g2_o21ai_1 _17263_ (.B1(net4603),
    .Y(_02648_),
    .A1(net3637),
    .A2(_02647_));
 sg13g2_nor2b_1 _17264_ (.A(net3638),
    .B_N(_00132_),
    .Y(_02649_));
 sg13g2_a21oi_1 _17265_ (.A1(net4284),
    .A2(net3638),
    .Y(_02650_),
    .B1(_02649_));
 sg13g2_nand2_1 _17266_ (.Y(_02651_),
    .A(net363),
    .B(_02648_));
 sg13g2_o21ai_1 _17267_ (.B1(_02651_),
    .Y(_00992_),
    .A1(_02648_),
    .A2(_02650_));
 sg13g2_xor2_1 _17268_ (.B(net363),
    .A(net382),
    .X(_02652_));
 sg13g2_nor2_1 _17269_ (.A(net3638),
    .B(_02652_),
    .Y(_02653_));
 sg13g2_a21oi_1 _17270_ (.A1(net4281),
    .A2(net3637),
    .Y(_02654_),
    .B1(_02653_));
 sg13g2_nand2_1 _17271_ (.Y(_02655_),
    .A(net382),
    .B(_02648_));
 sg13g2_o21ai_1 _17272_ (.B1(_02655_),
    .Y(_00993_),
    .A1(_02648_),
    .A2(_02654_));
 sg13g2_o21ai_1 _17273_ (.B1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[2] ),
    .Y(_02656_),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[1] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[0] ));
 sg13g2_nor2b_1 _17274_ (.A(_02644_),
    .B_N(_02656_),
    .Y(_02657_));
 sg13g2_nor2_1 _17275_ (.A(net3637),
    .B(_02657_),
    .Y(_02658_));
 sg13g2_a21oi_1 _17276_ (.A1(net4277),
    .A2(net3637),
    .Y(_02659_),
    .B1(_02658_));
 sg13g2_nand2_1 _17277_ (.Y(_02660_),
    .A(net244),
    .B(_02648_));
 sg13g2_o21ai_1 _17278_ (.B1(_02660_),
    .Y(_00994_),
    .A1(_02648_),
    .A2(_02659_));
 sg13g2_nand2_1 _17279_ (.Y(_02661_),
    .A(net4274),
    .B(net3637));
 sg13g2_xnor2_1 _17280_ (.Y(_02662_),
    .A(net439),
    .B(_02644_));
 sg13g2_o21ai_1 _17281_ (.B1(_02661_),
    .Y(_02663_),
    .A1(net3637),
    .A2(_02662_));
 sg13g2_mux2_1 _17282_ (.A0(_02663_),
    .A1(net439),
    .S(_02648_),
    .X(_00995_));
 sg13g2_nand2_1 _17283_ (.Y(_02664_),
    .A(net3947),
    .B(net266));
 sg13g2_nand2b_1 _17284_ (.Y(_02665_),
    .B(net266),
    .A_N(_02645_));
 sg13g2_a21oi_1 _17285_ (.A1(_02647_),
    .A2(_02665_),
    .Y(_02666_),
    .B1(net3637));
 sg13g2_a21oi_1 _17286_ (.A1(net4270),
    .A2(net3637),
    .Y(_02667_),
    .B1(_02666_));
 sg13g2_o21ai_1 _17287_ (.B1(_02664_),
    .Y(_00996_),
    .A1(_02648_),
    .A2(_02667_));
 sg13g2_mux2_1 _17288_ (.A0(net345),
    .A1(net171),
    .S(net4646),
    .X(_00997_));
 sg13g2_nor2_1 _17289_ (.A(_00127_),
    .B(net3740),
    .Y(_02668_));
 sg13g2_nor3_2 _17290_ (.A(_00127_),
    .B(net3744),
    .C(_05090_),
    .Y(_02669_));
 sg13g2_nand2_1 _17291_ (.Y(_02670_),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ),
    .B(_00127_));
 sg13g2_a21oi_1 _17292_ (.A1(net3916),
    .A2(net3740),
    .Y(_02671_),
    .B1(_00127_));
 sg13g2_nor2_1 _17293_ (.A(_03463_),
    .B(_02671_),
    .Y(_02672_));
 sg13g2_nand2_1 _17294_ (.Y(_02673_),
    .A(_00128_),
    .B(net3744));
 sg13g2_o21ai_1 _17295_ (.B1(_02673_),
    .Y(_02674_),
    .A1(net3744),
    .A2(_02668_));
 sg13g2_nor2_1 _17296_ (.A(_00128_),
    .B(net3903),
    .Y(_02675_));
 sg13g2_a221oi_1 _17297_ (.B2(_02668_),
    .C1(_02675_),
    .B1(net3903),
    .A1(_03505_),
    .Y(_02676_),
    .A2(net3744));
 sg13g2_nand2_1 _17298_ (.Y(_02677_),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ),
    .B(_02676_));
 sg13g2_o21ai_1 _17299_ (.B1(net3916),
    .Y(_02678_),
    .A1(_00127_),
    .A2(net3909));
 sg13g2_a221oi_1 _17300_ (.B2(_03504_),
    .C1(_02678_),
    .B1(net3901),
    .A1(_03505_),
    .Y(_02679_),
    .A2(net3738));
 sg13g2_a21oi_1 _17301_ (.A1(_00131_),
    .A2(net3744),
    .Y(_02680_),
    .B1(_02679_));
 sg13g2_and2_1 _17302_ (.A(_00130_),
    .B(_02680_),
    .X(_02681_));
 sg13g2_xnor2_1 _17303_ (.Y(_02682_),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ),
    .B(_02676_));
 sg13g2_o21ai_1 _17304_ (.B1(_02677_),
    .Y(_02683_),
    .A1(_02681_),
    .A2(_02682_));
 sg13g2_xnor2_1 _17305_ (.Y(_02684_),
    .A(_03505_),
    .B(_02674_));
 sg13g2_nor2b_1 _17306_ (.A(_02684_),
    .B_N(_02683_),
    .Y(_02685_));
 sg13g2_a21o_1 _17307_ (.A2(_02674_),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ),
    .B1(_02685_),
    .X(_02686_));
 sg13g2_xnor2_1 _17308_ (.Y(_02687_),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ),
    .B(_02671_));
 sg13g2_a21oi_1 _17309_ (.A1(_02686_),
    .A2(_02687_),
    .Y(_02688_),
    .B1(_02672_));
 sg13g2_nor2b_1 _17310_ (.A(_02669_),
    .B_N(_02688_),
    .Y(_02689_));
 sg13g2_a22oi_1 _17311_ (.Y(_02690_),
    .B1(_02670_),
    .B2(_02689_),
    .A2(_02669_),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ));
 sg13g2_inv_1 _17312_ (.Y(_02691_),
    .A(_02690_));
 sg13g2_mux2_2 _17313_ (.A0(net4492),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[515] ),
    .X(_02692_));
 sg13g2_nand2_1 _17314_ (.Y(_02693_),
    .A(\spiking_network_top_uut.all_data_out[129] ),
    .B(_02692_));
 sg13g2_mux2_2 _17315_ (.A0(net4491),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[519] ),
    .X(_02694_));
 sg13g2_nand2_1 _17316_ (.Y(_02695_),
    .A(\spiking_network_top_uut.all_data_out[131] ),
    .B(_02694_));
 sg13g2_nor2_1 _17317_ (.A(_02693_),
    .B(_02695_),
    .Y(_02696_));
 sg13g2_nand4_1 _17318_ (.B(\spiking_network_top_uut.all_data_out[130] ),
    .C(_02692_),
    .A(\spiking_network_top_uut.all_data_out[128] ),
    .Y(_02697_),
    .D(_02694_));
 sg13g2_inv_1 _17319_ (.Y(_02698_),
    .A(_02697_));
 sg13g2_xor2_1 _17320_ (.B(_02695_),
    .A(_02693_),
    .X(_02699_));
 sg13g2_a21oi_2 _17321_ (.B1(_02696_),
    .Y(_02700_),
    .A2(_02699_),
    .A1(_02697_));
 sg13g2_mux2_2 _17322_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.din ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[527] ),
    .X(_02701_));
 sg13g2_nand2_1 _17323_ (.Y(_02702_),
    .A(\spiking_network_top_uut.all_data_out[135] ),
    .B(_02701_));
 sg13g2_mux2_2 _17324_ (.A0(net4490),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[523] ),
    .X(_02703_));
 sg13g2_nand2_1 _17325_ (.Y(_02704_),
    .A(\spiking_network_top_uut.all_data_out[133] ),
    .B(_02703_));
 sg13g2_nor2_1 _17326_ (.A(_02702_),
    .B(_02704_),
    .Y(_02705_));
 sg13g2_nand2_1 _17327_ (.Y(_02706_),
    .A(\spiking_network_top_uut.all_data_out[134] ),
    .B(_02701_));
 sg13g2_nand2_1 _17328_ (.Y(_02707_),
    .A(\spiking_network_top_uut.all_data_out[132] ),
    .B(_02703_));
 sg13g2_or2_2 _17329_ (.X(_02708_),
    .B(_02707_),
    .A(_02706_));
 sg13g2_xor2_1 _17330_ (.B(_02704_),
    .A(_02702_),
    .X(_02709_));
 sg13g2_a21oi_2 _17331_ (.B1(_02705_),
    .Y(_02710_),
    .A2(_02709_),
    .A1(_02708_));
 sg13g2_mux2_2 _17332_ (.A0(net4487),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[535] ),
    .X(_02711_));
 sg13g2_mux2_2 _17333_ (.A0(net4488),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[531] ),
    .X(_02712_));
 sg13g2_a22oi_1 _17334_ (.Y(_02713_),
    .B1(_02712_),
    .B2(\spiking_network_top_uut.all_data_out[137] ),
    .A2(_02711_),
    .A1(\spiking_network_top_uut.all_data_out[139] ));
 sg13g2_and4_1 _17335_ (.A(\spiking_network_top_uut.all_data_out[139] ),
    .B(\spiking_network_top_uut.all_data_out[137] ),
    .C(_02711_),
    .D(_02712_),
    .X(_02714_));
 sg13g2_nand4_1 _17336_ (.B(\spiking_network_top_uut.all_data_out[137] ),
    .C(_02711_),
    .A(\spiking_network_top_uut.all_data_out[139] ),
    .Y(_02715_),
    .D(_02712_));
 sg13g2_and4_2 _17337_ (.A(\spiking_network_top_uut.all_data_out[138] ),
    .B(\spiking_network_top_uut.all_data_out[136] ),
    .C(_02711_),
    .D(_02712_),
    .X(_02716_));
 sg13g2_a21oi_2 _17338_ (.B1(_02713_),
    .Y(_02717_),
    .A2(_02716_),
    .A1(_02715_));
 sg13g2_mux2_2 _17339_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.din ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[543] ),
    .X(_02718_));
 sg13g2_mux2_2 _17340_ (.A0(net4486),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[539] ),
    .X(_02719_));
 sg13g2_and4_1 _17341_ (.A(\spiking_network_top_uut.all_data_out[143] ),
    .B(\spiking_network_top_uut.all_data_out[141] ),
    .C(_02718_),
    .D(_02719_),
    .X(_02720_));
 sg13g2_nand4_1 _17342_ (.B(\spiking_network_top_uut.all_data_out[141] ),
    .C(_02718_),
    .A(\spiking_network_top_uut.all_data_out[143] ),
    .Y(_02721_),
    .D(_02719_));
 sg13g2_and4_1 _17343_ (.A(\spiking_network_top_uut.all_data_out[142] ),
    .B(\spiking_network_top_uut.all_data_out[140] ),
    .C(_02718_),
    .D(_02719_),
    .X(_02722_));
 sg13g2_a22oi_1 _17344_ (.Y(_02723_),
    .B1(_02719_),
    .B2(\spiking_network_top_uut.all_data_out[141] ),
    .A2(_02718_),
    .A1(\spiking_network_top_uut.all_data_out[143] ));
 sg13g2_or3_1 _17345_ (.A(_02720_),
    .B(_02722_),
    .C(_02723_),
    .X(_02724_));
 sg13g2_o21ai_1 _17346_ (.B1(_02721_),
    .Y(_02725_),
    .A1(_02722_),
    .A2(_02723_));
 sg13g2_nand3b_1 _17347_ (.B(_02717_),
    .C(_02725_),
    .Y(_02726_),
    .A_N(_02710_));
 sg13g2_inv_1 _17348_ (.Y(_02727_),
    .A(_02726_));
 sg13g2_or2_1 _17349_ (.X(_02728_),
    .B(_02726_),
    .A(_02700_));
 sg13g2_inv_1 _17350_ (.Y(_02729_),
    .A(_02728_));
 sg13g2_nor2_1 _17351_ (.A(_02717_),
    .B(_02725_),
    .Y(_02730_));
 sg13g2_and2_2 _17352_ (.A(_02710_),
    .B(_02730_),
    .X(_02731_));
 sg13g2_a21oi_2 _17353_ (.B1(_02729_),
    .Y(_02732_),
    .A2(_02731_),
    .A1(_02700_));
 sg13g2_xor2_1 _17354_ (.B(_02688_),
    .A(_02669_),
    .X(_02733_));
 sg13g2_a21o_1 _17355_ (.A2(_02733_),
    .A1(_02732_),
    .B1(_02729_),
    .X(_02734_));
 sg13g2_xor2_1 _17356_ (.B(_02732_),
    .A(_02690_),
    .X(_02735_));
 sg13g2_nor2b_1 _17357_ (.A(_02735_),
    .B_N(_02734_),
    .Y(_02736_));
 sg13g2_xnor2_1 _17358_ (.Y(_02737_),
    .A(_02734_),
    .B(_02735_));
 sg13g2_o21ai_1 _17359_ (.B1(_02722_),
    .Y(_02738_),
    .A1(_02720_),
    .A2(_02723_));
 sg13g2_o21ai_1 _17360_ (.B1(_02716_),
    .Y(_02739_),
    .A1(_02713_),
    .A2(_02714_));
 sg13g2_or3_1 _17361_ (.A(_02713_),
    .B(_02714_),
    .C(_02716_),
    .X(_02740_));
 sg13g2_a22oi_1 _17362_ (.Y(_02741_),
    .B1(_02739_),
    .B2(_02740_),
    .A2(_02738_),
    .A1(_02724_));
 sg13g2_xor2_1 _17363_ (.B(_02709_),
    .A(_02708_),
    .X(_02742_));
 sg13g2_xnor2_1 _17364_ (.Y(_02743_),
    .A(_02708_),
    .B(_02709_));
 sg13g2_and4_1 _17365_ (.A(_02724_),
    .B(_02738_),
    .C(_02739_),
    .D(_02740_),
    .X(_02744_));
 sg13g2_nand4_1 _17366_ (.B(_02738_),
    .C(_02739_),
    .A(_02724_),
    .Y(_02745_),
    .D(_02740_));
 sg13g2_nand3b_1 _17367_ (.B(_02743_),
    .C(_02745_),
    .Y(_02746_),
    .A_N(_02741_));
 sg13g2_a21oi_2 _17368_ (.B1(_02741_),
    .Y(_02747_),
    .A2(_02745_),
    .A1(_02743_));
 sg13g2_xor2_1 _17369_ (.B(_02725_),
    .A(_02717_),
    .X(_02748_));
 sg13g2_xnor2_1 _17370_ (.Y(_02749_),
    .A(_02710_),
    .B(_02748_));
 sg13g2_nor2b_1 _17371_ (.A(_02747_),
    .B_N(_02749_),
    .Y(_02750_));
 sg13g2_xnor2_1 _17372_ (.Y(_02751_),
    .A(_02747_),
    .B(_02749_));
 sg13g2_nor2b_1 _17373_ (.A(_02700_),
    .B_N(_02751_),
    .Y(_02752_));
 sg13g2_nor2_2 _17374_ (.A(_02750_),
    .B(_02752_),
    .Y(_02753_));
 sg13g2_nor2_1 _17375_ (.A(_02727_),
    .B(_02731_),
    .Y(_02754_));
 sg13g2_xnor2_1 _17376_ (.Y(_02755_),
    .A(_02700_),
    .B(_02754_));
 sg13g2_nor2b_1 _17377_ (.A(_02753_),
    .B_N(_02755_),
    .Y(_02756_));
 sg13g2_xnor2_1 _17378_ (.Y(_02757_),
    .A(_02753_),
    .B(_02755_));
 sg13g2_xor2_1 _17379_ (.B(_02687_),
    .A(_02686_),
    .X(_02758_));
 sg13g2_a21oi_1 _17380_ (.A1(_02757_),
    .A2(_02758_),
    .Y(_02759_),
    .B1(_02756_));
 sg13g2_xor2_1 _17381_ (.B(_02733_),
    .A(_02732_),
    .X(_02760_));
 sg13g2_nor2b_1 _17382_ (.A(_02759_),
    .B_N(_02760_),
    .Y(_02761_));
 sg13g2_xnor2_1 _17383_ (.Y(_02762_),
    .A(_02757_),
    .B(_02758_));
 sg13g2_a22oi_1 _17384_ (.Y(_02763_),
    .B1(_02719_),
    .B2(\spiking_network_top_uut.all_data_out[140] ),
    .A2(_02718_),
    .A1(\spiking_network_top_uut.all_data_out[142] ));
 sg13g2_nor2_1 _17385_ (.A(_02722_),
    .B(_02763_),
    .Y(_02764_));
 sg13g2_a22oi_1 _17386_ (.Y(_02765_),
    .B1(_02712_),
    .B2(\spiking_network_top_uut.all_data_out[136] ),
    .A2(_02711_),
    .A1(\spiking_network_top_uut.all_data_out[138] ));
 sg13g2_nor2_1 _17387_ (.A(_02716_),
    .B(_02765_),
    .Y(_02766_));
 sg13g2_and2_1 _17388_ (.A(_02764_),
    .B(_02766_),
    .X(_02767_));
 sg13g2_xor2_1 _17389_ (.B(_02707_),
    .A(_02706_),
    .X(_02768_));
 sg13g2_xor2_1 _17390_ (.B(_02766_),
    .A(_02764_),
    .X(_02769_));
 sg13g2_a21o_1 _17391_ (.A2(_02769_),
    .A1(_02768_),
    .B1(_02767_),
    .X(_02770_));
 sg13g2_o21ai_1 _17392_ (.B1(_02742_),
    .Y(_02771_),
    .A1(_02741_),
    .A2(_02744_));
 sg13g2_and3_1 _17393_ (.X(_02772_),
    .A(_02746_),
    .B(_02770_),
    .C(_02771_));
 sg13g2_nand3_1 _17394_ (.B(_02770_),
    .C(_02771_),
    .A(_02746_),
    .Y(_02773_));
 sg13g2_xnor2_1 _17395_ (.Y(_02774_),
    .A(_02698_),
    .B(_02699_));
 sg13g2_a21oi_1 _17396_ (.A1(_02746_),
    .A2(_02771_),
    .Y(_02775_),
    .B1(_02770_));
 sg13g2_or3_2 _17397_ (.A(_02772_),
    .B(_02774_),
    .C(_02775_),
    .X(_02776_));
 sg13g2_o21ai_1 _17398_ (.B1(_02773_),
    .Y(_02777_),
    .A1(_02774_),
    .A2(_02775_));
 sg13g2_xnor2_1 _17399_ (.Y(_02778_),
    .A(_02700_),
    .B(_02751_));
 sg13g2_nand2_1 _17400_ (.Y(_02779_),
    .A(_02777_),
    .B(_02778_));
 sg13g2_xnor2_1 _17401_ (.Y(_02780_),
    .A(_02777_),
    .B(_02778_));
 sg13g2_xor2_1 _17402_ (.B(_02684_),
    .A(_02683_),
    .X(_02781_));
 sg13g2_o21ai_1 _17403_ (.B1(_02779_),
    .Y(_02782_),
    .A1(_02780_),
    .A2(_02781_));
 sg13g2_nand2b_1 _17404_ (.Y(_02783_),
    .B(_02782_),
    .A_N(_02762_));
 sg13g2_a22oi_1 _17405_ (.Y(_02784_),
    .B1(_02694_),
    .B2(\spiking_network_top_uut.all_data_out[130] ),
    .A2(_02692_),
    .A1(\spiking_network_top_uut.all_data_out[128] ));
 sg13g2_nor2_2 _17406_ (.A(_02698_),
    .B(_02784_),
    .Y(_02785_));
 sg13g2_inv_1 _17407_ (.Y(_02786_),
    .A(_02785_));
 sg13g2_xnor2_1 _17408_ (.Y(_02787_),
    .A(_02768_),
    .B(_02769_));
 sg13g2_nor2_1 _17409_ (.A(_02786_),
    .B(_02787_),
    .Y(_02788_));
 sg13g2_o21ai_1 _17410_ (.B1(_02774_),
    .Y(_02789_),
    .A1(_02772_),
    .A2(_02775_));
 sg13g2_nand3_1 _17411_ (.B(_02788_),
    .C(_02789_),
    .A(_02776_),
    .Y(_02790_));
 sg13g2_a21oi_2 _17412_ (.B1(_02788_),
    .Y(_02791_),
    .A2(_02789_),
    .A1(_02776_));
 sg13g2_a21o_2 _17413_ (.A2(_02789_),
    .A1(_02776_),
    .B1(_02788_),
    .X(_02792_));
 sg13g2_xnor2_1 _17414_ (.Y(_02793_),
    .A(_02681_),
    .B(_02682_));
 sg13g2_inv_1 _17415_ (.Y(_02794_),
    .A(_02793_));
 sg13g2_and3_1 _17416_ (.X(_02795_),
    .A(_02790_),
    .B(_02792_),
    .C(_02794_));
 sg13g2_o21ai_1 _17417_ (.B1(_02790_),
    .Y(_02796_),
    .A1(_02791_),
    .A2(_02793_));
 sg13g2_xor2_1 _17418_ (.B(_02781_),
    .A(_02780_),
    .X(_02797_));
 sg13g2_and2_1 _17419_ (.A(_02796_),
    .B(_02797_),
    .X(_02798_));
 sg13g2_a21oi_1 _17420_ (.A1(_02790_),
    .A2(_02792_),
    .Y(_02799_),
    .B1(_02794_));
 sg13g2_xnor2_1 _17421_ (.Y(_02800_),
    .A(_02786_),
    .B(_02787_));
 sg13g2_xnor2_1 _17422_ (.Y(_02801_),
    .A(_00130_),
    .B(_02680_));
 sg13g2_nand2b_1 _17423_ (.Y(_02802_),
    .B(_02801_),
    .A_N(_02800_));
 sg13g2_nor3_2 _17424_ (.A(_02795_),
    .B(_02799_),
    .C(_02802_),
    .Y(_02803_));
 sg13g2_or2_1 _17425_ (.X(_02804_),
    .B(_02797_),
    .A(_02796_));
 sg13g2_nand2b_1 _17426_ (.Y(_02805_),
    .B(_02804_),
    .A_N(_02798_));
 sg13g2_a21oi_1 _17427_ (.A1(_02803_),
    .A2(_02804_),
    .Y(_02806_),
    .B1(_02798_));
 sg13g2_xor2_1 _17428_ (.B(_02782_),
    .A(_02762_),
    .X(_02807_));
 sg13g2_o21ai_1 _17429_ (.B1(_02783_),
    .Y(_02808_),
    .A1(_02806_),
    .A2(_02807_));
 sg13g2_xnor2_1 _17430_ (.Y(_02809_),
    .A(_02759_),
    .B(_02760_));
 sg13g2_a21o_1 _17431_ (.A2(_02809_),
    .A1(_02808_),
    .B1(_02761_),
    .X(_02810_));
 sg13g2_a21oi_1 _17432_ (.A1(_02737_),
    .A2(_02810_),
    .Y(_02811_),
    .B1(_02736_));
 sg13g2_nand3_1 _17433_ (.B(_02700_),
    .C(_02731_),
    .A(_02690_),
    .Y(_02812_));
 sg13g2_a221oi_1 _17434_ (.B2(_02812_),
    .C1(_02647_),
    .B1(_02811_),
    .A1(_02691_),
    .Y(_02813_),
    .A2(_02729_));
 sg13g2_a21oi_2 _17435_ (.B1(_02813_),
    .Y(_02814_),
    .A2(_02690_),
    .A1(_02647_));
 sg13g2_xor2_1 _17436_ (.B(_02810_),
    .A(_02737_),
    .X(_02815_));
 sg13g2_mux2_1 _17437_ (.A0(_02691_),
    .A1(_02815_),
    .S(_02646_),
    .X(_02816_));
 sg13g2_nand2_1 _17438_ (.Y(_02817_),
    .A(_02647_),
    .B(_02733_));
 sg13g2_xnor2_1 _17439_ (.Y(_02818_),
    .A(_02808_),
    .B(_02809_));
 sg13g2_o21ai_1 _17440_ (.B1(_02817_),
    .Y(_02819_),
    .A1(_02647_),
    .A2(_02818_));
 sg13g2_nand2_1 _17441_ (.Y(_02820_),
    .A(_02816_),
    .B(_02819_));
 sg13g2_a21oi_2 _17442_ (.B1(net3639),
    .Y(_02821_),
    .A2(_02820_),
    .A1(_02814_));
 sg13g2_nor2_1 _17443_ (.A(_02816_),
    .B(_02819_),
    .Y(_02822_));
 sg13g2_nor2_2 _17444_ (.A(_02814_),
    .B(_02822_),
    .Y(_02823_));
 sg13g2_nor2_1 _17445_ (.A(_02647_),
    .B(_02800_),
    .Y(_02824_));
 sg13g2_xor2_1 _17446_ (.B(_02824_),
    .A(_02801_),
    .X(_02825_));
 sg13g2_o21ai_1 _17447_ (.B1(_02821_),
    .Y(_02826_),
    .A1(_02823_),
    .A2(_02825_));
 sg13g2_xor2_1 _17448_ (.B(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[0] ),
    .A(net4313),
    .X(_02827_));
 sg13g2_a21oi_1 _17449_ (.A1(net3639),
    .A2(_02827_),
    .Y(_02828_),
    .B1(net3948));
 sg13g2_a22oi_1 _17450_ (.Y(_00998_),
    .B1(_02826_),
    .B2(_02828_),
    .A2(_03465_),
    .A1(net3948));
 sg13g2_o21ai_1 _17451_ (.B1(_02802_),
    .Y(_02829_),
    .A1(_02795_),
    .A2(_02799_));
 sg13g2_nand3b_1 _17452_ (.B(_02829_),
    .C(_02646_),
    .Y(_02830_),
    .A_N(_02803_));
 sg13g2_o21ai_1 _17453_ (.B1(_02830_),
    .Y(_02831_),
    .A1(_02646_),
    .A2(_02793_));
 sg13g2_o21ai_1 _17454_ (.B1(_02821_),
    .Y(_02832_),
    .A1(_02823_),
    .A2(_02831_));
 sg13g2_xor2_1 _17455_ (.B(_04945_),
    .A(_04944_),
    .X(_02833_));
 sg13g2_a21oi_1 _17456_ (.A1(net3639),
    .A2(_02833_),
    .Y(_02834_),
    .B1(net3949));
 sg13g2_a22oi_1 _17457_ (.Y(_00999_),
    .B1(_02832_),
    .B2(_02834_),
    .A2(_03464_),
    .A1(net3948));
 sg13g2_xnor2_1 _17458_ (.Y(_02835_),
    .A(_02803_),
    .B(_02805_));
 sg13g2_nand2_1 _17459_ (.Y(_02836_),
    .A(_02646_),
    .B(_02835_));
 sg13g2_o21ai_1 _17460_ (.B1(_02836_),
    .Y(_02837_),
    .A1(_02646_),
    .A2(_02781_));
 sg13g2_nor2_1 _17461_ (.A(_02823_),
    .B(_02837_),
    .Y(_02838_));
 sg13g2_nand2_1 _17462_ (.Y(_02839_),
    .A(net4603),
    .B(_02821_));
 sg13g2_xor2_1 _17463_ (.B(_04947_),
    .A(_04946_),
    .X(_02840_));
 sg13g2_a22oi_1 _17464_ (.Y(_02841_),
    .B1(_00007_),
    .B2(_02840_),
    .A2(net519),
    .A1(net3948));
 sg13g2_o21ai_1 _17465_ (.B1(_02841_),
    .Y(_01000_),
    .A1(_02838_),
    .A2(_02839_));
 sg13g2_nor2_1 _17466_ (.A(_02646_),
    .B(_02758_),
    .Y(_02842_));
 sg13g2_xnor2_1 _17467_ (.Y(_02843_),
    .A(_02806_),
    .B(_02807_));
 sg13g2_a21oi_1 _17468_ (.A1(_02646_),
    .A2(_02843_),
    .Y(_02844_),
    .B1(_02842_));
 sg13g2_o21ai_1 _17469_ (.B1(_02821_),
    .Y(_02845_),
    .A1(_02823_),
    .A2(_02844_));
 sg13g2_or3_1 _17470_ (.A(_04941_),
    .B(_04942_),
    .C(_04948_),
    .X(_02846_));
 sg13g2_and2_1 _17471_ (.A(_04949_),
    .B(_02846_),
    .X(_02847_));
 sg13g2_a21oi_1 _17472_ (.A1(net3639),
    .A2(_02847_),
    .Y(_02848_),
    .B1(net3947));
 sg13g2_a22oi_1 _17473_ (.Y(_01001_),
    .B1(_02845_),
    .B2(_02848_),
    .A2(_03463_),
    .A1(net3948));
 sg13g2_o21ai_1 _17474_ (.B1(net4603),
    .Y(_02849_),
    .A1(_04939_),
    .A2(_04950_));
 sg13g2_a21oi_1 _17475_ (.A1(_04952_),
    .A2(_02814_),
    .Y(_02850_),
    .B1(_02849_));
 sg13g2_a21oi_1 _17476_ (.A1(net3948),
    .A2(_03462_),
    .Y(_01002_),
    .B1(_02850_));
 sg13g2_mux4_1 _17477_ (.S0(\spiking_network_top_uut.all_data_out[572] ),
    .A0(net3789),
    .A1(net3788),
    .A2(net3787),
    .A3(net3786),
    .S1(\spiking_network_top_uut.all_data_out[573] ),
    .X(_02851_));
 sg13g2_mux2_1 _17478_ (.A0(net3783),
    .A1(net3899),
    .S(\spiking_network_top_uut.all_data_out[572] ),
    .X(_02852_));
 sg13g2_nor2b_1 _17479_ (.A(\spiking_network_top_uut.all_data_out[572] ),
    .B_N(net3785),
    .Y(_02853_));
 sg13g2_a21oi_1 _17480_ (.A1(\spiking_network_top_uut.all_data_out[572] ),
    .A2(net3784),
    .Y(_02854_),
    .B1(_02853_));
 sg13g2_o21ai_1 _17481_ (.B1(\spiking_network_top_uut.all_data_out[574] ),
    .Y(_02855_),
    .A1(\spiking_network_top_uut.all_data_out[573] ),
    .A2(_02854_));
 sg13g2_a21oi_1 _17482_ (.A1(\spiking_network_top_uut.all_data_out[573] ),
    .A2(_02852_),
    .Y(_02856_),
    .B1(_02855_));
 sg13g2_o21ai_1 _17483_ (.B1(net4638),
    .Y(_02857_),
    .A1(\spiking_network_top_uut.all_data_out[574] ),
    .A2(_02851_));
 sg13g2_nand2_1 _17484_ (.Y(_02858_),
    .A(net3962),
    .B(net246));
 sg13g2_o21ai_1 _17485_ (.B1(_02858_),
    .Y(_01003_),
    .A1(_02856_),
    .A2(_02857_));
 sg13g2_mux2_1 _17486_ (.A0(net3840),
    .A1(net4486),
    .S(net4636),
    .X(_01004_));
 sg13g2_mux2_1 _17487_ (.A0(net3839),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[0] ),
    .S(net4641),
    .X(_01005_));
 sg13g2_mux2_1 _17488_ (.A0(net3838),
    .A1(net3839),
    .S(net4640),
    .X(_01006_));
 sg13g2_mux2_1 _17489_ (.A0(net3837),
    .A1(net3838),
    .S(net4640),
    .X(_01007_));
 sg13g2_mux2_1 _17490_ (.A0(net3836),
    .A1(net3837),
    .S(net4643),
    .X(_01008_));
 sg13g2_nand2_1 _17491_ (.Y(_02859_),
    .A(net4642),
    .B(net3836));
 sg13g2_o21ai_1 _17492_ (.B1(_02859_),
    .Y(_01009_),
    .A1(net4642),
    .A2(_03662_));
 sg13g2_nor2_1 _17493_ (.A(net4642),
    .B(net3835),
    .Y(_02860_));
 sg13g2_a21oi_1 _17494_ (.A1(net4642),
    .A2(_03662_),
    .Y(_01010_),
    .B1(_02860_));
 sg13g2_mux2_1 _17495_ (.A0(net3834),
    .A1(net3835),
    .S(net4641),
    .X(_01011_));
 sg13g2_mux2_1 _17496_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_dout ),
    .A1(net246),
    .S(net4639),
    .X(_01012_));
 sg13g2_mux4_1 _17497_ (.S0(\spiking_network_top_uut.all_data_out[568] ),
    .A0(net3840),
    .A1(net3839),
    .A2(net3838),
    .A3(net3837),
    .S1(\spiking_network_top_uut.all_data_out[569] ),
    .X(_02861_));
 sg13g2_mux2_1 _17498_ (.A0(net3835),
    .A1(net3834),
    .S(\spiking_network_top_uut.all_data_out[568] ),
    .X(_02862_));
 sg13g2_nor2b_1 _17499_ (.A(\spiking_network_top_uut.all_data_out[568] ),
    .B_N(net3836),
    .Y(_02863_));
 sg13g2_a21oi_1 _17500_ (.A1(\spiking_network_top_uut.all_data_out[568] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[5] ),
    .Y(_02864_),
    .B1(_02863_));
 sg13g2_o21ai_1 _17501_ (.B1(\spiking_network_top_uut.all_data_out[570] ),
    .Y(_02865_),
    .A1(\spiking_network_top_uut.all_data_out[569] ),
    .A2(_02864_));
 sg13g2_a21oi_1 _17502_ (.A1(\spiking_network_top_uut.all_data_out[569] ),
    .A2(_02862_),
    .Y(_02866_),
    .B1(_02865_));
 sg13g2_o21ai_1 _17503_ (.B1(net4641),
    .Y(_02867_),
    .A1(\spiking_network_top_uut.all_data_out[570] ),
    .A2(_02861_));
 sg13g2_nand2_1 _17504_ (.Y(_02868_),
    .A(net3963),
    .B(net47));
 sg13g2_o21ai_1 _17505_ (.B1(_02868_),
    .Y(_01013_),
    .A1(_02866_),
    .A2(_02867_));
 sg13g2_mux2_1 _17506_ (.A0(net3833),
    .A1(net4487),
    .S(net4607),
    .X(_01014_));
 sg13g2_mux2_1 _17507_ (.A0(net3832),
    .A1(net3833),
    .S(net4609),
    .X(_01015_));
 sg13g2_mux2_1 _17508_ (.A0(net3831),
    .A1(net3832),
    .S(net4609),
    .X(_01016_));
 sg13g2_mux2_1 _17509_ (.A0(net3830),
    .A1(net3831),
    .S(net4610),
    .X(_01017_));
 sg13g2_mux2_1 _17510_ (.A0(net3829),
    .A1(net3830),
    .S(net4609),
    .X(_01018_));
 sg13g2_nand2_1 _17511_ (.Y(_02869_),
    .A(net4607),
    .B(net3829));
 sg13g2_o21ai_1 _17512_ (.B1(_02869_),
    .Y(_01019_),
    .A1(net4607),
    .A2(_03661_));
 sg13g2_nor2_1 _17513_ (.A(net4607),
    .B(net3828),
    .Y(_02870_));
 sg13g2_a21oi_1 _17514_ (.A1(net4607),
    .A2(_03661_),
    .Y(_01020_),
    .B1(_02870_));
 sg13g2_mux2_1 _17515_ (.A0(net3827),
    .A1(net3828),
    .S(net4609),
    .X(_01021_));
 sg13g2_mux2_1 _17516_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_dout ),
    .A1(net47),
    .S(net4636),
    .X(_01022_));
 sg13g2_mux4_1 _17517_ (.S0(\spiking_network_top_uut.all_data_out[564] ),
    .A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[0] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[1] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[2] ),
    .A3(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[3] ),
    .S1(\spiking_network_top_uut.all_data_out[565] ),
    .X(_02871_));
 sg13g2_mux2_1 _17518_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[6] ),
    .A1(net3827),
    .S(\spiking_network_top_uut.all_data_out[564] ),
    .X(_02872_));
 sg13g2_nor2b_1 _17519_ (.A(\spiking_network_top_uut.all_data_out[564] ),
    .B_N(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[4] ),
    .Y(_02873_));
 sg13g2_a21oi_1 _17520_ (.A1(\spiking_network_top_uut.all_data_out[564] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[5] ),
    .Y(_02874_),
    .B1(_02873_));
 sg13g2_o21ai_1 _17521_ (.B1(\spiking_network_top_uut.all_data_out[566] ),
    .Y(_02875_),
    .A1(\spiking_network_top_uut.all_data_out[565] ),
    .A2(_02874_));
 sg13g2_a21oi_1 _17522_ (.A1(\spiking_network_top_uut.all_data_out[565] ),
    .A2(_02872_),
    .Y(_02876_),
    .B1(_02875_));
 sg13g2_o21ai_1 _17523_ (.B1(net4609),
    .Y(_02877_),
    .A1(\spiking_network_top_uut.all_data_out[566] ),
    .A2(_02871_));
 sg13g2_nand2_1 _17524_ (.Y(_02878_),
    .A(net3966),
    .B(net369));
 sg13g2_o21ai_1 _17525_ (.B1(_02878_),
    .Y(_01023_),
    .A1(_02876_),
    .A2(_02877_));
 sg13g2_mux2_1 _17526_ (.A0(net3826),
    .A1(net4488),
    .S(net4613),
    .X(_01024_));
 sg13g2_mux2_1 _17527_ (.A0(net3825),
    .A1(net3826),
    .S(net4614),
    .X(_01025_));
 sg13g2_mux2_1 _17528_ (.A0(net3824),
    .A1(net3825),
    .S(net4614),
    .X(_01026_));
 sg13g2_mux2_1 _17529_ (.A0(net3823),
    .A1(net3824),
    .S(net4620),
    .X(_01027_));
 sg13g2_mux2_1 _17530_ (.A0(net3822),
    .A1(net3823),
    .S(net4620),
    .X(_01028_));
 sg13g2_nand2_1 _17531_ (.Y(_02879_),
    .A(net4613),
    .B(net3822));
 sg13g2_o21ai_1 _17532_ (.B1(_02879_),
    .Y(_01029_),
    .A1(net4613),
    .A2(_03660_));
 sg13g2_nor2_1 _17533_ (.A(net4614),
    .B(net3821),
    .Y(_02880_));
 sg13g2_a21oi_1 _17534_ (.A1(net4614),
    .A2(_03660_),
    .Y(_01030_),
    .B1(_02880_));
 sg13g2_mux2_1 _17535_ (.A0(net3820),
    .A1(net3821),
    .S(net4614),
    .X(_01031_));
 sg13g2_mux2_1 _17536_ (.A0(net271),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_reg1 ),
    .S(net4612),
    .X(_01032_));
 sg13g2_a21oi_1 _17537_ (.A1(\spiking_network_top_uut.all_data_out[560] ),
    .A2(_03660_),
    .Y(_02881_),
    .B1(\spiking_network_top_uut.all_data_out[561] ));
 sg13g2_o21ai_1 _17538_ (.B1(_02881_),
    .Y(_02882_),
    .A1(\spiking_network_top_uut.all_data_out[560] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[4] ));
 sg13g2_mux2_1 _17539_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[6] ),
    .A1(net3820),
    .S(\spiking_network_top_uut.all_data_out[560] ),
    .X(_02883_));
 sg13g2_nand2_1 _17540_ (.Y(_02884_),
    .A(\spiking_network_top_uut.all_data_out[561] ),
    .B(_02883_));
 sg13g2_nand3_1 _17541_ (.B(_02882_),
    .C(_02884_),
    .A(\spiking_network_top_uut.all_data_out[562] ),
    .Y(_02885_));
 sg13g2_mux2_1 _17542_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[2] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[3] ),
    .S(\spiking_network_top_uut.all_data_out[560] ),
    .X(_02886_));
 sg13g2_nor2b_1 _17543_ (.A(\spiking_network_top_uut.all_data_out[560] ),
    .B_N(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[0] ),
    .Y(_02887_));
 sg13g2_a21oi_1 _17544_ (.A1(\spiking_network_top_uut.all_data_out[560] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[1] ),
    .Y(_02888_),
    .B1(_02887_));
 sg13g2_a21oi_1 _17545_ (.A1(\spiking_network_top_uut.all_data_out[561] ),
    .A2(_02886_),
    .Y(_02889_),
    .B1(\spiking_network_top_uut.all_data_out[562] ));
 sg13g2_o21ai_1 _17546_ (.B1(_02889_),
    .Y(_02890_),
    .A1(\spiking_network_top_uut.all_data_out[561] ),
    .A2(_02888_));
 sg13g2_nand3_1 _17547_ (.B(_02885_),
    .C(_02890_),
    .A(net4615),
    .Y(_02891_));
 sg13g2_o21ai_1 _17548_ (.B1(_02891_),
    .Y(_01033_),
    .A1(net4620),
    .A2(_03691_));
 sg13g2_mux2_1 _17549_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[0] ),
    .A1(net4489),
    .S(net4626),
    .X(_01034_));
 sg13g2_mux2_1 _17550_ (.A0(net3818),
    .A1(net3819),
    .S(net4625),
    .X(_01035_));
 sg13g2_mux2_1 _17551_ (.A0(net3817),
    .A1(net3818),
    .S(net4625),
    .X(_01036_));
 sg13g2_mux2_1 _17552_ (.A0(net3816),
    .A1(net3817),
    .S(net4625),
    .X(_01037_));
 sg13g2_mux2_1 _17553_ (.A0(net3815),
    .A1(net3816),
    .S(net4626),
    .X(_01038_));
 sg13g2_nand2_1 _17554_ (.Y(_02892_),
    .A(net4625),
    .B(net3815));
 sg13g2_o21ai_1 _17555_ (.B1(_02892_),
    .Y(_01039_),
    .A1(net4625),
    .A2(_03659_));
 sg13g2_nor2_1 _17556_ (.A(net4626),
    .B(net3814),
    .Y(_02893_));
 sg13g2_a21oi_1 _17557_ (.A1(net4626),
    .A2(_03659_),
    .Y(_01040_),
    .B1(_02893_));
 sg13g2_mux2_1 _17558_ (.A0(net3813),
    .A1(net3814),
    .S(net4625),
    .X(_01041_));
 sg13g2_nor2_1 _17559_ (.A(net4620),
    .B(net111),
    .Y(_02894_));
 sg13g2_a21oi_1 _17560_ (.A1(net4620),
    .A2(_03691_),
    .Y(_01042_),
    .B1(_02894_));
 sg13g2_mux2_1 _17561_ (.A0(net3817),
    .A1(net3816),
    .S(\spiking_network_top_uut.all_data_out[556] ),
    .X(_02895_));
 sg13g2_nor2b_1 _17562_ (.A(\spiking_network_top_uut.all_data_out[556] ),
    .B_N(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[0] ),
    .Y(_02896_));
 sg13g2_a21oi_1 _17563_ (.A1(\spiking_network_top_uut.all_data_out[556] ),
    .A2(net3818),
    .Y(_02897_),
    .B1(_02896_));
 sg13g2_a21oi_1 _17564_ (.A1(\spiking_network_top_uut.all_data_out[557] ),
    .A2(_02895_),
    .Y(_02898_),
    .B1(\spiking_network_top_uut.all_data_out[558] ));
 sg13g2_o21ai_1 _17565_ (.B1(_02898_),
    .Y(_02899_),
    .A1(\spiking_network_top_uut.all_data_out[557] ),
    .A2(_02897_));
 sg13g2_mux2_1 _17566_ (.A0(net3814),
    .A1(net3813),
    .S(\spiking_network_top_uut.all_data_out[556] ),
    .X(_02900_));
 sg13g2_nand2_1 _17567_ (.Y(_02901_),
    .A(\spiking_network_top_uut.all_data_out[557] ),
    .B(_02900_));
 sg13g2_a21oi_1 _17568_ (.A1(\spiking_network_top_uut.all_data_out[556] ),
    .A2(_03659_),
    .Y(_02902_),
    .B1(\spiking_network_top_uut.all_data_out[557] ));
 sg13g2_o21ai_1 _17569_ (.B1(_02902_),
    .Y(_02903_),
    .A1(\spiking_network_top_uut.all_data_out[556] ),
    .A2(net3815));
 sg13g2_nand3_1 _17570_ (.B(_02901_),
    .C(_02903_),
    .A(\spiking_network_top_uut.all_data_out[558] ),
    .Y(_02904_));
 sg13g2_nand3_1 _17571_ (.B(_02899_),
    .C(_02904_),
    .A(net4627),
    .Y(_02905_));
 sg13g2_o21ai_1 _17572_ (.B1(_02905_),
    .Y(_01043_),
    .A1(net4628),
    .A2(_03692_));
 sg13g2_mux2_1 _17573_ (.A0(net3812),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.din ),
    .S(net4624),
    .X(_01044_));
 sg13g2_mux2_1 _17574_ (.A0(net3811),
    .A1(net3812),
    .S(net4621),
    .X(_01045_));
 sg13g2_mux2_1 _17575_ (.A0(net3810),
    .A1(net3811),
    .S(net4621),
    .X(_01046_));
 sg13g2_mux2_1 _17576_ (.A0(net3809),
    .A1(net3810),
    .S(net4621),
    .X(_01047_));
 sg13g2_mux2_1 _17577_ (.A0(net3808),
    .A1(net3809),
    .S(net4621),
    .X(_01048_));
 sg13g2_mux2_1 _17578_ (.A0(net3807),
    .A1(net3808),
    .S(net4622),
    .X(_01049_));
 sg13g2_mux2_1 _17579_ (.A0(net3806),
    .A1(net3807),
    .S(net4622),
    .X(_01050_));
 sg13g2_mux2_1 _17580_ (.A0(net3805),
    .A1(net3806),
    .S(net4622),
    .X(_01051_));
 sg13g2_mux2_1 _17581_ (.A0(net301),
    .A1(net106),
    .S(net4628),
    .X(_01052_));
 sg13g2_mux2_1 _17582_ (.A0(net3810),
    .A1(net3809),
    .S(\spiking_network_top_uut.all_data_out[552] ),
    .X(_02906_));
 sg13g2_nor2b_1 _17583_ (.A(\spiking_network_top_uut.all_data_out[552] ),
    .B_N(net3812),
    .Y(_02907_));
 sg13g2_a21oi_1 _17584_ (.A1(\spiking_network_top_uut.all_data_out[552] ),
    .A2(net3811),
    .Y(_02908_),
    .B1(_02907_));
 sg13g2_a21oi_1 _17585_ (.A1(\spiking_network_top_uut.all_data_out[553] ),
    .A2(_02906_),
    .Y(_02909_),
    .B1(\spiking_network_top_uut.all_data_out[554] ));
 sg13g2_o21ai_1 _17586_ (.B1(_02909_),
    .Y(_02910_),
    .A1(\spiking_network_top_uut.all_data_out[553] ),
    .A2(_02908_));
 sg13g2_mux2_1 _17587_ (.A0(net3806),
    .A1(net3805),
    .S(\spiking_network_top_uut.all_data_out[552] ),
    .X(_02911_));
 sg13g2_nor2b_1 _17588_ (.A(\spiking_network_top_uut.all_data_out[552] ),
    .B_N(net3808),
    .Y(_02912_));
 sg13g2_a21oi_1 _17589_ (.A1(\spiking_network_top_uut.all_data_out[552] ),
    .A2(net3807),
    .Y(_02913_),
    .B1(_02912_));
 sg13g2_o21ai_1 _17590_ (.B1(\spiking_network_top_uut.all_data_out[554] ),
    .Y(_02914_),
    .A1(\spiking_network_top_uut.all_data_out[553] ),
    .A2(_02913_));
 sg13g2_a21oi_1 _17591_ (.A1(\spiking_network_top_uut.all_data_out[553] ),
    .A2(_02911_),
    .Y(_02915_),
    .B1(_02914_));
 sg13g2_nand2_1 _17592_ (.Y(_02916_),
    .A(net4624),
    .B(_02910_));
 sg13g2_nand2_1 _17593_ (.Y(_02917_),
    .A(net3959),
    .B(net67));
 sg13g2_o21ai_1 _17594_ (.B1(_02917_),
    .Y(_01053_),
    .A1(_02915_),
    .A2(_02916_));
 sg13g2_mux2_1 _17595_ (.A0(net3804),
    .A1(net4491),
    .S(net4632),
    .X(_01054_));
 sg13g2_mux2_1 _17596_ (.A0(net3803),
    .A1(net3804),
    .S(net4631),
    .X(_01055_));
 sg13g2_mux2_1 _17597_ (.A0(net3802),
    .A1(net3803),
    .S(net4631),
    .X(_01056_));
 sg13g2_mux2_1 _17598_ (.A0(net3801),
    .A1(net3802),
    .S(net4631),
    .X(_01057_));
 sg13g2_mux2_1 _17599_ (.A0(net3800),
    .A1(net3801),
    .S(net4631),
    .X(_01058_));
 sg13g2_mux2_1 _17600_ (.A0(net3799),
    .A1(net3800),
    .S(net4632),
    .X(_01059_));
 sg13g2_mux2_1 _17601_ (.A0(net3798),
    .A1(net3799),
    .S(net4633),
    .X(_01060_));
 sg13g2_mux2_1 _17602_ (.A0(net3797),
    .A1(net3798),
    .S(net4633),
    .X(_01061_));
 sg13g2_mux2_1 _17603_ (.A0(net322),
    .A1(net67),
    .S(net4624),
    .X(_01062_));
 sg13g2_mux4_1 _17604_ (.S0(\spiking_network_top_uut.all_data_out[548] ),
    .A0(net3804),
    .A1(net3803),
    .A2(net3802),
    .A3(net3801),
    .S1(\spiking_network_top_uut.all_data_out[549] ),
    .X(_02918_));
 sg13g2_mux2_1 _17605_ (.A0(net3798),
    .A1(net3797),
    .S(\spiking_network_top_uut.all_data_out[548] ),
    .X(_02919_));
 sg13g2_nor2b_1 _17606_ (.A(\spiking_network_top_uut.all_data_out[548] ),
    .B_N(net3800),
    .Y(_02920_));
 sg13g2_a21oi_1 _17607_ (.A1(\spiking_network_top_uut.all_data_out[548] ),
    .A2(net3799),
    .Y(_02921_),
    .B1(_02920_));
 sg13g2_o21ai_1 _17608_ (.B1(\spiking_network_top_uut.all_data_out[550] ),
    .Y(_02922_),
    .A1(\spiking_network_top_uut.all_data_out[549] ),
    .A2(_02921_));
 sg13g2_a21oi_1 _17609_ (.A1(\spiking_network_top_uut.all_data_out[549] ),
    .A2(_02919_),
    .Y(_02923_),
    .B1(_02922_));
 sg13g2_o21ai_1 _17610_ (.B1(net4631),
    .Y(_02924_),
    .A1(\spiking_network_top_uut.all_data_out[550] ),
    .A2(_02918_));
 sg13g2_nand2_1 _17611_ (.Y(_02925_),
    .A(net3961),
    .B(net119));
 sg13g2_o21ai_1 _17612_ (.B1(_02925_),
    .Y(_01063_),
    .A1(_02923_),
    .A2(_02924_));
 sg13g2_mux2_1 _17613_ (.A0(net3796),
    .A1(net4492),
    .S(net4620),
    .X(_01064_));
 sg13g2_mux2_1 _17614_ (.A0(net3795),
    .A1(net3796),
    .S(net4618),
    .X(_01065_));
 sg13g2_mux2_1 _17615_ (.A0(net3794),
    .A1(net3795),
    .S(net4634),
    .X(_01066_));
 sg13g2_mux2_1 _17616_ (.A0(net3793),
    .A1(net3794),
    .S(net4634),
    .X(_01067_));
 sg13g2_mux2_1 _17617_ (.A0(net3792),
    .A1(net3793),
    .S(net4634),
    .X(_01068_));
 sg13g2_nand2_1 _17618_ (.Y(_02926_),
    .A(net4617),
    .B(net3792));
 sg13g2_o21ai_1 _17619_ (.B1(_02926_),
    .Y(_01069_),
    .A1(net4617),
    .A2(_03658_));
 sg13g2_nor2_1 _17620_ (.A(net4617),
    .B(net3791),
    .Y(_02927_));
 sg13g2_a21oi_1 _17621_ (.A1(net4617),
    .A2(_03658_),
    .Y(_01070_),
    .B1(_02927_));
 sg13g2_mux2_1 _17622_ (.A0(net3790),
    .A1(net3791),
    .S(net4617),
    .X(_01071_));
 sg13g2_mux2_1 _17623_ (.A0(net233),
    .A1(net119),
    .S(net4631),
    .X(_01072_));
 sg13g2_a21oi_1 _17624_ (.A1(\spiking_network_top_uut.all_data_out[544] ),
    .A2(_03658_),
    .Y(_02928_),
    .B1(\spiking_network_top_uut.all_data_out[545] ));
 sg13g2_o21ai_1 _17625_ (.B1(_02928_),
    .Y(_02929_),
    .A1(\spiking_network_top_uut.all_data_out[544] ),
    .A2(net3792));
 sg13g2_mux2_1 _17626_ (.A0(net3791),
    .A1(net3790),
    .S(\spiking_network_top_uut.all_data_out[544] ),
    .X(_02930_));
 sg13g2_nand2_1 _17627_ (.Y(_02931_),
    .A(\spiking_network_top_uut.all_data_out[545] ),
    .B(_02930_));
 sg13g2_nand3_1 _17628_ (.B(_02929_),
    .C(_02931_),
    .A(\spiking_network_top_uut.all_data_out[546] ),
    .Y(_02932_));
 sg13g2_mux2_1 _17629_ (.A0(net3794),
    .A1(net3793),
    .S(\spiking_network_top_uut.all_data_out[544] ),
    .X(_02933_));
 sg13g2_nor2b_1 _17630_ (.A(\spiking_network_top_uut.all_data_out[544] ),
    .B_N(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[0] ),
    .Y(_02934_));
 sg13g2_a21oi_1 _17631_ (.A1(\spiking_network_top_uut.all_data_out[544] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[1] ),
    .Y(_02935_),
    .B1(_02934_));
 sg13g2_a21oi_1 _17632_ (.A1(\spiking_network_top_uut.all_data_out[545] ),
    .A2(_02933_),
    .Y(_02936_),
    .B1(\spiking_network_top_uut.all_data_out[546] ));
 sg13g2_o21ai_1 _17633_ (.B1(_02936_),
    .Y(_02937_),
    .A1(\spiking_network_top_uut.all_data_out[545] ),
    .A2(_02935_));
 sg13g2_nand3_1 _17634_ (.B(_02932_),
    .C(_02937_),
    .A(net4634),
    .Y(_02938_));
 sg13g2_o21ai_1 _17635_ (.B1(_02938_),
    .Y(_01073_),
    .A1(net4636),
    .A2(_03693_));
 sg13g2_nor3_2 _17636_ (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[2] ),
    .B(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[1] ),
    .C(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[0] ),
    .Y(_02939_));
 sg13g2_nor2b_2 _17637_ (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[3] ),
    .B_N(_02939_),
    .Y(_02940_));
 sg13g2_nor2b_2 _17638_ (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[4] ),
    .B_N(_02940_),
    .Y(_02941_));
 sg13g2_nand2b_2 _17639_ (.Y(_02942_),
    .B(_02940_),
    .A_N(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[4] ));
 sg13g2_o21ai_1 _17640_ (.B1(net4603),
    .Y(_02943_),
    .A1(net3636),
    .A2(net3699));
 sg13g2_nor2b_1 _17641_ (.A(net3635),
    .B_N(net390),
    .Y(_02944_));
 sg13g2_a21oi_1 _17642_ (.A1(net4284),
    .A2(net3635),
    .Y(_02945_),
    .B1(_02944_));
 sg13g2_nand2_1 _17643_ (.Y(_02946_),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[0] ),
    .B(_02943_));
 sg13g2_o21ai_1 _17644_ (.B1(_02946_),
    .Y(_01074_),
    .A1(_02943_),
    .A2(_02945_));
 sg13g2_xor2_1 _17645_ (.B(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[0] ),
    .A(net407),
    .X(_02947_));
 sg13g2_nor2_1 _17646_ (.A(net3635),
    .B(_02947_),
    .Y(_02948_));
 sg13g2_a21oi_1 _17647_ (.A1(net4281),
    .A2(net3635),
    .Y(_02949_),
    .B1(_02948_));
 sg13g2_nand2_1 _17648_ (.Y(_02950_),
    .A(net407),
    .B(_02943_));
 sg13g2_o21ai_1 _17649_ (.B1(_02950_),
    .Y(_01075_),
    .A1(_02943_),
    .A2(_02949_));
 sg13g2_o21ai_1 _17650_ (.B1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[2] ),
    .Y(_02951_),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[1] ),
    .A2(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[0] ));
 sg13g2_nor2b_1 _17651_ (.A(_02939_),
    .B_N(_02951_),
    .Y(_02952_));
 sg13g2_nor2_1 _17652_ (.A(net3635),
    .B(_02952_),
    .Y(_02953_));
 sg13g2_a21oi_1 _17653_ (.A1(net4277),
    .A2(net3635),
    .Y(_02954_),
    .B1(_02953_));
 sg13g2_nand2_1 _17654_ (.Y(_02955_),
    .A(net201),
    .B(_02943_));
 sg13g2_o21ai_1 _17655_ (.B1(_02955_),
    .Y(_01076_),
    .A1(_02943_),
    .A2(_02954_));
 sg13g2_nand2_1 _17656_ (.Y(_02956_),
    .A(net4274),
    .B(net3635));
 sg13g2_xnor2_1 _17657_ (.Y(_02957_),
    .A(net433),
    .B(_02939_));
 sg13g2_o21ai_1 _17658_ (.B1(_02956_),
    .Y(_02958_),
    .A1(net3635),
    .A2(_02957_));
 sg13g2_mux2_1 _17659_ (.A0(_02958_),
    .A1(net433),
    .S(_02943_),
    .X(_01077_));
 sg13g2_nand2_1 _17660_ (.Y(_02959_),
    .A(net3947),
    .B(net250));
 sg13g2_nor2_2 _17661_ (.A(net4271),
    .B(_04967_),
    .Y(_02960_));
 sg13g2_nor2b_1 _17662_ (.A(_02940_),
    .B_N(net250),
    .Y(_02961_));
 sg13g2_o21ai_1 _17663_ (.B1(net4603),
    .Y(_02962_),
    .A1(net3636),
    .A2(_02961_));
 sg13g2_o21ai_1 _17664_ (.B1(_02959_),
    .Y(_01078_),
    .A1(_02960_),
    .A2(_02962_));
 sg13g2_nor2_1 _17665_ (.A(net4636),
    .B(net184),
    .Y(_02963_));
 sg13g2_a21oi_1 _17666_ (.A1(net4636),
    .A2(_03693_),
    .Y(_01079_),
    .B1(_02963_));
 sg13g2_mux2_1 _17667_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[0] ),
    .A1(net4485),
    .S(net4644),
    .X(_01080_));
 sg13g2_mux2_1 _17668_ (.A0(net3788),
    .A1(net3789),
    .S(net4637),
    .X(_01081_));
 sg13g2_mux2_1 _17669_ (.A0(net3787),
    .A1(net3788),
    .S(net4628),
    .X(_01082_));
 sg13g2_mux2_1 _17670_ (.A0(net3786),
    .A1(net3787),
    .S(net4628),
    .X(_01083_));
 sg13g2_mux2_1 _17671_ (.A0(net3785),
    .A1(net3786),
    .S(net4628),
    .X(_01084_));
 sg13g2_mux2_1 _17672_ (.A0(net3784),
    .A1(net3785),
    .S(net4628),
    .X(_01085_));
 sg13g2_mux2_1 _17673_ (.A0(net3783),
    .A1(net3784),
    .S(net4637),
    .X(_01086_));
 sg13g2_a21oi_1 _17674_ (.A1(net3915),
    .A2(net3911),
    .Y(_02964_),
    .B1(_00133_));
 sg13g2_nor2_2 _17675_ (.A(net3751),
    .B(_02964_),
    .Y(_02965_));
 sg13g2_nor2_1 _17676_ (.A(_00133_),
    .B(_02965_),
    .Y(_02966_));
 sg13g2_nand2b_1 _17677_ (.Y(_02967_),
    .B(_02965_),
    .A_N(_00133_));
 sg13g2_o21ai_1 _17678_ (.B1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ),
    .Y(_02968_),
    .A1(_00133_),
    .A2(_02965_));
 sg13g2_inv_1 _17679_ (.Y(_02969_),
    .A(_02968_));
 sg13g2_a21o_1 _17680_ (.A2(net3751),
    .A1(_00134_),
    .B1(_02965_),
    .X(_02970_));
 sg13g2_nor2_1 _17681_ (.A(_00134_),
    .B(net3907),
    .Y(_02971_));
 sg13g2_a221oi_1 _17682_ (.B2(_02964_),
    .C1(_02971_),
    .B1(net3907),
    .A1(_03506_),
    .Y(_02972_),
    .A2(net3751));
 sg13g2_nand2_1 _17683_ (.Y(_02973_),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ),
    .B(_02972_));
 sg13g2_or2_1 _17684_ (.X(_02974_),
    .B(net3911),
    .A(_00133_));
 sg13g2_a21oi_1 _17685_ (.A1(net4266),
    .A2(_00134_),
    .Y(_02975_),
    .B1(_05084_));
 sg13g2_a21oi_1 _17686_ (.A1(_03506_),
    .A2(net3739),
    .Y(_02976_),
    .B1(_02975_));
 sg13g2_and2_1 _17687_ (.A(_00137_),
    .B(net3751),
    .X(_02977_));
 sg13g2_a21o_1 _17688_ (.A2(_02976_),
    .A1(_02974_),
    .B1(_02977_),
    .X(_02978_));
 sg13g2_a221oi_1 _17689_ (.B2(_02976_),
    .C1(_03507_),
    .B1(_02974_),
    .A1(_00137_),
    .Y(_02979_),
    .A2(net3751));
 sg13g2_xnor2_1 _17690_ (.Y(_02980_),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ),
    .B(_02972_));
 sg13g2_o21ai_1 _17691_ (.B1(_02973_),
    .Y(_02981_),
    .A1(_02979_),
    .A2(_02980_));
 sg13g2_xnor2_1 _17692_ (.Y(_02982_),
    .A(_03506_),
    .B(_02970_));
 sg13g2_nor2b_1 _17693_ (.A(_02982_),
    .B_N(_02981_),
    .Y(_02983_));
 sg13g2_a21o_1 _17694_ (.A2(_02970_),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ),
    .B1(_02983_),
    .X(_02984_));
 sg13g2_xnor2_1 _17695_ (.Y(_02985_),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ),
    .B(_02966_));
 sg13g2_a21oi_1 _17696_ (.A1(_02984_),
    .A2(_02985_),
    .Y(_02986_),
    .B1(_02969_));
 sg13g2_a22oi_1 _17697_ (.Y(_02987_),
    .B1(_02967_),
    .B2(_02986_),
    .A2(_02965_),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ));
 sg13g2_a21oi_2 _17698_ (.B1(_02987_),
    .Y(_02988_),
    .A2(_00133_),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ));
 sg13g2_mux2_2 _17699_ (.A0(net4491),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[551] ),
    .X(_02989_));
 sg13g2_nand2_1 _17700_ (.Y(_02990_),
    .A(\spiking_network_top_uut.all_data_out[147] ),
    .B(_02989_));
 sg13g2_mux2_2 _17701_ (.A0(net4492),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[547] ),
    .X(_02991_));
 sg13g2_nand2_1 _17702_ (.Y(_02992_),
    .A(\spiking_network_top_uut.all_data_out[145] ),
    .B(_02991_));
 sg13g2_nor2_1 _17703_ (.A(_02990_),
    .B(_02992_),
    .Y(_02993_));
 sg13g2_nand4_1 _17704_ (.B(\spiking_network_top_uut.all_data_out[144] ),
    .C(_02989_),
    .A(\spiking_network_top_uut.all_data_out[146] ),
    .Y(_02994_),
    .D(_02991_));
 sg13g2_inv_1 _17705_ (.Y(_02995_),
    .A(_02994_));
 sg13g2_xor2_1 _17706_ (.B(_02992_),
    .A(_02990_),
    .X(_02996_));
 sg13g2_a21oi_2 _17707_ (.B1(_02993_),
    .Y(_02997_),
    .A2(_02996_),
    .A1(_02994_));
 sg13g2_mux2_2 _17708_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.din ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[555] ),
    .X(_02998_));
 sg13g2_nand2_2 _17709_ (.Y(_02999_),
    .A(\spiking_network_top_uut.all_data_out[149] ),
    .B(_02998_));
 sg13g2_mux2_2 _17710_ (.A0(net4489),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[559] ),
    .X(_03000_));
 sg13g2_nand2_2 _17711_ (.Y(_03001_),
    .A(\spiking_network_top_uut.all_data_out[151] ),
    .B(_03000_));
 sg13g2_nor2_1 _17712_ (.A(_02999_),
    .B(_03001_),
    .Y(_03002_));
 sg13g2_nand2_2 _17713_ (.Y(_03003_),
    .A(\spiking_network_top_uut.all_data_out[148] ),
    .B(_02998_));
 sg13g2_nand2_2 _17714_ (.Y(_03004_),
    .A(\spiking_network_top_uut.all_data_out[150] ),
    .B(_03000_));
 sg13g2_or2_2 _17715_ (.X(_03005_),
    .B(_03004_),
    .A(_03003_));
 sg13g2_xor2_1 _17716_ (.B(_03001_),
    .A(_02999_),
    .X(_03006_));
 sg13g2_a21oi_2 _17717_ (.B1(_03002_),
    .Y(_03007_),
    .A2(_03006_),
    .A1(_03005_));
 sg13g2_mux2_2 _17718_ (.A0(net4487),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[567] ),
    .X(_03008_));
 sg13g2_mux2_2 _17719_ (.A0(net4488),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[563] ),
    .X(_03009_));
 sg13g2_a22oi_1 _17720_ (.Y(_03010_),
    .B1(_03009_),
    .B2(\spiking_network_top_uut.all_data_out[153] ),
    .A2(_03008_),
    .A1(\spiking_network_top_uut.all_data_out[155] ));
 sg13g2_and4_1 _17721_ (.A(\spiking_network_top_uut.all_data_out[155] ),
    .B(\spiking_network_top_uut.all_data_out[153] ),
    .C(_03008_),
    .D(_03009_),
    .X(_03011_));
 sg13g2_nand4_1 _17722_ (.B(\spiking_network_top_uut.all_data_out[153] ),
    .C(_03008_),
    .A(\spiking_network_top_uut.all_data_out[155] ),
    .Y(_03012_),
    .D(_03009_));
 sg13g2_and4_2 _17723_ (.A(\spiking_network_top_uut.all_data_out[154] ),
    .B(\spiking_network_top_uut.all_data_out[152] ),
    .C(_03008_),
    .D(_03009_),
    .X(_03013_));
 sg13g2_nand4_1 _17724_ (.B(\spiking_network_top_uut.all_data_out[152] ),
    .C(_03008_),
    .A(\spiking_network_top_uut.all_data_out[154] ),
    .Y(_03014_),
    .D(_03009_));
 sg13g2_nand3b_1 _17725_ (.B(_03012_),
    .C(_03013_),
    .Y(_03015_),
    .A_N(_03010_));
 sg13g2_a21oi_2 _17726_ (.B1(_03010_),
    .Y(_03016_),
    .A2(_03013_),
    .A1(_03012_));
 sg13g2_mux2_2 _17727_ (.A0(net4485),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[575] ),
    .X(_03017_));
 sg13g2_mux2_2 _17728_ (.A0(net4486),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_dout ),
    .S(\spiking_network_top_uut.all_data_out[571] ),
    .X(_03018_));
 sg13g2_and4_1 _17729_ (.A(\spiking_network_top_uut.all_data_out[159] ),
    .B(\spiking_network_top_uut.all_data_out[157] ),
    .C(_03017_),
    .D(_03018_),
    .X(_03019_));
 sg13g2_nand4_1 _17730_ (.B(\spiking_network_top_uut.all_data_out[157] ),
    .C(_03017_),
    .A(\spiking_network_top_uut.all_data_out[159] ),
    .Y(_03020_),
    .D(_03018_));
 sg13g2_and4_1 _17731_ (.A(\spiking_network_top_uut.all_data_out[158] ),
    .B(\spiking_network_top_uut.all_data_out[156] ),
    .C(_03017_),
    .D(_03018_),
    .X(_03021_));
 sg13g2_a22oi_1 _17732_ (.Y(_03022_),
    .B1(_03018_),
    .B2(\spiking_network_top_uut.all_data_out[157] ),
    .A2(_03017_),
    .A1(\spiking_network_top_uut.all_data_out[159] ));
 sg13g2_or3_2 _17733_ (.A(_03019_),
    .B(_03021_),
    .C(_03022_),
    .X(_03023_));
 sg13g2_o21ai_1 _17734_ (.B1(_03020_),
    .Y(_03024_),
    .A1(_03021_),
    .A2(_03022_));
 sg13g2_nand3b_1 _17735_ (.B(_03016_),
    .C(_03024_),
    .Y(_03025_),
    .A_N(_03007_));
 sg13g2_inv_1 _17736_ (.Y(_03026_),
    .A(_03025_));
 sg13g2_nor2_2 _17737_ (.A(_02997_),
    .B(_03025_),
    .Y(_03027_));
 sg13g2_nor2_1 _17738_ (.A(_03016_),
    .B(_03024_),
    .Y(_03028_));
 sg13g2_and2_1 _17739_ (.A(_03007_),
    .B(_03028_),
    .X(_03029_));
 sg13g2_a21oi_2 _17740_ (.B1(_03027_),
    .Y(_03030_),
    .A2(_03029_),
    .A1(_02997_));
 sg13g2_xor2_1 _17741_ (.B(_02986_),
    .A(_02967_),
    .X(_03031_));
 sg13g2_inv_1 _17742_ (.Y(_03032_),
    .A(_03031_));
 sg13g2_xnor2_1 _17743_ (.Y(_03033_),
    .A(_03030_),
    .B(_03031_));
 sg13g2_o21ai_1 _17744_ (.B1(_03021_),
    .Y(_03034_),
    .A1(_03019_),
    .A2(_03022_));
 sg13g2_o21ai_1 _17745_ (.B1(_03014_),
    .Y(_03035_),
    .A1(_03010_),
    .A2(_03011_));
 sg13g2_o21ai_1 _17746_ (.B1(_03013_),
    .Y(_03036_),
    .A1(_03010_),
    .A2(_03011_));
 sg13g2_nand3b_1 _17747_ (.B(_03012_),
    .C(_03014_),
    .Y(_03037_),
    .A_N(_03010_));
 sg13g2_a22oi_1 _17748_ (.Y(_03038_),
    .B1(_03036_),
    .B2(_03037_),
    .A2(_03034_),
    .A1(_03023_));
 sg13g2_xor2_1 _17749_ (.B(_03006_),
    .A(_03005_),
    .X(_03039_));
 sg13g2_xnor2_1 _17750_ (.Y(_03040_),
    .A(_03005_),
    .B(_03006_));
 sg13g2_and4_1 _17751_ (.A(_03023_),
    .B(_03034_),
    .C(_03036_),
    .D(_03037_),
    .X(_03041_));
 sg13g2_nand4_1 _17752_ (.B(_03034_),
    .C(_03036_),
    .A(_03023_),
    .Y(_03042_),
    .D(_03037_));
 sg13g2_and4_1 _17753_ (.A(_03015_),
    .B(_03023_),
    .C(_03034_),
    .D(_03035_),
    .X(_03043_));
 sg13g2_a22oi_1 _17754_ (.Y(_03044_),
    .B1(_03035_),
    .B2(_03015_),
    .A2(_03034_),
    .A1(_03023_));
 sg13g2_nor3_2 _17755_ (.A(_03038_),
    .B(_03039_),
    .C(_03041_),
    .Y(_03045_));
 sg13g2_a21oi_2 _17756_ (.B1(_03038_),
    .Y(_03046_),
    .A2(_03042_),
    .A1(_03040_));
 sg13g2_xor2_1 _17757_ (.B(_03024_),
    .A(_03016_),
    .X(_03047_));
 sg13g2_xnor2_1 _17758_ (.Y(_03048_),
    .A(_03007_),
    .B(_03047_));
 sg13g2_nor2b_1 _17759_ (.A(_03046_),
    .B_N(_03048_),
    .Y(_03049_));
 sg13g2_xnor2_1 _17760_ (.Y(_03050_),
    .A(_03046_),
    .B(_03048_));
 sg13g2_nor2b_1 _17761_ (.A(_02997_),
    .B_N(_03050_),
    .Y(_03051_));
 sg13g2_nor2_1 _17762_ (.A(_03049_),
    .B(_03051_),
    .Y(_03052_));
 sg13g2_nor2_1 _17763_ (.A(_03026_),
    .B(_03029_),
    .Y(_03053_));
 sg13g2_xnor2_1 _17764_ (.Y(_03054_),
    .A(_02997_),
    .B(_03053_));
 sg13g2_nor2b_1 _17765_ (.A(_03052_),
    .B_N(_03054_),
    .Y(_03055_));
 sg13g2_xnor2_1 _17766_ (.Y(_03056_),
    .A(_03052_),
    .B(_03054_));
 sg13g2_xnor2_1 _17767_ (.Y(_03057_),
    .A(_02984_),
    .B(_02985_));
 sg13g2_inv_1 _17768_ (.Y(_03058_),
    .A(_03057_));
 sg13g2_a21oi_1 _17769_ (.A1(_03056_),
    .A2(_03058_),
    .Y(_03059_),
    .B1(_03055_));
 sg13g2_nand2b_1 _17770_ (.Y(_03060_),
    .B(_03033_),
    .A_N(_03059_));
 sg13g2_xnor2_1 _17771_ (.Y(_03061_),
    .A(_03056_),
    .B(_03058_));
 sg13g2_a22oi_1 _17772_ (.Y(_03062_),
    .B1(_03018_),
    .B2(\spiking_network_top_uut.all_data_out[156] ),
    .A2(_03017_),
    .A1(\spiking_network_top_uut.all_data_out[158] ));
 sg13g2_nor2_2 _17773_ (.A(_03021_),
    .B(_03062_),
    .Y(_03063_));
 sg13g2_a22oi_1 _17774_ (.Y(_03064_),
    .B1(_03009_),
    .B2(\spiking_network_top_uut.all_data_out[152] ),
    .A2(_03008_),
    .A1(\spiking_network_top_uut.all_data_out[154] ));
 sg13g2_nor2_1 _17775_ (.A(_03013_),
    .B(_03064_),
    .Y(_03065_));
 sg13g2_and2_1 _17776_ (.A(_03063_),
    .B(_03065_),
    .X(_03066_));
 sg13g2_xor2_1 _17777_ (.B(_03004_),
    .A(_03003_),
    .X(_03067_));
 sg13g2_xor2_1 _17778_ (.B(_03065_),
    .A(_03063_),
    .X(_03068_));
 sg13g2_a21oi_2 _17779_ (.B1(_03066_),
    .Y(_03069_),
    .A2(_03068_),
    .A1(_03067_));
 sg13g2_nor3_2 _17780_ (.A(_03040_),
    .B(_03043_),
    .C(_03044_),
    .Y(_03070_));
 sg13g2_nor3_1 _17781_ (.A(_03045_),
    .B(_03069_),
    .C(_03070_),
    .Y(_03071_));
 sg13g2_or3_1 _17782_ (.A(_03045_),
    .B(_03069_),
    .C(_03070_),
    .X(_03072_));
 sg13g2_xnor2_1 _17783_ (.Y(_03073_),
    .A(_02994_),
    .B(_02996_));
 sg13g2_o21ai_1 _17784_ (.B1(_03069_),
    .Y(_03074_),
    .A1(_03045_),
    .A2(_03070_));
 sg13g2_nand3_1 _17785_ (.B(_03073_),
    .C(_03074_),
    .A(_03072_),
    .Y(_03075_));
 sg13g2_a21o_2 _17786_ (.A2(_03074_),
    .A1(_03073_),
    .B1(_03071_),
    .X(_03076_));
 sg13g2_xnor2_1 _17787_ (.Y(_03077_),
    .A(_02997_),
    .B(_03050_));
 sg13g2_nand2_1 _17788_ (.Y(_03078_),
    .A(_03076_),
    .B(_03077_));
 sg13g2_xnor2_1 _17789_ (.Y(_03079_),
    .A(_03076_),
    .B(_03077_));
 sg13g2_xor2_1 _17790_ (.B(_02982_),
    .A(_02981_),
    .X(_03080_));
 sg13g2_o21ai_1 _17791_ (.B1(_03078_),
    .Y(_03081_),
    .A1(_03079_),
    .A2(_03080_));
 sg13g2_nor2b_1 _17792_ (.A(_03061_),
    .B_N(_03081_),
    .Y(_03082_));
 sg13g2_a22oi_1 _17793_ (.Y(_03083_),
    .B1(_02991_),
    .B2(\spiking_network_top_uut.all_data_out[144] ),
    .A2(_02989_),
    .A1(\spiking_network_top_uut.all_data_out[146] ));
 sg13g2_nor2_1 _17794_ (.A(_02995_),
    .B(_03083_),
    .Y(_03084_));
 sg13g2_inv_1 _17795_ (.Y(_03085_),
    .A(_03084_));
 sg13g2_xnor2_1 _17796_ (.Y(_03086_),
    .A(_03067_),
    .B(_03068_));
 sg13g2_nor2_2 _17797_ (.A(_03085_),
    .B(_03086_),
    .Y(_03087_));
 sg13g2_a21o_2 _17798_ (.A2(_03074_),
    .A1(_03072_),
    .B1(_03073_),
    .X(_03088_));
 sg13g2_and3_1 _17799_ (.X(_03089_),
    .A(_03075_),
    .B(_03087_),
    .C(_03088_));
 sg13g2_nand3_1 _17800_ (.B(_03087_),
    .C(_03088_),
    .A(_03075_),
    .Y(_03090_));
 sg13g2_a21oi_1 _17801_ (.A1(_03075_),
    .A2(_03088_),
    .Y(_03091_),
    .B1(_03087_));
 sg13g2_xor2_1 _17802_ (.B(_02980_),
    .A(_02979_),
    .X(_03092_));
 sg13g2_inv_1 _17803_ (.Y(_03093_),
    .A(_03092_));
 sg13g2_nor3_1 _17804_ (.A(_03089_),
    .B(_03091_),
    .C(_03093_),
    .Y(_03094_));
 sg13g2_o21ai_1 _17805_ (.B1(_03090_),
    .Y(_03095_),
    .A1(_03091_),
    .A2(_03093_));
 sg13g2_xor2_1 _17806_ (.B(_03080_),
    .A(_03079_),
    .X(_03096_));
 sg13g2_nand2_1 _17807_ (.Y(_03097_),
    .A(_03095_),
    .B(_03096_));
 sg13g2_o21ai_1 _17808_ (.B1(_03093_),
    .Y(_03098_),
    .A1(_03089_),
    .A2(_03091_));
 sg13g2_nand2b_1 _17809_ (.Y(_03099_),
    .B(_03098_),
    .A_N(_03094_));
 sg13g2_xnor2_1 _17810_ (.Y(_03100_),
    .A(_03085_),
    .B(_03086_));
 sg13g2_xnor2_1 _17811_ (.Y(_03101_),
    .A(_00136_),
    .B(_02978_));
 sg13g2_nor2_1 _17812_ (.A(_03100_),
    .B(_03101_),
    .Y(_03102_));
 sg13g2_nand3b_1 _17813_ (.B(_03098_),
    .C(_03102_),
    .Y(_03103_),
    .A_N(_03094_));
 sg13g2_xnor2_1 _17814_ (.Y(_03104_),
    .A(_03095_),
    .B(_03096_));
 sg13g2_or2_1 _17815_ (.X(_03105_),
    .B(_03104_),
    .A(_03103_));
 sg13g2_o21ai_1 _17816_ (.B1(_03097_),
    .Y(_03106_),
    .A1(_03103_),
    .A2(_03104_));
 sg13g2_nand2b_1 _17817_ (.Y(_03107_),
    .B(_03061_),
    .A_N(_03081_));
 sg13g2_nand2b_1 _17818_ (.Y(_03108_),
    .B(_03107_),
    .A_N(_03082_));
 sg13g2_nor2b_1 _17819_ (.A(_03108_),
    .B_N(_03106_),
    .Y(_03109_));
 sg13g2_a21oi_1 _17820_ (.A1(_03106_),
    .A2(_03107_),
    .Y(_03110_),
    .B1(_03082_));
 sg13g2_xor2_1 _17821_ (.B(_03059_),
    .A(_03033_),
    .X(_03111_));
 sg13g2_nor2_1 _17822_ (.A(_03110_),
    .B(_03111_),
    .Y(_03112_));
 sg13g2_o21ai_1 _17823_ (.B1(_03060_),
    .Y(_03113_),
    .A1(_03110_),
    .A2(_03111_));
 sg13g2_a21oi_1 _17824_ (.A1(_03030_),
    .A2(_03032_),
    .Y(_03114_),
    .B1(_03027_));
 sg13g2_xor2_1 _17825_ (.B(_03030_),
    .A(_02988_),
    .X(_03115_));
 sg13g2_nand2b_1 _17826_ (.Y(_03116_),
    .B(_03115_),
    .A_N(_03114_));
 sg13g2_xnor2_1 _17827_ (.Y(_03117_),
    .A(_03114_),
    .B(_03115_));
 sg13g2_nand2_1 _17828_ (.Y(_03118_),
    .A(_03113_),
    .B(_03117_));
 sg13g2_xor2_1 _17829_ (.B(_03117_),
    .A(_03113_),
    .X(_03119_));
 sg13g2_or2_1 _17830_ (.X(_03120_),
    .B(_02988_),
    .A(_02941_));
 sg13g2_o21ai_1 _17831_ (.B1(_03120_),
    .Y(_03121_),
    .A1(_02942_),
    .A2(_03119_));
 sg13g2_nand2_1 _17832_ (.Y(_03122_),
    .A(_03110_),
    .B(_03111_));
 sg13g2_nor2_1 _17833_ (.A(net3699),
    .B(_03112_),
    .Y(_03123_));
 sg13g2_a22oi_1 _17834_ (.Y(_03124_),
    .B1(_03122_),
    .B2(_03123_),
    .A2(_03032_),
    .A1(net3699));
 sg13g2_or2_1 _17835_ (.X(_03125_),
    .B(_03124_),
    .A(_03121_));
 sg13g2_o21ai_1 _17836_ (.B1(_02988_),
    .Y(_03126_),
    .A1(net3699),
    .A2(_03027_));
 sg13g2_or3_1 _17837_ (.A(_02988_),
    .B(_03027_),
    .C(_03030_),
    .X(_03127_));
 sg13g2_nand3_1 _17838_ (.B(_03118_),
    .C(_03127_),
    .A(_03116_),
    .Y(_03128_));
 sg13g2_o21ai_1 _17839_ (.B1(_03126_),
    .Y(_03129_),
    .A1(net3699),
    .A2(_03128_));
 sg13g2_a21oi_1 _17840_ (.A1(_03125_),
    .A2(_03129_),
    .Y(_03130_),
    .B1(net3636));
 sg13g2_nand2_1 _17841_ (.Y(_03131_),
    .A(net4605),
    .B(_03130_));
 sg13g2_a21oi_2 _17842_ (.B1(_03129_),
    .Y(_03132_),
    .A2(_03124_),
    .A1(_03121_));
 sg13g2_nor2_1 _17843_ (.A(net3699),
    .B(_03100_),
    .Y(_03133_));
 sg13g2_xnor2_1 _17844_ (.Y(_03134_),
    .A(_03101_),
    .B(_03133_));
 sg13g2_nor2_1 _17845_ (.A(_03132_),
    .B(_03134_),
    .Y(_03135_));
 sg13g2_o21ai_1 _17846_ (.B1(net4605),
    .Y(_03136_),
    .A1(net4315),
    .A2(_04967_));
 sg13g2_a22oi_1 _17847_ (.Y(_03137_),
    .B1(_03136_),
    .B2(net447),
    .A2(_00008_),
    .A1(_04960_));
 sg13g2_o21ai_1 _17848_ (.B1(_03137_),
    .Y(_01087_),
    .A1(_03131_),
    .A2(_03135_));
 sg13g2_nor2_1 _17849_ (.A(_02941_),
    .B(_03092_),
    .Y(_03138_));
 sg13g2_xor2_1 _17850_ (.B(_03102_),
    .A(_03099_),
    .X(_03139_));
 sg13g2_a21oi_1 _17851_ (.A1(_02941_),
    .A2(_03139_),
    .Y(_03140_),
    .B1(_03138_));
 sg13g2_o21ai_1 _17852_ (.B1(_03130_),
    .Y(_03141_),
    .A1(_03132_),
    .A2(_03140_));
 sg13g2_xnor2_1 _17853_ (.Y(_03142_),
    .A(_04959_),
    .B(_04960_));
 sg13g2_a21oi_1 _17854_ (.A1(net3636),
    .A2(_03142_),
    .Y(_03143_),
    .B1(net3953));
 sg13g2_a22oi_1 _17855_ (.Y(_01088_),
    .B1(_03141_),
    .B2(_03143_),
    .A2(_03435_),
    .A1(net3952));
 sg13g2_nand2_1 _17856_ (.Y(_03144_),
    .A(_03103_),
    .B(_03104_));
 sg13g2_nand3_1 _17857_ (.B(_03105_),
    .C(_03144_),
    .A(_02941_),
    .Y(_03145_));
 sg13g2_o21ai_1 _17858_ (.B1(_03145_),
    .Y(_03146_),
    .A1(_02941_),
    .A2(_03080_));
 sg13g2_o21ai_1 _17859_ (.B1(_03130_),
    .Y(_03147_),
    .A1(_03132_),
    .A2(_03146_));
 sg13g2_xnor2_1 _17860_ (.Y(_03148_),
    .A(_04958_),
    .B(_04962_));
 sg13g2_a21oi_1 _17861_ (.A1(net3636),
    .A2(_03148_),
    .Y(_03149_),
    .B1(net3953));
 sg13g2_a22oi_1 _17862_ (.Y(_01089_),
    .B1(_03147_),
    .B2(_03149_),
    .A2(_03434_),
    .A1(net3953));
 sg13g2_nand2b_1 _17863_ (.Y(_03150_),
    .B(_03108_),
    .A_N(_03106_));
 sg13g2_nor2_1 _17864_ (.A(net3699),
    .B(_03109_),
    .Y(_03151_));
 sg13g2_a221oi_1 _17865_ (.B2(_03151_),
    .C1(_03132_),
    .B1(_03150_),
    .A1(net3699),
    .Y(_03152_),
    .A2(_03058_));
 sg13g2_or3_1 _17866_ (.A(_04956_),
    .B(_04957_),
    .C(_04963_),
    .X(_03153_));
 sg13g2_and2_1 _17867_ (.A(_04964_),
    .B(_03153_),
    .X(_03154_));
 sg13g2_a22oi_1 _17868_ (.Y(_03155_),
    .B1(_00008_),
    .B2(_03154_),
    .A2(net536),
    .A1(net3952));
 sg13g2_o21ai_1 _17869_ (.B1(_03155_),
    .Y(_01090_),
    .A1(_03131_),
    .A2(_03152_));
 sg13g2_o21ai_1 _17870_ (.B1(net4605),
    .Y(_03156_),
    .A1(_04954_),
    .A2(_04965_));
 sg13g2_a21oi_1 _17871_ (.A1(_04967_),
    .A2(_03129_),
    .Y(_03157_),
    .B1(_03156_));
 sg13g2_a21oi_1 _17872_ (.A1(net3952),
    .A2(_03433_),
    .Y(_01091_),
    .B1(_03157_));
 sg13g2_nand2b_1 _17873_ (.Y(_03158_),
    .B(\spiking_network_top_uut.clk_div_inst.counter[3] ),
    .A_N(\spiking_network_top_uut.all_data_out[27] ));
 sg13g2_a22oi_1 _17874_ (.Y(_03159_),
    .B1(\spiking_network_top_uut.all_data_out[24] ),
    .B2(_03398_),
    .A2(\spiking_network_top_uut.all_data_out[25] ),
    .A1(_03397_));
 sg13g2_nand2b_1 _17875_ (.Y(_03160_),
    .B(\spiking_network_top_uut.clk_div_inst.counter[2] ),
    .A_N(\spiking_network_top_uut.all_data_out[26] ));
 sg13g2_o21ai_1 _17876_ (.B1(_03160_),
    .Y(_03161_),
    .A1(_03397_),
    .A2(\spiking_network_top_uut.all_data_out[25] ));
 sg13g2_a22oi_1 _17877_ (.Y(_03162_),
    .B1(_03396_),
    .B2(\spiking_network_top_uut.all_data_out[26] ),
    .A2(\spiking_network_top_uut.all_data_out[27] ),
    .A1(_03395_));
 sg13g2_o21ai_1 _17878_ (.B1(_03162_),
    .Y(_03163_),
    .A1(_03159_),
    .A2(_03161_));
 sg13g2_a22oi_1 _17879_ (.Y(_03164_),
    .B1(_03158_),
    .B2(_03163_),
    .A2(\spiking_network_top_uut.all_data_out[28] ),
    .A1(_03393_));
 sg13g2_a22oi_1 _17880_ (.Y(_03165_),
    .B1(\spiking_network_top_uut.clk_div_inst.counter[4] ),
    .B2(_03394_),
    .A2(_03392_),
    .A1(\spiking_network_top_uut.clk_div_inst.counter[5] ));
 sg13g2_nand2b_1 _17881_ (.Y(_03166_),
    .B(_03165_),
    .A_N(_03164_));
 sg13g2_o21ai_1 _17882_ (.B1(_03166_),
    .Y(_03167_),
    .A1(\spiking_network_top_uut.clk_div_inst.counter[5] ),
    .A2(_03392_));
 sg13g2_o21ai_1 _17883_ (.B1(_03167_),
    .Y(_03168_),
    .A1(_03391_),
    .A2(\spiking_network_top_uut.all_data_out[30] ));
 sg13g2_a22oi_1 _17884_ (.Y(_03169_),
    .B1(_03391_),
    .B2(\spiking_network_top_uut.all_data_out[30] ),
    .A2(\spiking_network_top_uut.all_data_out[31] ),
    .A1(_03389_));
 sg13g2_a22oi_1 _17885_ (.Y(_03170_),
    .B1(_03168_),
    .B2(_03169_),
    .A2(_03390_),
    .A1(\spiking_network_top_uut.clk_div_inst.counter[7] ));
 sg13g2_nor2b_1 _17886_ (.A(_03170_),
    .B_N(\spiking_network_top_uut.clk_div_inst.enable ),
    .Y(_03171_));
 sg13g2_xnor2_1 _17887_ (.Y(_03172_),
    .A(net429),
    .B(\spiking_network_top_uut.clk_div_inst.enable ));
 sg13g2_nor2_1 _17888_ (.A(net3616),
    .B(net430),
    .Y(_01092_));
 sg13g2_and3_1 _17889_ (.X(_03173_),
    .A(net100),
    .B(\spiking_network_top_uut.clk_div_inst.counter[0] ),
    .C(\spiking_network_top_uut.clk_div_inst.enable ));
 sg13g2_a21oi_1 _17890_ (.A1(\spiking_network_top_uut.clk_div_inst.counter[0] ),
    .A2(\spiking_network_top_uut.clk_div_inst.enable ),
    .Y(_03174_),
    .B1(net100));
 sg13g2_nor3_1 _17891_ (.A(net3616),
    .B(_03173_),
    .C(net101),
    .Y(_01093_));
 sg13g2_and2_1 _17892_ (.A(net371),
    .B(_03173_),
    .X(_03175_));
 sg13g2_nor2_1 _17893_ (.A(net371),
    .B(_03173_),
    .Y(_03176_));
 sg13g2_nor3_1 _17894_ (.A(net3616),
    .B(_03175_),
    .C(net372),
    .Y(_01094_));
 sg13g2_and2_1 _17895_ (.A(net386),
    .B(_03175_),
    .X(_03177_));
 sg13g2_nor2_1 _17896_ (.A(net386),
    .B(_03175_),
    .Y(_03178_));
 sg13g2_nor3_1 _17897_ (.A(net3616),
    .B(_03177_),
    .C(_03178_),
    .Y(_01095_));
 sg13g2_xnor2_1 _17898_ (.Y(_03179_),
    .A(net448),
    .B(_03177_));
 sg13g2_nor2_1 _17899_ (.A(net3616),
    .B(_03179_),
    .Y(_01096_));
 sg13g2_nand3_1 _17900_ (.B(net448),
    .C(_03177_),
    .A(net468),
    .Y(_03180_));
 sg13g2_a21oi_1 _17901_ (.A1(net448),
    .A2(_03177_),
    .Y(_03181_),
    .B1(net468));
 sg13g2_nor2_1 _17902_ (.A(net3616),
    .B(_03181_),
    .Y(_03182_));
 sg13g2_and2_1 _17903_ (.A(_03180_),
    .B(_03182_),
    .X(_01097_));
 sg13g2_or2_1 _17904_ (.X(_03183_),
    .B(_03180_),
    .A(_03391_));
 sg13g2_xnor2_1 _17905_ (.Y(_03184_),
    .A(_03391_),
    .B(_03180_));
 sg13g2_nor2_1 _17906_ (.A(net3616),
    .B(_03184_),
    .Y(_01098_));
 sg13g2_xnor2_1 _17907_ (.Y(_03185_),
    .A(_03389_),
    .B(_03183_));
 sg13g2_nor2_1 _17908_ (.A(net3616),
    .B(_03185_),
    .Y(_01099_));
 sg13g2_mux2_1 _17909_ (.A0(net4505),
    .A1(net40),
    .S(_03171_),
    .X(_01100_));
 sg13g2_mux2_1 _17910_ (.A0(net4492),
    .A1(net2),
    .S(\spiking_network_top_uut.input_ready_sync ),
    .X(_01101_));
 sg13g2_mux2_1 _17911_ (.A0(net4491),
    .A1(net3),
    .S(\spiking_network_top_uut.input_ready_sync ),
    .X(_01102_));
 sg13g2_mux2_1 _17912_ (.A0(net4490),
    .A1(net4),
    .S(\spiking_network_top_uut.input_ready_sync ),
    .X(_01103_));
 sg13g2_mux2_1 _17913_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.din ),
    .A1(net5),
    .S(\spiking_network_top_uut.input_ready_sync ),
    .X(_01104_));
 sg13g2_mux2_1 _17914_ (.A0(net399),
    .A1(net6),
    .S(\spiking_network_top_uut.input_ready_sync ),
    .X(_01105_));
 sg13g2_mux2_1 _17915_ (.A0(net281),
    .A1(net7),
    .S(\spiking_network_top_uut.input_ready_sync ),
    .X(_01106_));
 sg13g2_mux2_1 _17916_ (.A0(net4486),
    .A1(net8),
    .S(\spiking_network_top_uut.input_ready_sync ),
    .X(_01107_));
 sg13g2_mux2_1 _17917_ (.A0(net4485),
    .A1(net9),
    .S(\spiking_network_top_uut.input_ready_sync ),
    .X(_01108_));
 sg13g2_mux2_1 _17918_ (.A0(\spiking_network_top_uut.clk_div_ready_reg_out ),
    .A1(\spiking_network_top_uut.spi_inst.clk_div_ready_reg_in ),
    .S(\spiking_network_top_uut.spi_inst.clk_div_ready_reg_en ),
    .X(_01109_));
 sg13g2_mux2_1 _17919_ (.A0(\spiking_network_top_uut.spi_inst.LSB_Address_reg[0] ),
    .A1(net4473),
    .S(\spiking_network_top_uut.spi_inst.SPI_address_LSB_reg_en ),
    .X(_01110_));
 sg13g2_mux2_1 _17920_ (.A0(\spiking_network_top_uut.spi_inst.LSB_Address_reg[1] ),
    .A1(net4452),
    .S(\spiking_network_top_uut.spi_inst.SPI_address_LSB_reg_en ),
    .X(_01111_));
 sg13g2_nand2_1 _17921_ (.Y(_03186_),
    .A(net4432),
    .B(\spiking_network_top_uut.spi_inst.SPI_address_LSB_reg_en ));
 sg13g2_o21ai_1 _17922_ (.B1(_03186_),
    .Y(_01112_),
    .A1(_03405_),
    .A2(\spiking_network_top_uut.spi_inst.SPI_address_LSB_reg_en ));
 sg13g2_mux2_1 _17923_ (.A0(\spiking_network_top_uut.spi_inst.LSB_Address_reg[3] ),
    .A1(net4413),
    .S(\spiking_network_top_uut.spi_inst.SPI_address_LSB_reg_en ),
    .X(_01113_));
 sg13g2_mux2_1 _17924_ (.A0(\spiking_network_top_uut.spi_inst.LSB_Address_reg[4] ),
    .A1(net4392),
    .S(\spiking_network_top_uut.spi_inst.SPI_address_LSB_reg_en ),
    .X(_01114_));
 sg13g2_mux2_1 _17925_ (.A0(\spiking_network_top_uut.spi_inst.LSB_Address_reg[5] ),
    .A1(net4370),
    .S(\spiking_network_top_uut.spi_inst.SPI_address_LSB_reg_en ),
    .X(_01115_));
 sg13g2_mux2_1 _17926_ (.A0(\spiking_network_top_uut.spi_inst.LSB_Address_reg[6] ),
    .A1(net4347),
    .S(\spiking_network_top_uut.spi_inst.SPI_address_LSB_reg_en ),
    .X(_01116_));
 sg13g2_mux2_1 _17927_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[0] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.spike_out ),
    .S(net4585),
    .X(_01117_));
 sg13g2_mux2_1 _17928_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[1] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[0] ),
    .S(net4584),
    .X(_01118_));
 sg13g2_mux2_1 _17929_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[2] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[1] ),
    .S(net4584),
    .X(_01119_));
 sg13g2_mux2_1 _17930_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[3] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[2] ),
    .S(net4584),
    .X(_01120_));
 sg13g2_mux2_1 _17931_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[4] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[3] ),
    .S(net4584),
    .X(_01121_));
 sg13g2_mux2_1 _17932_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[5] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[4] ),
    .S(net4584),
    .X(_01122_));
 sg13g2_mux2_1 _17933_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[6] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[5] ),
    .S(net4584),
    .X(_01123_));
 sg13g2_mux2_1 _17934_ (.A0(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[7] ),
    .A1(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[6] ),
    .S(net4584),
    .X(_01124_));
 sg13g2_mux2_1 _17935_ (.A0(\spiking_network_top_uut.spi_inst.SPI_instruction_reg[0] ),
    .A1(net4464),
    .S(net4318),
    .X(_01125_));
 sg13g2_mux2_1 _17936_ (.A0(\spiking_network_top_uut.spi_inst.SPI_instruction_reg[1] ),
    .A1(net4443),
    .S(net4318),
    .X(_01126_));
 sg13g2_mux2_1 _17937_ (.A0(\spiking_network_top_uut.spi_inst.SPI_instruction_reg[2] ),
    .A1(net4424),
    .S(\spiking_network_top_uut.spi_inst.SPI_instruction_reg_en ),
    .X(_01127_));
 sg13g2_nand2_1 _17938_ (.Y(_03187_),
    .A(net4403),
    .B(net4318));
 sg13g2_o21ai_1 _17939_ (.B1(_03187_),
    .Y(_01128_),
    .A1(_03472_),
    .A2(net4318));
 sg13g2_mux2_1 _17940_ (.A0(\spiking_network_top_uut.spi_inst.SPI_instruction_reg[4] ),
    .A1(net4380),
    .S(net4318),
    .X(_01129_));
 sg13g2_mux2_1 _17941_ (.A0(\spiking_network_top_uut.spi_inst.SPI_instruction_reg[5] ),
    .A1(net4361),
    .S(net4318),
    .X(_01130_));
 sg13g2_mux2_1 _17942_ (.A0(\spiking_network_top_uut.spi_inst.SPI_instruction_reg[6] ),
    .A1(net4339),
    .S(net4318),
    .X(_01131_));
 sg13g2_mux2_1 _17943_ (.A0(\spiking_network_top_uut.spi_inst.SPI_instruction_reg[7] ),
    .A1(net4320),
    .S(net4318),
    .X(_01132_));
 sg13g2_o21ai_1 _17944_ (.B1(_00028_),
    .Y(_03188_),
    .A1(\spiking_network_top_uut.spi_inst.spi_control_unit_inst.current_state[1] ),
    .A2(\spiking_network_top_uut.spi_inst.spi_control_unit_inst.current_state[0] ));
 sg13g2_inv_1 _17945_ (.Y(_03189_),
    .A(_03188_));
 sg13g2_nor2_1 _17946_ (.A(\spiking_network_top_uut.data_valid_out ),
    .B(_03188_),
    .Y(_03190_));
 sg13g2_nor2_1 _17947_ (.A(_03470_),
    .B(_04968_),
    .Y(_03191_));
 sg13g2_a221oi_1 _17948_ (.B2(_03469_),
    .C1(_03190_),
    .B1(_03191_),
    .A1(_00029_),
    .Y(_03192_),
    .A2(_04971_));
 sg13g2_a21o_1 _17949_ (.A2(_03701_),
    .A1(_03698_),
    .B1(_04972_),
    .X(_03193_));
 sg13g2_nand3_1 _17950_ (.B(_03192_),
    .C(_03193_),
    .A(_04968_),
    .Y(_03194_));
 sg13g2_o21ai_1 _17951_ (.B1(_03194_),
    .Y(_03195_),
    .A1(\spiking_network_top_uut.spi_inst.spi_control_unit_inst.current_state[0] ),
    .A2(_03192_));
 sg13g2_inv_1 _17952_ (.Y(_01133_),
    .A(_03195_));
 sg13g2_nand3_1 _17953_ (.B(_03189_),
    .C(_03192_),
    .A(_04594_),
    .Y(_03196_));
 sg13g2_o21ai_1 _17954_ (.B1(_03196_),
    .Y(_01134_),
    .A1(_03469_),
    .A2(_03192_));
 sg13g2_nand3_1 _17955_ (.B(_03192_),
    .C(_03193_),
    .A(_04595_),
    .Y(_03197_));
 sg13g2_o21ai_1 _17956_ (.B1(_03197_),
    .Y(_03198_),
    .A1(\spiking_network_top_uut.spi_inst.spi_control_unit_inst.current_state[2] ),
    .A2(_03192_));
 sg13g2_inv_1 _17957_ (.Y(_01135_),
    .A(_03198_));
 sg13g2_mux2_1 _17958_ (.A0(net4470),
    .A1(net11),
    .S(net3722),
    .X(_01136_));
 sg13g2_mux2_1 _17959_ (.A0(net4447),
    .A1(\spiking_network_top_uut.spi_inst.spi_slave_inst.shift_reg[0] ),
    .S(net3722),
    .X(_01137_));
 sg13g2_mux2_1 _17960_ (.A0(net4429),
    .A1(\spiking_network_top_uut.spi_inst.spi_slave_inst.shift_reg[1] ),
    .S(net3720),
    .X(_01138_));
 sg13g2_mux2_1 _17961_ (.A0(net4408),
    .A1(\spiking_network_top_uut.spi_inst.spi_slave_inst.shift_reg[2] ),
    .S(net3720),
    .X(_01139_));
 sg13g2_mux2_1 _17962_ (.A0(net4385),
    .A1(\spiking_network_top_uut.spi_inst.spi_slave_inst.shift_reg[3] ),
    .S(net3721),
    .X(_01140_));
 sg13g2_mux2_1 _17963_ (.A0(net4367),
    .A1(\spiking_network_top_uut.spi_inst.spi_slave_inst.shift_reg[4] ),
    .S(net3720),
    .X(_01141_));
 sg13g2_mux2_1 _17964_ (.A0(net4343),
    .A1(\spiking_network_top_uut.spi_inst.spi_slave_inst.shift_reg[5] ),
    .S(net3720),
    .X(_01142_));
 sg13g2_mux2_1 _17965_ (.A0(net4323),
    .A1(\spiking_network_top_uut.spi_inst.spi_slave_inst.shift_reg[6] ),
    .S(net3720),
    .X(_01143_));
 sg13g2_nor3_2 _17966_ (.A(\spiking_network_top_uut.spi_inst.LSB_Address_reg[2] ),
    .B(\spiking_network_top_uut.spi_inst.LSB_Address_reg[3] ),
    .C(_03406_),
    .Y(_03199_));
 sg13g2_nor2_2 _17967_ (.A(net4484),
    .B(net4483),
    .Y(_03200_));
 sg13g2_nand2_2 _17968_ (.Y(_03201_),
    .A(net3737),
    .B(_03200_));
 sg13g2_nand2_1 _17969_ (.Y(_03202_),
    .A(\spiking_network_top_uut.spi_inst.LSB_Address_reg[4] ),
    .B(\spiking_network_top_uut.spi_inst.LSB_Address_reg[5] ));
 sg13g2_nor3_2 _17970_ (.A(_00027_),
    .B(_03201_),
    .C(_03202_),
    .Y(_03203_));
 sg13g2_mux2_1 _17971_ (.A0(\spiking_network_top_uut.all_data_out[896] ),
    .A1(net4462),
    .S(_03203_),
    .X(_01144_));
 sg13g2_mux2_1 _17972_ (.A0(\spiking_network_top_uut.all_data_out[897] ),
    .A1(net4442),
    .S(_03203_),
    .X(_01145_));
 sg13g2_mux2_1 _17973_ (.A0(\spiking_network_top_uut.all_data_out[898] ),
    .A1(net4423),
    .S(_03203_),
    .X(_01146_));
 sg13g2_mux2_1 _17974_ (.A0(\spiking_network_top_uut.all_data_out[899] ),
    .A1(net4401),
    .S(_03203_),
    .X(_01147_));
 sg13g2_mux2_1 _17975_ (.A0(\spiking_network_top_uut.all_data_out[900] ),
    .A1(net4381),
    .S(_03203_),
    .X(_01148_));
 sg13g2_mux2_1 _17976_ (.A0(\spiking_network_top_uut.all_data_out[901] ),
    .A1(net4360),
    .S(_03203_),
    .X(_01149_));
 sg13g2_mux2_1 _17977_ (.A0(\spiking_network_top_uut.all_data_out[902] ),
    .A1(net4340),
    .S(_03203_),
    .X(_01150_));
 sg13g2_mux2_1 _17978_ (.A0(\spiking_network_top_uut.all_data_out[903] ),
    .A1(net4319),
    .S(_03203_),
    .X(_01151_));
 sg13g2_and4_1 _17979_ (.A(\spiking_network_top_uut.data_valid_out ),
    .B(_03698_),
    .C(_03701_),
    .D(_04971_),
    .X(_03204_));
 sg13g2_a21oi_1 _17980_ (.A1(spi_instruction_done),
    .A2(_04972_),
    .Y(_03205_),
    .B1(_03204_));
 sg13g2_o21ai_1 _17981_ (.B1(_03695_),
    .Y(_01152_),
    .A1(_03189_),
    .A2(_03205_));
 sg13g2_or2_2 _17982_ (.X(_03206_),
    .B(_03202_),
    .A(\spiking_network_top_uut.spi_inst.LSB_Address_reg[6] ));
 sg13g2_nor3_2 _17983_ (.A(_03405_),
    .B(\spiking_network_top_uut.spi_inst.LSB_Address_reg[3] ),
    .C(_03406_),
    .Y(_03207_));
 sg13g2_nand3_1 _17984_ (.B(\spiking_network_top_uut.spi_inst.LSB_Address_reg[1] ),
    .C(_03207_),
    .A(\spiking_network_top_uut.spi_inst.LSB_Address_reg[0] ),
    .Y(_03208_));
 sg13g2_nor2_2 _17985_ (.A(net3735),
    .B(_03208_),
    .Y(_03209_));
 sg13g2_mux2_1 _17986_ (.A0(\spiking_network_top_uut.all_data_out[440] ),
    .A1(net4479),
    .S(_03209_),
    .X(_01153_));
 sg13g2_mux2_1 _17987_ (.A0(\spiking_network_top_uut.all_data_out[441] ),
    .A1(net4458),
    .S(_03209_),
    .X(_01154_));
 sg13g2_mux2_1 _17988_ (.A0(\spiking_network_top_uut.all_data_out[442] ),
    .A1(net4437),
    .S(_03209_),
    .X(_01155_));
 sg13g2_mux2_1 _17989_ (.A0(\spiking_network_top_uut.all_data_out[443] ),
    .A1(net4414),
    .S(_03209_),
    .X(_01156_));
 sg13g2_mux2_1 _17990_ (.A0(\spiking_network_top_uut.all_data_out[444] ),
    .A1(net4399),
    .S(_03209_),
    .X(_01157_));
 sg13g2_mux2_1 _17991_ (.A0(\spiking_network_top_uut.all_data_out[445] ),
    .A1(net4379),
    .S(_03209_),
    .X(_01158_));
 sg13g2_mux2_1 _17992_ (.A0(\spiking_network_top_uut.all_data_out[446] ),
    .A1(net4358),
    .S(_03209_),
    .X(_01159_));
 sg13g2_mux2_1 _17993_ (.A0(\spiking_network_top_uut.all_data_out[447] ),
    .A1(net4330),
    .S(_03209_),
    .X(_01160_));
 sg13g2_nor2_2 _17994_ (.A(\spiking_network_top_uut.spi_inst.LSB_Address_reg[4] ),
    .B(\spiking_network_top_uut.spi_inst.LSB_Address_reg[5] ),
    .Y(_03210_));
 sg13g2_nand2b_2 _17995_ (.Y(_03211_),
    .B(_03210_),
    .A_N(_00027_));
 sg13g2_nand2_2 _17996_ (.Y(_03212_),
    .A(\spiking_network_top_uut.spi_inst.LSB_Address_reg[3] ),
    .B(net4317));
 sg13g2_nor2_2 _17997_ (.A(_03405_),
    .B(_03212_),
    .Y(_03213_));
 sg13g2_nor2b_2 _17998_ (.A(net4483),
    .B_N(net4484),
    .Y(_03214_));
 sg13g2_nand2_2 _17999_ (.Y(_03215_),
    .A(_03213_),
    .B(_03214_));
 sg13g2_nor2_2 _18000_ (.A(net3733),
    .B(_03215_),
    .Y(_03216_));
 sg13g2_mux2_1 _18001_ (.A0(\spiking_network_top_uut.all_data_out[616] ),
    .A1(net4477),
    .S(_03216_),
    .X(_01161_));
 sg13g2_mux2_1 _18002_ (.A0(\spiking_network_top_uut.all_data_out[617] ),
    .A1(net4457),
    .S(_03216_),
    .X(_01162_));
 sg13g2_mux2_1 _18003_ (.A0(\spiking_network_top_uut.all_data_out[618] ),
    .A1(net4436),
    .S(_03216_),
    .X(_01163_));
 sg13g2_mux2_1 _18004_ (.A0(\spiking_network_top_uut.all_data_out[619] ),
    .A1(net4417),
    .S(_03216_),
    .X(_01164_));
 sg13g2_mux2_1 _18005_ (.A0(\spiking_network_top_uut.all_data_out[620] ),
    .A1(net4394),
    .S(_03216_),
    .X(_01165_));
 sg13g2_mux2_1 _18006_ (.A0(\spiking_network_top_uut.all_data_out[621] ),
    .A1(net4378),
    .S(_03216_),
    .X(_01166_));
 sg13g2_mux2_1 _18007_ (.A0(\spiking_network_top_uut.all_data_out[622] ),
    .A1(net4353),
    .S(_03216_),
    .X(_01167_));
 sg13g2_mux2_1 _18008_ (.A0(\spiking_network_top_uut.all_data_out[623] ),
    .A1(net4335),
    .S(_03216_),
    .X(_01168_));
 sg13g2_nor2b_2 _18009_ (.A(net4484),
    .B_N(net4483),
    .Y(_03217_));
 sg13g2_nand2_2 _18010_ (.Y(_03218_),
    .A(_03207_),
    .B(_03217_));
 sg13g2_nor2_1 _18011_ (.A(net3735),
    .B(_03218_),
    .Y(_03219_));
 sg13g2_mux2_1 _18012_ (.A0(\spiking_network_top_uut.all_data_out[432] ),
    .A1(net4475),
    .S(net3692),
    .X(_01169_));
 sg13g2_mux2_1 _18013_ (.A0(\spiking_network_top_uut.all_data_out[433] ),
    .A1(net4455),
    .S(net3692),
    .X(_01170_));
 sg13g2_mux2_1 _18014_ (.A0(\spiking_network_top_uut.all_data_out[434] ),
    .A1(net4433),
    .S(net3692),
    .X(_01171_));
 sg13g2_mux2_1 _18015_ (.A0(\spiking_network_top_uut.all_data_out[435] ),
    .A1(net4415),
    .S(_03219_),
    .X(_01172_));
 sg13g2_mux2_1 _18016_ (.A0(\spiking_network_top_uut.all_data_out[436] ),
    .A1(net4391),
    .S(net3692),
    .X(_01173_));
 sg13g2_mux2_1 _18017_ (.A0(\spiking_network_top_uut.all_data_out[437] ),
    .A1(net4370),
    .S(net3692),
    .X(_01174_));
 sg13g2_nand2_1 _18018_ (.Y(_03220_),
    .A(net4350),
    .B(net3692));
 sg13g2_o21ai_1 _18019_ (.B1(_03220_),
    .Y(_01175_),
    .A1(_03539_),
    .A2(net3692));
 sg13g2_mux2_1 _18020_ (.A0(\spiking_network_top_uut.all_data_out[439] ),
    .A1(net4329),
    .S(net3692),
    .X(_01176_));
 sg13g2_nor2b_1 _18021_ (.A(\spiking_network_top_uut.spi_inst.LSB_Address_reg[5] ),
    .B_N(\spiking_network_top_uut.spi_inst.LSB_Address_reg[4] ),
    .Y(_03221_));
 sg13g2_nand2b_1 _18022_ (.Y(_03222_),
    .B(\spiking_network_top_uut.spi_inst.LSB_Address_reg[4] ),
    .A_N(\spiking_network_top_uut.spi_inst.LSB_Address_reg[5] ));
 sg13g2_nor2_2 _18023_ (.A(_00027_),
    .B(_03222_),
    .Y(_03223_));
 sg13g2_nand2b_1 _18024_ (.Y(_03224_),
    .B(_03221_),
    .A_N(_00027_));
 sg13g2_nand2_2 _18025_ (.Y(_03225_),
    .A(_03207_),
    .B(_03214_));
 sg13g2_nor2_2 _18026_ (.A(net3732),
    .B(_03225_),
    .Y(_03226_));
 sg13g2_mux2_1 _18027_ (.A0(\spiking_network_top_uut.all_data_out[680] ),
    .A1(net4476),
    .S(_03226_),
    .X(_01177_));
 sg13g2_mux2_1 _18028_ (.A0(\spiking_network_top_uut.all_data_out[681] ),
    .A1(net4456),
    .S(net3691),
    .X(_01178_));
 sg13g2_nand2_1 _18029_ (.Y(_03227_),
    .A(net4435),
    .B(net3691));
 sg13g2_o21ai_1 _18030_ (.B1(_03227_),
    .Y(_01179_),
    .A1(_03596_),
    .A2(net3691));
 sg13g2_mux2_1 _18031_ (.A0(\spiking_network_top_uut.all_data_out[683] ),
    .A1(net4413),
    .S(net3691),
    .X(_01180_));
 sg13g2_mux2_1 _18032_ (.A0(\spiking_network_top_uut.all_data_out[684] ),
    .A1(net4395),
    .S(net3691),
    .X(_01181_));
 sg13g2_mux2_1 _18033_ (.A0(\spiking_network_top_uut.all_data_out[685] ),
    .A1(net4374),
    .S(net3691),
    .X(_01182_));
 sg13g2_mux2_1 _18034_ (.A0(\spiking_network_top_uut.all_data_out[686] ),
    .A1(net4354),
    .S(net3691),
    .X(_01183_));
 sg13g2_mux2_1 _18035_ (.A0(\spiking_network_top_uut.all_data_out[687] ),
    .A1(net4333),
    .S(net3691),
    .X(_01184_));
 sg13g2_nor2_2 _18036_ (.A(_03206_),
    .B(_03225_),
    .Y(_03228_));
 sg13g2_mux2_1 _18037_ (.A0(\spiking_network_top_uut.all_data_out[424] ),
    .A1(net4477),
    .S(_03228_),
    .X(_01185_));
 sg13g2_mux2_1 _18038_ (.A0(\spiking_network_top_uut.all_data_out[425] ),
    .A1(net4457),
    .S(net3690),
    .X(_01186_));
 sg13g2_mux2_1 _18039_ (.A0(\spiking_network_top_uut.all_data_out[426] ),
    .A1(net4436),
    .S(net3690),
    .X(_01187_));
 sg13g2_mux2_1 _18040_ (.A0(\spiking_network_top_uut.all_data_out[427] ),
    .A1(net4418),
    .S(net3690),
    .X(_01188_));
 sg13g2_mux2_1 _18041_ (.A0(\spiking_network_top_uut.all_data_out[428] ),
    .A1(net4396),
    .S(net3690),
    .X(_01189_));
 sg13g2_mux2_1 _18042_ (.A0(\spiking_network_top_uut.all_data_out[429] ),
    .A1(net4375),
    .S(net3690),
    .X(_01190_));
 sg13g2_nand2_1 _18043_ (.Y(_03229_),
    .A(net4355),
    .B(net3690));
 sg13g2_o21ai_1 _18044_ (.B1(_03229_),
    .Y(_01191_),
    .A1(_03540_),
    .A2(net3690));
 sg13g2_mux2_1 _18045_ (.A0(\spiking_network_top_uut.all_data_out[431] ),
    .A1(net4336),
    .S(net3690),
    .X(_01192_));
 sg13g2_nor2_2 _18046_ (.A(net3734),
    .B(_03225_),
    .Y(_03230_));
 sg13g2_mux2_1 _18047_ (.A0(\spiking_network_top_uut.all_data_out[552] ),
    .A1(net4477),
    .S(_03230_),
    .X(_01193_));
 sg13g2_mux2_1 _18048_ (.A0(\spiking_network_top_uut.all_data_out[553] ),
    .A1(net4460),
    .S(_03230_),
    .X(_01194_));
 sg13g2_mux2_1 _18049_ (.A0(\spiking_network_top_uut.all_data_out[554] ),
    .A1(net4436),
    .S(_03230_),
    .X(_01195_));
 sg13g2_mux2_1 _18050_ (.A0(\spiking_network_top_uut.all_data_out[555] ),
    .A1(net4417),
    .S(_03230_),
    .X(_01196_));
 sg13g2_mux2_1 _18051_ (.A0(\spiking_network_top_uut.all_data_out[556] ),
    .A1(net4396),
    .S(_03230_),
    .X(_01197_));
 sg13g2_mux2_1 _18052_ (.A0(\spiking_network_top_uut.all_data_out[557] ),
    .A1(net4375),
    .S(_03230_),
    .X(_01198_));
 sg13g2_mux2_1 _18053_ (.A0(\spiking_network_top_uut.all_data_out[558] ),
    .A1(net4355),
    .S(_03230_),
    .X(_01199_));
 sg13g2_mux2_1 _18054_ (.A0(\spiking_network_top_uut.all_data_out[559] ),
    .A1(net4335),
    .S(_03230_),
    .X(_01200_));
 sg13g2_nand2_2 _18055_ (.Y(_03231_),
    .A(_03200_),
    .B(_03207_));
 sg13g2_nor2_2 _18056_ (.A(net3736),
    .B(_03231_),
    .Y(_03232_));
 sg13g2_mux2_1 _18057_ (.A0(\spiking_network_top_uut.all_data_out[416] ),
    .A1(net4475),
    .S(_03232_),
    .X(_01201_));
 sg13g2_mux2_1 _18058_ (.A0(\spiking_network_top_uut.all_data_out[417] ),
    .A1(net4456),
    .S(_03232_),
    .X(_01202_));
 sg13g2_mux2_1 _18059_ (.A0(\spiking_network_top_uut.all_data_out[418] ),
    .A1(net4439),
    .S(_03232_),
    .X(_01203_));
 sg13g2_mux2_1 _18060_ (.A0(\spiking_network_top_uut.all_data_out[419] ),
    .A1(net4419),
    .S(_03232_),
    .X(_01204_));
 sg13g2_mux2_1 _18061_ (.A0(\spiking_network_top_uut.all_data_out[420] ),
    .A1(net4395),
    .S(_03232_),
    .X(_01205_));
 sg13g2_mux2_1 _18062_ (.A0(\spiking_network_top_uut.all_data_out[421] ),
    .A1(net4378),
    .S(_03232_),
    .X(_01206_));
 sg13g2_mux2_1 _18063_ (.A0(\spiking_network_top_uut.all_data_out[422] ),
    .A1(net4354),
    .S(_03232_),
    .X(_01207_));
 sg13g2_mux2_1 _18064_ (.A0(\spiking_network_top_uut.all_data_out[423] ),
    .A1(net4336),
    .S(_03232_),
    .X(_01208_));
 sg13g2_nor2_2 _18065_ (.A(_03218_),
    .B(net3732),
    .Y(_03233_));
 sg13g2_mux2_1 _18066_ (.A0(\spiking_network_top_uut.all_data_out[688] ),
    .A1(net4473),
    .S(_03233_),
    .X(_01209_));
 sg13g2_mux2_1 _18067_ (.A0(\spiking_network_top_uut.all_data_out[689] ),
    .A1(net4452),
    .S(_03233_),
    .X(_01210_));
 sg13g2_mux2_1 _18068_ (.A0(\spiking_network_top_uut.all_data_out[690] ),
    .A1(net4432),
    .S(_03233_),
    .X(_01211_));
 sg13g2_mux2_1 _18069_ (.A0(\spiking_network_top_uut.all_data_out[691] ),
    .A1(net4411),
    .S(_03233_),
    .X(_01212_));
 sg13g2_mux2_1 _18070_ (.A0(\spiking_network_top_uut.all_data_out[692] ),
    .A1(net4394),
    .S(_03233_),
    .X(_01213_));
 sg13g2_mux2_1 _18071_ (.A0(\spiking_network_top_uut.all_data_out[693] ),
    .A1(net4372),
    .S(_03233_),
    .X(_01214_));
 sg13g2_mux2_1 _18072_ (.A0(\spiking_network_top_uut.all_data_out[694] ),
    .A1(net4353),
    .S(_03233_),
    .X(_01215_));
 sg13g2_mux2_1 _18073_ (.A0(\spiking_network_top_uut.all_data_out[695] ),
    .A1(net4334),
    .S(_03233_),
    .X(_01216_));
 sg13g2_and3_2 _18074_ (.X(_03234_),
    .A(net4484),
    .B(net4483),
    .C(_03199_));
 sg13g2_nand3_1 _18075_ (.B(net4483),
    .C(_03199_),
    .A(net4484),
    .Y(_03235_));
 sg13g2_nor2_2 _18076_ (.A(net3736),
    .B(_03235_),
    .Y(_03236_));
 sg13g2_mux2_1 _18077_ (.A0(\spiking_network_top_uut.all_data_out[408] ),
    .A1(net4479),
    .S(_03236_),
    .X(_01217_));
 sg13g2_mux2_1 _18078_ (.A0(\spiking_network_top_uut.all_data_out[409] ),
    .A1(net4459),
    .S(_03236_),
    .X(_01218_));
 sg13g2_mux2_1 _18079_ (.A0(\spiking_network_top_uut.all_data_out[410] ),
    .A1(net4438),
    .S(_03236_),
    .X(_01219_));
 sg13g2_mux2_1 _18080_ (.A0(\spiking_network_top_uut.all_data_out[411] ),
    .A1(net4414),
    .S(_03236_),
    .X(_01220_));
 sg13g2_mux2_1 _18081_ (.A0(\spiking_network_top_uut.all_data_out[412] ),
    .A1(net4398),
    .S(_03236_),
    .X(_01221_));
 sg13g2_mux2_1 _18082_ (.A0(\spiking_network_top_uut.all_data_out[413] ),
    .A1(net4377),
    .S(_03236_),
    .X(_01222_));
 sg13g2_mux2_1 _18083_ (.A0(\spiking_network_top_uut.all_data_out[414] ),
    .A1(net4356),
    .S(_03236_),
    .X(_01223_));
 sg13g2_mux2_1 _18084_ (.A0(\spiking_network_top_uut.all_data_out[415] ),
    .A1(net4332),
    .S(_03236_),
    .X(_01224_));
 sg13g2_nor2_2 _18085_ (.A(\spiking_network_top_uut.spi_inst.LSB_Address_reg[2] ),
    .B(_03212_),
    .Y(_03237_));
 sg13g2_nand2_2 _18086_ (.Y(_03238_),
    .A(_03214_),
    .B(_03237_));
 sg13g2_nor2_2 _18087_ (.A(net3733),
    .B(_03238_),
    .Y(_03239_));
 sg13g2_mux2_1 _18088_ (.A0(\spiking_network_top_uut.all_data_out[584] ),
    .A1(net4476),
    .S(_03239_),
    .X(_01225_));
 sg13g2_mux2_1 _18089_ (.A0(\spiking_network_top_uut.all_data_out[585] ),
    .A1(net4456),
    .S(_03239_),
    .X(_01226_));
 sg13g2_mux2_1 _18090_ (.A0(\spiking_network_top_uut.all_data_out[586] ),
    .A1(net4435),
    .S(_03239_),
    .X(_01227_));
 sg13g2_mux2_1 _18091_ (.A0(\spiking_network_top_uut.all_data_out[587] ),
    .A1(net4417),
    .S(_03239_),
    .X(_01228_));
 sg13g2_mux2_1 _18092_ (.A0(\spiking_network_top_uut.all_data_out[588] ),
    .A1(net4394),
    .S(_03239_),
    .X(_01229_));
 sg13g2_mux2_1 _18093_ (.A0(\spiking_network_top_uut.all_data_out[589] ),
    .A1(net4378),
    .S(_03239_),
    .X(_01230_));
 sg13g2_mux2_1 _18094_ (.A0(\spiking_network_top_uut.all_data_out[590] ),
    .A1(net4353),
    .S(_03239_),
    .X(_01231_));
 sg13g2_mux2_1 _18095_ (.A0(\spiking_network_top_uut.all_data_out[591] ),
    .A1(net4336),
    .S(_03239_),
    .X(_01232_));
 sg13g2_and2_2 _18096_ (.A(net3737),
    .B(_03217_),
    .X(_03240_));
 sg13g2_nand2_2 _18097_ (.Y(_03241_),
    .A(net3737),
    .B(_03217_));
 sg13g2_nor2_2 _18098_ (.A(net3735),
    .B(_03241_),
    .Y(_03242_));
 sg13g2_mux2_1 _18099_ (.A0(\spiking_network_top_uut.all_data_out[400] ),
    .A1(net4475),
    .S(_03242_),
    .X(_01233_));
 sg13g2_mux2_1 _18100_ (.A0(\spiking_network_top_uut.all_data_out[401] ),
    .A1(net4455),
    .S(_03242_),
    .X(_01234_));
 sg13g2_mux2_1 _18101_ (.A0(\spiking_network_top_uut.all_data_out[402] ),
    .A1(net4434),
    .S(_03242_),
    .X(_01235_));
 sg13g2_mux2_1 _18102_ (.A0(\spiking_network_top_uut.all_data_out[403] ),
    .A1(net4414),
    .S(_03242_),
    .X(_01236_));
 sg13g2_mux2_1 _18103_ (.A0(\spiking_network_top_uut.all_data_out[404] ),
    .A1(net4392),
    .S(_03242_),
    .X(_01237_));
 sg13g2_mux2_1 _18104_ (.A0(\spiking_network_top_uut.all_data_out[405] ),
    .A1(net4373),
    .S(_03242_),
    .X(_01238_));
 sg13g2_mux2_1 _18105_ (.A0(\spiking_network_top_uut.all_data_out[406] ),
    .A1(net4351),
    .S(_03242_),
    .X(_01239_));
 sg13g2_mux2_1 _18106_ (.A0(\spiking_network_top_uut.all_data_out[407] ),
    .A1(net4332),
    .S(_03242_),
    .X(_01240_));
 sg13g2_nor2_2 _18107_ (.A(_03208_),
    .B(net3732),
    .Y(_03243_));
 sg13g2_mux2_1 _18108_ (.A0(\spiking_network_top_uut.all_data_out[696] ),
    .A1(net4471),
    .S(_03243_),
    .X(_01241_));
 sg13g2_mux2_1 _18109_ (.A0(\spiking_network_top_uut.all_data_out[697] ),
    .A1(net4450),
    .S(_03243_),
    .X(_01242_));
 sg13g2_mux2_1 _18110_ (.A0(\spiking_network_top_uut.all_data_out[698] ),
    .A1(net4430),
    .S(_03243_),
    .X(_01243_));
 sg13g2_mux2_1 _18111_ (.A0(\spiking_network_top_uut.all_data_out[699] ),
    .A1(net4411),
    .S(_03243_),
    .X(_01244_));
 sg13g2_mux2_1 _18112_ (.A0(\spiking_network_top_uut.all_data_out[700] ),
    .A1(net4388),
    .S(_03243_),
    .X(_01245_));
 sg13g2_mux2_1 _18113_ (.A0(\spiking_network_top_uut.all_data_out[701] ),
    .A1(net4369),
    .S(_03243_),
    .X(_01246_));
 sg13g2_mux2_1 _18114_ (.A0(\spiking_network_top_uut.all_data_out[702] ),
    .A1(net4348),
    .S(_03243_),
    .X(_01247_));
 sg13g2_mux2_1 _18115_ (.A0(\spiking_network_top_uut.all_data_out[703] ),
    .A1(net4331),
    .S(_03243_),
    .X(_01248_));
 sg13g2_and2_2 _18116_ (.A(net3737),
    .B(_03214_),
    .X(_03244_));
 sg13g2_nand2_2 _18117_ (.Y(_03245_),
    .A(_03199_),
    .B(_03214_));
 sg13g2_nor2_2 _18118_ (.A(net3736),
    .B(_03245_),
    .Y(_03246_));
 sg13g2_mux2_1 _18119_ (.A0(\spiking_network_top_uut.all_data_out[392] ),
    .A1(net4480),
    .S(_03246_),
    .X(_01249_));
 sg13g2_mux2_1 _18120_ (.A0(\spiking_network_top_uut.all_data_out[393] ),
    .A1(net4457),
    .S(net3689),
    .X(_01250_));
 sg13g2_mux2_1 _18121_ (.A0(\spiking_network_top_uut.all_data_out[394] ),
    .A1(net4436),
    .S(net3689),
    .X(_01251_));
 sg13g2_mux2_1 _18122_ (.A0(\spiking_network_top_uut.all_data_out[395] ),
    .A1(net4418),
    .S(net3689),
    .X(_01252_));
 sg13g2_mux2_1 _18123_ (.A0(\spiking_network_top_uut.all_data_out[396] ),
    .A1(net4396),
    .S(net3689),
    .X(_01253_));
 sg13g2_mux2_1 _18124_ (.A0(\spiking_network_top_uut.all_data_out[397] ),
    .A1(net4375),
    .S(net3689),
    .X(_01254_));
 sg13g2_nand2_1 _18125_ (.Y(_03247_),
    .A(net4355),
    .B(net3689));
 sg13g2_o21ai_1 _18126_ (.B1(_03247_),
    .Y(_01255_),
    .A1(_03542_),
    .A2(net3689));
 sg13g2_mux2_1 _18127_ (.A0(\spiking_network_top_uut.all_data_out[399] ),
    .A1(net4335),
    .S(net3689),
    .X(_01256_));
 sg13g2_nor2_2 _18128_ (.A(net3733),
    .B(_03231_),
    .Y(_03248_));
 sg13g2_mux2_1 _18129_ (.A0(\spiking_network_top_uut.all_data_out[544] ),
    .A1(net4478),
    .S(_03248_),
    .X(_01257_));
 sg13g2_mux2_1 _18130_ (.A0(\spiking_network_top_uut.all_data_out[545] ),
    .A1(net4458),
    .S(_03248_),
    .X(_01258_));
 sg13g2_mux2_1 _18131_ (.A0(\spiking_network_top_uut.all_data_out[546] ),
    .A1(net4439),
    .S(_03248_),
    .X(_01259_));
 sg13g2_mux2_1 _18132_ (.A0(\spiking_network_top_uut.all_data_out[547] ),
    .A1(net4420),
    .S(_03248_),
    .X(_01260_));
 sg13g2_mux2_1 _18133_ (.A0(\spiking_network_top_uut.all_data_out[548] ),
    .A1(net4395),
    .S(_03248_),
    .X(_01261_));
 sg13g2_mux2_1 _18134_ (.A0(\spiking_network_top_uut.all_data_out[549] ),
    .A1(net4378),
    .S(_03248_),
    .X(_01262_));
 sg13g2_mux2_1 _18135_ (.A0(\spiking_network_top_uut.all_data_out[550] ),
    .A1(net4354),
    .S(_03248_),
    .X(_01263_));
 sg13g2_mux2_1 _18136_ (.A0(\spiking_network_top_uut.all_data_out[551] ),
    .A1(net4336),
    .S(_03248_),
    .X(_01264_));
 sg13g2_nor2_2 _18137_ (.A(_03201_),
    .B(net3735),
    .Y(_03249_));
 sg13g2_mux2_1 _18138_ (.A0(\spiking_network_top_uut.all_data_out[384] ),
    .A1(net4478),
    .S(_03249_),
    .X(_01265_));
 sg13g2_mux2_1 _18139_ (.A0(\spiking_network_top_uut.all_data_out[385] ),
    .A1(net4458),
    .S(_03249_),
    .X(_01266_));
 sg13g2_mux2_1 _18140_ (.A0(\spiking_network_top_uut.all_data_out[386] ),
    .A1(net4437),
    .S(_03249_),
    .X(_01267_));
 sg13g2_mux2_1 _18141_ (.A0(\spiking_network_top_uut.all_data_out[387] ),
    .A1(net4408),
    .S(_03249_),
    .X(_01268_));
 sg13g2_mux2_1 _18142_ (.A0(\spiking_network_top_uut.all_data_out[388] ),
    .A1(net4397),
    .S(_03249_),
    .X(_01269_));
 sg13g2_mux2_1 _18143_ (.A0(\spiking_network_top_uut.all_data_out[389] ),
    .A1(net4376),
    .S(_03249_),
    .X(_01270_));
 sg13g2_mux2_1 _18144_ (.A0(\spiking_network_top_uut.all_data_out[390] ),
    .A1(net4357),
    .S(_03249_),
    .X(_01271_));
 sg13g2_mux2_1 _18145_ (.A0(\spiking_network_top_uut.all_data_out[391] ),
    .A1(net4326),
    .S(_03249_),
    .X(_01272_));
 sg13g2_nand2_2 _18146_ (.Y(_03250_),
    .A(_03200_),
    .B(_03237_));
 sg13g2_nor2_2 _18147_ (.A(net3731),
    .B(_03250_),
    .Y(_03251_));
 sg13g2_mux2_1 _18148_ (.A0(\spiking_network_top_uut.all_data_out[704] ),
    .A1(net4465),
    .S(_03251_),
    .X(_01273_));
 sg13g2_mux2_1 _18149_ (.A0(\spiking_network_top_uut.all_data_out[705] ),
    .A1(net4445),
    .S(_03251_),
    .X(_01274_));
 sg13g2_mux2_1 _18150_ (.A0(\spiking_network_top_uut.all_data_out[706] ),
    .A1(net4424),
    .S(_03251_),
    .X(_01275_));
 sg13g2_mux2_1 _18151_ (.A0(\spiking_network_top_uut.all_data_out[707] ),
    .A1(net4406),
    .S(_03251_),
    .X(_01276_));
 sg13g2_mux2_1 _18152_ (.A0(\spiking_network_top_uut.all_data_out[708] ),
    .A1(net4382),
    .S(_03251_),
    .X(_01277_));
 sg13g2_mux2_1 _18153_ (.A0(\spiking_network_top_uut.all_data_out[709] ),
    .A1(net4362),
    .S(_03251_),
    .X(_01278_));
 sg13g2_mux2_1 _18154_ (.A0(\spiking_network_top_uut.all_data_out[710] ),
    .A1(net4342),
    .S(_03251_),
    .X(_01279_));
 sg13g2_mux2_1 _18155_ (.A0(\spiking_network_top_uut.all_data_out[711] ),
    .A1(net4321),
    .S(_03251_),
    .X(_01280_));
 sg13g2_nor2b_1 _18156_ (.A(\spiking_network_top_uut.spi_inst.LSB_Address_reg[4] ),
    .B_N(\spiking_network_top_uut.spi_inst.LSB_Address_reg[5] ),
    .Y(_03252_));
 sg13g2_nand2b_1 _18157_ (.Y(_03253_),
    .B(\spiking_network_top_uut.spi_inst.LSB_Address_reg[5] ),
    .A_N(\spiking_network_top_uut.spi_inst.LSB_Address_reg[4] ));
 sg13g2_nor2_2 _18158_ (.A(\spiking_network_top_uut.spi_inst.LSB_Address_reg[6] ),
    .B(_03253_),
    .Y(_03254_));
 sg13g2_nand2b_2 _18159_ (.Y(_03255_),
    .B(_03252_),
    .A_N(\spiking_network_top_uut.spi_inst.LSB_Address_reg[6] ));
 sg13g2_nand3_1 _18160_ (.B(net4483),
    .C(_03213_),
    .A(net4484),
    .Y(_03256_));
 sg13g2_nor2_2 _18161_ (.A(net3729),
    .B(net15),
    .Y(_03257_));
 sg13g2_mux2_1 _18162_ (.A0(\spiking_network_top_uut.all_data_out[376] ),
    .A1(net4478),
    .S(_03257_),
    .X(_01281_));
 sg13g2_mux2_1 _18163_ (.A0(\spiking_network_top_uut.all_data_out[377] ),
    .A1(net4459),
    .S(_03257_),
    .X(_01282_));
 sg13g2_mux2_1 _18164_ (.A0(\spiking_network_top_uut.all_data_out[378] ),
    .A1(net4437),
    .S(_03257_),
    .X(_01283_));
 sg13g2_mux2_1 _18165_ (.A0(\spiking_network_top_uut.all_data_out[379] ),
    .A1(net4408),
    .S(_03257_),
    .X(_01284_));
 sg13g2_mux2_1 _18166_ (.A0(\spiking_network_top_uut.all_data_out[380] ),
    .A1(net4398),
    .S(_03257_),
    .X(_01285_));
 sg13g2_mux2_1 _18167_ (.A0(\spiking_network_top_uut.all_data_out[381] ),
    .A1(net4377),
    .S(_03257_),
    .X(_01286_));
 sg13g2_mux2_1 _18168_ (.A0(\spiking_network_top_uut.all_data_out[382] ),
    .A1(net4358),
    .S(_03257_),
    .X(_01287_));
 sg13g2_mux2_1 _18169_ (.A0(\spiking_network_top_uut.all_data_out[383] ),
    .A1(net4326),
    .S(_03257_),
    .X(_01288_));
 sg13g2_nand2_2 _18170_ (.Y(_03258_),
    .A(_03213_),
    .B(_03217_));
 sg13g2_nor2_1 _18171_ (.A(net3733),
    .B(_03258_),
    .Y(_03259_));
 sg13g2_mux2_1 _18172_ (.A0(\spiking_network_top_uut.all_data_out[624] ),
    .A1(net4473),
    .S(net3688),
    .X(_01289_));
 sg13g2_mux2_1 _18173_ (.A0(\spiking_network_top_uut.all_data_out[625] ),
    .A1(net4456),
    .S(_03259_),
    .X(_01290_));
 sg13g2_mux2_1 _18174_ (.A0(\spiking_network_top_uut.all_data_out[626] ),
    .A1(net4432),
    .S(net3688),
    .X(_01291_));
 sg13g2_mux2_1 _18175_ (.A0(\spiking_network_top_uut.all_data_out[627] ),
    .A1(net4416),
    .S(net3688),
    .X(_01292_));
 sg13g2_mux2_1 _18176_ (.A0(\spiking_network_top_uut.all_data_out[628] ),
    .A1(net4394),
    .S(net3688),
    .X(_01293_));
 sg13g2_mux2_1 _18177_ (.A0(\spiking_network_top_uut.all_data_out[629] ),
    .A1(net4378),
    .S(net3688),
    .X(_01294_));
 sg13g2_nand2_1 _18178_ (.Y(_03260_),
    .A(net4353),
    .B(net3688));
 sg13g2_o21ai_1 _18179_ (.B1(_03260_),
    .Y(_01295_),
    .A1(_03530_),
    .A2(net3688));
 sg13g2_mux2_1 _18180_ (.A0(\spiking_network_top_uut.all_data_out[631] ),
    .A1(net4334),
    .S(net3688),
    .X(_01296_));
 sg13g2_nor2_1 _18181_ (.A(net3730),
    .B(_03258_),
    .Y(_03261_));
 sg13g2_mux2_1 _18182_ (.A0(\spiking_network_top_uut.all_data_out[368] ),
    .A1(net4475),
    .S(net3687),
    .X(_01297_));
 sg13g2_mux2_1 _18183_ (.A0(\spiking_network_top_uut.all_data_out[369] ),
    .A1(net4455),
    .S(net3687),
    .X(_01298_));
 sg13g2_mux2_1 _18184_ (.A0(\spiking_network_top_uut.all_data_out[370] ),
    .A1(net4434),
    .S(net3687),
    .X(_01299_));
 sg13g2_mux2_1 _18185_ (.A0(\spiking_network_top_uut.all_data_out[371] ),
    .A1(net4419),
    .S(_03261_),
    .X(_01300_));
 sg13g2_mux2_1 _18186_ (.A0(\spiking_network_top_uut.all_data_out[372] ),
    .A1(net4392),
    .S(net3687),
    .X(_01301_));
 sg13g2_mux2_1 _18187_ (.A0(\spiking_network_top_uut.all_data_out[373] ),
    .A1(net4373),
    .S(net3687),
    .X(_01302_));
 sg13g2_nand2_1 _18188_ (.Y(_03262_),
    .A(net4351),
    .B(net3687));
 sg13g2_o21ai_1 _18189_ (.B1(_03262_),
    .Y(_01303_),
    .A1(_03545_),
    .A2(net3687));
 sg13g2_mux2_1 _18190_ (.A0(\spiking_network_top_uut.all_data_out[375] ),
    .A1(net4332),
    .S(net3687),
    .X(_01304_));
 sg13g2_nor2_2 _18191_ (.A(net3731),
    .B(_03238_),
    .Y(_03263_));
 sg13g2_mux2_1 _18192_ (.A0(\spiking_network_top_uut.all_data_out[712] ),
    .A1(net4476),
    .S(net3686),
    .X(_01305_));
 sg13g2_mux2_1 _18193_ (.A0(\spiking_network_top_uut.all_data_out[713] ),
    .A1(net4457),
    .S(_03263_),
    .X(_01306_));
 sg13g2_mux2_1 _18194_ (.A0(\spiking_network_top_uut.all_data_out[714] ),
    .A1(net4435),
    .S(net3686),
    .X(_01307_));
 sg13g2_mux2_1 _18195_ (.A0(\spiking_network_top_uut.all_data_out[715] ),
    .A1(net4413),
    .S(net3686),
    .X(_01308_));
 sg13g2_mux2_1 _18196_ (.A0(\spiking_network_top_uut.all_data_out[716] ),
    .A1(net4395),
    .S(net3686),
    .X(_01309_));
 sg13g2_mux2_1 _18197_ (.A0(\spiking_network_top_uut.all_data_out[717] ),
    .A1(net4372),
    .S(net3686),
    .X(_01310_));
 sg13g2_nand2_1 _18198_ (.Y(_03264_),
    .A(net4354),
    .B(net3686));
 sg13g2_o21ai_1 _18199_ (.B1(_03264_),
    .Y(_01311_),
    .A1(_03523_),
    .A2(net3686));
 sg13g2_mux2_1 _18200_ (.A0(\spiking_network_top_uut.all_data_out[719] ),
    .A1(net4333),
    .S(net3686),
    .X(_01312_));
 sg13g2_nor2_2 _18201_ (.A(_03215_),
    .B(net3730),
    .Y(_03265_));
 sg13g2_mux2_1 _18202_ (.A0(\spiking_network_top_uut.all_data_out[360] ),
    .A1(net4477),
    .S(_03265_),
    .X(_01313_));
 sg13g2_mux2_1 _18203_ (.A0(\spiking_network_top_uut.all_data_out[361] ),
    .A1(net4460),
    .S(_03265_),
    .X(_01314_));
 sg13g2_mux2_1 _18204_ (.A0(\spiking_network_top_uut.all_data_out[362] ),
    .A1(net4438),
    .S(_03265_),
    .X(_01315_));
 sg13g2_mux2_1 _18205_ (.A0(\spiking_network_top_uut.all_data_out[363] ),
    .A1(net4417),
    .S(_03265_),
    .X(_01316_));
 sg13g2_mux2_1 _18206_ (.A0(\spiking_network_top_uut.all_data_out[364] ),
    .A1(net4396),
    .S(_03265_),
    .X(_01317_));
 sg13g2_mux2_1 _18207_ (.A0(\spiking_network_top_uut.all_data_out[365] ),
    .A1(net4375),
    .S(_03265_),
    .X(_01318_));
 sg13g2_mux2_1 _18208_ (.A0(\spiking_network_top_uut.all_data_out[366] ),
    .A1(net4355),
    .S(_03265_),
    .X(_01319_));
 sg13g2_mux2_1 _18209_ (.A0(\spiking_network_top_uut.all_data_out[367] ),
    .A1(net4335),
    .S(_03265_),
    .X(_01320_));
 sg13g2_nor2_2 _18210_ (.A(net3733),
    .B(_03235_),
    .Y(_03266_));
 sg13g2_mux2_1 _18211_ (.A0(\spiking_network_top_uut.all_data_out[536] ),
    .A1(net4479),
    .S(_03266_),
    .X(_01321_));
 sg13g2_mux2_1 _18212_ (.A0(\spiking_network_top_uut.all_data_out[537] ),
    .A1(net4459),
    .S(net3685),
    .X(_01322_));
 sg13g2_nand2_1 _18213_ (.Y(_03267_),
    .A(net4437),
    .B(net3685));
 sg13g2_o21ai_1 _18214_ (.B1(_03267_),
    .Y(_01323_),
    .A1(_03612_),
    .A2(net3685));
 sg13g2_mux2_1 _18215_ (.A0(\spiking_network_top_uut.all_data_out[539] ),
    .A1(net4414),
    .S(net3685),
    .X(_01324_));
 sg13g2_mux2_1 _18216_ (.A0(\spiking_network_top_uut.all_data_out[540] ),
    .A1(net4397),
    .S(net3685),
    .X(_01325_));
 sg13g2_mux2_1 _18217_ (.A0(\spiking_network_top_uut.all_data_out[541] ),
    .A1(net4376),
    .S(net3685),
    .X(_01326_));
 sg13g2_mux2_1 _18218_ (.A0(\spiking_network_top_uut.all_data_out[542] ),
    .A1(net4356),
    .S(net3685),
    .X(_01327_));
 sg13g2_mux2_1 _18219_ (.A0(\spiking_network_top_uut.all_data_out[543] ),
    .A1(net4332),
    .S(net3685),
    .X(_01328_));
 sg13g2_nand2_2 _18220_ (.Y(_03268_),
    .A(_03200_),
    .B(_03213_));
 sg13g2_nor2_2 _18221_ (.A(net3730),
    .B(_03268_),
    .Y(_03269_));
 sg13g2_mux2_1 _18222_ (.A0(\spiking_network_top_uut.all_data_out[352] ),
    .A1(net4478),
    .S(_03269_),
    .X(_01329_));
 sg13g2_mux2_1 _18223_ (.A0(\spiking_network_top_uut.all_data_out[353] ),
    .A1(net4458),
    .S(_03269_),
    .X(_01330_));
 sg13g2_mux2_1 _18224_ (.A0(\spiking_network_top_uut.all_data_out[354] ),
    .A1(net4434),
    .S(_03269_),
    .X(_01331_));
 sg13g2_mux2_1 _18225_ (.A0(\spiking_network_top_uut.all_data_out[355] ),
    .A1(net4419),
    .S(_03269_),
    .X(_01332_));
 sg13g2_mux2_1 _18226_ (.A0(\spiking_network_top_uut.all_data_out[356] ),
    .A1(net4398),
    .S(_03269_),
    .X(_01333_));
 sg13g2_mux2_1 _18227_ (.A0(\spiking_network_top_uut.all_data_out[357] ),
    .A1(net4377),
    .S(_03269_),
    .X(_01334_));
 sg13g2_mux2_1 _18228_ (.A0(\spiking_network_top_uut.all_data_out[358] ),
    .A1(net4358),
    .S(_03269_),
    .X(_01335_));
 sg13g2_mux2_1 _18229_ (.A0(\spiking_network_top_uut.all_data_out[359] ),
    .A1(net4329),
    .S(_03269_),
    .X(_01336_));
 sg13g2_nand2_2 _18230_ (.Y(_03270_),
    .A(_03217_),
    .B(_03237_));
 sg13g2_nor2_2 _18231_ (.A(net3732),
    .B(_03270_),
    .Y(_03271_));
 sg13g2_mux2_1 _18232_ (.A0(\spiking_network_top_uut.all_data_out[720] ),
    .A1(net4473),
    .S(_03271_),
    .X(_01337_));
 sg13g2_mux2_1 _18233_ (.A0(\spiking_network_top_uut.all_data_out[721] ),
    .A1(net4452),
    .S(_03271_),
    .X(_01338_));
 sg13g2_mux2_1 _18234_ (.A0(\spiking_network_top_uut.all_data_out[722] ),
    .A1(net4432),
    .S(_03271_),
    .X(_01339_));
 sg13g2_mux2_1 _18235_ (.A0(\spiking_network_top_uut.all_data_out[723] ),
    .A1(net4413),
    .S(_03271_),
    .X(_01340_));
 sg13g2_mux2_1 _18236_ (.A0(\spiking_network_top_uut.all_data_out[724] ),
    .A1(net4392),
    .S(_03271_),
    .X(_01341_));
 sg13g2_mux2_1 _18237_ (.A0(\spiking_network_top_uut.all_data_out[725] ),
    .A1(net4373),
    .S(_03271_),
    .X(_01342_));
 sg13g2_mux2_1 _18238_ (.A0(\spiking_network_top_uut.all_data_out[726] ),
    .A1(net4351),
    .S(_03271_),
    .X(_01343_));
 sg13g2_mux2_1 _18239_ (.A0(\spiking_network_top_uut.all_data_out[727] ),
    .A1(net4334),
    .S(_03271_),
    .X(_01344_));
 sg13g2_nand3_1 _18240_ (.B(net4483),
    .C(_03237_),
    .A(net4484),
    .Y(_03272_));
 sg13g2_nor2_2 _18241_ (.A(net3730),
    .B(_03272_),
    .Y(_03273_));
 sg13g2_mux2_1 _18242_ (.A0(\spiking_network_top_uut.all_data_out[344] ),
    .A1(net4479),
    .S(_03273_),
    .X(_01345_));
 sg13g2_mux2_1 _18243_ (.A0(\spiking_network_top_uut.all_data_out[345] ),
    .A1(net4459),
    .S(_03273_),
    .X(_01346_));
 sg13g2_mux2_1 _18244_ (.A0(\spiking_network_top_uut.all_data_out[346] ),
    .A1(net4438),
    .S(_03273_),
    .X(_01347_));
 sg13g2_mux2_1 _18245_ (.A0(\spiking_network_top_uut.all_data_out[347] ),
    .A1(net4419),
    .S(_03273_),
    .X(_01348_));
 sg13g2_mux2_1 _18246_ (.A0(\spiking_network_top_uut.all_data_out[348] ),
    .A1(net4397),
    .S(_03273_),
    .X(_01349_));
 sg13g2_mux2_1 _18247_ (.A0(\spiking_network_top_uut.all_data_out[349] ),
    .A1(net4376),
    .S(_03273_),
    .X(_01350_));
 sg13g2_mux2_1 _18248_ (.A0(\spiking_network_top_uut.all_data_out[350] ),
    .A1(net4356),
    .S(_03273_),
    .X(_01351_));
 sg13g2_mux2_1 _18249_ (.A0(\spiking_network_top_uut.all_data_out[351] ),
    .A1(net4336),
    .S(_03273_),
    .X(_01352_));
 sg13g2_nor2_2 _18250_ (.A(net3733),
    .B(_03270_),
    .Y(_03274_));
 sg13g2_mux2_1 _18251_ (.A0(\spiking_network_top_uut.all_data_out[592] ),
    .A1(net4473),
    .S(_03274_),
    .X(_01353_));
 sg13g2_mux2_1 _18252_ (.A0(\spiking_network_top_uut.all_data_out[593] ),
    .A1(net4452),
    .S(_03274_),
    .X(_01354_));
 sg13g2_mux2_1 _18253_ (.A0(\spiking_network_top_uut.all_data_out[594] ),
    .A1(net4432),
    .S(_03274_),
    .X(_01355_));
 sg13g2_mux2_1 _18254_ (.A0(\spiking_network_top_uut.all_data_out[595] ),
    .A1(net4413),
    .S(_03274_),
    .X(_01356_));
 sg13g2_mux2_1 _18255_ (.A0(\spiking_network_top_uut.all_data_out[596] ),
    .A1(net4394),
    .S(_03274_),
    .X(_01357_));
 sg13g2_mux2_1 _18256_ (.A0(\spiking_network_top_uut.all_data_out[597] ),
    .A1(net4372),
    .S(_03274_),
    .X(_01358_));
 sg13g2_mux2_1 _18257_ (.A0(\spiking_network_top_uut.all_data_out[598] ),
    .A1(net4353),
    .S(_03274_),
    .X(_01359_));
 sg13g2_mux2_1 _18258_ (.A0(\spiking_network_top_uut.all_data_out[599] ),
    .A1(net4331),
    .S(_03274_),
    .X(_01360_));
 sg13g2_nor2_2 _18259_ (.A(net3729),
    .B(_03270_),
    .Y(_03275_));
 sg13g2_mux2_1 _18260_ (.A0(\spiking_network_top_uut.all_data_out[336] ),
    .A1(net4475),
    .S(_03275_),
    .X(_01361_));
 sg13g2_mux2_1 _18261_ (.A0(\spiking_network_top_uut.all_data_out[337] ),
    .A1(net4455),
    .S(_03275_),
    .X(_01362_));
 sg13g2_mux2_1 _18262_ (.A0(\spiking_network_top_uut.all_data_out[338] ),
    .A1(net4434),
    .S(_03275_),
    .X(_01363_));
 sg13g2_mux2_1 _18263_ (.A0(\spiking_network_top_uut.all_data_out[339] ),
    .A1(net4419),
    .S(_03275_),
    .X(_01364_));
 sg13g2_mux2_1 _18264_ (.A0(\spiking_network_top_uut.all_data_out[340] ),
    .A1(net4390),
    .S(_03275_),
    .X(_01365_));
 sg13g2_mux2_1 _18265_ (.A0(\spiking_network_top_uut.all_data_out[341] ),
    .A1(net4370),
    .S(_03275_),
    .X(_01366_));
 sg13g2_mux2_1 _18266_ (.A0(\spiking_network_top_uut.all_data_out[342] ),
    .A1(net4349),
    .S(_03275_),
    .X(_01367_));
 sg13g2_mux2_1 _18267_ (.A0(\spiking_network_top_uut.all_data_out[343] ),
    .A1(net4330),
    .S(_03275_),
    .X(_01368_));
 sg13g2_nor2_1 _18268_ (.A(net3731),
    .B(net14),
    .Y(_03276_));
 sg13g2_mux2_1 _18269_ (.A0(\spiking_network_top_uut.all_data_out[728] ),
    .A1(net4471),
    .S(net3684),
    .X(_01369_));
 sg13g2_mux2_1 _18270_ (.A0(\spiking_network_top_uut.all_data_out[729] ),
    .A1(net4450),
    .S(net3684),
    .X(_01370_));
 sg13g2_mux2_1 _18271_ (.A0(\spiking_network_top_uut.all_data_out[730] ),
    .A1(net4430),
    .S(net3684),
    .X(_01371_));
 sg13g2_mux2_1 _18272_ (.A0(\spiking_network_top_uut.all_data_out[731] ),
    .A1(net4411),
    .S(net3684),
    .X(_01372_));
 sg13g2_mux2_1 _18273_ (.A0(\spiking_network_top_uut.all_data_out[732] ),
    .A1(net4389),
    .S(_03276_),
    .X(_01373_));
 sg13g2_mux2_1 _18274_ (.A0(\spiking_network_top_uut.all_data_out[733] ),
    .A1(net4369),
    .S(net3684),
    .X(_01374_));
 sg13g2_nand2_1 _18275_ (.Y(_03277_),
    .A(net4347),
    .B(net3684));
 sg13g2_o21ai_1 _18276_ (.B1(_03277_),
    .Y(_01375_),
    .A1(_03520_),
    .A2(net3684));
 sg13g2_mux2_1 _18277_ (.A0(\spiking_network_top_uut.all_data_out[735] ),
    .A1(net4325),
    .S(net3684),
    .X(_01376_));
 sg13g2_nor2_2 _18278_ (.A(_03238_),
    .B(net3729),
    .Y(_03278_));
 sg13g2_mux2_1 _18279_ (.A0(\spiking_network_top_uut.all_data_out[328] ),
    .A1(net4477),
    .S(_03278_),
    .X(_01377_));
 sg13g2_mux2_1 _18280_ (.A0(\spiking_network_top_uut.all_data_out[329] ),
    .A1(net4457),
    .S(_03278_),
    .X(_01378_));
 sg13g2_mux2_1 _18281_ (.A0(\spiking_network_top_uut.all_data_out[330] ),
    .A1(net4436),
    .S(_03278_),
    .X(_01379_));
 sg13g2_mux2_1 _18282_ (.A0(\spiking_network_top_uut.all_data_out[331] ),
    .A1(net4417),
    .S(_03278_),
    .X(_01380_));
 sg13g2_mux2_1 _18283_ (.A0(\spiking_network_top_uut.all_data_out[332] ),
    .A1(net4396),
    .S(_03278_),
    .X(_01381_));
 sg13g2_mux2_1 _18284_ (.A0(\spiking_network_top_uut.all_data_out[333] ),
    .A1(net4375),
    .S(_03278_),
    .X(_01382_));
 sg13g2_mux2_1 _18285_ (.A0(\spiking_network_top_uut.all_data_out[334] ),
    .A1(net4355),
    .S(_03278_),
    .X(_01383_));
 sg13g2_mux2_1 _18286_ (.A0(\spiking_network_top_uut.all_data_out[335] ),
    .A1(net4335),
    .S(_03278_),
    .X(_01384_));
 sg13g2_nor2_2 _18287_ (.A(net3733),
    .B(_03241_),
    .Y(_03279_));
 sg13g2_mux2_1 _18288_ (.A0(\spiking_network_top_uut.all_data_out[528] ),
    .A1(net4474),
    .S(_03279_),
    .X(_01385_));
 sg13g2_mux2_1 _18289_ (.A0(\spiking_network_top_uut.all_data_out[529] ),
    .A1(net4453),
    .S(_03279_),
    .X(_01386_));
 sg13g2_mux2_1 _18290_ (.A0(\spiking_network_top_uut.all_data_out[530] ),
    .A1(net4433),
    .S(_03279_),
    .X(_01387_));
 sg13g2_mux2_1 _18291_ (.A0(\spiking_network_top_uut.all_data_out[531] ),
    .A1(net4410),
    .S(_03279_),
    .X(_01388_));
 sg13g2_mux2_1 _18292_ (.A0(\spiking_network_top_uut.all_data_out[532] ),
    .A1(net4393),
    .S(_03279_),
    .X(_01389_));
 sg13g2_mux2_1 _18293_ (.A0(\spiking_network_top_uut.all_data_out[533] ),
    .A1(net4373),
    .S(_03279_),
    .X(_01390_));
 sg13g2_mux2_1 _18294_ (.A0(\spiking_network_top_uut.all_data_out[534] ),
    .A1(net4351),
    .S(_03279_),
    .X(_01391_));
 sg13g2_mux2_1 _18295_ (.A0(\spiking_network_top_uut.all_data_out[535] ),
    .A1(net4330),
    .S(_03279_),
    .X(_01392_));
 sg13g2_nor2_2 _18296_ (.A(_03250_),
    .B(net3729),
    .Y(_03280_));
 sg13g2_mux2_1 _18297_ (.A0(\spiking_network_top_uut.all_data_out[320] ),
    .A1(net4478),
    .S(_03280_),
    .X(_01393_));
 sg13g2_mux2_1 _18298_ (.A0(\spiking_network_top_uut.all_data_out[321] ),
    .A1(net4458),
    .S(_03280_),
    .X(_01394_));
 sg13g2_mux2_1 _18299_ (.A0(\spiking_network_top_uut.all_data_out[322] ),
    .A1(net4437),
    .S(_03280_),
    .X(_01395_));
 sg13g2_mux2_1 _18300_ (.A0(\spiking_network_top_uut.all_data_out[323] ),
    .A1(net4419),
    .S(_03280_),
    .X(_01396_));
 sg13g2_mux2_1 _18301_ (.A0(\spiking_network_top_uut.all_data_out[324] ),
    .A1(net4398),
    .S(_03280_),
    .X(_01397_));
 sg13g2_mux2_1 _18302_ (.A0(\spiking_network_top_uut.all_data_out[325] ),
    .A1(net4377),
    .S(_03280_),
    .X(_01398_));
 sg13g2_mux2_1 _18303_ (.A0(\spiking_network_top_uut.all_data_out[326] ),
    .A1(net4358),
    .S(_03280_),
    .X(_01399_));
 sg13g2_mux2_1 _18304_ (.A0(\spiking_network_top_uut.all_data_out[327] ),
    .A1(net4336),
    .S(_03280_),
    .X(_01400_));
 sg13g2_nor2_2 _18305_ (.A(net3731),
    .B(_03268_),
    .Y(_03281_));
 sg13g2_mux2_1 _18306_ (.A0(\spiking_network_top_uut.all_data_out[736] ),
    .A1(net4468),
    .S(_03281_),
    .X(_01401_));
 sg13g2_mux2_1 _18307_ (.A0(\spiking_network_top_uut.all_data_out[737] ),
    .A1(net4446),
    .S(_03281_),
    .X(_01402_));
 sg13g2_mux2_1 _18308_ (.A0(\spiking_network_top_uut.all_data_out[738] ),
    .A1(net4426),
    .S(_03281_),
    .X(_01403_));
 sg13g2_mux2_1 _18309_ (.A0(\spiking_network_top_uut.all_data_out[739] ),
    .A1(net4403),
    .S(_03281_),
    .X(_01404_));
 sg13g2_mux2_1 _18310_ (.A0(\spiking_network_top_uut.all_data_out[740] ),
    .A1(net4383),
    .S(_03281_),
    .X(_01405_));
 sg13g2_mux2_1 _18311_ (.A0(\spiking_network_top_uut.all_data_out[741] ),
    .A1(net4362),
    .S(_03281_),
    .X(_01406_));
 sg13g2_mux2_1 _18312_ (.A0(\spiking_network_top_uut.all_data_out[742] ),
    .A1(net4346),
    .S(_03281_),
    .X(_01407_));
 sg13g2_mux2_1 _18313_ (.A0(\spiking_network_top_uut.all_data_out[743] ),
    .A1(net4321),
    .S(_03281_),
    .X(_01408_));
 sg13g2_nor2_2 _18314_ (.A(_03208_),
    .B(net3729),
    .Y(_03282_));
 sg13g2_mux2_1 _18315_ (.A0(\spiking_network_top_uut.all_data_out[312] ),
    .A1(net4462),
    .S(_03282_),
    .X(_01409_));
 sg13g2_mux2_1 _18316_ (.A0(\spiking_network_top_uut.all_data_out[313] ),
    .A1(net4441),
    .S(_03282_),
    .X(_01410_));
 sg13g2_mux2_1 _18317_ (.A0(\spiking_network_top_uut.all_data_out[314] ),
    .A1(net4422),
    .S(_03282_),
    .X(_01411_));
 sg13g2_mux2_1 _18318_ (.A0(\spiking_network_top_uut.all_data_out[315] ),
    .A1(net4402),
    .S(_03282_),
    .X(_01412_));
 sg13g2_mux2_1 _18319_ (.A0(\spiking_network_top_uut.all_data_out[316] ),
    .A1(net4380),
    .S(_03282_),
    .X(_01413_));
 sg13g2_mux2_1 _18320_ (.A0(\spiking_network_top_uut.all_data_out[317] ),
    .A1(net4360),
    .S(_03282_),
    .X(_01414_));
 sg13g2_mux2_1 _18321_ (.A0(\spiking_network_top_uut.all_data_out[318] ),
    .A1(net4339),
    .S(_03282_),
    .X(_01415_));
 sg13g2_mux2_1 _18322_ (.A0(\spiking_network_top_uut.all_data_out[319] ),
    .A1(net4324),
    .S(_03282_),
    .X(_01416_));
 sg13g2_nor2_2 _18323_ (.A(net3734),
    .B(_03256_),
    .Y(_03283_));
 sg13g2_mux2_1 _18324_ (.A0(\spiking_network_top_uut.all_data_out[632] ),
    .A1(net4467),
    .S(net3683),
    .X(_01417_));
 sg13g2_mux2_1 _18325_ (.A0(\spiking_network_top_uut.all_data_out[633] ),
    .A1(net4446),
    .S(net3683),
    .X(_01418_));
 sg13g2_nand2_1 _18326_ (.Y(_03284_),
    .A(net4427),
    .B(net3683));
 sg13g2_o21ai_1 _18327_ (.B1(_03284_),
    .Y(_01419_),
    .A1(_03603_),
    .A2(net3683));
 sg13g2_mux2_1 _18328_ (.A0(\spiking_network_top_uut.all_data_out[635] ),
    .A1(net4409),
    .S(net3683),
    .X(_01420_));
 sg13g2_mux2_1 _18329_ (.A0(\spiking_network_top_uut.all_data_out[636] ),
    .A1(net4389),
    .S(_03283_),
    .X(_01421_));
 sg13g2_mux2_1 _18330_ (.A0(\spiking_network_top_uut.all_data_out[637] ),
    .A1(net4370),
    .S(net3683),
    .X(_01422_));
 sg13g2_mux2_1 _18331_ (.A0(\spiking_network_top_uut.all_data_out[638] ),
    .A1(net4348),
    .S(net3683),
    .X(_01423_));
 sg13g2_mux2_1 _18332_ (.A0(\spiking_network_top_uut.all_data_out[639] ),
    .A1(net4323),
    .S(net3683),
    .X(_01424_));
 sg13g2_nor2_2 _18333_ (.A(_03218_),
    .B(net3729),
    .Y(_03285_));
 sg13g2_mux2_1 _18334_ (.A0(\spiking_network_top_uut.all_data_out[304] ),
    .A1(net4462),
    .S(_03285_),
    .X(_01425_));
 sg13g2_mux2_1 _18335_ (.A0(\spiking_network_top_uut.all_data_out[305] ),
    .A1(net4442),
    .S(_03285_),
    .X(_01426_));
 sg13g2_mux2_1 _18336_ (.A0(\spiking_network_top_uut.all_data_out[306] ),
    .A1(net4423),
    .S(_03285_),
    .X(_01427_));
 sg13g2_mux2_1 _18337_ (.A0(\spiking_network_top_uut.all_data_out[307] ),
    .A1(net4401),
    .S(_03285_),
    .X(_01428_));
 sg13g2_mux2_1 _18338_ (.A0(\spiking_network_top_uut.all_data_out[308] ),
    .A1(net4380),
    .S(_03285_),
    .X(_01429_));
 sg13g2_mux2_1 _18339_ (.A0(\spiking_network_top_uut.all_data_out[309] ),
    .A1(net4360),
    .S(_03285_),
    .X(_01430_));
 sg13g2_mux2_1 _18340_ (.A0(\spiking_network_top_uut.all_data_out[310] ),
    .A1(net4340),
    .S(_03285_),
    .X(_01431_));
 sg13g2_mux2_1 _18341_ (.A0(\spiking_network_top_uut.all_data_out[311] ),
    .A1(net4324),
    .S(_03285_),
    .X(_01432_));
 sg13g2_nor2_2 _18342_ (.A(_03215_),
    .B(net3731),
    .Y(_03286_));
 sg13g2_mux2_1 _18343_ (.A0(\spiking_network_top_uut.all_data_out[744] ),
    .A1(net4476),
    .S(_03286_),
    .X(_01433_));
 sg13g2_mux2_1 _18344_ (.A0(\spiking_network_top_uut.all_data_out[745] ),
    .A1(net4457),
    .S(_03286_),
    .X(_01434_));
 sg13g2_mux2_1 _18345_ (.A0(\spiking_network_top_uut.all_data_out[746] ),
    .A1(net4435),
    .S(_03286_),
    .X(_01435_));
 sg13g2_mux2_1 _18346_ (.A0(\spiking_network_top_uut.all_data_out[747] ),
    .A1(net4414),
    .S(_03286_),
    .X(_01436_));
 sg13g2_mux2_1 _18347_ (.A0(\spiking_network_top_uut.all_data_out[748] ),
    .A1(net4395),
    .S(_03286_),
    .X(_01437_));
 sg13g2_mux2_1 _18348_ (.A0(\spiking_network_top_uut.all_data_out[749] ),
    .A1(net4373),
    .S(_03286_),
    .X(_01438_));
 sg13g2_mux2_1 _18349_ (.A0(\spiking_network_top_uut.all_data_out[750] ),
    .A1(net4354),
    .S(_03286_),
    .X(_01439_));
 sg13g2_mux2_1 _18350_ (.A0(\spiking_network_top_uut.all_data_out[751] ),
    .A1(net4332),
    .S(_03286_),
    .X(_01440_));
 sg13g2_nor2_2 _18351_ (.A(_03225_),
    .B(net3729),
    .Y(_03287_));
 sg13g2_mux2_1 _18352_ (.A0(\spiking_network_top_uut.all_data_out[296] ),
    .A1(net4462),
    .S(_03287_),
    .X(_01441_));
 sg13g2_mux2_1 _18353_ (.A0(\spiking_network_top_uut.all_data_out[297] ),
    .A1(net4441),
    .S(_03287_),
    .X(_01442_));
 sg13g2_mux2_1 _18354_ (.A0(\spiking_network_top_uut.all_data_out[298] ),
    .A1(net4423),
    .S(_03287_),
    .X(_01443_));
 sg13g2_mux2_1 _18355_ (.A0(\spiking_network_top_uut.all_data_out[299] ),
    .A1(net4402),
    .S(_03287_),
    .X(_01444_));
 sg13g2_mux2_1 _18356_ (.A0(\spiking_network_top_uut.all_data_out[300] ),
    .A1(net4380),
    .S(_03287_),
    .X(_01445_));
 sg13g2_mux2_1 _18357_ (.A0(\spiking_network_top_uut.all_data_out[301] ),
    .A1(net4360),
    .S(_03287_),
    .X(_01446_));
 sg13g2_mux2_1 _18358_ (.A0(\spiking_network_top_uut.all_data_out[302] ),
    .A1(net4339),
    .S(_03287_),
    .X(_01447_));
 sg13g2_mux2_1 _18359_ (.A0(\spiking_network_top_uut.all_data_out[303] ),
    .A1(net4324),
    .S(_03287_),
    .X(_01448_));
 sg13g2_nor2_2 _18360_ (.A(_03211_),
    .B(_03245_),
    .Y(_03288_));
 sg13g2_mux2_1 _18361_ (.A0(\spiking_network_top_uut.all_data_out[520] ),
    .A1(net4477),
    .S(_03288_),
    .X(_01449_));
 sg13g2_mux2_1 _18362_ (.A0(\spiking_network_top_uut.all_data_out[521] ),
    .A1(net4460),
    .S(_03288_),
    .X(_01450_));
 sg13g2_mux2_1 _18363_ (.A0(\spiking_network_top_uut.all_data_out[522] ),
    .A1(net4436),
    .S(_03288_),
    .X(_01451_));
 sg13g2_mux2_1 _18364_ (.A0(\spiking_network_top_uut.all_data_out[523] ),
    .A1(net4417),
    .S(_03288_),
    .X(_01452_));
 sg13g2_mux2_1 _18365_ (.A0(\spiking_network_top_uut.all_data_out[524] ),
    .A1(net4396),
    .S(_03288_),
    .X(_01453_));
 sg13g2_mux2_1 _18366_ (.A0(\spiking_network_top_uut.all_data_out[525] ),
    .A1(net4375),
    .S(_03288_),
    .X(_01454_));
 sg13g2_mux2_1 _18367_ (.A0(\spiking_network_top_uut.all_data_out[526] ),
    .A1(net4355),
    .S(_03288_),
    .X(_01455_));
 sg13g2_mux2_1 _18368_ (.A0(\spiking_network_top_uut.all_data_out[527] ),
    .A1(net4335),
    .S(_03288_),
    .X(_01456_));
 sg13g2_nor2_2 _18369_ (.A(_03231_),
    .B(net3729),
    .Y(_03289_));
 sg13g2_mux2_1 _18370_ (.A0(\spiking_network_top_uut.all_data_out[288] ),
    .A1(net4462),
    .S(_03289_),
    .X(_01457_));
 sg13g2_mux2_1 _18371_ (.A0(\spiking_network_top_uut.all_data_out[289] ),
    .A1(net4442),
    .S(_03289_),
    .X(_01458_));
 sg13g2_mux2_1 _18372_ (.A0(\spiking_network_top_uut.all_data_out[290] ),
    .A1(net4423),
    .S(_03289_),
    .X(_01459_));
 sg13g2_mux2_1 _18373_ (.A0(\spiking_network_top_uut.all_data_out[291] ),
    .A1(net4401),
    .S(_03289_),
    .X(_01460_));
 sg13g2_mux2_1 _18374_ (.A0(\spiking_network_top_uut.all_data_out[292] ),
    .A1(net4381),
    .S(_03289_),
    .X(_01461_));
 sg13g2_mux2_1 _18375_ (.A0(\spiking_network_top_uut.all_data_out[293] ),
    .A1(net4360),
    .S(_03289_),
    .X(_01462_));
 sg13g2_mux2_1 _18376_ (.A0(\spiking_network_top_uut.all_data_out[294] ),
    .A1(net4340),
    .S(_03289_),
    .X(_01463_));
 sg13g2_mux2_1 _18377_ (.A0(\spiking_network_top_uut.all_data_out[295] ),
    .A1(net4319),
    .S(_03289_),
    .X(_01464_));
 sg13g2_nor2_2 _18378_ (.A(net3731),
    .B(_03258_),
    .Y(_03290_));
 sg13g2_mux2_1 _18379_ (.A0(\spiking_network_top_uut.all_data_out[752] ),
    .A1(net4474),
    .S(_03290_),
    .X(_01465_));
 sg13g2_mux2_1 _18380_ (.A0(\spiking_network_top_uut.all_data_out[753] ),
    .A1(net4452),
    .S(_03290_),
    .X(_01466_));
 sg13g2_mux2_1 _18381_ (.A0(\spiking_network_top_uut.all_data_out[754] ),
    .A1(net4433),
    .S(_03290_),
    .X(_01467_));
 sg13g2_mux2_1 _18382_ (.A0(\spiking_network_top_uut.all_data_out[755] ),
    .A1(net4416),
    .S(_03290_),
    .X(_01468_));
 sg13g2_mux2_1 _18383_ (.A0(\spiking_network_top_uut.all_data_out[756] ),
    .A1(net4392),
    .S(_03290_),
    .X(_01469_));
 sg13g2_mux2_1 _18384_ (.A0(\spiking_network_top_uut.all_data_out[757] ),
    .A1(net4372),
    .S(_03290_),
    .X(_01470_));
 sg13g2_mux2_1 _18385_ (.A0(\spiking_network_top_uut.all_data_out[758] ),
    .A1(net4351),
    .S(_03290_),
    .X(_01471_));
 sg13g2_mux2_1 _18386_ (.A0(\spiking_network_top_uut.all_data_out[759] ),
    .A1(net4334),
    .S(_03290_),
    .X(_01472_));
 sg13g2_nand2_2 _18387_ (.Y(_03291_),
    .A(_03234_),
    .B(_03254_));
 sg13g2_mux2_1 _18388_ (.A0(net4471),
    .A1(\spiking_network_top_uut.all_data_out[280] ),
    .S(_03291_),
    .X(_01473_));
 sg13g2_mux2_1 _18389_ (.A0(net4450),
    .A1(\spiking_network_top_uut.all_data_out[281] ),
    .S(_03291_),
    .X(_01474_));
 sg13g2_mux2_1 _18390_ (.A0(net4430),
    .A1(\spiking_network_top_uut.all_data_out[282] ),
    .S(_03291_),
    .X(_01475_));
 sg13g2_mux2_1 _18391_ (.A0(net4411),
    .A1(\spiking_network_top_uut.all_data_out[283] ),
    .S(_03291_),
    .X(_01476_));
 sg13g2_mux2_1 _18392_ (.A0(net4388),
    .A1(\spiking_network_top_uut.all_data_out[284] ),
    .S(_03291_),
    .X(_01477_));
 sg13g2_mux2_1 _18393_ (.A0(net4366),
    .A1(\spiking_network_top_uut.all_data_out[285] ),
    .S(_03291_),
    .X(_01478_));
 sg13g2_mux2_1 _18394_ (.A0(net4344),
    .A1(\spiking_network_top_uut.all_data_out[286] ),
    .S(_03291_),
    .X(_01479_));
 sg13g2_mux2_1 _18395_ (.A0(net4331),
    .A1(\spiking_network_top_uut.all_data_out[287] ),
    .S(_03291_),
    .X(_01480_));
 sg13g2_nor2_2 _18396_ (.A(net3734),
    .B(_03250_),
    .Y(_03292_));
 sg13g2_mux2_1 _18397_ (.A0(\spiking_network_top_uut.all_data_out[576] ),
    .A1(net4468),
    .S(_03292_),
    .X(_01481_));
 sg13g2_mux2_1 _18398_ (.A0(\spiking_network_top_uut.all_data_out[577] ),
    .A1(net4445),
    .S(_03292_),
    .X(_01482_));
 sg13g2_mux2_1 _18399_ (.A0(\spiking_network_top_uut.all_data_out[578] ),
    .A1(net4426),
    .S(_03292_),
    .X(_01483_));
 sg13g2_mux2_1 _18400_ (.A0(\spiking_network_top_uut.all_data_out[579] ),
    .A1(net4405),
    .S(_03292_),
    .X(_01484_));
 sg13g2_mux2_1 _18401_ (.A0(\spiking_network_top_uut.all_data_out[580] ),
    .A1(net4382),
    .S(_03292_),
    .X(_01485_));
 sg13g2_mux2_1 _18402_ (.A0(\spiking_network_top_uut.all_data_out[581] ),
    .A1(net4364),
    .S(_03292_),
    .X(_01486_));
 sg13g2_mux2_1 _18403_ (.A0(\spiking_network_top_uut.all_data_out[582] ),
    .A1(net4341),
    .S(_03292_),
    .X(_01487_));
 sg13g2_mux2_1 _18404_ (.A0(\spiking_network_top_uut.all_data_out[583] ),
    .A1(net4323),
    .S(_03292_),
    .X(_01488_));
 sg13g2_nand2_2 _18405_ (.Y(_03293_),
    .A(_03240_),
    .B(_03254_));
 sg13g2_mux2_1 _18406_ (.A0(net4462),
    .A1(\spiking_network_top_uut.all_data_out[272] ),
    .S(_03293_),
    .X(_01489_));
 sg13g2_mux2_1 _18407_ (.A0(net4441),
    .A1(\spiking_network_top_uut.all_data_out[273] ),
    .S(_03293_),
    .X(_01490_));
 sg13g2_mux2_1 _18408_ (.A0(net4423),
    .A1(\spiking_network_top_uut.all_data_out[274] ),
    .S(_03293_),
    .X(_01491_));
 sg13g2_mux2_1 _18409_ (.A0(net4404),
    .A1(\spiking_network_top_uut.all_data_out[275] ),
    .S(_03293_),
    .X(_01492_));
 sg13g2_mux2_1 _18410_ (.A0(net4386),
    .A1(\spiking_network_top_uut.all_data_out[276] ),
    .S(_03293_),
    .X(_01493_));
 sg13g2_mux2_1 _18411_ (.A0(net4369),
    .A1(\spiking_network_top_uut.all_data_out[277] ),
    .S(_03293_),
    .X(_01494_));
 sg13g2_mux2_1 _18412_ (.A0(net4347),
    .A1(\spiking_network_top_uut.all_data_out[278] ),
    .S(_03293_),
    .X(_01495_));
 sg13g2_mux2_1 _18413_ (.A0(net4328),
    .A1(\spiking_network_top_uut.all_data_out[279] ),
    .S(_03293_),
    .X(_01496_));
 sg13g2_nor2_2 _18414_ (.A(net3731),
    .B(_03256_),
    .Y(_03294_));
 sg13g2_mux2_1 _18415_ (.A0(\spiking_network_top_uut.all_data_out[760] ),
    .A1(net4467),
    .S(net3682),
    .X(_01497_));
 sg13g2_mux2_1 _18416_ (.A0(\spiking_network_top_uut.all_data_out[761] ),
    .A1(net4450),
    .S(_03294_),
    .X(_01498_));
 sg13g2_mux2_1 _18417_ (.A0(\spiking_network_top_uut.all_data_out[762] ),
    .A1(net4430),
    .S(net3682),
    .X(_01499_));
 sg13g2_mux2_1 _18418_ (.A0(\spiking_network_top_uut.all_data_out[763] ),
    .A1(net4408),
    .S(net3682),
    .X(_01500_));
 sg13g2_mux2_1 _18419_ (.A0(\spiking_network_top_uut.all_data_out[764] ),
    .A1(net4388),
    .S(net3682),
    .X(_01501_));
 sg13g2_mux2_1 _18420_ (.A0(\spiking_network_top_uut.all_data_out[765] ),
    .A1(net4366),
    .S(net3682),
    .X(_01502_));
 sg13g2_nand2_1 _18421_ (.Y(_03295_),
    .A(net4347),
    .B(net3682));
 sg13g2_o21ai_1 _18422_ (.B1(_03295_),
    .Y(_01503_),
    .A1(_03515_),
    .A2(net3682));
 sg13g2_mux2_1 _18423_ (.A0(\spiking_network_top_uut.all_data_out[767] ),
    .A1(net4326),
    .S(net3682),
    .X(_01504_));
 sg13g2_nand2_2 _18424_ (.Y(_03296_),
    .A(_03244_),
    .B(_03254_));
 sg13g2_mux2_1 _18425_ (.A0(net4471),
    .A1(\spiking_network_top_uut.all_data_out[264] ),
    .S(_03296_),
    .X(_01505_));
 sg13g2_mux2_1 _18426_ (.A0(net4450),
    .A1(\spiking_network_top_uut.all_data_out[265] ),
    .S(_03296_),
    .X(_01506_));
 sg13g2_mux2_1 _18427_ (.A0(net4430),
    .A1(\spiking_network_top_uut.all_data_out[266] ),
    .S(_03296_),
    .X(_01507_));
 sg13g2_mux2_1 _18428_ (.A0(net4409),
    .A1(\spiking_network_top_uut.all_data_out[267] ),
    .S(_03296_),
    .X(_01508_));
 sg13g2_mux2_1 _18429_ (.A0(net4386),
    .A1(\spiking_network_top_uut.all_data_out[268] ),
    .S(_03296_),
    .X(_01509_));
 sg13g2_mux2_1 _18430_ (.A0(net4369),
    .A1(\spiking_network_top_uut.all_data_out[269] ),
    .S(_03296_),
    .X(_01510_));
 sg13g2_mux2_1 _18431_ (.A0(net4344),
    .A1(\spiking_network_top_uut.all_data_out[270] ),
    .S(_03296_),
    .X(_01511_));
 sg13g2_mux2_1 _18432_ (.A0(net4325),
    .A1(\spiking_network_top_uut.all_data_out[271] ),
    .S(_03296_),
    .X(_01512_));
 sg13g2_nor2_2 _18433_ (.A(_03201_),
    .B(net3734),
    .Y(_03297_));
 sg13g2_mux2_1 _18434_ (.A0(\spiking_network_top_uut.all_data_out[512] ),
    .A1(net4478),
    .S(_03297_),
    .X(_01513_));
 sg13g2_mux2_1 _18435_ (.A0(\spiking_network_top_uut.all_data_out[513] ),
    .A1(net4455),
    .S(_03297_),
    .X(_01514_));
 sg13g2_mux2_1 _18436_ (.A0(\spiking_network_top_uut.all_data_out[514] ),
    .A1(net4434),
    .S(_03297_),
    .X(_01515_));
 sg13g2_mux2_1 _18437_ (.A0(\spiking_network_top_uut.all_data_out[515] ),
    .A1(net4410),
    .S(_03297_),
    .X(_01516_));
 sg13g2_mux2_1 _18438_ (.A0(\spiking_network_top_uut.all_data_out[516] ),
    .A1(net4397),
    .S(_03297_),
    .X(_01517_));
 sg13g2_mux2_1 _18439_ (.A0(\spiking_network_top_uut.all_data_out[517] ),
    .A1(net4376),
    .S(_03297_),
    .X(_01518_));
 sg13g2_mux2_1 _18440_ (.A0(\spiking_network_top_uut.all_data_out[518] ),
    .A1(net4357),
    .S(_03297_),
    .X(_01519_));
 sg13g2_mux2_1 _18441_ (.A0(\spiking_network_top_uut.all_data_out[519] ),
    .A1(net4334),
    .S(_03297_),
    .X(_01520_));
 sg13g2_nand3_1 _18442_ (.B(_03200_),
    .C(_03254_),
    .A(net3737),
    .Y(_03298_));
 sg13g2_mux2_1 _18443_ (.A0(net4464),
    .A1(\spiking_network_top_uut.all_data_out[256] ),
    .S(_03298_),
    .X(_01521_));
 sg13g2_mux2_1 _18444_ (.A0(net4443),
    .A1(\spiking_network_top_uut.all_data_out[257] ),
    .S(_03298_),
    .X(_01522_));
 sg13g2_mux2_1 _18445_ (.A0(net4424),
    .A1(\spiking_network_top_uut.all_data_out[258] ),
    .S(_03298_),
    .X(_01523_));
 sg13g2_mux2_1 _18446_ (.A0(net4403),
    .A1(\spiking_network_top_uut.all_data_out[259] ),
    .S(_03298_),
    .X(_01524_));
 sg13g2_mux2_1 _18447_ (.A0(net4388),
    .A1(\spiking_network_top_uut.all_data_out[260] ),
    .S(_03298_),
    .X(_01525_));
 sg13g2_mux2_1 _18448_ (.A0(net4366),
    .A1(\spiking_network_top_uut.all_data_out[261] ),
    .S(_03298_),
    .X(_01526_));
 sg13g2_mux2_1 _18449_ (.A0(net4347),
    .A1(\spiking_network_top_uut.all_data_out[262] ),
    .S(_03298_),
    .X(_01527_));
 sg13g2_mux2_1 _18450_ (.A0(net4325),
    .A1(\spiking_network_top_uut.all_data_out[263] ),
    .S(_03298_),
    .X(_01528_));
 sg13g2_nor2_2 _18451_ (.A(_00027_),
    .B(_03253_),
    .Y(_03299_));
 sg13g2_nand2b_1 _18452_ (.Y(_03300_),
    .B(_03252_),
    .A_N(_00027_));
 sg13g2_nand3_1 _18453_ (.B(_03200_),
    .C(_03299_),
    .A(net3737),
    .Y(_03301_));
 sg13g2_mux2_1 _18454_ (.A0(net4464),
    .A1(\spiking_network_top_uut.all_data_out[768] ),
    .S(_03301_),
    .X(_01529_));
 sg13g2_mux2_1 _18455_ (.A0(net4445),
    .A1(\spiking_network_top_uut.all_data_out[769] ),
    .S(net3698),
    .X(_01530_));
 sg13g2_mux2_1 _18456_ (.A0(net4427),
    .A1(\spiking_network_top_uut.all_data_out[770] ),
    .S(net3698),
    .X(_01531_));
 sg13g2_mux2_1 _18457_ (.A0(net4403),
    .A1(\spiking_network_top_uut.all_data_out[771] ),
    .S(net3698),
    .X(_01532_));
 sg13g2_mux2_1 _18458_ (.A0(net4387),
    .A1(\spiking_network_top_uut.all_data_out[772] ),
    .S(net3698),
    .X(_01533_));
 sg13g2_mux2_1 _18459_ (.A0(net4362),
    .A1(\spiking_network_top_uut.all_data_out[773] ),
    .S(net3698),
    .X(_01534_));
 sg13g2_nor2_1 _18460_ (.A(net4339),
    .B(net3698),
    .Y(_03302_));
 sg13g2_a21oi_1 _18461_ (.A1(_03513_),
    .A2(net3698),
    .Y(_01535_),
    .B1(_03302_));
 sg13g2_mux2_1 _18462_ (.A0(net4320),
    .A1(\spiking_network_top_uut.all_data_out[775] ),
    .S(net3698),
    .X(_01536_));
 sg13g2_nor2_2 _18463_ (.A(\spiking_network_top_uut.spi_inst.LSB_Address_reg[6] ),
    .B(_03222_),
    .Y(_03303_));
 sg13g2_nand2b_1 _18464_ (.Y(_03304_),
    .B(_03221_),
    .A_N(\spiking_network_top_uut.spi_inst.LSB_Address_reg[6] ));
 sg13g2_nor2_2 _18465_ (.A(net15),
    .B(net3725),
    .Y(_03305_));
 sg13g2_mux2_1 _18466_ (.A0(\spiking_network_top_uut.all_data_out[248] ),
    .A1(net4469),
    .S(_03305_),
    .X(_01537_));
 sg13g2_mux2_1 _18467_ (.A0(\spiking_network_top_uut.all_data_out[249] ),
    .A1(net4447),
    .S(_03305_),
    .X(_01538_));
 sg13g2_mux2_1 _18468_ (.A0(\spiking_network_top_uut.all_data_out[250] ),
    .A1(net4428),
    .S(_03305_),
    .X(_01539_));
 sg13g2_mux2_1 _18469_ (.A0(\spiking_network_top_uut.all_data_out[251] ),
    .A1(net4406),
    .S(_03305_),
    .X(_01540_));
 sg13g2_mux2_1 _18470_ (.A0(\spiking_network_top_uut.all_data_out[252] ),
    .A1(net4382),
    .S(_03305_),
    .X(_01541_));
 sg13g2_mux2_1 _18471_ (.A0(\spiking_network_top_uut.all_data_out[253] ),
    .A1(net4364),
    .S(_03305_),
    .X(_01542_));
 sg13g2_mux2_1 _18472_ (.A0(\spiking_network_top_uut.all_data_out[254] ),
    .A1(net4341),
    .S(_03305_),
    .X(_01543_));
 sg13g2_mux2_1 _18473_ (.A0(\spiking_network_top_uut.all_data_out[255] ),
    .A1(net4323),
    .S(_03305_),
    .X(_01544_));
 sg13g2_nand3_1 _18474_ (.B(_03200_),
    .C(_03223_),
    .A(net3737),
    .Y(_03306_));
 sg13g2_mux2_1 _18475_ (.A0(net4468),
    .A1(\spiking_network_top_uut.all_data_out[640] ),
    .S(net3697),
    .X(_01545_));
 sg13g2_mux2_1 _18476_ (.A0(net4445),
    .A1(\spiking_network_top_uut.all_data_out[641] ),
    .S(_03306_),
    .X(_01546_));
 sg13g2_mux2_1 _18477_ (.A0(net4424),
    .A1(\spiking_network_top_uut.all_data_out[642] ),
    .S(net3697),
    .X(_01547_));
 sg13g2_mux2_1 _18478_ (.A0(net4401),
    .A1(\spiking_network_top_uut.all_data_out[643] ),
    .S(net3697),
    .X(_01548_));
 sg13g2_mux2_1 _18479_ (.A0(net4380),
    .A1(\spiking_network_top_uut.all_data_out[644] ),
    .S(net3697),
    .X(_01549_));
 sg13g2_mux2_1 _18480_ (.A0(net4362),
    .A1(\spiking_network_top_uut.all_data_out[645] ),
    .S(net3697),
    .X(_01550_));
 sg13g2_nor2_1 _18481_ (.A(net4346),
    .B(net3697),
    .Y(_03307_));
 sg13g2_a21oi_1 _18482_ (.A1(_03528_),
    .A2(net3697),
    .Y(_01551_),
    .B1(_03307_));
 sg13g2_mux2_1 _18483_ (.A0(net4319),
    .A1(\spiking_network_top_uut.all_data_out[647] ),
    .S(net3697),
    .X(_01552_));
 sg13g2_nor2_2 _18484_ (.A(_03258_),
    .B(net3725),
    .Y(_03308_));
 sg13g2_mux2_1 _18485_ (.A0(\spiking_network_top_uut.all_data_out[240] ),
    .A1(net4466),
    .S(_03308_),
    .X(_01553_));
 sg13g2_mux2_1 _18486_ (.A0(\spiking_network_top_uut.all_data_out[241] ),
    .A1(net4449),
    .S(_03308_),
    .X(_01554_));
 sg13g2_mux2_1 _18487_ (.A0(\spiking_network_top_uut.all_data_out[242] ),
    .A1(net4425),
    .S(_03308_),
    .X(_01555_));
 sg13g2_mux2_1 _18488_ (.A0(\spiking_network_top_uut.all_data_out[243] ),
    .A1(net4404),
    .S(_03308_),
    .X(_01556_));
 sg13g2_mux2_1 _18489_ (.A0(\spiking_network_top_uut.all_data_out[244] ),
    .A1(net4383),
    .S(_03308_),
    .X(_01557_));
 sg13g2_mux2_1 _18490_ (.A0(\spiking_network_top_uut.all_data_out[245] ),
    .A1(net4364),
    .S(_03308_),
    .X(_01558_));
 sg13g2_mux2_1 _18491_ (.A0(\spiking_network_top_uut.all_data_out[246] ),
    .A1(net4345),
    .S(_03308_),
    .X(_01559_));
 sg13g2_mux2_1 _18492_ (.A0(\spiking_network_top_uut.all_data_out[247] ),
    .A1(net4322),
    .S(_03308_),
    .X(_01560_));
 sg13g2_nand2_2 _18493_ (.Y(_03309_),
    .A(_03244_),
    .B(_03299_));
 sg13g2_mux2_1 _18494_ (.A0(net4476),
    .A1(\spiking_network_top_uut.all_data_out[776] ),
    .S(_03309_),
    .X(_01561_));
 sg13g2_mux2_1 _18495_ (.A0(net4456),
    .A1(\spiking_network_top_uut.all_data_out[777] ),
    .S(_03309_),
    .X(_01562_));
 sg13g2_mux2_1 _18496_ (.A0(net4435),
    .A1(\spiking_network_top_uut.all_data_out[778] ),
    .S(_03309_),
    .X(_01563_));
 sg13g2_mux2_1 _18497_ (.A0(net4413),
    .A1(\spiking_network_top_uut.all_data_out[779] ),
    .S(_03309_),
    .X(_01564_));
 sg13g2_mux2_1 _18498_ (.A0(net4394),
    .A1(\spiking_network_top_uut.all_data_out[780] ),
    .S(_03309_),
    .X(_01565_));
 sg13g2_mux2_1 _18499_ (.A0(net4378),
    .A1(\spiking_network_top_uut.all_data_out[781] ),
    .S(_03309_),
    .X(_01566_));
 sg13g2_mux2_1 _18500_ (.A0(net4353),
    .A1(\spiking_network_top_uut.all_data_out[782] ),
    .S(_03309_),
    .X(_01567_));
 sg13g2_mux2_1 _18501_ (.A0(net4334),
    .A1(\spiking_network_top_uut.all_data_out[783] ),
    .S(_03309_),
    .X(_01568_));
 sg13g2_nor2_2 _18502_ (.A(_03215_),
    .B(net3725),
    .Y(_03310_));
 sg13g2_mux2_1 _18503_ (.A0(\spiking_network_top_uut.all_data_out[232] ),
    .A1(net4466),
    .S(_03310_),
    .X(_01569_));
 sg13g2_mux2_1 _18504_ (.A0(\spiking_network_top_uut.all_data_out[233] ),
    .A1(net4444),
    .S(_03310_),
    .X(_01570_));
 sg13g2_mux2_1 _18505_ (.A0(\spiking_network_top_uut.all_data_out[234] ),
    .A1(net4428),
    .S(_03310_),
    .X(_01571_));
 sg13g2_mux2_1 _18506_ (.A0(\spiking_network_top_uut.all_data_out[235] ),
    .A1(net4406),
    .S(_03310_),
    .X(_01572_));
 sg13g2_mux2_1 _18507_ (.A0(\spiking_network_top_uut.all_data_out[236] ),
    .A1(net4382),
    .S(_03310_),
    .X(_01573_));
 sg13g2_mux2_1 _18508_ (.A0(\spiking_network_top_uut.all_data_out[237] ),
    .A1(net4365),
    .S(_03310_),
    .X(_01574_));
 sg13g2_mux2_1 _18509_ (.A0(\spiking_network_top_uut.all_data_out[238] ),
    .A1(net4341),
    .S(_03310_),
    .X(_01575_));
 sg13g2_mux2_1 _18510_ (.A0(\spiking_network_top_uut.all_data_out[239] ),
    .A1(net4321),
    .S(_03310_),
    .X(_01576_));
 sg13g2_nor2_2 _18511_ (.A(net3735),
    .B(net15),
    .Y(_03311_));
 sg13g2_mux2_1 _18512_ (.A0(\spiking_network_top_uut.all_data_out[504] ),
    .A1(net4479),
    .S(_03311_),
    .X(_01577_));
 sg13g2_mux2_1 _18513_ (.A0(\spiking_network_top_uut.all_data_out[505] ),
    .A1(net4459),
    .S(_03311_),
    .X(_01578_));
 sg13g2_mux2_1 _18514_ (.A0(\spiking_network_top_uut.all_data_out[506] ),
    .A1(net4438),
    .S(_03311_),
    .X(_01579_));
 sg13g2_mux2_1 _18515_ (.A0(\spiking_network_top_uut.all_data_out[507] ),
    .A1(net4414),
    .S(_03311_),
    .X(_01580_));
 sg13g2_mux2_1 _18516_ (.A0(\spiking_network_top_uut.all_data_out[508] ),
    .A1(net4397),
    .S(_03311_),
    .X(_01581_));
 sg13g2_mux2_1 _18517_ (.A0(\spiking_network_top_uut.all_data_out[509] ),
    .A1(net4376),
    .S(_03311_),
    .X(_01582_));
 sg13g2_mux2_1 _18518_ (.A0(\spiking_network_top_uut.all_data_out[510] ),
    .A1(net4356),
    .S(_03311_),
    .X(_01583_));
 sg13g2_mux2_1 _18519_ (.A0(\spiking_network_top_uut.all_data_out[511] ),
    .A1(net4330),
    .S(_03311_),
    .X(_01584_));
 sg13g2_nor2_2 _18520_ (.A(_03268_),
    .B(net3725),
    .Y(_03312_));
 sg13g2_mux2_1 _18521_ (.A0(\spiking_network_top_uut.all_data_out[224] ),
    .A1(net4466),
    .S(_03312_),
    .X(_01585_));
 sg13g2_mux2_1 _18522_ (.A0(\spiking_network_top_uut.all_data_out[225] ),
    .A1(net4444),
    .S(_03312_),
    .X(_01586_));
 sg13g2_mux2_1 _18523_ (.A0(\spiking_network_top_uut.all_data_out[226] ),
    .A1(net4425),
    .S(_03312_),
    .X(_01587_));
 sg13g2_mux2_1 _18524_ (.A0(\spiking_network_top_uut.all_data_out[227] ),
    .A1(net4406),
    .S(_03312_),
    .X(_01588_));
 sg13g2_mux2_1 _18525_ (.A0(\spiking_network_top_uut.all_data_out[228] ),
    .A1(net4385),
    .S(_03312_),
    .X(_01589_));
 sg13g2_mux2_1 _18526_ (.A0(\spiking_network_top_uut.all_data_out[229] ),
    .A1(net4367),
    .S(_03312_),
    .X(_01590_));
 sg13g2_mux2_1 _18527_ (.A0(\spiking_network_top_uut.all_data_out[230] ),
    .A1(net4344),
    .S(_03312_),
    .X(_01591_));
 sg13g2_mux2_1 _18528_ (.A0(\spiking_network_top_uut.all_data_out[231] ),
    .A1(net4326),
    .S(_03312_),
    .X(_01592_));
 sg13g2_nand2_2 _18529_ (.Y(_03313_),
    .A(_03240_),
    .B(_03299_));
 sg13g2_mux2_1 _18530_ (.A0(net4473),
    .A1(\spiking_network_top_uut.all_data_out[784] ),
    .S(_03313_),
    .X(_01593_));
 sg13g2_mux2_1 _18531_ (.A0(net4452),
    .A1(\spiking_network_top_uut.all_data_out[785] ),
    .S(_03313_),
    .X(_01594_));
 sg13g2_mux2_1 _18532_ (.A0(net4432),
    .A1(\spiking_network_top_uut.all_data_out[786] ),
    .S(_03313_),
    .X(_01595_));
 sg13g2_mux2_1 _18533_ (.A0(net4413),
    .A1(\spiking_network_top_uut.all_data_out[787] ),
    .S(_03313_),
    .X(_01596_));
 sg13g2_mux2_1 _18534_ (.A0(net4392),
    .A1(\spiking_network_top_uut.all_data_out[788] ),
    .S(_03313_),
    .X(_01597_));
 sg13g2_mux2_1 _18535_ (.A0(net4372),
    .A1(\spiking_network_top_uut.all_data_out[789] ),
    .S(_03313_),
    .X(_01598_));
 sg13g2_mux2_1 _18536_ (.A0(net4351),
    .A1(\spiking_network_top_uut.all_data_out[790] ),
    .S(_03313_),
    .X(_01599_));
 sg13g2_mux2_1 _18537_ (.A0(net4334),
    .A1(\spiking_network_top_uut.all_data_out[791] ),
    .S(_03313_),
    .X(_01600_));
 sg13g2_nor2_2 _18538_ (.A(net14),
    .B(net3726),
    .Y(_03314_));
 sg13g2_mux2_1 _18539_ (.A0(\spiking_network_top_uut.all_data_out[216] ),
    .A1(net4471),
    .S(_03314_),
    .X(_01601_));
 sg13g2_mux2_1 _18540_ (.A0(\spiking_network_top_uut.all_data_out[217] ),
    .A1(net4450),
    .S(_03314_),
    .X(_01602_));
 sg13g2_mux2_1 _18541_ (.A0(\spiking_network_top_uut.all_data_out[218] ),
    .A1(net4430),
    .S(_03314_),
    .X(_01603_));
 sg13g2_mux2_1 _18542_ (.A0(\spiking_network_top_uut.all_data_out[219] ),
    .A1(net4411),
    .S(_03314_),
    .X(_01604_));
 sg13g2_mux2_1 _18543_ (.A0(\spiking_network_top_uut.all_data_out[220] ),
    .A1(net4389),
    .S(_03314_),
    .X(_01605_));
 sg13g2_mux2_1 _18544_ (.A0(\spiking_network_top_uut.all_data_out[221] ),
    .A1(net4369),
    .S(_03314_),
    .X(_01606_));
 sg13g2_mux2_1 _18545_ (.A0(\spiking_network_top_uut.all_data_out[222] ),
    .A1(net4348),
    .S(_03314_),
    .X(_01607_));
 sg13g2_mux2_1 _18546_ (.A0(\spiking_network_top_uut.all_data_out[223] ),
    .A1(net4331),
    .S(_03314_),
    .X(_01608_));
 sg13g2_nor2_1 _18547_ (.A(net3734),
    .B(_03268_),
    .Y(_03315_));
 sg13g2_mux2_1 _18548_ (.A0(\spiking_network_top_uut.all_data_out[608] ),
    .A1(net4468),
    .S(net3681),
    .X(_01609_));
 sg13g2_mux2_1 _18549_ (.A0(\spiking_network_top_uut.all_data_out[609] ),
    .A1(net4445),
    .S(_03315_),
    .X(_01610_));
 sg13g2_mux2_1 _18550_ (.A0(\spiking_network_top_uut.all_data_out[610] ),
    .A1(net4426),
    .S(net3681),
    .X(_01611_));
 sg13g2_mux2_1 _18551_ (.A0(\spiking_network_top_uut.all_data_out[611] ),
    .A1(net4405),
    .S(net3681),
    .X(_01612_));
 sg13g2_mux2_1 _18552_ (.A0(\spiking_network_top_uut.all_data_out[612] ),
    .A1(net4382),
    .S(net3681),
    .X(_01613_));
 sg13g2_mux2_1 _18553_ (.A0(\spiking_network_top_uut.all_data_out[613] ),
    .A1(net4362),
    .S(net3681),
    .X(_01614_));
 sg13g2_nand2_1 _18554_ (.Y(_03316_),
    .A(net4341),
    .B(net3681));
 sg13g2_o21ai_1 _18555_ (.B1(_03316_),
    .Y(_01615_),
    .A1(_03531_),
    .A2(net3681));
 sg13g2_mux2_1 _18556_ (.A0(\spiking_network_top_uut.all_data_out[615] ),
    .A1(net4322),
    .S(net3681),
    .X(_01616_));
 sg13g2_nor2_2 _18557_ (.A(_03270_),
    .B(net3725),
    .Y(_03317_));
 sg13g2_mux2_1 _18558_ (.A0(\spiking_network_top_uut.all_data_out[208] ),
    .A1(net4464),
    .S(_03317_),
    .X(_01617_));
 sg13g2_mux2_1 _18559_ (.A0(\spiking_network_top_uut.all_data_out[209] ),
    .A1(net4445),
    .S(_03317_),
    .X(_01618_));
 sg13g2_mux2_1 _18560_ (.A0(\spiking_network_top_uut.all_data_out[210] ),
    .A1(net4426),
    .S(_03317_),
    .X(_01619_));
 sg13g2_mux2_1 _18561_ (.A0(\spiking_network_top_uut.all_data_out[211] ),
    .A1(net4405),
    .S(_03317_),
    .X(_01620_));
 sg13g2_mux2_1 _18562_ (.A0(\spiking_network_top_uut.all_data_out[212] ),
    .A1(net4388),
    .S(_03317_),
    .X(_01621_));
 sg13g2_mux2_1 _18563_ (.A0(\spiking_network_top_uut.all_data_out[213] ),
    .A1(net4369),
    .S(_03317_),
    .X(_01622_));
 sg13g2_mux2_1 _18564_ (.A0(\spiking_network_top_uut.all_data_out[214] ),
    .A1(net4349),
    .S(_03317_),
    .X(_01623_));
 sg13g2_mux2_1 _18565_ (.A0(\spiking_network_top_uut.all_data_out[215] ),
    .A1(net4331),
    .S(_03317_),
    .X(_01624_));
 sg13g2_nand2_2 _18566_ (.Y(_03318_),
    .A(_03234_),
    .B(_03299_));
 sg13g2_mux2_1 _18567_ (.A0(net4471),
    .A1(\spiking_network_top_uut.all_data_out[792] ),
    .S(_03318_),
    .X(_01625_));
 sg13g2_mux2_1 _18568_ (.A0(net4450),
    .A1(\spiking_network_top_uut.all_data_out[793] ),
    .S(_03318_),
    .X(_01626_));
 sg13g2_mux2_1 _18569_ (.A0(net4430),
    .A1(\spiking_network_top_uut.all_data_out[794] ),
    .S(_03318_),
    .X(_01627_));
 sg13g2_mux2_1 _18570_ (.A0(net4411),
    .A1(\spiking_network_top_uut.all_data_out[795] ),
    .S(_03318_),
    .X(_01628_));
 sg13g2_mux2_1 _18571_ (.A0(net4389),
    .A1(\spiking_network_top_uut.all_data_out[796] ),
    .S(_03318_),
    .X(_01629_));
 sg13g2_mux2_1 _18572_ (.A0(net4370),
    .A1(\spiking_network_top_uut.all_data_out[797] ),
    .S(_03318_),
    .X(_01630_));
 sg13g2_mux2_1 _18573_ (.A0(net4348),
    .A1(\spiking_network_top_uut.all_data_out[798] ),
    .S(_03318_),
    .X(_01631_));
 sg13g2_mux2_1 _18574_ (.A0(net4328),
    .A1(\spiking_network_top_uut.all_data_out[799] ),
    .S(_03318_),
    .X(_01632_));
 sg13g2_nor2_2 _18575_ (.A(_03238_),
    .B(net3725),
    .Y(_03319_));
 sg13g2_mux2_1 _18576_ (.A0(\spiking_network_top_uut.all_data_out[200] ),
    .A1(net4470),
    .S(_03319_),
    .X(_01633_));
 sg13g2_mux2_1 _18577_ (.A0(\spiking_network_top_uut.all_data_out[201] ),
    .A1(net4444),
    .S(_03319_),
    .X(_01634_));
 sg13g2_mux2_1 _18578_ (.A0(\spiking_network_top_uut.all_data_out[202] ),
    .A1(net4424),
    .S(_03319_),
    .X(_01635_));
 sg13g2_mux2_1 _18579_ (.A0(\spiking_network_top_uut.all_data_out[203] ),
    .A1(net4404),
    .S(_03319_),
    .X(_01636_));
 sg13g2_mux2_1 _18580_ (.A0(\spiking_network_top_uut.all_data_out[204] ),
    .A1(net4387),
    .S(_03319_),
    .X(_01637_));
 sg13g2_mux2_1 _18581_ (.A0(\spiking_network_top_uut.all_data_out[205] ),
    .A1(net4361),
    .S(_03319_),
    .X(_01638_));
 sg13g2_mux2_1 _18582_ (.A0(\spiking_network_top_uut.all_data_out[206] ),
    .A1(net4339),
    .S(_03319_),
    .X(_01639_));
 sg13g2_mux2_1 _18583_ (.A0(\spiking_network_top_uut.all_data_out[207] ),
    .A1(net4320),
    .S(_03319_),
    .X(_01640_));
 sg13g2_nor2_2 _18584_ (.A(net3735),
    .B(_03258_),
    .Y(_03320_));
 sg13g2_mux2_1 _18585_ (.A0(\spiking_network_top_uut.all_data_out[496] ),
    .A1(net4474),
    .S(_03320_),
    .X(_01641_));
 sg13g2_mux2_1 _18586_ (.A0(\spiking_network_top_uut.all_data_out[497] ),
    .A1(net4453),
    .S(_03320_),
    .X(_01642_));
 sg13g2_mux2_1 _18587_ (.A0(\spiking_network_top_uut.all_data_out[498] ),
    .A1(net4433),
    .S(_03320_),
    .X(_01643_));
 sg13g2_mux2_1 _18588_ (.A0(\spiking_network_top_uut.all_data_out[499] ),
    .A1(net4415),
    .S(_03320_),
    .X(_01644_));
 sg13g2_mux2_1 _18589_ (.A0(\spiking_network_top_uut.all_data_out[500] ),
    .A1(net4393),
    .S(_03320_),
    .X(_01645_));
 sg13g2_mux2_1 _18590_ (.A0(\spiking_network_top_uut.all_data_out[501] ),
    .A1(net4370),
    .S(_03320_),
    .X(_01646_));
 sg13g2_mux2_1 _18591_ (.A0(\spiking_network_top_uut.all_data_out[502] ),
    .A1(net4352),
    .S(_03320_),
    .X(_01647_));
 sg13g2_mux2_1 _18592_ (.A0(\spiking_network_top_uut.all_data_out[503] ),
    .A1(net4332),
    .S(_03320_),
    .X(_01648_));
 sg13g2_nor2_2 _18593_ (.A(_03250_),
    .B(net3725),
    .Y(_03321_));
 sg13g2_mux2_1 _18594_ (.A0(\spiking_network_top_uut.all_data_out[192] ),
    .A1(net4462),
    .S(_03321_),
    .X(_01649_));
 sg13g2_mux2_1 _18595_ (.A0(\spiking_network_top_uut.all_data_out[193] ),
    .A1(net4441),
    .S(_03321_),
    .X(_01650_));
 sg13g2_mux2_1 _18596_ (.A0(\spiking_network_top_uut.all_data_out[194] ),
    .A1(net4422),
    .S(_03321_),
    .X(_01651_));
 sg13g2_mux2_1 _18597_ (.A0(\spiking_network_top_uut.all_data_out[195] ),
    .A1(net4401),
    .S(_03321_),
    .X(_01652_));
 sg13g2_mux2_1 _18598_ (.A0(\spiking_network_top_uut.all_data_out[196] ),
    .A1(net4380),
    .S(_03321_),
    .X(_01653_));
 sg13g2_mux2_1 _18599_ (.A0(\spiking_network_top_uut.all_data_out[197] ),
    .A1(net4361),
    .S(_03321_),
    .X(_01654_));
 sg13g2_mux2_1 _18600_ (.A0(\spiking_network_top_uut.all_data_out[198] ),
    .A1(net4339),
    .S(_03321_),
    .X(_01655_));
 sg13g2_mux2_1 _18601_ (.A0(\spiking_network_top_uut.all_data_out[199] ),
    .A1(net4320),
    .S(_03321_),
    .X(_01656_));
 sg13g2_nor2_2 _18602_ (.A(_03231_),
    .B(net3728),
    .Y(_03322_));
 sg13g2_mux2_1 _18603_ (.A0(\spiking_network_top_uut.all_data_out[800] ),
    .A1(net4468),
    .S(net3680),
    .X(_01657_));
 sg13g2_mux2_1 _18604_ (.A0(\spiking_network_top_uut.all_data_out[801] ),
    .A1(net4445),
    .S(_03322_),
    .X(_01658_));
 sg13g2_nand2_1 _18605_ (.Y(_03323_),
    .A(net4426),
    .B(net3680));
 sg13g2_o21ai_1 _18606_ (.B1(_03323_),
    .Y(_01659_),
    .A1(_03585_),
    .A2(net3680));
 sg13g2_mux2_1 _18607_ (.A0(\spiking_network_top_uut.all_data_out[803] ),
    .A1(net4402),
    .S(net3680),
    .X(_01660_));
 sg13g2_mux2_1 _18608_ (.A0(\spiking_network_top_uut.all_data_out[804] ),
    .A1(net4387),
    .S(net3680),
    .X(_01661_));
 sg13g2_mux2_1 _18609_ (.A0(\spiking_network_top_uut.all_data_out[805] ),
    .A1(net4362),
    .S(net3680),
    .X(_01662_));
 sg13g2_mux2_1 _18610_ (.A0(\spiking_network_top_uut.all_data_out[806] ),
    .A1(net4339),
    .S(net3680),
    .X(_01663_));
 sg13g2_mux2_1 _18611_ (.A0(\spiking_network_top_uut.all_data_out[807] ),
    .A1(net4319),
    .S(net3680),
    .X(_01664_));
 sg13g2_nor2_2 _18612_ (.A(_03208_),
    .B(net3726),
    .Y(_03324_));
 sg13g2_mux2_1 _18613_ (.A0(\spiking_network_top_uut.all_data_out[184] ),
    .A1(net4467),
    .S(_03324_),
    .X(_01665_));
 sg13g2_mux2_1 _18614_ (.A0(\spiking_network_top_uut.all_data_out[185] ),
    .A1(net4446),
    .S(_03324_),
    .X(_01666_));
 sg13g2_mux2_1 _18615_ (.A0(\spiking_network_top_uut.all_data_out[186] ),
    .A1(net4427),
    .S(_03324_),
    .X(_01667_));
 sg13g2_mux2_1 _18616_ (.A0(\spiking_network_top_uut.all_data_out[187] ),
    .A1(net4409),
    .S(_03324_),
    .X(_01668_));
 sg13g2_mux2_1 _18617_ (.A0(\spiking_network_top_uut.all_data_out[188] ),
    .A1(net4386),
    .S(_03324_),
    .X(_01669_));
 sg13g2_mux2_1 _18618_ (.A0(\spiking_network_top_uut.all_data_out[189] ),
    .A1(net4366),
    .S(_03324_),
    .X(_01670_));
 sg13g2_mux2_1 _18619_ (.A0(\spiking_network_top_uut.all_data_out[190] ),
    .A1(net4343),
    .S(_03324_),
    .X(_01671_));
 sg13g2_mux2_1 _18620_ (.A0(\spiking_network_top_uut.all_data_out[191] ),
    .A1(net4326),
    .S(_03324_),
    .X(_01672_));
 sg13g2_nand2_2 _18621_ (.Y(_03325_),
    .A(_03223_),
    .B(_03244_));
 sg13g2_mux2_1 _18622_ (.A0(net4476),
    .A1(\spiking_network_top_uut.all_data_out[648] ),
    .S(_03325_),
    .X(_01673_));
 sg13g2_mux2_1 _18623_ (.A0(net4456),
    .A1(\spiking_network_top_uut.all_data_out[649] ),
    .S(net3679),
    .X(_01674_));
 sg13g2_nor2_1 _18624_ (.A(net4435),
    .B(net3679),
    .Y(_03326_));
 sg13g2_a21oi_1 _18625_ (.A1(_03600_),
    .A2(net3679),
    .Y(_01675_),
    .B1(_03326_));
 sg13g2_mux2_1 _18626_ (.A0(net4417),
    .A1(\spiking_network_top_uut.all_data_out[651] ),
    .S(net3679),
    .X(_01676_));
 sg13g2_mux2_1 _18627_ (.A0(net4395),
    .A1(\spiking_network_top_uut.all_data_out[652] ),
    .S(net3679),
    .X(_01677_));
 sg13g2_mux2_1 _18628_ (.A0(net4378),
    .A1(\spiking_network_top_uut.all_data_out[653] ),
    .S(net3679),
    .X(_01678_));
 sg13g2_mux2_1 _18629_ (.A0(net4354),
    .A1(\spiking_network_top_uut.all_data_out[654] ),
    .S(net3679),
    .X(_01679_));
 sg13g2_mux2_1 _18630_ (.A0(net4333),
    .A1(\spiking_network_top_uut.all_data_out[655] ),
    .S(net3679),
    .X(_01680_));
 sg13g2_nor2_2 _18631_ (.A(_03218_),
    .B(net3725),
    .Y(_03327_));
 sg13g2_mux2_1 _18632_ (.A0(\spiking_network_top_uut.all_data_out[176] ),
    .A1(net4467),
    .S(_03327_),
    .X(_01681_));
 sg13g2_mux2_1 _18633_ (.A0(\spiking_network_top_uut.all_data_out[177] ),
    .A1(net4447),
    .S(_03327_),
    .X(_01682_));
 sg13g2_mux2_1 _18634_ (.A0(\spiking_network_top_uut.all_data_out[178] ),
    .A1(net4427),
    .S(_03327_),
    .X(_01683_));
 sg13g2_mux2_1 _18635_ (.A0(\spiking_network_top_uut.all_data_out[179] ),
    .A1(net4409),
    .S(_03327_),
    .X(_01684_));
 sg13g2_mux2_1 _18636_ (.A0(\spiking_network_top_uut.all_data_out[180] ),
    .A1(net4385),
    .S(_03327_),
    .X(_01685_));
 sg13g2_mux2_1 _18637_ (.A0(\spiking_network_top_uut.all_data_out[181] ),
    .A1(net4366),
    .S(_03327_),
    .X(_01686_));
 sg13g2_mux2_1 _18638_ (.A0(\spiking_network_top_uut.all_data_out[182] ),
    .A1(net4343),
    .S(_03327_),
    .X(_01687_));
 sg13g2_mux2_1 _18639_ (.A0(\spiking_network_top_uut.all_data_out[183] ),
    .A1(net4325),
    .S(_03327_),
    .X(_01688_));
 sg13g2_nor2_1 _18640_ (.A(_03225_),
    .B(net3728),
    .Y(_03328_));
 sg13g2_mux2_1 _18641_ (.A0(\spiking_network_top_uut.all_data_out[808] ),
    .A1(net4476),
    .S(net3678),
    .X(_01689_));
 sg13g2_mux2_1 _18642_ (.A0(\spiking_network_top_uut.all_data_out[809] ),
    .A1(net4456),
    .S(net3678),
    .X(_01690_));
 sg13g2_mux2_1 _18643_ (.A0(\spiking_network_top_uut.all_data_out[810] ),
    .A1(net4435),
    .S(net3678),
    .X(_01691_));
 sg13g2_mux2_1 _18644_ (.A0(\spiking_network_top_uut.all_data_out[811] ),
    .A1(net4417),
    .S(net3678),
    .X(_01692_));
 sg13g2_mux2_1 _18645_ (.A0(\spiking_network_top_uut.all_data_out[812] ),
    .A1(net4394),
    .S(_03328_),
    .X(_01693_));
 sg13g2_mux2_1 _18646_ (.A0(\spiking_network_top_uut.all_data_out[813] ),
    .A1(net4372),
    .S(net3678),
    .X(_01694_));
 sg13g2_nand2_1 _18647_ (.Y(_03329_),
    .A(net4353),
    .B(net3678));
 sg13g2_o21ai_1 _18648_ (.B1(_03329_),
    .Y(_01695_),
    .A1(_03511_),
    .A2(net3678));
 sg13g2_mux2_1 _18649_ (.A0(\spiking_network_top_uut.all_data_out[815] ),
    .A1(net4334),
    .S(net3678),
    .X(_01696_));
 sg13g2_nor2_2 _18650_ (.A(_03225_),
    .B(net3726),
    .Y(_03330_));
 sg13g2_mux2_1 _18651_ (.A0(\spiking_network_top_uut.all_data_out[168] ),
    .A1(net4468),
    .S(_03330_),
    .X(_01697_));
 sg13g2_mux2_1 _18652_ (.A0(\spiking_network_top_uut.all_data_out[169] ),
    .A1(net4446),
    .S(_03330_),
    .X(_01698_));
 sg13g2_mux2_1 _18653_ (.A0(\spiking_network_top_uut.all_data_out[170] ),
    .A1(net4427),
    .S(_03330_),
    .X(_01699_));
 sg13g2_mux2_1 _18654_ (.A0(\spiking_network_top_uut.all_data_out[171] ),
    .A1(net4409),
    .S(_03330_),
    .X(_01700_));
 sg13g2_mux2_1 _18655_ (.A0(\spiking_network_top_uut.all_data_out[172] ),
    .A1(net4386),
    .S(_03330_),
    .X(_01701_));
 sg13g2_mux2_1 _18656_ (.A0(\spiking_network_top_uut.all_data_out[173] ),
    .A1(net4366),
    .S(_03330_),
    .X(_01702_));
 sg13g2_mux2_1 _18657_ (.A0(\spiking_network_top_uut.all_data_out[174] ),
    .A1(net4344),
    .S(_03330_),
    .X(_01703_));
 sg13g2_mux2_1 _18658_ (.A0(\spiking_network_top_uut.all_data_out[175] ),
    .A1(net4325),
    .S(_03330_),
    .X(_01704_));
 sg13g2_nor2_2 _18659_ (.A(net3736),
    .B(_03215_),
    .Y(_03331_));
 sg13g2_mux2_1 _18660_ (.A0(\spiking_network_top_uut.all_data_out[488] ),
    .A1(net4477),
    .S(_03331_),
    .X(_01705_));
 sg13g2_mux2_1 _18661_ (.A0(\spiking_network_top_uut.all_data_out[489] ),
    .A1(net4457),
    .S(net3677),
    .X(_01706_));
 sg13g2_nand2_1 _18662_ (.Y(_03332_),
    .A(net4436),
    .B(net3677));
 sg13g2_o21ai_1 _18663_ (.B1(_03332_),
    .Y(_01707_),
    .A1(_03617_),
    .A2(net3677));
 sg13g2_mux2_1 _18664_ (.A0(\spiking_network_top_uut.all_data_out[491] ),
    .A1(net4418),
    .S(net3677),
    .X(_01708_));
 sg13g2_mux2_1 _18665_ (.A0(\spiking_network_top_uut.all_data_out[492] ),
    .A1(net4396),
    .S(net3677),
    .X(_01709_));
 sg13g2_mux2_1 _18666_ (.A0(\spiking_network_top_uut.all_data_out[493] ),
    .A1(net4375),
    .S(net3677),
    .X(_01710_));
 sg13g2_mux2_1 _18667_ (.A0(\spiking_network_top_uut.all_data_out[494] ),
    .A1(net4355),
    .S(net3677),
    .X(_01711_));
 sg13g2_mux2_1 _18668_ (.A0(\spiking_network_top_uut.all_data_out[495] ),
    .A1(net4335),
    .S(net3677),
    .X(_01712_));
 sg13g2_nor2_2 _18669_ (.A(_03231_),
    .B(net3726),
    .Y(_03333_));
 sg13g2_mux2_1 _18670_ (.A0(\spiking_network_top_uut.all_data_out[160] ),
    .A1(net4467),
    .S(_03333_),
    .X(_01713_));
 sg13g2_mux2_1 _18671_ (.A0(\spiking_network_top_uut.all_data_out[161] ),
    .A1(net4447),
    .S(_03333_),
    .X(_01714_));
 sg13g2_mux2_1 _18672_ (.A0(\spiking_network_top_uut.all_data_out[162] ),
    .A1(net4426),
    .S(_03333_),
    .X(_01715_));
 sg13g2_mux2_1 _18673_ (.A0(\spiking_network_top_uut.all_data_out[163] ),
    .A1(net4405),
    .S(_03333_),
    .X(_01716_));
 sg13g2_mux2_1 _18674_ (.A0(\spiking_network_top_uut.all_data_out[164] ),
    .A1(net4385),
    .S(_03333_),
    .X(_01717_));
 sg13g2_mux2_1 _18675_ (.A0(\spiking_network_top_uut.all_data_out[165] ),
    .A1(net4364),
    .S(_03333_),
    .X(_01718_));
 sg13g2_mux2_1 _18676_ (.A0(\spiking_network_top_uut.all_data_out[166] ),
    .A1(net4343),
    .S(_03333_),
    .X(_01719_));
 sg13g2_mux2_1 _18677_ (.A0(\spiking_network_top_uut.all_data_out[167] ),
    .A1(net4322),
    .S(_03333_),
    .X(_01720_));
 sg13g2_nor2_1 _18678_ (.A(_03218_),
    .B(net3728),
    .Y(_03334_));
 sg13g2_mux2_1 _18679_ (.A0(\spiking_network_top_uut.all_data_out[816] ),
    .A1(net4473),
    .S(net3676),
    .X(_01721_));
 sg13g2_mux2_1 _18680_ (.A0(\spiking_network_top_uut.all_data_out[817] ),
    .A1(net4452),
    .S(net3676),
    .X(_01722_));
 sg13g2_nand2_1 _18681_ (.Y(_03335_),
    .A(net4432),
    .B(net3676));
 sg13g2_o21ai_1 _18682_ (.B1(_03335_),
    .Y(_01723_),
    .A1(_03583_),
    .A2(net3676));
 sg13g2_mux2_1 _18683_ (.A0(\spiking_network_top_uut.all_data_out[819] ),
    .A1(net4413),
    .S(net3676),
    .X(_01724_));
 sg13g2_mux2_1 _18684_ (.A0(\spiking_network_top_uut.all_data_out[820] ),
    .A1(net4394),
    .S(_03334_),
    .X(_01725_));
 sg13g2_mux2_1 _18685_ (.A0(\spiking_network_top_uut.all_data_out[821] ),
    .A1(net4372),
    .S(net3676),
    .X(_01726_));
 sg13g2_mux2_1 _18686_ (.A0(\spiking_network_top_uut.all_data_out[822] ),
    .A1(net4353),
    .S(net3676),
    .X(_01727_));
 sg13g2_mux2_1 _18687_ (.A0(\spiking_network_top_uut.all_data_out[823] ),
    .A1(net4331),
    .S(net3676),
    .X(_01728_));
 sg13g2_nand2_2 _18688_ (.Y(_03336_),
    .A(_03234_),
    .B(_03303_));
 sg13g2_mux2_1 _18689_ (.A0(net4469),
    .A1(\spiking_network_top_uut.all_data_out[152] ),
    .S(_03336_),
    .X(_01729_));
 sg13g2_mux2_1 _18690_ (.A0(net4444),
    .A1(\spiking_network_top_uut.all_data_out[153] ),
    .S(_03336_),
    .X(_01730_));
 sg13g2_mux2_1 _18691_ (.A0(net4428),
    .A1(\spiking_network_top_uut.all_data_out[154] ),
    .S(_03336_),
    .X(_01731_));
 sg13g2_mux2_1 _18692_ (.A0(net4406),
    .A1(\spiking_network_top_uut.all_data_out[155] ),
    .S(_03336_),
    .X(_01732_));
 sg13g2_mux2_1 _18693_ (.A0(net4382),
    .A1(\spiking_network_top_uut.all_data_out[156] ),
    .S(_03336_),
    .X(_01733_));
 sg13g2_mux2_1 _18694_ (.A0(net4365),
    .A1(\spiking_network_top_uut.all_data_out[157] ),
    .S(_03336_),
    .X(_01734_));
 sg13g2_mux2_1 _18695_ (.A0(net4345),
    .A1(\spiking_network_top_uut.all_data_out[158] ),
    .S(_03336_),
    .X(_01735_));
 sg13g2_mux2_1 _18696_ (.A0(net4322),
    .A1(\spiking_network_top_uut.all_data_out[159] ),
    .S(_03336_),
    .X(_01736_));
 sg13g2_nor2_2 _18697_ (.A(_03208_),
    .B(net3733),
    .Y(_03337_));
 sg13g2_mux2_1 _18698_ (.A0(\spiking_network_top_uut.all_data_out[568] ),
    .A1(net4478),
    .S(_03337_),
    .X(_01737_));
 sg13g2_mux2_1 _18699_ (.A0(\spiking_network_top_uut.all_data_out[569] ),
    .A1(net4458),
    .S(_03337_),
    .X(_01738_));
 sg13g2_mux2_1 _18700_ (.A0(\spiking_network_top_uut.all_data_out[570] ),
    .A1(net4437),
    .S(_03337_),
    .X(_01739_));
 sg13g2_mux2_1 _18701_ (.A0(\spiking_network_top_uut.all_data_out[571] ),
    .A1(net4414),
    .S(_03337_),
    .X(_01740_));
 sg13g2_mux2_1 _18702_ (.A0(\spiking_network_top_uut.all_data_out[572] ),
    .A1(net4398),
    .S(_03337_),
    .X(_01741_));
 sg13g2_mux2_1 _18703_ (.A0(\spiking_network_top_uut.all_data_out[573] ),
    .A1(net4377),
    .S(_03337_),
    .X(_01742_));
 sg13g2_mux2_1 _18704_ (.A0(\spiking_network_top_uut.all_data_out[574] ),
    .A1(net4358),
    .S(_03337_),
    .X(_01743_));
 sg13g2_mux2_1 _18705_ (.A0(\spiking_network_top_uut.all_data_out[575] ),
    .A1(net4329),
    .S(_03337_),
    .X(_01744_));
 sg13g2_nand2_2 _18706_ (.Y(_03338_),
    .A(_03240_),
    .B(_03303_));
 sg13g2_mux2_1 _18707_ (.A0(net4466),
    .A1(\spiking_network_top_uut.all_data_out[144] ),
    .S(_03338_),
    .X(_01745_));
 sg13g2_mux2_1 _18708_ (.A0(net4444),
    .A1(\spiking_network_top_uut.all_data_out[145] ),
    .S(_03338_),
    .X(_01746_));
 sg13g2_mux2_1 _18709_ (.A0(net4424),
    .A1(\spiking_network_top_uut.all_data_out[146] ),
    .S(_03338_),
    .X(_01747_));
 sg13g2_mux2_1 _18710_ (.A0(net4403),
    .A1(\spiking_network_top_uut.all_data_out[147] ),
    .S(_03338_),
    .X(_01748_));
 sg13g2_mux2_1 _18711_ (.A0(net4384),
    .A1(\spiking_network_top_uut.all_data_out[148] ),
    .S(_03338_),
    .X(_01749_));
 sg13g2_mux2_1 _18712_ (.A0(net4365),
    .A1(\spiking_network_top_uut.all_data_out[149] ),
    .S(_03338_),
    .X(_01750_));
 sg13g2_mux2_1 _18713_ (.A0(net4341),
    .A1(\spiking_network_top_uut.all_data_out[150] ),
    .S(_03338_),
    .X(_01751_));
 sg13g2_mux2_1 _18714_ (.A0(net4322),
    .A1(\spiking_network_top_uut.all_data_out[151] ),
    .S(_03338_),
    .X(_01752_));
 sg13g2_nor2_2 _18715_ (.A(_03208_),
    .B(net3728),
    .Y(_03339_));
 sg13g2_mux2_1 _18716_ (.A0(\spiking_network_top_uut.all_data_out[824] ),
    .A1(net4467),
    .S(_03339_),
    .X(_01753_));
 sg13g2_mux2_1 _18717_ (.A0(\spiking_network_top_uut.all_data_out[825] ),
    .A1(net4446),
    .S(_03339_),
    .X(_01754_));
 sg13g2_mux2_1 _18718_ (.A0(\spiking_network_top_uut.all_data_out[826] ),
    .A1(net4427),
    .S(_03339_),
    .X(_01755_));
 sg13g2_mux2_1 _18719_ (.A0(\spiking_network_top_uut.all_data_out[827] ),
    .A1(net4409),
    .S(_03339_),
    .X(_01756_));
 sg13g2_mux2_1 _18720_ (.A0(\spiking_network_top_uut.all_data_out[828] ),
    .A1(net4388),
    .S(_03339_),
    .X(_01757_));
 sg13g2_mux2_1 _18721_ (.A0(\spiking_network_top_uut.all_data_out[829] ),
    .A1(net4366),
    .S(_03339_),
    .X(_01758_));
 sg13g2_mux2_1 _18722_ (.A0(\spiking_network_top_uut.all_data_out[830] ),
    .A1(net4347),
    .S(_03339_),
    .X(_01759_));
 sg13g2_mux2_1 _18723_ (.A0(\spiking_network_top_uut.all_data_out[831] ),
    .A1(net4325),
    .S(_03339_),
    .X(_01760_));
 sg13g2_nand2_2 _18724_ (.Y(_03340_),
    .A(_03244_),
    .B(_03303_));
 sg13g2_mux2_1 _18725_ (.A0(net4472),
    .A1(\spiking_network_top_uut.all_data_out[136] ),
    .S(_03340_),
    .X(_01761_));
 sg13g2_mux2_1 _18726_ (.A0(net4451),
    .A1(\spiking_network_top_uut.all_data_out[137] ),
    .S(_03340_),
    .X(_01762_));
 sg13g2_mux2_1 _18727_ (.A0(net4433),
    .A1(\spiking_network_top_uut.all_data_out[138] ),
    .S(_03340_),
    .X(_01763_));
 sg13g2_mux2_1 _18728_ (.A0(net4410),
    .A1(\spiking_network_top_uut.all_data_out[139] ),
    .S(_03340_),
    .X(_01764_));
 sg13g2_mux2_1 _18729_ (.A0(net4390),
    .A1(\spiking_network_top_uut.all_data_out[140] ),
    .S(_03340_),
    .X(_01765_));
 sg13g2_mux2_1 _18730_ (.A0(net4371),
    .A1(\spiking_network_top_uut.all_data_out[141] ),
    .S(_03340_),
    .X(_01766_));
 sg13g2_mux2_1 _18731_ (.A0(net4349),
    .A1(\spiking_network_top_uut.all_data_out[142] ),
    .S(_03340_),
    .X(_01767_));
 sg13g2_mux2_1 _18732_ (.A0(net4327),
    .A1(\spiking_network_top_uut.all_data_out[143] ),
    .S(_03340_),
    .X(_01768_));
 sg13g2_nor2_2 _18733_ (.A(net3735),
    .B(_03268_),
    .Y(_03341_));
 sg13g2_mux2_1 _18734_ (.A0(\spiking_network_top_uut.all_data_out[480] ),
    .A1(net4478),
    .S(_03341_),
    .X(_01769_));
 sg13g2_mux2_1 _18735_ (.A0(\spiking_network_top_uut.all_data_out[481] ),
    .A1(net4458),
    .S(net3675),
    .X(_01770_));
 sg13g2_mux2_1 _18736_ (.A0(\spiking_network_top_uut.all_data_out[482] ),
    .A1(net4437),
    .S(net3675),
    .X(_01771_));
 sg13g2_mux2_1 _18737_ (.A0(\spiking_network_top_uut.all_data_out[483] ),
    .A1(net4410),
    .S(net3675),
    .X(_01772_));
 sg13g2_mux2_1 _18738_ (.A0(\spiking_network_top_uut.all_data_out[484] ),
    .A1(net4398),
    .S(net3675),
    .X(_01773_));
 sg13g2_mux2_1 _18739_ (.A0(\spiking_network_top_uut.all_data_out[485] ),
    .A1(net4377),
    .S(net3675),
    .X(_01774_));
 sg13g2_nand2_1 _18740_ (.Y(_03342_),
    .A(net4358),
    .B(net3675));
 sg13g2_o21ai_1 _18741_ (.B1(_03342_),
    .Y(_01775_),
    .A1(_03538_),
    .A2(net3675));
 sg13g2_mux2_1 _18742_ (.A0(\spiking_network_top_uut.all_data_out[487] ),
    .A1(net4329),
    .S(net3675),
    .X(_01776_));
 sg13g2_nand3_1 _18743_ (.B(_03200_),
    .C(_03303_),
    .A(net3737),
    .Y(_03343_));
 sg13g2_mux2_1 _18744_ (.A0(net4471),
    .A1(\spiking_network_top_uut.all_data_out[128] ),
    .S(_03343_),
    .X(_01777_));
 sg13g2_mux2_1 _18745_ (.A0(net4451),
    .A1(\spiking_network_top_uut.all_data_out[129] ),
    .S(_03343_),
    .X(_01778_));
 sg13g2_mux2_1 _18746_ (.A0(net4431),
    .A1(\spiking_network_top_uut.all_data_out[130] ),
    .S(_03343_),
    .X(_01779_));
 sg13g2_mux2_1 _18747_ (.A0(net4410),
    .A1(\spiking_network_top_uut.all_data_out[131] ),
    .S(_03343_),
    .X(_01780_));
 sg13g2_mux2_1 _18748_ (.A0(net4390),
    .A1(\spiking_network_top_uut.all_data_out[132] ),
    .S(_03343_),
    .X(_01781_));
 sg13g2_mux2_1 _18749_ (.A0(net4371),
    .A1(\spiking_network_top_uut.all_data_out[133] ),
    .S(_03343_),
    .X(_01782_));
 sg13g2_mux2_1 _18750_ (.A0(net4349),
    .A1(\spiking_network_top_uut.all_data_out[134] ),
    .S(_03343_),
    .X(_01783_));
 sg13g2_mux2_1 _18751_ (.A0(net4329),
    .A1(\spiking_network_top_uut.all_data_out[135] ),
    .S(_03343_),
    .X(_01784_));
 sg13g2_nor2_2 _18752_ (.A(_03250_),
    .B(net3727),
    .Y(_03344_));
 sg13g2_mux2_1 _18753_ (.A0(\spiking_network_top_uut.all_data_out[832] ),
    .A1(net4463),
    .S(_03344_),
    .X(_01785_));
 sg13g2_mux2_1 _18754_ (.A0(\spiking_network_top_uut.all_data_out[833] ),
    .A1(net4441),
    .S(_03344_),
    .X(_01786_));
 sg13g2_mux2_1 _18755_ (.A0(\spiking_network_top_uut.all_data_out[834] ),
    .A1(net4422),
    .S(_03344_),
    .X(_01787_));
 sg13g2_mux2_1 _18756_ (.A0(\spiking_network_top_uut.all_data_out[835] ),
    .A1(net4402),
    .S(_03344_),
    .X(_01788_));
 sg13g2_mux2_1 _18757_ (.A0(\spiking_network_top_uut.all_data_out[836] ),
    .A1(net4381),
    .S(_03344_),
    .X(_01789_));
 sg13g2_mux2_1 _18758_ (.A0(\spiking_network_top_uut.all_data_out[837] ),
    .A1(net4360),
    .S(_03344_),
    .X(_01790_));
 sg13g2_mux2_1 _18759_ (.A0(\spiking_network_top_uut.all_data_out[838] ),
    .A1(net4340),
    .S(_03344_),
    .X(_01791_));
 sg13g2_mux2_1 _18760_ (.A0(\spiking_network_top_uut.all_data_out[839] ),
    .A1(net4319),
    .S(_03344_),
    .X(_01792_));
 sg13g2_nand2b_2 _18761_ (.Y(_03345_),
    .B(_03210_),
    .A_N(\spiking_network_top_uut.spi_inst.LSB_Address_reg[6] ));
 sg13g2_nor2_2 _18762_ (.A(net15),
    .B(net3723),
    .Y(_03346_));
 sg13g2_mux2_1 _18763_ (.A0(\spiking_network_top_uut.all_data_out[120] ),
    .A1(net4472),
    .S(_03346_),
    .X(_01793_));
 sg13g2_mux2_1 _18764_ (.A0(\spiking_network_top_uut.all_data_out[121] ),
    .A1(net4451),
    .S(_03346_),
    .X(_01794_));
 sg13g2_mux2_1 _18765_ (.A0(\spiking_network_top_uut.all_data_out[122] ),
    .A1(net4431),
    .S(_03346_),
    .X(_01795_));
 sg13g2_mux2_1 _18766_ (.A0(\spiking_network_top_uut.all_data_out[123] ),
    .A1(net4410),
    .S(_03346_),
    .X(_01796_));
 sg13g2_mux2_1 _18767_ (.A0(\spiking_network_top_uut.all_data_out[124] ),
    .A1(net4390),
    .S(_03346_),
    .X(_01797_));
 sg13g2_mux2_1 _18768_ (.A0(\spiking_network_top_uut.all_data_out[125] ),
    .A1(net4367),
    .S(_03346_),
    .X(_01798_));
 sg13g2_mux2_1 _18769_ (.A0(\spiking_network_top_uut.all_data_out[126] ),
    .A1(net4349),
    .S(_03346_),
    .X(_01799_));
 sg13g2_mux2_1 _18770_ (.A0(\spiking_network_top_uut.all_data_out[127] ),
    .A1(net4327),
    .S(_03346_),
    .X(_01800_));
 sg13g2_nand2_2 _18771_ (.Y(_03347_),
    .A(_03223_),
    .B(_03240_));
 sg13g2_mux2_1 _18772_ (.A0(net4473),
    .A1(\spiking_network_top_uut.all_data_out[656] ),
    .S(_03347_),
    .X(_01801_));
 sg13g2_mux2_1 _18773_ (.A0(net4452),
    .A1(\spiking_network_top_uut.all_data_out[657] ),
    .S(_03347_),
    .X(_01802_));
 sg13g2_mux2_1 _18774_ (.A0(net4432),
    .A1(\spiking_network_top_uut.all_data_out[658] ),
    .S(_03347_),
    .X(_01803_));
 sg13g2_mux2_1 _18775_ (.A0(net4415),
    .A1(\spiking_network_top_uut.all_data_out[659] ),
    .S(_03347_),
    .X(_01804_));
 sg13g2_mux2_1 _18776_ (.A0(net4392),
    .A1(\spiking_network_top_uut.all_data_out[660] ),
    .S(_03347_),
    .X(_01805_));
 sg13g2_mux2_1 _18777_ (.A0(net4372),
    .A1(\spiking_network_top_uut.all_data_out[661] ),
    .S(_03347_),
    .X(_01806_));
 sg13g2_mux2_1 _18778_ (.A0(net4351),
    .A1(\spiking_network_top_uut.all_data_out[662] ),
    .S(_03347_),
    .X(_01807_));
 sg13g2_mux2_1 _18779_ (.A0(net4333),
    .A1(\spiking_network_top_uut.all_data_out[663] ),
    .S(_03347_),
    .X(_01808_));
 sg13g2_nor2_2 _18780_ (.A(_03258_),
    .B(net3723),
    .Y(_03348_));
 sg13g2_mux2_1 _18781_ (.A0(\spiking_network_top_uut.all_data_out[112] ),
    .A1(net4472),
    .S(_03348_),
    .X(_01809_));
 sg13g2_mux2_1 _18782_ (.A0(\spiking_network_top_uut.all_data_out[113] ),
    .A1(net4451),
    .S(_03348_),
    .X(_01810_));
 sg13g2_mux2_1 _18783_ (.A0(\spiking_network_top_uut.all_data_out[114] ),
    .A1(net4431),
    .S(_03348_),
    .X(_01811_));
 sg13g2_mux2_1 _18784_ (.A0(\spiking_network_top_uut.all_data_out[115] ),
    .A1(net4412),
    .S(_03348_),
    .X(_01812_));
 sg13g2_mux2_1 _18785_ (.A0(\spiking_network_top_uut.all_data_out[116] ),
    .A1(net4390),
    .S(_03348_),
    .X(_01813_));
 sg13g2_mux2_1 _18786_ (.A0(\spiking_network_top_uut.all_data_out[117] ),
    .A1(net4371),
    .S(_03348_),
    .X(_01814_));
 sg13g2_mux2_1 _18787_ (.A0(\spiking_network_top_uut.all_data_out[118] ),
    .A1(net4349),
    .S(_03348_),
    .X(_01815_));
 sg13g2_mux2_1 _18788_ (.A0(\spiking_network_top_uut.all_data_out[119] ),
    .A1(net4327),
    .S(_03348_),
    .X(_01816_));
 sg13g2_nor2_2 _18789_ (.A(_03238_),
    .B(net3727),
    .Y(_03349_));
 sg13g2_mux2_1 _18790_ (.A0(\spiking_network_top_uut.all_data_out[840] ),
    .A1(net4463),
    .S(_03349_),
    .X(_01817_));
 sg13g2_mux2_1 _18791_ (.A0(\spiking_network_top_uut.all_data_out[841] ),
    .A1(net4441),
    .S(net3674),
    .X(_01818_));
 sg13g2_nand2_1 _18792_ (.Y(_03350_),
    .A(net4422),
    .B(net3674));
 sg13g2_o21ai_1 _18793_ (.B1(_03350_),
    .Y(_01819_),
    .A1(_03581_),
    .A2(net3674));
 sg13g2_mux2_1 _18794_ (.A0(\spiking_network_top_uut.all_data_out[843] ),
    .A1(net4401),
    .S(net3674),
    .X(_01820_));
 sg13g2_mux2_1 _18795_ (.A0(\spiking_network_top_uut.all_data_out[844] ),
    .A1(net4381),
    .S(net3674),
    .X(_01821_));
 sg13g2_mux2_1 _18796_ (.A0(\spiking_network_top_uut.all_data_out[845] ),
    .A1(net4363),
    .S(net3674),
    .X(_01822_));
 sg13g2_mux2_1 _18797_ (.A0(\spiking_network_top_uut.all_data_out[846] ),
    .A1(net4340),
    .S(net3674),
    .X(_01823_));
 sg13g2_mux2_1 _18798_ (.A0(\spiking_network_top_uut.all_data_out[847] ),
    .A1(net4319),
    .S(net3674),
    .X(_01824_));
 sg13g2_nor2_2 _18799_ (.A(_03215_),
    .B(net3723),
    .Y(_03351_));
 sg13g2_mux2_1 _18800_ (.A0(\spiking_network_top_uut.all_data_out[104] ),
    .A1(net4471),
    .S(_03351_),
    .X(_01825_));
 sg13g2_mux2_1 _18801_ (.A0(\spiking_network_top_uut.all_data_out[105] ),
    .A1(net4451),
    .S(_03351_),
    .X(_01826_));
 sg13g2_mux2_1 _18802_ (.A0(\spiking_network_top_uut.all_data_out[106] ),
    .A1(net4431),
    .S(_03351_),
    .X(_01827_));
 sg13g2_mux2_1 _18803_ (.A0(\spiking_network_top_uut.all_data_out[107] ),
    .A1(net4410),
    .S(_03351_),
    .X(_01828_));
 sg13g2_mux2_1 _18804_ (.A0(\spiking_network_top_uut.all_data_out[108] ),
    .A1(net4390),
    .S(_03351_),
    .X(_01829_));
 sg13g2_mux2_1 _18805_ (.A0(\spiking_network_top_uut.all_data_out[109] ),
    .A1(net4366),
    .S(_03351_),
    .X(_01830_));
 sg13g2_mux2_1 _18806_ (.A0(\spiking_network_top_uut.all_data_out[110] ),
    .A1(net4349),
    .S(_03351_),
    .X(_01831_));
 sg13g2_mux2_1 _18807_ (.A0(\spiking_network_top_uut.all_data_out[111] ),
    .A1(net4329),
    .S(_03351_),
    .X(_01832_));
 sg13g2_nor2_2 _18808_ (.A(net3736),
    .B(_03272_),
    .Y(_03352_));
 sg13g2_mux2_1 _18809_ (.A0(\spiking_network_top_uut.all_data_out[472] ),
    .A1(net4479),
    .S(_03352_),
    .X(_01833_));
 sg13g2_mux2_1 _18810_ (.A0(\spiking_network_top_uut.all_data_out[473] ),
    .A1(net4458),
    .S(_03352_),
    .X(_01834_));
 sg13g2_mux2_1 _18811_ (.A0(\spiking_network_top_uut.all_data_out[474] ),
    .A1(net4437),
    .S(_03352_),
    .X(_01835_));
 sg13g2_mux2_1 _18812_ (.A0(\spiking_network_top_uut.all_data_out[475] ),
    .A1(net4420),
    .S(_03352_),
    .X(_01836_));
 sg13g2_mux2_1 _18813_ (.A0(\spiking_network_top_uut.all_data_out[476] ),
    .A1(net4398),
    .S(_03352_),
    .X(_01837_));
 sg13g2_mux2_1 _18814_ (.A0(\spiking_network_top_uut.all_data_out[477] ),
    .A1(net4377),
    .S(_03352_),
    .X(_01838_));
 sg13g2_mux2_1 _18815_ (.A0(\spiking_network_top_uut.all_data_out[478] ),
    .A1(net4358),
    .S(_03352_),
    .X(_01839_));
 sg13g2_mux2_1 _18816_ (.A0(\spiking_network_top_uut.all_data_out[479] ),
    .A1(net4337),
    .S(_03352_),
    .X(_01840_));
 sg13g2_nor2_2 _18817_ (.A(_03268_),
    .B(net3723),
    .Y(_03353_));
 sg13g2_mux2_1 _18818_ (.A0(\spiking_network_top_uut.all_data_out[96] ),
    .A1(net4472),
    .S(_03353_),
    .X(_01841_));
 sg13g2_mux2_1 _18819_ (.A0(\spiking_network_top_uut.all_data_out[97] ),
    .A1(net4450),
    .S(_03353_),
    .X(_01842_));
 sg13g2_mux2_1 _18820_ (.A0(\spiking_network_top_uut.all_data_out[98] ),
    .A1(net4431),
    .S(_03353_),
    .X(_01843_));
 sg13g2_mux2_1 _18821_ (.A0(\spiking_network_top_uut.all_data_out[99] ),
    .A1(net4410),
    .S(_03353_),
    .X(_01844_));
 sg13g2_mux2_1 _18822_ (.A0(\spiking_network_top_uut.all_data_out[100] ),
    .A1(net4390),
    .S(_03353_),
    .X(_01845_));
 sg13g2_mux2_1 _18823_ (.A0(\spiking_network_top_uut.all_data_out[101] ),
    .A1(net4367),
    .S(_03353_),
    .X(_01846_));
 sg13g2_mux2_1 _18824_ (.A0(\spiking_network_top_uut.all_data_out[102] ),
    .A1(net4349),
    .S(_03353_),
    .X(_01847_));
 sg13g2_mux2_1 _18825_ (.A0(\spiking_network_top_uut.all_data_out[103] ),
    .A1(net4327),
    .S(_03353_),
    .X(_01848_));
 sg13g2_nor2_2 _18826_ (.A(_03270_),
    .B(net3727),
    .Y(_03354_));
 sg13g2_mux2_1 _18827_ (.A0(\spiking_network_top_uut.all_data_out[848] ),
    .A1(net4464),
    .S(_03354_),
    .X(_01849_));
 sg13g2_mux2_1 _18828_ (.A0(\spiking_network_top_uut.all_data_out[849] ),
    .A1(net4443),
    .S(_03354_),
    .X(_01850_));
 sg13g2_mux2_1 _18829_ (.A0(\spiking_network_top_uut.all_data_out[850] ),
    .A1(net4425),
    .S(_03354_),
    .X(_01851_));
 sg13g2_mux2_1 _18830_ (.A0(\spiking_network_top_uut.all_data_out[851] ),
    .A1(net4403),
    .S(_03354_),
    .X(_01852_));
 sg13g2_mux2_1 _18831_ (.A0(\spiking_network_top_uut.all_data_out[852] ),
    .A1(net4380),
    .S(_03354_),
    .X(_01853_));
 sg13g2_mux2_1 _18832_ (.A0(\spiking_network_top_uut.all_data_out[853] ),
    .A1(net4361),
    .S(_03354_),
    .X(_01854_));
 sg13g2_mux2_1 _18833_ (.A0(\spiking_network_top_uut.all_data_out[854] ),
    .A1(net4342),
    .S(_03354_),
    .X(_01855_));
 sg13g2_mux2_1 _18834_ (.A0(\spiking_network_top_uut.all_data_out[855] ),
    .A1(net4321),
    .S(_03354_),
    .X(_01856_));
 sg13g2_nor2_2 _18835_ (.A(net14),
    .B(net3724),
    .Y(_03355_));
 sg13g2_mux2_1 _18836_ (.A0(\spiking_network_top_uut.all_data_out[88] ),
    .A1(net4466),
    .S(_03355_),
    .X(_01857_));
 sg13g2_mux2_1 _18837_ (.A0(\spiking_network_top_uut.all_data_out[89] ),
    .A1(net4447),
    .S(_03355_),
    .X(_01858_));
 sg13g2_mux2_1 _18838_ (.A0(\spiking_network_top_uut.all_data_out[90] ),
    .A1(net4425),
    .S(_03355_),
    .X(_01859_));
 sg13g2_mux2_1 _18839_ (.A0(\spiking_network_top_uut.all_data_out[91] ),
    .A1(net4406),
    .S(_03355_),
    .X(_01860_));
 sg13g2_mux2_1 _18840_ (.A0(\spiking_network_top_uut.all_data_out[92] ),
    .A1(net4382),
    .S(_03355_),
    .X(_01861_));
 sg13g2_mux2_1 _18841_ (.A0(\spiking_network_top_uut.all_data_out[93] ),
    .A1(net4364),
    .S(_03355_),
    .X(_01862_));
 sg13g2_mux2_1 _18842_ (.A0(\spiking_network_top_uut.all_data_out[94] ),
    .A1(net4341),
    .S(_03355_),
    .X(_01863_));
 sg13g2_mux2_1 _18843_ (.A0(\spiking_network_top_uut.all_data_out[95] ),
    .A1(net4322),
    .S(_03355_),
    .X(_01864_));
 sg13g2_nor2_2 _18844_ (.A(net3734),
    .B(net14),
    .Y(_03356_));
 sg13g2_mux2_1 _18845_ (.A0(\spiking_network_top_uut.all_data_out[600] ),
    .A1(net4467),
    .S(_03356_),
    .X(_01865_));
 sg13g2_mux2_1 _18846_ (.A0(\spiking_network_top_uut.all_data_out[601] ),
    .A1(net4446),
    .S(_03356_),
    .X(_01866_));
 sg13g2_mux2_1 _18847_ (.A0(\spiking_network_top_uut.all_data_out[602] ),
    .A1(net4427),
    .S(_03356_),
    .X(_01867_));
 sg13g2_mux2_1 _18848_ (.A0(\spiking_network_top_uut.all_data_out[603] ),
    .A1(net4409),
    .S(_03356_),
    .X(_01868_));
 sg13g2_mux2_1 _18849_ (.A0(\spiking_network_top_uut.all_data_out[604] ),
    .A1(net4388),
    .S(_03356_),
    .X(_01869_));
 sg13g2_mux2_1 _18850_ (.A0(\spiking_network_top_uut.all_data_out[605] ),
    .A1(net4369),
    .S(_03356_),
    .X(_01870_));
 sg13g2_mux2_1 _18851_ (.A0(\spiking_network_top_uut.all_data_out[606] ),
    .A1(net4347),
    .S(_03356_),
    .X(_01871_));
 sg13g2_mux2_1 _18852_ (.A0(\spiking_network_top_uut.all_data_out[607] ),
    .A1(net4328),
    .S(_03356_),
    .X(_01872_));
 sg13g2_nor2_2 _18853_ (.A(_03270_),
    .B(net3724),
    .Y(_03357_));
 sg13g2_mux2_1 _18854_ (.A0(\spiking_network_top_uut.all_data_out[80] ),
    .A1(net4466),
    .S(_03357_),
    .X(_01873_));
 sg13g2_mux2_1 _18855_ (.A0(\spiking_network_top_uut.all_data_out[81] ),
    .A1(net4444),
    .S(_03357_),
    .X(_01874_));
 sg13g2_mux2_1 _18856_ (.A0(\spiking_network_top_uut.all_data_out[82] ),
    .A1(net4425),
    .S(_03357_),
    .X(_01875_));
 sg13g2_mux2_1 _18857_ (.A0(\spiking_network_top_uut.all_data_out[83] ),
    .A1(net4406),
    .S(_03357_),
    .X(_01876_));
 sg13g2_mux2_1 _18858_ (.A0(\spiking_network_top_uut.all_data_out[84] ),
    .A1(net4382),
    .S(_03357_),
    .X(_01877_));
 sg13g2_mux2_1 _18859_ (.A0(\spiking_network_top_uut.all_data_out[85] ),
    .A1(net4364),
    .S(_03357_),
    .X(_01878_));
 sg13g2_mux2_1 _18860_ (.A0(\spiking_network_top_uut.all_data_out[86] ),
    .A1(net4341),
    .S(_03357_),
    .X(_01879_));
 sg13g2_mux2_1 _18861_ (.A0(\spiking_network_top_uut.all_data_out[87] ),
    .A1(net4321),
    .S(_03357_),
    .X(_01880_));
 sg13g2_nor2_2 _18862_ (.A(net14),
    .B(net3727),
    .Y(_03358_));
 sg13g2_mux2_1 _18863_ (.A0(\spiking_network_top_uut.all_data_out[856] ),
    .A1(net4465),
    .S(_03358_),
    .X(_01881_));
 sg13g2_mux2_1 _18864_ (.A0(\spiking_network_top_uut.all_data_out[857] ),
    .A1(net4443),
    .S(_03358_),
    .X(_01882_));
 sg13g2_mux2_1 _18865_ (.A0(\spiking_network_top_uut.all_data_out[858] ),
    .A1(net4425),
    .S(_03358_),
    .X(_01883_));
 sg13g2_mux2_1 _18866_ (.A0(\spiking_network_top_uut.all_data_out[859] ),
    .A1(net4405),
    .S(_03358_),
    .X(_01884_));
 sg13g2_mux2_1 _18867_ (.A0(\spiking_network_top_uut.all_data_out[860] ),
    .A1(net4384),
    .S(_03358_),
    .X(_01885_));
 sg13g2_mux2_1 _18868_ (.A0(\spiking_network_top_uut.all_data_out[861] ),
    .A1(net4361),
    .S(_03358_),
    .X(_01886_));
 sg13g2_mux2_1 _18869_ (.A0(\spiking_network_top_uut.all_data_out[862] ),
    .A1(net4342),
    .S(_03358_),
    .X(_01887_));
 sg13g2_mux2_1 _18870_ (.A0(\spiking_network_top_uut.all_data_out[863] ),
    .A1(net4320),
    .S(_03358_),
    .X(_01888_));
 sg13g2_nor2_2 _18871_ (.A(_03238_),
    .B(net3724),
    .Y(_03359_));
 sg13g2_mux2_1 _18872_ (.A0(\spiking_network_top_uut.all_data_out[72] ),
    .A1(net4469),
    .S(_03359_),
    .X(_01889_));
 sg13g2_mux2_1 _18873_ (.A0(\spiking_network_top_uut.all_data_out[73] ),
    .A1(net4447),
    .S(_03359_),
    .X(_01890_));
 sg13g2_mux2_1 _18874_ (.A0(\spiking_network_top_uut.all_data_out[74] ),
    .A1(net4428),
    .S(_03359_),
    .X(_01891_));
 sg13g2_mux2_1 _18875_ (.A0(\spiking_network_top_uut.all_data_out[75] ),
    .A1(net4408),
    .S(_03359_),
    .X(_01892_));
 sg13g2_mux2_1 _18876_ (.A0(\spiking_network_top_uut.all_data_out[76] ),
    .A1(net4385),
    .S(_03359_),
    .X(_01893_));
 sg13g2_mux2_1 _18877_ (.A0(\spiking_network_top_uut.all_data_out[77] ),
    .A1(net4364),
    .S(_03359_),
    .X(_01894_));
 sg13g2_mux2_1 _18878_ (.A0(\spiking_network_top_uut.all_data_out[78] ),
    .A1(net4343),
    .S(_03359_),
    .X(_01895_));
 sg13g2_mux2_1 _18879_ (.A0(\spiking_network_top_uut.all_data_out[79] ),
    .A1(net4326),
    .S(_03359_),
    .X(_01896_));
 sg13g2_nor2_1 _18880_ (.A(net3735),
    .B(_03270_),
    .Y(_03360_));
 sg13g2_mux2_1 _18881_ (.A0(\spiking_network_top_uut.all_data_out[464] ),
    .A1(net4475),
    .S(net3673),
    .X(_01897_));
 sg13g2_mux2_1 _18882_ (.A0(\spiking_network_top_uut.all_data_out[465] ),
    .A1(net4455),
    .S(net3673),
    .X(_01898_));
 sg13g2_nand2_1 _18883_ (.Y(_03361_),
    .A(net4434),
    .B(net3673));
 sg13g2_o21ai_1 _18884_ (.B1(_03361_),
    .Y(_01899_),
    .A1(_03621_),
    .A2(net3673));
 sg13g2_mux2_1 _18885_ (.A0(\spiking_network_top_uut.all_data_out[467] ),
    .A1(net4419),
    .S(_03360_),
    .X(_01900_));
 sg13g2_mux2_1 _18886_ (.A0(\spiking_network_top_uut.all_data_out[468] ),
    .A1(net4390),
    .S(net3673),
    .X(_01901_));
 sg13g2_mux2_1 _18887_ (.A0(\spiking_network_top_uut.all_data_out[469] ),
    .A1(net4373),
    .S(net3673),
    .X(_01902_));
 sg13g2_mux2_1 _18888_ (.A0(\spiking_network_top_uut.all_data_out[470] ),
    .A1(net4350),
    .S(net3673),
    .X(_01903_));
 sg13g2_mux2_1 _18889_ (.A0(\spiking_network_top_uut.all_data_out[471] ),
    .A1(net4329),
    .S(net3673),
    .X(_01904_));
 sg13g2_nor2_2 _18890_ (.A(_03250_),
    .B(net3724),
    .Y(_03362_));
 sg13g2_mux2_1 _18891_ (.A0(\spiking_network_top_uut.all_data_out[64] ),
    .A1(net4469),
    .S(_03362_),
    .X(_01905_));
 sg13g2_mux2_1 _18892_ (.A0(\spiking_network_top_uut.all_data_out[65] ),
    .A1(net4447),
    .S(_03362_),
    .X(_01906_));
 sg13g2_mux2_1 _18893_ (.A0(\spiking_network_top_uut.all_data_out[66] ),
    .A1(net4428),
    .S(_03362_),
    .X(_01907_));
 sg13g2_mux2_1 _18894_ (.A0(\spiking_network_top_uut.all_data_out[67] ),
    .A1(net4408),
    .S(_03362_),
    .X(_01908_));
 sg13g2_mux2_1 _18895_ (.A0(\spiking_network_top_uut.all_data_out[68] ),
    .A1(net4385),
    .S(_03362_),
    .X(_01909_));
 sg13g2_mux2_1 _18896_ (.A0(\spiking_network_top_uut.all_data_out[69] ),
    .A1(net4364),
    .S(_03362_),
    .X(_01910_));
 sg13g2_mux2_1 _18897_ (.A0(\spiking_network_top_uut.all_data_out[70] ),
    .A1(net4343),
    .S(_03362_),
    .X(_01911_));
 sg13g2_mux2_1 _18898_ (.A0(\spiking_network_top_uut.all_data_out[71] ),
    .A1(net4326),
    .S(_03362_),
    .X(_01912_));
 sg13g2_nor2_2 _18899_ (.A(_03268_),
    .B(net3727),
    .Y(_03363_));
 sg13g2_mux2_1 _18900_ (.A0(\spiking_network_top_uut.all_data_out[864] ),
    .A1(net4463),
    .S(_03363_),
    .X(_01913_));
 sg13g2_mux2_1 _18901_ (.A0(\spiking_network_top_uut.all_data_out[865] ),
    .A1(net4441),
    .S(_03363_),
    .X(_01914_));
 sg13g2_mux2_1 _18902_ (.A0(\spiking_network_top_uut.all_data_out[866] ),
    .A1(net4422),
    .S(_03363_),
    .X(_01915_));
 sg13g2_mux2_1 _18903_ (.A0(\spiking_network_top_uut.all_data_out[867] ),
    .A1(net4401),
    .S(_03363_),
    .X(_01916_));
 sg13g2_mux2_1 _18904_ (.A0(\spiking_network_top_uut.all_data_out[868] ),
    .A1(net4381),
    .S(_03363_),
    .X(_01917_));
 sg13g2_mux2_1 _18905_ (.A0(\spiking_network_top_uut.all_data_out[869] ),
    .A1(net4360),
    .S(_03363_),
    .X(_01918_));
 sg13g2_mux2_1 _18906_ (.A0(\spiking_network_top_uut.all_data_out[870] ),
    .A1(net4340),
    .S(_03363_),
    .X(_01919_));
 sg13g2_mux2_1 _18907_ (.A0(\spiking_network_top_uut.all_data_out[871] ),
    .A1(net4319),
    .S(_03363_),
    .X(_01920_));
 sg13g2_nor2_2 _18908_ (.A(_03208_),
    .B(net3724),
    .Y(_03364_));
 sg13g2_mux2_1 _18909_ (.A0(\spiking_network_top_uut.all_data_out[56] ),
    .A1(net4469),
    .S(_03364_),
    .X(_01921_));
 sg13g2_mux2_1 _18910_ (.A0(\spiking_network_top_uut.all_data_out[57] ),
    .A1(net4451),
    .S(_03364_),
    .X(_01922_));
 sg13g2_mux2_1 _18911_ (.A0(\spiking_network_top_uut.all_data_out[58] ),
    .A1(net4431),
    .S(_03364_),
    .X(_01923_));
 sg13g2_mux2_1 _18912_ (.A0(\spiking_network_top_uut.all_data_out[59] ),
    .A1(net4408),
    .S(_03364_),
    .X(_01924_));
 sg13g2_mux2_1 _18913_ (.A0(\spiking_network_top_uut.all_data_out[60] ),
    .A1(net4386),
    .S(_03364_),
    .X(_01925_));
 sg13g2_mux2_1 _18914_ (.A0(\spiking_network_top_uut.all_data_out[61] ),
    .A1(net4367),
    .S(_03364_),
    .X(_01926_));
 sg13g2_mux2_1 _18915_ (.A0(\spiking_network_top_uut.all_data_out[62] ),
    .A1(net4343),
    .S(_03364_),
    .X(_01927_));
 sg13g2_mux2_1 _18916_ (.A0(\spiking_network_top_uut.all_data_out[63] ),
    .A1(net4326),
    .S(_03364_),
    .X(_01928_));
 sg13g2_nand2_2 _18917_ (.Y(_03365_),
    .A(_03223_),
    .B(_03234_));
 sg13g2_mux2_1 _18918_ (.A0(net4467),
    .A1(\spiking_network_top_uut.all_data_out[664] ),
    .S(_03365_),
    .X(_01929_));
 sg13g2_mux2_1 _18919_ (.A0(net4446),
    .A1(\spiking_network_top_uut.all_data_out[665] ),
    .S(_03365_),
    .X(_01930_));
 sg13g2_mux2_1 _18920_ (.A0(net4430),
    .A1(\spiking_network_top_uut.all_data_out[666] ),
    .S(_03365_),
    .X(_01931_));
 sg13g2_mux2_1 _18921_ (.A0(net4409),
    .A1(\spiking_network_top_uut.all_data_out[667] ),
    .S(_03365_),
    .X(_01932_));
 sg13g2_mux2_1 _18922_ (.A0(net4388),
    .A1(\spiking_network_top_uut.all_data_out[668] ),
    .S(_03365_),
    .X(_01933_));
 sg13g2_mux2_1 _18923_ (.A0(net4369),
    .A1(\spiking_network_top_uut.all_data_out[669] ),
    .S(_03365_),
    .X(_01934_));
 sg13g2_mux2_1 _18924_ (.A0(net4347),
    .A1(\spiking_network_top_uut.all_data_out[670] ),
    .S(_03365_),
    .X(_01935_));
 sg13g2_mux2_1 _18925_ (.A0(net4325),
    .A1(\spiking_network_top_uut.all_data_out[671] ),
    .S(_03365_),
    .X(_01936_));
 sg13g2_nor2_2 _18926_ (.A(_03218_),
    .B(net3724),
    .Y(_03366_));
 sg13g2_mux2_1 _18927_ (.A0(\spiking_network_top_uut.all_data_out[48] ),
    .A1(net4469),
    .S(_03366_),
    .X(_01937_));
 sg13g2_mux2_1 _18928_ (.A0(\spiking_network_top_uut.all_data_out[49] ),
    .A1(net4447),
    .S(_03366_),
    .X(_01938_));
 sg13g2_mux2_1 _18929_ (.A0(\spiking_network_top_uut.all_data_out[50] ),
    .A1(net4428),
    .S(_03366_),
    .X(_01939_));
 sg13g2_mux2_1 _18930_ (.A0(\spiking_network_top_uut.all_data_out[51] ),
    .A1(net4408),
    .S(_03366_),
    .X(_01940_));
 sg13g2_mux2_1 _18931_ (.A0(\spiking_network_top_uut.all_data_out[52] ),
    .A1(net4385),
    .S(_03366_),
    .X(_01941_));
 sg13g2_mux2_1 _18932_ (.A0(\spiking_network_top_uut.all_data_out[53] ),
    .A1(net4367),
    .S(_03366_),
    .X(_01942_));
 sg13g2_mux2_1 _18933_ (.A0(\spiking_network_top_uut.all_data_out[54] ),
    .A1(net4343),
    .S(_03366_),
    .X(_01943_));
 sg13g2_mux2_1 _18934_ (.A0(\spiking_network_top_uut.all_data_out[55] ),
    .A1(net4327),
    .S(_03366_),
    .X(_01944_));
 sg13g2_nor2_2 _18935_ (.A(_03215_),
    .B(net3727),
    .Y(_03367_));
 sg13g2_mux2_1 _18936_ (.A0(\spiking_network_top_uut.all_data_out[872] ),
    .A1(net4462),
    .S(_03367_),
    .X(_01945_));
 sg13g2_mux2_1 _18937_ (.A0(\spiking_network_top_uut.all_data_out[873] ),
    .A1(net4441),
    .S(_03367_),
    .X(_01946_));
 sg13g2_mux2_1 _18938_ (.A0(\spiking_network_top_uut.all_data_out[874] ),
    .A1(net4422),
    .S(_03367_),
    .X(_01947_));
 sg13g2_mux2_1 _18939_ (.A0(\spiking_network_top_uut.all_data_out[875] ),
    .A1(net4401),
    .S(_03367_),
    .X(_01948_));
 sg13g2_mux2_1 _18940_ (.A0(\spiking_network_top_uut.all_data_out[876] ),
    .A1(net4381),
    .S(_03367_),
    .X(_01949_));
 sg13g2_mux2_1 _18941_ (.A0(\spiking_network_top_uut.all_data_out[877] ),
    .A1(net4360),
    .S(_03367_),
    .X(_01950_));
 sg13g2_mux2_1 _18942_ (.A0(\spiking_network_top_uut.all_data_out[878] ),
    .A1(net4340),
    .S(_03367_),
    .X(_01951_));
 sg13g2_mux2_1 _18943_ (.A0(\spiking_network_top_uut.all_data_out[879] ),
    .A1(net4319),
    .S(_03367_),
    .X(_01952_));
 sg13g2_nor2_2 _18944_ (.A(_03225_),
    .B(net3723),
    .Y(_03368_));
 sg13g2_mux2_1 _18945_ (.A0(\spiking_network_top_uut.all_data_out[40] ),
    .A1(net4474),
    .S(_03368_),
    .X(_01953_));
 sg13g2_mux2_1 _18946_ (.A0(\spiking_network_top_uut.all_data_out[41] ),
    .A1(net4453),
    .S(_03368_),
    .X(_01954_));
 sg13g2_mux2_1 _18947_ (.A0(\spiking_network_top_uut.all_data_out[42] ),
    .A1(net4433),
    .S(_03368_),
    .X(_01955_));
 sg13g2_mux2_1 _18948_ (.A0(\spiking_network_top_uut.all_data_out[43] ),
    .A1(net4414),
    .S(_03368_),
    .X(_01956_));
 sg13g2_mux2_1 _18949_ (.A0(\spiking_network_top_uut.all_data_out[44] ),
    .A1(net4393),
    .S(_03368_),
    .X(_01957_));
 sg13g2_mux2_1 _18950_ (.A0(\spiking_network_top_uut.all_data_out[45] ),
    .A1(net4374),
    .S(_03368_),
    .X(_01958_));
 sg13g2_mux2_1 _18951_ (.A0(\spiking_network_top_uut.all_data_out[46] ),
    .A1(net4352),
    .S(_03368_),
    .X(_01959_));
 sg13g2_mux2_1 _18952_ (.A0(\spiking_network_top_uut.all_data_out[47] ),
    .A1(net4332),
    .S(_03368_),
    .X(_01960_));
 sg13g2_nor2_2 _18953_ (.A(net3736),
    .B(_03238_),
    .Y(_03369_));
 sg13g2_mux2_1 _18954_ (.A0(\spiking_network_top_uut.all_data_out[456] ),
    .A1(net4477),
    .S(_03369_),
    .X(_01961_));
 sg13g2_mux2_1 _18955_ (.A0(\spiking_network_top_uut.all_data_out[457] ),
    .A1(net4457),
    .S(_03369_),
    .X(_01962_));
 sg13g2_mux2_1 _18956_ (.A0(\spiking_network_top_uut.all_data_out[458] ),
    .A1(net4436),
    .S(_03369_),
    .X(_01963_));
 sg13g2_mux2_1 _18957_ (.A0(\spiking_network_top_uut.all_data_out[459] ),
    .A1(net4418),
    .S(_03369_),
    .X(_01964_));
 sg13g2_mux2_1 _18958_ (.A0(\spiking_network_top_uut.all_data_out[460] ),
    .A1(net4396),
    .S(_03369_),
    .X(_01965_));
 sg13g2_mux2_1 _18959_ (.A0(\spiking_network_top_uut.all_data_out[461] ),
    .A1(net4375),
    .S(_03369_),
    .X(_01966_));
 sg13g2_mux2_1 _18960_ (.A0(\spiking_network_top_uut.all_data_out[462] ),
    .A1(net4355),
    .S(_03369_),
    .X(_01967_));
 sg13g2_mux2_1 _18961_ (.A0(\spiking_network_top_uut.all_data_out[463] ),
    .A1(net4335),
    .S(_03369_),
    .X(_01968_));
 sg13g2_nor2_2 _18962_ (.A(_03231_),
    .B(net3723),
    .Y(_03370_));
 sg13g2_mux2_1 _18963_ (.A0(\spiking_network_top_uut.all_data_out[32] ),
    .A1(net4474),
    .S(_03370_),
    .X(_01969_));
 sg13g2_mux2_1 _18964_ (.A0(\spiking_network_top_uut.all_data_out[33] ),
    .A1(net4453),
    .S(_03370_),
    .X(_01970_));
 sg13g2_mux2_1 _18965_ (.A0(\spiking_network_top_uut.all_data_out[34] ),
    .A1(net4433),
    .S(_03370_),
    .X(_01971_));
 sg13g2_mux2_1 _18966_ (.A0(\spiking_network_top_uut.all_data_out[35] ),
    .A1(net4411),
    .S(_03370_),
    .X(_01972_));
 sg13g2_mux2_1 _18967_ (.A0(\spiking_network_top_uut.all_data_out[36] ),
    .A1(net4393),
    .S(_03370_),
    .X(_01973_));
 sg13g2_mux2_1 _18968_ (.A0(\spiking_network_top_uut.all_data_out[37] ),
    .A1(net4371),
    .S(_03370_),
    .X(_01974_));
 sg13g2_mux2_1 _18969_ (.A0(\spiking_network_top_uut.all_data_out[38] ),
    .A1(net4352),
    .S(_03370_),
    .X(_01975_));
 sg13g2_mux2_1 _18970_ (.A0(\spiking_network_top_uut.all_data_out[39] ),
    .A1(net4332),
    .S(_03370_),
    .X(_01976_));
 sg13g2_nor2_2 _18971_ (.A(_03258_),
    .B(net3727),
    .Y(_03371_));
 sg13g2_mux2_1 _18972_ (.A0(\spiking_network_top_uut.all_data_out[880] ),
    .A1(net4464),
    .S(net3672),
    .X(_01977_));
 sg13g2_mux2_1 _18973_ (.A0(\spiking_network_top_uut.all_data_out[881] ),
    .A1(net4443),
    .S(_03371_),
    .X(_01978_));
 sg13g2_nand2_1 _18974_ (.Y(_03372_),
    .A(net4424),
    .B(net3672));
 sg13g2_o21ai_1 _18975_ (.B1(_03372_),
    .Y(_01979_),
    .A1(_03577_),
    .A2(net3672));
 sg13g2_mux2_1 _18976_ (.A0(\spiking_network_top_uut.all_data_out[883] ),
    .A1(net4403),
    .S(net3672),
    .X(_01980_));
 sg13g2_mux2_1 _18977_ (.A0(\spiking_network_top_uut.all_data_out[884] ),
    .A1(net4380),
    .S(net3672),
    .X(_01981_));
 sg13g2_mux2_1 _18978_ (.A0(\spiking_network_top_uut.all_data_out[885] ),
    .A1(net4361),
    .S(net3672),
    .X(_01982_));
 sg13g2_mux2_1 _18979_ (.A0(\spiking_network_top_uut.all_data_out[886] ),
    .A1(net4339),
    .S(net3672),
    .X(_01983_));
 sg13g2_mux2_1 _18980_ (.A0(\spiking_network_top_uut.all_data_out[887] ),
    .A1(net4320),
    .S(net3672),
    .X(_01984_));
 sg13g2_nor2_2 _18981_ (.A(_03235_),
    .B(net3724),
    .Y(_03373_));
 sg13g2_mux2_1 _18982_ (.A0(\spiking_network_top_uut.all_data_out[24] ),
    .A1(net4464),
    .S(_03373_),
    .X(_01985_));
 sg13g2_mux2_1 _18983_ (.A0(\spiking_network_top_uut.all_data_out[25] ),
    .A1(net4443),
    .S(net3671),
    .X(_01986_));
 sg13g2_mux2_1 _18984_ (.A0(\spiking_network_top_uut.all_data_out[26] ),
    .A1(net4424),
    .S(net3671),
    .X(_01987_));
 sg13g2_mux2_1 _18985_ (.A0(\spiking_network_top_uut.all_data_out[27] ),
    .A1(net4405),
    .S(_03373_),
    .X(_01988_));
 sg13g2_nand2_1 _18986_ (.Y(_03374_),
    .A(net4384),
    .B(net3671));
 sg13g2_o21ai_1 _18987_ (.B1(_03374_),
    .Y(_01989_),
    .A1(_03394_),
    .A2(net3671));
 sg13g2_nand2_1 _18988_ (.Y(_03375_),
    .A(net4361),
    .B(net3671));
 sg13g2_o21ai_1 _18989_ (.B1(_03375_),
    .Y(_01990_),
    .A1(_03392_),
    .A2(net3671));
 sg13g2_mux2_1 _18990_ (.A0(\spiking_network_top_uut.all_data_out[30] ),
    .A1(net4342),
    .S(_03373_),
    .X(_01991_));
 sg13g2_nand2_1 _18991_ (.Y(_03376_),
    .A(net4321),
    .B(net3671));
 sg13g2_o21ai_1 _18992_ (.B1(_03376_),
    .Y(_01992_),
    .A1(_03390_),
    .A2(net3671));
 sg13g2_nor2_2 _18993_ (.A(net3734),
    .B(_03218_),
    .Y(_03377_));
 sg13g2_mux2_1 _18994_ (.A0(\spiking_network_top_uut.all_data_out[560] ),
    .A1(net4475),
    .S(_03377_),
    .X(_01993_));
 sg13g2_mux2_1 _18995_ (.A0(\spiking_network_top_uut.all_data_out[561] ),
    .A1(net4455),
    .S(_03377_),
    .X(_01994_));
 sg13g2_mux2_1 _18996_ (.A0(\spiking_network_top_uut.all_data_out[562] ),
    .A1(net4434),
    .S(_03377_),
    .X(_01995_));
 sg13g2_mux2_1 _18997_ (.A0(\spiking_network_top_uut.all_data_out[563] ),
    .A1(net4415),
    .S(_03377_),
    .X(_01996_));
 sg13g2_mux2_1 _18998_ (.A0(\spiking_network_top_uut.all_data_out[564] ),
    .A1(net4392),
    .S(_03377_),
    .X(_01997_));
 sg13g2_mux2_1 _18999_ (.A0(\spiking_network_top_uut.all_data_out[565] ),
    .A1(net4370),
    .S(_03377_),
    .X(_01998_));
 sg13g2_mux2_1 _19000_ (.A0(\spiking_network_top_uut.all_data_out[566] ),
    .A1(net4351),
    .S(_03377_),
    .X(_01999_));
 sg13g2_mux2_1 _19001_ (.A0(\spiking_network_top_uut.all_data_out[567] ),
    .A1(net4329),
    .S(_03377_),
    .X(_02000_));
 sg13g2_nor2_2 _19002_ (.A(_03241_),
    .B(_03345_),
    .Y(_03378_));
 sg13g2_mux2_1 _19003_ (.A0(\spiking_network_top_uut.all_data_out[16] ),
    .A1(net4463),
    .S(net3670),
    .X(_02001_));
 sg13g2_nand2_1 _19004_ (.Y(_03379_),
    .A(net4442),
    .B(net3670));
 sg13g2_o21ai_1 _19005_ (.B1(_03379_),
    .Y(_02002_),
    .A1(_03401_),
    .A2(net3670));
 sg13g2_mux2_1 _19006_ (.A0(net4305),
    .A1(net4423),
    .S(net3670),
    .X(_02003_));
 sg13g2_mux2_1 _19007_ (.A0(\spiking_network_top_uut.all_data_out[19] ),
    .A1(net4404),
    .S(net3670),
    .X(_02004_));
 sg13g2_mux2_1 _19008_ (.A0(net4292),
    .A1(net4381),
    .S(net3670),
    .X(_02005_));
 sg13g2_mux2_1 _19009_ (.A0(\spiking_network_top_uut.all_data_out[21] ),
    .A1(net4365),
    .S(net3670),
    .X(_02006_));
 sg13g2_mux2_1 _19010_ (.A0(\spiking_network_top_uut.all_data_out[22] ),
    .A1(net4352),
    .S(_03378_),
    .X(_02007_));
 sg13g2_mux2_1 _19011_ (.A0(\spiking_network_top_uut.all_data_out[23] ),
    .A1(net4320),
    .S(net3670),
    .X(_02008_));
 sg13g2_nor2_2 _19012_ (.A(_03256_),
    .B(net3727),
    .Y(_03380_));
 sg13g2_mux2_1 _19013_ (.A0(\spiking_network_top_uut.all_data_out[888] ),
    .A1(net4465),
    .S(_03380_),
    .X(_02009_));
 sg13g2_mux2_1 _19014_ (.A0(\spiking_network_top_uut.all_data_out[889] ),
    .A1(net4443),
    .S(_03380_),
    .X(_02010_));
 sg13g2_mux2_1 _19015_ (.A0(\spiking_network_top_uut.all_data_out[890] ),
    .A1(net4426),
    .S(_03380_),
    .X(_02011_));
 sg13g2_mux2_1 _19016_ (.A0(\spiking_network_top_uut.all_data_out[891] ),
    .A1(net4405),
    .S(_03380_),
    .X(_02012_));
 sg13g2_mux2_1 _19017_ (.A0(\spiking_network_top_uut.all_data_out[892] ),
    .A1(net4384),
    .S(_03380_),
    .X(_02013_));
 sg13g2_mux2_1 _19018_ (.A0(\spiking_network_top_uut.all_data_out[893] ),
    .A1(net4361),
    .S(_03380_),
    .X(_02014_));
 sg13g2_mux2_1 _19019_ (.A0(\spiking_network_top_uut.all_data_out[894] ),
    .A1(net4342),
    .S(_03380_),
    .X(_02015_));
 sg13g2_mux2_1 _19020_ (.A0(\spiking_network_top_uut.all_data_out[895] ),
    .A1(net4320),
    .S(_03380_),
    .X(_02016_));
 sg13g2_nor2_2 _19021_ (.A(_03245_),
    .B(net3723),
    .Y(_03381_));
 sg13g2_mux2_1 _19022_ (.A0(net4286),
    .A1(net4464),
    .S(_03381_),
    .X(_02017_));
 sg13g2_mux2_1 _19023_ (.A0(net4282),
    .A1(net4443),
    .S(_03381_),
    .X(_02018_));
 sg13g2_mux2_1 _19024_ (.A0(net4279),
    .A1(net4425),
    .S(_03381_),
    .X(_02019_));
 sg13g2_mux2_1 _19025_ (.A0(net4275),
    .A1(net4403),
    .S(_03381_),
    .X(_02020_));
 sg13g2_mux2_1 _19026_ (.A0(net4272),
    .A1(net4384),
    .S(_03381_),
    .X(_02021_));
 sg13g2_mux2_1 _19027_ (.A0(\spiking_network_top_uut.all_data_out[13] ),
    .A1(net4373),
    .S(_03381_),
    .X(_02022_));
 sg13g2_mux2_1 _19028_ (.A0(\spiking_network_top_uut.all_data_out[14] ),
    .A1(net4342),
    .S(_03381_),
    .X(_02023_));
 sg13g2_mux2_1 _19029_ (.A0(\spiking_network_top_uut.all_data_out[15] ),
    .A1(net4325),
    .S(_03381_),
    .X(_02024_));
 sg13g2_nor2_2 _19030_ (.A(net3736),
    .B(_03250_),
    .Y(_03382_));
 sg13g2_mux2_1 _19031_ (.A0(\spiking_network_top_uut.all_data_out[448] ),
    .A1(net4475),
    .S(net3669),
    .X(_02025_));
 sg13g2_mux2_1 _19032_ (.A0(\spiking_network_top_uut.all_data_out[449] ),
    .A1(net4455),
    .S(net3669),
    .X(_02026_));
 sg13g2_nand2_1 _19033_ (.Y(_03383_),
    .A(net4434),
    .B(net3669));
 sg13g2_o21ai_1 _19034_ (.B1(_03383_),
    .Y(_02027_),
    .A1(_03623_),
    .A2(net3669));
 sg13g2_mux2_1 _19035_ (.A0(\spiking_network_top_uut.all_data_out[451] ),
    .A1(net4419),
    .S(_03382_),
    .X(_02028_));
 sg13g2_mux2_1 _19036_ (.A0(\spiking_network_top_uut.all_data_out[452] ),
    .A1(net4395),
    .S(net3669),
    .X(_02029_));
 sg13g2_mux2_1 _19037_ (.A0(\spiking_network_top_uut.all_data_out[453] ),
    .A1(net4378),
    .S(net3669),
    .X(_02030_));
 sg13g2_mux2_1 _19038_ (.A0(\spiking_network_top_uut.all_data_out[454] ),
    .A1(net4354),
    .S(net3669),
    .X(_02031_));
 sg13g2_mux2_1 _19039_ (.A0(\spiking_network_top_uut.all_data_out[455] ),
    .A1(net4336),
    .S(net3669),
    .X(_02032_));
 sg13g2_nor2_2 _19040_ (.A(_03201_),
    .B(net3723),
    .Y(_03384_));
 sg13g2_mux2_1 _19041_ (.A0(net4268),
    .A1(net4469),
    .S(net3668),
    .X(_02033_));
 sg13g2_mux2_1 _19042_ (.A0(net4267),
    .A1(net4448),
    .S(net3668),
    .X(_02034_));
 sg13g2_nand2_1 _19043_ (.Y(_03385_),
    .A(net4429),
    .B(net3668));
 sg13g2_o21ai_1 _19044_ (.B1(_03385_),
    .Y(_02035_),
    .A1(_03473_),
    .A2(net3668));
 sg13g2_mux2_1 _19045_ (.A0(\spiking_network_top_uut.all_data_out[3] ),
    .A1(net4412),
    .S(_03384_),
    .X(_02036_));
 sg13g2_nand2_1 _19046_ (.Y(_03386_),
    .A(net4385),
    .B(net3668));
 sg13g2_o21ai_1 _19047_ (.B1(_03386_),
    .Y(_02037_),
    .A1(_03575_),
    .A2(net3668));
 sg13g2_mux2_1 _19048_ (.A0(\spiking_network_top_uut.all_data_out[5] ),
    .A1(net4367),
    .S(_03384_),
    .X(_02038_));
 sg13g2_mux2_1 _19049_ (.A0(\spiking_network_top_uut.all_data_out[6] ),
    .A1(net4344),
    .S(net3668),
    .X(_02039_));
 sg13g2_mux2_1 _19050_ (.A0(\spiking_network_top_uut.all_data_out[7] ),
    .A1(net4327),
    .S(net3668),
    .X(_02040_));
 sg13g2_mux2_1 _19051_ (.A0(net4265),
    .A1(net4484),
    .S(\spiking_network_top_uut.spi_inst.memory_inst.write_enable ),
    .X(_02041_));
 sg13g2_mux2_1 _19052_ (.A0(net4263),
    .A1(net4483),
    .S(net4317),
    .X(_02042_));
 sg13g2_nor2_1 _19053_ (.A(net4317),
    .B(\spiking_network_top_uut.spi_inst.memory_inst.addr_reg_out[2] ),
    .Y(_03387_));
 sg13g2_a21oi_1 _19054_ (.A1(_03405_),
    .A2(net4317),
    .Y(_02043_),
    .B1(_03387_));
 sg13g2_o21ai_1 _19055_ (.B1(_03212_),
    .Y(_02044_),
    .A1(net4317),
    .A2(_03508_));
 sg13g2_mux2_1 _19056_ (.A0(\spiking_network_top_uut.spi_inst.memory_inst.addr_reg_out[4] ),
    .A1(\spiking_network_top_uut.spi_inst.LSB_Address_reg[4] ),
    .S(net4317),
    .X(_02045_));
 sg13g2_mux2_1 _19057_ (.A0(\spiking_network_top_uut.spi_inst.memory_inst.addr_reg_out[5] ),
    .A1(\spiking_network_top_uut.spi_inst.LSB_Address_reg[5] ),
    .S(net4317),
    .X(_02046_));
 sg13g2_mux2_1 _19058_ (.A0(\spiking_network_top_uut.spi_inst.memory_inst.addr_reg_out[6] ),
    .A1(\spiking_network_top_uut.spi_inst.LSB_Address_reg[6] ),
    .S(\spiking_network_top_uut.spi_inst.memory_inst.write_enable ),
    .X(_02047_));
 sg13g2_nor2_2 _19059_ (.A(net3731),
    .B(_03231_),
    .Y(_03388_));
 sg13g2_mux2_1 _19060_ (.A0(\spiking_network_top_uut.all_data_out[672] ),
    .A1(net4468),
    .S(_03388_),
    .X(_02048_));
 sg13g2_mux2_1 _19061_ (.A0(\spiking_network_top_uut.all_data_out[673] ),
    .A1(net4445),
    .S(_03388_),
    .X(_02049_));
 sg13g2_mux2_1 _19062_ (.A0(\spiking_network_top_uut.all_data_out[674] ),
    .A1(net4426),
    .S(_03388_),
    .X(_02050_));
 sg13g2_mux2_1 _19063_ (.A0(\spiking_network_top_uut.all_data_out[675] ),
    .A1(net4405),
    .S(_03388_),
    .X(_02051_));
 sg13g2_mux2_1 _19064_ (.A0(\spiking_network_top_uut.all_data_out[676] ),
    .A1(net4383),
    .S(_03388_),
    .X(_02052_));
 sg13g2_mux2_1 _19065_ (.A0(\spiking_network_top_uut.all_data_out[677] ),
    .A1(net4362),
    .S(_03388_),
    .X(_02053_));
 sg13g2_mux2_1 _19066_ (.A0(\spiking_network_top_uut.all_data_out[678] ),
    .A1(net4341),
    .S(_03388_),
    .X(_02054_));
 sg13g2_mux2_1 _19067_ (.A0(\spiking_network_top_uut.all_data_out[679] ),
    .A1(net4322),
    .S(_03388_),
    .X(_02055_));
 sg13g2_mux2_1 _19068_ (.A0(\spiking_network_top_uut.debug_config_ready_reg_out ),
    .A1(\spiking_network_top_uut.spi_inst.debug_config_ready_reg_in ),
    .S(\spiking_network_top_uut.spi_inst.debug_config_ready_reg_en ),
    .X(_02056_));
 sg13g2_inv_1 _19069_ (.Y(_00422_),
    .A(net4704));
 sg13g2_inv_1 _19070_ (.Y(_00423_),
    .A(net4708));
 sg13g2_inv_1 _19071_ (.Y(_00424_),
    .A(net4704));
 sg13g2_dfrbp_1 _19072_ (.CLK(net4703),
    .RESET_B(net4023),
    .D(_00425_),
    .Q_N(_10326_),
    .Q(\spiking_network_top_uut.spi_inst.spi_slave_inst.shift_reg[0] ));
 sg13g2_dfrbp_1 _19073_ (.CLK(net4707),
    .RESET_B(net4027),
    .D(_00426_),
    .Q_N(_10325_),
    .Q(\spiking_network_top_uut.spi_inst.spi_slave_inst.shift_reg[1] ));
 sg13g2_dfrbp_1 _19074_ (.CLK(net4707),
    .RESET_B(net4027),
    .D(_00427_),
    .Q_N(_10324_),
    .Q(\spiking_network_top_uut.spi_inst.spi_slave_inst.shift_reg[2] ));
 sg13g2_dfrbp_1 _19075_ (.CLK(net4704),
    .RESET_B(net4025),
    .D(_00428_),
    .Q_N(_10323_),
    .Q(\spiking_network_top_uut.spi_inst.spi_slave_inst.shift_reg[3] ));
 sg13g2_dfrbp_1 _19076_ (.CLK(net4705),
    .RESET_B(net4025),
    .D(_00429_),
    .Q_N(_10322_),
    .Q(\spiking_network_top_uut.spi_inst.spi_slave_inst.shift_reg[4] ));
 sg13g2_dfrbp_1 _19077_ (.CLK(net4705),
    .RESET_B(net4024),
    .D(_00430_),
    .Q_N(_10321_),
    .Q(\spiking_network_top_uut.spi_inst.spi_slave_inst.shift_reg[5] ));
 sg13g2_dfrbp_1 _19078_ (.CLK(net4704),
    .RESET_B(net4024),
    .D(_00431_),
    .Q_N(_10327_),
    .Q(\spiking_network_top_uut.spi_inst.spi_slave_inst.shift_reg[6] ));
 sg13g2_dfrbp_1 _19079_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net4140),
    .D(net33),
    .Q_N(_10328_),
    .Q(\spiking_network_top_uut.debug_config_ready_sync ));
 sg13g2_dfrbp_1 _19080_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net4194),
    .D(net31),
    .Q_N(_10329_),
    .Q(\spiking_network_top_uut.clk_div_inst.enable ));
 sg13g2_dfrbp_1 _19081_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net4171),
    .D(net34),
    .Q_N(_10330_),
    .Q(\spiking_network_top_uut.SNN_en_sync ));
 sg13g2_dfrbp_1 _19082_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net4192),
    .D(net32),
    .Q_N(_10320_),
    .Q(\spiking_network_top_uut.input_ready_sync ));
 sg13g2_dfrbp_1 _19083_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net4184),
    .D(_00432_),
    .Q_N(_10319_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19084_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net4184),
    .D(_00433_),
    .Q_N(_10318_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19085_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net4194),
    .D(_00434_),
    .Q_N(_10317_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19086_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net4182),
    .D(_00435_),
    .Q_N(_10316_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19087_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net4180),
    .D(_00436_),
    .Q_N(_10315_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19088_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net4180),
    .D(_00437_),
    .Q_N(_10314_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19089_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net4184),
    .D(_00438_),
    .Q_N(_10313_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19090_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net4185),
    .D(net92),
    .Q_N(_10312_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19091_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net4163),
    .D(_00440_),
    .Q_N(_10311_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19092_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net4164),
    .D(_00441_),
    .Q_N(_10310_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19093_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net4166),
    .D(_00442_),
    .Q_N(_10309_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19094_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net4177),
    .D(_00443_),
    .Q_N(_10308_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19095_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net4167),
    .D(_00444_),
    .Q_N(_10307_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19096_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net4165),
    .D(_00445_),
    .Q_N(_10306_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19097_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net4177),
    .D(_00446_),
    .Q_N(_10305_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19098_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net4139),
    .D(net378),
    .Q_N(_00036_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[0] ));
 sg13g2_dfrbp_1 _19099_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net4139),
    .D(net352),
    .Q_N(_10304_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[1] ));
 sg13g2_dfrbp_1 _19100_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net4139),
    .D(_00449_),
    .Q_N(_10303_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[2] ));
 sg13g2_dfrbp_1 _19101_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net4139),
    .D(_00450_),
    .Q_N(_10302_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[3] ));
 sg13g2_dfrbp_1 _19102_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net4139),
    .D(_00451_),
    .Q_N(_10301_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[4] ));
 sg13g2_dfrbp_1 _19103_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net4164),
    .D(_00452_),
    .Q_N(_10300_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19104_ (.CLK(net4510),
    .RESET_B(net4210),
    .D(_00453_),
    .Q_N(_10331_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[7] ));
 sg13g2_dfrbp_1 _19105_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net4148),
    .D(_00017_),
    .Q_N(_10299_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.spike_out ));
 sg13g2_dfrbp_1 _19106_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net4147),
    .D(_00454_),
    .Q_N(_00034_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[0] ));
 sg13g2_dfrbp_1 _19107_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net4147),
    .D(_00455_),
    .Q_N(_00035_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ));
 sg13g2_dfrbp_1 _19108_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net4147),
    .D(_00456_),
    .Q_N(_00033_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ));
 sg13g2_dfrbp_1 _19109_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net4146),
    .D(_00457_),
    .Q_N(_00032_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ));
 sg13g2_dfrbp_1 _19110_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net4146),
    .D(_00458_),
    .Q_N(_00030_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ));
 sg13g2_dfrbp_1 _19111_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net4184),
    .D(_00459_),
    .Q_N(_10298_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[1].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19112_ (.CLK(net4503),
    .RESET_B(net4194),
    .D(_00460_),
    .Q_N(_10297_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[0] ));
 sg13g2_dfrbp_1 _19113_ (.CLK(net4503),
    .RESET_B(net4194),
    .D(_00461_),
    .Q_N(_10296_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[1] ));
 sg13g2_dfrbp_1 _19114_ (.CLK(net4503),
    .RESET_B(net4194),
    .D(_00462_),
    .Q_N(_10295_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[2] ));
 sg13g2_dfrbp_1 _19115_ (.CLK(net4503),
    .RESET_B(net4194),
    .D(_00463_),
    .Q_N(_10294_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[3] ));
 sg13g2_dfrbp_1 _19116_ (.CLK(net4503),
    .RESET_B(net4195),
    .D(_00464_),
    .Q_N(_10293_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[4] ));
 sg13g2_dfrbp_1 _19117_ (.CLK(net4503),
    .RESET_B(net4195),
    .D(_00465_),
    .Q_N(_10292_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[5] ));
 sg13g2_dfrbp_1 _19118_ (.CLK(net4503),
    .RESET_B(net4195),
    .D(_00466_),
    .Q_N(_10291_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[6] ));
 sg13g2_dfrbp_1 _19119_ (.CLK(net4503),
    .RESET_B(net4195),
    .D(_00467_),
    .Q_N(_10290_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[7] ));
 sg13g2_dfrbp_1 _19120_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net4184),
    .D(_00468_),
    .Q_N(_10289_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[1].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19121_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net4194),
    .D(_00469_),
    .Q_N(_10288_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[1].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19122_ (.CLK(net4499),
    .RESET_B(net4181),
    .D(_00470_),
    .Q_N(_10287_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[0] ));
 sg13g2_dfrbp_1 _19123_ (.CLK(net4498),
    .RESET_B(net4179),
    .D(_00471_),
    .Q_N(_10286_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[1] ));
 sg13g2_dfrbp_1 _19124_ (.CLK(net4497),
    .RESET_B(net4179),
    .D(_00472_),
    .Q_N(_10285_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[2] ));
 sg13g2_dfrbp_1 _19125_ (.CLK(net4498),
    .RESET_B(net4178),
    .D(_00473_),
    .Q_N(_10284_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[3] ));
 sg13g2_dfrbp_1 _19126_ (.CLK(net4498),
    .RESET_B(net4179),
    .D(_00474_),
    .Q_N(_10283_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[4] ));
 sg13g2_dfrbp_1 _19127_ (.CLK(net4495),
    .RESET_B(net4176),
    .D(_00475_),
    .Q_N(_10282_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[5] ));
 sg13g2_dfrbp_1 _19128_ (.CLK(net4495),
    .RESET_B(net4176),
    .D(_00476_),
    .Q_N(_10281_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[6] ));
 sg13g2_dfrbp_1 _19129_ (.CLK(net4496),
    .RESET_B(net4176),
    .D(_00477_),
    .Q_N(_10280_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[7] ));
 sg13g2_dfrbp_1 _19130_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net4194),
    .D(_00478_),
    .Q_N(_10279_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[1].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19131_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net4181),
    .D(_00479_),
    .Q_N(_10278_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[1].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19132_ (.CLK(net4499),
    .RESET_B(net4185),
    .D(_00480_),
    .Q_N(_10277_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[0] ));
 sg13g2_dfrbp_1 _19133_ (.CLK(net4502),
    .RESET_B(net4182),
    .D(_00481_),
    .Q_N(_10276_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[1] ));
 sg13g2_dfrbp_1 _19134_ (.CLK(net4502),
    .RESET_B(net4182),
    .D(_00482_),
    .Q_N(_10275_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[2] ));
 sg13g2_dfrbp_1 _19135_ (.CLK(net4502),
    .RESET_B(net4182),
    .D(_00483_),
    .Q_N(_10274_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[3] ));
 sg13g2_dfrbp_1 _19136_ (.CLK(net4502),
    .RESET_B(net4184),
    .D(_00484_),
    .Q_N(_10273_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[4] ));
 sg13g2_dfrbp_1 _19137_ (.CLK(net4502),
    .RESET_B(net4182),
    .D(_00485_),
    .Q_N(_10272_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[5] ));
 sg13g2_dfrbp_1 _19138_ (.CLK(net4502),
    .RESET_B(net4182),
    .D(_00486_),
    .Q_N(_10271_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[6] ));
 sg13g2_dfrbp_1 _19139_ (.CLK(net4502),
    .RESET_B(net4182),
    .D(_00487_),
    .Q_N(_10270_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[7] ));
 sg13g2_dfrbp_1 _19140_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net4180),
    .D(_00488_),
    .Q_N(_10269_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[1].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19141_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net4185),
    .D(_00489_),
    .Q_N(_10268_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[1].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19142_ (.CLK(net4493),
    .RESET_B(net4145),
    .D(_00490_),
    .Q_N(_10267_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[0] ));
 sg13g2_dfrbp_1 _19143_ (.CLK(net4493),
    .RESET_B(net4145),
    .D(_00491_),
    .Q_N(_10266_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[1] ));
 sg13g2_dfrbp_1 _19144_ (.CLK(net4493),
    .RESET_B(net4145),
    .D(_00492_),
    .Q_N(_10265_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[2] ));
 sg13g2_dfrbp_1 _19145_ (.CLK(net4493),
    .RESET_B(net4145),
    .D(_00493_),
    .Q_N(_10264_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[3] ));
 sg13g2_dfrbp_1 _19146_ (.CLK(net4493),
    .RESET_B(net4145),
    .D(_00494_),
    .Q_N(_10263_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[4] ));
 sg13g2_dfrbp_1 _19147_ (.CLK(net4493),
    .RESET_B(net4163),
    .D(_00495_),
    .Q_N(_10262_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[5] ));
 sg13g2_dfrbp_1 _19148_ (.CLK(net4493),
    .RESET_B(net4163),
    .D(_00496_),
    .Q_N(_10261_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[6] ));
 sg13g2_dfrbp_1 _19149_ (.CLK(net4493),
    .RESET_B(net4163),
    .D(_00497_),
    .Q_N(_10260_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[7] ));
 sg13g2_dfrbp_1 _19150_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net4185),
    .D(_00498_),
    .Q_N(_10259_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[1].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19151_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net4163),
    .D(_00499_),
    .Q_N(_10258_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[1].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19152_ (.CLK(net4495),
    .RESET_B(net4166),
    .D(_00500_),
    .Q_N(_10257_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[0] ));
 sg13g2_dfrbp_1 _19153_ (.CLK(net4495),
    .RESET_B(net4166),
    .D(_00501_),
    .Q_N(_10256_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[1] ));
 sg13g2_dfrbp_1 _19154_ (.CLK(net4495),
    .RESET_B(net4166),
    .D(_00502_),
    .Q_N(_10255_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[2] ));
 sg13g2_dfrbp_1 _19155_ (.CLK(net4495),
    .RESET_B(net4166),
    .D(_00503_),
    .Q_N(_10254_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[3] ));
 sg13g2_dfrbp_1 _19156_ (.CLK(net4496),
    .RESET_B(net4176),
    .D(_00504_),
    .Q_N(_10253_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[4] ));
 sg13g2_dfrbp_1 _19157_ (.CLK(net4496),
    .RESET_B(net4176),
    .D(_00505_),
    .Q_N(_10252_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[5] ));
 sg13g2_dfrbp_1 _19158_ (.CLK(net4496),
    .RESET_B(net4176),
    .D(_00506_),
    .Q_N(_10251_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[6] ));
 sg13g2_dfrbp_1 _19159_ (.CLK(net4496),
    .RESET_B(net4176),
    .D(_00507_),
    .Q_N(_10250_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[7] ));
 sg13g2_dfrbp_1 _19160_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net4163),
    .D(_00508_),
    .Q_N(_10249_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[1].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19161_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net4176),
    .D(_00509_),
    .Q_N(_10248_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[1].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19162_ (.CLK(net4494),
    .RESET_B(net4165),
    .D(_00510_),
    .Q_N(_10247_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[0] ));
 sg13g2_dfrbp_1 _19163_ (.CLK(net4494),
    .RESET_B(net4165),
    .D(_00511_),
    .Q_N(_10246_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[1] ));
 sg13g2_dfrbp_1 _19164_ (.CLK(net4494),
    .RESET_B(net4165),
    .D(_00512_),
    .Q_N(_10245_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[2] ));
 sg13g2_dfrbp_1 _19165_ (.CLK(net4494),
    .RESET_B(net4165),
    .D(_00513_),
    .Q_N(_10244_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[3] ));
 sg13g2_dfrbp_1 _19166_ (.CLK(net4494),
    .RESET_B(net4165),
    .D(_00514_),
    .Q_N(_10243_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[4] ));
 sg13g2_dfrbp_1 _19167_ (.CLK(net4494),
    .RESET_B(net4166),
    .D(_00515_),
    .Q_N(_10242_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[5] ));
 sg13g2_dfrbp_1 _19168_ (.CLK(net4495),
    .RESET_B(net4166),
    .D(_00516_),
    .Q_N(_10241_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[6] ));
 sg13g2_dfrbp_1 _19169_ (.CLK(net4495),
    .RESET_B(net4166),
    .D(_00517_),
    .Q_N(_10240_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[7] ));
 sg13g2_dfrbp_1 _19170_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net4177),
    .D(_00518_),
    .Q_N(_10239_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[1].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19171_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net4167),
    .D(_00519_),
    .Q_N(_10238_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[1].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19172_ (.CLK(net4494),
    .RESET_B(net4165),
    .D(_00520_),
    .Q_N(_10237_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[0] ));
 sg13g2_dfrbp_1 _19173_ (.CLK(net4497),
    .RESET_B(net4178),
    .D(_00521_),
    .Q_N(_10236_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[1] ));
 sg13g2_dfrbp_1 _19174_ (.CLK(net4497),
    .RESET_B(net4178),
    .D(_00522_),
    .Q_N(_10235_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[2] ));
 sg13g2_dfrbp_1 _19175_ (.CLK(net4497),
    .RESET_B(net4178),
    .D(_00523_),
    .Q_N(_10234_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[3] ));
 sg13g2_dfrbp_1 _19176_ (.CLK(net4497),
    .RESET_B(net4178),
    .D(_00524_),
    .Q_N(_10233_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[4] ));
 sg13g2_dfrbp_1 _19177_ (.CLK(net4497),
    .RESET_B(net4178),
    .D(_00525_),
    .Q_N(_10232_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[5] ));
 sg13g2_dfrbp_1 _19178_ (.CLK(net4497),
    .RESET_B(net4178),
    .D(_00526_),
    .Q_N(_10231_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[6] ));
 sg13g2_dfrbp_1 _19179_ (.CLK(net4497),
    .RESET_B(net4178),
    .D(_00527_),
    .Q_N(_10230_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[7] ));
 sg13g2_dfrbp_1 _19180_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net4167),
    .D(_00528_),
    .Q_N(_10229_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[1].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19181_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net4177),
    .D(_00529_),
    .Q_N(_10228_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[1].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19182_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net4137),
    .D(net338),
    .Q_N(_00042_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[0] ));
 sg13g2_dfrbp_1 _19183_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net4137),
    .D(net410),
    .Q_N(_10227_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[1] ));
 sg13g2_dfrbp_1 _19184_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net4137),
    .D(_00532_),
    .Q_N(_10226_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[2] ));
 sg13g2_dfrbp_1 _19185_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net4137),
    .D(_00533_),
    .Q_N(_10225_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[3] ));
 sg13g2_dfrbp_1 _19186_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net4139),
    .D(_00534_),
    .Q_N(_10224_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[4] ));
 sg13g2_dfrbp_1 _19187_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net4165),
    .D(_00535_),
    .Q_N(_10332_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[1].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19188_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net4148),
    .D(_00018_),
    .Q_N(_10223_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.spike_out ));
 sg13g2_dfrbp_1 _19189_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net4142),
    .D(_00536_),
    .Q_N(_00040_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[0] ));
 sg13g2_dfrbp_1 _19190_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net4142),
    .D(_00537_),
    .Q_N(_00041_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ));
 sg13g2_dfrbp_1 _19191_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net4142),
    .D(_00538_),
    .Q_N(_00039_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ));
 sg13g2_dfrbp_1 _19192_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net4142),
    .D(_00539_),
    .Q_N(_00038_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ));
 sg13g2_dfrbp_1 _19193_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net4142),
    .D(_00540_),
    .Q_N(_00037_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ));
 sg13g2_dfrbp_1 _19194_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net4207),
    .D(_00541_),
    .Q_N(_10222_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19195_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net4207),
    .D(_00542_),
    .Q_N(_10221_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19196_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net4205),
    .D(_00543_),
    .Q_N(_10220_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19197_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net4199),
    .D(_00544_),
    .Q_N(_10219_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19198_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net4220),
    .D(_00545_),
    .Q_N(_10218_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19199_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net4219),
    .D(_00546_),
    .Q_N(_10217_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19200_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net4213),
    .D(_00547_),
    .Q_N(_10216_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19201_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net4213),
    .D(_00548_),
    .Q_N(_10215_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19202_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net4233),
    .D(_00549_),
    .Q_N(_10214_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19203_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net4232),
    .D(_00550_),
    .Q_N(_10213_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19204_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net4224),
    .D(_00551_),
    .Q_N(_10212_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19205_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net4226),
    .D(_00552_),
    .Q_N(_10211_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19206_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net4201),
    .D(_00553_),
    .Q_N(_10210_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19207_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net4201),
    .D(_00554_),
    .Q_N(_10209_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19208_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net4198),
    .D(_00555_),
    .Q_N(_10208_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19209_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net4140),
    .D(net376),
    .Q_N(_00048_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[0] ));
 sg13g2_dfrbp_1 _19210_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net4139),
    .D(_00557_),
    .Q_N(_10207_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[1] ));
 sg13g2_dfrbp_1 _19211_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net4139),
    .D(net154),
    .Q_N(_10206_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[2] ));
 sg13g2_dfrbp_1 _19212_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net4140),
    .D(_00559_),
    .Q_N(_10205_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[3] ));
 sg13g2_dfrbp_1 _19213_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net4140),
    .D(_00560_),
    .Q_N(_10204_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[4] ));
 sg13g2_dfrbp_1 _19214_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net4198),
    .D(_00561_),
    .Q_N(_10203_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19215_ (.CLK(net4523),
    .RESET_B(net4254),
    .D(_00562_),
    .Q_N(_10333_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[7] ));
 sg13g2_dfrbp_1 _19216_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net4163),
    .D(_00009_),
    .Q_N(_10202_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.spike_out ));
 sg13g2_dfrbp_1 _19217_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net4164),
    .D(_00563_),
    .Q_N(_00046_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[0] ));
 sg13g2_dfrbp_1 _19218_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net4164),
    .D(_00564_),
    .Q_N(_00047_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ));
 sg13g2_dfrbp_1 _19219_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net4164),
    .D(_00565_),
    .Q_N(_00045_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ));
 sg13g2_dfrbp_1 _19220_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net4164),
    .D(_00566_),
    .Q_N(_00044_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ));
 sg13g2_dfrbp_1 _19221_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net4164),
    .D(_00567_),
    .Q_N(_00043_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ));
 sg13g2_dfrbp_1 _19222_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net4210),
    .D(_00568_),
    .Q_N(_10201_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19223_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net4199),
    .D(net481),
    .Q_N(_10200_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19224_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net4199),
    .D(_00570_),
    .Q_N(_10199_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19225_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net4199),
    .D(_00571_),
    .Q_N(_10198_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19226_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net4220),
    .D(_00572_),
    .Q_N(_10197_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19227_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net4211),
    .D(_00573_),
    .Q_N(_10196_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19228_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net4221),
    .D(_00574_),
    .Q_N(_10195_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19229_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net4221),
    .D(_00575_),
    .Q_N(_10194_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19230_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net4227),
    .D(_00576_),
    .Q_N(_10193_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19231_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net4226),
    .D(_00577_),
    .Q_N(_10192_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19232_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net4239),
    .D(_00578_),
    .Q_N(_10191_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19233_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net4239),
    .D(_00579_),
    .Q_N(_10190_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19234_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net4201),
    .D(_00580_),
    .Q_N(_10189_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19235_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net4201),
    .D(_00581_),
    .Q_N(_10188_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19236_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net4200),
    .D(_00582_),
    .Q_N(_10187_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19237_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net4138),
    .D(net332),
    .Q_N(_00054_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[0] ));
 sg13g2_dfrbp_1 _19238_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net4138),
    .D(_00584_),
    .Q_N(_10186_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[1] ));
 sg13g2_dfrbp_1 _19239_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net4138),
    .D(_00585_),
    .Q_N(_10185_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[2] ));
 sg13g2_dfrbp_1 _19240_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net4138),
    .D(_00586_),
    .Q_N(_10184_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[3] ));
 sg13g2_dfrbp_1 _19241_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net4141),
    .D(_00587_),
    .Q_N(_10183_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[4] ));
 sg13g2_dfrbp_1 _19242_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net4196),
    .D(_00588_),
    .Q_N(_10334_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19243_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net4148),
    .D(_00010_),
    .Q_N(_10182_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.spike_out ));
 sg13g2_dfrbp_1 _19244_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net4148),
    .D(_00589_),
    .Q_N(_00052_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[0] ));
 sg13g2_dfrbp_1 _19245_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net4148),
    .D(_00590_),
    .Q_N(_00053_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ));
 sg13g2_dfrbp_1 _19246_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net4147),
    .D(_00591_),
    .Q_N(_00051_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ));
 sg13g2_dfrbp_1 _19247_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net4147),
    .D(_00592_),
    .Q_N(_00050_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ));
 sg13g2_dfrbp_1 _19248_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net4147),
    .D(_00593_),
    .Q_N(_00049_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ));
 sg13g2_dfrbp_1 _19249_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net4206),
    .D(_00594_),
    .Q_N(_10181_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19250_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net4206),
    .D(_00595_),
    .Q_N(_10180_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19251_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net4205),
    .D(_00596_),
    .Q_N(_10179_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19252_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net4206),
    .D(_00597_),
    .Q_N(_10178_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19253_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net4222),
    .D(_00598_),
    .Q_N(_10177_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19254_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net4222),
    .D(_00599_),
    .Q_N(_10176_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19255_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net4212),
    .D(_00600_),
    .Q_N(_10175_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19256_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net4214),
    .D(_00601_),
    .Q_N(_10174_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19257_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net4228),
    .D(_00602_),
    .Q_N(_10173_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19258_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net4231),
    .D(_00603_),
    .Q_N(_10172_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19259_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net4225),
    .D(_00604_),
    .Q_N(_10171_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19260_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net4226),
    .D(_00605_),
    .Q_N(_10170_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19261_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net4187),
    .D(_00606_),
    .Q_N(_10169_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19262_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net4187),
    .D(_00607_),
    .Q_N(_10168_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19263_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net4180),
    .D(_00608_),
    .Q_N(_10167_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19264_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net4137),
    .D(net317),
    .Q_N(_00060_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[0] ));
 sg13g2_dfrbp_1 _19265_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net4137),
    .D(net415),
    .Q_N(_10166_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[1] ));
 sg13g2_dfrbp_1 _19266_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net4137),
    .D(_00611_),
    .Q_N(_10165_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[2] ));
 sg13g2_dfrbp_1 _19267_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net4138),
    .D(_00612_),
    .Q_N(_10164_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[3] ));
 sg13g2_dfrbp_1 _19268_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net4137),
    .D(_00613_),
    .Q_N(_10163_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[4] ));
 sg13g2_dfrbp_1 _19269_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net4180),
    .D(_00614_),
    .Q_N(_10335_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19270_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net4169),
    .D(_00011_),
    .Q_N(_10162_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.spike_out ));
 sg13g2_dfrbp_1 _19271_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net4168),
    .D(_00615_),
    .Q_N(_00058_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[0] ));
 sg13g2_dfrbp_1 _19272_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net4168),
    .D(_00616_),
    .Q_N(_00059_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ));
 sg13g2_dfrbp_1 _19273_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net4159),
    .D(_00617_),
    .Q_N(_00057_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ));
 sg13g2_dfrbp_1 _19274_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net4168),
    .D(_00618_),
    .Q_N(_00056_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ));
 sg13g2_dfrbp_1 _19275_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net4168),
    .D(_00619_),
    .Q_N(_00055_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ));
 sg13g2_dfrbp_1 _19276_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net4210),
    .D(_00620_),
    .Q_N(_10161_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19277_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net4207),
    .D(net350),
    .Q_N(_10160_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19278_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net4204),
    .D(_00622_),
    .Q_N(_10159_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19279_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net4208),
    .D(net63),
    .Q_N(_10158_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19280_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net4223),
    .D(_00624_),
    .Q_N(_10157_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19281_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net4223),
    .D(_00625_),
    .Q_N(_10156_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19282_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net4213),
    .D(_00626_),
    .Q_N(_10155_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19283_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net4214),
    .D(_00627_),
    .Q_N(_10154_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19284_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net4228),
    .D(_00628_),
    .Q_N(_10153_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19285_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net4228),
    .D(net37),
    .Q_N(_10152_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19286_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net4225),
    .D(_00630_),
    .Q_N(_10151_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19287_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net4226),
    .D(_00631_),
    .Q_N(_10150_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19288_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net4191),
    .D(_00632_),
    .Q_N(_10149_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19289_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net4201),
    .D(_00633_),
    .Q_N(_10148_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19290_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net4196),
    .D(_00634_),
    .Q_N(_10147_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19291_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net4141),
    .D(net334),
    .Q_N(_00066_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[0] ));
 sg13g2_dfrbp_1 _19292_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net4141),
    .D(net344),
    .Q_N(_10146_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[1] ));
 sg13g2_dfrbp_1 _19293_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net4141),
    .D(net209),
    .Q_N(_10145_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[2] ));
 sg13g2_dfrbp_1 _19294_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net4141),
    .D(_00638_),
    .Q_N(_10144_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[3] ));
 sg13g2_dfrbp_1 _19295_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net4141),
    .D(_00639_),
    .Q_N(_10143_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[4] ));
 sg13g2_dfrbp_1 _19296_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net4196),
    .D(_00640_),
    .Q_N(_10336_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19297_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net4148),
    .D(_00012_),
    .Q_N(_10142_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.spike_out ));
 sg13g2_dfrbp_1 _19298_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net4152),
    .D(_00641_),
    .Q_N(_00064_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[0] ));
 sg13g2_dfrbp_1 _19299_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net4152),
    .D(_00642_),
    .Q_N(_00065_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ));
 sg13g2_dfrbp_1 _19300_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net4150),
    .D(_00643_),
    .Q_N(_00063_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ));
 sg13g2_dfrbp_1 _19301_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net4150),
    .D(_00644_),
    .Q_N(_00062_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ));
 sg13g2_dfrbp_1 _19302_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net4150),
    .D(_00645_),
    .Q_N(_00061_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ));
 sg13g2_dfrbp_1 _19303_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net4207),
    .D(_00646_),
    .Q_N(_10141_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19304_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net4208),
    .D(_00647_),
    .Q_N(_10140_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19305_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net4205),
    .D(_00648_),
    .Q_N(_10139_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19306_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net4206),
    .D(_00649_),
    .Q_N(_10138_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19307_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net4222),
    .D(_00650_),
    .Q_N(_10137_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19308_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net4222),
    .D(_00651_),
    .Q_N(_10136_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19309_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net4211),
    .D(_00652_),
    .Q_N(_10135_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19310_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net4213),
    .D(_00653_),
    .Q_N(_10134_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19311_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net4231),
    .D(_00654_),
    .Q_N(_10133_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19312_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net4231),
    .D(_00655_),
    .Q_N(_10132_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19313_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net4226),
    .D(_00656_),
    .Q_N(_10131_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19314_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net4241),
    .D(_00657_),
    .Q_N(_10130_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19315_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net4201),
    .D(_00658_),
    .Q_N(_10129_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19316_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net4201),
    .D(_00659_),
    .Q_N(_10128_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19317_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net4196),
    .D(_00660_),
    .Q_N(_10127_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19318_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net4156),
    .D(net347),
    .Q_N(_00072_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[0] ));
 sg13g2_dfrbp_1 _19319_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net4156),
    .D(net420),
    .Q_N(_10126_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[1] ));
 sg13g2_dfrbp_1 _19320_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net4156),
    .D(_00663_),
    .Q_N(_10125_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[2] ));
 sg13g2_dfrbp_1 _19321_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net4156),
    .D(_00664_),
    .Q_N(_10124_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[3] ));
 sg13g2_dfrbp_1 _19322_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net4157),
    .D(_00665_),
    .Q_N(_10123_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[4] ));
 sg13g2_dfrbp_1 _19323_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net4201),
    .D(net167),
    .Q_N(_10337_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19324_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net4158),
    .D(_00013_),
    .Q_N(_10122_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.spike_out ));
 sg13g2_dfrbp_1 _19325_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net4158),
    .D(_00667_),
    .Q_N(_00070_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[0] ));
 sg13g2_dfrbp_1 _19326_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net4158),
    .D(_00668_),
    .Q_N(_00071_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ));
 sg13g2_dfrbp_1 _19327_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net4160),
    .D(_00669_),
    .Q_N(_00069_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ));
 sg13g2_dfrbp_1 _19328_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net4158),
    .D(_00670_),
    .Q_N(_00068_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ));
 sg13g2_dfrbp_1 _19329_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net4158),
    .D(_00671_),
    .Q_N(_00067_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ));
 sg13g2_dfrbp_1 _19330_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net4208),
    .D(_00672_),
    .Q_N(_10121_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19331_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net4206),
    .D(_00673_),
    .Q_N(_10120_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19332_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net4199),
    .D(_00674_),
    .Q_N(_10119_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19333_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net4198),
    .D(_00675_),
    .Q_N(_10118_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19334_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net4222),
    .D(_00676_),
    .Q_N(_10117_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19335_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net4222),
    .D(_00677_),
    .Q_N(_10116_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19336_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net4212),
    .D(_00678_),
    .Q_N(_10115_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19337_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net4212),
    .D(_00679_),
    .Q_N(_10114_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19338_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net4228),
    .D(_00680_),
    .Q_N(_10113_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19339_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net4228),
    .D(_00681_),
    .Q_N(_10112_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19340_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net4227),
    .D(_00682_),
    .Q_N(_10111_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19341_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net4226),
    .D(net384),
    .Q_N(_10110_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19342_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net4191),
    .D(_00684_),
    .Q_N(_10109_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19343_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net4191),
    .D(_00685_),
    .Q_N(_10108_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19344_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net4200),
    .D(_00686_),
    .Q_N(_10107_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19345_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net4154),
    .D(net354),
    .Q_N(_00078_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[0] ));
 sg13g2_dfrbp_1 _19346_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net4154),
    .D(net324),
    .Q_N(_10106_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[1] ));
 sg13g2_dfrbp_1 _19347_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net4154),
    .D(_00689_),
    .Q_N(_10105_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[2] ));
 sg13g2_dfrbp_1 _19348_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net4155),
    .D(_00690_),
    .Q_N(_10104_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[3] ));
 sg13g2_dfrbp_1 _19349_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net4156),
    .D(_00691_),
    .Q_N(_10103_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[4] ));
 sg13g2_dfrbp_1 _19350_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net4185),
    .D(net292),
    .Q_N(_10338_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19351_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net4159),
    .D(_00014_),
    .Q_N(_10102_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.spike_out ));
 sg13g2_dfrbp_1 _19352_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net4159),
    .D(_00693_),
    .Q_N(_00076_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[0] ));
 sg13g2_dfrbp_1 _19353_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net4160),
    .D(_00694_),
    .Q_N(_00077_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ));
 sg13g2_dfrbp_1 _19354_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net4160),
    .D(_00695_),
    .Q_N(_00075_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ));
 sg13g2_dfrbp_1 _19355_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net4161),
    .D(_00696_),
    .Q_N(_00074_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ));
 sg13g2_dfrbp_1 _19356_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net4159),
    .D(_00697_),
    .Q_N(_00073_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ));
 sg13g2_dfrbp_1 _19357_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net4214),
    .D(_00698_),
    .Q_N(_10101_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19358_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net4210),
    .D(net59),
    .Q_N(_10100_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19359_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net4204),
    .D(_00700_),
    .Q_N(_10099_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19360_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net4208),
    .D(_00701_),
    .Q_N(_10098_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19361_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net4219),
    .D(_00702_),
    .Q_N(_10097_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19362_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net4220),
    .D(_00703_),
    .Q_N(_10096_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19363_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net4211),
    .D(_00704_),
    .Q_N(_10095_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19364_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net4211),
    .D(_00705_),
    .Q_N(_10094_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19365_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net4223),
    .D(_00706_),
    .Q_N(_10093_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19366_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net4223),
    .D(_00707_),
    .Q_N(_10092_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19367_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net4224),
    .D(_00708_),
    .Q_N(_10091_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19368_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net4225),
    .D(_00709_),
    .Q_N(_10090_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19369_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net4190),
    .D(_00710_),
    .Q_N(_10089_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19370_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net4180),
    .D(_00711_),
    .Q_N(_10088_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19371_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net4187),
    .D(_00712_),
    .Q_N(_10087_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19372_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net4146),
    .D(net321),
    .Q_N(_00084_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[0] ));
 sg13g2_dfrbp_1 _19373_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net4146),
    .D(_00714_),
    .Q_N(_10086_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[1] ));
 sg13g2_dfrbp_1 _19374_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net4146),
    .D(net214),
    .Q_N(_10085_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[2] ));
 sg13g2_dfrbp_1 _19375_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net4146),
    .D(_00716_),
    .Q_N(_10084_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[3] ));
 sg13g2_dfrbp_1 _19376_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net4146),
    .D(_00717_),
    .Q_N(_10083_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[4] ));
 sg13g2_dfrbp_1 _19377_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net4187),
    .D(_00718_),
    .Q_N(_10339_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19378_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net4163),
    .D(_00015_),
    .Q_N(_10082_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.spike_out ));
 sg13g2_dfrbp_1 _19379_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net4148),
    .D(_00719_),
    .Q_N(_00082_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[0] ));
 sg13g2_dfrbp_1 _19380_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net4149),
    .D(_00720_),
    .Q_N(_00083_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ));
 sg13g2_dfrbp_1 _19381_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net4145),
    .D(_00721_),
    .Q_N(_00081_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ));
 sg13g2_dfrbp_1 _19382_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net4145),
    .D(_00722_),
    .Q_N(_00080_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ));
 sg13g2_dfrbp_1 _19383_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net4149),
    .D(_00723_),
    .Q_N(_00079_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ));
 sg13g2_dfrbp_1 _19384_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net4207),
    .D(_00724_),
    .Q_N(_10081_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19385_ (.CLK(net4506),
    .RESET_B(net4205),
    .D(_00725_),
    .Q_N(_10080_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[0] ));
 sg13g2_dfrbp_1 _19386_ (.CLK(net4507),
    .RESET_B(net4205),
    .D(_00726_),
    .Q_N(_10079_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[1] ));
 sg13g2_dfrbp_1 _19387_ (.CLK(net4507),
    .RESET_B(net4204),
    .D(_00727_),
    .Q_N(_10078_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[2] ));
 sg13g2_dfrbp_1 _19388_ (.CLK(net4507),
    .RESET_B(net4204),
    .D(_00728_),
    .Q_N(_10077_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[3] ));
 sg13g2_dfrbp_1 _19389_ (.CLK(net4507),
    .RESET_B(net4204),
    .D(_00729_),
    .Q_N(_10076_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[4] ));
 sg13g2_dfrbp_1 _19390_ (.CLK(net4506),
    .RESET_B(net4205),
    .D(_00730_),
    .Q_N(_10075_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[5] ));
 sg13g2_dfrbp_1 _19391_ (.CLK(net4506),
    .RESET_B(net4205),
    .D(_00731_),
    .Q_N(_10074_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[6] ));
 sg13g2_dfrbp_1 _19392_ (.CLK(net4506),
    .RESET_B(net4204),
    .D(_00732_),
    .Q_N(_10073_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[7] ));
 sg13g2_dfrbp_1 _19393_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net4208),
    .D(_00733_),
    .Q_N(_10072_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19394_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net4204),
    .D(_00734_),
    .Q_N(_10071_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19395_ (.CLK(net4513),
    .RESET_B(net4222),
    .D(_00735_),
    .Q_N(_10070_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[0] ));
 sg13g2_dfrbp_1 _19396_ (.CLK(net4514),
    .RESET_B(net4219),
    .D(_00736_),
    .Q_N(_10069_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[1] ));
 sg13g2_dfrbp_1 _19397_ (.CLK(net4514),
    .RESET_B(net4219),
    .D(_00737_),
    .Q_N(_10068_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[2] ));
 sg13g2_dfrbp_1 _19398_ (.CLK(net4514),
    .RESET_B(net4219),
    .D(_00738_),
    .Q_N(_10067_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[3] ));
 sg13g2_dfrbp_1 _19399_ (.CLK(net4514),
    .RESET_B(net4219),
    .D(_00739_),
    .Q_N(_10066_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[4] ));
 sg13g2_dfrbp_1 _19400_ (.CLK(net4514),
    .RESET_B(net4220),
    .D(_00740_),
    .Q_N(_10065_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[5] ));
 sg13g2_dfrbp_1 _19401_ (.CLK(net4514),
    .RESET_B(net4219),
    .D(_00741_),
    .Q_N(_10064_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[6] ));
 sg13g2_dfrbp_1 _19402_ (.CLK(net4514),
    .RESET_B(net4219),
    .D(_00742_),
    .Q_N(_10063_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[7] ));
 sg13g2_dfrbp_1 _19403_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net4204),
    .D(_00743_),
    .Q_N(_10062_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19404_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net4223),
    .D(_00744_),
    .Q_N(_10061_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19405_ (.CLK(net4511),
    .RESET_B(net4212),
    .D(_00745_),
    .Q_N(_10060_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[0] ));
 sg13g2_dfrbp_1 _19406_ (.CLK(net4511),
    .RESET_B(net4211),
    .D(_00746_),
    .Q_N(_10059_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[1] ));
 sg13g2_dfrbp_1 _19407_ (.CLK(net4511),
    .RESET_B(net4211),
    .D(_00747_),
    .Q_N(_10058_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[2] ));
 sg13g2_dfrbp_1 _19408_ (.CLK(net4511),
    .RESET_B(net4211),
    .D(_00748_),
    .Q_N(_10057_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[3] ));
 sg13g2_dfrbp_1 _19409_ (.CLK(net4511),
    .RESET_B(net4211),
    .D(_00749_),
    .Q_N(_10056_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[4] ));
 sg13g2_dfrbp_1 _19410_ (.CLK(net4511),
    .RESET_B(net4221),
    .D(_00750_),
    .Q_N(_10055_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[5] ));
 sg13g2_dfrbp_1 _19411_ (.CLK(net4511),
    .RESET_B(net4221),
    .D(_00751_),
    .Q_N(_10054_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[6] ));
 sg13g2_dfrbp_1 _19412_ (.CLK(net4511),
    .RESET_B(net4221),
    .D(_00752_),
    .Q_N(_10053_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[7] ));
 sg13g2_dfrbp_1 _19413_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net4222),
    .D(_00753_),
    .Q_N(_10052_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19414_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net4213),
    .D(_00754_),
    .Q_N(_10051_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19415_ (.CLK(net4513),
    .RESET_B(net4228),
    .D(_00755_),
    .Q_N(_10050_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[0] ));
 sg13g2_dfrbp_1 _19416_ (.CLK(net4516),
    .RESET_B(net4232),
    .D(_00756_),
    .Q_N(_10049_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[1] ));
 sg13g2_dfrbp_1 _19417_ (.CLK(net4516),
    .RESET_B(net4232),
    .D(_00757_),
    .Q_N(_10048_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[2] ));
 sg13g2_dfrbp_1 _19418_ (.CLK(net4516),
    .RESET_B(net4232),
    .D(_00758_),
    .Q_N(_10047_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[3] ));
 sg13g2_dfrbp_1 _19419_ (.CLK(net4516),
    .RESET_B(net4232),
    .D(_00759_),
    .Q_N(_10046_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[4] ));
 sg13g2_dfrbp_1 _19420_ (.CLK(net4517),
    .RESET_B(net4232),
    .D(_00760_),
    .Q_N(_10045_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[5] ));
 sg13g2_dfrbp_1 _19421_ (.CLK(net4517),
    .RESET_B(net4232),
    .D(_00761_),
    .Q_N(_10044_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[6] ));
 sg13g2_dfrbp_1 _19422_ (.CLK(net4517),
    .RESET_B(net4232),
    .D(_00762_),
    .Q_N(_10043_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[7] ));
 sg13g2_dfrbp_1 _19423_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net4213),
    .D(_00763_),
    .Q_N(_10042_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19424_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net4228),
    .D(_00764_),
    .Q_N(_10041_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19425_ (.CLK(net4515),
    .RESET_B(net4227),
    .D(_00765_),
    .Q_N(_10040_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[0] ));
 sg13g2_dfrbp_1 _19426_ (.CLK(net4515),
    .RESET_B(net4224),
    .D(_00766_),
    .Q_N(_10039_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[1] ));
 sg13g2_dfrbp_1 _19427_ (.CLK(net4515),
    .RESET_B(net4224),
    .D(_00767_),
    .Q_N(_10038_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[2] ));
 sg13g2_dfrbp_1 _19428_ (.CLK(net4514),
    .RESET_B(net4224),
    .D(_00768_),
    .Q_N(_10037_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[3] ));
 sg13g2_dfrbp_1 _19429_ (.CLK(net4515),
    .RESET_B(net4225),
    .D(_00769_),
    .Q_N(_10036_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[4] ));
 sg13g2_dfrbp_1 _19430_ (.CLK(net4515),
    .RESET_B(net4225),
    .D(_00770_),
    .Q_N(_10035_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[5] ));
 sg13g2_dfrbp_1 _19431_ (.CLK(net4515),
    .RESET_B(net4224),
    .D(_00771_),
    .Q_N(_10034_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[6] ));
 sg13g2_dfrbp_1 _19432_ (.CLK(net4515),
    .RESET_B(net4224),
    .D(_00772_),
    .Q_N(_10033_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[7] ));
 sg13g2_dfrbp_1 _19433_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net4228),
    .D(_00773_),
    .Q_N(_10032_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19434_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net4224),
    .D(_00774_),
    .Q_N(_10031_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19435_ (.CLK(net4500),
    .RESET_B(net4187),
    .D(_00775_),
    .Q_N(_10030_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[0] ));
 sg13g2_dfrbp_1 _19436_ (.CLK(net4500),
    .RESET_B(net4187),
    .D(_00776_),
    .Q_N(_10029_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[1] ));
 sg13g2_dfrbp_1 _19437_ (.CLK(net4500),
    .RESET_B(net4187),
    .D(_00777_),
    .Q_N(_10028_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[2] ));
 sg13g2_dfrbp_1 _19438_ (.CLK(net4500),
    .RESET_B(net4191),
    .D(_00778_),
    .Q_N(_10027_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[3] ));
 sg13g2_dfrbp_1 _19439_ (.CLK(net4500),
    .RESET_B(net4187),
    .D(_00779_),
    .Q_N(_10026_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[4] ));
 sg13g2_dfrbp_1 _19440_ (.CLK(net4508),
    .RESET_B(net4191),
    .D(_00780_),
    .Q_N(_10025_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[5] ));
 sg13g2_dfrbp_1 _19441_ (.CLK(net4500),
    .RESET_B(net4190),
    .D(_00781_),
    .Q_N(_10024_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[6] ));
 sg13g2_dfrbp_1 _19442_ (.CLK(net4500),
    .RESET_B(net4191),
    .D(_00782_),
    .Q_N(_10023_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[7] ));
 sg13g2_dfrbp_1 _19443_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net4226),
    .D(_00783_),
    .Q_N(_10022_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19444_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net4180),
    .D(_00784_),
    .Q_N(_10021_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19445_ (.CLK(net4506),
    .RESET_B(net4200),
    .D(_00785_),
    .Q_N(_10020_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[0] ));
 sg13g2_dfrbp_1 _19446_ (.CLK(net4506),
    .RESET_B(net4198),
    .D(_00786_),
    .Q_N(_10019_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[1] ));
 sg13g2_dfrbp_1 _19447_ (.CLK(net4506),
    .RESET_B(net4198),
    .D(_00787_),
    .Q_N(_10018_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[2] ));
 sg13g2_dfrbp_1 _19448_ (.CLK(net4506),
    .RESET_B(net4198),
    .D(_00788_),
    .Q_N(_10017_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[3] ));
 sg13g2_dfrbp_1 _19449_ (.CLK(net4504),
    .RESET_B(net4198),
    .D(_00789_),
    .Q_N(_10016_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[4] ));
 sg13g2_dfrbp_1 _19450_ (.CLK(net4504),
    .RESET_B(net4195),
    .D(_00790_),
    .Q_N(_10015_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[5] ));
 sg13g2_dfrbp_1 _19451_ (.CLK(net4504),
    .RESET_B(net4195),
    .D(_00791_),
    .Q_N(_10014_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[6] ));
 sg13g2_dfrbp_1 _19452_ (.CLK(net4504),
    .RESET_B(net4198),
    .D(_00792_),
    .Q_N(_10013_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[7] ));
 sg13g2_dfrbp_1 _19453_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net4180),
    .D(_00793_),
    .Q_N(_10012_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19454_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net4200),
    .D(_00794_),
    .Q_N(_10011_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19455_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net4143),
    .D(net366),
    .Q_N(_00090_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[0] ));
 sg13g2_dfrbp_1 _19456_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net4143),
    .D(_00796_),
    .Q_N(_10010_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[1] ));
 sg13g2_dfrbp_1 _19457_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net4141),
    .D(net211),
    .Q_N(_10009_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[2] ));
 sg13g2_dfrbp_1 _19458_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net4141),
    .D(net442),
    .Q_N(_10008_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[3] ));
 sg13g2_dfrbp_1 _19459_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net4150),
    .D(_00799_),
    .Q_N(_10007_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[4] ));
 sg13g2_dfrbp_1 _19460_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net4191),
    .D(net197),
    .Q_N(_10006_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19461_ (.CLK(net4510),
    .RESET_B(net4207),
    .D(_00801_),
    .Q_N(_10005_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[0] ));
 sg13g2_dfrbp_1 _19462_ (.CLK(net4510),
    .RESET_B(net4210),
    .D(_00802_),
    .Q_N(_10004_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[1] ));
 sg13g2_dfrbp_1 _19463_ (.CLK(net4510),
    .RESET_B(net4210),
    .D(_00803_),
    .Q_N(_10003_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[2] ));
 sg13g2_dfrbp_1 _19464_ (.CLK(net4510),
    .RESET_B(net4210),
    .D(_00804_),
    .Q_N(_10002_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[3] ));
 sg13g2_dfrbp_1 _19465_ (.CLK(net4510),
    .RESET_B(net4210),
    .D(_00805_),
    .Q_N(_10001_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[4] ));
 sg13g2_dfrbp_1 _19466_ (.CLK(net4510),
    .RESET_B(net4207),
    .D(_00806_),
    .Q_N(_10000_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[5] ));
 sg13g2_dfrbp_1 _19467_ (.CLK(net4510),
    .RESET_B(net4207),
    .D(_00807_),
    .Q_N(_10340_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[6] ));
 sg13g2_dfrbp_1 _19468_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net4173),
    .D(_00016_),
    .Q_N(_09999_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.spike_out ));
 sg13g2_dfrbp_1 _19469_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net4173),
    .D(_00808_),
    .Q_N(_00088_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[0] ));
 sg13g2_dfrbp_1 _19470_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net4173),
    .D(_00809_),
    .Q_N(_00089_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ));
 sg13g2_dfrbp_1 _19471_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net4173),
    .D(_00810_),
    .Q_N(_00087_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ));
 sg13g2_dfrbp_1 _19472_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net4173),
    .D(_00811_),
    .Q_N(_00086_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ));
 sg13g2_dfrbp_1 _19473_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net4173),
    .D(_00812_),
    .Q_N(_00085_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ));
 sg13g2_dfrbp_1 _19474_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net4254),
    .D(_00813_),
    .Q_N(_09998_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19475_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net4252),
    .D(_00814_),
    .Q_N(_09997_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19476_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net4256),
    .D(_00815_),
    .Q_N(_09996_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19477_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net4255),
    .D(_00816_),
    .Q_N(_09995_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19478_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net4218),
    .D(_00817_),
    .Q_N(_09994_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19479_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net4215),
    .D(_00818_),
    .Q_N(_09993_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19480_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net4230),
    .D(_00819_),
    .Q_N(_09992_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19481_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net4230),
    .D(_00820_),
    .Q_N(_09991_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19482_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net4243),
    .D(_00821_),
    .Q_N(_09990_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19483_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net4243),
    .D(_00822_),
    .Q_N(_09989_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19484_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net4240),
    .D(_00823_),
    .Q_N(_09988_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19485_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net4240),
    .D(_00824_),
    .Q_N(_09987_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19486_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net4251),
    .D(_00825_),
    .Q_N(_09986_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19487_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net4247),
    .D(_00826_),
    .Q_N(_09985_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19488_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net4248),
    .D(_00827_),
    .Q_N(_09984_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19489_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net4188),
    .D(net358),
    .Q_N(_00096_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[0] ));
 sg13g2_dfrbp_1 _19490_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net4188),
    .D(_00829_),
    .Q_N(_09983_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[1] ));
 sg13g2_dfrbp_1 _19491_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net4188),
    .D(net174),
    .Q_N(_09982_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[2] ));
 sg13g2_dfrbp_1 _19492_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net4188),
    .D(_00831_),
    .Q_N(_09981_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[3] ));
 sg13g2_dfrbp_1 _19493_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net4188),
    .D(_00832_),
    .Q_N(_09980_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[4] ));
 sg13g2_dfrbp_1 _19494_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net4248),
    .D(_00833_),
    .Q_N(_09979_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19495_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net4159),
    .D(_00834_),
    .Q_N(_09978_),
    .Q(\spiking_network_top_uut.debug_inst.debug_config[0] ));
 sg13g2_dfrbp_1 _19496_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net4147),
    .D(_00835_),
    .Q_N(_09977_),
    .Q(\spiking_network_top_uut.debug_inst.debug_config[1] ));
 sg13g2_dfrbp_1 _19497_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net4158),
    .D(_00836_),
    .Q_N(_09976_),
    .Q(\spiking_network_top_uut.debug_inst.debug_config[2] ));
 sg13g2_dfrbp_1 _19498_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net4147),
    .D(_00837_),
    .Q_N(_09975_),
    .Q(\spiking_network_top_uut.debug_inst.debug_config[3] ));
 sg13g2_dfrbp_1 _19499_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net4143),
    .D(_00838_),
    .Q_N(_09974_),
    .Q(\spiking_network_top_uut.debug_inst.debug_config[4] ));
 sg13g2_dfrbp_1 _19500_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net4142),
    .D(_00839_),
    .Q_N(_09973_),
    .Q(\spiking_network_top_uut.debug_inst.debug_config[5] ));
 sg13g2_dfrbp_1 _19501_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net4142),
    .D(_00840_),
    .Q_N(_09972_),
    .Q(\spiking_network_top_uut.debug_inst.debug_config[6] ));
 sg13g2_dfrbp_1 _19502_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net4142),
    .D(_00841_),
    .Q_N(_10341_),
    .Q(\spiking_network_top_uut.debug_inst.debug_config[7] ));
 sg13g2_dfrbp_1 _19503_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net4189),
    .D(_00001_),
    .Q_N(_09971_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.spike_out ));
 sg13g2_dfrbp_1 _19504_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net4188),
    .D(_00842_),
    .Q_N(_00094_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[0] ));
 sg13g2_dfrbp_1 _19505_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net4189),
    .D(_00843_),
    .Q_N(_00095_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ));
 sg13g2_dfrbp_1 _19506_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net4189),
    .D(_00844_),
    .Q_N(_00093_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ));
 sg13g2_dfrbp_1 _19507_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net4174),
    .D(_00845_),
    .Q_N(_00092_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ));
 sg13g2_dfrbp_1 _19508_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net4189),
    .D(_00846_),
    .Q_N(_00091_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ));
 sg13g2_dfrbp_1 _19509_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net4253),
    .D(_00847_),
    .Q_N(_09970_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19510_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net4257),
    .D(_00848_),
    .Q_N(_09969_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19511_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net4255),
    .D(_00849_),
    .Q_N(_09968_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19512_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net4250),
    .D(_00850_),
    .Q_N(_09967_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19513_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net4217),
    .D(_00851_),
    .Q_N(_09966_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19514_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net4216),
    .D(net126),
    .Q_N(_09965_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19515_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net4229),
    .D(_00853_),
    .Q_N(_09964_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19516_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net4230),
    .D(_00854_),
    .Q_N(_09963_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19517_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net4244),
    .D(_00855_),
    .Q_N(_09962_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19518_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net4244),
    .D(net39),
    .Q_N(_09961_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19519_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net4240),
    .D(_00857_),
    .Q_N(_09960_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19520_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net4240),
    .D(_00858_),
    .Q_N(_09959_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19521_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net4250),
    .D(_00859_),
    .Q_N(_09958_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19522_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net4250),
    .D(net44),
    .Q_N(_09957_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19523_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net4248),
    .D(_00861_),
    .Q_N(_09956_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19524_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net4154),
    .D(net380),
    .Q_N(_00102_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[0] ));
 sg13g2_dfrbp_1 _19525_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net4154),
    .D(_00863_),
    .Q_N(_09955_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[1] ));
 sg13g2_dfrbp_1 _19526_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net4154),
    .D(_00864_),
    .Q_N(_09954_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[2] ));
 sg13g2_dfrbp_1 _19527_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net4154),
    .D(_00865_),
    .Q_N(_09953_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[3] ));
 sg13g2_dfrbp_1 _19528_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net4154),
    .D(_00866_),
    .Q_N(_09952_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[4] ));
 sg13g2_dfrbp_1 _19529_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net4249),
    .D(_00867_),
    .Q_N(_10342_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19530_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net4173),
    .D(_00002_),
    .Q_N(_09951_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.spike_out ));
 sg13g2_dfrbp_1 _19531_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net4170),
    .D(_00868_),
    .Q_N(_00100_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[0] ));
 sg13g2_dfrbp_1 _19532_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net4170),
    .D(_00869_),
    .Q_N(_00101_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ));
 sg13g2_dfrbp_1 _19533_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net4172),
    .D(_00870_),
    .Q_N(_00099_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ));
 sg13g2_dfrbp_1 _19534_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net4172),
    .D(_00871_),
    .Q_N(_00098_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ));
 sg13g2_dfrbp_1 _19535_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net4172),
    .D(_00872_),
    .Q_N(_00097_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ));
 sg13g2_dfrbp_1 _19536_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net4254),
    .D(_00873_),
    .Q_N(_09950_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19537_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net4252),
    .D(_00874_),
    .Q_N(_09949_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19538_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net4257),
    .D(_00875_),
    .Q_N(_09948_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19539_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net4253),
    .D(_00876_),
    .Q_N(_09947_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19540_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net4217),
    .D(_00877_),
    .Q_N(_09946_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19541_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net4217),
    .D(_00878_),
    .Q_N(_09945_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19542_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net4217),
    .D(_00879_),
    .Q_N(_09944_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19543_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net4217),
    .D(_00880_),
    .Q_N(_09943_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19544_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net4245),
    .D(_00881_),
    .Q_N(_09942_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19545_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net4245),
    .D(_00882_),
    .Q_N(_09941_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19546_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net4238),
    .D(_00883_),
    .Q_N(_09940_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19547_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net4238),
    .D(_00884_),
    .Q_N(_09939_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19548_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net4246),
    .D(_00885_),
    .Q_N(_09938_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19549_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net4247),
    .D(_00886_),
    .Q_N(_09937_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19550_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net4249),
    .D(_00887_),
    .Q_N(_09936_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19551_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net4171),
    .D(net304),
    .Q_N(_00108_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[0] ));
 sg13g2_dfrbp_1 _19552_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net4170),
    .D(_00889_),
    .Q_N(_09935_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[1] ));
 sg13g2_dfrbp_1 _19553_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net4170),
    .D(net195),
    .Q_N(_09934_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[2] ));
 sg13g2_dfrbp_1 _19554_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net4170),
    .D(_00891_),
    .Q_N(_09933_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[3] ));
 sg13g2_dfrbp_1 _19555_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net4171),
    .D(_00892_),
    .Q_N(_09932_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[4] ));
 sg13g2_dfrbp_1 _19556_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net4249),
    .D(_00893_),
    .Q_N(_10343_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19557_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net4169),
    .D(_00003_),
    .Q_N(_09931_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.spike_out ));
 sg13g2_dfrbp_1 _19558_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net4168),
    .D(_00894_),
    .Q_N(_00106_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[0] ));
 sg13g2_dfrbp_1 _19559_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net4169),
    .D(_00895_),
    .Q_N(_00107_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ));
 sg13g2_dfrbp_1 _19560_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net4168),
    .D(_00896_),
    .Q_N(_00105_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ));
 sg13g2_dfrbp_1 _19561_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net4168),
    .D(_00897_),
    .Q_N(_00104_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ));
 sg13g2_dfrbp_1 _19562_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net4168),
    .D(_00898_),
    .Q_N(_00103_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ));
 sg13g2_dfrbp_1 _19563_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net4252),
    .D(_00899_),
    .Q_N(_09930_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19564_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net4252),
    .D(_00900_),
    .Q_N(_09929_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19565_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net4255),
    .D(_00901_),
    .Q_N(_09928_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19566_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net4250),
    .D(_00902_),
    .Q_N(_09927_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19567_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net4215),
    .D(_00903_),
    .Q_N(_09926_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19568_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net4215),
    .D(net163),
    .Q_N(_09925_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19569_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net4229),
    .D(_00905_),
    .Q_N(_09924_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19570_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net4229),
    .D(_00906_),
    .Q_N(_09923_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19571_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net4242),
    .D(_00907_),
    .Q_N(_09922_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19572_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net4242),
    .D(_00908_),
    .Q_N(_09921_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19573_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net4237),
    .D(_00909_),
    .Q_N(_09920_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19574_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net4239),
    .D(_00910_),
    .Q_N(_09919_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19575_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net4249),
    .D(_00911_),
    .Q_N(_09918_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19576_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net4249),
    .D(net42),
    .Q_N(_09917_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19577_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net4234),
    .D(_00913_),
    .Q_N(_09916_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19578_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net4155),
    .D(net395),
    .Q_N(_00114_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[0] ));
 sg13g2_dfrbp_1 _19579_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net4155),
    .D(net413),
    .Q_N(_09915_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[1] ));
 sg13g2_dfrbp_1 _19580_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net4155),
    .D(_00916_),
    .Q_N(_09914_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[2] ));
 sg13g2_dfrbp_1 _19581_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net4157),
    .D(_00917_),
    .Q_N(_09913_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[3] ));
 sg13g2_dfrbp_1 _19582_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net4157),
    .D(_00918_),
    .Q_N(_09912_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[4] ));
 sg13g2_dfrbp_1 _19583_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net4248),
    .D(_00919_),
    .Q_N(_10344_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19584_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net4159),
    .D(_00004_),
    .Q_N(_09911_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.spike_out ));
 sg13g2_dfrbp_1 _19585_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net4160),
    .D(_00920_),
    .Q_N(_00112_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[0] ));
 sg13g2_dfrbp_1 _19586_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net4160),
    .D(_00921_),
    .Q_N(_00113_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ));
 sg13g2_dfrbp_1 _19587_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net4160),
    .D(_00922_),
    .Q_N(_00111_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ));
 sg13g2_dfrbp_1 _19588_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net4160),
    .D(_00923_),
    .Q_N(_00110_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ));
 sg13g2_dfrbp_1 _19589_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net4160),
    .D(_00924_),
    .Q_N(_00109_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ));
 sg13g2_dfrbp_1 _19590_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net4253),
    .D(_00925_),
    .Q_N(_09910_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19591_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net4258),
    .D(_00926_),
    .Q_N(_09909_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19592_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net4255),
    .D(_00927_),
    .Q_N(_09908_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19593_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net4255),
    .D(_00928_),
    .Q_N(_09907_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19594_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net4215),
    .D(_00929_),
    .Q_N(_09906_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19595_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net4209),
    .D(net56),
    .Q_N(_09905_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19596_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net4234),
    .D(_00931_),
    .Q_N(_09904_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19597_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net4234),
    .D(_00932_),
    .Q_N(_09903_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19598_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net4242),
    .D(_00933_),
    .Q_N(_09902_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19599_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net4243),
    .D(_00934_),
    .Q_N(_09901_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19600_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net4237),
    .D(_00935_),
    .Q_N(_09900_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19601_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net4243),
    .D(_00936_),
    .Q_N(_09899_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19602_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net4246),
    .D(_00937_),
    .Q_N(_09898_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19603_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net4249),
    .D(net152),
    .Q_N(_09897_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19604_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net4235),
    .D(_00939_),
    .Q_N(_09896_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19605_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net4192),
    .D(net330),
    .Q_N(_00120_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[0] ));
 sg13g2_dfrbp_1 _19606_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net4192),
    .D(_00941_),
    .Q_N(_09895_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[1] ));
 sg13g2_dfrbp_1 _19607_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net4192),
    .D(_00942_),
    .Q_N(_09894_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[2] ));
 sg13g2_dfrbp_1 _19608_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net4192),
    .D(_00943_),
    .Q_N(_09893_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[3] ));
 sg13g2_dfrbp_1 _19609_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net4192),
    .D(_00944_),
    .Q_N(_09892_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[4] ));
 sg13g2_dfrbp_1 _19610_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net4235),
    .D(_00945_),
    .Q_N(_10345_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19611_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net4191),
    .D(_00005_),
    .Q_N(_09891_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.spike_out ));
 sg13g2_dfrbp_1 _19612_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net4189),
    .D(_00946_),
    .Q_N(_00118_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[0] ));
 sg13g2_dfrbp_1 _19613_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net4188),
    .D(_00947_),
    .Q_N(_00119_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ));
 sg13g2_dfrbp_1 _19614_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net4189),
    .D(_00948_),
    .Q_N(_00117_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ));
 sg13g2_dfrbp_1 _19615_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net4188),
    .D(_00949_),
    .Q_N(_00116_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ));
 sg13g2_dfrbp_1 _19616_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net4189),
    .D(_00950_),
    .Q_N(_00115_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ));
 sg13g2_dfrbp_1 _19617_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net4254),
    .D(_00951_),
    .Q_N(_09890_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19618_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net4253),
    .D(_00952_),
    .Q_N(_09889_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19619_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net4257),
    .D(_00953_),
    .Q_N(_09888_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19620_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net4257),
    .D(_00954_),
    .Q_N(_09887_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19621_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net4216),
    .D(_00955_),
    .Q_N(_09886_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19622_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net4217),
    .D(_00956_),
    .Q_N(_09885_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19623_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net4229),
    .D(_00957_),
    .Q_N(_09884_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19624_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net4229),
    .D(_00958_),
    .Q_N(_09883_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19625_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net4245),
    .D(_00959_),
    .Q_N(_09882_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19626_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net4245),
    .D(_00960_),
    .Q_N(_09881_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19627_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net4237),
    .D(_00961_),
    .Q_N(_09880_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19628_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net4237),
    .D(_00962_),
    .Q_N(_09879_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19629_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net4246),
    .D(_00963_),
    .Q_N(_09878_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19630_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net4246),
    .D(net50),
    .Q_N(_09877_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19631_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net4249),
    .D(_00965_),
    .Q_N(_09876_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19632_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net4155),
    .D(net341),
    .Q_N(_00126_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[0] ));
 sg13g2_dfrbp_1 _19633_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net4157),
    .D(net388),
    .Q_N(_09875_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[1] ));
 sg13g2_dfrbp_1 _19634_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net4155),
    .D(_00968_),
    .Q_N(_09874_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[2] ));
 sg13g2_dfrbp_1 _19635_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net4157),
    .D(_00969_),
    .Q_N(_09873_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[3] ));
 sg13g2_dfrbp_1 _19636_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net4156),
    .D(_00970_),
    .Q_N(_09872_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[4] ));
 sg13g2_dfrbp_1 _19637_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net4250),
    .D(_00971_),
    .Q_N(_10346_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19638_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net4159),
    .D(_00006_),
    .Q_N(_09871_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.spike_out ));
 sg13g2_dfrbp_1 _19639_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net4152),
    .D(_00972_),
    .Q_N(_00124_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[0] ));
 sg13g2_dfrbp_1 _19640_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net4152),
    .D(_00973_),
    .Q_N(_00125_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ));
 sg13g2_dfrbp_1 _19641_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net4153),
    .D(_00974_),
    .Q_N(_00123_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ));
 sg13g2_dfrbp_1 _19642_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net4153),
    .D(_00975_),
    .Q_N(_00122_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ));
 sg13g2_dfrbp_1 _19643_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net4150),
    .D(_00976_),
    .Q_N(_00121_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ));
 sg13g2_dfrbp_1 _19644_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net4254),
    .D(_00977_),
    .Q_N(_09870_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19645_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net4252),
    .D(_00978_),
    .Q_N(_09869_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19646_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net4257),
    .D(_00979_),
    .Q_N(_09868_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19647_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net4252),
    .D(_00980_),
    .Q_N(_09867_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19648_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net4218),
    .D(_00981_),
    .Q_N(_09866_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19649_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net4215),
    .D(net308),
    .Q_N(_09865_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19650_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net4218),
    .D(_00983_),
    .Q_N(_09864_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19651_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net4217),
    .D(_00984_),
    .Q_N(_09863_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19652_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net4245),
    .D(_00985_),
    .Q_N(_09862_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19653_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net4244),
    .D(net46),
    .Q_N(_09861_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19654_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net4241),
    .D(_00987_),
    .Q_N(_09860_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19655_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net4240),
    .D(_00988_),
    .Q_N(_09859_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19656_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net4240),
    .D(_00989_),
    .Q_N(_09858_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19657_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net4251),
    .D(_00990_),
    .Q_N(_09857_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19658_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net4233),
    .D(_00991_),
    .Q_N(_09856_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19659_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net4151),
    .D(net364),
    .Q_N(_00132_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[0] ));
 sg13g2_dfrbp_1 _19660_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net4151),
    .D(_00993_),
    .Q_N(_09855_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[1] ));
 sg13g2_dfrbp_1 _19661_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net4151),
    .D(_00994_),
    .Q_N(_09854_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[2] ));
 sg13g2_dfrbp_1 _19662_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net4150),
    .D(net440),
    .Q_N(_09853_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[3] ));
 sg13g2_dfrbp_1 _19663_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net4150),
    .D(_00996_),
    .Q_N(_09852_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[4] ));
 sg13g2_dfrbp_1 _19664_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net4233),
    .D(_00997_),
    .Q_N(_10347_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19665_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net4159),
    .D(_00007_),
    .Q_N(_09851_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.spike_out ));
 sg13g2_dfrbp_1 _19666_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net4158),
    .D(_00998_),
    .Q_N(_00130_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[0] ));
 sg13g2_dfrbp_1 _19667_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net4152),
    .D(_00999_),
    .Q_N(_00131_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ));
 sg13g2_dfrbp_1 _19668_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net4158),
    .D(_01000_),
    .Q_N(_00129_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ));
 sg13g2_dfrbp_1 _19669_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net4152),
    .D(_01001_),
    .Q_N(_00128_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ));
 sg13g2_dfrbp_1 _19670_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net4152),
    .D(_01002_),
    .Q_N(_00127_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ));
 sg13g2_dfrbp_1 _19671_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net4252),
    .D(_01003_),
    .Q_N(_09850_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19672_ (.CLK(net4524),
    .RESET_B(net4250),
    .D(_01004_),
    .Q_N(_09849_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[0] ));
 sg13g2_dfrbp_1 _19673_ (.CLK(net4525),
    .RESET_B(net4256),
    .D(_01005_),
    .Q_N(_09848_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[1] ));
 sg13g2_dfrbp_1 _19674_ (.CLK(net4525),
    .RESET_B(net4255),
    .D(_01006_),
    .Q_N(_09847_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[2] ));
 sg13g2_dfrbp_1 _19675_ (.CLK(net4523),
    .RESET_B(net4255),
    .D(_01007_),
    .Q_N(_09846_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[3] ));
 sg13g2_dfrbp_1 _19676_ (.CLK(net4523),
    .RESET_B(net4257),
    .D(_01008_),
    .Q_N(_09845_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[4] ));
 sg13g2_dfrbp_1 _19677_ (.CLK(net4525),
    .RESET_B(net4258),
    .D(_01009_),
    .Q_N(_09844_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[5] ));
 sg13g2_dfrbp_1 _19678_ (.CLK(net4523),
    .RESET_B(net4257),
    .D(_01010_),
    .Q_N(_09843_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[6] ));
 sg13g2_dfrbp_1 _19679_ (.CLK(net4523),
    .RESET_B(net4255),
    .D(_01011_),
    .Q_N(_09842_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[7] ));
 sg13g2_dfrbp_1 _19680_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net4252),
    .D(_01012_),
    .Q_N(_09841_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19681_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net4256),
    .D(_01013_),
    .Q_N(_09840_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19682_ (.CLK(net4528),
    .RESET_B(net4215),
    .D(_01014_),
    .Q_N(_09839_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[0] ));
 sg13g2_dfrbp_1 _19683_ (.CLK(net4512),
    .RESET_B(net4216),
    .D(_01015_),
    .Q_N(_09838_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[1] ));
 sg13g2_dfrbp_1 _19684_ (.CLK(net4512),
    .RESET_B(net4216),
    .D(_01016_),
    .Q_N(_09837_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[2] ));
 sg13g2_dfrbp_1 _19685_ (.CLK(net4512),
    .RESET_B(net4216),
    .D(_01017_),
    .Q_N(_09836_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[3] ));
 sg13g2_dfrbp_1 _19686_ (.CLK(net4512),
    .RESET_B(net4216),
    .D(_01018_),
    .Q_N(_09835_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[4] ));
 sg13g2_dfrbp_1 _19687_ (.CLK(net4512),
    .RESET_B(net4215),
    .D(_01019_),
    .Q_N(_09834_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[5] ));
 sg13g2_dfrbp_1 _19688_ (.CLK(net4512),
    .RESET_B(net4215),
    .D(_01020_),
    .Q_N(_09833_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[6] ));
 sg13g2_dfrbp_1 _19689_ (.CLK(net4512),
    .RESET_B(net4216),
    .D(_01021_),
    .Q_N(_09832_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[7] ));
 sg13g2_dfrbp_1 _19690_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net4250),
    .D(net48),
    .Q_N(_09831_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19691_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net4216),
    .D(_01023_),
    .Q_N(_09830_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19692_ (.CLK(net4512),
    .RESET_B(net4229),
    .D(_01024_),
    .Q_N(_09829_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[0] ));
 sg13g2_dfrbp_1 _19693_ (.CLK(net4519),
    .RESET_B(net4229),
    .D(_01025_),
    .Q_N(_09828_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[1] ));
 sg13g2_dfrbp_1 _19694_ (.CLK(net4519),
    .RESET_B(net4234),
    .D(_01026_),
    .Q_N(_09827_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[2] ));
 sg13g2_dfrbp_1 _19695_ (.CLK(net4519),
    .RESET_B(net4234),
    .D(_01027_),
    .Q_N(_09826_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[3] ));
 sg13g2_dfrbp_1 _19696_ (.CLK(net4516),
    .RESET_B(net4234),
    .D(_01028_),
    .Q_N(_09825_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[4] ));
 sg13g2_dfrbp_1 _19697_ (.CLK(net4516),
    .RESET_B(net4229),
    .D(_01029_),
    .Q_N(_09824_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[5] ));
 sg13g2_dfrbp_1 _19698_ (.CLK(net4516),
    .RESET_B(net4230),
    .D(_01030_),
    .Q_N(_09823_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[6] ));
 sg13g2_dfrbp_1 _19699_ (.CLK(net4516),
    .RESET_B(net4230),
    .D(_01031_),
    .Q_N(_09822_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[7] ));
 sg13g2_dfrbp_1 _19700_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net4209),
    .D(net272),
    .Q_N(_09821_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19701_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net4234),
    .D(_01033_),
    .Q_N(_09820_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19702_ (.CLK(net4520),
    .RESET_B(net4243),
    .D(_01034_),
    .Q_N(_09819_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[0] ));
 sg13g2_dfrbp_1 _19703_ (.CLK(net4520),
    .RESET_B(net4242),
    .D(_01035_),
    .Q_N(_09818_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[1] ));
 sg13g2_dfrbp_1 _19704_ (.CLK(net4520),
    .RESET_B(net4242),
    .D(_01036_),
    .Q_N(_09817_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[2] ));
 sg13g2_dfrbp_1 _19705_ (.CLK(net4520),
    .RESET_B(net4242),
    .D(_01037_),
    .Q_N(_09816_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[3] ));
 sg13g2_dfrbp_1 _19706_ (.CLK(net4520),
    .RESET_B(net4243),
    .D(_01038_),
    .Q_N(_09815_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[4] ));
 sg13g2_dfrbp_1 _19707_ (.CLK(net4520),
    .RESET_B(net4242),
    .D(_01039_),
    .Q_N(_09814_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[5] ));
 sg13g2_dfrbp_1 _19708_ (.CLK(net4520),
    .RESET_B(net4243),
    .D(_01040_),
    .Q_N(_09813_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[6] ));
 sg13g2_dfrbp_1 _19709_ (.CLK(net4520),
    .RESET_B(net4242),
    .D(_01041_),
    .Q_N(_09812_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[7] ));
 sg13g2_dfrbp_1 _19710_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net4234),
    .D(_01042_),
    .Q_N(_09811_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19711_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net4244),
    .D(_01043_),
    .Q_N(_09810_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19712_ (.CLK(net4522),
    .RESET_B(net4239),
    .D(_01044_),
    .Q_N(_09809_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[0] ));
 sg13g2_dfrbp_1 _19713_ (.CLK(net4522),
    .RESET_B(net4237),
    .D(_01045_),
    .Q_N(_09808_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[1] ));
 sg13g2_dfrbp_1 _19714_ (.CLK(net4522),
    .RESET_B(net4237),
    .D(_01046_),
    .Q_N(_09807_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[2] ));
 sg13g2_dfrbp_1 _19715_ (.CLK(net4522),
    .RESET_B(net4238),
    .D(_01047_),
    .Q_N(_09806_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[3] ));
 sg13g2_dfrbp_1 _19716_ (.CLK(net4522),
    .RESET_B(net4237),
    .D(_01048_),
    .Q_N(_09805_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[4] ));
 sg13g2_dfrbp_1 _19717_ (.CLK(net4522),
    .RESET_B(net4238),
    .D(_01049_),
    .Q_N(_09804_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[5] ));
 sg13g2_dfrbp_1 _19718_ (.CLK(net4522),
    .RESET_B(net4238),
    .D(_01050_),
    .Q_N(_09803_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[6] ));
 sg13g2_dfrbp_1 _19719_ (.CLK(net4522),
    .RESET_B(net4237),
    .D(_01051_),
    .Q_N(_09802_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[7] ));
 sg13g2_dfrbp_1 _19720_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net4244),
    .D(_01052_),
    .Q_N(_09801_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19721_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net4240),
    .D(_01053_),
    .Q_N(_09800_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19722_ (.CLK(net4517),
    .RESET_B(net4247),
    .D(_01054_),
    .Q_N(_09799_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[0] ));
 sg13g2_dfrbp_1 _19723_ (.CLK(net4524),
    .RESET_B(net4246),
    .D(_01055_),
    .Q_N(_09798_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[1] ));
 sg13g2_dfrbp_1 _19724_ (.CLK(net4524),
    .RESET_B(net4247),
    .D(_01056_),
    .Q_N(_09797_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[2] ));
 sg13g2_dfrbp_1 _19725_ (.CLK(net4524),
    .RESET_B(net4247),
    .D(_01057_),
    .Q_N(_09796_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[3] ));
 sg13g2_dfrbp_1 _19726_ (.CLK(net4524),
    .RESET_B(net4246),
    .D(_01058_),
    .Q_N(_09795_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[4] ));
 sg13g2_dfrbp_1 _19727_ (.CLK(net4524),
    .RESET_B(net4251),
    .D(_01059_),
    .Q_N(_09794_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[5] ));
 sg13g2_dfrbp_1 _19728_ (.CLK(net4524),
    .RESET_B(net4247),
    .D(_01060_),
    .Q_N(_09793_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[6] ));
 sg13g2_dfrbp_1 _19729_ (.CLK(net4524),
    .RESET_B(net4247),
    .D(_01061_),
    .Q_N(_09792_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[7] ));
 sg13g2_dfrbp_1 _19730_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net4240),
    .D(_01062_),
    .Q_N(_09791_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19731_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net4246),
    .D(_01063_),
    .Q_N(_09790_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19732_ (.CLK(net4517),
    .RESET_B(net4235),
    .D(_01064_),
    .Q_N(_09789_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[0] ));
 sg13g2_dfrbp_1 _19733_ (.CLK(net4518),
    .RESET_B(net4248),
    .D(_01065_),
    .Q_N(_09788_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[1] ));
 sg13g2_dfrbp_1 _19734_ (.CLK(net4517),
    .RESET_B(net4248),
    .D(_01066_),
    .Q_N(_09787_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[2] ));
 sg13g2_dfrbp_1 _19735_ (.CLK(net4517),
    .RESET_B(net4248),
    .D(_01067_),
    .Q_N(_09786_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[3] ));
 sg13g2_dfrbp_1 _19736_ (.CLK(net4518),
    .RESET_B(net4248),
    .D(_01068_),
    .Q_N(_09785_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[4] ));
 sg13g2_dfrbp_1 _19737_ (.CLK(net4517),
    .RESET_B(net4235),
    .D(_01069_),
    .Q_N(_09784_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[5] ));
 sg13g2_dfrbp_1 _19738_ (.CLK(net4518),
    .RESET_B(net4235),
    .D(_01070_),
    .Q_N(_09783_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[6] ));
 sg13g2_dfrbp_1 _19739_ (.CLK(net4518),
    .RESET_B(net4235),
    .D(_01071_),
    .Q_N(_09782_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[7] ));
 sg13g2_dfrbp_1 _19740_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net4246),
    .D(_01072_),
    .Q_N(_09781_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19741_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net4250),
    .D(_01073_),
    .Q_N(_09780_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_reg1 ));
 sg13g2_dfrbp_1 _19742_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net4151),
    .D(net391),
    .Q_N(_00138_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[0] ));
 sg13g2_dfrbp_1 _19743_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net4151),
    .D(net408),
    .Q_N(_09779_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[1] ));
 sg13g2_dfrbp_1 _19744_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net4151),
    .D(_01076_),
    .Q_N(_09778_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[2] ));
 sg13g2_dfrbp_1 _19745_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net4150),
    .D(_01077_),
    .Q_N(_09777_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[3] ));
 sg13g2_dfrbp_1 _19746_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net4152),
    .D(_01078_),
    .Q_N(_09776_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[4] ));
 sg13g2_dfrbp_1 _19747_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net4251),
    .D(_01079_),
    .Q_N(_09775_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_dout ));
 sg13g2_dfrbp_1 _19748_ (.CLK(net4523),
    .RESET_B(net4258),
    .D(_01080_),
    .Q_N(_09774_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[0] ));
 sg13g2_dfrbp_1 _19749_ (.CLK(net4523),
    .RESET_B(net4254),
    .D(_01081_),
    .Q_N(_09773_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[1] ));
 sg13g2_dfrbp_1 _19750_ (.CLK(net4521),
    .RESET_B(net4245),
    .D(_01082_),
    .Q_N(_09772_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[2] ));
 sg13g2_dfrbp_1 _19751_ (.CLK(net4521),
    .RESET_B(net4244),
    .D(_01083_),
    .Q_N(_09771_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[3] ));
 sg13g2_dfrbp_1 _19752_ (.CLK(net4521),
    .RESET_B(net4244),
    .D(_01084_),
    .Q_N(_09770_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[4] ));
 sg13g2_dfrbp_1 _19753_ (.CLK(net4521),
    .RESET_B(net4244),
    .D(_01085_),
    .Q_N(_09769_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[5] ));
 sg13g2_dfrbp_1 _19754_ (.CLK(net4523),
    .RESET_B(net4254),
    .D(_01086_),
    .Q_N(_10348_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[6] ));
 sg13g2_dfrbp_1 _19755_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net4173),
    .D(_00008_),
    .Q_N(_09768_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.spike_out ));
 sg13g2_dfrbp_1 _19756_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net4169),
    .D(_01087_),
    .Q_N(_00136_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[0] ));
 sg13g2_dfrbp_1 _19757_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net4170),
    .D(_01088_),
    .Q_N(_00137_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ));
 sg13g2_dfrbp_1 _19758_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net4170),
    .D(_01089_),
    .Q_N(_00135_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ));
 sg13g2_dfrbp_1 _19759_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net4170),
    .D(_01090_),
    .Q_N(_00134_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ));
 sg13g2_dfrbp_1 _19760_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net4169),
    .D(_01091_),
    .Q_N(_00133_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ));
 sg13g2_dfrbp_1 _19761_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net4145),
    .D(net4529),
    .Q_N(_10349_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.enable_LYR_3 ));
 sg13g2_dfrbp_1 _19762_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net4146),
    .D(net4574),
    .Q_N(_10350_),
    .Q(\spiking_network_top_uut.output_data_ready ));
 sg13g2_dfrbp_1 _19763_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net4235),
    .D(net4617),
    .Q_N(_09767_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.enable_LYR_2 ));
 sg13g2_dfrbp_1 _19764_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net4196),
    .D(_01092_),
    .Q_N(_09766_),
    .Q(\spiking_network_top_uut.clk_div_inst.counter[0] ));
 sg13g2_dfrbp_1 _19765_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net4196),
    .D(net102),
    .Q_N(_09765_),
    .Q(\spiking_network_top_uut.clk_div_inst.counter[1] ));
 sg13g2_dfrbp_1 _19766_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net4196),
    .D(_01094_),
    .Q_N(_09764_),
    .Q(\spiking_network_top_uut.clk_div_inst.counter[2] ));
 sg13g2_dfrbp_1 _19767_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net4185),
    .D(_01095_),
    .Q_N(_09763_),
    .Q(\spiking_network_top_uut.clk_div_inst.counter[3] ));
 sg13g2_dfrbp_1 _19768_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net4186),
    .D(_01096_),
    .Q_N(_09762_),
    .Q(\spiking_network_top_uut.clk_div_inst.counter[4] ));
 sg13g2_dfrbp_1 _19769_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net4185),
    .D(_01097_),
    .Q_N(_09761_),
    .Q(\spiking_network_top_uut.clk_div_inst.counter[5] ));
 sg13g2_dfrbp_1 _19770_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net4185),
    .D(_01098_),
    .Q_N(_09760_),
    .Q(\spiking_network_top_uut.clk_div_inst.counter[6] ));
 sg13g2_dfrbp_1 _19771_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net4196),
    .D(_01099_),
    .Q_N(_09759_),
    .Q(\spiking_network_top_uut.clk_div_inst.counter[7] ));
 sg13g2_dfrbp_1 _19772_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net4197),
    .D(_01100_),
    .Q_N(_00000_),
    .Q(\spiking_network_top_uut.clk_div_inst.clk_out ));
 sg13g2_dfrbp_1 _19773_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net4202),
    .D(_01101_),
    .Q_N(_09758_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.din ));
 sg13g2_dfrbp_1 _19774_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net4202),
    .D(_01102_),
    .Q_N(_09757_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.din ));
 sg13g2_dfrbp_1 _19775_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net4202),
    .D(_01103_),
    .Q_N(_09756_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.din ));
 sg13g2_dfrbp_1 _19776_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net4203),
    .D(_01104_),
    .Q_N(_09755_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.din ));
 sg13g2_dfrbp_1 _19777_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net4202),
    .D(_01105_),
    .Q_N(_09754_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.din ));
 sg13g2_dfrbp_1 _19778_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net4202),
    .D(_01106_),
    .Q_N(_09753_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.din ));
 sg13g2_dfrbp_1 _19779_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net4202),
    .D(_01107_),
    .Q_N(_09752_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.din ));
 sg13g2_dfrbp_1 _19780_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net4202),
    .D(_01108_),
    .Q_N(_09751_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.din ));
 sg13g2_dfrbp_1 _19781_ (.CLK(net4663),
    .RESET_B(net3983),
    .D(_01109_),
    .Q_N(_09750_),
    .Q(\spiking_network_top_uut.clk_div_ready_reg_out ));
 sg13g2_dfrbp_1 _19782_ (.CLK(net4740),
    .RESET_B(net4062),
    .D(_01110_),
    .Q_N(_09749_),
    .Q(\spiking_network_top_uut.spi_inst.LSB_Address_reg[0] ));
 sg13g2_dfrbp_1 _19783_ (.CLK(net4743),
    .RESET_B(net4063),
    .D(_01111_),
    .Q_N(_09748_),
    .Q(\spiking_network_top_uut.spi_inst.LSB_Address_reg[1] ));
 sg13g2_dfrbp_1 _19784_ (.CLK(net4743),
    .RESET_B(net4062),
    .D(_01112_),
    .Q_N(_09747_),
    .Q(\spiking_network_top_uut.spi_inst.LSB_Address_reg[2] ));
 sg13g2_dfrbp_1 _19785_ (.CLK(net4740),
    .RESET_B(net4061),
    .D(_01113_),
    .Q_N(_09746_),
    .Q(\spiking_network_top_uut.spi_inst.LSB_Address_reg[3] ));
 sg13g2_dfrbp_1 _19786_ (.CLK(net4741),
    .RESET_B(net4061),
    .D(_01114_),
    .Q_N(_09745_),
    .Q(\spiking_network_top_uut.spi_inst.LSB_Address_reg[4] ));
 sg13g2_dfrbp_1 _19787_ (.CLK(net4740),
    .RESET_B(net4064),
    .D(_01115_),
    .Q_N(_09744_),
    .Q(\spiking_network_top_uut.spi_inst.LSB_Address_reg[5] ));
 sg13g2_dfrbp_1 _19788_ (.CLK(net4742),
    .RESET_B(net4063),
    .D(_01116_),
    .Q_N(_00027_),
    .Q(\spiking_network_top_uut.spi_inst.LSB_Address_reg[6] ));
 sg13g2_dfrbp_1 _19789_ (.CLK(net4501),
    .RESET_B(net4182),
    .D(_01117_),
    .Q_N(_09743_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[0] ));
 sg13g2_dfrbp_1 _19790_ (.CLK(net4501),
    .RESET_B(net4184),
    .D(_01118_),
    .Q_N(_09742_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[1] ));
 sg13g2_dfrbp_1 _19791_ (.CLK(net4501),
    .RESET_B(net4183),
    .D(_01119_),
    .Q_N(_09741_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[2] ));
 sg13g2_dfrbp_1 _19792_ (.CLK(net4501),
    .RESET_B(net4183),
    .D(_01120_),
    .Q_N(_09740_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[3] ));
 sg13g2_dfrbp_1 _19793_ (.CLK(net4501),
    .RESET_B(net4183),
    .D(_01121_),
    .Q_N(_09739_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[4] ));
 sg13g2_dfrbp_1 _19794_ (.CLK(net4501),
    .RESET_B(net4183),
    .D(_01122_),
    .Q_N(_09738_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[5] ));
 sg13g2_dfrbp_1 _19795_ (.CLK(net4501),
    .RESET_B(net4183),
    .D(_01123_),
    .Q_N(_09737_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[6] ));
 sg13g2_dfrbp_1 _19796_ (.CLK(net4501),
    .RESET_B(net4183),
    .D(_01124_),
    .Q_N(_09736_),
    .Q(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[7] ));
 sg13g2_dfrbp_1 _19797_ (.CLK(net4664),
    .RESET_B(net3984),
    .D(_01125_),
    .Q_N(_09735_),
    .Q(\spiking_network_top_uut.spi_inst.SPI_instruction_reg[0] ));
 sg13g2_dfrbp_1 _19798_ (.CLK(net4664),
    .RESET_B(net3984),
    .D(_01126_),
    .Q_N(_09734_),
    .Q(\spiking_network_top_uut.spi_inst.SPI_instruction_reg[1] ));
 sg13g2_dfrbp_1 _19799_ (.CLK(net4664),
    .RESET_B(net3984),
    .D(_01127_),
    .Q_N(_09733_),
    .Q(\spiking_network_top_uut.spi_inst.SPI_instruction_reg[2] ));
 sg13g2_dfrbp_1 _19800_ (.CLK(net4665),
    .RESET_B(net3985),
    .D(_01128_),
    .Q_N(_09732_),
    .Q(\spiking_network_top_uut.spi_inst.SPI_instruction_reg[3] ));
 sg13g2_dfrbp_1 _19801_ (.CLK(net4665),
    .RESET_B(net3985),
    .D(_01129_),
    .Q_N(_09731_),
    .Q(\spiking_network_top_uut.spi_inst.SPI_instruction_reg[4] ));
 sg13g2_dfrbp_1 _19802_ (.CLK(net4665),
    .RESET_B(net3985),
    .D(_01130_),
    .Q_N(_09730_),
    .Q(\spiking_network_top_uut.spi_inst.SPI_instruction_reg[5] ));
 sg13g2_dfrbp_1 _19803_ (.CLK(net4665),
    .RESET_B(net3985),
    .D(_01131_),
    .Q_N(_09729_),
    .Q(\spiking_network_top_uut.spi_inst.SPI_instruction_reg[6] ));
 sg13g2_dfrbp_1 _19804_ (.CLK(net4665),
    .RESET_B(net3985),
    .D(_01132_),
    .Q_N(_10351_),
    .Q(\spiking_network_top_uut.spi_inst.SPI_instruction_reg[7] ));
 sg13g2_dfrbp_1 _19805_ (.CLK(net4680),
    .RESET_B(net3999),
    .D(_00026_),
    .Q_N(_00029_),
    .Q(\spiking_network_top_uut.data_valid_out ));
 sg13g2_dfrbp_1 _19806_ (.CLK(_00421_),
    .RESET_B(net4025),
    .D(_00023_),
    .Q_N(_09728_),
    .Q(\spiking_network_top_uut.spi_inst.spi_slave_inst.bit_cnt[0] ));
 sg13g2_dfrbp_1 _19807_ (.CLK(_00422_),
    .RESET_B(net4024),
    .D(_00024_),
    .Q_N(_09727_),
    .Q(\spiking_network_top_uut.spi_inst.spi_slave_inst.bit_cnt[1] ));
 sg13g2_dfrbp_1 _19808_ (.CLK(_00423_),
    .RESET_B(net4015),
    .D(_00025_),
    .Q_N(_00140_),
    .Q(\spiking_network_top_uut.spi_inst.spi_slave_inst.bit_cnt[2] ));
 sg13g2_dfrbp_1 _19809_ (.CLK(net4680),
    .RESET_B(net3999),
    .D(_01133_),
    .Q_N(_09726_),
    .Q(\spiking_network_top_uut.spi_inst.spi_control_unit_inst.current_state[0] ));
 sg13g2_dfrbp_1 _19810_ (.CLK(net4680),
    .RESET_B(net3999),
    .D(_01134_),
    .Q_N(_09725_),
    .Q(\spiking_network_top_uut.spi_inst.spi_control_unit_inst.current_state[1] ));
 sg13g2_dfrbp_1 _19811_ (.CLK(net4680),
    .RESET_B(net3999),
    .D(_01135_),
    .Q_N(_00028_),
    .Q(\spiking_network_top_uut.spi_inst.spi_control_unit_inst.current_state[2] ));
 sg13g2_dfrbp_1 _19812_ (.CLK(_00424_),
    .RESET_B(net4024),
    .D(_00022_),
    .Q_N(_09724_),
    .Q(MISO));
 sg13g2_dfrbp_1 _19813_ (.CLK(net4696),
    .RESET_B(net4017),
    .D(_01136_),
    .Q_N(_09723_),
    .Q(\spiking_network_top_uut.spi_inst.SPI_instruction_reg_in[0] ));
 sg13g2_dfrbp_1 _19814_ (.CLK(net4703),
    .RESET_B(net4023),
    .D(_01137_),
    .Q_N(_09722_),
    .Q(\spiking_network_top_uut.spi_inst.SPI_instruction_reg_in[1] ));
 sg13g2_dfrbp_1 _19815_ (.CLK(net4707),
    .RESET_B(net4027),
    .D(_01138_),
    .Q_N(_09721_),
    .Q(\spiking_network_top_uut.spi_inst.SPI_instruction_reg_in[2] ));
 sg13g2_dfrbp_1 _19816_ (.CLK(net4704),
    .RESET_B(net4024),
    .D(_01139_),
    .Q_N(_09720_),
    .Q(\spiking_network_top_uut.spi_inst.SPI_instruction_reg_in[3] ));
 sg13g2_dfrbp_1 _19817_ (.CLK(net4705),
    .RESET_B(net4025),
    .D(_01140_),
    .Q_N(_09719_),
    .Q(\spiking_network_top_uut.spi_inst.SPI_instruction_reg_in[4] ));
 sg13g2_dfrbp_1 _19818_ (.CLK(net4728),
    .RESET_B(net4048),
    .D(_01141_),
    .Q_N(_09718_),
    .Q(\spiking_network_top_uut.spi_inst.SPI_instruction_reg_in[5] ));
 sg13g2_dfrbp_1 _19819_ (.CLK(net4704),
    .RESET_B(net4024),
    .D(_01142_),
    .Q_N(_09717_),
    .Q(\spiking_network_top_uut.spi_inst.SPI_instruction_reg_in[6] ));
 sg13g2_dfrbp_1 _19820_ (.CLK(net4704),
    .RESET_B(net4024),
    .D(_01143_),
    .Q_N(_10352_),
    .Q(\spiking_network_top_uut.spi_inst.SPI_instruction_reg_in[7] ));
 sg13g2_dfrbp_1 _19821_ (.CLK(net4686),
    .RESET_B(net4005),
    .D(_00019_),
    .Q_N(_10353_),
    .Q(\spiking_network_top_uut.spi_inst.SPI_address_LSB_reg_en ));
 sg13g2_dfrbp_1 _19822_ (.CLK(net4647),
    .RESET_B(net3967),
    .D(_02057_),
    .Q_N(_10354_),
    .Q(\spiking_network_top_uut.spi_inst.debug_config_ready_reg_in ));
 sg13g2_dfrbp_1 _19823_ (.CLK(net4663),
    .RESET_B(net3983),
    .D(_02058_),
    .Q_N(_10355_),
    .Q(\spiking_network_top_uut.spi_inst.clk_div_ready_reg_in ));
 sg13g2_dfrbp_1 _19824_ (.CLK(net4691),
    .RESET_B(net4010),
    .D(_00020_),
    .Q_N(_10356_),
    .Q(\spiking_network_top_uut.spi_inst.SPI_instruction_reg_en ));
 sg13g2_dfrbp_1 _19825_ (.CLK(net4647),
    .RESET_B(net3967),
    .D(_10369_),
    .Q_N(_10357_),
    .Q(\spiking_network_top_uut.spi_inst.debug_config_ready_reg_en ));
 sg13g2_dfrbp_1 _19826_ (.CLK(net4686),
    .RESET_B(net4005),
    .D(_00021_),
    .Q_N(_10358_),
    .Q(\spiking_network_top_uut.spi_inst.memory_inst.write_enable ));
 sg13g2_dfrbp_1 _19827_ (.CLK(net4663),
    .RESET_B(net3983),
    .D(_10370_),
    .Q_N(_09716_),
    .Q(\spiking_network_top_uut.spi_inst.clk_div_ready_reg_en ));
 sg13g2_dfrbp_1 _19828_ (.CLK(net4647),
    .RESET_B(net3967),
    .D(_01144_),
    .Q_N(_09715_),
    .Q(\spiking_network_top_uut.all_data_out[896] ));
 sg13g2_dfrbp_1 _19829_ (.CLK(net4647),
    .RESET_B(net3967),
    .D(_01145_),
    .Q_N(_09714_),
    .Q(\spiking_network_top_uut.all_data_out[897] ));
 sg13g2_dfrbp_1 _19830_ (.CLK(net4647),
    .RESET_B(net3967),
    .D(_01146_),
    .Q_N(_09713_),
    .Q(\spiking_network_top_uut.all_data_out[898] ));
 sg13g2_dfrbp_1 _19831_ (.CLK(net4647),
    .RESET_B(net3967),
    .D(_01147_),
    .Q_N(_09712_),
    .Q(\spiking_network_top_uut.all_data_out[899] ));
 sg13g2_dfrbp_1 _19832_ (.CLK(net4651),
    .RESET_B(net3970),
    .D(_01148_),
    .Q_N(_09711_),
    .Q(\spiking_network_top_uut.all_data_out[900] ));
 sg13g2_dfrbp_1 _19833_ (.CLK(net4652),
    .RESET_B(net3971),
    .D(_01149_),
    .Q_N(_09710_),
    .Q(\spiking_network_top_uut.all_data_out[901] ));
 sg13g2_dfrbp_1 _19834_ (.CLK(net4651),
    .RESET_B(net3970),
    .D(_01150_),
    .Q_N(_09709_),
    .Q(\spiking_network_top_uut.all_data_out[902] ));
 sg13g2_dfrbp_1 _19835_ (.CLK(net4647),
    .RESET_B(net3967),
    .D(_01151_),
    .Q_N(_09708_),
    .Q(\spiking_network_top_uut.all_data_out[903] ));
 sg13g2_dfrbp_1 _19836_ (.CLK(net4678),
    .RESET_B(net3997),
    .D(_01152_),
    .Q_N(_09707_),
    .Q(spi_instruction_done));
 sg13g2_dfrbp_1 _19837_ (.CLK(net4812),
    .RESET_B(net4133),
    .D(_01153_),
    .Q_N(_09706_),
    .Q(\spiking_network_top_uut.all_data_out[440] ));
 sg13g2_dfrbp_1 _19838_ (.CLK(net4811),
    .RESET_B(net4133),
    .D(_01154_),
    .Q_N(_00407_),
    .Q(\spiking_network_top_uut.all_data_out[441] ));
 sg13g2_dfrbp_1 _19839_ (.CLK(net4811),
    .RESET_B(net4133),
    .D(_01155_),
    .Q_N(_00337_),
    .Q(\spiking_network_top_uut.all_data_out[442] ));
 sg13g2_dfrbp_1 _19840_ (.CLK(net4758),
    .RESET_B(net4079),
    .D(_01156_),
    .Q_N(_09705_),
    .Q(\spiking_network_top_uut.all_data_out[443] ));
 sg13g2_dfrbp_1 _19841_ (.CLK(net4810),
    .RESET_B(net4130),
    .D(_01157_),
    .Q_N(_09704_),
    .Q(\spiking_network_top_uut.all_data_out[444] ));
 sg13g2_dfrbp_1 _19842_ (.CLK(net4808),
    .RESET_B(net4129),
    .D(_01158_),
    .Q_N(_00267_),
    .Q(\spiking_network_top_uut.all_data_out[445] ));
 sg13g2_dfrbp_1 _19843_ (.CLK(net4808),
    .RESET_B(net4129),
    .D(_01159_),
    .Q_N(_00197_),
    .Q(\spiking_network_top_uut.all_data_out[446] ));
 sg13g2_dfrbp_1 _19844_ (.CLK(net4750),
    .RESET_B(net4071),
    .D(_01160_),
    .Q_N(_09703_),
    .Q(\spiking_network_top_uut.all_data_out[447] ));
 sg13g2_dfrbp_1 _19845_ (.CLK(net4790),
    .RESET_B(net4112),
    .D(_01161_),
    .Q_N(_09702_),
    .Q(\spiking_network_top_uut.all_data_out[616] ));
 sg13g2_dfrbp_1 _19846_ (.CLK(net4770),
    .RESET_B(net4091),
    .D(_01162_),
    .Q_N(_00385_),
    .Q(\spiking_network_top_uut.all_data_out[617] ));
 sg13g2_dfrbp_1 _19847_ (.CLK(net4790),
    .RESET_B(net4112),
    .D(_01163_),
    .Q_N(_00315_),
    .Q(\spiking_network_top_uut.all_data_out[618] ));
 sg13g2_dfrbp_1 _19848_ (.CLK(net4774),
    .RESET_B(net4095),
    .D(_01164_),
    .Q_N(_09701_),
    .Q(\spiking_network_top_uut.all_data_out[619] ));
 sg13g2_dfrbp_1 _19849_ (.CLK(net4774),
    .RESET_B(net4095),
    .D(_01165_),
    .Q_N(_09700_),
    .Q(\spiking_network_top_uut.all_data_out[620] ));
 sg13g2_dfrbp_1 _19850_ (.CLK(net4774),
    .RESET_B(net4095),
    .D(_01166_),
    .Q_N(_00245_),
    .Q(\spiking_network_top_uut.all_data_out[621] ));
 sg13g2_dfrbp_1 _19851_ (.CLK(net4774),
    .RESET_B(net4095),
    .D(_01167_),
    .Q_N(_00175_),
    .Q(\spiking_network_top_uut.all_data_out[622] ));
 sg13g2_dfrbp_1 _19852_ (.CLK(net4793),
    .RESET_B(net4115),
    .D(_01168_),
    .Q_N(_09699_),
    .Q(\spiking_network_top_uut.all_data_out[623] ));
 sg13g2_dfrbp_1 _19853_ (.CLK(net4780),
    .RESET_B(net4102),
    .D(_01169_),
    .Q_N(_09698_),
    .Q(\spiking_network_top_uut.all_data_out[432] ));
 sg13g2_dfrbp_1 _19854_ (.CLK(net4780),
    .RESET_B(net4101),
    .D(_01170_),
    .Q_N(_00408_),
    .Q(\spiking_network_top_uut.all_data_out[433] ));
 sg13g2_dfrbp_1 _19855_ (.CLK(net4780),
    .RESET_B(net4101),
    .D(_01171_),
    .Q_N(_00338_),
    .Q(\spiking_network_top_uut.all_data_out[434] ));
 sg13g2_dfrbp_1 _19856_ (.CLK(net4782),
    .RESET_B(net4102),
    .D(_01172_),
    .Q_N(_09697_),
    .Q(\spiking_network_top_uut.all_data_out[435] ));
 sg13g2_dfrbp_1 _19857_ (.CLK(net4752),
    .RESET_B(net4073),
    .D(_01173_),
    .Q_N(_09696_),
    .Q(\spiking_network_top_uut.all_data_out[436] ));
 sg13g2_dfrbp_1 _19858_ (.CLK(net4752),
    .RESET_B(net4073),
    .D(_01174_),
    .Q_N(_00268_),
    .Q(\spiking_network_top_uut.all_data_out[437] ));
 sg13g2_dfrbp_1 _19859_ (.CLK(net4753),
    .RESET_B(net4074),
    .D(_01175_),
    .Q_N(_00198_),
    .Q(\spiking_network_top_uut.all_data_out[438] ));
 sg13g2_dfrbp_1 _19860_ (.CLK(net4752),
    .RESET_B(net4073),
    .D(_01176_),
    .Q_N(_09695_),
    .Q(\spiking_network_top_uut.all_data_out[439] ));
 sg13g2_dfrbp_1 _19861_ (.CLK(net4770),
    .RESET_B(net4091),
    .D(_01177_),
    .Q_N(_09694_),
    .Q(\spiking_network_top_uut.all_data_out[680] ));
 sg13g2_dfrbp_1 _19862_ (.CLK(net4771),
    .RESET_B(net4092),
    .D(_01178_),
    .Q_N(_00377_),
    .Q(\spiking_network_top_uut.all_data_out[681] ));
 sg13g2_dfrbp_1 _19863_ (.CLK(net4770),
    .RESET_B(net4091),
    .D(_01179_),
    .Q_N(_00307_),
    .Q(\spiking_network_top_uut.all_data_out[682] ));
 sg13g2_dfrbp_1 _19864_ (.CLK(net4768),
    .RESET_B(net4089),
    .D(_01180_),
    .Q_N(_09693_),
    .Q(\spiking_network_top_uut.all_data_out[683] ));
 sg13g2_dfrbp_1 _19865_ (.CLK(net4784),
    .RESET_B(net4106),
    .D(_01181_),
    .Q_N(_09692_),
    .Q(\spiking_network_top_uut.all_data_out[684] ));
 sg13g2_dfrbp_1 _19866_ (.CLK(net4778),
    .RESET_B(net4099),
    .D(_01182_),
    .Q_N(_00237_),
    .Q(\spiking_network_top_uut.all_data_out[685] ));
 sg13g2_dfrbp_1 _19867_ (.CLK(net4778),
    .RESET_B(net4099),
    .D(_01183_),
    .Q_N(_00167_),
    .Q(\spiking_network_top_uut.all_data_out[686] ));
 sg13g2_dfrbp_1 _19868_ (.CLK(net4778),
    .RESET_B(net4099),
    .D(_01184_),
    .Q_N(_09691_),
    .Q(\spiking_network_top_uut.all_data_out[687] ));
 sg13g2_dfrbp_1 _19869_ (.CLK(net4789),
    .RESET_B(net4111),
    .D(_01185_),
    .Q_N(_09690_),
    .Q(\spiking_network_top_uut.all_data_out[424] ));
 sg13g2_dfrbp_1 _19870_ (.CLK(net4789),
    .RESET_B(net4111),
    .D(_01186_),
    .Q_N(_00409_),
    .Q(\spiking_network_top_uut.all_data_out[425] ));
 sg13g2_dfrbp_1 _19871_ (.CLK(net4789),
    .RESET_B(net4111),
    .D(_01187_),
    .Q_N(_00339_),
    .Q(\spiking_network_top_uut.all_data_out[426] ));
 sg13g2_dfrbp_1 _19872_ (.CLK(net4772),
    .RESET_B(net4093),
    .D(_01188_),
    .Q_N(_09689_),
    .Q(\spiking_network_top_uut.all_data_out[427] ));
 sg13g2_dfrbp_1 _19873_ (.CLK(net4795),
    .RESET_B(net4117),
    .D(_01189_),
    .Q_N(_09688_),
    .Q(\spiking_network_top_uut.all_data_out[428] ));
 sg13g2_dfrbp_1 _19874_ (.CLK(net4795),
    .RESET_B(net4119),
    .D(_01190_),
    .Q_N(_00269_),
    .Q(\spiking_network_top_uut.all_data_out[429] ));
 sg13g2_dfrbp_1 _19875_ (.CLK(net4795),
    .RESET_B(net4123),
    .D(_01191_),
    .Q_N(_00199_),
    .Q(\spiking_network_top_uut.all_data_out[430] ));
 sg13g2_dfrbp_1 _19876_ (.CLK(net4772),
    .RESET_B(net4093),
    .D(_01192_),
    .Q_N(_09687_),
    .Q(\spiking_network_top_uut.all_data_out[431] ));
 sg13g2_dfrbp_1 _19877_ (.CLK(net4793),
    .RESET_B(net4115),
    .D(_01193_),
    .Q_N(_09686_),
    .Q(\spiking_network_top_uut.all_data_out[552] ));
 sg13g2_dfrbp_1 _19878_ (.CLK(net4791),
    .RESET_B(net4113),
    .D(_01194_),
    .Q_N(_00393_),
    .Q(\spiking_network_top_uut.all_data_out[553] ));
 sg13g2_dfrbp_1 _19879_ (.CLK(net4791),
    .RESET_B(net4113),
    .D(_01195_),
    .Q_N(_00323_),
    .Q(\spiking_network_top_uut.all_data_out[554] ));
 sg13g2_dfrbp_1 _19880_ (.CLK(net4773),
    .RESET_B(net4094),
    .D(_01196_),
    .Q_N(_09685_),
    .Q(\spiking_network_top_uut.all_data_out[555] ));
 sg13g2_dfrbp_1 _19881_ (.CLK(net4797),
    .RESET_B(net4118),
    .D(_01197_),
    .Q_N(_09684_),
    .Q(\spiking_network_top_uut.all_data_out[556] ));
 sg13g2_dfrbp_1 _19882_ (.CLK(net4799),
    .RESET_B(net4119),
    .D(_01198_),
    .Q_N(_00253_),
    .Q(\spiking_network_top_uut.all_data_out[557] ));
 sg13g2_dfrbp_1 _19883_ (.CLK(net4800),
    .RESET_B(net4122),
    .D(_01199_),
    .Q_N(_00183_),
    .Q(\spiking_network_top_uut.all_data_out[558] ));
 sg13g2_dfrbp_1 _19884_ (.CLK(net4793),
    .RESET_B(net4115),
    .D(_01200_),
    .Q_N(_09683_),
    .Q(\spiking_network_top_uut.all_data_out[559] ));
 sg13g2_dfrbp_1 _19885_ (.CLK(net4783),
    .RESET_B(net4105),
    .D(_01201_),
    .Q_N(_09682_),
    .Q(\spiking_network_top_uut.all_data_out[416] ));
 sg13g2_dfrbp_1 _19886_ (.CLK(net4785),
    .RESET_B(net4107),
    .D(_01202_),
    .Q_N(_00410_),
    .Q(\spiking_network_top_uut.all_data_out[417] ));
 sg13g2_dfrbp_1 _19887_ (.CLK(net4786),
    .RESET_B(net4108),
    .D(_01203_),
    .Q_N(_00340_),
    .Q(\spiking_network_top_uut.all_data_out[418] ));
 sg13g2_dfrbp_1 _19888_ (.CLK(net4785),
    .RESET_B(net4107),
    .D(_01204_),
    .Q_N(_09681_),
    .Q(\spiking_network_top_uut.all_data_out[419] ));
 sg13g2_dfrbp_1 _19889_ (.CLK(net4783),
    .RESET_B(net4105),
    .D(_01205_),
    .Q_N(_09680_),
    .Q(\spiking_network_top_uut.all_data_out[420] ));
 sg13g2_dfrbp_1 _19890_ (.CLK(net4803),
    .RESET_B(net4125),
    .D(_01206_),
    .Q_N(_00270_),
    .Q(\spiking_network_top_uut.all_data_out[421] ));
 sg13g2_dfrbp_1 _19891_ (.CLK(net4803),
    .RESET_B(net4125),
    .D(_01207_),
    .Q_N(_00200_),
    .Q(\spiking_network_top_uut.all_data_out[422] ));
 sg13g2_dfrbp_1 _19892_ (.CLK(net4785),
    .RESET_B(net4107),
    .D(_01208_),
    .Q_N(_09679_),
    .Q(\spiking_network_top_uut.all_data_out[423] ));
 sg13g2_dfrbp_1 _19893_ (.CLK(net4746),
    .RESET_B(net4067),
    .D(_01209_),
    .Q_N(_09678_),
    .Q(\spiking_network_top_uut.all_data_out[688] ));
 sg13g2_dfrbp_1 _19894_ (.CLK(net4744),
    .RESET_B(net4065),
    .D(_01210_),
    .Q_N(_00376_),
    .Q(\spiking_network_top_uut.all_data_out[689] ));
 sg13g2_dfrbp_1 _19895_ (.CLK(net4740),
    .RESET_B(net4061),
    .D(_01211_),
    .Q_N(_00306_),
    .Q(\spiking_network_top_uut.all_data_out[690] ));
 sg13g2_dfrbp_1 _19896_ (.CLK(net4740),
    .RESET_B(net4061),
    .D(_01212_),
    .Q_N(_09677_),
    .Q(\spiking_network_top_uut.all_data_out[691] ));
 sg13g2_dfrbp_1 _19897_ (.CLK(net4777),
    .RESET_B(net4098),
    .D(_01213_),
    .Q_N(_09676_),
    .Q(\spiking_network_top_uut.all_data_out[692] ));
 sg13g2_dfrbp_1 _19898_ (.CLK(net4767),
    .RESET_B(net4088),
    .D(_01214_),
    .Q_N(_00236_),
    .Q(\spiking_network_top_uut.all_data_out[693] ));
 sg13g2_dfrbp_1 _19899_ (.CLK(net4766),
    .RESET_B(net4087),
    .D(_01215_),
    .Q_N(_00166_),
    .Q(\spiking_network_top_uut.all_data_out[694] ));
 sg13g2_dfrbp_1 _19900_ (.CLK(net4744),
    .RESET_B(net4065),
    .D(_01216_),
    .Q_N(_09675_),
    .Q(\spiking_network_top_uut.all_data_out[695] ));
 sg13g2_dfrbp_1 _19901_ (.CLK(net4809),
    .RESET_B(net4131),
    .D(_01217_),
    .Q_N(_09674_),
    .Q(\spiking_network_top_uut.all_data_out[408] ));
 sg13g2_dfrbp_1 _19902_ (.CLK(net4809),
    .RESET_B(net4130),
    .D(_01218_),
    .Q_N(_00411_),
    .Q(\spiking_network_top_uut.all_data_out[409] ));
 sg13g2_dfrbp_1 _19903_ (.CLK(net4809),
    .RESET_B(net4130),
    .D(_01219_),
    .Q_N(_00341_),
    .Q(\spiking_network_top_uut.all_data_out[410] ));
 sg13g2_dfrbp_1 _19904_ (.CLK(net4755),
    .RESET_B(net4076),
    .D(_01220_),
    .Q_N(_09673_),
    .Q(\spiking_network_top_uut.all_data_out[411] ));
 sg13g2_dfrbp_1 _19905_ (.CLK(net4808),
    .RESET_B(net4129),
    .D(_01221_),
    .Q_N(_09672_),
    .Q(\spiking_network_top_uut.all_data_out[412] ));
 sg13g2_dfrbp_1 _19906_ (.CLK(net4810),
    .RESET_B(net4131),
    .D(_01222_),
    .Q_N(_00271_),
    .Q(\spiking_network_top_uut.all_data_out[413] ));
 sg13g2_dfrbp_1 _19907_ (.CLK(net4798),
    .RESET_B(net4120),
    .D(_01223_),
    .Q_N(_00201_),
    .Q(\spiking_network_top_uut.all_data_out[414] ));
 sg13g2_dfrbp_1 _19908_ (.CLK(net4755),
    .RESET_B(net4076),
    .D(_01224_),
    .Q_N(_09671_),
    .Q(\spiking_network_top_uut.all_data_out[415] ));
 sg13g2_dfrbp_1 _19909_ (.CLK(net4770),
    .RESET_B(net4091),
    .D(_01225_),
    .Q_N(_09670_),
    .Q(\spiking_network_top_uut.all_data_out[584] ));
 sg13g2_dfrbp_1 _19910_ (.CLK(net4770),
    .RESET_B(net4091),
    .D(_01226_),
    .Q_N(_00389_),
    .Q(\spiking_network_top_uut.all_data_out[585] ));
 sg13g2_dfrbp_1 _19911_ (.CLK(net4770),
    .RESET_B(net4091),
    .D(_01227_),
    .Q_N(_00319_),
    .Q(\spiking_network_top_uut.all_data_out[586] ));
 sg13g2_dfrbp_1 _19912_ (.CLK(net4775),
    .RESET_B(net4096),
    .D(_01228_),
    .Q_N(_09669_),
    .Q(\spiking_network_top_uut.all_data_out[587] ));
 sg13g2_dfrbp_1 _19913_ (.CLK(net4772),
    .RESET_B(net4093),
    .D(_01229_),
    .Q_N(_09668_),
    .Q(\spiking_network_top_uut.all_data_out[588] ));
 sg13g2_dfrbp_1 _19914_ (.CLK(net4775),
    .RESET_B(net4093),
    .D(_01230_),
    .Q_N(_00249_),
    .Q(\spiking_network_top_uut.all_data_out[589] ));
 sg13g2_dfrbp_1 _19915_ (.CLK(net4772),
    .RESET_B(net4093),
    .D(_01231_),
    .Q_N(_00179_),
    .Q(\spiking_network_top_uut.all_data_out[590] ));
 sg13g2_dfrbp_1 _19916_ (.CLK(net4774),
    .RESET_B(net4095),
    .D(_01232_),
    .Q_N(_09667_),
    .Q(\spiking_network_top_uut.all_data_out[591] ));
 sg13g2_dfrbp_1 _19917_ (.CLK(net4780),
    .RESET_B(net4101),
    .D(_01233_),
    .Q_N(_09666_),
    .Q(\spiking_network_top_uut.all_data_out[400] ));
 sg13g2_dfrbp_1 _19918_ (.CLK(net4778),
    .RESET_B(net4101),
    .D(_01234_),
    .Q_N(_00412_),
    .Q(\spiking_network_top_uut.all_data_out[401] ));
 sg13g2_dfrbp_1 _19919_ (.CLK(net4779),
    .RESET_B(net4100),
    .D(_01235_),
    .Q_N(_00342_),
    .Q(\spiking_network_top_uut.all_data_out[402] ));
 sg13g2_dfrbp_1 _19920_ (.CLK(net4758),
    .RESET_B(net4079),
    .D(_01236_),
    .Q_N(_09665_),
    .Q(\spiking_network_top_uut.all_data_out[403] ));
 sg13g2_dfrbp_1 _19921_ (.CLK(net4762),
    .RESET_B(net4083),
    .D(_01237_),
    .Q_N(_09664_),
    .Q(\spiking_network_top_uut.all_data_out[404] ));
 sg13g2_dfrbp_1 _19922_ (.CLK(net4760),
    .RESET_B(net4081),
    .D(_01238_),
    .Q_N(_00272_),
    .Q(\spiking_network_top_uut.all_data_out[405] ));
 sg13g2_dfrbp_1 _19923_ (.CLK(net4760),
    .RESET_B(net4081),
    .D(_01239_),
    .Q_N(_00202_),
    .Q(\spiking_network_top_uut.all_data_out[406] ));
 sg13g2_dfrbp_1 _19924_ (.CLK(net4758),
    .RESET_B(net4079),
    .D(_01240_),
    .Q_N(_09663_),
    .Q(\spiking_network_top_uut.all_data_out[407] ));
 sg13g2_dfrbp_1 _19925_ (.CLK(net4715),
    .RESET_B(net4035),
    .D(_01241_),
    .Q_N(_09662_),
    .Q(\spiking_network_top_uut.all_data_out[696] ));
 sg13g2_dfrbp_1 _19926_ (.CLK(net4715),
    .RESET_B(net4035),
    .D(_01242_),
    .Q_N(_00375_),
    .Q(\spiking_network_top_uut.all_data_out[697] ));
 sg13g2_dfrbp_1 _19927_ (.CLK(net4710),
    .RESET_B(net4030),
    .D(_01243_),
    .Q_N(_00305_),
    .Q(\spiking_network_top_uut.all_data_out[698] ));
 sg13g2_dfrbp_1 _19928_ (.CLK(net4716),
    .RESET_B(net4036),
    .D(_01244_),
    .Q_N(_09661_),
    .Q(\spiking_network_top_uut.all_data_out[699] ));
 sg13g2_dfrbp_1 _19929_ (.CLK(net4718),
    .RESET_B(net4037),
    .D(_01245_),
    .Q_N(_09660_),
    .Q(\spiking_network_top_uut.all_data_out[700] ));
 sg13g2_dfrbp_1 _19930_ (.CLK(net4739),
    .RESET_B(net4060),
    .D(_01246_),
    .Q_N(_00235_),
    .Q(\spiking_network_top_uut.all_data_out[701] ));
 sg13g2_dfrbp_1 _19931_ (.CLK(net4739),
    .RESET_B(net4060),
    .D(_01247_),
    .Q_N(_00165_),
    .Q(\spiking_network_top_uut.all_data_out[702] ));
 sg13g2_dfrbp_1 _19932_ (.CLK(net4717),
    .RESET_B(net4038),
    .D(_01248_),
    .Q_N(_09659_),
    .Q(\spiking_network_top_uut.all_data_out[703] ));
 sg13g2_dfrbp_1 _19933_ (.CLK(net4789),
    .RESET_B(net4111),
    .D(_01249_),
    .Q_N(_09658_),
    .Q(\spiking_network_top_uut.all_data_out[392] ));
 sg13g2_dfrbp_1 _19934_ (.CLK(net4791),
    .RESET_B(net4113),
    .D(_01250_),
    .Q_N(_00413_),
    .Q(\spiking_network_top_uut.all_data_out[393] ));
 sg13g2_dfrbp_1 _19935_ (.CLK(net4790),
    .RESET_B(net4112),
    .D(_01251_),
    .Q_N(_00343_),
    .Q(\spiking_network_top_uut.all_data_out[394] ));
 sg13g2_dfrbp_1 _19936_ (.CLK(net4772),
    .RESET_B(net4093),
    .D(_01252_),
    .Q_N(_09657_),
    .Q(\spiking_network_top_uut.all_data_out[395] ));
 sg13g2_dfrbp_1 _19937_ (.CLK(net4795),
    .RESET_B(net4117),
    .D(_01253_),
    .Q_N(_09656_),
    .Q(\spiking_network_top_uut.all_data_out[396] ));
 sg13g2_dfrbp_1 _19938_ (.CLK(net4797),
    .RESET_B(net4118),
    .D(_01254_),
    .Q_N(_00273_),
    .Q(\spiking_network_top_uut.all_data_out[397] ));
 sg13g2_dfrbp_1 _19939_ (.CLK(net4799),
    .RESET_B(net4119),
    .D(_01255_),
    .Q_N(_00203_),
    .Q(\spiking_network_top_uut.all_data_out[398] ));
 sg13g2_dfrbp_1 _19940_ (.CLK(net4793),
    .RESET_B(net4115),
    .D(_01256_),
    .Q_N(_09655_),
    .Q(\spiking_network_top_uut.all_data_out[399] ));
 sg13g2_dfrbp_1 _19941_ (.CLK(net4805),
    .RESET_B(net4127),
    .D(_01257_),
    .Q_N(_09654_),
    .Q(\spiking_network_top_uut.all_data_out[544] ));
 sg13g2_dfrbp_1 _19942_ (.CLK(net4786),
    .RESET_B(net4108),
    .D(_01258_),
    .Q_N(_00394_),
    .Q(\spiking_network_top_uut.all_data_out[545] ));
 sg13g2_dfrbp_1 _19943_ (.CLK(net4787),
    .RESET_B(net4105),
    .D(_01259_),
    .Q_N(_00324_),
    .Q(\spiking_network_top_uut.all_data_out[546] ));
 sg13g2_dfrbp_1 _19944_ (.CLK(net4783),
    .RESET_B(net4109),
    .D(_01260_),
    .Q_N(_09653_),
    .Q(\spiking_network_top_uut.all_data_out[547] ));
 sg13g2_dfrbp_1 _19945_ (.CLK(net4802),
    .RESET_B(net4124),
    .D(_01261_),
    .Q_N(_09652_),
    .Q(\spiking_network_top_uut.all_data_out[548] ));
 sg13g2_dfrbp_1 _19946_ (.CLK(net4802),
    .RESET_B(net4124),
    .D(_01262_),
    .Q_N(_00254_),
    .Q(\spiking_network_top_uut.all_data_out[549] ));
 sg13g2_dfrbp_1 _19947_ (.CLK(net4802),
    .RESET_B(net4124),
    .D(_01263_),
    .Q_N(_00184_),
    .Q(\spiking_network_top_uut.all_data_out[550] ));
 sg13g2_dfrbp_1 _19948_ (.CLK(net4783),
    .RESET_B(net4105),
    .D(_01264_),
    .Q_N(_09651_),
    .Q(\spiking_network_top_uut.all_data_out[551] ));
 sg13g2_dfrbp_1 _19949_ (.CLK(net4805),
    .RESET_B(net4128),
    .D(_01265_),
    .Q_N(_09650_),
    .Q(\spiking_network_top_uut.all_data_out[384] ));
 sg13g2_dfrbp_1 _19950_ (.CLK(net4805),
    .RESET_B(net4127),
    .D(_01266_),
    .Q_N(_00414_),
    .Q(\spiking_network_top_uut.all_data_out[385] ));
 sg13g2_dfrbp_1 _19951_ (.CLK(net4805),
    .RESET_B(net4127),
    .D(_01267_),
    .Q_N(_00344_),
    .Q(\spiking_network_top_uut.all_data_out[386] ));
 sg13g2_dfrbp_1 _19952_ (.CLK(net4727),
    .RESET_B(net4047),
    .D(_01268_),
    .Q_N(_09649_),
    .Q(\spiking_network_top_uut.all_data_out[387] ));
 sg13g2_dfrbp_1 _19953_ (.CLK(net4791),
    .RESET_B(net4114),
    .D(_01269_),
    .Q_N(_09648_),
    .Q(\spiking_network_top_uut.all_data_out[388] ));
 sg13g2_dfrbp_1 _19954_ (.CLK(net4792),
    .RESET_B(net4113),
    .D(_01270_),
    .Q_N(_00274_),
    .Q(\spiking_network_top_uut.all_data_out[389] ));
 sg13g2_dfrbp_1 _19955_ (.CLK(net4792),
    .RESET_B(net4114),
    .D(_01271_),
    .Q_N(_00204_),
    .Q(\spiking_network_top_uut.all_data_out[390] ));
 sg13g2_dfrbp_1 _19956_ (.CLK(net4725),
    .RESET_B(net4045),
    .D(_01272_),
    .Q_N(_09647_),
    .Q(\spiking_network_top_uut.all_data_out[391] ));
 sg13g2_dfrbp_1 _19957_ (.CLK(net4680),
    .RESET_B(net3999),
    .D(_01273_),
    .Q_N(_09646_),
    .Q(\spiking_network_top_uut.all_data_out[704] ));
 sg13g2_dfrbp_1 _19958_ (.CLK(net4683),
    .RESET_B(net4002),
    .D(_01274_),
    .Q_N(_00374_),
    .Q(\spiking_network_top_uut.all_data_out[705] ));
 sg13g2_dfrbp_1 _19959_ (.CLK(net4681),
    .RESET_B(net4000),
    .D(_01275_),
    .Q_N(_00304_),
    .Q(\spiking_network_top_uut.all_data_out[706] ));
 sg13g2_dfrbp_1 _19960_ (.CLK(net4693),
    .RESET_B(net4017),
    .D(_01276_),
    .Q_N(_09645_),
    .Q(\spiking_network_top_uut.all_data_out[707] ));
 sg13g2_dfrbp_1 _19961_ (.CLK(net4693),
    .RESET_B(net4013),
    .D(_01277_),
    .Q_N(_09644_),
    .Q(\spiking_network_top_uut.all_data_out[708] ));
 sg13g2_dfrbp_1 _19962_ (.CLK(net4674),
    .RESET_B(net3994),
    .D(_01278_),
    .Q_N(_00234_),
    .Q(\spiking_network_top_uut.all_data_out[709] ));
 sg13g2_dfrbp_1 _19963_ (.CLK(net4692),
    .RESET_B(net4011),
    .D(_01279_),
    .Q_N(_00164_),
    .Q(\spiking_network_top_uut.all_data_out[710] ));
 sg13g2_dfrbp_1 _19964_ (.CLK(net4674),
    .RESET_B(net3993),
    .D(_01280_),
    .Q_N(_09643_),
    .Q(\spiking_network_top_uut.all_data_out[711] ));
 sg13g2_dfrbp_1 _19965_ (.CLK(net4811),
    .RESET_B(net4133),
    .D(_01281_),
    .Q_N(_09642_),
    .Q(\spiking_network_top_uut.all_data_out[376] ));
 sg13g2_dfrbp_1 _19966_ (.CLK(net4811),
    .RESET_B(net4133),
    .D(_01282_),
    .Q_N(_00415_),
    .Q(\spiking_network_top_uut.all_data_out[377] ));
 sg13g2_dfrbp_1 _19967_ (.CLK(net4811),
    .RESET_B(net4133),
    .D(_01283_),
    .Q_N(_00345_),
    .Q(\spiking_network_top_uut.all_data_out[378] ));
 sg13g2_dfrbp_1 _19968_ (.CLK(net4729),
    .RESET_B(net4049),
    .D(_01284_),
    .Q_N(_09641_),
    .Q(\spiking_network_top_uut.all_data_out[379] ));
 sg13g2_dfrbp_1 _19969_ (.CLK(net4807),
    .RESET_B(net4132),
    .D(_01285_),
    .Q_N(_09640_),
    .Q(\spiking_network_top_uut.all_data_out[380] ));
 sg13g2_dfrbp_1 _19970_ (.CLK(net4807),
    .RESET_B(net4132),
    .D(_01286_),
    .Q_N(_00275_),
    .Q(\spiking_network_top_uut.all_data_out[381] ));
 sg13g2_dfrbp_1 _19971_ (.CLK(net4808),
    .RESET_B(net4129),
    .D(_01287_),
    .Q_N(_00205_),
    .Q(\spiking_network_top_uut.all_data_out[382] ));
 sg13g2_dfrbp_1 _19972_ (.CLK(net4729),
    .RESET_B(net4049),
    .D(_01288_),
    .Q_N(_09639_),
    .Q(\spiking_network_top_uut.all_data_out[383] ));
 sg13g2_dfrbp_1 _19973_ (.CLK(net4766),
    .RESET_B(net4087),
    .D(_01289_),
    .Q_N(_09638_),
    .Q(\spiking_network_top_uut.all_data_out[624] ));
 sg13g2_dfrbp_1 _19974_ (.CLK(net4766),
    .RESET_B(net4087),
    .D(_01290_),
    .Q_N(_00384_),
    .Q(\spiking_network_top_uut.all_data_out[625] ));
 sg13g2_dfrbp_1 _19975_ (.CLK(net4766),
    .RESET_B(net4087),
    .D(_01291_),
    .Q_N(_00314_),
    .Q(\spiking_network_top_uut.all_data_out[626] ));
 sg13g2_dfrbp_1 _19976_ (.CLK(net4748),
    .RESET_B(net4069),
    .D(_01292_),
    .Q_N(_09637_),
    .Q(\spiking_network_top_uut.all_data_out[627] ));
 sg13g2_dfrbp_1 _19977_ (.CLK(net4765),
    .RESET_B(net4086),
    .D(_01293_),
    .Q_N(_09636_),
    .Q(\spiking_network_top_uut.all_data_out[628] ));
 sg13g2_dfrbp_1 _19978_ (.CLK(net4765),
    .RESET_B(net4086),
    .D(_01294_),
    .Q_N(_00244_),
    .Q(\spiking_network_top_uut.all_data_out[629] ));
 sg13g2_dfrbp_1 _19979_ (.CLK(net4765),
    .RESET_B(net4086),
    .D(_01295_),
    .Q_N(_00174_),
    .Q(\spiking_network_top_uut.all_data_out[630] ));
 sg13g2_dfrbp_1 _19980_ (.CLK(net4747),
    .RESET_B(net4068),
    .D(_01296_),
    .Q_N(_09635_),
    .Q(\spiking_network_top_uut.all_data_out[631] ));
 sg13g2_dfrbp_1 _19981_ (.CLK(net4778),
    .RESET_B(net4099),
    .D(_01297_),
    .Q_N(_09634_),
    .Q(\spiking_network_top_uut.all_data_out[368] ));
 sg13g2_dfrbp_1 _19982_ (.CLK(net4779),
    .RESET_B(net4101),
    .D(_01298_),
    .Q_N(_00416_),
    .Q(\spiking_network_top_uut.all_data_out[369] ));
 sg13g2_dfrbp_1 _19983_ (.CLK(net4778),
    .RESET_B(net4099),
    .D(_01299_),
    .Q_N(_00346_),
    .Q(\spiking_network_top_uut.all_data_out[370] ));
 sg13g2_dfrbp_1 _19984_ (.CLK(net4780),
    .RESET_B(net4101),
    .D(_01300_),
    .Q_N(_09633_),
    .Q(\spiking_network_top_uut.all_data_out[371] ));
 sg13g2_dfrbp_1 _19985_ (.CLK(net4760),
    .RESET_B(net4081),
    .D(_01301_),
    .Q_N(_09632_),
    .Q(\spiking_network_top_uut.all_data_out[372] ));
 sg13g2_dfrbp_1 _19986_ (.CLK(net4760),
    .RESET_B(net4081),
    .D(_01302_),
    .Q_N(_00276_),
    .Q(\spiking_network_top_uut.all_data_out[373] ));
 sg13g2_dfrbp_1 _19987_ (.CLK(net4760),
    .RESET_B(net4081),
    .D(_01303_),
    .Q_N(_00206_),
    .Q(\spiking_network_top_uut.all_data_out[374] ));
 sg13g2_dfrbp_1 _19988_ (.CLK(net4762),
    .RESET_B(net4083),
    .D(_01304_),
    .Q_N(_09631_),
    .Q(\spiking_network_top_uut.all_data_out[375] ));
 sg13g2_dfrbp_1 _19989_ (.CLK(net4790),
    .RESET_B(net4112),
    .D(_01305_),
    .Q_N(_09630_),
    .Q(\spiking_network_top_uut.all_data_out[712] ));
 sg13g2_dfrbp_1 _19990_ (.CLK(net4776),
    .RESET_B(net4097),
    .D(_01306_),
    .Q_N(_00373_),
    .Q(\spiking_network_top_uut.all_data_out[713] ));
 sg13g2_dfrbp_1 _19991_ (.CLK(net4773),
    .RESET_B(net4094),
    .D(_01307_),
    .Q_N(_00303_),
    .Q(\spiking_network_top_uut.all_data_out[714] ));
 sg13g2_dfrbp_1 _19992_ (.CLK(net4748),
    .RESET_B(net4068),
    .D(_01308_),
    .Q_N(_09629_),
    .Q(\spiking_network_top_uut.all_data_out[715] ));
 sg13g2_dfrbp_1 _19993_ (.CLK(net4784),
    .RESET_B(net4106),
    .D(_01309_),
    .Q_N(_09628_),
    .Q(\spiking_network_top_uut.all_data_out[716] ));
 sg13g2_dfrbp_1 _19994_ (.CLK(net4768),
    .RESET_B(net4099),
    .D(_01310_),
    .Q_N(_00233_),
    .Q(\spiking_network_top_uut.all_data_out[717] ));
 sg13g2_dfrbp_1 _19995_ (.CLK(net4779),
    .RESET_B(net4100),
    .D(_01311_),
    .Q_N(_00163_),
    .Q(\spiking_network_top_uut.all_data_out[718] ));
 sg13g2_dfrbp_1 _19996_ (.CLK(net4757),
    .RESET_B(net4078),
    .D(_01312_),
    .Q_N(_09627_),
    .Q(\spiking_network_top_uut.all_data_out[719] ));
 sg13g2_dfrbp_1 _19997_ (.CLK(net4792),
    .RESET_B(net4114),
    .D(_01313_),
    .Q_N(_09626_),
    .Q(\spiking_network_top_uut.all_data_out[360] ));
 sg13g2_dfrbp_1 _19998_ (.CLK(net4800),
    .RESET_B(net4122),
    .D(_01314_),
    .Q_N(_00417_),
    .Q(\spiking_network_top_uut.all_data_out[361] ));
 sg13g2_dfrbp_1 _19999_ (.CLK(net4791),
    .RESET_B(net4113),
    .D(_01315_),
    .Q_N(_00347_),
    .Q(\spiking_network_top_uut.all_data_out[362] ));
 sg13g2_dfrbp_1 _20000_ (.CLK(net4773),
    .RESET_B(net4094),
    .D(_01316_),
    .Q_N(_09625_),
    .Q(\spiking_network_top_uut.all_data_out[363] ));
 sg13g2_dfrbp_1 _20001_ (.CLK(net4797),
    .RESET_B(net4118),
    .D(_01317_),
    .Q_N(_09624_),
    .Q(\spiking_network_top_uut.all_data_out[364] ));
 sg13g2_dfrbp_1 _20002_ (.CLK(net4799),
    .RESET_B(net4119),
    .D(_01318_),
    .Q_N(_00277_),
    .Q(\spiking_network_top_uut.all_data_out[365] ));
 sg13g2_dfrbp_1 _20003_ (.CLK(net4797),
    .RESET_B(net4118),
    .D(_01319_),
    .Q_N(_00207_),
    .Q(\spiking_network_top_uut.all_data_out[366] ));
 sg13g2_dfrbp_1 _20004_ (.CLK(net4793),
    .RESET_B(net4115),
    .D(_01320_),
    .Q_N(_09623_),
    .Q(\spiking_network_top_uut.all_data_out[367] ));
 sg13g2_dfrbp_1 _20005_ (.CLK(net4811),
    .RESET_B(net4134),
    .D(_01321_),
    .Q_N(_09622_),
    .Q(\spiking_network_top_uut.all_data_out[536] ));
 sg13g2_dfrbp_1 _20006_ (.CLK(net4809),
    .RESET_B(net4130),
    .D(_01322_),
    .Q_N(_00395_),
    .Q(\spiking_network_top_uut.all_data_out[537] ));
 sg13g2_dfrbp_1 _20007_ (.CLK(net4810),
    .RESET_B(net4131),
    .D(_01323_),
    .Q_N(_00325_),
    .Q(\spiking_network_top_uut.all_data_out[538] ));
 sg13g2_dfrbp_1 _20008_ (.CLK(net4755),
    .RESET_B(net4076),
    .D(_01324_),
    .Q_N(_09621_),
    .Q(\spiking_network_top_uut.all_data_out[539] ));
 sg13g2_dfrbp_1 _20009_ (.CLK(net4798),
    .RESET_B(net4120),
    .D(_01325_),
    .Q_N(_09620_),
    .Q(\spiking_network_top_uut.all_data_out[540] ));
 sg13g2_dfrbp_1 _20010_ (.CLK(net4798),
    .RESET_B(net4121),
    .D(_01326_),
    .Q_N(_00255_),
    .Q(\spiking_network_top_uut.all_data_out[541] ));
 sg13g2_dfrbp_1 _20011_ (.CLK(net4798),
    .RESET_B(net4120),
    .D(_01327_),
    .Q_N(_00185_),
    .Q(\spiking_network_top_uut.all_data_out[542] ));
 sg13g2_dfrbp_1 _20012_ (.CLK(net4755),
    .RESET_B(net4076),
    .D(_01328_),
    .Q_N(_09619_),
    .Q(\spiking_network_top_uut.all_data_out[543] ));
 sg13g2_dfrbp_1 _20013_ (.CLK(net4805),
    .RESET_B(net4127),
    .D(_01329_),
    .Q_N(_09618_),
    .Q(\spiking_network_top_uut.all_data_out[352] ));
 sg13g2_dfrbp_1 _20014_ (.CLK(net4786),
    .RESET_B(net4108),
    .D(_01330_),
    .Q_N(_00418_),
    .Q(\spiking_network_top_uut.all_data_out[353] ));
 sg13g2_dfrbp_1 _20015_ (.CLK(net4786),
    .RESET_B(net4107),
    .D(_01331_),
    .Q_N(_00348_),
    .Q(\spiking_network_top_uut.all_data_out[354] ));
 sg13g2_dfrbp_1 _20016_ (.CLK(net4780),
    .RESET_B(net4101),
    .D(_01332_),
    .Q_N(_09617_),
    .Q(\spiking_network_top_uut.all_data_out[355] ));
 sg13g2_dfrbp_1 _20017_ (.CLK(net4804),
    .RESET_B(net4127),
    .D(_01333_),
    .Q_N(_09616_),
    .Q(\spiking_network_top_uut.all_data_out[356] ));
 sg13g2_dfrbp_1 _20018_ (.CLK(net4804),
    .RESET_B(net4126),
    .D(_01334_),
    .Q_N(_00278_),
    .Q(\spiking_network_top_uut.all_data_out[357] ));
 sg13g2_dfrbp_1 _20019_ (.CLK(net4804),
    .RESET_B(net4126),
    .D(_01335_),
    .Q_N(_00208_),
    .Q(\spiking_network_top_uut.all_data_out[358] ));
 sg13g2_dfrbp_1 _20020_ (.CLK(net4753),
    .RESET_B(net4074),
    .D(_01336_),
    .Q_N(_09615_),
    .Q(\spiking_network_top_uut.all_data_out[359] ));
 sg13g2_dfrbp_1 _20021_ (.CLK(net4745),
    .RESET_B(net4066),
    .D(_01337_),
    .Q_N(_09614_),
    .Q(\spiking_network_top_uut.all_data_out[720] ));
 sg13g2_dfrbp_1 _20022_ (.CLK(net4745),
    .RESET_B(net4066),
    .D(_01338_),
    .Q_N(_00372_),
    .Q(\spiking_network_top_uut.all_data_out[721] ));
 sg13g2_dfrbp_1 _20023_ (.CLK(net4746),
    .RESET_B(net4067),
    .D(_01339_),
    .Q_N(_00302_),
    .Q(\spiking_network_top_uut.all_data_out[722] ));
 sg13g2_dfrbp_1 _20024_ (.CLK(net4744),
    .RESET_B(net4065),
    .D(_01340_),
    .Q_N(_09613_),
    .Q(\spiking_network_top_uut.all_data_out[723] ));
 sg13g2_dfrbp_1 _20025_ (.CLK(net4767),
    .RESET_B(net4088),
    .D(_01341_),
    .Q_N(_09612_),
    .Q(\spiking_network_top_uut.all_data_out[724] ));
 sg13g2_dfrbp_1 _20026_ (.CLK(net4767),
    .RESET_B(net4088),
    .D(_01342_),
    .Q_N(_00232_),
    .Q(\spiking_network_top_uut.all_data_out[725] ));
 sg13g2_dfrbp_1 _20027_ (.CLK(net4767),
    .RESET_B(net4088),
    .D(_01343_),
    .Q_N(_00162_),
    .Q(\spiking_network_top_uut.all_data_out[726] ));
 sg13g2_dfrbp_1 _20028_ (.CLK(net4747),
    .RESET_B(net4069),
    .D(_01344_),
    .Q_N(_09611_),
    .Q(\spiking_network_top_uut.all_data_out[727] ));
 sg13g2_dfrbp_1 _20029_ (.CLK(net4809),
    .RESET_B(net4130),
    .D(_01345_),
    .Q_N(_09610_),
    .Q(\spiking_network_top_uut.all_data_out[344] ));
 sg13g2_dfrbp_1 _20030_ (.CLK(net4807),
    .RESET_B(net4133),
    .D(_01346_),
    .Q_N(_00419_),
    .Q(\spiking_network_top_uut.all_data_out[345] ));
 sg13g2_dfrbp_1 _20031_ (.CLK(net4812),
    .RESET_B(net4132),
    .D(_01347_),
    .Q_N(_00349_),
    .Q(\spiking_network_top_uut.all_data_out[346] ));
 sg13g2_dfrbp_1 _20032_ (.CLK(net4784),
    .RESET_B(net4106),
    .D(_01348_),
    .Q_N(_09609_),
    .Q(\spiking_network_top_uut.all_data_out[347] ));
 sg13g2_dfrbp_1 _20033_ (.CLK(net4798),
    .RESET_B(net4120),
    .D(_01349_),
    .Q_N(_09608_),
    .Q(\spiking_network_top_uut.all_data_out[348] ));
 sg13g2_dfrbp_1 _20034_ (.CLK(net4798),
    .RESET_B(net4120),
    .D(_01350_),
    .Q_N(_00279_),
    .Q(\spiking_network_top_uut.all_data_out[349] ));
 sg13g2_dfrbp_1 _20035_ (.CLK(net4798),
    .RESET_B(net4120),
    .D(_01351_),
    .Q_N(_00209_),
    .Q(\spiking_network_top_uut.all_data_out[350] ));
 sg13g2_dfrbp_1 _20036_ (.CLK(net4784),
    .RESET_B(net4106),
    .D(_01352_),
    .Q_N(_09607_),
    .Q(\spiking_network_top_uut.all_data_out[351] ));
 sg13g2_dfrbp_1 _20037_ (.CLK(net4744),
    .RESET_B(net4065),
    .D(_01353_),
    .Q_N(_09606_),
    .Q(\spiking_network_top_uut.all_data_out[592] ));
 sg13g2_dfrbp_1 _20038_ (.CLK(net4746),
    .RESET_B(net4065),
    .D(_01354_),
    .Q_N(_00388_),
    .Q(\spiking_network_top_uut.all_data_out[593] ));
 sg13g2_dfrbp_1 _20039_ (.CLK(net4744),
    .RESET_B(net4065),
    .D(_01355_),
    .Q_N(_00318_),
    .Q(\spiking_network_top_uut.all_data_out[594] ));
 sg13g2_dfrbp_1 _20040_ (.CLK(net4747),
    .RESET_B(net4068),
    .D(_01356_),
    .Q_N(_09605_),
    .Q(\spiking_network_top_uut.all_data_out[595] ));
 sg13g2_dfrbp_1 _20041_ (.CLK(net4765),
    .RESET_B(net4086),
    .D(_01357_),
    .Q_N(_09604_),
    .Q(\spiking_network_top_uut.all_data_out[596] ));
 sg13g2_dfrbp_1 _20042_ (.CLK(net4765),
    .RESET_B(net4086),
    .D(_01358_),
    .Q_N(_00248_),
    .Q(\spiking_network_top_uut.all_data_out[597] ));
 sg13g2_dfrbp_1 _20043_ (.CLK(net4765),
    .RESET_B(net4086),
    .D(_01359_),
    .Q_N(_00178_),
    .Q(\spiking_network_top_uut.all_data_out[598] ));
 sg13g2_dfrbp_1 _20044_ (.CLK(net4742),
    .RESET_B(net4063),
    .D(_01360_),
    .Q_N(_09603_),
    .Q(\spiking_network_top_uut.all_data_out[599] ));
 sg13g2_dfrbp_1 _20045_ (.CLK(net4781),
    .RESET_B(net4103),
    .D(_01361_),
    .Q_N(_09602_),
    .Q(\spiking_network_top_uut.all_data_out[336] ));
 sg13g2_dfrbp_1 _20046_ (.CLK(net4781),
    .RESET_B(net4103),
    .D(_01362_),
    .Q_N(_09601_),
    .Q(\spiking_network_top_uut.all_data_out[337] ));
 sg13g2_dfrbp_1 _20047_ (.CLK(net4781),
    .RESET_B(net4103),
    .D(_01363_),
    .Q_N(_09600_),
    .Q(\spiking_network_top_uut.all_data_out[338] ));
 sg13g2_dfrbp_1 _20048_ (.CLK(net4779),
    .RESET_B(net4102),
    .D(_01364_),
    .Q_N(_09599_),
    .Q(\spiking_network_top_uut.all_data_out[339] ));
 sg13g2_dfrbp_1 _20049_ (.CLK(net4752),
    .RESET_B(net4073),
    .D(_01365_),
    .Q_N(_09598_),
    .Q(\spiking_network_top_uut.all_data_out[340] ));
 sg13g2_dfrbp_1 _20050_ (.CLK(net4752),
    .RESET_B(net4073),
    .D(_01366_),
    .Q_N(_09597_),
    .Q(\spiking_network_top_uut.all_data_out[341] ));
 sg13g2_dfrbp_1 _20051_ (.CLK(net4754),
    .RESET_B(net4075),
    .D(_01367_),
    .Q_N(_09596_),
    .Q(\spiking_network_top_uut.all_data_out[342] ));
 sg13g2_dfrbp_1 _20052_ (.CLK(net4752),
    .RESET_B(net4073),
    .D(_01368_),
    .Q_N(_09595_),
    .Q(\spiking_network_top_uut.all_data_out[343] ));
 sg13g2_dfrbp_1 _20053_ (.CLK(net4710),
    .RESET_B(net4030),
    .D(_01369_),
    .Q_N(_09594_),
    .Q(\spiking_network_top_uut.all_data_out[728] ));
 sg13g2_dfrbp_1 _20054_ (.CLK(net4710),
    .RESET_B(net4030),
    .D(_01370_),
    .Q_N(_00371_),
    .Q(\spiking_network_top_uut.all_data_out[729] ));
 sg13g2_dfrbp_1 _20055_ (.CLK(net4710),
    .RESET_B(net4030),
    .D(_01371_),
    .Q_N(_00301_),
    .Q(\spiking_network_top_uut.all_data_out[730] ));
 sg13g2_dfrbp_1 _20056_ (.CLK(net4716),
    .RESET_B(net4036),
    .D(_01372_),
    .Q_N(_09593_),
    .Q(\spiking_network_top_uut.all_data_out[731] ));
 sg13g2_dfrbp_1 _20057_ (.CLK(net4717),
    .RESET_B(net4037),
    .D(_01373_),
    .Q_N(_09592_),
    .Q(\spiking_network_top_uut.all_data_out[732] ));
 sg13g2_dfrbp_1 _20058_ (.CLK(net4741),
    .RESET_B(net4060),
    .D(_01374_),
    .Q_N(_00231_),
    .Q(\spiking_network_top_uut.all_data_out[733] ));
 sg13g2_dfrbp_1 _20059_ (.CLK(net4717),
    .RESET_B(net4037),
    .D(_01375_),
    .Q_N(_00161_),
    .Q(\spiking_network_top_uut.all_data_out[734] ));
 sg13g2_dfrbp_1 _20060_ (.CLK(net4713),
    .RESET_B(net4033),
    .D(_01376_),
    .Q_N(_09591_),
    .Q(\spiking_network_top_uut.all_data_out[735] ));
 sg13g2_dfrbp_1 _20061_ (.CLK(net4789),
    .RESET_B(net4111),
    .D(_01377_),
    .Q_N(_09590_),
    .Q(\spiking_network_top_uut.all_data_out[328] ));
 sg13g2_dfrbp_1 _20062_ (.CLK(net4795),
    .RESET_B(net4117),
    .D(_01378_),
    .Q_N(_09589_),
    .Q(\spiking_network_top_uut.all_data_out[329] ));
 sg13g2_dfrbp_1 _20063_ (.CLK(net4791),
    .RESET_B(net4113),
    .D(_01379_),
    .Q_N(_09588_),
    .Q(\spiking_network_top_uut.all_data_out[330] ));
 sg13g2_dfrbp_1 _20064_ (.CLK(net4773),
    .RESET_B(net4094),
    .D(_01380_),
    .Q_N(_09587_),
    .Q(\spiking_network_top_uut.all_data_out[331] ));
 sg13g2_dfrbp_1 _20065_ (.CLK(net4796),
    .RESET_B(net4123),
    .D(_01381_),
    .Q_N(_09586_),
    .Q(\spiking_network_top_uut.all_data_out[332] ));
 sg13g2_dfrbp_1 _20066_ (.CLK(net4796),
    .RESET_B(net4117),
    .D(_01382_),
    .Q_N(_09585_),
    .Q(\spiking_network_top_uut.all_data_out[333] ));
 sg13g2_dfrbp_1 _20067_ (.CLK(net4795),
    .RESET_B(net4117),
    .D(_01383_),
    .Q_N(_09584_),
    .Q(\spiking_network_top_uut.all_data_out[334] ));
 sg13g2_dfrbp_1 _20068_ (.CLK(net4790),
    .RESET_B(net4112),
    .D(_01384_),
    .Q_N(_09583_),
    .Q(\spiking_network_top_uut.all_data_out[335] ));
 sg13g2_dfrbp_1 _20069_ (.CLK(net4762),
    .RESET_B(net4083),
    .D(_01385_),
    .Q_N(_09582_),
    .Q(\spiking_network_top_uut.all_data_out[528] ));
 sg13g2_dfrbp_1 _20070_ (.CLK(net4780),
    .RESET_B(net4101),
    .D(_01386_),
    .Q_N(_00396_),
    .Q(\spiking_network_top_uut.all_data_out[529] ));
 sg13g2_dfrbp_1 _20071_ (.CLK(net4758),
    .RESET_B(net4079),
    .D(_01387_),
    .Q_N(_00326_),
    .Q(\spiking_network_top_uut.all_data_out[530] ));
 sg13g2_dfrbp_1 _20072_ (.CLK(net4736),
    .RESET_B(net4057),
    .D(_01388_),
    .Q_N(_09581_),
    .Q(\spiking_network_top_uut.all_data_out[531] ));
 sg13g2_dfrbp_1 _20073_ (.CLK(net4753),
    .RESET_B(net4074),
    .D(_01389_),
    .Q_N(_09580_),
    .Q(\spiking_network_top_uut.all_data_out[532] ));
 sg13g2_dfrbp_1 _20074_ (.CLK(net4760),
    .RESET_B(net4081),
    .D(_01390_),
    .Q_N(_00256_),
    .Q(\spiking_network_top_uut.all_data_out[533] ));
 sg13g2_dfrbp_1 _20075_ (.CLK(net4760),
    .RESET_B(net4081),
    .D(_01391_),
    .Q_N(_00186_),
    .Q(\spiking_network_top_uut.all_data_out[534] ));
 sg13g2_dfrbp_1 _20076_ (.CLK(net4752),
    .RESET_B(net4073),
    .D(_01392_),
    .Q_N(_09579_),
    .Q(\spiking_network_top_uut.all_data_out[535] ));
 sg13g2_dfrbp_1 _20077_ (.CLK(net4805),
    .RESET_B(net4127),
    .D(_01393_),
    .Q_N(_09578_),
    .Q(\spiking_network_top_uut.all_data_out[320] ));
 sg13g2_dfrbp_1 _20078_ (.CLK(net4805),
    .RESET_B(net4127),
    .D(_01394_),
    .Q_N(_00420_),
    .Q(\spiking_network_top_uut.all_data_out[321] ));
 sg13g2_dfrbp_1 _20079_ (.CLK(net4803),
    .RESET_B(net4125),
    .D(_01395_),
    .Q_N(_00350_),
    .Q(\spiking_network_top_uut.all_data_out[322] ));
 sg13g2_dfrbp_1 _20080_ (.CLK(net4784),
    .RESET_B(net4106),
    .D(_01396_),
    .Q_N(_09577_),
    .Q(\spiking_network_top_uut.all_data_out[323] ));
 sg13g2_dfrbp_1 _20081_ (.CLK(net4802),
    .RESET_B(net4124),
    .D(_01397_),
    .Q_N(_09576_),
    .Q(\spiking_network_top_uut.all_data_out[324] ));
 sg13g2_dfrbp_1 _20082_ (.CLK(net4802),
    .RESET_B(net4124),
    .D(_01398_),
    .Q_N(_00280_),
    .Q(\spiking_network_top_uut.all_data_out[325] ));
 sg13g2_dfrbp_1 _20083_ (.CLK(net4802),
    .RESET_B(net4124),
    .D(_01399_),
    .Q_N(_00210_),
    .Q(\spiking_network_top_uut.all_data_out[326] ));
 sg13g2_dfrbp_1 _20084_ (.CLK(net4802),
    .RESET_B(net4124),
    .D(_01400_),
    .Q_N(_09575_),
    .Q(\spiking_network_top_uut.all_data_out[327] ));
 sg13g2_dfrbp_1 _20085_ (.CLK(net4686),
    .RESET_B(net4005),
    .D(_01401_),
    .Q_N(_09574_),
    .Q(\spiking_network_top_uut.all_data_out[736] ));
 sg13g2_dfrbp_1 _20086_ (.CLK(net4690),
    .RESET_B(net4005),
    .D(_01402_),
    .Q_N(_00370_),
    .Q(\spiking_network_top_uut.all_data_out[737] ));
 sg13g2_dfrbp_1 _20087_ (.CLK(net4687),
    .RESET_B(net4006),
    .D(_01403_),
    .Q_N(_00300_),
    .Q(\spiking_network_top_uut.all_data_out[738] ));
 sg13g2_dfrbp_1 _20088_ (.CLK(net4668),
    .RESET_B(net3988),
    .D(_01404_),
    .Q_N(_09573_),
    .Q(\spiking_network_top_uut.all_data_out[739] ));
 sg13g2_dfrbp_1 _20089_ (.CLK(net4675),
    .RESET_B(net3993),
    .D(_01405_),
    .Q_N(_09572_),
    .Q(\spiking_network_top_uut.all_data_out[740] ));
 sg13g2_dfrbp_1 _20090_ (.CLK(net4675),
    .RESET_B(net3994),
    .D(_01406_),
    .Q_N(_00230_),
    .Q(\spiking_network_top_uut.all_data_out[741] ));
 sg13g2_dfrbp_1 _20091_ (.CLK(net4673),
    .RESET_B(net3992),
    .D(_01407_),
    .Q_N(_00160_),
    .Q(\spiking_network_top_uut.all_data_out[742] ));
 sg13g2_dfrbp_1 _20092_ (.CLK(net4674),
    .RESET_B(net3994),
    .D(_01408_),
    .Q_N(_09571_),
    .Q(\spiking_network_top_uut.all_data_out[743] ));
 sg13g2_dfrbp_1 _20093_ (.CLK(net4656),
    .RESET_B(net3975),
    .D(_01409_),
    .Q_N(_09570_),
    .Q(\spiking_network_top_uut.all_data_out[312] ));
 sg13g2_dfrbp_1 _20094_ (.CLK(net4657),
    .RESET_B(net3976),
    .D(_01410_),
    .Q_N(_09569_),
    .Q(\spiking_network_top_uut.all_data_out[313] ));
 sg13g2_dfrbp_1 _20095_ (.CLK(net4657),
    .RESET_B(net3976),
    .D(_01411_),
    .Q_N(_09568_),
    .Q(\spiking_network_top_uut.all_data_out[314] ));
 sg13g2_dfrbp_1 _20096_ (.CLK(net4657),
    .RESET_B(net3976),
    .D(_01412_),
    .Q_N(_09567_),
    .Q(\spiking_network_top_uut.all_data_out[315] ));
 sg13g2_dfrbp_1 _20097_ (.CLK(net4662),
    .RESET_B(net3982),
    .D(_01413_),
    .Q_N(_09566_),
    .Q(\spiking_network_top_uut.all_data_out[316] ));
 sg13g2_dfrbp_1 _20098_ (.CLK(net4661),
    .RESET_B(net3981),
    .D(_01414_),
    .Q_N(_09565_),
    .Q(\spiking_network_top_uut.all_data_out[317] ));
 sg13g2_dfrbp_1 _20099_ (.CLK(net4661),
    .RESET_B(net3981),
    .D(_01415_),
    .Q_N(_09564_),
    .Q(\spiking_network_top_uut.all_data_out[318] ));
 sg13g2_dfrbp_1 _20100_ (.CLK(net4658),
    .RESET_B(net3977),
    .D(_01416_),
    .Q_N(_09563_),
    .Q(\spiking_network_top_uut.all_data_out[319] ));
 sg13g2_dfrbp_1 _20101_ (.CLK(net4685),
    .RESET_B(net4004),
    .D(_01417_),
    .Q_N(_09562_),
    .Q(\spiking_network_top_uut.all_data_out[632] ));
 sg13g2_dfrbp_1 _20102_ (.CLK(net4685),
    .RESET_B(net4004),
    .D(_01418_),
    .Q_N(_00383_),
    .Q(\spiking_network_top_uut.all_data_out[633] ));
 sg13g2_dfrbp_1 _20103_ (.CLK(net4685),
    .RESET_B(net4004),
    .D(_01419_),
    .Q_N(_00313_),
    .Q(\spiking_network_top_uut.all_data_out[634] ));
 sg13g2_dfrbp_1 _20104_ (.CLK(net4724),
    .RESET_B(net4044),
    .D(_01420_),
    .Q_N(_09561_),
    .Q(\spiking_network_top_uut.all_data_out[635] ));
 sg13g2_dfrbp_1 _20105_ (.CLK(net4739),
    .RESET_B(net4060),
    .D(_01421_),
    .Q_N(_09560_),
    .Q(\spiking_network_top_uut.all_data_out[636] ));
 sg13g2_dfrbp_1 _20106_ (.CLK(net4739),
    .RESET_B(net4060),
    .D(_01422_),
    .Q_N(_00243_),
    .Q(\spiking_network_top_uut.all_data_out[637] ));
 sg13g2_dfrbp_1 _20107_ (.CLK(net4739),
    .RESET_B(net4060),
    .D(_01423_),
    .Q_N(_00173_),
    .Q(\spiking_network_top_uut.all_data_out[638] ));
 sg13g2_dfrbp_1 _20108_ (.CLK(net4700),
    .RESET_B(net4020),
    .D(_01424_),
    .Q_N(_09559_),
    .Q(\spiking_network_top_uut.all_data_out[639] ));
 sg13g2_dfrbp_1 _20109_ (.CLK(net4651),
    .RESET_B(net3970),
    .D(_01425_),
    .Q_N(_09558_),
    .Q(\spiking_network_top_uut.all_data_out[304] ));
 sg13g2_dfrbp_1 _20110_ (.CLK(net4651),
    .RESET_B(net3970),
    .D(_01426_),
    .Q_N(_09557_),
    .Q(\spiking_network_top_uut.all_data_out[305] ));
 sg13g2_dfrbp_1 _20111_ (.CLK(net4651),
    .RESET_B(net3970),
    .D(_01427_),
    .Q_N(_09556_),
    .Q(\spiking_network_top_uut.all_data_out[306] ));
 sg13g2_dfrbp_1 _20112_ (.CLK(net4651),
    .RESET_B(net3970),
    .D(_01428_),
    .Q_N(_09555_),
    .Q(\spiking_network_top_uut.all_data_out[307] ));
 sg13g2_dfrbp_1 _20113_ (.CLK(net4662),
    .RESET_B(net3982),
    .D(_01429_),
    .Q_N(_09554_),
    .Q(\spiking_network_top_uut.all_data_out[308] ));
 sg13g2_dfrbp_1 _20114_ (.CLK(net4658),
    .RESET_B(net3977),
    .D(_01430_),
    .Q_N(_09553_),
    .Q(\spiking_network_top_uut.all_data_out[309] ));
 sg13g2_dfrbp_1 _20115_ (.CLK(net4656),
    .RESET_B(net3975),
    .D(_01431_),
    .Q_N(_09552_),
    .Q(\spiking_network_top_uut.all_data_out[310] ));
 sg13g2_dfrbp_1 _20116_ (.CLK(net4656),
    .RESET_B(net3975),
    .D(_01432_),
    .Q_N(_09551_),
    .Q(\spiking_network_top_uut.all_data_out[311] ));
 sg13g2_dfrbp_1 _20117_ (.CLK(net4783),
    .RESET_B(net4105),
    .D(_01433_),
    .Q_N(_09550_),
    .Q(\spiking_network_top_uut.all_data_out[744] ));
 sg13g2_dfrbp_1 _20118_ (.CLK(net4793),
    .RESET_B(net4115),
    .D(_01434_),
    .Q_N(_00369_),
    .Q(\spiking_network_top_uut.all_data_out[745] ));
 sg13g2_dfrbp_1 _20119_ (.CLK(net4793),
    .RESET_B(net4115),
    .D(_01435_),
    .Q_N(_00299_),
    .Q(\spiking_network_top_uut.all_data_out[746] ));
 sg13g2_dfrbp_1 _20120_ (.CLK(net4757),
    .RESET_B(net4078),
    .D(_01436_),
    .Q_N(_09549_),
    .Q(\spiking_network_top_uut.all_data_out[747] ));
 sg13g2_dfrbp_1 _20121_ (.CLK(net4784),
    .RESET_B(net4106),
    .D(_01437_),
    .Q_N(_09548_),
    .Q(\spiking_network_top_uut.all_data_out[748] ));
 sg13g2_dfrbp_1 _20122_ (.CLK(net4778),
    .RESET_B(net4099),
    .D(_01438_),
    .Q_N(_00229_),
    .Q(\spiking_network_top_uut.all_data_out[749] ));
 sg13g2_dfrbp_1 _20123_ (.CLK(net4779),
    .RESET_B(net4100),
    .D(_01439_),
    .Q_N(_00159_),
    .Q(\spiking_network_top_uut.all_data_out[750] ));
 sg13g2_dfrbp_1 _20124_ (.CLK(net4755),
    .RESET_B(net4076),
    .D(_01440_),
    .Q_N(_09547_),
    .Q(\spiking_network_top_uut.all_data_out[751] ));
 sg13g2_dfrbp_1 _20125_ (.CLK(net4652),
    .RESET_B(net3971),
    .D(_01441_),
    .Q_N(_09546_),
    .Q(\spiking_network_top_uut.all_data_out[296] ));
 sg13g2_dfrbp_1 _20126_ (.CLK(net4652),
    .RESET_B(net3971),
    .D(_01442_),
    .Q_N(_09545_),
    .Q(\spiking_network_top_uut.all_data_out[297] ));
 sg13g2_dfrbp_1 _20127_ (.CLK(net4652),
    .RESET_B(net3971),
    .D(_01443_),
    .Q_N(_09544_),
    .Q(\spiking_network_top_uut.all_data_out[298] ));
 sg13g2_dfrbp_1 _20128_ (.CLK(net4652),
    .RESET_B(net3971),
    .D(_01444_),
    .Q_N(_09543_),
    .Q(\spiking_network_top_uut.all_data_out[299] ));
 sg13g2_dfrbp_1 _20129_ (.CLK(net4661),
    .RESET_B(net3981),
    .D(_01445_),
    .Q_N(_09542_),
    .Q(\spiking_network_top_uut.all_data_out[300] ));
 sg13g2_dfrbp_1 _20130_ (.CLK(net4661),
    .RESET_B(net3981),
    .D(_01446_),
    .Q_N(_09541_),
    .Q(\spiking_network_top_uut.all_data_out[301] ));
 sg13g2_dfrbp_1 _20131_ (.CLK(net4661),
    .RESET_B(net3981),
    .D(_01447_),
    .Q_N(_09540_),
    .Q(\spiking_network_top_uut.all_data_out[302] ));
 sg13g2_dfrbp_1 _20132_ (.CLK(net4656),
    .RESET_B(net3975),
    .D(_01448_),
    .Q_N(_09539_),
    .Q(\spiking_network_top_uut.all_data_out[303] ));
 sg13g2_dfrbp_1 _20133_ (.CLK(net4797),
    .RESET_B(net4118),
    .D(_01449_),
    .Q_N(_09538_),
    .Q(\spiking_network_top_uut.all_data_out[520] ));
 sg13g2_dfrbp_1 _20134_ (.CLK(net4791),
    .RESET_B(net4113),
    .D(_01450_),
    .Q_N(_00397_),
    .Q(\spiking_network_top_uut.all_data_out[521] ));
 sg13g2_dfrbp_1 _20135_ (.CLK(net4797),
    .RESET_B(net4118),
    .D(_01451_),
    .Q_N(_00327_),
    .Q(\spiking_network_top_uut.all_data_out[522] ));
 sg13g2_dfrbp_1 _20136_ (.CLK(net4773),
    .RESET_B(net4094),
    .D(_01452_),
    .Q_N(_09537_),
    .Q(\spiking_network_top_uut.all_data_out[523] ));
 sg13g2_dfrbp_1 _20137_ (.CLK(net4800),
    .RESET_B(net4120),
    .D(_01453_),
    .Q_N(_09536_),
    .Q(\spiking_network_top_uut.all_data_out[524] ));
 sg13g2_dfrbp_1 _20138_ (.CLK(net4799),
    .RESET_B(net4119),
    .D(_01454_),
    .Q_N(_00257_),
    .Q(\spiking_network_top_uut.all_data_out[525] ));
 sg13g2_dfrbp_1 _20139_ (.CLK(net4799),
    .RESET_B(net4121),
    .D(_01455_),
    .Q_N(_00187_),
    .Q(\spiking_network_top_uut.all_data_out[526] ));
 sg13g2_dfrbp_1 _20140_ (.CLK(net4774),
    .RESET_B(net4095),
    .D(_01456_),
    .Q_N(_09535_),
    .Q(\spiking_network_top_uut.all_data_out[527] ));
 sg13g2_dfrbp_1 _20141_ (.CLK(net4650),
    .RESET_B(net3969),
    .D(_01457_),
    .Q_N(_09534_),
    .Q(\spiking_network_top_uut.all_data_out[288] ));
 sg13g2_dfrbp_1 _20142_ (.CLK(net4649),
    .RESET_B(net3968),
    .D(_01458_),
    .Q_N(_09533_),
    .Q(\spiking_network_top_uut.all_data_out[289] ));
 sg13g2_dfrbp_1 _20143_ (.CLK(net4650),
    .RESET_B(net3969),
    .D(_01459_),
    .Q_N(_09532_),
    .Q(\spiking_network_top_uut.all_data_out[290] ));
 sg13g2_dfrbp_1 _20144_ (.CLK(net4650),
    .RESET_B(net3969),
    .D(_01460_),
    .Q_N(_09531_),
    .Q(\spiking_network_top_uut.all_data_out[291] ));
 sg13g2_dfrbp_1 _20145_ (.CLK(net4656),
    .RESET_B(net3975),
    .D(_01461_),
    .Q_N(_09530_),
    .Q(\spiking_network_top_uut.all_data_out[292] ));
 sg13g2_dfrbp_1 _20146_ (.CLK(net4652),
    .RESET_B(net3971),
    .D(_01462_),
    .Q_N(_09529_),
    .Q(\spiking_network_top_uut.all_data_out[293] ));
 sg13g2_dfrbp_1 _20147_ (.CLK(net4657),
    .RESET_B(net3976),
    .D(_01463_),
    .Q_N(_09528_),
    .Q(\spiking_network_top_uut.all_data_out[294] ));
 sg13g2_dfrbp_1 _20148_ (.CLK(net4657),
    .RESET_B(net3976),
    .D(_01464_),
    .Q_N(_09527_),
    .Q(\spiking_network_top_uut.all_data_out[295] ));
 sg13g2_dfrbp_1 _20149_ (.CLK(net4745),
    .RESET_B(net4066),
    .D(_01465_),
    .Q_N(_09526_),
    .Q(\spiking_network_top_uut.all_data_out[752] ));
 sg13g2_dfrbp_1 _20150_ (.CLK(net4746),
    .RESET_B(net4067),
    .D(_01466_),
    .Q_N(_00368_),
    .Q(\spiking_network_top_uut.all_data_out[753] ));
 sg13g2_dfrbp_1 _20151_ (.CLK(net4745),
    .RESET_B(net4066),
    .D(_01467_),
    .Q_N(_00298_),
    .Q(\spiking_network_top_uut.all_data_out[754] ));
 sg13g2_dfrbp_1 _20152_ (.CLK(net4748),
    .RESET_B(net4069),
    .D(_01468_),
    .Q_N(_09525_),
    .Q(\spiking_network_top_uut.all_data_out[755] ));
 sg13g2_dfrbp_1 _20153_ (.CLK(net4767),
    .RESET_B(net4088),
    .D(_01469_),
    .Q_N(_09524_),
    .Q(\spiking_network_top_uut.all_data_out[756] ));
 sg13g2_dfrbp_1 _20154_ (.CLK(net4768),
    .RESET_B(net4088),
    .D(_01470_),
    .Q_N(_00228_),
    .Q(\spiking_network_top_uut.all_data_out[757] ));
 sg13g2_dfrbp_1 _20155_ (.CLK(net4767),
    .RESET_B(net4089),
    .D(_01471_),
    .Q_N(_00158_),
    .Q(\spiking_network_top_uut.all_data_out[758] ));
 sg13g2_dfrbp_1 _20156_ (.CLK(net4748),
    .RESET_B(net4069),
    .D(_01472_),
    .Q_N(_09523_),
    .Q(\spiking_network_top_uut.all_data_out[759] ));
 sg13g2_dfrbp_1 _20157_ (.CLK(net4720),
    .RESET_B(net4041),
    .D(_01473_),
    .Q_N(_09522_),
    .Q(\spiking_network_top_uut.all_data_out[280] ));
 sg13g2_dfrbp_1 _20158_ (.CLK(net4713),
    .RESET_B(net4033),
    .D(_01474_),
    .Q_N(_09521_),
    .Q(\spiking_network_top_uut.all_data_out[281] ));
 sg13g2_dfrbp_1 _20159_ (.CLK(net4720),
    .RESET_B(net4052),
    .D(_01475_),
    .Q_N(_09520_),
    .Q(\spiking_network_top_uut.all_data_out[282] ));
 sg13g2_dfrbp_1 _20160_ (.CLK(net4720),
    .RESET_B(net4041),
    .D(_01476_),
    .Q_N(_09519_),
    .Q(\spiking_network_top_uut.all_data_out[283] ));
 sg13g2_dfrbp_1 _20161_ (.CLK(net4719),
    .RESET_B(net4040),
    .D(_01477_),
    .Q_N(_09518_),
    .Q(\spiking_network_top_uut.all_data_out[284] ));
 sg13g2_dfrbp_1 _20162_ (.CLK(net4720),
    .RESET_B(net4041),
    .D(_01478_),
    .Q_N(_09517_),
    .Q(\spiking_network_top_uut.all_data_out[285] ));
 sg13g2_dfrbp_1 _20163_ (.CLK(net4713),
    .RESET_B(net4033),
    .D(_01479_),
    .Q_N(_09516_),
    .Q(\spiking_network_top_uut.all_data_out[286] ));
 sg13g2_dfrbp_1 _20164_ (.CLK(net4719),
    .RESET_B(net4040),
    .D(_01480_),
    .Q_N(_09515_),
    .Q(\spiking_network_top_uut.all_data_out[287] ));
 sg13g2_dfrbp_1 _20165_ (.CLK(net4686),
    .RESET_B(net4005),
    .D(_01481_),
    .Q_N(_09514_),
    .Q(\spiking_network_top_uut.all_data_out[576] ));
 sg13g2_dfrbp_1 _20166_ (.CLK(net4686),
    .RESET_B(net4005),
    .D(_01482_),
    .Q_N(_00390_),
    .Q(\spiking_network_top_uut.all_data_out[577] ));
 sg13g2_dfrbp_1 _20167_ (.CLK(net4686),
    .RESET_B(net4005),
    .D(_01483_),
    .Q_N(_00320_),
    .Q(\spiking_network_top_uut.all_data_out[578] ));
 sg13g2_dfrbp_1 _20168_ (.CLK(net4689),
    .RESET_B(net4018),
    .D(_01484_),
    .Q_N(_09513_),
    .Q(\spiking_network_top_uut.all_data_out[579] ));
 sg13g2_dfrbp_1 _20169_ (.CLK(net4692),
    .RESET_B(net4011),
    .D(_01485_),
    .Q_N(_09512_),
    .Q(\spiking_network_top_uut.all_data_out[580] ));
 sg13g2_dfrbp_1 _20170_ (.CLK(net4698),
    .RESET_B(net4018),
    .D(_01486_),
    .Q_N(_00250_),
    .Q(\spiking_network_top_uut.all_data_out[581] ));
 sg13g2_dfrbp_1 _20171_ (.CLK(net4692),
    .RESET_B(net4011),
    .D(_01487_),
    .Q_N(_00180_),
    .Q(\spiking_network_top_uut.all_data_out[582] ));
 sg13g2_dfrbp_1 _20172_ (.CLK(net4698),
    .RESET_B(net4018),
    .D(_01488_),
    .Q_N(_09511_),
    .Q(\spiking_network_top_uut.all_data_out[583] ));
 sg13g2_dfrbp_1 _20173_ (.CLK(net4662),
    .RESET_B(net3982),
    .D(_01489_),
    .Q_N(_09510_),
    .Q(\spiking_network_top_uut.all_data_out[272] ));
 sg13g2_dfrbp_1 _20174_ (.CLK(net4671),
    .RESET_B(net3990),
    .D(_01490_),
    .Q_N(_09509_),
    .Q(\spiking_network_top_uut.all_data_out[273] ));
 sg13g2_dfrbp_1 _20175_ (.CLK(net4671),
    .RESET_B(net3990),
    .D(_01491_),
    .Q_N(_09508_),
    .Q(\spiking_network_top_uut.all_data_out[274] ));
 sg13g2_dfrbp_1 _20176_ (.CLK(net4671),
    .RESET_B(net3990),
    .D(_01492_),
    .Q_N(_09507_),
    .Q(\spiking_network_top_uut.all_data_out[275] ));
 sg13g2_dfrbp_1 _20177_ (.CLK(net4725),
    .RESET_B(net4045),
    .D(_01493_),
    .Q_N(_09506_),
    .Q(\spiking_network_top_uut.all_data_out[276] ));
 sg13g2_dfrbp_1 _20178_ (.CLK(net4719),
    .RESET_B(net4053),
    .D(_01494_),
    .Q_N(_09505_),
    .Q(\spiking_network_top_uut.all_data_out[277] ));
 sg13g2_dfrbp_1 _20179_ (.CLK(net4721),
    .RESET_B(net4053),
    .D(_01495_),
    .Q_N(_09504_),
    .Q(\spiking_network_top_uut.all_data_out[278] ));
 sg13g2_dfrbp_1 _20180_ (.CLK(net4714),
    .RESET_B(net4034),
    .D(_01496_),
    .Q_N(_09503_),
    .Q(\spiking_network_top_uut.all_data_out[279] ));
 sg13g2_dfrbp_1 _20181_ (.CLK(net4685),
    .RESET_B(net4004),
    .D(_01497_),
    .Q_N(_09502_),
    .Q(\spiking_network_top_uut.all_data_out[760] ));
 sg13g2_dfrbp_1 _20182_ (.CLK(net4710),
    .RESET_B(net4030),
    .D(_01498_),
    .Q_N(_00367_),
    .Q(\spiking_network_top_uut.all_data_out[761] ));
 sg13g2_dfrbp_1 _20183_ (.CLK(net4715),
    .RESET_B(net4035),
    .D(_01499_),
    .Q_N(_00297_),
    .Q(\spiking_network_top_uut.all_data_out[762] ));
 sg13g2_dfrbp_1 _20184_ (.CLK(net4700),
    .RESET_B(net4020),
    .D(_01500_),
    .Q_N(_09501_),
    .Q(\spiking_network_top_uut.all_data_out[763] ));
 sg13g2_dfrbp_1 _20185_ (.CLK(net4716),
    .RESET_B(net4036),
    .D(_01501_),
    .Q_N(_09500_),
    .Q(\spiking_network_top_uut.all_data_out[764] ));
 sg13g2_dfrbp_1 _20186_ (.CLK(net4716),
    .RESET_B(net4036),
    .D(_01502_),
    .Q_N(_00227_),
    .Q(\spiking_network_top_uut.all_data_out[765] ));
 sg13g2_dfrbp_1 _20187_ (.CLK(net4717),
    .RESET_B(net4038),
    .D(_01503_),
    .Q_N(_00157_),
    .Q(\spiking_network_top_uut.all_data_out[766] ));
 sg13g2_dfrbp_1 _20188_ (.CLK(net4724),
    .RESET_B(net4044),
    .D(_01504_),
    .Q_N(_09499_),
    .Q(\spiking_network_top_uut.all_data_out[767] ));
 sg13g2_dfrbp_1 _20189_ (.CLK(net4717),
    .RESET_B(net4038),
    .D(_01505_),
    .Q_N(_09498_),
    .Q(\spiking_network_top_uut.all_data_out[264] ));
 sg13g2_dfrbp_1 _20190_ (.CLK(net4717),
    .RESET_B(net4038),
    .D(_01506_),
    .Q_N(_09497_),
    .Q(\spiking_network_top_uut.all_data_out[265] ));
 sg13g2_dfrbp_1 _20191_ (.CLK(net4710),
    .RESET_B(net4030),
    .D(_01507_),
    .Q_N(_09496_),
    .Q(\spiking_network_top_uut.all_data_out[266] ));
 sg13g2_dfrbp_1 _20192_ (.CLK(net4711),
    .RESET_B(net4031),
    .D(_01508_),
    .Q_N(_09495_),
    .Q(\spiking_network_top_uut.all_data_out[267] ));
 sg13g2_dfrbp_1 _20193_ (.CLK(net4710),
    .RESET_B(net4030),
    .D(_01509_),
    .Q_N(_09494_),
    .Q(\spiking_network_top_uut.all_data_out[268] ));
 sg13g2_dfrbp_1 _20194_ (.CLK(net4719),
    .RESET_B(net4040),
    .D(_01510_),
    .Q_N(_09493_),
    .Q(\spiking_network_top_uut.all_data_out[269] ));
 sg13g2_dfrbp_1 _20195_ (.CLK(net4722),
    .RESET_B(net4031),
    .D(_01511_),
    .Q_N(_09492_),
    .Q(\spiking_network_top_uut.all_data_out[270] ));
 sg13g2_dfrbp_1 _20196_ (.CLK(net4711),
    .RESET_B(net4033),
    .D(_01512_),
    .Q_N(_09491_),
    .Q(\spiking_network_top_uut.all_data_out[271] ));
 sg13g2_dfrbp_1 _20197_ (.CLK(net4803),
    .RESET_B(net4125),
    .D(_01513_),
    .Q_N(_09490_),
    .Q(\spiking_network_top_uut.all_data_out[512] ));
 sg13g2_dfrbp_1 _20198_ (.CLK(net4787),
    .RESET_B(net4109),
    .D(_01514_),
    .Q_N(_00398_),
    .Q(\spiking_network_top_uut.all_data_out[513] ));
 sg13g2_dfrbp_1 _20199_ (.CLK(net4787),
    .RESET_B(net4109),
    .D(_01515_),
    .Q_N(_00328_),
    .Q(\spiking_network_top_uut.all_data_out[514] ));
 sg13g2_dfrbp_1 _20200_ (.CLK(net4751),
    .RESET_B(net4072),
    .D(_01516_),
    .Q_N(_09489_),
    .Q(\spiking_network_top_uut.all_data_out[515] ));
 sg13g2_dfrbp_1 _20201_ (.CLK(net4791),
    .RESET_B(net4113),
    .D(_01517_),
    .Q_N(_09488_),
    .Q(\spiking_network_top_uut.all_data_out[516] ));
 sg13g2_dfrbp_1 _20202_ (.CLK(net4792),
    .RESET_B(net4114),
    .D(_01518_),
    .Q_N(_00258_),
    .Q(\spiking_network_top_uut.all_data_out[517] ));
 sg13g2_dfrbp_1 _20203_ (.CLK(net4792),
    .RESET_B(net4114),
    .D(_01519_),
    .Q_N(_00188_),
    .Q(\spiking_network_top_uut.all_data_out[518] ));
 sg13g2_dfrbp_1 _20204_ (.CLK(net4757),
    .RESET_B(net4078),
    .D(_01520_),
    .Q_N(_09487_),
    .Q(\spiking_network_top_uut.all_data_out[519] ));
 sg13g2_dfrbp_1 _20205_ (.CLK(net4667),
    .RESET_B(net3986),
    .D(_01521_),
    .Q_N(_09486_),
    .Q(\spiking_network_top_uut.all_data_out[256] ));
 sg13g2_dfrbp_1 _20206_ (.CLK(net4666),
    .RESET_B(net3986),
    .D(_01522_),
    .Q_N(_09485_),
    .Q(\spiking_network_top_uut.all_data_out[257] ));
 sg13g2_dfrbp_1 _20207_ (.CLK(net4662),
    .RESET_B(net3982),
    .D(_01523_),
    .Q_N(_09484_),
    .Q(\spiking_network_top_uut.all_data_out[258] ));
 sg13g2_dfrbp_1 _20208_ (.CLK(net4662),
    .RESET_B(net3982),
    .D(_01524_),
    .Q_N(_09483_),
    .Q(\spiking_network_top_uut.all_data_out[259] ));
 sg13g2_dfrbp_1 _20209_ (.CLK(net4720),
    .RESET_B(net4041),
    .D(_01525_),
    .Q_N(_09482_),
    .Q(\spiking_network_top_uut.all_data_out[260] ));
 sg13g2_dfrbp_1 _20210_ (.CLK(net4713),
    .RESET_B(net4033),
    .D(_01526_),
    .Q_N(_09481_),
    .Q(\spiking_network_top_uut.all_data_out[261] ));
 sg13g2_dfrbp_1 _20211_ (.CLK(net4720),
    .RESET_B(net4041),
    .D(_01527_),
    .Q_N(_09480_),
    .Q(\spiking_network_top_uut.all_data_out[262] ));
 sg13g2_dfrbp_1 _20212_ (.CLK(net4713),
    .RESET_B(net4033),
    .D(_01528_),
    .Q_N(_09479_),
    .Q(\spiking_network_top_uut.all_data_out[263] ));
 sg13g2_dfrbp_1 _20213_ (.CLK(net4681),
    .RESET_B(net4000),
    .D(_01529_),
    .Q_N(_09478_),
    .Q(\spiking_network_top_uut.all_data_out[768] ));
 sg13g2_dfrbp_1 _20214_ (.CLK(net4684),
    .RESET_B(net4002),
    .D(_01530_),
    .Q_N(_00366_),
    .Q(\spiking_network_top_uut.all_data_out[769] ));
 sg13g2_dfrbp_1 _20215_ (.CLK(net4687),
    .RESET_B(net4006),
    .D(_01531_),
    .Q_N(_00296_),
    .Q(\spiking_network_top_uut.all_data_out[770] ));
 sg13g2_dfrbp_1 _20216_ (.CLK(net4662),
    .RESET_B(net3982),
    .D(_01532_),
    .Q_N(_09477_),
    .Q(\spiking_network_top_uut.all_data_out[771] ));
 sg13g2_dfrbp_1 _20217_ (.CLK(net4672),
    .RESET_B(net3991),
    .D(_01533_),
    .Q_N(_09476_),
    .Q(\spiking_network_top_uut.all_data_out[772] ));
 sg13g2_dfrbp_1 _20218_ (.CLK(net4672),
    .RESET_B(net3991),
    .D(_01534_),
    .Q_N(_00226_),
    .Q(\spiking_network_top_uut.all_data_out[773] ));
 sg13g2_dfrbp_1 _20219_ (.CLK(net4671),
    .RESET_B(net3990),
    .D(_01535_),
    .Q_N(_00156_),
    .Q(\spiking_network_top_uut.all_data_out[774] ));
 sg13g2_dfrbp_1 _20220_ (.CLK(net4662),
    .RESET_B(net3982),
    .D(_01536_),
    .Q_N(_09475_),
    .Q(\spiking_network_top_uut.all_data_out[775] ));
 sg13g2_dfrbp_1 _20221_ (.CLK(net4699),
    .RESET_B(net4019),
    .D(_01537_),
    .Q_N(_09474_),
    .Q(\spiking_network_top_uut.all_data_out[248] ));
 sg13g2_dfrbp_1 _20222_ (.CLK(net4693),
    .RESET_B(net4012),
    .D(_01538_),
    .Q_N(_09473_),
    .Q(\spiking_network_top_uut.all_data_out[249] ));
 sg13g2_dfrbp_1 _20223_ (.CLK(net4699),
    .RESET_B(net4019),
    .D(_01539_),
    .Q_N(_09472_),
    .Q(\spiking_network_top_uut.all_data_out[250] ));
 sg13g2_dfrbp_1 _20224_ (.CLK(net4693),
    .RESET_B(net4012),
    .D(_01540_),
    .Q_N(_09471_),
    .Q(\spiking_network_top_uut.all_data_out[251] ));
 sg13g2_dfrbp_1 _20225_ (.CLK(net4693),
    .RESET_B(net4012),
    .D(_01541_),
    .Q_N(_09470_),
    .Q(\spiking_network_top_uut.all_data_out[252] ));
 sg13g2_dfrbp_1 _20226_ (.CLK(net4693),
    .RESET_B(net4012),
    .D(_01542_),
    .Q_N(_09469_),
    .Q(\spiking_network_top_uut.all_data_out[253] ));
 sg13g2_dfrbp_1 _20227_ (.CLK(net4693),
    .RESET_B(net4012),
    .D(_01543_),
    .Q_N(_09468_),
    .Q(\spiking_network_top_uut.all_data_out[254] ));
 sg13g2_dfrbp_1 _20228_ (.CLK(net4699),
    .RESET_B(net4019),
    .D(_01544_),
    .Q_N(_09467_),
    .Q(\spiking_network_top_uut.all_data_out[255] ));
 sg13g2_dfrbp_1 _20229_ (.CLK(net4689),
    .RESET_B(net4008),
    .D(_01545_),
    .Q_N(_09466_),
    .Q(\spiking_network_top_uut.all_data_out[640] ));
 sg13g2_dfrbp_1 _20230_ (.CLK(net4683),
    .RESET_B(net4002),
    .D(_01546_),
    .Q_N(_00382_),
    .Q(\spiking_network_top_uut.all_data_out[641] ));
 sg13g2_dfrbp_1 _20231_ (.CLK(net4683),
    .RESET_B(net4011),
    .D(_01547_),
    .Q_N(_00312_),
    .Q(\spiking_network_top_uut.all_data_out[642] ));
 sg13g2_dfrbp_1 _20232_ (.CLK(net4656),
    .RESET_B(net3975),
    .D(_01548_),
    .Q_N(_09465_),
    .Q(\spiking_network_top_uut.all_data_out[643] ));
 sg13g2_dfrbp_1 _20233_ (.CLK(net4671),
    .RESET_B(net3990),
    .D(_01549_),
    .Q_N(_09464_),
    .Q(\spiking_network_top_uut.all_data_out[644] ));
 sg13g2_dfrbp_1 _20234_ (.CLK(net4672),
    .RESET_B(net3991),
    .D(_01550_),
    .Q_N(_00242_),
    .Q(\spiking_network_top_uut.all_data_out[645] ));
 sg13g2_dfrbp_1 _20235_ (.CLK(net4659),
    .RESET_B(net3978),
    .D(_01551_),
    .Q_N(_00172_),
    .Q(\spiking_network_top_uut.all_data_out[646] ));
 sg13g2_dfrbp_1 _20236_ (.CLK(net4659),
    .RESET_B(net3978),
    .D(_01552_),
    .Q_N(_09463_),
    .Q(\spiking_network_top_uut.all_data_out[647] ));
 sg13g2_dfrbp_1 _20237_ (.CLK(net4673),
    .RESET_B(net3992),
    .D(_01553_),
    .Q_N(_09462_),
    .Q(\spiking_network_top_uut.all_data_out[240] ));
 sg13g2_dfrbp_1 _20238_ (.CLK(net4676),
    .RESET_B(net3996),
    .D(_01554_),
    .Q_N(_09461_),
    .Q(\spiking_network_top_uut.all_data_out[241] ));
 sg13g2_dfrbp_1 _20239_ (.CLK(net4673),
    .RESET_B(net3992),
    .D(_01555_),
    .Q_N(_09460_),
    .Q(\spiking_network_top_uut.all_data_out[242] ));
 sg13g2_dfrbp_1 _20240_ (.CLK(net4673),
    .RESET_B(net3995),
    .D(_01556_),
    .Q_N(_09459_),
    .Q(\spiking_network_top_uut.all_data_out[243] ));
 sg13g2_dfrbp_1 _20241_ (.CLK(net4696),
    .RESET_B(net4015),
    .D(_01557_),
    .Q_N(_09458_),
    .Q(\spiking_network_top_uut.all_data_out[244] ));
 sg13g2_dfrbp_1 _20242_ (.CLK(net4699),
    .RESET_B(net4019),
    .D(_01558_),
    .Q_N(_09457_),
    .Q(\spiking_network_top_uut.all_data_out[245] ));
 sg13g2_dfrbp_1 _20243_ (.CLK(net4699),
    .RESET_B(net4019),
    .D(_01559_),
    .Q_N(_09456_),
    .Q(\spiking_network_top_uut.all_data_out[246] ));
 sg13g2_dfrbp_1 _20244_ (.CLK(net4699),
    .RESET_B(net4019),
    .D(_01560_),
    .Q_N(_09455_),
    .Q(\spiking_network_top_uut.all_data_out[247] ));
 sg13g2_dfrbp_1 _20245_ (.CLK(net4771),
    .RESET_B(net4092),
    .D(_01561_),
    .Q_N(_09454_),
    .Q(\spiking_network_top_uut.all_data_out[776] ));
 sg13g2_dfrbp_1 _20246_ (.CLK(net4771),
    .RESET_B(net4092),
    .D(_01562_),
    .Q_N(_00365_),
    .Q(\spiking_network_top_uut.all_data_out[777] ));
 sg13g2_dfrbp_1 _20247_ (.CLK(net4771),
    .RESET_B(net4092),
    .D(_01563_),
    .Q_N(_00295_),
    .Q(\spiking_network_top_uut.all_data_out[778] ));
 sg13g2_dfrbp_1 _20248_ (.CLK(net4747),
    .RESET_B(net4068),
    .D(_01564_),
    .Q_N(_09453_),
    .Q(\spiking_network_top_uut.all_data_out[779] ));
 sg13g2_dfrbp_1 _20249_ (.CLK(net4769),
    .RESET_B(net4090),
    .D(_01565_),
    .Q_N(_09452_),
    .Q(\spiking_network_top_uut.all_data_out[780] ));
 sg13g2_dfrbp_1 _20250_ (.CLK(net4769),
    .RESET_B(net4090),
    .D(_01566_),
    .Q_N(_00225_),
    .Q(\spiking_network_top_uut.all_data_out[781] ));
 sg13g2_dfrbp_1 _20251_ (.CLK(net4769),
    .RESET_B(net4090),
    .D(_01567_),
    .Q_N(_00155_),
    .Q(\spiking_network_top_uut.all_data_out[782] ));
 sg13g2_dfrbp_1 _20252_ (.CLK(net4768),
    .RESET_B(net4089),
    .D(_01568_),
    .Q_N(_09451_),
    .Q(\spiking_network_top_uut.all_data_out[783] ));
 sg13g2_dfrbp_1 _20253_ (.CLK(net4694),
    .RESET_B(net4013),
    .D(_01569_),
    .Q_N(_09450_),
    .Q(\spiking_network_top_uut.all_data_out[232] ));
 sg13g2_dfrbp_1 _20254_ (.CLK(net4694),
    .RESET_B(net4013),
    .D(_01570_),
    .Q_N(_09449_),
    .Q(\spiking_network_top_uut.all_data_out[233] ));
 sg13g2_dfrbp_1 _20255_ (.CLK(net4698),
    .RESET_B(net4018),
    .D(_01571_),
    .Q_N(_09448_),
    .Q(\spiking_network_top_uut.all_data_out[234] ));
 sg13g2_dfrbp_1 _20256_ (.CLK(net4694),
    .RESET_B(net4013),
    .D(_01572_),
    .Q_N(_09447_),
    .Q(\spiking_network_top_uut.all_data_out[235] ));
 sg13g2_dfrbp_1 _20257_ (.CLK(net4692),
    .RESET_B(net4011),
    .D(_01573_),
    .Q_N(_09446_),
    .Q(\spiking_network_top_uut.all_data_out[236] ));
 sg13g2_dfrbp_1 _20258_ (.CLK(net4698),
    .RESET_B(net4019),
    .D(_01574_),
    .Q_N(_09445_),
    .Q(\spiking_network_top_uut.all_data_out[237] ));
 sg13g2_dfrbp_1 _20259_ (.CLK(net4698),
    .RESET_B(net4018),
    .D(_01575_),
    .Q_N(_09444_),
    .Q(\spiking_network_top_uut.all_data_out[238] ));
 sg13g2_dfrbp_1 _20260_ (.CLK(net4694),
    .RESET_B(net4013),
    .D(_01576_),
    .Q_N(_09443_),
    .Q(\spiking_network_top_uut.all_data_out[239] ));
 sg13g2_dfrbp_1 _20261_ (.CLK(net4812),
    .RESET_B(net4134),
    .D(_01577_),
    .Q_N(_09442_),
    .Q(\spiking_network_top_uut.all_data_out[504] ));
 sg13g2_dfrbp_1 _20262_ (.CLK(net4809),
    .RESET_B(net4130),
    .D(_01578_),
    .Q_N(_00399_),
    .Q(\spiking_network_top_uut.all_data_out[505] ));
 sg13g2_dfrbp_1 _20263_ (.CLK(net4809),
    .RESET_B(net4130),
    .D(_01579_),
    .Q_N(_00329_),
    .Q(\spiking_network_top_uut.all_data_out[506] ));
 sg13g2_dfrbp_1 _20264_ (.CLK(net4750),
    .RESET_B(net4071),
    .D(_01580_),
    .Q_N(_09441_),
    .Q(\spiking_network_top_uut.all_data_out[507] ));
 sg13g2_dfrbp_1 _20265_ (.CLK(net4797),
    .RESET_B(net4118),
    .D(_01581_),
    .Q_N(_09440_),
    .Q(\spiking_network_top_uut.all_data_out[508] ));
 sg13g2_dfrbp_1 _20266_ (.CLK(net4797),
    .RESET_B(net4118),
    .D(_01582_),
    .Q_N(_00259_),
    .Q(\spiking_network_top_uut.all_data_out[509] ));
 sg13g2_dfrbp_1 _20267_ (.CLK(net4798),
    .RESET_B(net4120),
    .D(_01583_),
    .Q_N(_00189_),
    .Q(\spiking_network_top_uut.all_data_out[510] ));
 sg13g2_dfrbp_1 _20268_ (.CLK(net4750),
    .RESET_B(net4071),
    .D(_01584_),
    .Q_N(_09439_),
    .Q(\spiking_network_top_uut.all_data_out[511] ));
 sg13g2_dfrbp_1 _20269_ (.CLK(net4676),
    .RESET_B(net3995),
    .D(_01585_),
    .Q_N(_09438_),
    .Q(\spiking_network_top_uut.all_data_out[224] ));
 sg13g2_dfrbp_1 _20270_ (.CLK(net4676),
    .RESET_B(net3995),
    .D(_01586_),
    .Q_N(_09437_),
    .Q(\spiking_network_top_uut.all_data_out[225] ));
 sg13g2_dfrbp_1 _20271_ (.CLK(net4676),
    .RESET_B(net3995),
    .D(_01587_),
    .Q_N(_09436_),
    .Q(\spiking_network_top_uut.all_data_out[226] ));
 sg13g2_dfrbp_1 _20272_ (.CLK(net4676),
    .RESET_B(net3995),
    .D(_01588_),
    .Q_N(_09435_),
    .Q(\spiking_network_top_uut.all_data_out[227] ));
 sg13g2_dfrbp_1 _20273_ (.CLK(net4723),
    .RESET_B(net4043),
    .D(_01589_),
    .Q_N(_09434_),
    .Q(\spiking_network_top_uut.all_data_out[228] ));
 sg13g2_dfrbp_1 _20274_ (.CLK(net4701),
    .RESET_B(net4021),
    .D(_01590_),
    .Q_N(_09433_),
    .Q(\spiking_network_top_uut.all_data_out[229] ));
 sg13g2_dfrbp_1 _20275_ (.CLK(net4723),
    .RESET_B(net4043),
    .D(_01591_),
    .Q_N(_09432_),
    .Q(\spiking_network_top_uut.all_data_out[230] ));
 sg13g2_dfrbp_1 _20276_ (.CLK(net4726),
    .RESET_B(net4044),
    .D(_01592_),
    .Q_N(_09431_),
    .Q(\spiking_network_top_uut.all_data_out[231] ));
 sg13g2_dfrbp_1 _20277_ (.CLK(net4745),
    .RESET_B(net4066),
    .D(_01593_),
    .Q_N(_09430_),
    .Q(\spiking_network_top_uut.all_data_out[784] ));
 sg13g2_dfrbp_1 _20278_ (.CLK(net4745),
    .RESET_B(net4066),
    .D(_01594_),
    .Q_N(_00364_),
    .Q(\spiking_network_top_uut.all_data_out[785] ));
 sg13g2_dfrbp_1 _20279_ (.CLK(net4745),
    .RESET_B(net4066),
    .D(_01595_),
    .Q_N(_00294_),
    .Q(\spiking_network_top_uut.all_data_out[786] ));
 sg13g2_dfrbp_1 _20280_ (.CLK(net4748),
    .RESET_B(net4069),
    .D(_01596_),
    .Q_N(_09429_),
    .Q(\spiking_network_top_uut.all_data_out[787] ));
 sg13g2_dfrbp_1 _20281_ (.CLK(net4766),
    .RESET_B(net4087),
    .D(_01597_),
    .Q_N(_09428_),
    .Q(\spiking_network_top_uut.all_data_out[788] ));
 sg13g2_dfrbp_1 _20282_ (.CLK(net4766),
    .RESET_B(net4087),
    .D(_01598_),
    .Q_N(_00224_),
    .Q(\spiking_network_top_uut.all_data_out[789] ));
 sg13g2_dfrbp_1 _20283_ (.CLK(net4766),
    .RESET_B(net4087),
    .D(_01599_),
    .Q_N(_00154_),
    .Q(\spiking_network_top_uut.all_data_out[790] ));
 sg13g2_dfrbp_1 _20284_ (.CLK(net4747),
    .RESET_B(net4068),
    .D(_01600_),
    .Q_N(_09427_),
    .Q(\spiking_network_top_uut.all_data_out[791] ));
 sg13g2_dfrbp_1 _20285_ (.CLK(net4719),
    .RESET_B(net4040),
    .D(_01601_),
    .Q_N(_09426_),
    .Q(\spiking_network_top_uut.all_data_out[216] ));
 sg13g2_dfrbp_1 _20286_ (.CLK(net4742),
    .RESET_B(net4063),
    .D(_01602_),
    .Q_N(_09425_),
    .Q(\spiking_network_top_uut.all_data_out[217] ));
 sg13g2_dfrbp_1 _20287_ (.CLK(net4719),
    .RESET_B(net4040),
    .D(_01603_),
    .Q_N(_09424_),
    .Q(\spiking_network_top_uut.all_data_out[218] ));
 sg13g2_dfrbp_1 _20288_ (.CLK(net4719),
    .RESET_B(net4040),
    .D(_01604_),
    .Q_N(_09423_),
    .Q(\spiking_network_top_uut.all_data_out[219] ));
 sg13g2_dfrbp_1 _20289_ (.CLK(net4742),
    .RESET_B(net4063),
    .D(_01605_),
    .Q_N(_09422_),
    .Q(\spiking_network_top_uut.all_data_out[220] ));
 sg13g2_dfrbp_1 _20290_ (.CLK(net4719),
    .RESET_B(net4040),
    .D(_01606_),
    .Q_N(_09421_),
    .Q(\spiking_network_top_uut.all_data_out[221] ));
 sg13g2_dfrbp_1 _20291_ (.CLK(net4742),
    .RESET_B(net4063),
    .D(_01607_),
    .Q_N(_09420_),
    .Q(\spiking_network_top_uut.all_data_out[222] ));
 sg13g2_dfrbp_1 _20292_ (.CLK(net4743),
    .RESET_B(net4062),
    .D(_01608_),
    .Q_N(_09419_),
    .Q(\spiking_network_top_uut.all_data_out[223] ));
 sg13g2_dfrbp_1 _20293_ (.CLK(net4683),
    .RESET_B(net4002),
    .D(_01609_),
    .Q_N(_09418_),
    .Q(\spiking_network_top_uut.all_data_out[608] ));
 sg13g2_dfrbp_1 _20294_ (.CLK(net4689),
    .RESET_B(net4008),
    .D(_01610_),
    .Q_N(_00386_),
    .Q(\spiking_network_top_uut.all_data_out[609] ));
 sg13g2_dfrbp_1 _20295_ (.CLK(net4689),
    .RESET_B(net4008),
    .D(_01611_),
    .Q_N(_00316_),
    .Q(\spiking_network_top_uut.all_data_out[610] ));
 sg13g2_dfrbp_1 _20296_ (.CLK(net4683),
    .RESET_B(net4002),
    .D(_01612_),
    .Q_N(_09417_),
    .Q(\spiking_network_top_uut.all_data_out[611] ));
 sg13g2_dfrbp_1 _20297_ (.CLK(net4692),
    .RESET_B(net4011),
    .D(_01613_),
    .Q_N(_09416_),
    .Q(\spiking_network_top_uut.all_data_out[612] ));
 sg13g2_dfrbp_1 _20298_ (.CLK(net4674),
    .RESET_B(net3993),
    .D(_01614_),
    .Q_N(_00246_),
    .Q(\spiking_network_top_uut.all_data_out[613] ));
 sg13g2_dfrbp_1 _20299_ (.CLK(net4674),
    .RESET_B(net3993),
    .D(_01615_),
    .Q_N(_00176_),
    .Q(\spiking_network_top_uut.all_data_out[614] ));
 sg13g2_dfrbp_1 _20300_ (.CLK(net4694),
    .RESET_B(net4013),
    .D(_01616_),
    .Q_N(_09415_),
    .Q(\spiking_network_top_uut.all_data_out[615] ));
 sg13g2_dfrbp_1 _20301_ (.CLK(net4682),
    .RESET_B(net4001),
    .D(_01617_),
    .Q_N(_09414_),
    .Q(\spiking_network_top_uut.all_data_out[208] ));
 sg13g2_dfrbp_1 _20302_ (.CLK(net4684),
    .RESET_B(net4003),
    .D(_01618_),
    .Q_N(_09413_),
    .Q(\spiking_network_top_uut.all_data_out[209] ));
 sg13g2_dfrbp_1 _20303_ (.CLK(net4684),
    .RESET_B(net4002),
    .D(_01619_),
    .Q_N(_09412_),
    .Q(\spiking_network_top_uut.all_data_out[210] ));
 sg13g2_dfrbp_1 _20304_ (.CLK(net4681),
    .RESET_B(net4000),
    .D(_01620_),
    .Q_N(_09411_),
    .Q(\spiking_network_top_uut.all_data_out[211] ));
 sg13g2_dfrbp_1 _20305_ (.CLK(net4721),
    .RESET_B(net4042),
    .D(_01621_),
    .Q_N(_09410_),
    .Q(\spiking_network_top_uut.all_data_out[212] ));
 sg13g2_dfrbp_1 _20306_ (.CLK(net4721),
    .RESET_B(net4041),
    .D(_01622_),
    .Q_N(_09409_),
    .Q(\spiking_network_top_uut.all_data_out[213] ));
 sg13g2_dfrbp_1 _20307_ (.CLK(net4732),
    .RESET_B(net4052),
    .D(_01623_),
    .Q_N(_09408_),
    .Q(\spiking_network_top_uut.all_data_out[214] ));
 sg13g2_dfrbp_1 _20308_ (.CLK(net4733),
    .RESET_B(net4053),
    .D(_01624_),
    .Q_N(_09407_),
    .Q(\spiking_network_top_uut.all_data_out[215] ));
 sg13g2_dfrbp_1 _20309_ (.CLK(net4715),
    .RESET_B(net4035),
    .D(_01625_),
    .Q_N(_09406_),
    .Q(\spiking_network_top_uut.all_data_out[792] ));
 sg13g2_dfrbp_1 _20310_ (.CLK(net4715),
    .RESET_B(net4035),
    .D(_01626_),
    .Q_N(_00363_),
    .Q(\spiking_network_top_uut.all_data_out[793] ));
 sg13g2_dfrbp_1 _20311_ (.CLK(net4715),
    .RESET_B(net4035),
    .D(_01627_),
    .Q_N(_00293_),
    .Q(\spiking_network_top_uut.all_data_out[794] ));
 sg13g2_dfrbp_1 _20312_ (.CLK(net4739),
    .RESET_B(net4063),
    .D(_01628_),
    .Q_N(_09405_),
    .Q(\spiking_network_top_uut.all_data_out[795] ));
 sg13g2_dfrbp_1 _20313_ (.CLK(net4739),
    .RESET_B(net4060),
    .D(_01629_),
    .Q_N(_09404_),
    .Q(\spiking_network_top_uut.all_data_out[796] ));
 sg13g2_dfrbp_1 _20314_ (.CLK(net4741),
    .RESET_B(net4061),
    .D(_01630_),
    .Q_N(_00223_),
    .Q(\spiking_network_top_uut.all_data_out[797] ));
 sg13g2_dfrbp_1 _20315_ (.CLK(net4739),
    .RESET_B(net4060),
    .D(_01631_),
    .Q_N(_00153_),
    .Q(\spiking_network_top_uut.all_data_out[798] ));
 sg13g2_dfrbp_1 _20316_ (.CLK(net4720),
    .RESET_B(net4041),
    .D(_01632_),
    .Q_N(_09403_),
    .Q(\spiking_network_top_uut.all_data_out[799] ));
 sg13g2_dfrbp_1 _20317_ (.CLK(net4668),
    .RESET_B(net3993),
    .D(_01633_),
    .Q_N(_09402_),
    .Q(\spiking_network_top_uut.all_data_out[200] ));
 sg13g2_dfrbp_1 _20318_ (.CLK(net4674),
    .RESET_B(net3993),
    .D(_01634_),
    .Q_N(_09401_),
    .Q(\spiking_network_top_uut.all_data_out[201] ));
 sg13g2_dfrbp_1 _20319_ (.CLK(net4666),
    .RESET_B(net3986),
    .D(_01635_),
    .Q_N(_09400_),
    .Q(\spiking_network_top_uut.all_data_out[202] ));
 sg13g2_dfrbp_1 _20320_ (.CLK(net4672),
    .RESET_B(net3991),
    .D(_01636_),
    .Q_N(_09399_),
    .Q(\spiking_network_top_uut.all_data_out[203] ));
 sg13g2_dfrbp_1 _20321_ (.CLK(net4673),
    .RESET_B(net3992),
    .D(_01637_),
    .Q_N(_09398_),
    .Q(\spiking_network_top_uut.all_data_out[204] ));
 sg13g2_dfrbp_1 _20322_ (.CLK(net4672),
    .RESET_B(net3991),
    .D(_01638_),
    .Q_N(_09397_),
    .Q(\spiking_network_top_uut.all_data_out[205] ));
 sg13g2_dfrbp_1 _20323_ (.CLK(net4673),
    .RESET_B(net3992),
    .D(_01639_),
    .Q_N(_09396_),
    .Q(\spiking_network_top_uut.all_data_out[206] ));
 sg13g2_dfrbp_1 _20324_ (.CLK(net4666),
    .RESET_B(net3986),
    .D(_01640_),
    .Q_N(_09395_),
    .Q(\spiking_network_top_uut.all_data_out[207] ));
 sg13g2_dfrbp_1 _20325_ (.CLK(net4780),
    .RESET_B(net4102),
    .D(_01641_),
    .Q_N(_09394_),
    .Q(\spiking_network_top_uut.all_data_out[496] ));
 sg13g2_dfrbp_1 _20326_ (.CLK(net4762),
    .RESET_B(net4083),
    .D(_01642_),
    .Q_N(_00400_),
    .Q(\spiking_network_top_uut.all_data_out[497] ));
 sg13g2_dfrbp_1 _20327_ (.CLK(net4762),
    .RESET_B(net4083),
    .D(_01643_),
    .Q_N(_00330_),
    .Q(\spiking_network_top_uut.all_data_out[498] ));
 sg13g2_dfrbp_1 _20328_ (.CLK(net4762),
    .RESET_B(net4083),
    .D(_01644_),
    .Q_N(_09393_),
    .Q(\spiking_network_top_uut.all_data_out[499] ));
 sg13g2_dfrbp_1 _20329_ (.CLK(net4753),
    .RESET_B(net4074),
    .D(_01645_),
    .Q_N(_09392_),
    .Q(\spiking_network_top_uut.all_data_out[500] ));
 sg13g2_dfrbp_1 _20330_ (.CLK(net4754),
    .RESET_B(net4075),
    .D(_01646_),
    .Q_N(_00260_),
    .Q(\spiking_network_top_uut.all_data_out[501] ));
 sg13g2_dfrbp_1 _20331_ (.CLK(net4753),
    .RESET_B(net4075),
    .D(_01647_),
    .Q_N(_00190_),
    .Q(\spiking_network_top_uut.all_data_out[502] ));
 sg13g2_dfrbp_1 _20332_ (.CLK(net4761),
    .RESET_B(net4082),
    .D(_01648_),
    .Q_N(_09391_),
    .Q(\spiking_network_top_uut.all_data_out[503] ));
 sg13g2_dfrbp_1 _20333_ (.CLK(net4661),
    .RESET_B(net3981),
    .D(_01649_),
    .Q_N(_09390_),
    .Q(\spiking_network_top_uut.all_data_out[192] ));
 sg13g2_dfrbp_1 _20334_ (.CLK(net4656),
    .RESET_B(net3975),
    .D(_01650_),
    .Q_N(_09389_),
    .Q(\spiking_network_top_uut.all_data_out[193] ));
 sg13g2_dfrbp_1 _20335_ (.CLK(net4661),
    .RESET_B(net3981),
    .D(_01651_),
    .Q_N(_09388_),
    .Q(\spiking_network_top_uut.all_data_out[194] ));
 sg13g2_dfrbp_1 _20336_ (.CLK(net4661),
    .RESET_B(net3981),
    .D(_01652_),
    .Q_N(_09387_),
    .Q(\spiking_network_top_uut.all_data_out[195] ));
 sg13g2_dfrbp_1 _20337_ (.CLK(net4666),
    .RESET_B(net3986),
    .D(_01653_),
    .Q_N(_09386_),
    .Q(\spiking_network_top_uut.all_data_out[196] ));
 sg13g2_dfrbp_1 _20338_ (.CLK(net4667),
    .RESET_B(net3987),
    .D(_01654_),
    .Q_N(_09385_),
    .Q(\spiking_network_top_uut.all_data_out[197] ));
 sg13g2_dfrbp_1 _20339_ (.CLK(net4666),
    .RESET_B(net3986),
    .D(_01655_),
    .Q_N(_09384_),
    .Q(\spiking_network_top_uut.all_data_out[198] ));
 sg13g2_dfrbp_1 _20340_ (.CLK(net4666),
    .RESET_B(net3986),
    .D(_01656_),
    .Q_N(_09383_),
    .Q(\spiking_network_top_uut.all_data_out[199] ));
 sg13g2_dfrbp_1 _20341_ (.CLK(net4686),
    .RESET_B(net4008),
    .D(_01657_),
    .Q_N(_09382_),
    .Q(\spiking_network_top_uut.all_data_out[800] ));
 sg13g2_dfrbp_1 _20342_ (.CLK(net4689),
    .RESET_B(net4008),
    .D(_01658_),
    .Q_N(_00362_),
    .Q(\spiking_network_top_uut.all_data_out[801] ));
 sg13g2_dfrbp_1 _20343_ (.CLK(net4683),
    .RESET_B(net4002),
    .D(_01659_),
    .Q_N(_00292_),
    .Q(\spiking_network_top_uut.all_data_out[802] ));
 sg13g2_dfrbp_1 _20344_ (.CLK(net4671),
    .RESET_B(net3990),
    .D(_01660_),
    .Q_N(_09381_),
    .Q(\spiking_network_top_uut.all_data_out[803] ));
 sg13g2_dfrbp_1 _20345_ (.CLK(net4671),
    .RESET_B(net3990),
    .D(_01661_),
    .Q_N(_09380_),
    .Q(\spiking_network_top_uut.all_data_out[804] ));
 sg13g2_dfrbp_1 _20346_ (.CLK(net4672),
    .RESET_B(net3991),
    .D(_01662_),
    .Q_N(_00222_),
    .Q(\spiking_network_top_uut.all_data_out[805] ));
 sg13g2_dfrbp_1 _20347_ (.CLK(net4673),
    .RESET_B(net3992),
    .D(_01663_),
    .Q_N(_00152_),
    .Q(\spiking_network_top_uut.all_data_out[806] ));
 sg13g2_dfrbp_1 _20348_ (.CLK(net4656),
    .RESET_B(net3975),
    .D(_01664_),
    .Q_N(_09379_),
    .Q(\spiking_network_top_uut.all_data_out[807] ));
 sg13g2_dfrbp_1 _20349_ (.CLK(net4712),
    .RESET_B(net4032),
    .D(_01665_),
    .Q_N(_09378_),
    .Q(\spiking_network_top_uut.all_data_out[184] ));
 sg13g2_dfrbp_1 _20350_ (.CLK(net4687),
    .RESET_B(net4006),
    .D(_01666_),
    .Q_N(_09377_),
    .Q(\spiking_network_top_uut.all_data_out[185] ));
 sg13g2_dfrbp_1 _20351_ (.CLK(net4712),
    .RESET_B(net4032),
    .D(_01667_),
    .Q_N(_09376_),
    .Q(\spiking_network_top_uut.all_data_out[186] ));
 sg13g2_dfrbp_1 _20352_ (.CLK(net4687),
    .RESET_B(net4006),
    .D(_01668_),
    .Q_N(_09375_),
    .Q(\spiking_network_top_uut.all_data_out[187] ));
 sg13g2_dfrbp_1 _20353_ (.CLK(net4725),
    .RESET_B(net4045),
    .D(_01669_),
    .Q_N(_09374_),
    .Q(\spiking_network_top_uut.all_data_out[188] ));
 sg13g2_dfrbp_1 _20354_ (.CLK(net4724),
    .RESET_B(net4044),
    .D(_01670_),
    .Q_N(_09373_),
    .Q(\spiking_network_top_uut.all_data_out[189] ));
 sg13g2_dfrbp_1 _20355_ (.CLK(net4700),
    .RESET_B(net4020),
    .D(_01671_),
    .Q_N(_09372_),
    .Q(\spiking_network_top_uut.all_data_out[190] ));
 sg13g2_dfrbp_1 _20356_ (.CLK(net4724),
    .RESET_B(net4044),
    .D(_01672_),
    .Q_N(_09371_),
    .Q(\spiking_network_top_uut.all_data_out[191] ));
 sg13g2_dfrbp_1 _20357_ (.CLK(net4770),
    .RESET_B(net4091),
    .D(_01673_),
    .Q_N(_09370_),
    .Q(\spiking_network_top_uut.all_data_out[648] ));
 sg13g2_dfrbp_1 _20358_ (.CLK(net4776),
    .RESET_B(net4097),
    .D(_01674_),
    .Q_N(_00381_),
    .Q(\spiking_network_top_uut.all_data_out[649] ));
 sg13g2_dfrbp_1 _20359_ (.CLK(net4770),
    .RESET_B(net4091),
    .D(_01675_),
    .Q_N(_00311_),
    .Q(\spiking_network_top_uut.all_data_out[650] ));
 sg13g2_dfrbp_1 _20360_ (.CLK(net4772),
    .RESET_B(net4093),
    .D(_01676_),
    .Q_N(_09369_),
    .Q(\spiking_network_top_uut.all_data_out[651] ));
 sg13g2_dfrbp_1 _20361_ (.CLK(net4784),
    .RESET_B(net4106),
    .D(_01677_),
    .Q_N(_09368_),
    .Q(\spiking_network_top_uut.all_data_out[652] ));
 sg13g2_dfrbp_1 _20362_ (.CLK(net4779),
    .RESET_B(net4100),
    .D(_01678_),
    .Q_N(_00241_),
    .Q(\spiking_network_top_uut.all_data_out[653] ));
 sg13g2_dfrbp_1 _20363_ (.CLK(net4779),
    .RESET_B(net4100),
    .D(_01679_),
    .Q_N(_00171_),
    .Q(\spiking_network_top_uut.all_data_out[654] ));
 sg13g2_dfrbp_1 _20364_ (.CLK(net4778),
    .RESET_B(net4099),
    .D(_01680_),
    .Q_N(_09367_),
    .Q(\spiking_network_top_uut.all_data_out[655] ));
 sg13g2_dfrbp_1 _20365_ (.CLK(net4688),
    .RESET_B(net4007),
    .D(_01681_),
    .Q_N(_09366_),
    .Q(\spiking_network_top_uut.all_data_out[176] ));
 sg13g2_dfrbp_1 _20366_ (.CLK(net4698),
    .RESET_B(net4018),
    .D(_01682_),
    .Q_N(_09365_),
    .Q(\spiking_network_top_uut.all_data_out[177] ));
 sg13g2_dfrbp_1 _20367_ (.CLK(net4688),
    .RESET_B(net4007),
    .D(_01683_),
    .Q_N(_09364_),
    .Q(\spiking_network_top_uut.all_data_out[178] ));
 sg13g2_dfrbp_1 _20368_ (.CLK(net4688),
    .RESET_B(net4020),
    .D(_01684_),
    .Q_N(_09363_),
    .Q(\spiking_network_top_uut.all_data_out[179] ));
 sg13g2_dfrbp_1 _20369_ (.CLK(net4724),
    .RESET_B(net4044),
    .D(_01685_),
    .Q_N(_09362_),
    .Q(\spiking_network_top_uut.all_data_out[180] ));
 sg13g2_dfrbp_1 _20370_ (.CLK(net4712),
    .RESET_B(net4032),
    .D(_01686_),
    .Q_N(_09361_),
    .Q(\spiking_network_top_uut.all_data_out[181] ));
 sg13g2_dfrbp_1 _20371_ (.CLK(net4724),
    .RESET_B(net4044),
    .D(_01687_),
    .Q_N(_09360_),
    .Q(\spiking_network_top_uut.all_data_out[182] ));
 sg13g2_dfrbp_1 _20372_ (.CLK(net4688),
    .RESET_B(net4006),
    .D(_01688_),
    .Q_N(_09359_),
    .Q(\spiking_network_top_uut.all_data_out[183] ));
 sg13g2_dfrbp_1 _20373_ (.CLK(net4771),
    .RESET_B(net4092),
    .D(_01689_),
    .Q_N(_09358_),
    .Q(\spiking_network_top_uut.all_data_out[808] ));
 sg13g2_dfrbp_1 _20374_ (.CLK(net4771),
    .RESET_B(net4092),
    .D(_01690_),
    .Q_N(_00361_),
    .Q(\spiking_network_top_uut.all_data_out[809] ));
 sg13g2_dfrbp_1 _20375_ (.CLK(net4771),
    .RESET_B(net4092),
    .D(_01691_),
    .Q_N(_00291_),
    .Q(\spiking_network_top_uut.all_data_out[810] ));
 sg13g2_dfrbp_1 _20376_ (.CLK(net4772),
    .RESET_B(net4093),
    .D(_01692_),
    .Q_N(_09357_),
    .Q(\spiking_network_top_uut.all_data_out[811] ));
 sg13g2_dfrbp_1 _20377_ (.CLK(net4772),
    .RESET_B(net4096),
    .D(_01693_),
    .Q_N(_09356_),
    .Q(\spiking_network_top_uut.all_data_out[812] ));
 sg13g2_dfrbp_1 _20378_ (.CLK(net4769),
    .RESET_B(net4090),
    .D(_01694_),
    .Q_N(_00221_),
    .Q(\spiking_network_top_uut.all_data_out[813] ));
 sg13g2_dfrbp_1 _20379_ (.CLK(net4769),
    .RESET_B(net4090),
    .D(_01695_),
    .Q_N(_00151_),
    .Q(\spiking_network_top_uut.all_data_out[814] ));
 sg13g2_dfrbp_1 _20380_ (.CLK(net4757),
    .RESET_B(net4078),
    .D(_01696_),
    .Q_N(_09355_),
    .Q(\spiking_network_top_uut.all_data_out[815] ));
 sg13g2_dfrbp_1 _20381_ (.CLK(net4687),
    .RESET_B(net4006),
    .D(_01697_),
    .Q_N(_09354_),
    .Q(\spiking_network_top_uut.all_data_out[168] ));
 sg13g2_dfrbp_1 _20382_ (.CLK(net4687),
    .RESET_B(net4006),
    .D(_01698_),
    .Q_N(_09353_),
    .Q(\spiking_network_top_uut.all_data_out[169] ));
 sg13g2_dfrbp_1 _20383_ (.CLK(net4712),
    .RESET_B(net4032),
    .D(_01699_),
    .Q_N(_09352_),
    .Q(\spiking_network_top_uut.all_data_out[170] ));
 sg13g2_dfrbp_1 _20384_ (.CLK(net4688),
    .RESET_B(net4007),
    .D(_01700_),
    .Q_N(_09351_),
    .Q(\spiking_network_top_uut.all_data_out[171] ));
 sg13g2_dfrbp_1 _20385_ (.CLK(net4713),
    .RESET_B(net4034),
    .D(_01701_),
    .Q_N(_09350_),
    .Q(\spiking_network_top_uut.all_data_out[172] ));
 sg13g2_dfrbp_1 _20386_ (.CLK(net4712),
    .RESET_B(net4032),
    .D(_01702_),
    .Q_N(_09349_),
    .Q(\spiking_network_top_uut.all_data_out[173] ));
 sg13g2_dfrbp_1 _20387_ (.CLK(net4712),
    .RESET_B(net4032),
    .D(_01703_),
    .Q_N(_09348_),
    .Q(\spiking_network_top_uut.all_data_out[174] ));
 sg13g2_dfrbp_1 _20388_ (.CLK(net4713),
    .RESET_B(net4033),
    .D(_01704_),
    .Q_N(_09347_),
    .Q(\spiking_network_top_uut.all_data_out[175] ));
 sg13g2_dfrbp_1 _20389_ (.CLK(net4789),
    .RESET_B(net4111),
    .D(_01705_),
    .Q_N(_09346_),
    .Q(\spiking_network_top_uut.all_data_out[488] ));
 sg13g2_dfrbp_1 _20390_ (.CLK(net4789),
    .RESET_B(net4111),
    .D(_01706_),
    .Q_N(_00401_),
    .Q(\spiking_network_top_uut.all_data_out[489] ));
 sg13g2_dfrbp_1 _20391_ (.CLK(net4789),
    .RESET_B(net4112),
    .D(_01707_),
    .Q_N(_00331_),
    .Q(\spiking_network_top_uut.all_data_out[490] ));
 sg13g2_dfrbp_1 _20392_ (.CLK(net4773),
    .RESET_B(net4094),
    .D(_01708_),
    .Q_N(_09345_),
    .Q(\spiking_network_top_uut.all_data_out[491] ));
 sg13g2_dfrbp_1 _20393_ (.CLK(net4796),
    .RESET_B(net4117),
    .D(_01709_),
    .Q_N(_09344_),
    .Q(\spiking_network_top_uut.all_data_out[492] ));
 sg13g2_dfrbp_1 _20394_ (.CLK(net4799),
    .RESET_B(net4119),
    .D(_01710_),
    .Q_N(_00261_),
    .Q(\spiking_network_top_uut.all_data_out[493] ));
 sg13g2_dfrbp_1 _20395_ (.CLK(net4799),
    .RESET_B(net4119),
    .D(_01711_),
    .Q_N(_00191_),
    .Q(\spiking_network_top_uut.all_data_out[494] ));
 sg13g2_dfrbp_1 _20396_ (.CLK(net4793),
    .RESET_B(net4115),
    .D(_01712_),
    .Q_N(_09343_),
    .Q(\spiking_network_top_uut.all_data_out[495] ));
 sg13g2_dfrbp_1 _20397_ (.CLK(net4714),
    .RESET_B(net4034),
    .D(_01713_),
    .Q_N(_09342_),
    .Q(\spiking_network_top_uut.all_data_out[160] ));
 sg13g2_dfrbp_1 _20398_ (.CLK(net4692),
    .RESET_B(net4012),
    .D(_01714_),
    .Q_N(_09341_),
    .Q(\spiking_network_top_uut.all_data_out[161] ));
 sg13g2_dfrbp_1 _20399_ (.CLK(net4689),
    .RESET_B(net4008),
    .D(_01715_),
    .Q_N(_09340_),
    .Q(\spiking_network_top_uut.all_data_out[162] ));
 sg13g2_dfrbp_1 _20400_ (.CLK(net4692),
    .RESET_B(net4012),
    .D(_01716_),
    .Q_N(_09339_),
    .Q(\spiking_network_top_uut.all_data_out[163] ));
 sg13g2_dfrbp_1 _20401_ (.CLK(net4700),
    .RESET_B(net4020),
    .D(_01717_),
    .Q_N(_09338_),
    .Q(\spiking_network_top_uut.all_data_out[164] ));
 sg13g2_dfrbp_1 _20402_ (.CLK(net4700),
    .RESET_B(net4020),
    .D(_01718_),
    .Q_N(_09337_),
    .Q(\spiking_network_top_uut.all_data_out[165] ));
 sg13g2_dfrbp_1 _20403_ (.CLK(net4700),
    .RESET_B(net4020),
    .D(_01719_),
    .Q_N(_09336_),
    .Q(\spiking_network_top_uut.all_data_out[166] ));
 sg13g2_dfrbp_1 _20404_ (.CLK(net4687),
    .RESET_B(net4007),
    .D(_01720_),
    .Q_N(_09335_),
    .Q(\spiking_network_top_uut.all_data_out[167] ));
 sg13g2_dfrbp_1 _20405_ (.CLK(net4744),
    .RESET_B(net4065),
    .D(_01721_),
    .Q_N(_09334_),
    .Q(\spiking_network_top_uut.all_data_out[816] ));
 sg13g2_dfrbp_1 _20406_ (.CLK(net4740),
    .RESET_B(net4061),
    .D(_01722_),
    .Q_N(_00360_),
    .Q(\spiking_network_top_uut.all_data_out[817] ));
 sg13g2_dfrbp_1 _20407_ (.CLK(net4740),
    .RESET_B(net4061),
    .D(_01723_),
    .Q_N(_00290_),
    .Q(\spiking_network_top_uut.all_data_out[818] ));
 sg13g2_dfrbp_1 _20408_ (.CLK(net4747),
    .RESET_B(net4068),
    .D(_01724_),
    .Q_N(_09333_),
    .Q(\spiking_network_top_uut.all_data_out[819] ));
 sg13g2_dfrbp_1 _20409_ (.CLK(net4765),
    .RESET_B(net4086),
    .D(_01725_),
    .Q_N(_09332_),
    .Q(\spiking_network_top_uut.all_data_out[820] ));
 sg13g2_dfrbp_1 _20410_ (.CLK(net4769),
    .RESET_B(net4090),
    .D(_01726_),
    .Q_N(_00220_),
    .Q(\spiking_network_top_uut.all_data_out[821] ));
 sg13g2_dfrbp_1 _20411_ (.CLK(net4765),
    .RESET_B(net4086),
    .D(_01727_),
    .Q_N(_00150_),
    .Q(\spiking_network_top_uut.all_data_out[822] ));
 sg13g2_dfrbp_1 _20412_ (.CLK(net4740),
    .RESET_B(net4062),
    .D(_01728_),
    .Q_N(_09331_),
    .Q(\spiking_network_top_uut.all_data_out[823] ));
 sg13g2_dfrbp_1 _20413_ (.CLK(net4703),
    .RESET_B(net4023),
    .D(_01729_),
    .Q_N(_09330_),
    .Q(\spiking_network_top_uut.all_data_out[152] ));
 sg13g2_dfrbp_1 _20414_ (.CLK(net4695),
    .RESET_B(net4014),
    .D(_01730_),
    .Q_N(_09329_),
    .Q(\spiking_network_top_uut.all_data_out[153] ));
 sg13g2_dfrbp_1 _20415_ (.CLK(net4695),
    .RESET_B(net4015),
    .D(_01731_),
    .Q_N(_09328_),
    .Q(\spiking_network_top_uut.all_data_out[154] ));
 sg13g2_dfrbp_1 _20416_ (.CLK(net4696),
    .RESET_B(net4014),
    .D(_01732_),
    .Q_N(_09327_),
    .Q(\spiking_network_top_uut.all_data_out[155] ));
 sg13g2_dfrbp_1 _20417_ (.CLK(net4696),
    .RESET_B(net4014),
    .D(_01733_),
    .Q_N(_09326_),
    .Q(\spiking_network_top_uut.all_data_out[156] ));
 sg13g2_dfrbp_1 _20418_ (.CLK(net4703),
    .RESET_B(net4023),
    .D(_01734_),
    .Q_N(_09325_),
    .Q(\spiking_network_top_uut.all_data_out[157] ));
 sg13g2_dfrbp_1 _20419_ (.CLK(net4697),
    .RESET_B(net4016),
    .D(_01735_),
    .Q_N(_09324_),
    .Q(\spiking_network_top_uut.all_data_out[158] ));
 sg13g2_dfrbp_1 _20420_ (.CLK(net4695),
    .RESET_B(net4014),
    .D(_01736_),
    .Q_N(_09323_),
    .Q(\spiking_network_top_uut.all_data_out[159] ));
 sg13g2_dfrbp_1 _20421_ (.CLK(net4809),
    .RESET_B(net4130),
    .D(_01737_),
    .Q_N(_09322_),
    .Q(\spiking_network_top_uut.all_data_out[568] ));
 sg13g2_dfrbp_1 _20422_ (.CLK(net4807),
    .RESET_B(net4132),
    .D(_01738_),
    .Q_N(_00391_),
    .Q(\spiking_network_top_uut.all_data_out[569] ));
 sg13g2_dfrbp_1 _20423_ (.CLK(net4807),
    .RESET_B(net4132),
    .D(_01739_),
    .Q_N(_00321_),
    .Q(\spiking_network_top_uut.all_data_out[570] ));
 sg13g2_dfrbp_1 _20424_ (.CLK(net4750),
    .RESET_B(net4071),
    .D(_01740_),
    .Q_N(_09321_),
    .Q(\spiking_network_top_uut.all_data_out[571] ));
 sg13g2_dfrbp_1 _20425_ (.CLK(net4807),
    .RESET_B(net4132),
    .D(_01741_),
    .Q_N(_09320_),
    .Q(\spiking_network_top_uut.all_data_out[572] ));
 sg13g2_dfrbp_1 _20426_ (.CLK(net4807),
    .RESET_B(net4132),
    .D(_01742_),
    .Q_N(_00251_),
    .Q(\spiking_network_top_uut.all_data_out[573] ));
 sg13g2_dfrbp_1 _20427_ (.CLK(net4808),
    .RESET_B(net4129),
    .D(_01743_),
    .Q_N(_00181_),
    .Q(\spiking_network_top_uut.all_data_out[574] ));
 sg13g2_dfrbp_1 _20428_ (.CLK(net4750),
    .RESET_B(net4071),
    .D(_01744_),
    .Q_N(_09319_),
    .Q(\spiking_network_top_uut.all_data_out[575] ));
 sg13g2_dfrbp_1 _20429_ (.CLK(net4666),
    .RESET_B(net3992),
    .D(_01745_),
    .Q_N(_09318_),
    .Q(\spiking_network_top_uut.all_data_out[144] ));
 sg13g2_dfrbp_1 _20430_ (.CLK(net4673),
    .RESET_B(net3992),
    .D(_01746_),
    .Q_N(_09317_),
    .Q(\spiking_network_top_uut.all_data_out[145] ));
 sg13g2_dfrbp_1 _20431_ (.CLK(net4668),
    .RESET_B(net3988),
    .D(_01747_),
    .Q_N(_09316_),
    .Q(\spiking_network_top_uut.all_data_out[146] ));
 sg13g2_dfrbp_1 _20432_ (.CLK(net4671),
    .RESET_B(net3990),
    .D(_01748_),
    .Q_N(_09315_),
    .Q(\spiking_network_top_uut.all_data_out[147] ));
 sg13g2_dfrbp_1 _20433_ (.CLK(net4668),
    .RESET_B(net3988),
    .D(_01749_),
    .Q_N(_09314_),
    .Q(\spiking_network_top_uut.all_data_out[148] ));
 sg13g2_dfrbp_1 _20434_ (.CLK(net4683),
    .RESET_B(net4011),
    .D(_01750_),
    .Q_N(_09313_),
    .Q(\spiking_network_top_uut.all_data_out[149] ));
 sg13g2_dfrbp_1 _20435_ (.CLK(net4692),
    .RESET_B(net4011),
    .D(_01751_),
    .Q_N(_09312_),
    .Q(\spiking_network_top_uut.all_data_out[150] ));
 sg13g2_dfrbp_1 _20436_ (.CLK(net4698),
    .RESET_B(net4018),
    .D(_01752_),
    .Q_N(_09311_),
    .Q(\spiking_network_top_uut.all_data_out[151] ));
 sg13g2_dfrbp_1 _20437_ (.CLK(net4711),
    .RESET_B(net4031),
    .D(_01753_),
    .Q_N(_09310_),
    .Q(\spiking_network_top_uut.all_data_out[824] ));
 sg13g2_dfrbp_1 _20438_ (.CLK(net4711),
    .RESET_B(net4031),
    .D(_01754_),
    .Q_N(_00359_),
    .Q(\spiking_network_top_uut.all_data_out[825] ));
 sg13g2_dfrbp_1 _20439_ (.CLK(net4711),
    .RESET_B(net4031),
    .D(_01755_),
    .Q_N(_00289_),
    .Q(\spiking_network_top_uut.all_data_out[826] ));
 sg13g2_dfrbp_1 _20440_ (.CLK(net4710),
    .RESET_B(net4030),
    .D(_01756_),
    .Q_N(_09309_),
    .Q(\spiking_network_top_uut.all_data_out[827] ));
 sg13g2_dfrbp_1 _20441_ (.CLK(net4718),
    .RESET_B(net4037),
    .D(_01757_),
    .Q_N(_09308_),
    .Q(\spiking_network_top_uut.all_data_out[828] ));
 sg13g2_dfrbp_1 _20442_ (.CLK(net4715),
    .RESET_B(net4035),
    .D(_01758_),
    .Q_N(_00219_),
    .Q(\spiking_network_top_uut.all_data_out[829] ));
 sg13g2_dfrbp_1 _20443_ (.CLK(net4718),
    .RESET_B(net4037),
    .D(_01759_),
    .Q_N(_00149_),
    .Q(\spiking_network_top_uut.all_data_out[830] ));
 sg13g2_dfrbp_1 _20444_ (.CLK(net4713),
    .RESET_B(net4033),
    .D(_01760_),
    .Q_N(_09307_),
    .Q(\spiking_network_top_uut.all_data_out[831] ));
 sg13g2_dfrbp_1 _20445_ (.CLK(net4733),
    .RESET_B(net4053),
    .D(_01761_),
    .Q_N(_09306_),
    .Q(\spiking_network_top_uut.all_data_out[136] ));
 sg13g2_dfrbp_1 _20446_ (.CLK(net4732),
    .RESET_B(net4054),
    .D(_01762_),
    .Q_N(_09305_),
    .Q(\spiking_network_top_uut.all_data_out[137] ));
 sg13g2_dfrbp_1 _20447_ (.CLK(net4751),
    .RESET_B(net4072),
    .D(_01763_),
    .Q_N(_09304_),
    .Q(\spiking_network_top_uut.all_data_out[138] ));
 sg13g2_dfrbp_1 _20448_ (.CLK(net4732),
    .RESET_B(net4052),
    .D(_01764_),
    .Q_N(_09303_),
    .Q(\spiking_network_top_uut.all_data_out[139] ));
 sg13g2_dfrbp_1 _20449_ (.CLK(net4732),
    .RESET_B(net4052),
    .D(_01765_),
    .Q_N(_09302_),
    .Q(\spiking_network_top_uut.all_data_out[140] ));
 sg13g2_dfrbp_1 _20450_ (.CLK(net4751),
    .RESET_B(net4072),
    .D(_01766_),
    .Q_N(_09301_),
    .Q(\spiking_network_top_uut.all_data_out[141] ));
 sg13g2_dfrbp_1 _20451_ (.CLK(net4733),
    .RESET_B(net4053),
    .D(_01767_),
    .Q_N(_09300_),
    .Q(\spiking_network_top_uut.all_data_out[142] ));
 sg13g2_dfrbp_1 _20452_ (.CLK(net4734),
    .RESET_B(net4054),
    .D(_01768_),
    .Q_N(_09299_),
    .Q(\spiking_network_top_uut.all_data_out[143] ));
 sg13g2_dfrbp_1 _20453_ (.CLK(net4805),
    .RESET_B(net4127),
    .D(_01769_),
    .Q_N(_09298_),
    .Q(\spiking_network_top_uut.all_data_out[480] ));
 sg13g2_dfrbp_1 _20454_ (.CLK(net4806),
    .RESET_B(net4128),
    .D(_01770_),
    .Q_N(_00402_),
    .Q(\spiking_network_top_uut.all_data_out[481] ));
 sg13g2_dfrbp_1 _20455_ (.CLK(net4806),
    .RESET_B(net4128),
    .D(_01771_),
    .Q_N(_00332_),
    .Q(\spiking_network_top_uut.all_data_out[482] ));
 sg13g2_dfrbp_1 _20456_ (.CLK(net4736),
    .RESET_B(net4057),
    .D(_01772_),
    .Q_N(_09297_),
    .Q(\spiking_network_top_uut.all_data_out[483] ));
 sg13g2_dfrbp_1 _20457_ (.CLK(net4803),
    .RESET_B(net4125),
    .D(_01773_),
    .Q_N(_09296_),
    .Q(\spiking_network_top_uut.all_data_out[484] ));
 sg13g2_dfrbp_1 _20458_ (.CLK(net4803),
    .RESET_B(net4125),
    .D(_01774_),
    .Q_N(_00262_),
    .Q(\spiking_network_top_uut.all_data_out[485] ));
 sg13g2_dfrbp_1 _20459_ (.CLK(net4803),
    .RESET_B(net4125),
    .D(_01775_),
    .Q_N(_00192_),
    .Q(\spiking_network_top_uut.all_data_out[486] ));
 sg13g2_dfrbp_1 _20460_ (.CLK(net4733),
    .RESET_B(net4053),
    .D(_01776_),
    .Q_N(_09295_),
    .Q(\spiking_network_top_uut.all_data_out[487] ));
 sg13g2_dfrbp_1 _20461_ (.CLK(net4732),
    .RESET_B(net4052),
    .D(_01777_),
    .Q_N(_09294_),
    .Q(\spiking_network_top_uut.all_data_out[128] ));
 sg13g2_dfrbp_1 _20462_ (.CLK(net4732),
    .RESET_B(net4052),
    .D(_01778_),
    .Q_N(_09293_),
    .Q(\spiking_network_top_uut.all_data_out[129] ));
 sg13g2_dfrbp_1 _20463_ (.CLK(net4751),
    .RESET_B(net4072),
    .D(_01779_),
    .Q_N(_09292_),
    .Q(\spiking_network_top_uut.all_data_out[130] ));
 sg13g2_dfrbp_1 _20464_ (.CLK(net4732),
    .RESET_B(net4052),
    .D(_01780_),
    .Q_N(_09291_),
    .Q(\spiking_network_top_uut.all_data_out[131] ));
 sg13g2_dfrbp_1 _20465_ (.CLK(net4733),
    .RESET_B(net4054),
    .D(_01781_),
    .Q_N(_09290_),
    .Q(\spiking_network_top_uut.all_data_out[132] ));
 sg13g2_dfrbp_1 _20466_ (.CLK(net4750),
    .RESET_B(net4071),
    .D(_01782_),
    .Q_N(_09289_),
    .Q(\spiking_network_top_uut.all_data_out[133] ));
 sg13g2_dfrbp_1 _20467_ (.CLK(net4733),
    .RESET_B(net4053),
    .D(_01783_),
    .Q_N(_09288_),
    .Q(\spiking_network_top_uut.all_data_out[134] ));
 sg13g2_dfrbp_1 _20468_ (.CLK(net4733),
    .RESET_B(net4053),
    .D(_01784_),
    .Q_N(_09287_),
    .Q(\spiking_network_top_uut.all_data_out[135] ));
 sg13g2_dfrbp_1 _20469_ (.CLK(net4660),
    .RESET_B(net3980),
    .D(_01785_),
    .Q_N(_09286_),
    .Q(\spiking_network_top_uut.all_data_out[832] ));
 sg13g2_dfrbp_1 _20470_ (.CLK(net4660),
    .RESET_B(net3980),
    .D(_01786_),
    .Q_N(_00358_),
    .Q(\spiking_network_top_uut.all_data_out[833] ));
 sg13g2_dfrbp_1 _20471_ (.CLK(net4660),
    .RESET_B(net3980),
    .D(_01787_),
    .Q_N(_00288_),
    .Q(\spiking_network_top_uut.all_data_out[834] ));
 sg13g2_dfrbp_1 _20472_ (.CLK(net4654),
    .RESET_B(net3973),
    .D(_01788_),
    .Q_N(_09285_),
    .Q(\spiking_network_top_uut.all_data_out[835] ));
 sg13g2_dfrbp_1 _20473_ (.CLK(net4650),
    .RESET_B(net3969),
    .D(_01789_),
    .Q_N(_09284_),
    .Q(\spiking_network_top_uut.all_data_out[836] ));
 sg13g2_dfrbp_1 _20474_ (.CLK(net4654),
    .RESET_B(net3973),
    .D(_01790_),
    .Q_N(_00218_),
    .Q(\spiking_network_top_uut.all_data_out[837] ));
 sg13g2_dfrbp_1 _20475_ (.CLK(net4654),
    .RESET_B(net3973),
    .D(_01791_),
    .Q_N(_00148_),
    .Q(\spiking_network_top_uut.all_data_out[838] ));
 sg13g2_dfrbp_1 _20476_ (.CLK(net4657),
    .RESET_B(net3976),
    .D(_01792_),
    .Q_N(_09283_),
    .Q(\spiking_network_top_uut.all_data_out[839] ));
 sg13g2_dfrbp_1 _20477_ (.CLK(net4729),
    .RESET_B(net4049),
    .D(_01793_),
    .Q_N(_09282_),
    .Q(\spiking_network_top_uut.all_data_out[120] ));
 sg13g2_dfrbp_1 _20478_ (.CLK(net4735),
    .RESET_B(net4055),
    .D(_01794_),
    .Q_N(_09281_),
    .Q(\spiking_network_top_uut.all_data_out[121] ));
 sg13g2_dfrbp_1 _20479_ (.CLK(net4729),
    .RESET_B(net4049),
    .D(_01795_),
    .Q_N(_09280_),
    .Q(\spiking_network_top_uut.all_data_out[122] ));
 sg13g2_dfrbp_1 _20480_ (.CLK(net4735),
    .RESET_B(net4055),
    .D(_01796_),
    .Q_N(_09279_),
    .Q(\spiking_network_top_uut.all_data_out[123] ));
 sg13g2_dfrbp_1 _20481_ (.CLK(net4734),
    .RESET_B(net4057),
    .D(_01797_),
    .Q_N(_09278_),
    .Q(\spiking_network_top_uut.all_data_out[124] ));
 sg13g2_dfrbp_1 _20482_ (.CLK(net4725),
    .RESET_B(net4045),
    .D(_01798_),
    .Q_N(_09277_),
    .Q(\spiking_network_top_uut.all_data_out[125] ));
 sg13g2_dfrbp_1 _20483_ (.CLK(net4733),
    .RESET_B(net4057),
    .D(_01799_),
    .Q_N(_09276_),
    .Q(\spiking_network_top_uut.all_data_out[126] ));
 sg13g2_dfrbp_1 _20484_ (.CLK(net4725),
    .RESET_B(net4045),
    .D(_01800_),
    .Q_N(_09275_),
    .Q(\spiking_network_top_uut.all_data_out[127] ));
 sg13g2_dfrbp_1 _20485_ (.CLK(net4744),
    .RESET_B(net4067),
    .D(_01801_),
    .Q_N(_09274_),
    .Q(\spiking_network_top_uut.all_data_out[656] ));
 sg13g2_dfrbp_1 _20486_ (.CLK(net4745),
    .RESET_B(net4066),
    .D(_01802_),
    .Q_N(_00380_),
    .Q(\spiking_network_top_uut.all_data_out[657] ));
 sg13g2_dfrbp_1 _20487_ (.CLK(net4744),
    .RESET_B(net4065),
    .D(_01803_),
    .Q_N(_00310_),
    .Q(\spiking_network_top_uut.all_data_out[658] ));
 sg13g2_dfrbp_1 _20488_ (.CLK(net4757),
    .RESET_B(net4078),
    .D(_01804_),
    .Q_N(_09273_),
    .Q(\spiking_network_top_uut.all_data_out[659] ));
 sg13g2_dfrbp_1 _20489_ (.CLK(net4767),
    .RESET_B(net4088),
    .D(_01805_),
    .Q_N(_09272_),
    .Q(\spiking_network_top_uut.all_data_out[660] ));
 sg13g2_dfrbp_1 _20490_ (.CLK(net4767),
    .RESET_B(net4088),
    .D(_01806_),
    .Q_N(_00240_),
    .Q(\spiking_network_top_uut.all_data_out[661] ));
 sg13g2_dfrbp_1 _20491_ (.CLK(net4768),
    .RESET_B(net4089),
    .D(_01807_),
    .Q_N(_00170_),
    .Q(\spiking_network_top_uut.all_data_out[662] ));
 sg13g2_dfrbp_1 _20492_ (.CLK(net4757),
    .RESET_B(net4078),
    .D(_01808_),
    .Q_N(_09271_),
    .Q(\spiking_network_top_uut.all_data_out[663] ));
 sg13g2_dfrbp_1 _20493_ (.CLK(net4729),
    .RESET_B(net4049),
    .D(_01809_),
    .Q_N(_09270_),
    .Q(\spiking_network_top_uut.all_data_out[112] ));
 sg13g2_dfrbp_1 _20494_ (.CLK(net4725),
    .RESET_B(net4045),
    .D(_01810_),
    .Q_N(_09269_),
    .Q(\spiking_network_top_uut.all_data_out[113] ));
 sg13g2_dfrbp_1 _20495_ (.CLK(net4725),
    .RESET_B(net4045),
    .D(_01811_),
    .Q_N(_09268_),
    .Q(\spiking_network_top_uut.all_data_out[114] ));
 sg13g2_dfrbp_1 _20496_ (.CLK(net4726),
    .RESET_B(net4046),
    .D(_01812_),
    .Q_N(_09267_),
    .Q(\spiking_network_top_uut.all_data_out[115] ));
 sg13g2_dfrbp_1 _20497_ (.CLK(net4734),
    .RESET_B(net4052),
    .D(_01813_),
    .Q_N(_09266_),
    .Q(\spiking_network_top_uut.all_data_out[116] ));
 sg13g2_dfrbp_1 _20498_ (.CLK(net4734),
    .RESET_B(net4054),
    .D(_01814_),
    .Q_N(_09265_),
    .Q(\spiking_network_top_uut.all_data_out[117] ));
 sg13g2_dfrbp_1 _20499_ (.CLK(net4734),
    .RESET_B(net4054),
    .D(_01815_),
    .Q_N(_09264_),
    .Q(\spiking_network_top_uut.all_data_out[118] ));
 sg13g2_dfrbp_1 _20500_ (.CLK(net4732),
    .RESET_B(net4055),
    .D(_01816_),
    .Q_N(_09263_),
    .Q(\spiking_network_top_uut.all_data_out[119] ));
 sg13g2_dfrbp_1 _20501_ (.CLK(net4655),
    .RESET_B(net3974),
    .D(_01817_),
    .Q_N(_09262_),
    .Q(\spiking_network_top_uut.all_data_out[840] ));
 sg13g2_dfrbp_1 _20502_ (.CLK(net4654),
    .RESET_B(net3973),
    .D(_01818_),
    .Q_N(_00357_),
    .Q(\spiking_network_top_uut.all_data_out[841] ));
 sg13g2_dfrbp_1 _20503_ (.CLK(net4654),
    .RESET_B(net3973),
    .D(_01819_),
    .Q_N(_00287_),
    .Q(\spiking_network_top_uut.all_data_out[842] ));
 sg13g2_dfrbp_1 _20504_ (.CLK(net4649),
    .RESET_B(net3968),
    .D(_01820_),
    .Q_N(_09261_),
    .Q(\spiking_network_top_uut.all_data_out[843] ));
 sg13g2_dfrbp_1 _20505_ (.CLK(net4649),
    .RESET_B(net3968),
    .D(_01821_),
    .Q_N(_09260_),
    .Q(\spiking_network_top_uut.all_data_out[844] ));
 sg13g2_dfrbp_1 _20506_ (.CLK(net4654),
    .RESET_B(net3973),
    .D(_01822_),
    .Q_N(_00217_),
    .Q(\spiking_network_top_uut.all_data_out[845] ));
 sg13g2_dfrbp_1 _20507_ (.CLK(net4648),
    .RESET_B(net3979),
    .D(_01823_),
    .Q_N(_00147_),
    .Q(\spiking_network_top_uut.all_data_out[846] ));
 sg13g2_dfrbp_1 _20508_ (.CLK(net4649),
    .RESET_B(net3968),
    .D(_01824_),
    .Q_N(_09259_),
    .Q(\spiking_network_top_uut.all_data_out[847] ));
 sg13g2_dfrbp_1 _20509_ (.CLK(net4736),
    .RESET_B(net4057),
    .D(_01825_),
    .Q_N(_09258_),
    .Q(\spiking_network_top_uut.all_data_out[104] ));
 sg13g2_dfrbp_1 _20510_ (.CLK(net4737),
    .RESET_B(net4056),
    .D(_01826_),
    .Q_N(_09257_),
    .Q(\spiking_network_top_uut.all_data_out[105] ));
 sg13g2_dfrbp_1 _20511_ (.CLK(net4737),
    .RESET_B(net4056),
    .D(_01827_),
    .Q_N(_09256_),
    .Q(\spiking_network_top_uut.all_data_out[106] ));
 sg13g2_dfrbp_1 _20512_ (.CLK(net4737),
    .RESET_B(net4056),
    .D(_01828_),
    .Q_N(_09255_),
    .Q(\spiking_network_top_uut.all_data_out[107] ));
 sg13g2_dfrbp_1 _20513_ (.CLK(net4736),
    .RESET_B(net4058),
    .D(_01829_),
    .Q_N(_09254_),
    .Q(\spiking_network_top_uut.all_data_out[108] ));
 sg13g2_dfrbp_1 _20514_ (.CLK(net4735),
    .RESET_B(net4056),
    .D(_01830_),
    .Q_N(_09253_),
    .Q(\spiking_network_top_uut.all_data_out[109] ));
 sg13g2_dfrbp_1 _20515_ (.CLK(net4736),
    .RESET_B(net4057),
    .D(_01831_),
    .Q_N(_09252_),
    .Q(\spiking_network_top_uut.all_data_out[110] ));
 sg13g2_dfrbp_1 _20516_ (.CLK(net4736),
    .RESET_B(net4058),
    .D(_01832_),
    .Q_N(_09251_),
    .Q(\spiking_network_top_uut.all_data_out[111] ));
 sg13g2_dfrbp_1 _20517_ (.CLK(net4811),
    .RESET_B(net4134),
    .D(_01833_),
    .Q_N(_09250_),
    .Q(\spiking_network_top_uut.all_data_out[472] ));
 sg13g2_dfrbp_1 _20518_ (.CLK(net4807),
    .RESET_B(net4132),
    .D(_01834_),
    .Q_N(_00403_),
    .Q(\spiking_network_top_uut.all_data_out[473] ));
 sg13g2_dfrbp_1 _20519_ (.CLK(net4811),
    .RESET_B(net4133),
    .D(_01835_),
    .Q_N(_00333_),
    .Q(\spiking_network_top_uut.all_data_out[474] ));
 sg13g2_dfrbp_1 _20520_ (.CLK(net4785),
    .RESET_B(net4107),
    .D(_01836_),
    .Q_N(_09249_),
    .Q(\spiking_network_top_uut.all_data_out[475] ));
 sg13g2_dfrbp_1 _20521_ (.CLK(net4808),
    .RESET_B(net4129),
    .D(_01837_),
    .Q_N(_09248_),
    .Q(\spiking_network_top_uut.all_data_out[476] ));
 sg13g2_dfrbp_1 _20522_ (.CLK(net4808),
    .RESET_B(net4129),
    .D(_01838_),
    .Q_N(_00263_),
    .Q(\spiking_network_top_uut.all_data_out[477] ));
 sg13g2_dfrbp_1 _20523_ (.CLK(net4808),
    .RESET_B(net4129),
    .D(_01839_),
    .Q_N(_00193_),
    .Q(\spiking_network_top_uut.all_data_out[478] ));
 sg13g2_dfrbp_1 _20524_ (.CLK(net4802),
    .RESET_B(net4124),
    .D(_01840_),
    .Q_N(_09247_),
    .Q(\spiking_network_top_uut.all_data_out[479] ));
 sg13g2_dfrbp_1 _20525_ (.CLK(net4737),
    .RESET_B(net4058),
    .D(_01841_),
    .Q_N(_09246_),
    .Q(\spiking_network_top_uut.all_data_out[96] ));
 sg13g2_dfrbp_1 _20526_ (.CLK(net4736),
    .RESET_B(net4057),
    .D(_01842_),
    .Q_N(_09245_),
    .Q(\spiking_network_top_uut.all_data_out[97] ));
 sg13g2_dfrbp_1 _20527_ (.CLK(net4729),
    .RESET_B(net4049),
    .D(_01843_),
    .Q_N(_09244_),
    .Q(\spiking_network_top_uut.all_data_out[98] ));
 sg13g2_dfrbp_1 _20528_ (.CLK(net4735),
    .RESET_B(net4055),
    .D(_01844_),
    .Q_N(_09243_),
    .Q(\spiking_network_top_uut.all_data_out[99] ));
 sg13g2_dfrbp_1 _20529_ (.CLK(net4735),
    .RESET_B(net4055),
    .D(_01845_),
    .Q_N(_09242_),
    .Q(\spiking_network_top_uut.all_data_out[100] ));
 sg13g2_dfrbp_1 _20530_ (.CLK(net4735),
    .RESET_B(net4055),
    .D(_01846_),
    .Q_N(_09241_),
    .Q(\spiking_network_top_uut.all_data_out[101] ));
 sg13g2_dfrbp_1 _20531_ (.CLK(net4735),
    .RESET_B(net4055),
    .D(_01847_),
    .Q_N(_09240_),
    .Q(\spiking_network_top_uut.all_data_out[102] ));
 sg13g2_dfrbp_1 _20532_ (.CLK(net4735),
    .RESET_B(net4055),
    .D(_01848_),
    .Q_N(_09239_),
    .Q(\spiking_network_top_uut.all_data_out[103] ));
 sg13g2_dfrbp_1 _20533_ (.CLK(net4667),
    .RESET_B(net3987),
    .D(_01849_),
    .Q_N(_09238_),
    .Q(\spiking_network_top_uut.all_data_out[848] ));
 sg13g2_dfrbp_1 _20534_ (.CLK(net4670),
    .RESET_B(net3989),
    .D(_01850_),
    .Q_N(_00356_),
    .Q(\spiking_network_top_uut.all_data_out[849] ));
 sg13g2_dfrbp_1 _20535_ (.CLK(net4679),
    .RESET_B(net3998),
    .D(_01851_),
    .Q_N(_00286_),
    .Q(\spiking_network_top_uut.all_data_out[850] ));
 sg13g2_dfrbp_1 _20536_ (.CLK(net4667),
    .RESET_B(net3987),
    .D(_01852_),
    .Q_N(_09237_),
    .Q(\spiking_network_top_uut.all_data_out[851] ));
 sg13g2_dfrbp_1 _20537_ (.CLK(net4665),
    .RESET_B(net3985),
    .D(_01853_),
    .Q_N(_09236_),
    .Q(\spiking_network_top_uut.all_data_out[852] ));
 sg13g2_dfrbp_1 _20538_ (.CLK(net4660),
    .RESET_B(net3980),
    .D(_01854_),
    .Q_N(_00216_),
    .Q(\spiking_network_top_uut.all_data_out[853] ));
 sg13g2_dfrbp_1 _20539_ (.CLK(net4679),
    .RESET_B(net3998),
    .D(_01855_),
    .Q_N(_00146_),
    .Q(\spiking_network_top_uut.all_data_out[854] ));
 sg13g2_dfrbp_1 _20540_ (.CLK(net4668),
    .RESET_B(net3988),
    .D(_01856_),
    .Q_N(_09235_),
    .Q(\spiking_network_top_uut.all_data_out[855] ));
 sg13g2_dfrbp_1 _20541_ (.CLK(net4696),
    .RESET_B(net4015),
    .D(_01857_),
    .Q_N(_09234_),
    .Q(\spiking_network_top_uut.all_data_out[88] ));
 sg13g2_dfrbp_1 _20542_ (.CLK(net4696),
    .RESET_B(net4015),
    .D(_01858_),
    .Q_N(_09233_),
    .Q(\spiking_network_top_uut.all_data_out[89] ));
 sg13g2_dfrbp_1 _20543_ (.CLK(net4697),
    .RESET_B(net4016),
    .D(_01859_),
    .Q_N(_09232_),
    .Q(\spiking_network_top_uut.all_data_out[90] ));
 sg13g2_dfrbp_1 _20544_ (.CLK(net4696),
    .RESET_B(net4015),
    .D(_01860_),
    .Q_N(_09231_),
    .Q(\spiking_network_top_uut.all_data_out[91] ));
 sg13g2_dfrbp_1 _20545_ (.CLK(net4695),
    .RESET_B(net4014),
    .D(_01861_),
    .Q_N(_09230_),
    .Q(\spiking_network_top_uut.all_data_out[92] ));
 sg13g2_dfrbp_1 _20546_ (.CLK(net4697),
    .RESET_B(net4016),
    .D(_01862_),
    .Q_N(_09229_),
    .Q(\spiking_network_top_uut.all_data_out[93] ));
 sg13g2_dfrbp_1 _20547_ (.CLK(net4697),
    .RESET_B(net4016),
    .D(_01863_),
    .Q_N(_09228_),
    .Q(\spiking_network_top_uut.all_data_out[94] ));
 sg13g2_dfrbp_1 _20548_ (.CLK(net4695),
    .RESET_B(net4014),
    .D(_01864_),
    .Q_N(_09227_),
    .Q(\spiking_network_top_uut.all_data_out[95] ));
 sg13g2_dfrbp_1 _20549_ (.CLK(net4685),
    .RESET_B(net4004),
    .D(_01865_),
    .Q_N(_09226_),
    .Q(\spiking_network_top_uut.all_data_out[600] ));
 sg13g2_dfrbp_1 _20550_ (.CLK(net4685),
    .RESET_B(net4004),
    .D(_01866_),
    .Q_N(_00387_),
    .Q(\spiking_network_top_uut.all_data_out[601] ));
 sg13g2_dfrbp_1 _20551_ (.CLK(net4685),
    .RESET_B(net4004),
    .D(_01867_),
    .Q_N(_00317_),
    .Q(\spiking_network_top_uut.all_data_out[602] ));
 sg13g2_dfrbp_1 _20552_ (.CLK(net4685),
    .RESET_B(net4004),
    .D(_01868_),
    .Q_N(_09225_),
    .Q(\spiking_network_top_uut.all_data_out[603] ));
 sg13g2_dfrbp_1 _20553_ (.CLK(net4715),
    .RESET_B(net4035),
    .D(_01869_),
    .Q_N(_09224_),
    .Q(\spiking_network_top_uut.all_data_out[604] ));
 sg13g2_dfrbp_1 _20554_ (.CLK(net4718),
    .RESET_B(net4037),
    .D(_01870_),
    .Q_N(_00247_),
    .Q(\spiking_network_top_uut.all_data_out[605] ));
 sg13g2_dfrbp_1 _20555_ (.CLK(net4718),
    .RESET_B(net4037),
    .D(_01871_),
    .Q_N(_00177_),
    .Q(\spiking_network_top_uut.all_data_out[606] ));
 sg13g2_dfrbp_1 _20556_ (.CLK(net4716),
    .RESET_B(net4036),
    .D(_01872_),
    .Q_N(_09223_),
    .Q(\spiking_network_top_uut.all_data_out[607] ));
 sg13g2_dfrbp_1 _20557_ (.CLK(net4676),
    .RESET_B(net3995),
    .D(_01873_),
    .Q_N(_09222_),
    .Q(\spiking_network_top_uut.all_data_out[80] ));
 sg13g2_dfrbp_1 _20558_ (.CLK(net4697),
    .RESET_B(net4016),
    .D(_01874_),
    .Q_N(_09221_),
    .Q(\spiking_network_top_uut.all_data_out[81] ));
 sg13g2_dfrbp_1 _20559_ (.CLK(net4695),
    .RESET_B(net4015),
    .D(_01875_),
    .Q_N(_09220_),
    .Q(\spiking_network_top_uut.all_data_out[82] ));
 sg13g2_dfrbp_1 _20560_ (.CLK(net4697),
    .RESET_B(net4016),
    .D(_01876_),
    .Q_N(_09219_),
    .Q(\spiking_network_top_uut.all_data_out[83] ));
 sg13g2_dfrbp_1 _20561_ (.CLK(net4695),
    .RESET_B(net4014),
    .D(_01877_),
    .Q_N(_09218_),
    .Q(\spiking_network_top_uut.all_data_out[84] ));
 sg13g2_dfrbp_1 _20562_ (.CLK(net4695),
    .RESET_B(net4014),
    .D(_01878_),
    .Q_N(_09217_),
    .Q(\spiking_network_top_uut.all_data_out[85] ));
 sg13g2_dfrbp_1 _20563_ (.CLK(net4697),
    .RESET_B(net4016),
    .D(_01879_),
    .Q_N(_09216_),
    .Q(\spiking_network_top_uut.all_data_out[86] ));
 sg13g2_dfrbp_1 _20564_ (.CLK(net4676),
    .RESET_B(net3995),
    .D(_01880_),
    .Q_N(_09215_),
    .Q(\spiking_network_top_uut.all_data_out[87] ));
 sg13g2_dfrbp_1 _20565_ (.CLK(net4678),
    .RESET_B(net3997),
    .D(_01881_),
    .Q_N(_09214_),
    .Q(\spiking_network_top_uut.all_data_out[856] ));
 sg13g2_dfrbp_1 _20566_ (.CLK(net4678),
    .RESET_B(net3997),
    .D(_01882_),
    .Q_N(_00355_),
    .Q(\spiking_network_top_uut.all_data_out[857] ));
 sg13g2_dfrbp_1 _20567_ (.CLK(net4678),
    .RESET_B(net3997),
    .D(_01883_),
    .Q_N(_00285_),
    .Q(\spiking_network_top_uut.all_data_out[858] ));
 sg13g2_dfrbp_1 _20568_ (.CLK(net4679),
    .RESET_B(net3998),
    .D(_01884_),
    .Q_N(_09213_),
    .Q(\spiking_network_top_uut.all_data_out[859] ));
 sg13g2_dfrbp_1 _20569_ (.CLK(net4678),
    .RESET_B(net3997),
    .D(_01885_),
    .Q_N(_09212_),
    .Q(\spiking_network_top_uut.all_data_out[860] ));
 sg13g2_dfrbp_1 _20570_ (.CLK(net4664),
    .RESET_B(net3984),
    .D(_01886_),
    .Q_N(_00215_),
    .Q(\spiking_network_top_uut.all_data_out[861] ));
 sg13g2_dfrbp_1 _20571_ (.CLK(net4664),
    .RESET_B(net3984),
    .D(_01887_),
    .Q_N(_00145_),
    .Q(\spiking_network_top_uut.all_data_out[862] ));
 sg13g2_dfrbp_1 _20572_ (.CLK(net4679),
    .RESET_B(net3998),
    .D(_01888_),
    .Q_N(_09211_),
    .Q(\spiking_network_top_uut.all_data_out[863] ));
 sg13g2_dfrbp_1 _20573_ (.CLK(net4701),
    .RESET_B(net4026),
    .D(_01889_),
    .Q_N(_09210_),
    .Q(\spiking_network_top_uut.all_data_out[72] ));
 sg13g2_dfrbp_1 _20574_ (.CLK(net4723),
    .RESET_B(net4043),
    .D(_01890_),
    .Q_N(_09209_),
    .Q(\spiking_network_top_uut.all_data_out[73] ));
 sg13g2_dfrbp_1 _20575_ (.CLK(net4701),
    .RESET_B(net4021),
    .D(_01891_),
    .Q_N(_09208_),
    .Q(\spiking_network_top_uut.all_data_out[74] ));
 sg13g2_dfrbp_1 _20576_ (.CLK(net4701),
    .RESET_B(net4021),
    .D(_01892_),
    .Q_N(_09207_),
    .Q(\spiking_network_top_uut.all_data_out[75] ));
 sg13g2_dfrbp_1 _20577_ (.CLK(net4723),
    .RESET_B(net4043),
    .D(_01893_),
    .Q_N(_09206_),
    .Q(\spiking_network_top_uut.all_data_out[76] ));
 sg13g2_dfrbp_1 _20578_ (.CLK(net4700),
    .RESET_B(net4021),
    .D(_01894_),
    .Q_N(_09205_),
    .Q(\spiking_network_top_uut.all_data_out[77] ));
 sg13g2_dfrbp_1 _20579_ (.CLK(net4700),
    .RESET_B(net4020),
    .D(_01895_),
    .Q_N(_09204_),
    .Q(\spiking_network_top_uut.all_data_out[78] ));
 sg13g2_dfrbp_1 _20580_ (.CLK(net4724),
    .RESET_B(net4043),
    .D(_01896_),
    .Q_N(_09203_),
    .Q(\spiking_network_top_uut.all_data_out[79] ));
 sg13g2_dfrbp_1 _20581_ (.CLK(net4781),
    .RESET_B(net4103),
    .D(_01897_),
    .Q_N(_09202_),
    .Q(\spiking_network_top_uut.all_data_out[464] ));
 sg13g2_dfrbp_1 _20582_ (.CLK(net4781),
    .RESET_B(net4103),
    .D(_01898_),
    .Q_N(_00404_),
    .Q(\spiking_network_top_uut.all_data_out[465] ));
 sg13g2_dfrbp_1 _20583_ (.CLK(net4781),
    .RESET_B(net4103),
    .D(_01899_),
    .Q_N(_00334_),
    .Q(\spiking_network_top_uut.all_data_out[466] ));
 sg13g2_dfrbp_1 _20584_ (.CLK(net4782),
    .RESET_B(net4104),
    .D(_01900_),
    .Q_N(_09201_),
    .Q(\spiking_network_top_uut.all_data_out[467] ));
 sg13g2_dfrbp_1 _20585_ (.CLK(net4753),
    .RESET_B(net4074),
    .D(_01901_),
    .Q_N(_09200_),
    .Q(\spiking_network_top_uut.all_data_out[468] ));
 sg13g2_dfrbp_1 _20586_ (.CLK(net4761),
    .RESET_B(net4082),
    .D(_01902_),
    .Q_N(_00264_),
    .Q(\spiking_network_top_uut.all_data_out[469] ));
 sg13g2_dfrbp_1 _20587_ (.CLK(net4754),
    .RESET_B(net4074),
    .D(_01903_),
    .Q_N(_00194_),
    .Q(\spiking_network_top_uut.all_data_out[470] ));
 sg13g2_dfrbp_1 _20588_ (.CLK(net4736),
    .RESET_B(net4057),
    .D(_01904_),
    .Q_N(_09199_),
    .Q(\spiking_network_top_uut.all_data_out[471] ));
 sg13g2_dfrbp_1 _20589_ (.CLK(net4723),
    .RESET_B(net4046),
    .D(_01905_),
    .Q_N(_09198_),
    .Q(\spiking_network_top_uut.all_data_out[64] ));
 sg13g2_dfrbp_1 _20590_ (.CLK(net4723),
    .RESET_B(net4043),
    .D(_01906_),
    .Q_N(_09197_),
    .Q(\spiking_network_top_uut.all_data_out[65] ));
 sg13g2_dfrbp_1 _20591_ (.CLK(net4727),
    .RESET_B(net4047),
    .D(_01907_),
    .Q_N(_09196_),
    .Q(\spiking_network_top_uut.all_data_out[66] ));
 sg13g2_dfrbp_1 _20592_ (.CLK(net4706),
    .RESET_B(net4026),
    .D(_01908_),
    .Q_N(_09195_),
    .Q(\spiking_network_top_uut.all_data_out[67] ));
 sg13g2_dfrbp_1 _20593_ (.CLK(net4723),
    .RESET_B(net4043),
    .D(_01909_),
    .Q_N(_09194_),
    .Q(\spiking_network_top_uut.all_data_out[68] ));
 sg13g2_dfrbp_1 _20594_ (.CLK(net4701),
    .RESET_B(net4021),
    .D(_01910_),
    .Q_N(_09193_),
    .Q(\spiking_network_top_uut.all_data_out[69] ));
 sg13g2_dfrbp_1 _20595_ (.CLK(net4701),
    .RESET_B(net4021),
    .D(_01911_),
    .Q_N(_09192_),
    .Q(\spiking_network_top_uut.all_data_out[70] ));
 sg13g2_dfrbp_1 _20596_ (.CLK(net4723),
    .RESET_B(net4043),
    .D(_01912_),
    .Q_N(_09191_),
    .Q(\spiking_network_top_uut.all_data_out[71] ));
 sg13g2_dfrbp_1 _20597_ (.CLK(net4660),
    .RESET_B(net3980),
    .D(_01913_),
    .Q_N(_09190_),
    .Q(\spiking_network_top_uut.all_data_out[864] ));
 sg13g2_dfrbp_1 _20598_ (.CLK(net4660),
    .RESET_B(net3980),
    .D(_01914_),
    .Q_N(_00354_),
    .Q(\spiking_network_top_uut.all_data_out[865] ));
 sg13g2_dfrbp_1 _20599_ (.CLK(net4660),
    .RESET_B(net3980),
    .D(_01915_),
    .Q_N(_00284_),
    .Q(\spiking_network_top_uut.all_data_out[866] ));
 sg13g2_dfrbp_1 _20600_ (.CLK(net4649),
    .RESET_B(net3968),
    .D(_01916_),
    .Q_N(_09189_),
    .Q(\spiking_network_top_uut.all_data_out[867] ));
 sg13g2_dfrbp_1 _20601_ (.CLK(net4650),
    .RESET_B(net3969),
    .D(_01917_),
    .Q_N(_09188_),
    .Q(\spiking_network_top_uut.all_data_out[868] ));
 sg13g2_dfrbp_1 _20602_ (.CLK(net4654),
    .RESET_B(net3973),
    .D(_01918_),
    .Q_N(_00214_),
    .Q(\spiking_network_top_uut.all_data_out[869] ));
 sg13g2_dfrbp_1 _20603_ (.CLK(net4655),
    .RESET_B(net3974),
    .D(_01919_),
    .Q_N(_00144_),
    .Q(\spiking_network_top_uut.all_data_out[870] ));
 sg13g2_dfrbp_1 _20604_ (.CLK(net4649),
    .RESET_B(net3968),
    .D(_01920_),
    .Q_N(_09187_),
    .Q(\spiking_network_top_uut.all_data_out[871] ));
 sg13g2_dfrbp_1 _20605_ (.CLK(net4727),
    .RESET_B(net4047),
    .D(_01921_),
    .Q_N(_09186_),
    .Q(\spiking_network_top_uut.all_data_out[56] ));
 sg13g2_dfrbp_1 _20606_ (.CLK(net4729),
    .RESET_B(net4049),
    .D(_01922_),
    .Q_N(_09185_),
    .Q(\spiking_network_top_uut.all_data_out[57] ));
 sg13g2_dfrbp_1 _20607_ (.CLK(net4730),
    .RESET_B(net4050),
    .D(_01923_),
    .Q_N(_09184_),
    .Q(\spiking_network_top_uut.all_data_out[58] ));
 sg13g2_dfrbp_1 _20608_ (.CLK(net4730),
    .RESET_B(net4050),
    .D(_01924_),
    .Q_N(_09183_),
    .Q(\spiking_network_top_uut.all_data_out[59] ));
 sg13g2_dfrbp_1 _20609_ (.CLK(net4730),
    .RESET_B(net4050),
    .D(_01925_),
    .Q_N(_09182_),
    .Q(\spiking_network_top_uut.all_data_out[60] ));
 sg13g2_dfrbp_1 _20610_ (.CLK(net4727),
    .RESET_B(net4047),
    .D(_01926_),
    .Q_N(_09181_),
    .Q(\spiking_network_top_uut.all_data_out[61] ));
 sg13g2_dfrbp_1 _20611_ (.CLK(net4730),
    .RESET_B(net4050),
    .D(_01927_),
    .Q_N(_09180_),
    .Q(\spiking_network_top_uut.all_data_out[62] ));
 sg13g2_dfrbp_1 _20612_ (.CLK(net4730),
    .RESET_B(net4050),
    .D(_01928_),
    .Q_N(_09179_),
    .Q(\spiking_network_top_uut.all_data_out[63] ));
 sg13g2_dfrbp_1 _20613_ (.CLK(net4711),
    .RESET_B(net4031),
    .D(_01929_),
    .Q_N(_09178_),
    .Q(\spiking_network_top_uut.all_data_out[664] ));
 sg13g2_dfrbp_1 _20614_ (.CLK(net4711),
    .RESET_B(net4031),
    .D(_01930_),
    .Q_N(_00379_),
    .Q(\spiking_network_top_uut.all_data_out[665] ));
 sg13g2_dfrbp_1 _20615_ (.CLK(net4716),
    .RESET_B(net4036),
    .D(_01931_),
    .Q_N(_00309_),
    .Q(\spiking_network_top_uut.all_data_out[666] ));
 sg13g2_dfrbp_1 _20616_ (.CLK(net4712),
    .RESET_B(net4032),
    .D(_01932_),
    .Q_N(_09177_),
    .Q(\spiking_network_top_uut.all_data_out[667] ));
 sg13g2_dfrbp_1 _20617_ (.CLK(net4718),
    .RESET_B(net4038),
    .D(_01933_),
    .Q_N(_09176_),
    .Q(\spiking_network_top_uut.all_data_out[668] ));
 sg13g2_dfrbp_1 _20618_ (.CLK(net4717),
    .RESET_B(net4040),
    .D(_01934_),
    .Q_N(_00239_),
    .Q(\spiking_network_top_uut.all_data_out[669] ));
 sg13g2_dfrbp_1 _20619_ (.CLK(net4717),
    .RESET_B(net4037),
    .D(_01935_),
    .Q_N(_00169_),
    .Q(\spiking_network_top_uut.all_data_out[670] ));
 sg13g2_dfrbp_1 _20620_ (.CLK(net4712),
    .RESET_B(net4032),
    .D(_01936_),
    .Q_N(_09175_),
    .Q(\spiking_network_top_uut.all_data_out[671] ));
 sg13g2_dfrbp_1 _20621_ (.CLK(net4727),
    .RESET_B(net4048),
    .D(_01937_),
    .Q_N(_09174_),
    .Q(\spiking_network_top_uut.all_data_out[48] ));
 sg13g2_dfrbp_1 _20622_ (.CLK(net4703),
    .RESET_B(net4023),
    .D(_01938_),
    .Q_N(_09173_),
    .Q(\spiking_network_top_uut.all_data_out[49] ));
 sg13g2_dfrbp_1 _20623_ (.CLK(net4728),
    .RESET_B(net4048),
    .D(_01939_),
    .Q_N(_09172_),
    .Q(\spiking_network_top_uut.all_data_out[50] ));
 sg13g2_dfrbp_1 _20624_ (.CLK(net4706),
    .RESET_B(net4026),
    .D(_01940_),
    .Q_N(_09171_),
    .Q(\spiking_network_top_uut.all_data_out[51] ));
 sg13g2_dfrbp_1 _20625_ (.CLK(net4703),
    .RESET_B(net4023),
    .D(_01941_),
    .Q_N(_09170_),
    .Q(\spiking_network_top_uut.all_data_out[52] ));
 sg13g2_dfrbp_1 _20626_ (.CLK(net4727),
    .RESET_B(net4047),
    .D(_01942_),
    .Q_N(_09169_),
    .Q(\spiking_network_top_uut.all_data_out[53] ));
 sg13g2_dfrbp_1 _20627_ (.CLK(net4727),
    .RESET_B(net4047),
    .D(_01943_),
    .Q_N(_09168_),
    .Q(\spiking_network_top_uut.all_data_out[54] ));
 sg13g2_dfrbp_1 _20628_ (.CLK(net4706),
    .RESET_B(net4026),
    .D(_01944_),
    .Q_N(_09167_),
    .Q(\spiking_network_top_uut.all_data_out[55] ));
 sg13g2_dfrbp_1 _20629_ (.CLK(net4649),
    .RESET_B(net3968),
    .D(_01945_),
    .Q_N(_09166_),
    .Q(\spiking_network_top_uut.all_data_out[872] ));
 sg13g2_dfrbp_1 _20630_ (.CLK(net4654),
    .RESET_B(net3973),
    .D(_01946_),
    .Q_N(_00353_),
    .Q(\spiking_network_top_uut.all_data_out[873] ));
 sg13g2_dfrbp_1 _20631_ (.CLK(net4655),
    .RESET_B(net3974),
    .D(_01947_),
    .Q_N(_00283_),
    .Q(\spiking_network_top_uut.all_data_out[874] ));
 sg13g2_dfrbp_1 _20632_ (.CLK(net4651),
    .RESET_B(net3970),
    .D(_01948_),
    .Q_N(_09165_),
    .Q(\spiking_network_top_uut.all_data_out[875] ));
 sg13g2_dfrbp_1 _20633_ (.CLK(net4649),
    .RESET_B(net3968),
    .D(_01949_),
    .Q_N(_09164_),
    .Q(\spiking_network_top_uut.all_data_out[876] ));
 sg13g2_dfrbp_1 _20634_ (.CLK(net4655),
    .RESET_B(net3974),
    .D(_01950_),
    .Q_N(_00213_),
    .Q(\spiking_network_top_uut.all_data_out[877] ));
 sg13g2_dfrbp_1 _20635_ (.CLK(net4648),
    .RESET_B(net3979),
    .D(_01951_),
    .Q_N(_00143_),
    .Q(\spiking_network_top_uut.all_data_out[878] ));
 sg13g2_dfrbp_1 _20636_ (.CLK(net4651),
    .RESET_B(net3970),
    .D(_01952_),
    .Q_N(_09163_),
    .Q(\spiking_network_top_uut.all_data_out[879] ));
 sg13g2_dfrbp_1 _20637_ (.CLK(net4756),
    .RESET_B(net4077),
    .D(_01953_),
    .Q_N(_09162_),
    .Q(\spiking_network_top_uut.all_data_out[40] ));
 sg13g2_dfrbp_1 _20638_ (.CLK(net4750),
    .RESET_B(net4071),
    .D(_01954_),
    .Q_N(_09161_),
    .Q(\spiking_network_top_uut.all_data_out[41] ));
 sg13g2_dfrbp_1 _20639_ (.CLK(net4753),
    .RESET_B(net4074),
    .D(_01955_),
    .Q_N(_09160_),
    .Q(\spiking_network_top_uut.all_data_out[42] ));
 sg13g2_dfrbp_1 _20640_ (.CLK(net4763),
    .RESET_B(net4084),
    .D(_01956_),
    .Q_N(_09159_),
    .Q(\spiking_network_top_uut.all_data_out[43] ));
 sg13g2_dfrbp_1 _20641_ (.CLK(net4756),
    .RESET_B(net4077),
    .D(_01957_),
    .Q_N(_09158_),
    .Q(\spiking_network_top_uut.all_data_out[44] ));
 sg13g2_dfrbp_1 _20642_ (.CLK(net4756),
    .RESET_B(net4077),
    .D(_01958_),
    .Q_N(_09157_),
    .Q(\spiking_network_top_uut.all_data_out[45] ));
 sg13g2_dfrbp_1 _20643_ (.CLK(net4755),
    .RESET_B(net4076),
    .D(_01959_),
    .Q_N(_09156_),
    .Q(\spiking_network_top_uut.all_data_out[46] ));
 sg13g2_dfrbp_1 _20644_ (.CLK(net4756),
    .RESET_B(net4077),
    .D(_01960_),
    .Q_N(_09155_),
    .Q(\spiking_network_top_uut.all_data_out[47] ));
 sg13g2_dfrbp_1 _20645_ (.CLK(net4795),
    .RESET_B(net4117),
    .D(_01961_),
    .Q_N(_09154_),
    .Q(\spiking_network_top_uut.all_data_out[456] ));
 sg13g2_dfrbp_1 _20646_ (.CLK(net4790),
    .RESET_B(net4111),
    .D(_01962_),
    .Q_N(_00405_),
    .Q(\spiking_network_top_uut.all_data_out[457] ));
 sg13g2_dfrbp_1 _20647_ (.CLK(net4790),
    .RESET_B(net4112),
    .D(_01963_),
    .Q_N(_00335_),
    .Q(\spiking_network_top_uut.all_data_out[458] ));
 sg13g2_dfrbp_1 _20648_ (.CLK(net4773),
    .RESET_B(net4094),
    .D(_01964_),
    .Q_N(_09153_),
    .Q(\spiking_network_top_uut.all_data_out[459] ));
 sg13g2_dfrbp_1 _20649_ (.CLK(net4795),
    .RESET_B(net4117),
    .D(_01965_),
    .Q_N(_09152_),
    .Q(\spiking_network_top_uut.all_data_out[460] ));
 sg13g2_dfrbp_1 _20650_ (.CLK(net4796),
    .RESET_B(net4123),
    .D(_01966_),
    .Q_N(_00265_),
    .Q(\spiking_network_top_uut.all_data_out[461] ));
 sg13g2_dfrbp_1 _20651_ (.CLK(net4799),
    .RESET_B(net4119),
    .D(_01967_),
    .Q_N(_00195_),
    .Q(\spiking_network_top_uut.all_data_out[462] ));
 sg13g2_dfrbp_1 _20652_ (.CLK(net4773),
    .RESET_B(net4094),
    .D(_01968_),
    .Q_N(_09151_),
    .Q(\spiking_network_top_uut.all_data_out[463] ));
 sg13g2_dfrbp_1 _20653_ (.CLK(net4758),
    .RESET_B(net4079),
    .D(_01969_),
    .Q_N(_09150_),
    .Q(\spiking_network_top_uut.all_data_out[32] ));
 sg13g2_dfrbp_1 _20654_ (.CLK(net4751),
    .RESET_B(net4072),
    .D(_01970_),
    .Q_N(_09149_),
    .Q(\spiking_network_top_uut.all_data_out[33] ));
 sg13g2_dfrbp_1 _20655_ (.CLK(net4751),
    .RESET_B(net4072),
    .D(_01971_),
    .Q_N(_09148_),
    .Q(\spiking_network_top_uut.all_data_out[34] ));
 sg13g2_dfrbp_1 _20656_ (.CLK(net4751),
    .RESET_B(net4072),
    .D(_01972_),
    .Q_N(_09147_),
    .Q(\spiking_network_top_uut.all_data_out[35] ));
 sg13g2_dfrbp_1 _20657_ (.CLK(net4757),
    .RESET_B(net4078),
    .D(_01973_),
    .Q_N(_09146_),
    .Q(\spiking_network_top_uut.all_data_out[36] ));
 sg13g2_dfrbp_1 _20658_ (.CLK(net4755),
    .RESET_B(net4076),
    .D(_01974_),
    .Q_N(_09145_),
    .Q(\spiking_network_top_uut.all_data_out[37] ));
 sg13g2_dfrbp_1 _20659_ (.CLK(net4758),
    .RESET_B(net4079),
    .D(_01975_),
    .Q_N(_09144_),
    .Q(\spiking_network_top_uut.all_data_out[38] ));
 sg13g2_dfrbp_1 _20660_ (.CLK(net4757),
    .RESET_B(net4078),
    .D(_01976_),
    .Q_N(_09143_),
    .Q(\spiking_network_top_uut.all_data_out[39] ));
 sg13g2_dfrbp_1 _20661_ (.CLK(net4667),
    .RESET_B(net3987),
    .D(_01977_),
    .Q_N(_09142_),
    .Q(\spiking_network_top_uut.all_data_out[880] ));
 sg13g2_dfrbp_1 _20662_ (.CLK(net4668),
    .RESET_B(net3988),
    .D(_01978_),
    .Q_N(_00352_),
    .Q(\spiking_network_top_uut.all_data_out[881] ));
 sg13g2_dfrbp_1 _20663_ (.CLK(net4667),
    .RESET_B(net3987),
    .D(_01979_),
    .Q_N(_00282_),
    .Q(\spiking_network_top_uut.all_data_out[882] ));
 sg13g2_dfrbp_1 _20664_ (.CLK(net4668),
    .RESET_B(net3988),
    .D(_01980_),
    .Q_N(_09141_),
    .Q(\spiking_network_top_uut.all_data_out[883] ));
 sg13g2_dfrbp_1 _20665_ (.CLK(net4660),
    .RESET_B(net3980),
    .D(_01981_),
    .Q_N(_09140_),
    .Q(\spiking_network_top_uut.all_data_out[884] ));
 sg13g2_dfrbp_1 _20666_ (.CLK(net4663),
    .RESET_B(net3983),
    .D(_01982_),
    .Q_N(_00212_),
    .Q(\spiking_network_top_uut.all_data_out[885] ));
 sg13g2_dfrbp_1 _20667_ (.CLK(net4663),
    .RESET_B(net3983),
    .D(_01983_),
    .Q_N(_00142_),
    .Q(\spiking_network_top_uut.all_data_out[886] ));
 sg13g2_dfrbp_1 _20668_ (.CLK(net4667),
    .RESET_B(net3987),
    .D(_01984_),
    .Q_N(_09139_),
    .Q(\spiking_network_top_uut.all_data_out[887] ));
 sg13g2_dfrbp_1 _20669_ (.CLK(net4678),
    .RESET_B(net3997),
    .D(_01985_),
    .Q_N(_09138_),
    .Q(\spiking_network_top_uut.all_data_out[24] ));
 sg13g2_dfrbp_1 _20670_ (.CLK(net4681),
    .RESET_B(net4000),
    .D(_01986_),
    .Q_N(_09137_),
    .Q(\spiking_network_top_uut.all_data_out[25] ));
 sg13g2_dfrbp_1 _20671_ (.CLK(net4681),
    .RESET_B(net4000),
    .D(_01987_),
    .Q_N(_09136_),
    .Q(\spiking_network_top_uut.all_data_out[26] ));
 sg13g2_dfrbp_1 _20672_ (.CLK(net4681),
    .RESET_B(net4000),
    .D(_01988_),
    .Q_N(_09135_),
    .Q(\spiking_network_top_uut.all_data_out[27] ));
 sg13g2_dfrbp_1 _20673_ (.CLK(net4669),
    .RESET_B(net3989),
    .D(_01989_),
    .Q_N(_09134_),
    .Q(\spiking_network_top_uut.all_data_out[28] ));
 sg13g2_dfrbp_1 _20674_ (.CLK(net4669),
    .RESET_B(net3988),
    .D(_01990_),
    .Q_N(_09133_),
    .Q(\spiking_network_top_uut.all_data_out[29] ));
 sg13g2_dfrbp_1 _20675_ (.CLK(net4681),
    .RESET_B(net4000),
    .D(_01991_),
    .Q_N(_09132_),
    .Q(\spiking_network_top_uut.all_data_out[30] ));
 sg13g2_dfrbp_1 _20676_ (.CLK(net4668),
    .RESET_B(net3988),
    .D(_01992_),
    .Q_N(_09131_),
    .Q(\spiking_network_top_uut.all_data_out[31] ));
 sg13g2_dfrbp_1 _20677_ (.CLK(net4782),
    .RESET_B(net4104),
    .D(_01993_),
    .Q_N(_09130_),
    .Q(\spiking_network_top_uut.all_data_out[560] ));
 sg13g2_dfrbp_1 _20678_ (.CLK(net4781),
    .RESET_B(net4103),
    .D(_01994_),
    .Q_N(_00392_),
    .Q(\spiking_network_top_uut.all_data_out[561] ));
 sg13g2_dfrbp_1 _20679_ (.CLK(net4781),
    .RESET_B(net4103),
    .D(_01995_),
    .Q_N(_00322_),
    .Q(\spiking_network_top_uut.all_data_out[562] ));
 sg13g2_dfrbp_1 _20680_ (.CLK(net4762),
    .RESET_B(net4083),
    .D(_01996_),
    .Q_N(_09129_),
    .Q(\spiking_network_top_uut.all_data_out[563] ));
 sg13g2_dfrbp_1 _20681_ (.CLK(net4761),
    .RESET_B(net4082),
    .D(_01997_),
    .Q_N(_09128_),
    .Q(\spiking_network_top_uut.all_data_out[564] ));
 sg13g2_dfrbp_1 _20682_ (.CLK(net4753),
    .RESET_B(net4074),
    .D(_01998_),
    .Q_N(_00252_),
    .Q(\spiking_network_top_uut.all_data_out[565] ));
 sg13g2_dfrbp_1 _20683_ (.CLK(net4760),
    .RESET_B(net4081),
    .D(_01999_),
    .Q_N(_00182_),
    .Q(\spiking_network_top_uut.all_data_out[566] ));
 sg13g2_dfrbp_1 _20684_ (.CLK(net4752),
    .RESET_B(net4073),
    .D(_02000_),
    .Q_N(_09127_),
    .Q(\spiking_network_top_uut.all_data_out[567] ));
 sg13g2_dfrbp_1 _20685_ (.CLK(net4657),
    .RESET_B(net3976),
    .D(_02001_),
    .Q_N(_09126_),
    .Q(\spiking_network_top_uut.all_data_out[16] ));
 sg13g2_dfrbp_1 _20686_ (.CLK(net4659),
    .RESET_B(net3978),
    .D(_02002_),
    .Q_N(_09125_),
    .Q(\spiking_network_top_uut.all_data_out[17] ));
 sg13g2_dfrbp_1 _20687_ (.CLK(net4659),
    .RESET_B(net3978),
    .D(_02003_),
    .Q_N(_09124_),
    .Q(\spiking_network_top_uut.all_data_out[18] ));
 sg13g2_dfrbp_1 _20688_ (.CLK(net4672),
    .RESET_B(net3991),
    .D(_02004_),
    .Q_N(_09123_),
    .Q(\spiking_network_top_uut.all_data_out[19] ));
 sg13g2_dfrbp_1 _20689_ (.CLK(net4659),
    .RESET_B(net3978),
    .D(_02005_),
    .Q_N(_09122_),
    .Q(\spiking_network_top_uut.all_data_out[20] ));
 sg13g2_dfrbp_1 _20690_ (.CLK(net4683),
    .RESET_B(net4002),
    .D(_02006_),
    .Q_N(_09121_),
    .Q(\spiking_network_top_uut.all_data_out[21] ));
 sg13g2_dfrbp_1 _20691_ (.CLK(net4750),
    .RESET_B(net4071),
    .D(_02007_),
    .Q_N(_09120_),
    .Q(\spiking_network_top_uut.all_data_out[22] ));
 sg13g2_dfrbp_1 _20692_ (.CLK(net4666),
    .RESET_B(net3986),
    .D(_02008_),
    .Q_N(_09119_),
    .Q(\spiking_network_top_uut.all_data_out[23] ));
 sg13g2_dfrbp_1 _20693_ (.CLK(net4678),
    .RESET_B(net3997),
    .D(_02009_),
    .Q_N(_09118_),
    .Q(\spiking_network_top_uut.all_data_out[888] ));
 sg13g2_dfrbp_1 _20694_ (.CLK(net4678),
    .RESET_B(net3997),
    .D(_02010_),
    .Q_N(_00351_),
    .Q(\spiking_network_top_uut.all_data_out[889] ));
 sg13g2_dfrbp_1 _20695_ (.CLK(net4680),
    .RESET_B(net3999),
    .D(_02011_),
    .Q_N(_00281_),
    .Q(\spiking_network_top_uut.all_data_out[890] ));
 sg13g2_dfrbp_1 _20696_ (.CLK(net4682),
    .RESET_B(net4001),
    .D(_02012_),
    .Q_N(_09117_),
    .Q(\spiking_network_top_uut.all_data_out[891] ));
 sg13g2_dfrbp_1 _20697_ (.CLK(net4664),
    .RESET_B(net3984),
    .D(_02013_),
    .Q_N(_09116_),
    .Q(\spiking_network_top_uut.all_data_out[892] ));
 sg13g2_dfrbp_1 _20698_ (.CLK(net4664),
    .RESET_B(net3984),
    .D(_02014_),
    .Q_N(_00211_),
    .Q(\spiking_network_top_uut.all_data_out[893] ));
 sg13g2_dfrbp_1 _20699_ (.CLK(net4664),
    .RESET_B(net3984),
    .D(_02015_),
    .Q_N(_00141_),
    .Q(\spiking_network_top_uut.all_data_out[894] ));
 sg13g2_dfrbp_1 _20700_ (.CLK(net4681),
    .RESET_B(net4000),
    .D(_02016_),
    .Q_N(_09115_),
    .Q(\spiking_network_top_uut.all_data_out[895] ));
 sg13g2_dfrbp_1 _20701_ (.CLK(net4670),
    .RESET_B(net3989),
    .D(_02017_),
    .Q_N(_09114_),
    .Q(\spiking_network_top_uut.all_data_out[8] ));
 sg13g2_dfrbp_1 _20702_ (.CLK(net4679),
    .RESET_B(net3998),
    .D(_02018_),
    .Q_N(_09113_),
    .Q(\spiking_network_top_uut.all_data_out[9] ));
 sg13g2_dfrbp_1 _20703_ (.CLK(net4679),
    .RESET_B(net3998),
    .D(_02019_),
    .Q_N(_09112_),
    .Q(\spiking_network_top_uut.all_data_out[10] ));
 sg13g2_dfrbp_1 _20704_ (.CLK(net4665),
    .RESET_B(net3985),
    .D(_02020_),
    .Q_N(_09111_),
    .Q(\spiking_network_top_uut.all_data_out[11] ));
 sg13g2_dfrbp_1 _20705_ (.CLK(net4670),
    .RESET_B(net3989),
    .D(_02021_),
    .Q_N(_09110_),
    .Q(\spiking_network_top_uut.all_data_out[12] ));
 sg13g2_dfrbp_1 _20706_ (.CLK(net4755),
    .RESET_B(net4076),
    .D(_02022_),
    .Q_N(_09109_),
    .Q(\spiking_network_top_uut.all_data_out[13] ));
 sg13g2_dfrbp_1 _20707_ (.CLK(net4698),
    .RESET_B(net4018),
    .D(_02023_),
    .Q_N(_09108_),
    .Q(\spiking_network_top_uut.all_data_out[14] ));
 sg13g2_dfrbp_1 _20708_ (.CLK(net4725),
    .RESET_B(net4045),
    .D(_02024_),
    .Q_N(_09107_),
    .Q(\spiking_network_top_uut.all_data_out[15] ));
 sg13g2_dfrbp_1 _20709_ (.CLK(net4785),
    .RESET_B(net4107),
    .D(_02025_),
    .Q_N(_09106_),
    .Q(\spiking_network_top_uut.all_data_out[448] ));
 sg13g2_dfrbp_1 _20710_ (.CLK(net4785),
    .RESET_B(net4108),
    .D(_02026_),
    .Q_N(_00406_),
    .Q(\spiking_network_top_uut.all_data_out[449] ));
 sg13g2_dfrbp_1 _20711_ (.CLK(net4786),
    .RESET_B(net4108),
    .D(_02027_),
    .Q_N(_00336_),
    .Q(\spiking_network_top_uut.all_data_out[450] ));
 sg13g2_dfrbp_1 _20712_ (.CLK(net4785),
    .RESET_B(net4107),
    .D(_02028_),
    .Q_N(_09105_),
    .Q(\spiking_network_top_uut.all_data_out[451] ));
 sg13g2_dfrbp_1 _20713_ (.CLK(net4783),
    .RESET_B(net4105),
    .D(_02029_),
    .Q_N(_09104_),
    .Q(\spiking_network_top_uut.all_data_out[452] ));
 sg13g2_dfrbp_1 _20714_ (.CLK(net4783),
    .RESET_B(net4105),
    .D(_02030_),
    .Q_N(_00266_),
    .Q(\spiking_network_top_uut.all_data_out[453] ));
 sg13g2_dfrbp_1 _20715_ (.CLK(net4783),
    .RESET_B(net4105),
    .D(_02031_),
    .Q_N(_00196_),
    .Q(\spiking_network_top_uut.all_data_out[454] ));
 sg13g2_dfrbp_1 _20716_ (.CLK(net4785),
    .RESET_B(net4107),
    .D(_02032_),
    .Q_N(_09103_),
    .Q(\spiking_network_top_uut.all_data_out[455] ));
 sg13g2_dfrbp_1 _20717_ (.CLK(net4703),
    .RESET_B(net4023),
    .D(_02033_),
    .Q_N(_09102_),
    .Q(\spiking_network_top_uut.all_data_out[0] ));
 sg13g2_dfrbp_1 _20718_ (.CLK(net4706),
    .RESET_B(net4026),
    .D(_02034_),
    .Q_N(_09101_),
    .Q(\spiking_network_top_uut.all_data_out[1] ));
 sg13g2_dfrbp_1 _20719_ (.CLK(net4703),
    .RESET_B(net4023),
    .D(_02035_),
    .Q_N(_00031_),
    .Q(\spiking_network_top_uut.all_data_out[2] ));
 sg13g2_dfrbp_1 _20720_ (.CLK(net4727),
    .RESET_B(net4047),
    .D(_02036_),
    .Q_N(_09100_),
    .Q(\spiking_network_top_uut.all_data_out[3] ));
 sg13g2_dfrbp_1 _20721_ (.CLK(net4704),
    .RESET_B(net4024),
    .D(_02037_),
    .Q_N(_09099_),
    .Q(\spiking_network_top_uut.all_data_out[4] ));
 sg13g2_dfrbp_1 _20722_ (.CLK(net4728),
    .RESET_B(net4048),
    .D(_02038_),
    .Q_N(_09098_),
    .Q(\spiking_network_top_uut.all_data_out[5] ));
 sg13g2_dfrbp_1 _20723_ (.CLK(net4728),
    .RESET_B(net4047),
    .D(_02039_),
    .Q_N(_09097_),
    .Q(\spiking_network_top_uut.all_data_out[6] ));
 sg13g2_dfrbp_1 _20724_ (.CLK(net4729),
    .RESET_B(net4049),
    .D(_02040_),
    .Q_N(_09096_),
    .Q(\spiking_network_top_uut.all_data_out[7] ));
 sg13g2_dfrbp_1 _20725_ (.CLK(net4747),
    .RESET_B(net4068),
    .D(_02041_),
    .Q_N(_09095_),
    .Q(\spiking_network_top_uut.spi_inst.memory_inst.addr_reg_out[0] ));
 sg13g2_dfrbp_1 _20726_ (.CLK(net4747),
    .RESET_B(net4068),
    .D(_02042_),
    .Q_N(_09094_),
    .Q(\spiking_network_top_uut.spi_inst.memory_inst.addr_reg_out[1] ));
 sg13g2_dfrbp_1 _20727_ (.CLK(net4742),
    .RESET_B(net4062),
    .D(_02043_),
    .Q_N(_09093_),
    .Q(\spiking_network_top_uut.spi_inst.memory_inst.addr_reg_out[2] ));
 sg13g2_dfrbp_1 _20728_ (.CLK(net4743),
    .RESET_B(net4062),
    .D(_02044_),
    .Q_N(_09092_),
    .Q(\spiking_network_top_uut.spi_inst.memory_inst.addr_reg_out[3] ));
 sg13g2_dfrbp_1 _20729_ (.CLK(net4742),
    .RESET_B(net4062),
    .D(_02045_),
    .Q_N(_09091_),
    .Q(\spiking_network_top_uut.spi_inst.memory_inst.addr_reg_out[4] ));
 sg13g2_dfrbp_1 _20730_ (.CLK(net4742),
    .RESET_B(net4062),
    .D(_02046_),
    .Q_N(_09090_),
    .Q(\spiking_network_top_uut.spi_inst.memory_inst.addr_reg_out[5] ));
 sg13g2_dfrbp_1 _20731_ (.CLK(net4743),
    .RESET_B(net4063),
    .D(_02047_),
    .Q_N(_00139_),
    .Q(\spiking_network_top_uut.spi_inst.memory_inst.addr_reg_out[6] ));
 sg13g2_dfrbp_1 _20732_ (.CLK(net4687),
    .RESET_B(net4006),
    .D(_02048_),
    .Q_N(_09089_),
    .Q(\spiking_network_top_uut.all_data_out[672] ));
 sg13g2_dfrbp_1 _20733_ (.CLK(net4689),
    .RESET_B(net4008),
    .D(_02049_),
    .Q_N(_00378_),
    .Q(\spiking_network_top_uut.all_data_out[673] ));
 sg13g2_dfrbp_1 _20734_ (.CLK(net4689),
    .RESET_B(net4008),
    .D(_02050_),
    .Q_N(_00308_),
    .Q(\spiking_network_top_uut.all_data_out[674] ));
 sg13g2_dfrbp_1 _20735_ (.CLK(net4682),
    .RESET_B(net4001),
    .D(_02051_),
    .Q_N(_09088_),
    .Q(\spiking_network_top_uut.all_data_out[675] ));
 sg13g2_dfrbp_1 _20736_ (.CLK(net4674),
    .RESET_B(net3993),
    .D(_02052_),
    .Q_N(_09087_),
    .Q(\spiking_network_top_uut.all_data_out[676] ));
 sg13g2_dfrbp_1 _20737_ (.CLK(net4694),
    .RESET_B(net4013),
    .D(_02053_),
    .Q_N(_00238_),
    .Q(\spiking_network_top_uut.all_data_out[677] ));
 sg13g2_dfrbp_1 _20738_ (.CLK(net4674),
    .RESET_B(net3993),
    .D(_02054_),
    .Q_N(_00168_),
    .Q(\spiking_network_top_uut.all_data_out[678] ));
 sg13g2_dfrbp_1 _20739_ (.CLK(net4682),
    .RESET_B(net4001),
    .D(_02055_),
    .Q_N(_09086_),
    .Q(\spiking_network_top_uut.all_data_out[679] ));
 sg13g2_dfrbp_1 _20740_ (.CLK(net4647),
    .RESET_B(net3967),
    .D(_02056_),
    .Q_N(_10359_),
    .Q(\spiking_network_top_uut.debug_config_ready_reg_out ));
 sg13g2_dfrbp_1 _20741_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1),
    .D(net26),
    .Q_N(_10360_),
    .Q(\spiking_network_top_uut.u_sys_clk_reset.reset_ff1 ));
 sg13g2_dfrbp_1 _20742_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1),
    .D(net35),
    .Q_N(_10361_),
    .Q(\spiking_network_top_uut.sys_clk_reset_synchr ));
 sg13g2_dfrbp_1 _20743_ (.CLK(net4648),
    .RESET_B(net1),
    .D(net27),
    .Q_N(_10362_),
    .Q(\spiking_network_top_uut.u_SPI_reset.reset_ff1 ));
 sg13g2_dfrbp_1 _20744_ (.CLK(net4648),
    .RESET_B(net1),
    .D(\spiking_network_top_uut.u_SPI_reset.reset_ff1 ),
    .Q_N(_10363_),
    .Q(\spiking_network_top_uut.SPI_reset_synchr ));
 sg13g2_dfrbp_1 _20745_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net4140),
    .D(\spiking_network_top_uut.debug_config_ready_reg_out ),
    .Q_N(_10364_),
    .Q(\spiking_network_top_uut.debug_config_sync.sync_ff1 ));
 sg13g2_dfrbp_1 _20746_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net4183),
    .D(\spiking_network_top_uut.clk_div_ready_reg_out ),
    .Q_N(_10365_),
    .Q(\spiking_network_top_uut.clk_div_sync.sync_ff1 ));
 sg13g2_dfrbp_1 _20747_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net4171),
    .D(net13),
    .Q_N(_10366_),
    .Q(\spiking_network_top_uut.snn_en_sync_inst.sync_ff1 ));
 sg13g2_dfrbp_1 _20748_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net4192),
    .D(net12),
    .Q_N(_09085_),
    .Q(\spiking_network_top_uut.input_ready_sync_inst.sync_ff1 ));
 sg13g2_tiehi _20743__27 (.L_HI(net27));
 sg13g2_tiehi tt_um_snn_with_delays_paolaunisa_28 (.L_HI(net28));
 sg13g2_tiehi tt_um_snn_with_delays_paolaunisa_29 (.L_HI(net29));
 sg13g2_tiehi tt_um_snn_with_delays_paolaunisa_30 (.L_HI(net30));
 sg13g2_buf_2 clkbuf_leaf_0_clk (.A(clknet_4_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_tielo tt_um_snn_with_delays_paolaunisa_17 (.L_LO(net17));
 sg13g2_tielo tt_um_snn_with_delays_paolaunisa_18 (.L_LO(net18));
 sg13g2_tielo tt_um_snn_with_delays_paolaunisa_19 (.L_LO(net19));
 sg13g2_tielo tt_um_snn_with_delays_paolaunisa_20 (.L_LO(net20));
 sg13g2_tielo tt_um_snn_with_delays_paolaunisa_21 (.L_LO(net21));
 sg13g2_tielo tt_um_snn_with_delays_paolaunisa_22 (.L_LO(net22));
 sg13g2_tielo tt_um_snn_with_delays_paolaunisa_23 (.L_LO(net23));
 sg13g2_tielo tt_um_snn_with_delays_paolaunisa_24 (.L_LO(net24));
 sg13g2_tielo tt_um_snn_with_delays_paolaunisa_25 (.L_LO(net25));
 sg13g2_tiehi _20741__26 (.L_HI(net26));
 sg13g2_buf_8 _20764_ (.A(MISO),
    .X(uio_out[2]));
 sg13g2_buf_4 _20765_ (.X(uio_out[5]),
    .A(output_ready));
 sg13g2_buf_8 _20766_ (.A(spi_instruction_done),
    .X(uio_out[7]));
 sg13g2_buf_2 fanout3616 (.A(_03171_),
    .X(net3616));
 sg13g2_buf_2 fanout3617 (.A(net3618),
    .X(net3617));
 sg13g2_buf_1 fanout3618 (.A(net3619),
    .X(net3618));
 sg13g2_buf_2 fanout3619 (.A(_04907_),
    .X(net3619));
 sg13g2_buf_2 fanout3620 (.A(net3621),
    .X(net3620));
 sg13g2_buf_1 fanout3621 (.A(net3622),
    .X(net3621));
 sg13g2_buf_2 fanout3622 (.A(_04894_),
    .X(net3622));
 sg13g2_buf_2 fanout3623 (.A(net3624),
    .X(net3623));
 sg13g2_buf_1 fanout3624 (.A(net3625),
    .X(net3624));
 sg13g2_buf_4 fanout3625 (.X(net3625),
    .A(_04854_));
 sg13g2_buf_2 fanout3626 (.A(net3627),
    .X(net3626));
 sg13g2_buf_1 fanout3627 (.A(net3628),
    .X(net3627));
 sg13g2_buf_2 fanout3628 (.A(_04841_),
    .X(net3628));
 sg13g2_buf_2 fanout3629 (.A(net3630),
    .X(net3629));
 sg13g2_buf_1 fanout3630 (.A(net3631),
    .X(net3630));
 sg13g2_buf_4 fanout3631 (.X(net3631),
    .A(_04743_));
 sg13g2_buf_2 fanout3632 (.A(net3633),
    .X(net3632));
 sg13g2_buf_1 fanout3633 (.A(net3634),
    .X(net3633));
 sg13g2_buf_4 fanout3634 (.X(net3634),
    .A(_04730_));
 sg13g2_buf_2 fanout3635 (.A(net3636),
    .X(net3635));
 sg13g2_buf_4 fanout3636 (.X(net3636),
    .A(_04966_));
 sg13g2_buf_2 fanout3637 (.A(net3638),
    .X(net3637));
 sg13g2_buf_1 fanout3638 (.A(net3639),
    .X(net3638));
 sg13g2_buf_2 fanout3639 (.A(_04951_),
    .X(net3639));
 sg13g2_buf_2 fanout3640 (.A(net3641),
    .X(net3640));
 sg13g2_buf_1 fanout3641 (.A(net3642),
    .X(net3641));
 sg13g2_buf_2 fanout3642 (.A(_04936_),
    .X(net3642));
 sg13g2_buf_2 fanout3643 (.A(net3644),
    .X(net3643));
 sg13g2_buf_1 fanout3644 (.A(net3645),
    .X(net3644));
 sg13g2_buf_2 fanout3645 (.A(_04921_),
    .X(net3645));
 sg13g2_buf_2 fanout3646 (.A(net3647),
    .X(net3646));
 sg13g2_buf_2 fanout3647 (.A(_04867_),
    .X(net3647));
 sg13g2_buf_2 fanout3648 (.A(net3649),
    .X(net3648));
 sg13g2_buf_1 fanout3649 (.A(net3650),
    .X(net3649));
 sg13g2_buf_4 fanout3650 (.X(net3650),
    .A(_04827_));
 sg13g2_buf_2 fanout3651 (.A(net3652),
    .X(net3651));
 sg13g2_buf_4 fanout3652 (.X(net3652),
    .A(_04813_));
 sg13g2_buf_2 fanout3653 (.A(net3654),
    .X(net3653));
 sg13g2_buf_1 fanout3654 (.A(net3655),
    .X(net3654));
 sg13g2_buf_2 fanout3655 (.A(_04800_),
    .X(net3655));
 sg13g2_buf_2 fanout3656 (.A(net3657),
    .X(net3656));
 sg13g2_buf_1 fanout3657 (.A(net3658),
    .X(net3657));
 sg13g2_buf_4 fanout3658 (.X(net3658),
    .A(_04786_));
 sg13g2_buf_2 fanout3659 (.A(net3660),
    .X(net3659));
 sg13g2_buf_1 fanout3660 (.A(net3661),
    .X(net3660));
 sg13g2_buf_4 fanout3661 (.X(net3661),
    .A(_04756_));
 sg13g2_buf_2 fanout3662 (.A(net3663),
    .X(net3662));
 sg13g2_buf_1 fanout3663 (.A(net3664),
    .X(net3663));
 sg13g2_buf_4 fanout3664 (.X(net3664),
    .A(_04881_));
 sg13g2_buf_2 fanout3665 (.A(net3666),
    .X(net3665));
 sg13g2_buf_4 fanout3666 (.X(net3666),
    .A(_04771_));
 sg13g2_buf_4 fanout3667 (.X(net3667),
    .A(_04646_));
 sg13g2_buf_4 fanout3668 (.X(net3668),
    .A(_03384_));
 sg13g2_buf_4 fanout3669 (.X(net3669),
    .A(_03382_));
 sg13g2_buf_8 fanout3670 (.A(_03378_),
    .X(net3670));
 sg13g2_buf_2 fanout3671 (.A(_03373_),
    .X(net3671));
 sg13g2_buf_4 fanout3672 (.X(net3672),
    .A(_03371_));
 sg13g2_buf_4 fanout3673 (.X(net3673),
    .A(_03360_));
 sg13g2_buf_4 fanout3674 (.X(net3674),
    .A(_03349_));
 sg13g2_buf_8 fanout3675 (.A(_03341_),
    .X(net3675));
 sg13g2_buf_4 fanout3676 (.X(net3676),
    .A(_03334_));
 sg13g2_buf_4 fanout3677 (.X(net3677),
    .A(_03331_));
 sg13g2_buf_4 fanout3678 (.X(net3678),
    .A(_03328_));
 sg13g2_buf_8 fanout3679 (.A(_03325_),
    .X(net3679));
 sg13g2_buf_8 fanout3680 (.A(_03322_),
    .X(net3680));
 sg13g2_buf_4 fanout3681 (.X(net3681),
    .A(_03315_));
 sg13g2_buf_8 fanout3682 (.A(_03294_),
    .X(net3682));
 sg13g2_buf_8 fanout3683 (.A(_03283_),
    .X(net3683));
 sg13g2_buf_4 fanout3684 (.X(net3684),
    .A(_03276_));
 sg13g2_buf_8 fanout3685 (.A(_03266_),
    .X(net3685));
 sg13g2_buf_8 fanout3686 (.A(_03263_),
    .X(net3686));
 sg13g2_buf_4 fanout3687 (.X(net3687),
    .A(_03261_));
 sg13g2_buf_4 fanout3688 (.X(net3688),
    .A(_03259_));
 sg13g2_buf_4 fanout3689 (.X(net3689),
    .A(_03246_));
 sg13g2_buf_8 fanout3690 (.A(_03228_),
    .X(net3690));
 sg13g2_buf_8 fanout3691 (.A(_03226_),
    .X(net3691));
 sg13g2_buf_4 fanout3692 (.X(net3692),
    .A(_03219_));
 sg13g2_buf_8 fanout3693 (.A(_03750_),
    .X(net3693));
 sg13g2_buf_8 fanout3694 (.A(_03748_),
    .X(net3694));
 sg13g2_buf_8 fanout3695 (.A(_03747_),
    .X(net3695));
 sg13g2_buf_4 fanout3696 (.X(net3696),
    .A(_03740_));
 sg13g2_buf_8 fanout3697 (.A(_03306_),
    .X(net3697));
 sg13g2_buf_8 fanout3698 (.A(_03301_),
    .X(net3698));
 sg13g2_buf_4 fanout3699 (.X(net3699),
    .A(_02942_));
 sg13g2_buf_2 fanout3700 (.A(_02348_),
    .X(net3700));
 sg13g2_buf_2 fanout3701 (.A(_02065_),
    .X(net3701));
 sg13g2_buf_4 fanout3702 (.X(net3702),
    .A(_08230_));
 sg13g2_buf_2 fanout3703 (.A(_07663_),
    .X(net3703));
 sg13g2_buf_2 fanout3704 (.A(_07366_),
    .X(net3704));
 sg13g2_buf_4 fanout3705 (.X(net3705),
    .A(_06228_));
 sg13g2_buf_4 fanout3706 (.X(net3706),
    .A(_04613_));
 sg13g2_buf_4 fanout3707 (.X(net3707),
    .A(_03749_));
 sg13g2_buf_4 fanout3708 (.X(net3708),
    .A(_03746_));
 sg13g2_buf_8 fanout3709 (.A(_03742_),
    .X(net3709));
 sg13g2_buf_8 fanout3710 (.A(_03737_),
    .X(net3710));
 sg13g2_buf_4 fanout3711 (.X(net3711),
    .A(_03732_));
 sg13g2_buf_4 fanout3712 (.X(net3712),
    .A(_03730_));
 sg13g2_buf_4 fanout3713 (.X(net3713),
    .A(_03728_));
 sg13g2_buf_8 fanout3714 (.A(_03725_),
    .X(net3714));
 sg13g2_buf_8 fanout3715 (.A(_03723_),
    .X(net3715));
 sg13g2_buf_4 fanout3716 (.X(net3716),
    .A(_03715_));
 sg13g2_buf_4 fanout3717 (.X(net3717),
    .A(_03713_));
 sg13g2_buf_4 fanout3718 (.X(net3718),
    .A(_03709_));
 sg13g2_buf_8 fanout3719 (.A(_03706_),
    .X(net3719));
 sg13g2_buf_4 fanout3720 (.X(net3720),
    .A(net3722));
 sg13g2_buf_1 fanout3721 (.A(net3722),
    .X(net3721));
 sg13g2_buf_2 fanout3722 (.A(_00026_),
    .X(net3722));
 sg13g2_buf_8 fanout3723 (.A(net3724),
    .X(net3723));
 sg13g2_buf_8 fanout3724 (.A(_03345_),
    .X(net3724));
 sg13g2_buf_8 fanout3725 (.A(net3726),
    .X(net3725));
 sg13g2_buf_4 fanout3726 (.X(net3726),
    .A(_03304_));
 sg13g2_buf_4 fanout3727 (.X(net3727),
    .A(net3728));
 sg13g2_buf_8 fanout3728 (.A(_03300_),
    .X(net3728));
 sg13g2_buf_8 fanout3729 (.A(_03255_),
    .X(net3729));
 sg13g2_buf_4 fanout3730 (.X(net3730),
    .A(_03255_));
 sg13g2_buf_8 fanout3731 (.A(_03224_),
    .X(net3731));
 sg13g2_buf_4 fanout3732 (.X(net3732),
    .A(_03224_));
 sg13g2_buf_8 fanout3733 (.A(net3734),
    .X(net3733));
 sg13g2_buf_16 fanout3734 (.X(net3734),
    .A(_03211_));
 sg13g2_buf_4 fanout3735 (.X(net3735),
    .A(net3736));
 sg13g2_buf_8 fanout3736 (.A(_03206_),
    .X(net3736));
 sg13g2_buf_4 fanout3737 (.X(net3737),
    .A(_03199_));
 sg13g2_buf_8 fanout3738 (.A(net3739),
    .X(net3738));
 sg13g2_buf_8 fanout3739 (.A(_05097_),
    .X(net3739));
 sg13g2_buf_8 fanout3740 (.A(_05089_),
    .X(net3740));
 sg13g2_buf_4 fanout3741 (.X(net3741),
    .A(_05089_));
 sg13g2_buf_4 fanout3742 (.X(net3742),
    .A(net3750));
 sg13g2_buf_4 fanout3743 (.X(net3743),
    .A(net3750));
 sg13g2_buf_2 fanout3744 (.A(net3745),
    .X(net3744));
 sg13g2_buf_2 fanout3745 (.A(net3750),
    .X(net3745));
 sg13g2_buf_2 fanout3746 (.A(net3750),
    .X(net3746));
 sg13g2_buf_1 fanout3747 (.A(net3750),
    .X(net3747));
 sg13g2_buf_4 fanout3748 (.X(net3748),
    .A(net3749));
 sg13g2_buf_4 fanout3749 (.X(net3749),
    .A(net3750));
 sg13g2_buf_8 fanout3750 (.A(_05085_),
    .X(net3750));
 sg13g2_buf_2 fanout3751 (.A(net3752),
    .X(net3751));
 sg13g2_buf_2 fanout3752 (.A(net3755),
    .X(net3752));
 sg13g2_buf_2 fanout3753 (.A(net3754),
    .X(net3753));
 sg13g2_buf_2 fanout3754 (.A(net3755),
    .X(net3754));
 sg13g2_buf_2 fanout3755 (.A(_05085_),
    .X(net3755));
 sg13g2_buf_4 fanout3756 (.X(net3756),
    .A(_04603_));
 sg13g2_buf_4 fanout3757 (.X(net3757),
    .A(net3759));
 sg13g2_buf_2 fanout3758 (.A(net3759),
    .X(net3758));
 sg13g2_buf_4 fanout3759 (.X(net3759),
    .A(_03774_));
 sg13g2_buf_4 fanout3760 (.X(net3760),
    .A(net3761));
 sg13g2_buf_4 fanout3761 (.X(net3761),
    .A(net3762));
 sg13g2_buf_2 fanout3762 (.A(_03771_),
    .X(net3762));
 sg13g2_buf_4 fanout3763 (.X(net3763),
    .A(net3764));
 sg13g2_buf_2 fanout3764 (.A(_03766_),
    .X(net3764));
 sg13g2_buf_4 fanout3765 (.X(net3765),
    .A(_03766_));
 sg13g2_buf_4 fanout3766 (.X(net3766),
    .A(net3767));
 sg13g2_buf_4 fanout3767 (.X(net3767),
    .A(_03762_));
 sg13g2_buf_4 fanout3768 (.X(net3768),
    .A(net3770));
 sg13g2_buf_2 fanout3769 (.A(net3770),
    .X(net3769));
 sg13g2_buf_4 fanout3770 (.X(net3770),
    .A(_03759_));
 sg13g2_buf_4 fanout3771 (.X(net3771),
    .A(_03741_));
 sg13g2_buf_4 fanout3772 (.X(net3772),
    .A(_03733_));
 sg13g2_buf_4 fanout3773 (.X(net3773),
    .A(_03731_));
 sg13g2_buf_8 fanout3774 (.A(_03727_),
    .X(net3774));
 sg13g2_buf_4 fanout3775 (.X(net3775),
    .A(net3777));
 sg13g2_buf_4 fanout3776 (.X(net3776),
    .A(net3777));
 sg13g2_buf_4 fanout3777 (.X(net3777),
    .A(_03719_));
 sg13g2_buf_4 fanout3778 (.X(net3778),
    .A(_03714_));
 sg13g2_buf_4 fanout3779 (.X(net3779),
    .A(_03708_));
 sg13g2_buf_4 fanout3780 (.X(net3780),
    .A(_03705_));
 sg13g2_buf_4 fanout3781 (.X(net3781),
    .A(_03703_));
 sg13g2_buf_4 fanout3782 (.X(net3782),
    .A(_03703_));
 sg13g2_buf_2 fanout3783 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[6] ),
    .X(net3783));
 sg13g2_buf_2 fanout3784 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[5] ),
    .X(net3784));
 sg13g2_buf_2 fanout3785 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[4] ),
    .X(net3785));
 sg13g2_buf_2 fanout3786 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[3] ),
    .X(net3786));
 sg13g2_buf_2 fanout3787 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[2] ),
    .X(net3787));
 sg13g2_buf_2 fanout3788 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[1] ),
    .X(net3788));
 sg13g2_buf_2 fanout3789 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[0] ),
    .X(net3789));
 sg13g2_buf_4 fanout3790 (.X(net3790),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[7] ));
 sg13g2_buf_2 fanout3791 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[6] ),
    .X(net3791));
 sg13g2_buf_4 fanout3792 (.X(net3792),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[4] ));
 sg13g2_buf_4 fanout3793 (.X(net3793),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[3] ));
 sg13g2_buf_2 fanout3794 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[2] ),
    .X(net3794));
 sg13g2_buf_4 fanout3795 (.X(net3795),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[1] ));
 sg13g2_buf_2 fanout3796 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[0] ),
    .X(net3796));
 sg13g2_buf_4 fanout3797 (.X(net3797),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[7] ));
 sg13g2_buf_4 fanout3798 (.X(net3798),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[6] ));
 sg13g2_buf_4 fanout3799 (.X(net3799),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[5] ));
 sg13g2_buf_4 fanout3800 (.X(net3800),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[4] ));
 sg13g2_buf_2 fanout3801 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[3] ),
    .X(net3801));
 sg13g2_buf_2 fanout3802 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[2] ),
    .X(net3802));
 sg13g2_buf_2 fanout3803 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[1] ),
    .X(net3803));
 sg13g2_buf_2 fanout3804 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[0] ),
    .X(net3804));
 sg13g2_buf_4 fanout3805 (.X(net3805),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[7] ));
 sg13g2_buf_4 fanout3806 (.X(net3806),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[6] ));
 sg13g2_buf_2 fanout3807 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[5] ),
    .X(net3807));
 sg13g2_buf_2 fanout3808 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[4] ),
    .X(net3808));
 sg13g2_buf_2 fanout3809 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[3] ),
    .X(net3809));
 sg13g2_buf_2 fanout3810 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[2] ),
    .X(net3810));
 sg13g2_buf_2 fanout3811 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[1] ),
    .X(net3811));
 sg13g2_buf_2 fanout3812 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[0] ),
    .X(net3812));
 sg13g2_buf_4 fanout3813 (.X(net3813),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[7] ));
 sg13g2_buf_4 fanout3814 (.X(net3814),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[6] ));
 sg13g2_buf_2 fanout3815 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[4] ),
    .X(net3815));
 sg13g2_buf_2 fanout3816 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[3] ),
    .X(net3816));
 sg13g2_buf_2 fanout3817 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[2] ),
    .X(net3817));
 sg13g2_buf_2 fanout3818 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[1] ),
    .X(net3818));
 sg13g2_buf_2 fanout3819 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[0] ),
    .X(net3819));
 sg13g2_buf_4 fanout3820 (.X(net3820),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[7] ));
 sg13g2_buf_2 fanout3821 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[6] ),
    .X(net3821));
 sg13g2_buf_4 fanout3822 (.X(net3822),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[4] ));
 sg13g2_buf_2 fanout3823 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[3] ),
    .X(net3823));
 sg13g2_buf_2 fanout3824 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[2] ),
    .X(net3824));
 sg13g2_buf_2 fanout3825 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[1] ),
    .X(net3825));
 sg13g2_buf_2 fanout3826 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[0] ),
    .X(net3826));
 sg13g2_buf_4 fanout3827 (.X(net3827),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[7] ));
 sg13g2_buf_4 fanout3828 (.X(net3828),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[6] ));
 sg13g2_buf_2 fanout3829 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[4] ),
    .X(net3829));
 sg13g2_buf_2 fanout3830 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[3] ),
    .X(net3830));
 sg13g2_buf_2 fanout3831 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[2] ),
    .X(net3831));
 sg13g2_buf_2 fanout3832 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[1] ),
    .X(net3832));
 sg13g2_buf_2 fanout3833 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[0] ),
    .X(net3833));
 sg13g2_buf_2 fanout3834 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[7] ),
    .X(net3834));
 sg13g2_buf_2 fanout3835 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[6] ),
    .X(net3835));
 sg13g2_buf_2 fanout3836 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[4] ),
    .X(net3836));
 sg13g2_buf_4 fanout3837 (.X(net3837),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[3] ));
 sg13g2_buf_2 fanout3838 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[2] ),
    .X(net3838));
 sg13g2_buf_2 fanout3839 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[1] ),
    .X(net3839));
 sg13g2_buf_2 fanout3840 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[0] ),
    .X(net3840));
 sg13g2_buf_4 fanout3841 (.X(net3841),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[6] ));
 sg13g2_buf_2 fanout3842 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[4] ),
    .X(net3842));
 sg13g2_buf_4 fanout3843 (.X(net3843),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[3] ));
 sg13g2_buf_4 fanout3844 (.X(net3844),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[2] ));
 sg13g2_buf_2 fanout3845 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[1] ),
    .X(net3845));
 sg13g2_buf_2 fanout3846 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[0] ),
    .X(net3846));
 sg13g2_buf_4 fanout3847 (.X(net3847),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[7] ));
 sg13g2_buf_4 fanout3848 (.X(net3848),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[6] ));
 sg13g2_buf_4 fanout3849 (.X(net3849),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[4] ));
 sg13g2_buf_4 fanout3850 (.X(net3850),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[3] ));
 sg13g2_buf_4 fanout3851 (.X(net3851),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[2] ));
 sg13g2_buf_2 fanout3852 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[1] ),
    .X(net3852));
 sg13g2_buf_2 fanout3853 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.pd.shift_reg[0] ),
    .X(net3853));
 sg13g2_buf_4 fanout3854 (.X(net3854),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[7] ));
 sg13g2_buf_4 fanout3855 (.X(net3855),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[6] ));
 sg13g2_buf_4 fanout3856 (.X(net3856),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[4] ));
 sg13g2_buf_4 fanout3857 (.X(net3857),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[3] ));
 sg13g2_buf_4 fanout3858 (.X(net3858),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[2] ));
 sg13g2_buf_4 fanout3859 (.X(net3859),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[1] ));
 sg13g2_buf_4 fanout3860 (.X(net3860),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.pd.shift_reg[0] ));
 sg13g2_buf_4 fanout3861 (.X(net3861),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[7] ));
 sg13g2_buf_4 fanout3862 (.X(net3862),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[6] ));
 sg13g2_buf_2 fanout3863 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[5] ),
    .X(net3863));
 sg13g2_buf_4 fanout3864 (.X(net3864),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[4] ));
 sg13g2_buf_2 fanout3865 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[3] ),
    .X(net3865));
 sg13g2_buf_2 fanout3866 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[2] ),
    .X(net3866));
 sg13g2_buf_2 fanout3867 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[1] ),
    .X(net3867));
 sg13g2_buf_2 fanout3868 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.pd.shift_reg[0] ),
    .X(net3868));
 sg13g2_buf_4 fanout3869 (.X(net3869),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[7] ));
 sg13g2_buf_4 fanout3870 (.X(net3870),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[6] ));
 sg13g2_buf_4 fanout3871 (.X(net3871),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[5] ));
 sg13g2_buf_2 fanout3872 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[4] ),
    .X(net3872));
 sg13g2_buf_2 fanout3873 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[3] ),
    .X(net3873));
 sg13g2_buf_2 fanout3874 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[2] ),
    .X(net3874));
 sg13g2_buf_2 fanout3875 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[1] ),
    .X(net3875));
 sg13g2_buf_2 fanout3876 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.pd.shift_reg[0] ),
    .X(net3876));
 sg13g2_buf_4 fanout3877 (.X(net3877),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[7] ));
 sg13g2_buf_4 fanout3878 (.X(net3878),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[6] ));
 sg13g2_buf_4 fanout3879 (.X(net3879),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[5] ));
 sg13g2_buf_2 fanout3880 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[4] ),
    .X(net3880));
 sg13g2_buf_2 fanout3881 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[3] ),
    .X(net3881));
 sg13g2_buf_2 fanout3882 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[2] ),
    .X(net3882));
 sg13g2_buf_2 fanout3883 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[1] ),
    .X(net3883));
 sg13g2_buf_2 fanout3884 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.pd.shift_reg[0] ),
    .X(net3884));
 sg13g2_buf_4 fanout3885 (.X(net3885),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[7] ));
 sg13g2_buf_2 fanout3886 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[6] ),
    .X(net3886));
 sg13g2_buf_4 fanout3887 (.X(net3887),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[4] ));
 sg13g2_buf_2 fanout3888 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[3] ),
    .X(net3888));
 sg13g2_buf_2 fanout3889 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[2] ),
    .X(net3889));
 sg13g2_buf_2 fanout3890 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[1] ),
    .X(net3890));
 sg13g2_buf_2 fanout3891 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.pd.shift_reg[0] ),
    .X(net3891));
 sg13g2_buf_4 fanout3892 (.X(net3892),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[7] ));
 sg13g2_buf_4 fanout3893 (.X(net3893),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[6] ));
 sg13g2_buf_2 fanout3894 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[4] ),
    .X(net3894));
 sg13g2_buf_4 fanout3895 (.X(net3895),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[3] ));
 sg13g2_buf_2 fanout3896 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[2] ),
    .X(net3896));
 sg13g2_buf_4 fanout3897 (.X(net3897),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[1] ));
 sg13g2_buf_2 fanout3898 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.pd.shift_reg[0] ),
    .X(net3898));
 sg13g2_buf_4 fanout3899 (.X(net3899),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[7] ));
 sg13g2_buf_4 fanout3900 (.X(net3900),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.pd.shift_reg[7] ));
 sg13g2_buf_8 fanout3901 (.A(_05104_),
    .X(net3901));
 sg13g2_buf_4 fanout3902 (.X(net3902),
    .A(_05104_));
 sg13g2_buf_4 fanout3903 (.X(net3903),
    .A(net3906));
 sg13g2_buf_2 fanout3904 (.A(net3906),
    .X(net3904));
 sg13g2_buf_8 fanout3905 (.A(net3906),
    .X(net3905));
 sg13g2_buf_4 fanout3906 (.X(net3906),
    .A(_05098_));
 sg13g2_buf_4 fanout3907 (.X(net3907),
    .A(net3908));
 sg13g2_buf_4 fanout3908 (.X(net3908),
    .A(_05098_));
 sg13g2_buf_4 fanout3909 (.X(net3909),
    .A(net3910));
 sg13g2_buf_8 fanout3910 (.A(net3912),
    .X(net3910));
 sg13g2_buf_4 fanout3911 (.X(net3911),
    .A(net3912));
 sg13g2_buf_8 fanout3912 (.A(_05088_),
    .X(net3912));
 sg13g2_buf_4 fanout3913 (.X(net3913),
    .A(net3914));
 sg13g2_buf_4 fanout3914 (.X(net3914),
    .A(net3915));
 sg13g2_buf_8 fanout3915 (.A(_05087_),
    .X(net3915));
 sg13g2_buf_4 fanout3916 (.X(net3916),
    .A(net3917));
 sg13g2_buf_4 fanout3917 (.X(net3917),
    .A(net3918));
 sg13g2_buf_4 fanout3918 (.X(net3918),
    .A(_05086_));
 sg13g2_buf_4 fanout3919 (.X(net3919),
    .A(_03729_));
 sg13g2_buf_2 fanout3920 (.A(net3921),
    .X(net3920));
 sg13g2_buf_2 fanout3921 (.A(net3922),
    .X(net3921));
 sg13g2_buf_4 fanout3922 (.X(net3922),
    .A(net3931));
 sg13g2_buf_2 fanout3923 (.A(net3924),
    .X(net3923));
 sg13g2_buf_4 fanout3924 (.X(net3924),
    .A(net3931));
 sg13g2_buf_2 fanout3925 (.A(net3926),
    .X(net3925));
 sg13g2_buf_2 fanout3926 (.A(net3927),
    .X(net3926));
 sg13g2_buf_4 fanout3927 (.X(net3927),
    .A(net3931));
 sg13g2_buf_2 fanout3928 (.A(net3931),
    .X(net3928));
 sg13g2_buf_2 fanout3929 (.A(net3931),
    .X(net3929));
 sg13g2_buf_2 fanout3930 (.A(net3931),
    .X(net3930));
 sg13g2_buf_8 fanout3931 (.A(net3932),
    .X(net3931));
 sg13g2_buf_8 fanout3932 (.A(_03418_),
    .X(net3932));
 sg13g2_buf_4 fanout3933 (.X(net3933),
    .A(net3939));
 sg13g2_buf_4 fanout3934 (.X(net3934),
    .A(net3939));
 sg13g2_buf_4 fanout3935 (.X(net3935),
    .A(net3937));
 sg13g2_buf_2 fanout3936 (.A(net3937),
    .X(net3936));
 sg13g2_buf_4 fanout3937 (.X(net3937),
    .A(net3939));
 sg13g2_buf_4 fanout3938 (.X(net3938),
    .A(net3939));
 sg13g2_buf_8 fanout3939 (.A(_03418_),
    .X(net3939));
 sg13g2_buf_2 fanout3940 (.A(net3942),
    .X(net3940));
 sg13g2_buf_4 fanout3941 (.X(net3941),
    .A(net3942));
 sg13g2_buf_2 fanout3942 (.A(net3943),
    .X(net3942));
 sg13g2_buf_2 fanout3943 (.A(net3946),
    .X(net3943));
 sg13g2_buf_4 fanout3944 (.X(net3944),
    .A(net3946));
 sg13g2_buf_4 fanout3945 (.X(net3945),
    .A(net3946));
 sg13g2_buf_4 fanout3946 (.X(net3946),
    .A(_03412_));
 sg13g2_buf_4 fanout3947 (.X(net3947),
    .A(net3948));
 sg13g2_buf_2 fanout3948 (.A(net3949),
    .X(net3948));
 sg13g2_buf_4 fanout3949 (.X(net3949),
    .A(net3958));
 sg13g2_buf_2 fanout3950 (.A(net3951),
    .X(net3950));
 sg13g2_buf_2 fanout3951 (.A(net3958),
    .X(net3951));
 sg13g2_buf_2 fanout3952 (.A(net3954),
    .X(net3952));
 sg13g2_buf_2 fanout3953 (.A(net3954),
    .X(net3953));
 sg13g2_buf_2 fanout3954 (.A(net3955),
    .X(net3954));
 sg13g2_buf_2 fanout3955 (.A(net3958),
    .X(net3955));
 sg13g2_buf_4 fanout3956 (.X(net3956),
    .A(net3957));
 sg13g2_buf_2 fanout3957 (.A(net3958),
    .X(net3957));
 sg13g2_buf_8 fanout3958 (.A(_03402_),
    .X(net3958));
 sg13g2_buf_4 fanout3959 (.X(net3959),
    .A(net3960));
 sg13g2_buf_4 fanout3960 (.X(net3960),
    .A(net3965));
 sg13g2_buf_4 fanout3961 (.X(net3961),
    .A(net3964));
 sg13g2_buf_4 fanout3962 (.X(net3962),
    .A(net3964));
 sg13g2_buf_2 fanout3963 (.A(net3964),
    .X(net3963));
 sg13g2_buf_4 fanout3964 (.X(net3964),
    .A(net3965));
 sg13g2_buf_8 fanout3965 (.A(net3966),
    .X(net3965));
 sg13g2_buf_8 fanout3966 (.A(_03402_),
    .X(net3966));
 sg13g2_buf_8 fanout3967 (.A(net3979),
    .X(net3967));
 sg13g2_buf_4 fanout3968 (.X(net3968),
    .A(net3972));
 sg13g2_buf_2 fanout3969 (.A(net3972),
    .X(net3969));
 sg13g2_buf_4 fanout3970 (.X(net3970),
    .A(net3972));
 sg13g2_buf_4 fanout3971 (.X(net3971),
    .A(net3972));
 sg13g2_buf_2 fanout3972 (.A(net3978),
    .X(net3972));
 sg13g2_buf_4 fanout3973 (.X(net3973),
    .A(net3977));
 sg13g2_buf_2 fanout3974 (.A(net3977),
    .X(net3974));
 sg13g2_buf_4 fanout3975 (.X(net3975),
    .A(net3976));
 sg13g2_buf_4 fanout3976 (.X(net3976),
    .A(net3977));
 sg13g2_buf_2 fanout3977 (.A(net3978),
    .X(net3977));
 sg13g2_buf_4 fanout3978 (.X(net3978),
    .A(net3979));
 sg13g2_buf_2 fanout3979 (.A(net4136),
    .X(net3979));
 sg13g2_buf_4 fanout3980 (.X(net3980),
    .A(net3983));
 sg13g2_buf_4 fanout3981 (.X(net3981),
    .A(net3982));
 sg13g2_buf_4 fanout3982 (.X(net3982),
    .A(net3983));
 sg13g2_buf_4 fanout3983 (.X(net3983),
    .A(net4029));
 sg13g2_buf_4 fanout3984 (.X(net3984),
    .A(net3985));
 sg13g2_buf_4 fanout3985 (.X(net3985),
    .A(net3989));
 sg13g2_buf_4 fanout3986 (.X(net3986),
    .A(net3987));
 sg13g2_buf_4 fanout3987 (.X(net3987),
    .A(net3989));
 sg13g2_buf_4 fanout3988 (.X(net3988),
    .A(net3989));
 sg13g2_buf_4 fanout3989 (.X(net3989),
    .A(net4029));
 sg13g2_buf_4 fanout3990 (.X(net3990),
    .A(net3996));
 sg13g2_buf_4 fanout3991 (.X(net3991),
    .A(net3996));
 sg13g2_buf_4 fanout3992 (.X(net3992),
    .A(net3994));
 sg13g2_buf_4 fanout3993 (.X(net3993),
    .A(net3994));
 sg13g2_buf_2 fanout3994 (.A(net3995),
    .X(net3994));
 sg13g2_buf_4 fanout3995 (.X(net3995),
    .A(net3996));
 sg13g2_buf_2 fanout3996 (.A(net4029),
    .X(net3996));
 sg13g2_buf_4 fanout3997 (.X(net3997),
    .A(net3999));
 sg13g2_buf_4 fanout3998 (.X(net3998),
    .A(net3999));
 sg13g2_buf_4 fanout3999 (.X(net3999),
    .A(net4010));
 sg13g2_buf_4 fanout4000 (.X(net4000),
    .A(net4003));
 sg13g2_buf_2 fanout4001 (.A(net4003),
    .X(net4001));
 sg13g2_buf_4 fanout4002 (.X(net4002),
    .A(net4003));
 sg13g2_buf_2 fanout4003 (.A(net4010),
    .X(net4003));
 sg13g2_buf_4 fanout4004 (.X(net4004),
    .A(net4005));
 sg13g2_buf_4 fanout4005 (.X(net4005),
    .A(net4009));
 sg13g2_buf_4 fanout4006 (.X(net4006),
    .A(net4009));
 sg13g2_buf_2 fanout4007 (.A(net4009),
    .X(net4007));
 sg13g2_buf_4 fanout4008 (.X(net4008),
    .A(net4009));
 sg13g2_buf_2 fanout4009 (.A(net4010),
    .X(net4009));
 sg13g2_buf_2 fanout4010 (.A(net4028),
    .X(net4010));
 sg13g2_buf_4 fanout4011 (.X(net4011),
    .A(net4012));
 sg13g2_buf_4 fanout4012 (.X(net4012),
    .A(net4013));
 sg13g2_buf_4 fanout4013 (.X(net4013),
    .A(net4017));
 sg13g2_buf_4 fanout4014 (.X(net4014),
    .A(net4015));
 sg13g2_buf_4 fanout4015 (.X(net4015),
    .A(net4016));
 sg13g2_buf_4 fanout4016 (.X(net4016),
    .A(net4017));
 sg13g2_buf_2 fanout4017 (.A(net4028),
    .X(net4017));
 sg13g2_buf_4 fanout4018 (.X(net4018),
    .A(net4022));
 sg13g2_buf_4 fanout4019 (.X(net4019),
    .A(net4022));
 sg13g2_buf_4 fanout4020 (.X(net4020),
    .A(net4022));
 sg13g2_buf_4 fanout4021 (.X(net4021),
    .A(net4022));
 sg13g2_buf_2 fanout4022 (.A(net4028),
    .X(net4022));
 sg13g2_buf_4 fanout4023 (.X(net4023),
    .A(net4027));
 sg13g2_buf_4 fanout4024 (.X(net4024),
    .A(net4025));
 sg13g2_buf_2 fanout4025 (.A(net4026),
    .X(net4025));
 sg13g2_buf_4 fanout4026 (.X(net4026),
    .A(net4027));
 sg13g2_buf_2 fanout4027 (.A(net4028),
    .X(net4027));
 sg13g2_buf_4 fanout4028 (.X(net4028),
    .A(net4029));
 sg13g2_buf_2 fanout4029 (.A(net4136),
    .X(net4029));
 sg13g2_buf_4 fanout4030 (.X(net4030),
    .A(net4031));
 sg13g2_buf_4 fanout4031 (.X(net4031),
    .A(net4042));
 sg13g2_buf_4 fanout4032 (.X(net4032),
    .A(net4034));
 sg13g2_buf_4 fanout4033 (.X(net4033),
    .A(net4034));
 sg13g2_buf_2 fanout4034 (.A(net4042),
    .X(net4034));
 sg13g2_buf_4 fanout4035 (.X(net4035),
    .A(net4039));
 sg13g2_buf_4 fanout4036 (.X(net4036),
    .A(net4039));
 sg13g2_buf_4 fanout4037 (.X(net4037),
    .A(net4039));
 sg13g2_buf_4 fanout4038 (.X(net4038),
    .A(net4039));
 sg13g2_buf_2 fanout4039 (.A(net4042),
    .X(net4039));
 sg13g2_buf_4 fanout4040 (.X(net4040),
    .A(net4041));
 sg13g2_buf_4 fanout4041 (.X(net4041),
    .A(net4042));
 sg13g2_buf_2 fanout4042 (.A(net4085),
    .X(net4042));
 sg13g2_buf_4 fanout4043 (.X(net4043),
    .A(net4044));
 sg13g2_buf_4 fanout4044 (.X(net4044),
    .A(net4046));
 sg13g2_buf_4 fanout4045 (.X(net4045),
    .A(net4046));
 sg13g2_buf_2 fanout4046 (.A(net4059),
    .X(net4046));
 sg13g2_buf_4 fanout4047 (.X(net4047),
    .A(net4051));
 sg13g2_buf_2 fanout4048 (.A(net4051),
    .X(net4048));
 sg13g2_buf_4 fanout4049 (.X(net4049),
    .A(net4051));
 sg13g2_buf_2 fanout4050 (.A(net4051),
    .X(net4050));
 sg13g2_buf_2 fanout4051 (.A(net4059),
    .X(net4051));
 sg13g2_buf_4 fanout4052 (.X(net4052),
    .A(net4054));
 sg13g2_buf_4 fanout4053 (.X(net4053),
    .A(net4054));
 sg13g2_buf_4 fanout4054 (.X(net4054),
    .A(net4059));
 sg13g2_buf_4 fanout4055 (.X(net4055),
    .A(net4058));
 sg13g2_buf_2 fanout4056 (.A(net4058),
    .X(net4056));
 sg13g2_buf_4 fanout4057 (.X(net4057),
    .A(net4058));
 sg13g2_buf_2 fanout4058 (.A(net4059),
    .X(net4058));
 sg13g2_buf_2 fanout4059 (.A(net4085),
    .X(net4059));
 sg13g2_buf_4 fanout4060 (.X(net4060),
    .A(net4061));
 sg13g2_buf_4 fanout4061 (.X(net4061),
    .A(net4064));
 sg13g2_buf_4 fanout4062 (.X(net4062),
    .A(net4064));
 sg13g2_buf_4 fanout4063 (.X(net4063),
    .A(net4064));
 sg13g2_buf_2 fanout4064 (.A(net4070),
    .X(net4064));
 sg13g2_buf_4 fanout4065 (.X(net4065),
    .A(net4067));
 sg13g2_buf_4 fanout4066 (.X(net4066),
    .A(net4067));
 sg13g2_buf_4 fanout4067 (.X(net4067),
    .A(net4070));
 sg13g2_buf_4 fanout4068 (.X(net4068),
    .A(net4070));
 sg13g2_buf_2 fanout4069 (.A(net4070),
    .X(net4069));
 sg13g2_buf_2 fanout4070 (.A(net4085),
    .X(net4070));
 sg13g2_buf_4 fanout4071 (.X(net4071),
    .A(net4072));
 sg13g2_buf_4 fanout4072 (.X(net4072),
    .A(net4084));
 sg13g2_buf_4 fanout4073 (.X(net4073),
    .A(net4075));
 sg13g2_buf_4 fanout4074 (.X(net4074),
    .A(net4075));
 sg13g2_buf_2 fanout4075 (.A(net4084),
    .X(net4075));
 sg13g2_buf_4 fanout4076 (.X(net4076),
    .A(net4080));
 sg13g2_buf_2 fanout4077 (.A(net4080),
    .X(net4077));
 sg13g2_buf_4 fanout4078 (.X(net4078),
    .A(net4080));
 sg13g2_buf_4 fanout4079 (.X(net4079),
    .A(net4080));
 sg13g2_buf_2 fanout4080 (.A(net4084),
    .X(net4080));
 sg13g2_buf_4 fanout4081 (.X(net4081),
    .A(net4082));
 sg13g2_buf_2 fanout4082 (.A(net4083),
    .X(net4082));
 sg13g2_buf_4 fanout4083 (.X(net4083),
    .A(net4084));
 sg13g2_buf_2 fanout4084 (.A(net4085),
    .X(net4084));
 sg13g2_buf_8 fanout4085 (.A(net4136),
    .X(net4085));
 sg13g2_buf_4 fanout4086 (.X(net4086),
    .A(net4087));
 sg13g2_buf_4 fanout4087 (.X(net4087),
    .A(net4098));
 sg13g2_buf_4 fanout4088 (.X(net4088),
    .A(net4090));
 sg13g2_buf_2 fanout4089 (.A(net4090),
    .X(net4089));
 sg13g2_buf_4 fanout4090 (.X(net4090),
    .A(net4098));
 sg13g2_buf_4 fanout4091 (.X(net4091),
    .A(net4092));
 sg13g2_buf_4 fanout4092 (.X(net4092),
    .A(net4097));
 sg13g2_buf_4 fanout4093 (.X(net4093),
    .A(net4096));
 sg13g2_buf_4 fanout4094 (.X(net4094),
    .A(net4096));
 sg13g2_buf_4 fanout4095 (.X(net4095),
    .A(net4096));
 sg13g2_buf_2 fanout4096 (.A(net4097),
    .X(net4096));
 sg13g2_buf_2 fanout4097 (.A(net4098),
    .X(net4097));
 sg13g2_buf_2 fanout4098 (.A(net4110),
    .X(net4098));
 sg13g2_buf_4 fanout4099 (.X(net4099),
    .A(net4100));
 sg13g2_buf_4 fanout4100 (.X(net4100),
    .A(net4110));
 sg13g2_buf_4 fanout4101 (.X(net4101),
    .A(net4102));
 sg13g2_buf_2 fanout4102 (.A(net4104),
    .X(net4102));
 sg13g2_buf_4 fanout4103 (.X(net4103),
    .A(net4104));
 sg13g2_buf_2 fanout4104 (.A(net4110),
    .X(net4104));
 sg13g2_buf_4 fanout4105 (.X(net4105),
    .A(net4106));
 sg13g2_buf_4 fanout4106 (.X(net4106),
    .A(net4109));
 sg13g2_buf_4 fanout4107 (.X(net4107),
    .A(net4109));
 sg13g2_buf_4 fanout4108 (.X(net4108),
    .A(net4109));
 sg13g2_buf_2 fanout4109 (.A(net4110),
    .X(net4109));
 sg13g2_buf_4 fanout4110 (.X(net4110),
    .A(net4136));
 sg13g2_buf_4 fanout4111 (.X(net4111),
    .A(net4112));
 sg13g2_buf_4 fanout4112 (.X(net4112),
    .A(net4116));
 sg13g2_buf_4 fanout4113 (.X(net4113),
    .A(net4116));
 sg13g2_buf_2 fanout4114 (.A(net4116),
    .X(net4114));
 sg13g2_buf_4 fanout4115 (.X(net4115),
    .A(net4116));
 sg13g2_buf_2 fanout4116 (.A(net4135),
    .X(net4116));
 sg13g2_buf_4 fanout4117 (.X(net4117),
    .A(net4123));
 sg13g2_buf_4 fanout4118 (.X(net4118),
    .A(net4122));
 sg13g2_buf_4 fanout4119 (.X(net4119),
    .A(net4121));
 sg13g2_buf_4 fanout4120 (.X(net4120),
    .A(net4121));
 sg13g2_buf_2 fanout4121 (.A(net4122),
    .X(net4121));
 sg13g2_buf_2 fanout4122 (.A(net4123),
    .X(net4122));
 sg13g2_buf_4 fanout4123 (.X(net4123),
    .A(net4135));
 sg13g2_buf_4 fanout4124 (.X(net4124),
    .A(net4126));
 sg13g2_buf_4 fanout4125 (.X(net4125),
    .A(net4126));
 sg13g2_buf_2 fanout4126 (.A(net4128),
    .X(net4126));
 sg13g2_buf_4 fanout4127 (.X(net4127),
    .A(net4128));
 sg13g2_buf_2 fanout4128 (.A(net4135),
    .X(net4128));
 sg13g2_buf_4 fanout4129 (.X(net4129),
    .A(net4131));
 sg13g2_buf_4 fanout4130 (.X(net4130),
    .A(net4131));
 sg13g2_buf_2 fanout4131 (.A(net4134),
    .X(net4131));
 sg13g2_buf_4 fanout4132 (.X(net4132),
    .A(net4134));
 sg13g2_buf_4 fanout4133 (.X(net4133),
    .A(net4134));
 sg13g2_buf_4 fanout4134 (.X(net4134),
    .A(net4135));
 sg13g2_buf_4 fanout4135 (.X(net4135),
    .A(net4136));
 sg13g2_buf_16 fanout4136 (.X(net4136),
    .A(\spiking_network_top_uut.SPI_reset_synchr ));
 sg13g2_buf_4 fanout4137 (.X(net4137),
    .A(net4144));
 sg13g2_buf_2 fanout4138 (.A(net4144),
    .X(net4138));
 sg13g2_buf_4 fanout4139 (.X(net4139),
    .A(net4140));
 sg13g2_buf_4 fanout4140 (.X(net4140),
    .A(net4144));
 sg13g2_buf_4 fanout4141 (.X(net4141),
    .A(net4143));
 sg13g2_buf_4 fanout4142 (.X(net4142),
    .A(net4143));
 sg13g2_buf_4 fanout4143 (.X(net4143),
    .A(net4144));
 sg13g2_buf_2 fanout4144 (.A(net4162),
    .X(net4144));
 sg13g2_buf_4 fanout4145 (.X(net4145),
    .A(net4149));
 sg13g2_buf_8 fanout4146 (.A(net4149),
    .X(net4146));
 sg13g2_buf_8 fanout4147 (.A(net4148),
    .X(net4147));
 sg13g2_buf_4 fanout4148 (.X(net4148),
    .A(net4149));
 sg13g2_buf_4 fanout4149 (.X(net4149),
    .A(net4162));
 sg13g2_buf_4 fanout4150 (.X(net4150),
    .A(net4153));
 sg13g2_buf_4 fanout4151 (.X(net4151),
    .A(net4153));
 sg13g2_buf_4 fanout4152 (.X(net4152),
    .A(net4153));
 sg13g2_buf_2 fanout4153 (.A(net4162),
    .X(net4153));
 sg13g2_buf_4 fanout4154 (.X(net4154),
    .A(net4156));
 sg13g2_buf_4 fanout4155 (.X(net4155),
    .A(net4156));
 sg13g2_buf_4 fanout4156 (.X(net4156),
    .A(net4157));
 sg13g2_buf_4 fanout4157 (.X(net4157),
    .A(net4162));
 sg13g2_buf_8 fanout4158 (.A(net4161),
    .X(net4158));
 sg13g2_buf_4 fanout4159 (.X(net4159),
    .A(net4161));
 sg13g2_buf_4 fanout4160 (.X(net4160),
    .A(net4161));
 sg13g2_buf_2 fanout4161 (.A(net4162),
    .X(net4161));
 sg13g2_buf_4 fanout4162 (.X(net4162),
    .A(net4175));
 sg13g2_buf_4 fanout4163 (.X(net4163),
    .A(net4164));
 sg13g2_buf_4 fanout4164 (.X(net4164),
    .A(net4175));
 sg13g2_buf_4 fanout4165 (.X(net4165),
    .A(net4167));
 sg13g2_buf_4 fanout4166 (.X(net4166),
    .A(net4167));
 sg13g2_buf_2 fanout4167 (.A(net4175),
    .X(net4167));
 sg13g2_buf_8 fanout4168 (.A(net4169),
    .X(net4168));
 sg13g2_buf_4 fanout4169 (.X(net4169),
    .A(net4174));
 sg13g2_buf_4 fanout4170 (.X(net4170),
    .A(net4172));
 sg13g2_buf_4 fanout4171 (.X(net4171),
    .A(net4172));
 sg13g2_buf_2 fanout4172 (.A(net4174),
    .X(net4172));
 sg13g2_buf_4 fanout4173 (.X(net4173),
    .A(net4174));
 sg13g2_buf_4 fanout4174 (.X(net4174),
    .A(net4175));
 sg13g2_buf_8 fanout4175 (.A(net4261),
    .X(net4175));
 sg13g2_buf_4 fanout4176 (.X(net4176),
    .A(net4179));
 sg13g2_buf_2 fanout4177 (.A(net4179),
    .X(net4177));
 sg13g2_buf_4 fanout4178 (.X(net4178),
    .A(net4179));
 sg13g2_buf_2 fanout4179 (.A(net4181),
    .X(net4179));
 sg13g2_buf_8 fanout4180 (.A(net4181),
    .X(net4180));
 sg13g2_buf_2 fanout4181 (.A(net4186),
    .X(net4181));
 sg13g2_buf_4 fanout4182 (.X(net4182),
    .A(net4183));
 sg13g2_buf_4 fanout4183 (.X(net4183),
    .A(net4184));
 sg13g2_buf_4 fanout4184 (.X(net4184),
    .A(net4186));
 sg13g2_buf_4 fanout4185 (.X(net4185),
    .A(net4186));
 sg13g2_buf_4 fanout4186 (.X(net4186),
    .A(net4193));
 sg13g2_buf_4 fanout4187 (.X(net4187),
    .A(net4190));
 sg13g2_buf_4 fanout4188 (.X(net4188),
    .A(net4189));
 sg13g2_buf_4 fanout4189 (.X(net4189),
    .A(net4190));
 sg13g2_buf_2 fanout4190 (.A(net4193),
    .X(net4190));
 sg13g2_buf_8 fanout4191 (.A(net4193),
    .X(net4191));
 sg13g2_buf_4 fanout4192 (.X(net4192),
    .A(net4193));
 sg13g2_buf_2 fanout4193 (.A(net4261),
    .X(net4193));
 sg13g2_buf_4 fanout4194 (.X(net4194),
    .A(net4197));
 sg13g2_buf_4 fanout4195 (.X(net4195),
    .A(net4197));
 sg13g2_buf_4 fanout4196 (.X(net4196),
    .A(net4197));
 sg13g2_buf_2 fanout4197 (.A(net4203),
    .X(net4197));
 sg13g2_buf_4 fanout4198 (.X(net4198),
    .A(net4200));
 sg13g2_buf_2 fanout4199 (.A(net4200),
    .X(net4199));
 sg13g2_buf_4 fanout4200 (.X(net4200),
    .A(net4203));
 sg13g2_buf_4 fanout4201 (.X(net4201),
    .A(net4203));
 sg13g2_buf_4 fanout4202 (.X(net4202),
    .A(net4203));
 sg13g2_buf_8 fanout4203 (.A(net4261),
    .X(net4203));
 sg13g2_buf_4 fanout4204 (.X(net4204),
    .A(net4205));
 sg13g2_buf_4 fanout4205 (.X(net4205),
    .A(net4206));
 sg13g2_buf_4 fanout4206 (.X(net4206),
    .A(net4209));
 sg13g2_buf_4 fanout4207 (.X(net4207),
    .A(net4208));
 sg13g2_buf_4 fanout4208 (.X(net4208),
    .A(net4209));
 sg13g2_buf_8 fanout4209 (.A(net4260),
    .X(net4209));
 sg13g2_buf_4 fanout4210 (.X(net4210),
    .A(net4214));
 sg13g2_buf_4 fanout4211 (.X(net4211),
    .A(net4213));
 sg13g2_buf_2 fanout4212 (.A(net4213),
    .X(net4212));
 sg13g2_buf_4 fanout4213 (.X(net4213),
    .A(net4214));
 sg13g2_buf_2 fanout4214 (.A(net4260),
    .X(net4214));
 sg13g2_buf_4 fanout4215 (.X(net4215),
    .A(net4218));
 sg13g2_buf_4 fanout4216 (.X(net4216),
    .A(net4217));
 sg13g2_buf_4 fanout4217 (.X(net4217),
    .A(net4218));
 sg13g2_buf_4 fanout4218 (.X(net4218),
    .A(net4260));
 sg13g2_buf_4 fanout4219 (.X(net4219),
    .A(net4220));
 sg13g2_buf_2 fanout4220 (.A(net4221),
    .X(net4220));
 sg13g2_buf_4 fanout4221 (.X(net4221),
    .A(net4227));
 sg13g2_buf_4 fanout4222 (.X(net4222),
    .A(net4227));
 sg13g2_buf_4 fanout4223 (.X(net4223),
    .A(net4227));
 sg13g2_buf_4 fanout4224 (.X(net4224),
    .A(net4225));
 sg13g2_buf_4 fanout4225 (.X(net4225),
    .A(net4226));
 sg13g2_buf_8 fanout4226 (.A(net4227),
    .X(net4226));
 sg13g2_buf_8 fanout4227 (.A(net4260),
    .X(net4227));
 sg13g2_buf_4 fanout4228 (.X(net4228),
    .A(net4231));
 sg13g2_buf_4 fanout4229 (.X(net4229),
    .A(net4231));
 sg13g2_buf_4 fanout4230 (.X(net4230),
    .A(net4231));
 sg13g2_buf_4 fanout4231 (.X(net4231),
    .A(net4236));
 sg13g2_buf_4 fanout4232 (.X(net4232),
    .A(net4233));
 sg13g2_buf_4 fanout4233 (.X(net4233),
    .A(net4236));
 sg13g2_buf_4 fanout4234 (.X(net4234),
    .A(net4236));
 sg13g2_buf_4 fanout4235 (.X(net4235),
    .A(net4236));
 sg13g2_buf_1 fanout4236 (.A(net4260),
    .X(net4236));
 sg13g2_buf_4 fanout4237 (.X(net4237),
    .A(net4238));
 sg13g2_buf_4 fanout4238 (.X(net4238),
    .A(net4239));
 sg13g2_buf_4 fanout4239 (.X(net4239),
    .A(net4241));
 sg13g2_buf_4 fanout4240 (.X(net4240),
    .A(net4241));
 sg13g2_buf_2 fanout4241 (.A(net4259),
    .X(net4241));
 sg13g2_buf_4 fanout4242 (.X(net4242),
    .A(net4243));
 sg13g2_buf_4 fanout4243 (.X(net4243),
    .A(net4259));
 sg13g2_buf_4 fanout4244 (.X(net4244),
    .A(net4245));
 sg13g2_buf_4 fanout4245 (.X(net4245),
    .A(net4259));
 sg13g2_buf_4 fanout4246 (.X(net4246),
    .A(net4247));
 sg13g2_buf_4 fanout4247 (.X(net4247),
    .A(net4251));
 sg13g2_buf_4 fanout4248 (.X(net4248),
    .A(net4249));
 sg13g2_buf_4 fanout4249 (.X(net4249),
    .A(net4251));
 sg13g2_buf_4 fanout4250 (.X(net4250),
    .A(net4251));
 sg13g2_buf_4 fanout4251 (.X(net4251),
    .A(net4259));
 sg13g2_buf_4 fanout4252 (.X(net4252),
    .A(net4253));
 sg13g2_buf_2 fanout4253 (.A(net4254),
    .X(net4253));
 sg13g2_buf_4 fanout4254 (.X(net4254),
    .A(net4258));
 sg13g2_buf_4 fanout4255 (.X(net4255),
    .A(net4256));
 sg13g2_buf_2 fanout4256 (.A(net4257),
    .X(net4256));
 sg13g2_buf_4 fanout4257 (.X(net4257),
    .A(net4258));
 sg13g2_buf_2 fanout4258 (.A(net4259),
    .X(net4258));
 sg13g2_buf_8 fanout4259 (.A(net4260),
    .X(net4259));
 sg13g2_buf_16 fanout4260 (.X(net4260),
    .A(net4261));
 sg13g2_buf_8 fanout4261 (.A(\spiking_network_top_uut.sys_clk_reset_synchr ),
    .X(net4261));
 sg13g2_buf_2 fanout4262 (.A(net4263),
    .X(net4262));
 sg13g2_buf_2 fanout4263 (.A(\spiking_network_top_uut.spi_inst.memory_inst.addr_reg_out[1] ),
    .X(net4263));
 sg13g2_buf_2 fanout4264 (.A(net4265),
    .X(net4264));
 sg13g2_buf_1 fanout4265 (.A(\spiking_network_top_uut.spi_inst.memory_inst.addr_reg_out[0] ),
    .X(net4265));
 sg13g2_buf_4 fanout4266 (.X(net4266),
    .A(net4267));
 sg13g2_buf_8 fanout4267 (.A(\spiking_network_top_uut.all_data_out[1] ),
    .X(net4267));
 sg13g2_buf_8 fanout4268 (.A(\spiking_network_top_uut.all_data_out[0] ),
    .X(net4268));
 sg13g2_buf_8 fanout4269 (.A(net4271),
    .X(net4269));
 sg13g2_buf_4 fanout4270 (.X(net4270),
    .A(net4271));
 sg13g2_buf_8 fanout4271 (.A(net4272),
    .X(net4271));
 sg13g2_buf_8 fanout4272 (.A(\spiking_network_top_uut.all_data_out[12] ),
    .X(net4272));
 sg13g2_buf_8 fanout4273 (.A(net4275),
    .X(net4273));
 sg13g2_buf_4 fanout4274 (.X(net4274),
    .A(net4275));
 sg13g2_buf_16 fanout4275 (.X(net4275),
    .A(\spiking_network_top_uut.all_data_out[11] ));
 sg13g2_buf_8 fanout4276 (.A(net4278),
    .X(net4276));
 sg13g2_buf_4 fanout4277 (.X(net4277),
    .A(net4278));
 sg13g2_buf_8 fanout4278 (.A(net4279),
    .X(net4278));
 sg13g2_buf_8 fanout4279 (.A(\spiking_network_top_uut.all_data_out[10] ),
    .X(net4279));
 sg13g2_buf_8 fanout4280 (.A(net4282),
    .X(net4280));
 sg13g2_buf_4 fanout4281 (.X(net4281),
    .A(net4282));
 sg13g2_buf_16 fanout4282 (.X(net4282),
    .A(\spiking_network_top_uut.all_data_out[9] ));
 sg13g2_buf_8 fanout4283 (.A(net4285),
    .X(net4283));
 sg13g2_buf_4 fanout4284 (.X(net4284),
    .A(net4285));
 sg13g2_buf_8 fanout4285 (.A(net4286),
    .X(net4285));
 sg13g2_buf_8 fanout4286 (.A(\spiking_network_top_uut.all_data_out[8] ),
    .X(net4286));
 sg13g2_buf_4 fanout4287 (.X(net4287),
    .A(net4288));
 sg13g2_buf_4 fanout4288 (.X(net4288),
    .A(net4291));
 sg13g2_buf_4 fanout4289 (.X(net4289),
    .A(net4291));
 sg13g2_buf_2 fanout4290 (.A(net4291),
    .X(net4290));
 sg13g2_buf_4 fanout4291 (.X(net4291),
    .A(net4292));
 sg13g2_buf_8 fanout4292 (.A(\spiking_network_top_uut.all_data_out[20] ),
    .X(net4292));
 sg13g2_buf_8 fanout4293 (.A(net4294),
    .X(net4293));
 sg13g2_buf_8 fanout4294 (.A(net4297),
    .X(net4294));
 sg13g2_buf_4 fanout4295 (.X(net4295),
    .A(net4297));
 sg13g2_buf_2 fanout4296 (.A(net4297),
    .X(net4296));
 sg13g2_buf_4 fanout4297 (.X(net4297),
    .A(net4298));
 sg13g2_buf_8 fanout4298 (.A(\spiking_network_top_uut.all_data_out[19] ),
    .X(net4298));
 sg13g2_buf_4 fanout4299 (.X(net4299),
    .A(net4302));
 sg13g2_buf_2 fanout4300 (.A(net4302),
    .X(net4300));
 sg13g2_buf_4 fanout4301 (.X(net4301),
    .A(net4302));
 sg13g2_buf_4 fanout4302 (.X(net4302),
    .A(net4304));
 sg13g2_buf_4 fanout4303 (.X(net4303),
    .A(net4304));
 sg13g2_buf_2 fanout4304 (.A(net4305),
    .X(net4304));
 sg13g2_buf_8 fanout4305 (.A(\spiking_network_top_uut.all_data_out[18] ),
    .X(net4305));
 sg13g2_buf_4 fanout4306 (.X(net4306),
    .A(net4308));
 sg13g2_buf_4 fanout4307 (.X(net4307),
    .A(net4308));
 sg13g2_buf_4 fanout4308 (.X(net4308),
    .A(net4309));
 sg13g2_buf_4 fanout4309 (.X(net4309),
    .A(net4310));
 sg13g2_buf_4 fanout4310 (.X(net4310),
    .A(\spiking_network_top_uut.all_data_out[17] ));
 sg13g2_buf_4 fanout4311 (.X(net4311),
    .A(net4314));
 sg13g2_buf_2 fanout4312 (.A(net4314),
    .X(net4312));
 sg13g2_buf_4 fanout4313 (.X(net4313),
    .A(net4314));
 sg13g2_buf_4 fanout4314 (.X(net4314),
    .A(net4315));
 sg13g2_buf_4 fanout4315 (.X(net4315),
    .A(net4316));
 sg13g2_buf_8 fanout4316 (.A(\spiking_network_top_uut.all_data_out[16] ),
    .X(net4316));
 sg13g2_buf_4 fanout4317 (.X(net4317),
    .A(\spiking_network_top_uut.spi_inst.memory_inst.write_enable ));
 sg13g2_buf_4 fanout4318 (.X(net4318),
    .A(\spiking_network_top_uut.spi_inst.SPI_instruction_reg_en ));
 sg13g2_buf_4 fanout4319 (.X(net4319),
    .A(net4324));
 sg13g2_buf_4 fanout4320 (.X(net4320),
    .A(net4321));
 sg13g2_buf_4 fanout4321 (.X(net4321),
    .A(net4324));
 sg13g2_buf_8 fanout4322 (.A(net4324),
    .X(net4322));
 sg13g2_buf_4 fanout4323 (.X(net4323),
    .A(net4324));
 sg13g2_buf_8 fanout4324 (.A(net4338),
    .X(net4324));
 sg13g2_buf_4 fanout4325 (.X(net4325),
    .A(net4328));
 sg13g2_buf_4 fanout4326 (.X(net4326),
    .A(net4327));
 sg13g2_buf_4 fanout4327 (.X(net4327),
    .A(net4328));
 sg13g2_buf_2 fanout4328 (.A(net4338),
    .X(net4328));
 sg13g2_buf_4 fanout4329 (.X(net4329),
    .A(net4331));
 sg13g2_buf_2 fanout4330 (.A(net4331),
    .X(net4330));
 sg13g2_buf_8 fanout4331 (.A(net4338),
    .X(net4331));
 sg13g2_buf_4 fanout4332 (.X(net4332),
    .A(net4337));
 sg13g2_buf_1 fanout4333 (.A(net4337),
    .X(net4333));
 sg13g2_buf_4 fanout4334 (.X(net4334),
    .A(net4337));
 sg13g2_buf_4 fanout4335 (.X(net4335),
    .A(net4336));
 sg13g2_buf_4 fanout4336 (.X(net4336),
    .A(net4337));
 sg13g2_buf_2 fanout4337 (.A(net4338),
    .X(net4337));
 sg13g2_buf_8 fanout4338 (.A(\spiking_network_top_uut.spi_inst.SPI_instruction_reg_in[7] ),
    .X(net4338));
 sg13g2_buf_8 fanout4339 (.A(net4340),
    .X(net4339));
 sg13g2_buf_8 fanout4340 (.A(net4346),
    .X(net4340));
 sg13g2_buf_4 fanout4341 (.X(net4341),
    .A(net4342));
 sg13g2_buf_8 fanout4342 (.A(net4345),
    .X(net4342));
 sg13g2_buf_8 fanout4343 (.A(net4344),
    .X(net4343));
 sg13g2_buf_8 fanout4344 (.A(net4345),
    .X(net4344));
 sg13g2_buf_4 fanout4345 (.X(net4345),
    .A(net4346));
 sg13g2_buf_4 fanout4346 (.X(net4346),
    .A(\spiking_network_top_uut.spi_inst.SPI_instruction_reg_in[6] ));
 sg13g2_buf_4 fanout4347 (.X(net4347),
    .A(net4350));
 sg13g2_buf_2 fanout4348 (.A(net4350),
    .X(net4348));
 sg13g2_buf_4 fanout4349 (.X(net4349),
    .A(net4350));
 sg13g2_buf_4 fanout4350 (.X(net4350),
    .A(net4359));
 sg13g2_buf_4 fanout4351 (.X(net4351),
    .A(net4359));
 sg13g2_buf_2 fanout4352 (.A(net4359),
    .X(net4352));
 sg13g2_buf_4 fanout4353 (.X(net4353),
    .A(net4359));
 sg13g2_buf_4 fanout4354 (.X(net4354),
    .A(net4359));
 sg13g2_buf_4 fanout4355 (.X(net4355),
    .A(net4357));
 sg13g2_buf_1 fanout4356 (.A(net4357),
    .X(net4356));
 sg13g2_buf_2 fanout4357 (.A(net4358),
    .X(net4357));
 sg13g2_buf_4 fanout4358 (.X(net4358),
    .A(net4359));
 sg13g2_buf_8 fanout4359 (.A(\spiking_network_top_uut.spi_inst.SPI_instruction_reg_in[6] ),
    .X(net4359));
 sg13g2_buf_4 fanout4360 (.X(net4360),
    .A(net4363));
 sg13g2_buf_8 fanout4361 (.A(net4363),
    .X(net4361));
 sg13g2_buf_2 fanout4362 (.A(net4363),
    .X(net4362));
 sg13g2_buf_4 fanout4363 (.X(net4363),
    .A(net4368));
 sg13g2_buf_4 fanout4364 (.X(net4364),
    .A(net4365));
 sg13g2_buf_4 fanout4365 (.X(net4365),
    .A(net4368));
 sg13g2_buf_8 fanout4366 (.A(net4368),
    .X(net4366));
 sg13g2_buf_4 fanout4367 (.X(net4367),
    .A(net4368));
 sg13g2_buf_4 fanout4368 (.X(net4368),
    .A(\spiking_network_top_uut.spi_inst.SPI_instruction_reg_in[5] ));
 sg13g2_buf_4 fanout4369 (.X(net4369),
    .A(net4370));
 sg13g2_buf_8 fanout4370 (.A(net4374),
    .X(net4370));
 sg13g2_buf_2 fanout4371 (.A(net4374),
    .X(net4371));
 sg13g2_buf_4 fanout4372 (.X(net4372),
    .A(net4373));
 sg13g2_buf_4 fanout4373 (.X(net4373),
    .A(net4374));
 sg13g2_buf_4 fanout4374 (.X(net4374),
    .A(net4379));
 sg13g2_buf_4 fanout4375 (.X(net4375),
    .A(net4376));
 sg13g2_buf_4 fanout4376 (.X(net4376),
    .A(net4377));
 sg13g2_buf_4 fanout4377 (.X(net4377),
    .A(net4379));
 sg13g2_buf_4 fanout4378 (.X(net4378),
    .A(net4379));
 sg13g2_buf_8 fanout4379 (.A(\spiking_network_top_uut.spi_inst.SPI_instruction_reg_in[5] ),
    .X(net4379));
 sg13g2_buf_4 fanout4380 (.X(net4380),
    .A(net4381));
 sg13g2_buf_8 fanout4381 (.A(net4387),
    .X(net4381));
 sg13g2_buf_4 fanout4382 (.X(net4382),
    .A(net4383));
 sg13g2_buf_2 fanout4383 (.A(net4384),
    .X(net4383));
 sg13g2_buf_4 fanout4384 (.X(net4384),
    .A(net4387));
 sg13g2_buf_4 fanout4385 (.X(net4385),
    .A(net4386));
 sg13g2_buf_4 fanout4386 (.X(net4386),
    .A(net4387));
 sg13g2_buf_8 fanout4387 (.A(\spiking_network_top_uut.spi_inst.SPI_instruction_reg_in[4] ),
    .X(net4387));
 sg13g2_buf_4 fanout4388 (.X(net4388),
    .A(net4391));
 sg13g2_buf_2 fanout4389 (.A(net4391),
    .X(net4389));
 sg13g2_buf_4 fanout4390 (.X(net4390),
    .A(net4391));
 sg13g2_buf_4 fanout4391 (.X(net4391),
    .A(net4400));
 sg13g2_buf_8 fanout4392 (.A(net4400),
    .X(net4392));
 sg13g2_buf_2 fanout4393 (.A(net4400),
    .X(net4393));
 sg13g2_buf_4 fanout4394 (.X(net4394),
    .A(net4399));
 sg13g2_buf_2 fanout4395 (.A(net4399),
    .X(net4395));
 sg13g2_buf_4 fanout4396 (.X(net4396),
    .A(net4397));
 sg13g2_buf_2 fanout4397 (.A(net4398),
    .X(net4397));
 sg13g2_buf_4 fanout4398 (.X(net4398),
    .A(net4399));
 sg13g2_buf_2 fanout4399 (.A(net4400),
    .X(net4399));
 sg13g2_buf_4 fanout4400 (.X(net4400),
    .A(\spiking_network_top_uut.spi_inst.SPI_instruction_reg_in[4] ));
 sg13g2_buf_4 fanout4401 (.X(net4401),
    .A(net4421));
 sg13g2_buf_4 fanout4402 (.X(net4402),
    .A(net4421));
 sg13g2_buf_4 fanout4403 (.X(net4403),
    .A(net4407));
 sg13g2_buf_2 fanout4404 (.A(net4407),
    .X(net4404));
 sg13g2_buf_4 fanout4405 (.X(net4405),
    .A(net4407));
 sg13g2_buf_4 fanout4406 (.X(net4406),
    .A(net4407));
 sg13g2_buf_8 fanout4407 (.A(net4421),
    .X(net4407));
 sg13g2_buf_8 fanout4408 (.A(net4412),
    .X(net4408));
 sg13g2_buf_4 fanout4409 (.X(net4409),
    .A(net4412));
 sg13g2_buf_4 fanout4410 (.X(net4410),
    .A(net4411));
 sg13g2_buf_8 fanout4411 (.A(net4412),
    .X(net4411));
 sg13g2_buf_4 fanout4412 (.X(net4412),
    .A(net4421));
 sg13g2_buf_4 fanout4413 (.X(net4413),
    .A(net4416));
 sg13g2_buf_4 fanout4414 (.X(net4414),
    .A(net4416));
 sg13g2_buf_2 fanout4415 (.A(net4416),
    .X(net4415));
 sg13g2_buf_2 fanout4416 (.A(net4421),
    .X(net4416));
 sg13g2_buf_4 fanout4417 (.X(net4417),
    .A(net4418));
 sg13g2_buf_2 fanout4418 (.A(net4420),
    .X(net4418));
 sg13g2_buf_4 fanout4419 (.X(net4419),
    .A(net4420));
 sg13g2_buf_4 fanout4420 (.X(net4420),
    .A(net4421));
 sg13g2_buf_8 fanout4421 (.A(\spiking_network_top_uut.spi_inst.SPI_instruction_reg_in[3] ),
    .X(net4421));
 sg13g2_buf_4 fanout4422 (.X(net4422),
    .A(net4423));
 sg13g2_buf_8 fanout4423 (.A(\spiking_network_top_uut.spi_inst.SPI_instruction_reg_in[2] ),
    .X(net4423));
 sg13g2_buf_4 fanout4424 (.X(net4424),
    .A(net4425));
 sg13g2_buf_8 fanout4425 (.A(net4429),
    .X(net4425));
 sg13g2_buf_4 fanout4426 (.X(net4426),
    .A(net4428));
 sg13g2_buf_4 fanout4427 (.X(net4427),
    .A(net4428));
 sg13g2_buf_8 fanout4428 (.A(net4429),
    .X(net4428));
 sg13g2_buf_2 fanout4429 (.A(\spiking_network_top_uut.spi_inst.SPI_instruction_reg_in[2] ),
    .X(net4429));
 sg13g2_buf_4 fanout4430 (.X(net4430),
    .A(net4440));
 sg13g2_buf_4 fanout4431 (.X(net4431),
    .A(net4440));
 sg13g2_buf_4 fanout4432 (.X(net4432),
    .A(net4433));
 sg13g2_buf_8 fanout4433 (.A(net4440),
    .X(net4433));
 sg13g2_buf_4 fanout4434 (.X(net4434),
    .A(net4435));
 sg13g2_buf_8 fanout4435 (.A(net4439),
    .X(net4435));
 sg13g2_buf_4 fanout4436 (.X(net4436),
    .A(net4438));
 sg13g2_buf_4 fanout4437 (.X(net4437),
    .A(net4438));
 sg13g2_buf_8 fanout4438 (.A(net4439),
    .X(net4438));
 sg13g2_buf_4 fanout4439 (.X(net4439),
    .A(net4440));
 sg13g2_buf_8 fanout4440 (.A(\spiking_network_top_uut.spi_inst.SPI_instruction_reg_in[2] ),
    .X(net4440));
 sg13g2_buf_8 fanout4441 (.A(net4442),
    .X(net4441));
 sg13g2_buf_4 fanout4442 (.X(net4442),
    .A(net4449));
 sg13g2_buf_4 fanout4443 (.X(net4443),
    .A(net4444));
 sg13g2_buf_8 fanout4444 (.A(net4449),
    .X(net4444));
 sg13g2_buf_4 fanout4445 (.X(net4445),
    .A(net4448));
 sg13g2_buf_4 fanout4446 (.X(net4446),
    .A(net4448));
 sg13g2_buf_4 fanout4447 (.X(net4447),
    .A(net4448));
 sg13g2_buf_4 fanout4448 (.X(net4448),
    .A(net4449));
 sg13g2_buf_4 fanout4449 (.X(net4449),
    .A(net4461));
 sg13g2_buf_8 fanout4450 (.A(net4454),
    .X(net4450));
 sg13g2_buf_4 fanout4451 (.X(net4451),
    .A(net4454));
 sg13g2_buf_4 fanout4452 (.X(net4452),
    .A(net4454));
 sg13g2_buf_2 fanout4453 (.A(net4454),
    .X(net4453));
 sg13g2_buf_4 fanout4454 (.X(net4454),
    .A(net4461));
 sg13g2_buf_4 fanout4455 (.X(net4455),
    .A(net4456));
 sg13g2_buf_8 fanout4456 (.A(net4461),
    .X(net4456));
 sg13g2_buf_4 fanout4457 (.X(net4457),
    .A(net4460));
 sg13g2_buf_4 fanout4458 (.X(net4458),
    .A(net4460));
 sg13g2_buf_2 fanout4459 (.A(net4460),
    .X(net4459));
 sg13g2_buf_4 fanout4460 (.X(net4460),
    .A(net4461));
 sg13g2_buf_8 fanout4461 (.A(\spiking_network_top_uut.spi_inst.SPI_instruction_reg_in[1] ),
    .X(net4461));
 sg13g2_buf_8 fanout4462 (.A(net4482),
    .X(net4462));
 sg13g2_buf_2 fanout4463 (.A(net4482),
    .X(net4463));
 sg13g2_buf_4 fanout4464 (.X(net4464),
    .A(net4466));
 sg13g2_buf_2 fanout4465 (.A(net4466),
    .X(net4465));
 sg13g2_buf_8 fanout4466 (.A(net4470),
    .X(net4466));
 sg13g2_buf_4 fanout4467 (.X(net4467),
    .A(net4468));
 sg13g2_buf_4 fanout4468 (.X(net4468),
    .A(net4469));
 sg13g2_buf_4 fanout4469 (.X(net4469),
    .A(net4470));
 sg13g2_buf_4 fanout4470 (.X(net4470),
    .A(net4482));
 sg13g2_buf_4 fanout4471 (.X(net4471),
    .A(net4481));
 sg13g2_buf_2 fanout4472 (.A(net4481),
    .X(net4472));
 sg13g2_buf_4 fanout4473 (.X(net4473),
    .A(net4474));
 sg13g2_buf_4 fanout4474 (.X(net4474),
    .A(net4481));
 sg13g2_buf_4 fanout4475 (.X(net4475),
    .A(net4476));
 sg13g2_buf_8 fanout4476 (.A(net4481),
    .X(net4476));
 sg13g2_buf_4 fanout4477 (.X(net4477),
    .A(net4480));
 sg13g2_buf_4 fanout4478 (.X(net4478),
    .A(net4480));
 sg13g2_buf_2 fanout4479 (.A(net4480),
    .X(net4479));
 sg13g2_buf_2 fanout4480 (.A(net4481),
    .X(net4480));
 sg13g2_buf_8 fanout4481 (.A(net4482),
    .X(net4481));
 sg13g2_buf_8 fanout4482 (.A(\spiking_network_top_uut.spi_inst.SPI_instruction_reg_in[0] ),
    .X(net4482));
 sg13g2_buf_2 fanout4483 (.A(\spiking_network_top_uut.spi_inst.LSB_Address_reg[1] ),
    .X(net4483));
 sg13g2_buf_2 fanout4484 (.A(\spiking_network_top_uut.spi_inst.LSB_Address_reg[0] ),
    .X(net4484));
 sg13g2_buf_8 fanout4485 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.din ),
    .X(net4485));
 sg13g2_buf_8 fanout4486 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.din ),
    .X(net4486));
 sg13g2_buf_4 fanout4487 (.X(net4487),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.din ));
 sg13g2_buf_8 fanout4488 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.din ),
    .X(net4488));
 sg13g2_buf_4 fanout4489 (.X(net4489),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.din ));
 sg13g2_buf_8 fanout4490 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.din ),
    .X(net4490));
 sg13g2_buf_8 fanout4491 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.din ),
    .X(net4491));
 sg13g2_buf_8 fanout4492 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.din ),
    .X(net4492));
 sg13g2_buf_2 fanout4493 (.A(net4509),
    .X(net4493));
 sg13g2_buf_2 fanout4494 (.A(net4509),
    .X(net4494));
 sg13g2_buf_4 fanout4495 (.X(net4495),
    .A(net4499));
 sg13g2_buf_2 fanout4496 (.A(net4499),
    .X(net4496));
 sg13g2_buf_2 fanout4497 (.A(net4498),
    .X(net4497));
 sg13g2_buf_1 fanout4498 (.A(net4499),
    .X(net4498));
 sg13g2_buf_2 fanout4499 (.A(net4500),
    .X(net4499));
 sg13g2_buf_4 fanout4500 (.X(net4500),
    .A(net4509));
 sg13g2_buf_2 fanout4501 (.A(net4502),
    .X(net4501));
 sg13g2_buf_2 fanout4502 (.A(net4505),
    .X(net4502));
 sg13g2_buf_2 fanout4503 (.A(net4505),
    .X(net4503));
 sg13g2_buf_1 fanout4504 (.A(net4505),
    .X(net4504));
 sg13g2_buf_2 fanout4505 (.A(net4508),
    .X(net4505));
 sg13g2_buf_4 fanout4506 (.X(net4506),
    .A(net4508));
 sg13g2_buf_2 fanout4507 (.A(net4508),
    .X(net4507));
 sg13g2_buf_4 fanout4508 (.X(net4508),
    .A(net4509));
 sg13g2_buf_4 fanout4509 (.X(net4509),
    .A(\spiking_network_top_uut.clk_div_inst.clk_out ));
 sg13g2_buf_2 fanout4510 (.A(net4528),
    .X(net4510));
 sg13g2_buf_2 fanout4511 (.A(net4513),
    .X(net4511));
 sg13g2_buf_4 fanout4512 (.X(net4512),
    .A(net4513));
 sg13g2_buf_4 fanout4513 (.X(net4513),
    .A(net4528));
 sg13g2_buf_2 fanout4514 (.A(net4527),
    .X(net4514));
 sg13g2_buf_2 fanout4515 (.A(net4527),
    .X(net4515));
 sg13g2_buf_4 fanout4516 (.X(net4516),
    .A(net4519));
 sg13g2_buf_4 fanout4517 (.X(net4517),
    .A(net4519));
 sg13g2_buf_1 fanout4518 (.A(net4519),
    .X(net4518));
 sg13g2_buf_4 fanout4519 (.X(net4519),
    .A(net4527));
 sg13g2_buf_2 fanout4520 (.A(net4526),
    .X(net4520));
 sg13g2_buf_1 fanout4521 (.A(net4526),
    .X(net4521));
 sg13g2_buf_2 fanout4522 (.A(net4526),
    .X(net4522));
 sg13g2_buf_4 fanout4523 (.X(net4523),
    .A(net4525));
 sg13g2_buf_4 fanout4524 (.X(net4524),
    .A(net4526));
 sg13g2_buf_2 fanout4525 (.A(net4526),
    .X(net4525));
 sg13g2_buf_8 fanout4526 (.A(net4527),
    .X(net4526));
 sg13g2_buf_4 fanout4527 (.X(net4527),
    .A(net4528));
 sg13g2_buf_8 fanout4528 (.A(\spiking_network_top_uut.clk_div_inst.clk_out ),
    .X(net4528));
 sg13g2_buf_8 fanout4529 (.A(net4532),
    .X(net4529));
 sg13g2_buf_2 fanout4530 (.A(net4532),
    .X(net4530));
 sg13g2_buf_8 fanout4531 (.A(net4532),
    .X(net4531));
 sg13g2_buf_4 fanout4532 (.X(net4532),
    .A(net4533));
 sg13g2_buf_4 fanout4533 (.X(net4533),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.enable_LYR_2 ));
 sg13g2_buf_4 fanout4534 (.X(net4534),
    .A(net4537));
 sg13g2_buf_4 fanout4535 (.X(net4535),
    .A(net4536));
 sg13g2_buf_2 fanout4536 (.A(net4537),
    .X(net4536));
 sg13g2_buf_4 fanout4537 (.X(net4537),
    .A(net4542));
 sg13g2_buf_2 fanout4538 (.A(net4539),
    .X(net4538));
 sg13g2_buf_2 fanout4539 (.A(net4542),
    .X(net4539));
 sg13g2_buf_2 fanout4540 (.A(net4541),
    .X(net4540));
 sg13g2_buf_4 fanout4541 (.X(net4541),
    .A(net4542));
 sg13g2_buf_2 fanout4542 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.enable_LYR_2 ),
    .X(net4542));
 sg13g2_buf_4 fanout4543 (.X(net4543),
    .A(net4544));
 sg13g2_buf_4 fanout4544 (.X(net4544),
    .A(net4572));
 sg13g2_buf_2 fanout4545 (.A(net4547),
    .X(net4545));
 sg13g2_buf_4 fanout4546 (.X(net4546),
    .A(net4547));
 sg13g2_buf_2 fanout4547 (.A(net4548),
    .X(net4547));
 sg13g2_buf_2 fanout4548 (.A(net4572),
    .X(net4548));
 sg13g2_buf_4 fanout4549 (.X(net4549),
    .A(net4553));
 sg13g2_buf_4 fanout4550 (.X(net4550),
    .A(net4551));
 sg13g2_buf_2 fanout4551 (.A(net4552),
    .X(net4551));
 sg13g2_buf_2 fanout4552 (.A(net4553),
    .X(net4552));
 sg13g2_buf_2 fanout4553 (.A(net4572),
    .X(net4553));
 sg13g2_buf_4 fanout4554 (.X(net4554),
    .A(net4555));
 sg13g2_buf_4 fanout4555 (.X(net4555),
    .A(net4556));
 sg13g2_buf_4 fanout4556 (.X(net4556),
    .A(net4557));
 sg13g2_buf_4 fanout4557 (.X(net4557),
    .A(net4571));
 sg13g2_buf_2 fanout4558 (.A(net4560),
    .X(net4558));
 sg13g2_buf_1 fanout4559 (.A(net4560),
    .X(net4559));
 sg13g2_buf_2 fanout4560 (.A(net4565),
    .X(net4560));
 sg13g2_buf_4 fanout4561 (.X(net4561),
    .A(net4565));
 sg13g2_buf_4 fanout4562 (.X(net4562),
    .A(net4563));
 sg13g2_buf_4 fanout4563 (.X(net4563),
    .A(net4564));
 sg13g2_buf_4 fanout4564 (.X(net4564),
    .A(net4565));
 sg13g2_buf_4 fanout4565 (.X(net4565),
    .A(net4570));
 sg13g2_buf_4 fanout4566 (.X(net4566),
    .A(net4568));
 sg13g2_buf_2 fanout4567 (.A(net4568),
    .X(net4567));
 sg13g2_buf_2 fanout4568 (.A(net4570),
    .X(net4568));
 sg13g2_buf_4 fanout4569 (.X(net4569),
    .A(net4570));
 sg13g2_buf_2 fanout4570 (.A(net4571),
    .X(net4570));
 sg13g2_buf_4 fanout4571 (.X(net4571),
    .A(net4572));
 sg13g2_buf_8 fanout4572 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.enable_LYR_2 ),
    .X(net4572));
 sg13g2_buf_4 fanout4573 (.X(net4573),
    .A(net4574));
 sg13g2_buf_4 fanout4574 (.X(net4574),
    .A(net456));
 sg13g2_buf_4 fanout4575 (.X(net4575),
    .A(net4576));
 sg13g2_buf_2 fanout4576 (.A(net4577),
    .X(net4576));
 sg13g2_buf_2 fanout4577 (.A(net553),
    .X(net4577));
 sg13g2_buf_4 fanout4578 (.X(net4578),
    .A(net4591));
 sg13g2_buf_2 fanout4579 (.A(net4591),
    .X(net4579));
 sg13g2_buf_4 fanout4580 (.X(net4580),
    .A(net4583));
 sg13g2_buf_2 fanout4581 (.A(net4582),
    .X(net4581));
 sg13g2_buf_4 fanout4582 (.X(net4582),
    .A(net4583));
 sg13g2_buf_2 fanout4583 (.A(net4591),
    .X(net4583));
 sg13g2_buf_4 fanout4584 (.X(net4584),
    .A(net4585));
 sg13g2_buf_2 fanout4585 (.A(net4587),
    .X(net4585));
 sg13g2_buf_4 fanout4586 (.X(net4586),
    .A(net4587));
 sg13g2_buf_2 fanout4587 (.A(net4590),
    .X(net4587));
 sg13g2_buf_4 fanout4588 (.X(net4588),
    .A(net4589));
 sg13g2_buf_2 fanout4589 (.A(net4590),
    .X(net4589));
 sg13g2_buf_2 fanout4590 (.A(net4591),
    .X(net4590));
 sg13g2_buf_2 fanout4591 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.enable_LYR_3 ),
    .X(net4591));
 sg13g2_buf_4 fanout4592 (.X(net4592),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.spike_out ));
 sg13g2_buf_4 fanout4593 (.X(net4593),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.spike_out ));
 sg13g2_buf_8 fanout4594 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.spike_out ),
    .X(net4594));
 sg13g2_buf_4 fanout4595 (.X(net4595),
    .A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.spike_out ));
 sg13g2_buf_8 fanout4596 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.spike_out ),
    .X(net4596));
 sg13g2_buf_8 fanout4597 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.spike_out ),
    .X(net4597));
 sg13g2_buf_8 fanout4598 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.spike_out ),
    .X(net4598));
 sg13g2_buf_8 fanout4599 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.spike_out ),
    .X(net4599));
 sg13g2_buf_4 fanout4600 (.X(net4600),
    .A(net4601));
 sg13g2_buf_2 fanout4601 (.A(net518),
    .X(net4601));
 sg13g2_buf_4 fanout4602 (.X(net4602),
    .A(net533));
 sg13g2_buf_4 fanout4603 (.X(net4603),
    .A(net4604));
 sg13g2_buf_4 fanout4604 (.X(net4604),
    .A(net4605));
 sg13g2_buf_4 fanout4605 (.X(net4605),
    .A(net4606));
 sg13g2_buf_8 fanout4606 (.A(\spiking_network_top_uut.SNN_en_sync ),
    .X(net4606));
 sg13g2_buf_2 fanout4607 (.A(net4608),
    .X(net4607));
 sg13g2_buf_2 fanout4608 (.A(net4612),
    .X(net4608));
 sg13g2_buf_4 fanout4609 (.X(net4609),
    .A(net4610));
 sg13g2_buf_2 fanout4610 (.A(net4611),
    .X(net4610));
 sg13g2_buf_2 fanout4611 (.A(net4612),
    .X(net4611));
 sg13g2_buf_2 fanout4612 (.A(\spiking_network_top_uut.SNN_en_sync ),
    .X(net4612));
 sg13g2_buf_4 fanout4613 (.X(net4613),
    .A(net4616));
 sg13g2_buf_4 fanout4614 (.X(net4614),
    .A(net4615));
 sg13g2_buf_2 fanout4615 (.A(net4616),
    .X(net4615));
 sg13g2_buf_2 fanout4616 (.A(net4646),
    .X(net4616));
 sg13g2_buf_2 fanout4617 (.A(net4618),
    .X(net4617));
 sg13g2_buf_2 fanout4618 (.A(net4619),
    .X(net4618));
 sg13g2_buf_2 fanout4619 (.A(net4620),
    .X(net4619));
 sg13g2_buf_4 fanout4620 (.X(net4620),
    .A(net4646));
 sg13g2_buf_4 fanout4621 (.X(net4621),
    .A(net4623));
 sg13g2_buf_2 fanout4622 (.A(net4623),
    .X(net4622));
 sg13g2_buf_2 fanout4623 (.A(net4624),
    .X(net4623));
 sg13g2_buf_4 fanout4624 (.X(net4624),
    .A(net4630));
 sg13g2_buf_4 fanout4625 (.X(net4625),
    .A(net4629));
 sg13g2_buf_4 fanout4626 (.X(net4626),
    .A(net4629));
 sg13g2_buf_4 fanout4627 (.X(net4627),
    .A(net4629));
 sg13g2_buf_4 fanout4628 (.X(net4628),
    .A(net4629));
 sg13g2_buf_2 fanout4629 (.A(net4630),
    .X(net4629));
 sg13g2_buf_2 fanout4630 (.A(net4645),
    .X(net4630));
 sg13g2_buf_4 fanout4631 (.X(net4631),
    .A(net4633));
 sg13g2_buf_4 fanout4632 (.X(net4632),
    .A(net4633));
 sg13g2_buf_4 fanout4633 (.X(net4633),
    .A(net4645));
 sg13g2_buf_4 fanout4634 (.X(net4634),
    .A(net4635));
 sg13g2_buf_4 fanout4635 (.X(net4635),
    .A(net4636));
 sg13g2_buf_4 fanout4636 (.X(net4636),
    .A(net4645));
 sg13g2_buf_4 fanout4637 (.X(net4637),
    .A(net4638));
 sg13g2_buf_2 fanout4638 (.A(net4639),
    .X(net4638));
 sg13g2_buf_4 fanout4639 (.X(net4639),
    .A(net4644));
 sg13g2_buf_4 fanout4640 (.X(net4640),
    .A(net4641));
 sg13g2_buf_2 fanout4641 (.A(net4644),
    .X(net4641));
 sg13g2_buf_2 fanout4642 (.A(net4643),
    .X(net4642));
 sg13g2_buf_2 fanout4643 (.A(net4644),
    .X(net4643));
 sg13g2_buf_2 fanout4644 (.A(net4645),
    .X(net4644));
 sg13g2_buf_4 fanout4645 (.X(net4645),
    .A(net4646));
 sg13g2_buf_4 fanout4646 (.X(net4646),
    .A(\spiking_network_top_uut.SNN_en_sync ));
 sg13g2_buf_4 fanout4647 (.X(net4647),
    .A(net4648));
 sg13g2_buf_8 fanout4648 (.A(net4709),
    .X(net4648));
 sg13g2_buf_2 fanout4649 (.A(net4653),
    .X(net4649));
 sg13g2_buf_2 fanout4650 (.A(net4653),
    .X(net4650));
 sg13g2_buf_2 fanout4651 (.A(net4653),
    .X(net4651));
 sg13g2_buf_2 fanout4652 (.A(net4653),
    .X(net4652));
 sg13g2_buf_2 fanout4653 (.A(net4659),
    .X(net4653));
 sg13g2_buf_2 fanout4654 (.A(net4658),
    .X(net4654));
 sg13g2_buf_1 fanout4655 (.A(net4658),
    .X(net4655));
 sg13g2_buf_2 fanout4656 (.A(net4657),
    .X(net4656));
 sg13g2_buf_2 fanout4657 (.A(net4658),
    .X(net4657));
 sg13g2_buf_2 fanout4658 (.A(net4659),
    .X(net4658));
 sg13g2_buf_4 fanout4659 (.X(net4659),
    .A(net4709));
 sg13g2_buf_2 fanout4660 (.A(net4663),
    .X(net4660));
 sg13g2_buf_2 fanout4661 (.A(net4662),
    .X(net4661));
 sg13g2_buf_2 fanout4662 (.A(net4663),
    .X(net4662));
 sg13g2_buf_2 fanout4663 (.A(net4677),
    .X(net4663));
 sg13g2_buf_2 fanout4664 (.A(net4665),
    .X(net4664));
 sg13g2_buf_2 fanout4665 (.A(net4670),
    .X(net4665));
 sg13g2_buf_4 fanout4666 (.X(net4666),
    .A(net4667));
 sg13g2_buf_4 fanout4667 (.X(net4667),
    .A(net4669));
 sg13g2_buf_4 fanout4668 (.X(net4668),
    .A(net4669));
 sg13g2_buf_2 fanout4669 (.A(net4670),
    .X(net4669));
 sg13g2_buf_2 fanout4670 (.A(net4677),
    .X(net4670));
 sg13g2_buf_2 fanout4671 (.A(net4677),
    .X(net4671));
 sg13g2_buf_2 fanout4672 (.A(net4677),
    .X(net4672));
 sg13g2_buf_4 fanout4673 (.X(net4673),
    .A(net4675));
 sg13g2_buf_2 fanout4674 (.A(net4675),
    .X(net4674));
 sg13g2_buf_1 fanout4675 (.A(net4676),
    .X(net4675));
 sg13g2_buf_4 fanout4676 (.X(net4676),
    .A(net4677));
 sg13g2_buf_4 fanout4677 (.X(net4677),
    .A(net4709));
 sg13g2_buf_2 fanout4678 (.A(net4680),
    .X(net4678));
 sg13g2_buf_2 fanout4679 (.A(net4680),
    .X(net4679));
 sg13g2_buf_2 fanout4680 (.A(net4691),
    .X(net4680));
 sg13g2_buf_4 fanout4681 (.X(net4681),
    .A(net4684));
 sg13g2_buf_1 fanout4682 (.A(net4684),
    .X(net4682));
 sg13g2_buf_2 fanout4683 (.A(net4684),
    .X(net4683));
 sg13g2_buf_2 fanout4684 (.A(net4691),
    .X(net4684));
 sg13g2_buf_2 fanout4685 (.A(net4686),
    .X(net4685));
 sg13g2_buf_2 fanout4686 (.A(net4690),
    .X(net4686));
 sg13g2_buf_2 fanout4687 (.A(net4690),
    .X(net4687));
 sg13g2_buf_2 fanout4688 (.A(net4690),
    .X(net4688));
 sg13g2_buf_2 fanout4689 (.A(net4690),
    .X(net4689));
 sg13g2_buf_2 fanout4690 (.A(net4691),
    .X(net4690));
 sg13g2_buf_2 fanout4691 (.A(net4709),
    .X(net4691));
 sg13g2_buf_2 fanout4692 (.A(net4694),
    .X(net4692));
 sg13g2_buf_2 fanout4693 (.A(net4694),
    .X(net4693));
 sg13g2_buf_2 fanout4694 (.A(net4708),
    .X(net4694));
 sg13g2_buf_2 fanout4695 (.A(net4696),
    .X(net4695));
 sg13g2_buf_2 fanout4696 (.A(net4697),
    .X(net4696));
 sg13g2_buf_2 fanout4697 (.A(net4708),
    .X(net4697));
 sg13g2_buf_2 fanout4698 (.A(net4702),
    .X(net4698));
 sg13g2_buf_2 fanout4699 (.A(net4702),
    .X(net4699));
 sg13g2_buf_2 fanout4700 (.A(net4702),
    .X(net4700));
 sg13g2_buf_2 fanout4701 (.A(net4702),
    .X(net4701));
 sg13g2_buf_2 fanout4702 (.A(net4708),
    .X(net4702));
 sg13g2_buf_2 fanout4703 (.A(net4707),
    .X(net4703));
 sg13g2_buf_2 fanout4704 (.A(net4705),
    .X(net4704));
 sg13g2_buf_1 fanout4705 (.A(net4706),
    .X(net4705));
 sg13g2_buf_2 fanout4706 (.A(net4707),
    .X(net4706));
 sg13g2_buf_2 fanout4707 (.A(net4708),
    .X(net4707));
 sg13g2_buf_2 fanout4708 (.A(net4709),
    .X(net4708));
 sg13g2_buf_8 fanout4709 (.A(uio_in[3]),
    .X(net4709));
 sg13g2_buf_2 fanout4710 (.A(net4711),
    .X(net4710));
 sg13g2_buf_2 fanout4711 (.A(net4722),
    .X(net4711));
 sg13g2_buf_2 fanout4712 (.A(net4714),
    .X(net4712));
 sg13g2_buf_2 fanout4713 (.A(net4714),
    .X(net4713));
 sg13g2_buf_2 fanout4714 (.A(net4722),
    .X(net4714));
 sg13g2_buf_2 fanout4715 (.A(net4721),
    .X(net4715));
 sg13g2_buf_2 fanout4716 (.A(net4721),
    .X(net4716));
 sg13g2_buf_2 fanout4717 (.A(net4718),
    .X(net4717));
 sg13g2_buf_2 fanout4718 (.A(net4721),
    .X(net4718));
 sg13g2_buf_2 fanout4719 (.A(net4720),
    .X(net4719));
 sg13g2_buf_4 fanout4720 (.X(net4720),
    .A(net4721));
 sg13g2_buf_4 fanout4721 (.X(net4721),
    .A(net4722));
 sg13g2_buf_2 fanout4722 (.A(net4764),
    .X(net4722));
 sg13g2_buf_2 fanout4723 (.A(net4724),
    .X(net4723));
 sg13g2_buf_2 fanout4724 (.A(net4726),
    .X(net4724));
 sg13g2_buf_4 fanout4725 (.X(net4725),
    .A(net4726));
 sg13g2_buf_2 fanout4726 (.A(net4738),
    .X(net4726));
 sg13g2_buf_2 fanout4727 (.A(net4731),
    .X(net4727));
 sg13g2_buf_2 fanout4728 (.A(net4731),
    .X(net4728));
 sg13g2_buf_2 fanout4729 (.A(net4731),
    .X(net4729));
 sg13g2_buf_2 fanout4730 (.A(net4731),
    .X(net4730));
 sg13g2_buf_1 fanout4731 (.A(net4738),
    .X(net4731));
 sg13g2_buf_4 fanout4732 (.X(net4732),
    .A(net4734));
 sg13g2_buf_4 fanout4733 (.X(net4733),
    .A(net4734));
 sg13g2_buf_2 fanout4734 (.A(net4738),
    .X(net4734));
 sg13g2_buf_2 fanout4735 (.A(net4737),
    .X(net4735));
 sg13g2_buf_2 fanout4736 (.A(net4737),
    .X(net4736));
 sg13g2_buf_2 fanout4737 (.A(net4738),
    .X(net4737));
 sg13g2_buf_4 fanout4738 (.X(net4738),
    .A(net4764));
 sg13g2_buf_2 fanout4739 (.A(net4741),
    .X(net4739));
 sg13g2_buf_2 fanout4740 (.A(net4741),
    .X(net4740));
 sg13g2_buf_2 fanout4741 (.A(net4749),
    .X(net4741));
 sg13g2_buf_4 fanout4742 (.X(net4742),
    .A(net4749));
 sg13g2_buf_2 fanout4743 (.A(net4749),
    .X(net4743));
 sg13g2_buf_2 fanout4744 (.A(net4746),
    .X(net4744));
 sg13g2_buf_2 fanout4745 (.A(net4746),
    .X(net4745));
 sg13g2_buf_2 fanout4746 (.A(net4749),
    .X(net4746));
 sg13g2_buf_2 fanout4747 (.A(net4749),
    .X(net4747));
 sg13g2_buf_2 fanout4748 (.A(net4749),
    .X(net4748));
 sg13g2_buf_2 fanout4749 (.A(net4764),
    .X(net4749));
 sg13g2_buf_2 fanout4750 (.A(net4751),
    .X(net4750));
 sg13g2_buf_2 fanout4751 (.A(net4763),
    .X(net4751));
 sg13g2_buf_2 fanout4752 (.A(net4754),
    .X(net4752));
 sg13g2_buf_2 fanout4753 (.A(net4754),
    .X(net4753));
 sg13g2_buf_2 fanout4754 (.A(net4763),
    .X(net4754));
 sg13g2_buf_2 fanout4755 (.A(net4759),
    .X(net4755));
 sg13g2_buf_1 fanout4756 (.A(net4759),
    .X(net4756));
 sg13g2_buf_2 fanout4757 (.A(net4759),
    .X(net4757));
 sg13g2_buf_2 fanout4758 (.A(net4759),
    .X(net4758));
 sg13g2_buf_1 fanout4759 (.A(net4763),
    .X(net4759));
 sg13g2_buf_2 fanout4760 (.A(net4761),
    .X(net4760));
 sg13g2_buf_1 fanout4761 (.A(net4762),
    .X(net4761));
 sg13g2_buf_2 fanout4762 (.A(net4763),
    .X(net4762));
 sg13g2_buf_2 fanout4763 (.A(net4764),
    .X(net4763));
 sg13g2_buf_8 fanout4764 (.A(uio_in[3]),
    .X(net4764));
 sg13g2_buf_2 fanout4765 (.A(net4766),
    .X(net4765));
 sg13g2_buf_4 fanout4766 (.X(net4766),
    .A(net4777));
 sg13g2_buf_2 fanout4767 (.A(net4768),
    .X(net4767));
 sg13g2_buf_2 fanout4768 (.A(net4769),
    .X(net4768));
 sg13g2_buf_2 fanout4769 (.A(net4777),
    .X(net4769));
 sg13g2_buf_2 fanout4770 (.A(net4771),
    .X(net4770));
 sg13g2_buf_2 fanout4771 (.A(net4776),
    .X(net4771));
 sg13g2_buf_4 fanout4772 (.X(net4772),
    .A(net4775));
 sg13g2_buf_2 fanout4773 (.A(net4775),
    .X(net4773));
 sg13g2_buf_2 fanout4774 (.A(net4775),
    .X(net4774));
 sg13g2_buf_2 fanout4775 (.A(net4776),
    .X(net4775));
 sg13g2_buf_2 fanout4776 (.A(net4777),
    .X(net4776));
 sg13g2_buf_2 fanout4777 (.A(net4788),
    .X(net4777));
 sg13g2_buf_4 fanout4778 (.X(net4778),
    .A(net4779));
 sg13g2_buf_4 fanout4779 (.X(net4779),
    .A(net4788));
 sg13g2_buf_2 fanout4780 (.A(net4782),
    .X(net4780));
 sg13g2_buf_2 fanout4781 (.A(net4782),
    .X(net4781));
 sg13g2_buf_2 fanout4782 (.A(net4788),
    .X(net4782));
 sg13g2_buf_2 fanout4783 (.A(net4784),
    .X(net4783));
 sg13g2_buf_2 fanout4784 (.A(net4787),
    .X(net4784));
 sg13g2_buf_2 fanout4785 (.A(net4787),
    .X(net4785));
 sg13g2_buf_2 fanout4786 (.A(net4787),
    .X(net4786));
 sg13g2_buf_2 fanout4787 (.A(net4788),
    .X(net4787));
 sg13g2_buf_2 fanout4788 (.A(net4813),
    .X(net4788));
 sg13g2_buf_2 fanout4789 (.A(net4790),
    .X(net4789));
 sg13g2_buf_2 fanout4790 (.A(net4794),
    .X(net4790));
 sg13g2_buf_2 fanout4791 (.A(net4794),
    .X(net4791));
 sg13g2_buf_2 fanout4792 (.A(net4794),
    .X(net4792));
 sg13g2_buf_2 fanout4793 (.A(net4794),
    .X(net4793));
 sg13g2_buf_2 fanout4794 (.A(net4801),
    .X(net4794));
 sg13g2_buf_2 fanout4795 (.A(net4801),
    .X(net4795));
 sg13g2_buf_2 fanout4796 (.A(net4801),
    .X(net4796));
 sg13g2_buf_2 fanout4797 (.A(net4800),
    .X(net4797));
 sg13g2_buf_2 fanout4798 (.A(net4800),
    .X(net4798));
 sg13g2_buf_2 fanout4799 (.A(net4800),
    .X(net4799));
 sg13g2_buf_2 fanout4800 (.A(net4801),
    .X(net4800));
 sg13g2_buf_2 fanout4801 (.A(net4813),
    .X(net4801));
 sg13g2_buf_2 fanout4802 (.A(net4804),
    .X(net4802));
 sg13g2_buf_2 fanout4803 (.A(net4804),
    .X(net4803));
 sg13g2_buf_2 fanout4804 (.A(net4806),
    .X(net4804));
 sg13g2_buf_2 fanout4805 (.A(net4806),
    .X(net4805));
 sg13g2_buf_1 fanout4806 (.A(net4813),
    .X(net4806));
 sg13g2_buf_2 fanout4807 (.A(net4812),
    .X(net4807));
 sg13g2_buf_2 fanout4808 (.A(net4810),
    .X(net4808));
 sg13g2_buf_2 fanout4809 (.A(net4810),
    .X(net4809));
 sg13g2_buf_2 fanout4810 (.A(net4812),
    .X(net4810));
 sg13g2_buf_2 fanout4811 (.A(net4812),
    .X(net4811));
 sg13g2_buf_2 fanout4812 (.A(net4813),
    .X(net4812));
 sg13g2_buf_4 fanout4813 (.X(net4813),
    .A(uio_in[3]));
 sg13g2_buf_2 input1 (.A(rst_n),
    .X(net1));
 sg13g2_buf_8 input2 (.A(ui_in[0]),
    .X(net2));
 sg13g2_buf_8 input3 (.A(ui_in[1]),
    .X(net3));
 sg13g2_buf_8 input4 (.A(ui_in[2]),
    .X(net4));
 sg13g2_buf_4 input5 (.X(net5),
    .A(ui_in[3]));
 sg13g2_buf_8 input6 (.A(ui_in[4]),
    .X(net6));
 sg13g2_buf_8 input7 (.A(ui_in[5]),
    .X(net7));
 sg13g2_buf_8 input8 (.A(ui_in[6]),
    .X(net8));
 sg13g2_buf_8 input9 (.A(ui_in[7]),
    .X(net9));
 sg13g2_buf_8 input10 (.A(uio_in[0]),
    .X(net10));
 sg13g2_buf_8 input11 (.A(uio_in[1]),
    .X(net11));
 sg13g2_buf_4 input12 (.X(net12),
    .A(uio_in[4]));
 sg13g2_buf_4 input13 (.X(net13),
    .A(uio_in[6]));
 sg13g2_buf_16 max_cap14 (.X(net14),
    .A(_03272_));
 sg13g2_buf_16 max_cap15 (.X(net15),
    .A(_03256_));
 sg13g2_tielo tt_um_snn_with_delays_paolaunisa_16 (.L_LO(net16));
 sg13g2_buf_2 clkbuf_leaf_1_clk (.A(clknet_4_0__leaf_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_2 clkbuf_leaf_2_clk (.A(clknet_4_0__leaf_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_2 clkbuf_leaf_3_clk (.A(clknet_4_2__leaf_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_2 clkbuf_leaf_4_clk (.A(clknet_4_2__leaf_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_2 clkbuf_leaf_5_clk (.A(clknet_4_1__leaf_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_2 clkbuf_leaf_6_clk (.A(clknet_4_0__leaf_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_2 clkbuf_leaf_7_clk (.A(clknet_4_1__leaf_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_2 clkbuf_leaf_8_clk (.A(clknet_4_1__leaf_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_2 clkbuf_leaf_9_clk (.A(clknet_4_1__leaf_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_2 clkbuf_leaf_10_clk (.A(clknet_4_1__leaf_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_2 clkbuf_leaf_11_clk (.A(clknet_4_12__leaf_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_2 clkbuf_leaf_12_clk (.A(clknet_4_7__leaf_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_2 clkbuf_leaf_13_clk (.A(clknet_4_2__leaf_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_2 clkbuf_leaf_14_clk (.A(clknet_4_3__leaf_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_2 clkbuf_leaf_15_clk (.A(clknet_4_4__leaf_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_2 clkbuf_leaf_16_clk (.A(clknet_4_4__leaf_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_2 clkbuf_leaf_17_clk (.A(clknet_4_4__leaf_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_2 clkbuf_leaf_18_clk (.A(clknet_4_4__leaf_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_2 clkbuf_leaf_19_clk (.A(clknet_4_5__leaf_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_2 clkbuf_leaf_20_clk (.A(clknet_4_6__leaf_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_2 clkbuf_leaf_21_clk (.A(clknet_4_6__leaf_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_2 clkbuf_leaf_22_clk (.A(clknet_4_4__leaf_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_2 clkbuf_leaf_23_clk (.A(clknet_4_5__leaf_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_2 clkbuf_leaf_24_clk (.A(clknet_4_5__leaf_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_2 clkbuf_leaf_25_clk (.A(clknet_4_5__leaf_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_2 clkbuf_leaf_26_clk (.A(clknet_4_5__leaf_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_2 clkbuf_leaf_27_clk (.A(clknet_4_6__leaf_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_2 clkbuf_leaf_28_clk (.A(clknet_4_6__leaf_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_2 clkbuf_leaf_29_clk (.A(clknet_4_7__leaf_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_2 clkbuf_leaf_30_clk (.A(clknet_4_6__leaf_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_2 clkbuf_leaf_31_clk (.A(clknet_4_7__leaf_clk),
    .X(clknet_leaf_31_clk));
 sg13g2_buf_2 clkbuf_leaf_32_clk (.A(clknet_4_7__leaf_clk),
    .X(clknet_leaf_32_clk));
 sg13g2_buf_2 clkbuf_leaf_33_clk (.A(clknet_4_12__leaf_clk),
    .X(clknet_leaf_33_clk));
 sg13g2_buf_2 clkbuf_leaf_34_clk (.A(clknet_4_12__leaf_clk),
    .X(clknet_leaf_34_clk));
 sg13g2_buf_2 clkbuf_leaf_35_clk (.A(clknet_4_12__leaf_clk),
    .X(clknet_leaf_35_clk));
 sg13g2_buf_2 clkbuf_leaf_36_clk (.A(clknet_4_8__leaf_clk),
    .X(clknet_leaf_36_clk));
 sg13g2_buf_2 clkbuf_leaf_37_clk (.A(clknet_4_12__leaf_clk),
    .X(clknet_leaf_37_clk));
 sg13g2_buf_2 clkbuf_leaf_38_clk (.A(clknet_4_13__leaf_clk),
    .X(clknet_leaf_38_clk));
 sg13g2_buf_2 clkbuf_leaf_39_clk (.A(clknet_4_13__leaf_clk),
    .X(clknet_leaf_39_clk));
 sg13g2_buf_2 clkbuf_leaf_40_clk (.A(clknet_4_13__leaf_clk),
    .X(clknet_leaf_40_clk));
 sg13g2_buf_2 clkbuf_leaf_41_clk (.A(clknet_4_15__leaf_clk),
    .X(clknet_leaf_41_clk));
 sg13g2_buf_2 clkbuf_leaf_42_clk (.A(clknet_4_15__leaf_clk),
    .X(clknet_leaf_42_clk));
 sg13g2_buf_2 clkbuf_leaf_43_clk (.A(clknet_4_15__leaf_clk),
    .X(clknet_leaf_43_clk));
 sg13g2_buf_2 clkbuf_leaf_44_clk (.A(clknet_4_15__leaf_clk),
    .X(clknet_leaf_44_clk));
 sg13g2_buf_2 clkbuf_leaf_45_clk (.A(clknet_4_13__leaf_clk),
    .X(clknet_leaf_45_clk));
 sg13g2_buf_2 clkbuf_leaf_46_clk (.A(clknet_4_14__leaf_clk),
    .X(clknet_leaf_46_clk));
 sg13g2_buf_2 clkbuf_leaf_47_clk (.A(clknet_4_14__leaf_clk),
    .X(clknet_leaf_47_clk));
 sg13g2_buf_2 clkbuf_leaf_48_clk (.A(clknet_4_14__leaf_clk),
    .X(clknet_leaf_48_clk));
 sg13g2_buf_2 clkbuf_leaf_49_clk (.A(clknet_4_14__leaf_clk),
    .X(clknet_leaf_49_clk));
 sg13g2_buf_2 clkbuf_leaf_50_clk (.A(clknet_4_13__leaf_clk),
    .X(clknet_leaf_50_clk));
 sg13g2_buf_2 clkbuf_leaf_51_clk (.A(clknet_4_11__leaf_clk),
    .X(clknet_leaf_51_clk));
 sg13g2_buf_2 clkbuf_leaf_52_clk (.A(clknet_4_11__leaf_clk),
    .X(clknet_leaf_52_clk));
 sg13g2_buf_2 clkbuf_leaf_53_clk (.A(clknet_4_14__leaf_clk),
    .X(clknet_leaf_53_clk));
 sg13g2_buf_2 clkbuf_leaf_54_clk (.A(clknet_4_10__leaf_clk),
    .X(clknet_leaf_54_clk));
 sg13g2_buf_2 clkbuf_leaf_55_clk (.A(clknet_4_11__leaf_clk),
    .X(clknet_leaf_55_clk));
 sg13g2_buf_2 clkbuf_leaf_56_clk (.A(clknet_4_10__leaf_clk),
    .X(clknet_leaf_56_clk));
 sg13g2_buf_2 clkbuf_leaf_57_clk (.A(clknet_4_10__leaf_clk),
    .X(clknet_leaf_57_clk));
 sg13g2_buf_2 clkbuf_leaf_58_clk (.A(clknet_4_10__leaf_clk),
    .X(clknet_leaf_58_clk));
 sg13g2_buf_2 clkbuf_leaf_59_clk (.A(clknet_4_10__leaf_clk),
    .X(clknet_leaf_59_clk));
 sg13g2_buf_2 clkbuf_leaf_60_clk (.A(clknet_4_11__leaf_clk),
    .X(clknet_leaf_60_clk));
 sg13g2_buf_2 clkbuf_leaf_61_clk (.A(clknet_4_8__leaf_clk),
    .X(clknet_leaf_61_clk));
 sg13g2_buf_2 clkbuf_leaf_62_clk (.A(clknet_4_8__leaf_clk),
    .X(clknet_leaf_62_clk));
 sg13g2_buf_2 clkbuf_leaf_63_clk (.A(clknet_4_8__leaf_clk),
    .X(clknet_leaf_63_clk));
 sg13g2_buf_2 clkbuf_leaf_64_clk (.A(clknet_4_8__leaf_clk),
    .X(clknet_leaf_64_clk));
 sg13g2_buf_2 clkbuf_leaf_65_clk (.A(clknet_4_9__leaf_clk),
    .X(clknet_leaf_65_clk));
 sg13g2_buf_2 clkbuf_leaf_66_clk (.A(clknet_4_9__leaf_clk),
    .X(clknet_leaf_66_clk));
 sg13g2_buf_2 clkbuf_leaf_67_clk (.A(clknet_4_9__leaf_clk),
    .X(clknet_leaf_67_clk));
 sg13g2_buf_2 clkbuf_leaf_68_clk (.A(clknet_4_9__leaf_clk),
    .X(clknet_leaf_68_clk));
 sg13g2_buf_2 clkbuf_leaf_69_clk (.A(clknet_4_9__leaf_clk),
    .X(clknet_leaf_69_clk));
 sg13g2_buf_2 clkbuf_leaf_70_clk (.A(clknet_4_3__leaf_clk),
    .X(clknet_leaf_70_clk));
 sg13g2_buf_2 clkbuf_leaf_71_clk (.A(clknet_4_3__leaf_clk),
    .X(clknet_leaf_71_clk));
 sg13g2_buf_2 clkbuf_leaf_72_clk (.A(clknet_4_3__leaf_clk),
    .X(clknet_leaf_72_clk));
 sg13g2_buf_2 clkbuf_leaf_73_clk (.A(clknet_4_2__leaf_clk),
    .X(clknet_leaf_73_clk));
 sg13g2_buf_2 clkbuf_leaf_74_clk (.A(clknet_4_2__leaf_clk),
    .X(clknet_leaf_74_clk));
 sg13g2_buf_2 clkbuf_leaf_75_clk (.A(clknet_4_0__leaf_clk),
    .X(clknet_leaf_75_clk));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_2 clkbuf_2_0_0_clk (.A(clknet_0_clk),
    .X(clknet_2_0_0_clk));
 sg13g2_buf_2 clkbuf_2_1_0_clk (.A(clknet_0_clk),
    .X(clknet_2_1_0_clk));
 sg13g2_buf_2 clkbuf_2_2_0_clk (.A(clknet_0_clk),
    .X(clknet_2_2_0_clk));
 sg13g2_buf_2 clkbuf_2_3_0_clk (.A(clknet_0_clk),
    .X(clknet_2_3_0_clk));
 sg13g2_buf_2 clkbuf_4_0__f_clk (.A(clknet_2_0_0_clk),
    .X(clknet_4_0__leaf_clk));
 sg13g2_buf_2 clkbuf_4_1__f_clk (.A(clknet_2_0_0_clk),
    .X(clknet_4_1__leaf_clk));
 sg13g2_buf_2 clkbuf_4_2__f_clk (.A(clknet_2_0_0_clk),
    .X(clknet_4_2__leaf_clk));
 sg13g2_buf_2 clkbuf_4_3__f_clk (.A(clknet_2_0_0_clk),
    .X(clknet_4_3__leaf_clk));
 sg13g2_buf_2 clkbuf_4_4__f_clk (.A(clknet_2_1_0_clk),
    .X(clknet_4_4__leaf_clk));
 sg13g2_buf_2 clkbuf_4_5__f_clk (.A(clknet_2_1_0_clk),
    .X(clknet_4_5__leaf_clk));
 sg13g2_buf_2 clkbuf_4_6__f_clk (.A(clknet_2_1_0_clk),
    .X(clknet_4_6__leaf_clk));
 sg13g2_buf_2 clkbuf_4_7__f_clk (.A(clknet_2_1_0_clk),
    .X(clknet_4_7__leaf_clk));
 sg13g2_buf_2 clkbuf_4_8__f_clk (.A(clknet_2_2_0_clk),
    .X(clknet_4_8__leaf_clk));
 sg13g2_buf_2 clkbuf_4_9__f_clk (.A(clknet_2_2_0_clk),
    .X(clknet_4_9__leaf_clk));
 sg13g2_buf_2 clkbuf_4_10__f_clk (.A(clknet_2_2_0_clk),
    .X(clknet_4_10__leaf_clk));
 sg13g2_buf_2 clkbuf_4_11__f_clk (.A(clknet_2_2_0_clk),
    .X(clknet_4_11__leaf_clk));
 sg13g2_buf_2 clkbuf_4_12__f_clk (.A(clknet_2_3_0_clk),
    .X(clknet_4_12__leaf_clk));
 sg13g2_buf_2 clkbuf_4_13__f_clk (.A(clknet_2_3_0_clk),
    .X(clknet_4_13__leaf_clk));
 sg13g2_buf_2 clkbuf_4_14__f_clk (.A(clknet_2_3_0_clk),
    .X(clknet_4_14__leaf_clk));
 sg13g2_buf_2 clkbuf_4_15__f_clk (.A(clknet_2_3_0_clk),
    .X(clknet_4_15__leaf_clk));
 sg13g2_buf_2 clkload0 (.A(clknet_4_3__leaf_clk));
 sg13g2_buf_2 clkload1 (.A(clknet_4_7__leaf_clk));
 sg13g2_buf_2 clkload2 (.A(clknet_4_11__leaf_clk));
 sg13g2_buf_2 clkload3 (.A(clknet_4_15__leaf_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_leaf_2_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_leaf_6_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_leaf_75_clk));
 sg13g2_inv_1 clkload7 (.A(clknet_leaf_5_clk));
 sg13g2_inv_4 clkload8 (.A(clknet_leaf_7_clk));
 sg13g2_inv_8 clkload9 (.A(clknet_leaf_10_clk));
 sg13g2_inv_8 clkload10 (.A(clknet_leaf_3_clk));
 sg13g2_inv_2 clkload11 (.A(clknet_leaf_71_clk));
 sg13g2_inv_1 clkload12 (.A(clknet_leaf_72_clk));
 sg13g2_inv_8 clkload13 (.A(clknet_leaf_22_clk));
 sg13g2_inv_4 clkload14 (.A(clknet_leaf_21_clk));
 sg13g2_inv_2 clkload15 (.A(clknet_leaf_28_clk));
 sg13g2_inv_2 clkload16 (.A(clknet_leaf_12_clk));
 sg13g2_inv_4 clkload17 (.A(clknet_leaf_66_clk));
 sg13g2_inv_2 clkload18 (.A(clknet_leaf_54_clk));
 sg13g2_inv_4 clkload19 (.A(clknet_leaf_57_clk));
 sg13g2_inv_1 clkload20 (.A(clknet_leaf_51_clk));
 sg13g2_inv_4 clkload21 (.A(clknet_leaf_52_clk));
 sg13g2_inv_8 clkload22 (.A(clknet_leaf_33_clk));
 sg13g2_inv_4 clkload23 (.A(clknet_leaf_45_clk));
 sg13g2_inv_4 clkload24 (.A(clknet_leaf_50_clk));
 sg13g2_inv_4 clkload25 (.A(clknet_leaf_46_clk));
 sg13g2_inv_8 clkload26 (.A(clknet_leaf_48_clk));
 sg13g2_inv_2 clkload27 (.A(clknet_leaf_53_clk));
 sg13g2_inv_4 clkload28 (.A(clknet_leaf_42_clk));
 sg13g2_inv_4 clkload29 (.A(clknet_leaf_44_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\spiking_network_top_uut.clk_div_sync.sync_ff1 ),
    .X(net31));
 sg13g2_dlygate4sd3_1 hold2 (.A(\spiking_network_top_uut.input_ready_sync_inst.sync_ff1 ),
    .X(net32));
 sg13g2_dlygate4sd3_1 hold3 (.A(\spiking_network_top_uut.debug_config_sync.sync_ff1 ),
    .X(net33));
 sg13g2_dlygate4sd3_1 hold4 (.A(\spiking_network_top_uut.snn_en_sync_inst.sync_ff1 ),
    .X(net34));
 sg13g2_dlygate4sd3_1 hold5 (.A(\spiking_network_top_uut.u_sys_clk_reset.reset_ff1 ),
    .X(net35));
 sg13g2_dlygate4sd3_1 hold6 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_reg1 ),
    .X(net36));
 sg13g2_dlygate4sd3_1 hold7 (.A(_00629_),
    .X(net37));
 sg13g2_dlygate4sd3_1 hold8 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_reg1 ),
    .X(net38));
 sg13g2_dlygate4sd3_1 hold9 (.A(_00856_),
    .X(net39));
 sg13g2_dlygate4sd3_1 hold10 (.A(_00000_),
    .X(net40));
 sg13g2_dlygate4sd3_1 hold11 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_reg1 ),
    .X(net41));
 sg13g2_dlygate4sd3_1 hold12 (.A(_00912_),
    .X(net42));
 sg13g2_dlygate4sd3_1 hold13 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_reg1 ),
    .X(net43));
 sg13g2_dlygate4sd3_1 hold14 (.A(_00860_),
    .X(net44));
 sg13g2_dlygate4sd3_1 hold15 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_reg1 ),
    .X(net45));
 sg13g2_dlygate4sd3_1 hold16 (.A(_00986_),
    .X(net46));
 sg13g2_dlygate4sd3_1 hold17 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_reg1 ),
    .X(net47));
 sg13g2_dlygate4sd3_1 hold18 (.A(_01022_),
    .X(net48));
 sg13g2_dlygate4sd3_1 hold19 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_reg1 ),
    .X(net49));
 sg13g2_dlygate4sd3_1 hold20 (.A(_00964_),
    .X(net50));
 sg13g2_dlygate4sd3_1 hold21 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_reg1 ),
    .X(net51));
 sg13g2_dlygate4sd3_1 hold22 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_reg1 ),
    .X(net52));
 sg13g2_dlygate4sd3_1 hold23 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_reg1 ),
    .X(net53));
 sg13g2_dlygate4sd3_1 hold24 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[1].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_reg1 ),
    .X(net54));
 sg13g2_dlygate4sd3_1 hold25 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_dout ),
    .X(net55));
 sg13g2_dlygate4sd3_1 hold26 (.A(_00930_),
    .X(net56));
 sg13g2_dlygate4sd3_1 hold27 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_reg1 ),
    .X(net57));
 sg13g2_dlygate4sd3_1 hold28 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_reg1 ),
    .X(net58));
 sg13g2_dlygate4sd3_1 hold29 (.A(_00699_),
    .X(net59));
 sg13g2_dlygate4sd3_1 hold30 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[1].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_reg1 ),
    .X(net60));
 sg13g2_dlygate4sd3_1 hold31 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_reg1 ),
    .X(net61));
 sg13g2_dlygate4sd3_1 hold32 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_reg1 ),
    .X(net62));
 sg13g2_dlygate4sd3_1 hold33 (.A(_00623_),
    .X(net63));
 sg13g2_dlygate4sd3_1 hold34 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_reg1 ),
    .X(net64));
 sg13g2_dlygate4sd3_1 hold35 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_reg1 ),
    .X(net65));
 sg13g2_dlygate4sd3_1 hold36 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_reg1 ),
    .X(net66));
 sg13g2_dlygate4sd3_1 hold37 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_reg1 ),
    .X(net67));
 sg13g2_dlygate4sd3_1 hold38 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_reg1 ),
    .X(net68));
 sg13g2_dlygate4sd3_1 hold39 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_reg1 ),
    .X(net69));
 sg13g2_dlygate4sd3_1 hold40 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_reg1 ),
    .X(net70));
 sg13g2_dlygate4sd3_1 hold41 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_reg1 ),
    .X(net71));
 sg13g2_dlygate4sd3_1 hold42 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_reg1 ),
    .X(net72));
 sg13g2_dlygate4sd3_1 hold43 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_reg1 ),
    .X(net73));
 sg13g2_dlygate4sd3_1 hold44 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_reg1 ),
    .X(net74));
 sg13g2_dlygate4sd3_1 hold45 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_reg1 ),
    .X(net75));
 sg13g2_dlygate4sd3_1 hold46 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_reg1 ),
    .X(net76));
 sg13g2_dlygate4sd3_1 hold47 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_reg1 ),
    .X(net77));
 sg13g2_dlygate4sd3_1 hold48 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_reg1 ),
    .X(net78));
 sg13g2_dlygate4sd3_1 hold49 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_reg1 ),
    .X(net79));
 sg13g2_dlygate4sd3_1 hold50 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_reg1 ),
    .X(net80));
 sg13g2_dlygate4sd3_1 hold51 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_reg1 ),
    .X(net81));
 sg13g2_dlygate4sd3_1 hold52 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_reg1 ),
    .X(net82));
 sg13g2_dlygate4sd3_1 hold53 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[1].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_reg1 ),
    .X(net83));
 sg13g2_dlygate4sd3_1 hold54 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_dout ),
    .X(net84));
 sg13g2_dlygate4sd3_1 hold55 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_reg1 ),
    .X(net85));
 sg13g2_dlygate4sd3_1 hold56 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_reg1 ),
    .X(net86));
 sg13g2_dlygate4sd3_1 hold57 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_reg1 ),
    .X(net87));
 sg13g2_dlygate4sd3_1 hold58 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_reg1 ),
    .X(net88));
 sg13g2_dlygate4sd3_1 hold59 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_reg1 ),
    .X(net89));
 sg13g2_dlygate4sd3_1 hold60 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_reg1 ),
    .X(net90));
 sg13g2_dlygate4sd3_1 hold61 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_reg1 ),
    .X(net91));
 sg13g2_dlygate4sd3_1 hold62 (.A(_00439_),
    .X(net92));
 sg13g2_dlygate4sd3_1 hold63 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_reg1 ),
    .X(net93));
 sg13g2_dlygate4sd3_1 hold64 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_reg1 ),
    .X(net94));
 sg13g2_dlygate4sd3_1 hold65 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_reg1 ),
    .X(net95));
 sg13g2_dlygate4sd3_1 hold66 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_reg1 ),
    .X(net96));
 sg13g2_dlygate4sd3_1 hold67 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_reg1 ),
    .X(net97));
 sg13g2_dlygate4sd3_1 hold68 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_reg1 ),
    .X(net98));
 sg13g2_dlygate4sd3_1 hold69 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_reg1 ),
    .X(net99));
 sg13g2_dlygate4sd3_1 hold70 (.A(\spiking_network_top_uut.clk_div_inst.counter[1] ),
    .X(net100));
 sg13g2_dlygate4sd3_1 hold71 (.A(_03174_),
    .X(net101));
 sg13g2_dlygate4sd3_1 hold72 (.A(_01093_),
    .X(net102));
 sg13g2_dlygate4sd3_1 hold73 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_reg1 ),
    .X(net103));
 sg13g2_dlygate4sd3_1 hold74 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_reg1 ),
    .X(net104));
 sg13g2_dlygate4sd3_1 hold75 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_reg1 ),
    .X(net105));
 sg13g2_dlygate4sd3_1 hold76 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_reg1 ),
    .X(net106));
 sg13g2_dlygate4sd3_1 hold77 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_reg1 ),
    .X(net107));
 sg13g2_dlygate4sd3_1 hold78 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_reg1 ),
    .X(net108));
 sg13g2_dlygate4sd3_1 hold79 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_reg1 ),
    .X(net109));
 sg13g2_dlygate4sd3_1 hold80 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_reg1 ),
    .X(net110));
 sg13g2_dlygate4sd3_1 hold81 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_dout ),
    .X(net111));
 sg13g2_dlygate4sd3_1 hold82 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_reg1 ),
    .X(net112));
 sg13g2_dlygate4sd3_1 hold83 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_reg1 ),
    .X(net113));
 sg13g2_dlygate4sd3_1 hold84 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_reg1 ),
    .X(net114));
 sg13g2_dlygate4sd3_1 hold85 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_reg1 ),
    .X(net115));
 sg13g2_dlygate4sd3_1 hold86 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_reg1 ),
    .X(net116));
 sg13g2_dlygate4sd3_1 hold87 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_reg1 ),
    .X(net117));
 sg13g2_dlygate4sd3_1 hold88 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_reg1 ),
    .X(net118));
 sg13g2_dlygate4sd3_1 hold89 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_reg1 ),
    .X(net119));
 sg13g2_dlygate4sd3_1 hold90 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_reg1 ),
    .X(net120));
 sg13g2_dlygate4sd3_1 hold91 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_reg1 ),
    .X(net121));
 sg13g2_dlygate4sd3_1 hold92 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_reg1 ),
    .X(net122));
 sg13g2_dlygate4sd3_1 hold93 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_dout ),
    .X(net123));
 sg13g2_dlygate4sd3_1 hold94 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_dout ),
    .X(net124));
 sg13g2_dlygate4sd3_1 hold95 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_dout ),
    .X(net125));
 sg13g2_dlygate4sd3_1 hold96 (.A(_00852_),
    .X(net126));
 sg13g2_dlygate4sd3_1 hold97 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[1].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_reg1 ),
    .X(net127));
 sg13g2_dlygate4sd3_1 hold98 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_reg1 ),
    .X(net128));
 sg13g2_dlygate4sd3_1 hold99 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_reg1 ),
    .X(net129));
 sg13g2_dlygate4sd3_1 hold100 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_reg1 ),
    .X(net130));
 sg13g2_dlygate4sd3_1 hold101 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_reg1 ),
    .X(net131));
 sg13g2_dlygate4sd3_1 hold102 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_reg1 ),
    .X(net132));
 sg13g2_dlygate4sd3_1 hold103 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_reg1 ),
    .X(net133));
 sg13g2_dlygate4sd3_1 hold104 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_reg1 ),
    .X(net134));
 sg13g2_dlygate4sd3_1 hold105 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_reg1 ),
    .X(net135));
 sg13g2_dlygate4sd3_1 hold106 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_reg1 ),
    .X(net136));
 sg13g2_dlygate4sd3_1 hold107 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[1].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_reg1 ),
    .X(net137));
 sg13g2_dlygate4sd3_1 hold108 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_reg1 ),
    .X(net138));
 sg13g2_dlygate4sd3_1 hold109 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_reg1 ),
    .X(net139));
 sg13g2_dlygate4sd3_1 hold110 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_reg1 ),
    .X(net140));
 sg13g2_dlygate4sd3_1 hold111 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_reg1 ),
    .X(net141));
 sg13g2_dlygate4sd3_1 hold112 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_reg1 ),
    .X(net142));
 sg13g2_dlygate4sd3_1 hold113 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[1].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_reg1 ),
    .X(net143));
 sg13g2_dlygate4sd3_1 hold114 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_reg1 ),
    .X(net144));
 sg13g2_dlygate4sd3_1 hold115 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_reg1 ),
    .X(net145));
 sg13g2_dlygate4sd3_1 hold116 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_dout ),
    .X(net146));
 sg13g2_dlygate4sd3_1 hold117 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[1].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_dout ),
    .X(net147));
 sg13g2_dlygate4sd3_1 hold118 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_reg1 ),
    .X(net148));
 sg13g2_dlygate4sd3_1 hold119 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_reg1 ),
    .X(net149));
 sg13g2_dlygate4sd3_1 hold120 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_reg1 ),
    .X(net150));
 sg13g2_dlygate4sd3_1 hold121 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_reg1 ),
    .X(net151));
 sg13g2_dlygate4sd3_1 hold122 (.A(_00938_),
    .X(net152));
 sg13g2_dlygate4sd3_1 hold123 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[2] ),
    .X(net153));
 sg13g2_dlygate4sd3_1 hold124 (.A(_00558_),
    .X(net154));
 sg13g2_dlygate4sd3_1 hold125 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_reg1 ),
    .X(net155));
 sg13g2_dlygate4sd3_1 hold126 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[2] ),
    .X(net156));
 sg13g2_dlygate4sd3_1 hold127 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_dout ),
    .X(net157));
 sg13g2_dlygate4sd3_1 hold128 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_dout ),
    .X(net158));
 sg13g2_dlygate4sd3_1 hold129 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_reg1 ),
    .X(net159));
 sg13g2_dlygate4sd3_1 hold130 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[2] ),
    .X(net160));
 sg13g2_dlygate4sd3_1 hold131 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_reg1 ),
    .X(net161));
 sg13g2_dlygate4sd3_1 hold132 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_dout ),
    .X(net162));
 sg13g2_dlygate4sd3_1 hold133 (.A(_00904_),
    .X(net163));
 sg13g2_dlygate4sd3_1 hold134 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_reg1 ),
    .X(net164));
 sg13g2_dlygate4sd3_1 hold135 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_reg1 ),
    .X(net165));
 sg13g2_dlygate4sd3_1 hold136 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_dout ),
    .X(net166));
 sg13g2_dlygate4sd3_1 hold137 (.A(_00666_),
    .X(net167));
 sg13g2_dlygate4sd3_1 hold138 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_reg1 ),
    .X(net168));
 sg13g2_dlygate4sd3_1 hold139 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_reg1 ),
    .X(net169));
 sg13g2_dlygate4sd3_1 hold140 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_reg1 ),
    .X(net170));
 sg13g2_dlygate4sd3_1 hold141 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_reg1 ),
    .X(net171));
 sg13g2_dlygate4sd3_1 hold142 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_reg1 ),
    .X(net172));
 sg13g2_dlygate4sd3_1 hold143 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[2] ),
    .X(net173));
 sg13g2_dlygate4sd3_1 hold144 (.A(_00830_),
    .X(net174));
 sg13g2_dlygate4sd3_1 hold145 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_dout ),
    .X(net175));
 sg13g2_dlygate4sd3_1 hold146 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_reg1 ),
    .X(net176));
 sg13g2_dlygate4sd3_1 hold147 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_dout ),
    .X(net177));
 sg13g2_dlygate4sd3_1 hold148 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_reg1 ),
    .X(net178));
 sg13g2_dlygate4sd3_1 hold149 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_dout ),
    .X(net179));
 sg13g2_dlygate4sd3_1 hold150 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_reg1 ),
    .X(net180));
 sg13g2_dlygate4sd3_1 hold151 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_reg1 ),
    .X(net181));
 sg13g2_dlygate4sd3_1 hold152 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_dout ),
    .X(net182));
 sg13g2_dlygate4sd3_1 hold153 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[2] ),
    .X(net183));
 sg13g2_dlygate4sd3_1 hold154 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_dout ),
    .X(net184));
 sg13g2_dlygate4sd3_1 hold155 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_dout ),
    .X(net185));
 sg13g2_dlygate4sd3_1 hold156 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_reg1 ),
    .X(net186));
 sg13g2_dlygate4sd3_1 hold157 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_reg1 ),
    .X(net187));
 sg13g2_dlygate4sd3_1 hold158 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_reg1 ),
    .X(net188));
 sg13g2_dlygate4sd3_1 hold159 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_reg1 ),
    .X(net189));
 sg13g2_dlygate4sd3_1 hold160 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[2] ),
    .X(net190));
 sg13g2_dlygate4sd3_1 hold161 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_dout ),
    .X(net191));
 sg13g2_dlygate4sd3_1 hold162 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_reg1 ),
    .X(net192));
 sg13g2_dlygate4sd3_1 hold163 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_reg1 ),
    .X(net193));
 sg13g2_dlygate4sd3_1 hold164 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[2] ),
    .X(net194));
 sg13g2_dlygate4sd3_1 hold165 (.A(_00890_),
    .X(net195));
 sg13g2_dlygate4sd3_1 hold166 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_dout ),
    .X(net196));
 sg13g2_dlygate4sd3_1 hold167 (.A(_00800_),
    .X(net197));
 sg13g2_dlygate4sd3_1 hold168 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_reg1 ),
    .X(net198));
 sg13g2_dlygate4sd3_1 hold169 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_reg1 ),
    .X(net199));
 sg13g2_dlygate4sd3_1 hold170 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_dout ),
    .X(net200));
 sg13g2_dlygate4sd3_1 hold171 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[2] ),
    .X(net201));
 sg13g2_dlygate4sd3_1 hold172 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_dout ),
    .X(net202));
 sg13g2_dlygate4sd3_1 hold173 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[1].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_dout ),
    .X(net203));
 sg13g2_dlygate4sd3_1 hold174 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[1].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_reg1 ),
    .X(net204));
 sg13g2_dlygate4sd3_1 hold175 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_reg1 ),
    .X(net205));
 sg13g2_dlygate4sd3_1 hold176 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[2] ),
    .X(net206));
 sg13g2_dlygate4sd3_1 hold177 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_dout ),
    .X(net207));
 sg13g2_dlygate4sd3_1 hold178 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[2] ),
    .X(net208));
 sg13g2_dlygate4sd3_1 hold179 (.A(_00637_),
    .X(net209));
 sg13g2_dlygate4sd3_1 hold180 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[2] ),
    .X(net210));
 sg13g2_dlygate4sd3_1 hold181 (.A(_00797_),
    .X(net211));
 sg13g2_dlygate4sd3_1 hold182 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[2] ),
    .X(net212));
 sg13g2_dlygate4sd3_1 hold183 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[2] ),
    .X(net213));
 sg13g2_dlygate4sd3_1 hold184 (.A(_00715_),
    .X(net214));
 sg13g2_dlygate4sd3_1 hold185 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_reg1 ),
    .X(net215));
 sg13g2_dlygate4sd3_1 hold186 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_dout ),
    .X(net216));
 sg13g2_dlygate4sd3_1 hold187 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_reg1 ),
    .X(net217));
 sg13g2_dlygate4sd3_1 hold188 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[4] ),
    .X(net218));
 sg13g2_dlygate4sd3_1 hold189 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[1].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_reg1 ),
    .X(net219));
 sg13g2_dlygate4sd3_1 hold190 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_reg1 ),
    .X(net220));
 sg13g2_dlygate4sd3_1 hold191 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_dout ),
    .X(net221));
 sg13g2_dlygate4sd3_1 hold192 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_dout ),
    .X(net222));
 sg13g2_dlygate4sd3_1 hold193 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_dout ),
    .X(net223));
 sg13g2_dlygate4sd3_1 hold194 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_reg1 ),
    .X(net224));
 sg13g2_dlygate4sd3_1 hold195 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[4] ),
    .X(net225));
 sg13g2_dlygate4sd3_1 hold196 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_dout ),
    .X(net226));
 sg13g2_dlygate4sd3_1 hold197 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_reg1 ),
    .X(net227));
 sg13g2_dlygate4sd3_1 hold198 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_reg1 ),
    .X(net228));
 sg13g2_dlygate4sd3_1 hold199 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[2] ),
    .X(net229));
 sg13g2_dlygate4sd3_1 hold200 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_dout ),
    .X(net230));
 sg13g2_dlygate4sd3_1 hold201 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_dout ),
    .X(net231));
 sg13g2_dlygate4sd3_1 hold202 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_reg1 ),
    .X(net232));
 sg13g2_dlygate4sd3_1 hold203 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_dout ),
    .X(net233));
 sg13g2_dlygate4sd3_1 hold204 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_dout ),
    .X(net234));
 sg13g2_dlygate4sd3_1 hold205 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[2] ),
    .X(net235));
 sg13g2_dlygate4sd3_1 hold206 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_dout ),
    .X(net236));
 sg13g2_dlygate4sd3_1 hold207 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[1].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_dout ),
    .X(net237));
 sg13g2_dlygate4sd3_1 hold208 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_dout ),
    .X(net238));
 sg13g2_dlygate4sd3_1 hold209 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_dout ),
    .X(net239));
 sg13g2_dlygate4sd3_1 hold210 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_reg1 ),
    .X(net240));
 sg13g2_dlygate4sd3_1 hold211 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_dout ),
    .X(net241));
 sg13g2_dlygate4sd3_1 hold212 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_dout ),
    .X(net242));
 sg13g2_dlygate4sd3_1 hold213 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_dout ),
    .X(net243));
 sg13g2_dlygate4sd3_1 hold214 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[2] ),
    .X(net244));
 sg13g2_dlygate4sd3_1 hold215 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_dout ),
    .X(net245));
 sg13g2_dlygate4sd3_1 hold216 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_reg1 ),
    .X(net246));
 sg13g2_dlygate4sd3_1 hold217 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_dout ),
    .X(net247));
 sg13g2_dlygate4sd3_1 hold218 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_dout ),
    .X(net248));
 sg13g2_dlygate4sd3_1 hold219 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_reg1 ),
    .X(net249));
 sg13g2_dlygate4sd3_1 hold220 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[4] ),
    .X(net250));
 sg13g2_dlygate4sd3_1 hold221 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_reg1 ),
    .X(net251));
 sg13g2_dlygate4sd3_1 hold222 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_dout ),
    .X(net252));
 sg13g2_dlygate4sd3_1 hold223 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_dout ),
    .X(net253));
 sg13g2_dlygate4sd3_1 hold224 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_reg1 ),
    .X(net254));
 sg13g2_dlygate4sd3_1 hold225 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_dout ),
    .X(net255));
 sg13g2_dlygate4sd3_1 hold226 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_dout ),
    .X(net256));
 sg13g2_dlygate4sd3_1 hold227 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_dout ),
    .X(net257));
 sg13g2_dlygate4sd3_1 hold228 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[4] ),
    .X(net258));
 sg13g2_dlygate4sd3_1 hold229 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_dout ),
    .X(net259));
 sg13g2_dlygate4sd3_1 hold230 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_dout ),
    .X(net260));
 sg13g2_dlygate4sd3_1 hold231 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_dout ),
    .X(net261));
 sg13g2_dlygate4sd3_1 hold232 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_dout ),
    .X(net262));
 sg13g2_dlygate4sd3_1 hold233 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_dout ),
    .X(net263));
 sg13g2_dlygate4sd3_1 hold234 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_dout ),
    .X(net264));
 sg13g2_dlygate4sd3_1 hold235 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[4] ),
    .X(net265));
 sg13g2_dlygate4sd3_1 hold236 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[4] ),
    .X(net266));
 sg13g2_dlygate4sd3_1 hold237 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_dout ),
    .X(net267));
 sg13g2_dlygate4sd3_1 hold238 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_dout ),
    .X(net268));
 sg13g2_dlygate4sd3_1 hold239 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_dout ),
    .X(net269));
 sg13g2_dlygate4sd3_1 hold240 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_reg1 ),
    .X(net270));
 sg13g2_dlygate4sd3_1 hold241 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_dout ),
    .X(net271));
 sg13g2_dlygate4sd3_1 hold242 (.A(_01032_),
    .X(net272));
 sg13g2_dlygate4sd3_1 hold243 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_dout ),
    .X(net273));
 sg13g2_dlygate4sd3_1 hold244 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_dout ),
    .X(net274));
 sg13g2_dlygate4sd3_1 hold245 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[4] ),
    .X(net275));
 sg13g2_dlygate4sd3_1 hold246 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_dout ),
    .X(net276));
 sg13g2_dlygate4sd3_1 hold247 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_dout ),
    .X(net277));
 sg13g2_dlygate4sd3_1 hold248 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_dout ),
    .X(net278));
 sg13g2_dlygate4sd3_1 hold249 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_dout ),
    .X(net279));
 sg13g2_dlygate4sd3_1 hold250 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_dout ),
    .X(net280));
 sg13g2_dlygate4sd3_1 hold251 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.din ),
    .X(net281));
 sg13g2_dlygate4sd3_1 hold252 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[4] ),
    .X(net282));
 sg13g2_dlygate4sd3_1 hold253 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_dout ),
    .X(net283));
 sg13g2_dlygate4sd3_1 hold254 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_dout ),
    .X(net284));
 sg13g2_dlygate4sd3_1 hold255 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_dout ),
    .X(net285));
 sg13g2_dlygate4sd3_1 hold256 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_reg1 ),
    .X(net286));
 sg13g2_dlygate4sd3_1 hold257 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[4] ),
    .X(net287));
 sg13g2_dlygate4sd3_1 hold258 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_reg1 ),
    .X(net288));
 sg13g2_dlygate4sd3_1 hold259 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[1].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_dout ),
    .X(net289));
 sg13g2_dlygate4sd3_1 hold260 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_dout ),
    .X(net290));
 sg13g2_dlygate4sd3_1 hold261 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_dout ),
    .X(net291));
 sg13g2_dlygate4sd3_1 hold262 (.A(_00692_),
    .X(net292));
 sg13g2_dlygate4sd3_1 hold263 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[4] ),
    .X(net293));
 sg13g2_dlygate4sd3_1 hold264 (.A(\spiking_network_top_uut.debug_inst.debug_config[5] ),
    .X(net294));
 sg13g2_dlygate4sd3_1 hold265 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[4] ),
    .X(net295));
 sg13g2_dlygate4sd3_1 hold266 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_dout ),
    .X(net296));
 sg13g2_dlygate4sd3_1 hold267 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[4] ),
    .X(net297));
 sg13g2_dlygate4sd3_1 hold268 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[4] ),
    .X(net298));
 sg13g2_dlygate4sd3_1 hold269 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[1].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_dout ),
    .X(net299));
 sg13g2_dlygate4sd3_1 hold270 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_dout ),
    .X(net300));
 sg13g2_dlygate4sd3_1 hold271 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_dout ),
    .X(net301));
 sg13g2_dlygate4sd3_1 hold272 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[1].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_dout ),
    .X(net302));
 sg13g2_dlygate4sd3_1 hold273 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[0] ),
    .X(net303));
 sg13g2_dlygate4sd3_1 hold274 (.A(_00888_),
    .X(net304));
 sg13g2_dlygate4sd3_1 hold275 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_dout ),
    .X(net305));
 sg13g2_dlygate4sd3_1 hold276 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_dout ),
    .X(net306));
 sg13g2_dlygate4sd3_1 hold277 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_reg1 ),
    .X(net307));
 sg13g2_dlygate4sd3_1 hold278 (.A(_00982_),
    .X(net308));
 sg13g2_dlygate4sd3_1 hold279 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_dout ),
    .X(net309));
 sg13g2_dlygate4sd3_1 hold280 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_dout ),
    .X(net310));
 sg13g2_dlygate4sd3_1 hold281 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_dout ),
    .X(net311));
 sg13g2_dlygate4sd3_1 hold282 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[4] ),
    .X(net312));
 sg13g2_dlygate4sd3_1 hold283 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_dout ),
    .X(net313));
 sg13g2_dlygate4sd3_1 hold284 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_dout ),
    .X(net314));
 sg13g2_dlygate4sd3_1 hold285 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_dout ),
    .X(net315));
 sg13g2_dlygate4sd3_1 hold286 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[0] ),
    .X(net316));
 sg13g2_dlygate4sd3_1 hold287 (.A(_00609_),
    .X(net317));
 sg13g2_dlygate4sd3_1 hold288 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_dout ),
    .X(net318));
 sg13g2_dlygate4sd3_1 hold289 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_dout ),
    .X(net319));
 sg13g2_dlygate4sd3_1 hold290 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[0] ),
    .X(net320));
 sg13g2_dlygate4sd3_1 hold291 (.A(_00713_),
    .X(net321));
 sg13g2_dlygate4sd3_1 hold292 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_dout ),
    .X(net322));
 sg13g2_dlygate4sd3_1 hold293 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[1] ),
    .X(net323));
 sg13g2_dlygate4sd3_1 hold294 (.A(_00688_),
    .X(net324));
 sg13g2_dlygate4sd3_1 hold295 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[1].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_dout ),
    .X(net325));
 sg13g2_dlygate4sd3_1 hold296 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_dout ),
    .X(net326));
 sg13g2_dlygate4sd3_1 hold297 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_dout ),
    .X(net327));
 sg13g2_dlygate4sd3_1 hold298 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_dout ),
    .X(net328));
 sg13g2_dlygate4sd3_1 hold299 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[0] ),
    .X(net329));
 sg13g2_dlygate4sd3_1 hold300 (.A(_00940_),
    .X(net330));
 sg13g2_dlygate4sd3_1 hold301 (.A(_00054_),
    .X(net331));
 sg13g2_dlygate4sd3_1 hold302 (.A(_00583_),
    .X(net332));
 sg13g2_dlygate4sd3_1 hold303 (.A(_00066_),
    .X(net333));
 sg13g2_dlygate4sd3_1 hold304 (.A(_00635_),
    .X(net334));
 sg13g2_dlygate4sd3_1 hold305 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_dout ),
    .X(net335));
 sg13g2_dlygate4sd3_1 hold306 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_dout ),
    .X(net336));
 sg13g2_dlygate4sd3_1 hold307 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[0] ),
    .X(net337));
 sg13g2_dlygate4sd3_1 hold308 (.A(_00530_),
    .X(net338));
 sg13g2_dlygate4sd3_1 hold309 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[1] ),
    .X(net339));
 sg13g2_dlygate4sd3_1 hold310 (.A(_00126_),
    .X(net340));
 sg13g2_dlygate4sd3_1 hold311 (.A(_00966_),
    .X(net341));
 sg13g2_dlygate4sd3_1 hold312 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[1] ),
    .X(net342));
 sg13g2_dlygate4sd3_1 hold313 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[1] ),
    .X(net343));
 sg13g2_dlygate4sd3_1 hold314 (.A(_00636_),
    .X(net344));
 sg13g2_dlygate4sd3_1 hold315 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_dout ),
    .X(net345));
 sg13g2_dlygate4sd3_1 hold316 (.A(_00072_),
    .X(net346));
 sg13g2_dlygate4sd3_1 hold317 (.A(_00661_),
    .X(net347));
 sg13g2_dlygate4sd3_1 hold318 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[4] ),
    .X(net348));
 sg13g2_dlygate4sd3_1 hold319 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_reg1 ),
    .X(net349));
 sg13g2_dlygate4sd3_1 hold320 (.A(_00621_),
    .X(net350));
 sg13g2_dlygate4sd3_1 hold321 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[1] ),
    .X(net351));
 sg13g2_dlygate4sd3_1 hold322 (.A(_00448_),
    .X(net352));
 sg13g2_dlygate4sd3_1 hold323 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[0] ),
    .X(net353));
 sg13g2_dlygate4sd3_1 hold324 (.A(_00687_),
    .X(net354));
 sg13g2_dlygate4sd3_1 hold325 (.A(\spiking_network_top_uut.debug_inst.debug_config[7] ),
    .X(net355));
 sg13g2_dlygate4sd3_1 hold326 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_dout ),
    .X(net356));
 sg13g2_dlygate4sd3_1 hold327 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[0] ),
    .X(net357));
 sg13g2_dlygate4sd3_1 hold328 (.A(_00828_),
    .X(net358));
 sg13g2_dlygate4sd3_1 hold329 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[4] ),
    .X(net359));
 sg13g2_dlygate4sd3_1 hold330 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_dout ),
    .X(net360));
 sg13g2_dlygate4sd3_1 hold331 (.A(\spiking_network_top_uut.debug_inst.debug_config[4] ),
    .X(net361));
 sg13g2_dlygate4sd3_1 hold332 (.A(\spiking_network_top_uut.debug_inst.debug_config[6] ),
    .X(net362));
 sg13g2_dlygate4sd3_1 hold333 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[0] ),
    .X(net363));
 sg13g2_dlygate4sd3_1 hold334 (.A(_00992_),
    .X(net364));
 sg13g2_dlygate4sd3_1 hold335 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[0] ),
    .X(net365));
 sg13g2_dlygate4sd3_1 hold336 (.A(_00795_),
    .X(net366));
 sg13g2_dlygate4sd3_1 hold337 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[4] ),
    .X(net367));
 sg13g2_dlygate4sd3_1 hold338 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_dout ),
    .X(net368));
 sg13g2_dlygate4sd3_1 hold339 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_reg1 ),
    .X(net369));
 sg13g2_dlygate4sd3_1 hold340 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[1] ),
    .X(net370));
 sg13g2_dlygate4sd3_1 hold341 (.A(\spiking_network_top_uut.clk_div_inst.counter[2] ),
    .X(net371));
 sg13g2_dlygate4sd3_1 hold342 (.A(_03176_),
    .X(net372));
 sg13g2_dlygate4sd3_1 hold343 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_dout ),
    .X(net373));
 sg13g2_dlygate4sd3_1 hold344 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_dout ),
    .X(net374));
 sg13g2_dlygate4sd3_1 hold345 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[0] ),
    .X(net375));
 sg13g2_dlygate4sd3_1 hold346 (.A(_00556_),
    .X(net376));
 sg13g2_dlygate4sd3_1 hold347 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[0] ),
    .X(net377));
 sg13g2_dlygate4sd3_1 hold348 (.A(_00447_),
    .X(net378));
 sg13g2_dlygate4sd3_1 hold349 (.A(_00102_),
    .X(net379));
 sg13g2_dlygate4sd3_1 hold350 (.A(_00862_),
    .X(net380));
 sg13g2_dlygate4sd3_1 hold351 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[1] ),
    .X(net381));
 sg13g2_dlygate4sd3_1 hold352 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[1] ),
    .X(net382));
 sg13g2_dlygate4sd3_1 hold353 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_reg1 ),
    .X(net383));
 sg13g2_dlygate4sd3_1 hold354 (.A(_00683_),
    .X(net384));
 sg13g2_dlygate4sd3_1 hold355 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_reg1 ),
    .X(net385));
 sg13g2_dlygate4sd3_1 hold356 (.A(\spiking_network_top_uut.clk_div_inst.counter[3] ),
    .X(net386));
 sg13g2_dlygate4sd3_1 hold357 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[1] ),
    .X(net387));
 sg13g2_dlygate4sd3_1 hold358 (.A(_00967_),
    .X(net388));
 sg13g2_dlygate4sd3_1 hold359 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_reg1 ),
    .X(net389));
 sg13g2_dlygate4sd3_1 hold360 (.A(_00138_),
    .X(net390));
 sg13g2_dlygate4sd3_1 hold361 (.A(_01074_),
    .X(net391));
 sg13g2_dlygate4sd3_1 hold362 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[1] ),
    .X(net392));
 sg13g2_dlygate4sd3_1 hold363 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[1] ),
    .X(net393));
 sg13g2_dlygate4sd3_1 hold364 (.A(_00114_),
    .X(net394));
 sg13g2_dlygate4sd3_1 hold365 (.A(_00914_),
    .X(net395));
 sg13g2_dlygate4sd3_1 hold366 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[3] ),
    .X(net396));
 sg13g2_dlygate4sd3_1 hold367 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[1] ),
    .X(net397));
 sg13g2_dlygate4sd3_1 hold368 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[3] ),
    .X(net398));
 sg13g2_dlygate4sd3_1 hold369 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.din ),
    .X(net399));
 sg13g2_dlygate4sd3_1 hold370 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_dout ),
    .X(net400));
 sg13g2_dlygate4sd3_1 hold371 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[2] ),
    .X(net401));
 sg13g2_dlygate4sd3_1 hold372 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[1] ),
    .X(net402));
 sg13g2_dlygate4sd3_1 hold373 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[4] ),
    .X(net403));
 sg13g2_dlygate4sd3_1 hold374 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_reg1 ),
    .X(net404));
 sg13g2_dlygate4sd3_1 hold375 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_reg1 ),
    .X(net405));
 sg13g2_dlygate4sd3_1 hold376 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[3] ),
    .X(net406));
 sg13g2_dlygate4sd3_1 hold377 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[1] ),
    .X(net407));
 sg13g2_dlygate4sd3_1 hold378 (.A(_01075_),
    .X(net408));
 sg13g2_dlygate4sd3_1 hold379 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[1] ),
    .X(net409));
 sg13g2_dlygate4sd3_1 hold380 (.A(_00531_),
    .X(net410));
 sg13g2_dlygate4sd3_1 hold381 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_dout ),
    .X(net411));
 sg13g2_dlygate4sd3_1 hold382 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[1] ),
    .X(net412));
 sg13g2_dlygate4sd3_1 hold383 (.A(_00915_),
    .X(net413));
 sg13g2_dlygate4sd3_1 hold384 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[1] ),
    .X(net414));
 sg13g2_dlygate4sd3_1 hold385 (.A(_00610_),
    .X(net415));
 sg13g2_dlygate4sd3_1 hold386 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[3] ),
    .X(net416));
 sg13g2_dlygate4sd3_1 hold387 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[3] ),
    .X(net417));
 sg13g2_dlygate4sd3_1 hold388 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[0] ),
    .X(net418));
 sg13g2_dlygate4sd3_1 hold389 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[1] ),
    .X(net419));
 sg13g2_dlygate4sd3_1 hold390 (.A(_00662_),
    .X(net420));
 sg13g2_dlygate4sd3_1 hold391 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[3] ),
    .X(net421));
 sg13g2_dlygate4sd3_1 hold392 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[3] ),
    .X(net422));
 sg13g2_dlygate4sd3_1 hold393 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_dout ),
    .X(net423));
 sg13g2_dlygate4sd3_1 hold394 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_dout ),
    .X(net424));
 sg13g2_dlygate4sd3_1 hold395 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_dout ),
    .X(net425));
 sg13g2_dlygate4sd3_1 hold396 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[3] ),
    .X(net426));
 sg13g2_dlygate4sd3_1 hold397 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[3] ),
    .X(net427));
 sg13g2_dlygate4sd3_1 hold398 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[3] ),
    .X(net428));
 sg13g2_dlygate4sd3_1 hold399 (.A(\spiking_network_top_uut.clk_div_inst.counter[0] ),
    .X(net429));
 sg13g2_dlygate4sd3_1 hold400 (.A(_03172_),
    .X(net430));
 sg13g2_dlygate4sd3_1 hold401 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[3] ),
    .X(net431));
 sg13g2_dlygate4sd3_1 hold402 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_reg1 ),
    .X(net432));
 sg13g2_dlygate4sd3_1 hold403 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[3] ),
    .X(net433));
 sg13g2_dlygate4sd3_1 hold404 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[3] ),
    .X(net434));
 sg13g2_dlygate4sd3_1 hold405 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[2] ),
    .X(net435));
 sg13g2_dlygate4sd3_1 hold406 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[3] ),
    .X(net436));
 sg13g2_dlygate4sd3_1 hold407 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[1].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_dout ),
    .X(net437));
 sg13g2_dlygate4sd3_1 hold408 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[3] ),
    .X(net438));
 sg13g2_dlygate4sd3_1 hold409 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[3] ),
    .X(net439));
 sg13g2_dlygate4sd3_1 hold410 (.A(_00995_),
    .X(net440));
 sg13g2_dlygate4sd3_1 hold411 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[3] ),
    .X(net441));
 sg13g2_dlygate4sd3_1 hold412 (.A(_00798_),
    .X(net442));
 sg13g2_dlygate4sd3_1 hold413 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[3] ),
    .X(net443));
 sg13g2_dlygate4sd3_1 hold414 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_dout ),
    .X(net444));
 sg13g2_dlygate4sd3_1 hold415 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[0] ),
    .X(net445));
 sg13g2_dlygate4sd3_1 hold416 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_dout ),
    .X(net446));
 sg13g2_dlygate4sd3_1 hold417 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[0] ),
    .X(net447));
 sg13g2_dlygate4sd3_1 hold418 (.A(\spiking_network_top_uut.clk_div_inst.counter[4] ),
    .X(net448));
 sg13g2_dlygate4sd3_1 hold419 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ),
    .X(net449));
 sg13g2_dlygate4sd3_1 hold420 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ),
    .X(net450));
 sg13g2_dlygate4sd3_1 hold421 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[0] ),
    .X(net451));
 sg13g2_dlygate4sd3_1 hold422 (.A(\spiking_network_top_uut.clk_div_inst.counter[7] ),
    .X(net452));
 sg13g2_dlygate4sd3_1 hold423 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ),
    .X(net453));
 sg13g2_dlygate4sd3_1 hold424 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ),
    .X(net454));
 sg13g2_dlygate4sd3_1 hold425 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ),
    .X(net455));
 sg13g2_dlygate4sd3_1 hold426 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.enable_LYR_3 ),
    .X(net456));
 sg13g2_dlygate4sd3_1 hold427 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[0] ),
    .X(net457));
 sg13g2_dlygate4sd3_1 hold428 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_reg1 ),
    .X(net458));
 sg13g2_dlygate4sd3_1 hold429 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[0] ),
    .X(net459));
 sg13g2_dlygate4sd3_1 hold430 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ),
    .X(net460));
 sg13g2_dlygate4sd3_1 hold431 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ),
    .X(net461));
 sg13g2_dlygate4sd3_1 hold432 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_dout ),
    .X(net462));
 sg13g2_dlygate4sd3_1 hold433 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ),
    .X(net463));
 sg13g2_dlygate4sd3_1 hold434 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[0] ),
    .X(net464));
 sg13g2_dlygate4sd3_1 hold435 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[0] ),
    .X(net465));
 sg13g2_dlygate4sd3_1 hold436 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_dout ),
    .X(net466));
 sg13g2_dlygate4sd3_1 hold437 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[0] ),
    .X(net467));
 sg13g2_dlygate4sd3_1 hold438 (.A(\spiking_network_top_uut.clk_div_inst.counter[5] ),
    .X(net468));
 sg13g2_dlygate4sd3_1 hold439 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_dout ),
    .X(net469));
 sg13g2_dlygate4sd3_1 hold440 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_dout ),
    .X(net470));
 sg13g2_dlygate4sd3_1 hold441 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ),
    .X(net471));
 sg13g2_dlygate4sd3_1 hold442 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ),
    .X(net472));
 sg13g2_dlygate4sd3_1 hold443 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ),
    .X(net473));
 sg13g2_dlygate4sd3_1 hold444 (.A(\spiking_network_top_uut.clk_div_inst.counter[6] ),
    .X(net474));
 sg13g2_dlygate4sd3_1 hold445 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[0] ),
    .X(net475));
 sg13g2_dlygate4sd3_1 hold446 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_reg1 ),
    .X(net476));
 sg13g2_dlygate4sd3_1 hold447 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ),
    .X(net477));
 sg13g2_dlygate4sd3_1 hold448 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_dout ),
    .X(net478));
 sg13g2_dlygate4sd3_1 hold449 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_dout ),
    .X(net479));
 sg13g2_dlygate4sd3_1 hold450 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_dout ),
    .X(net480));
 sg13g2_dlygate4sd3_1 hold451 (.A(_00569_),
    .X(net481));
 sg13g2_dlygate4sd3_1 hold452 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ),
    .X(net482));
 sg13g2_dlygate4sd3_1 hold453 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ),
    .X(net483));
 sg13g2_dlygate4sd3_1 hold454 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[0] ),
    .X(net484));
 sg13g2_dlygate4sd3_1 hold455 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ),
    .X(net485));
 sg13g2_dlygate4sd3_1 hold456 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[0] ),
    .X(net486));
 sg13g2_dlygate4sd3_1 hold457 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ),
    .X(net487));
 sg13g2_dlygate4sd3_1 hold458 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ),
    .X(net488));
 sg13g2_dlygate4sd3_1 hold459 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ),
    .X(net489));
 sg13g2_dlygate4sd3_1 hold460 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ),
    .X(net490));
 sg13g2_dlygate4sd3_1 hold461 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[0] ),
    .X(net491));
 sg13g2_dlygate4sd3_1 hold462 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ),
    .X(net492));
 sg13g2_dlygate4sd3_1 hold463 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ),
    .X(net493));
 sg13g2_dlygate4sd3_1 hold464 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ),
    .X(net494));
 sg13g2_dlygate4sd3_1 hold465 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[0] ),
    .X(net495));
 sg13g2_dlygate4sd3_1 hold466 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[0] ),
    .X(net496));
 sg13g2_dlygate4sd3_1 hold467 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ),
    .X(net497));
 sg13g2_dlygate4sd3_1 hold468 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ),
    .X(net498));
 sg13g2_dlygate4sd3_1 hold469 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ),
    .X(net499));
 sg13g2_dlygate4sd3_1 hold470 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[0] ),
    .X(net500));
 sg13g2_dlygate4sd3_1 hold471 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ),
    .X(net501));
 sg13g2_dlygate4sd3_1 hold472 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ),
    .X(net502));
 sg13g2_dlygate4sd3_1 hold473 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ),
    .X(net503));
 sg13g2_dlygate4sd3_1 hold474 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ),
    .X(net504));
 sg13g2_dlygate4sd3_1 hold475 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ),
    .X(net505));
 sg13g2_dlygate4sd3_1 hold476 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[0] ),
    .X(net506));
 sg13g2_dlygate4sd3_1 hold477 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ),
    .X(net507));
 sg13g2_dlygate4sd3_1 hold478 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ),
    .X(net508));
 sg13g2_dlygate4sd3_1 hold479 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ),
    .X(net509));
 sg13g2_dlygate4sd3_1 hold480 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ),
    .X(net510));
 sg13g2_dlygate4sd3_1 hold481 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ),
    .X(net511));
 sg13g2_dlygate4sd3_1 hold482 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ),
    .X(net512));
 sg13g2_dlygate4sd3_1 hold483 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ),
    .X(net513));
 sg13g2_dlygate4sd3_1 hold484 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ),
    .X(net514));
 sg13g2_dlygate4sd3_1 hold485 (.A(\spiking_network_top_uut.debug_inst.debug_config[3] ),
    .X(net515));
 sg13g2_dlygate4sd3_1 hold486 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ),
    .X(net516));
 sg13g2_dlygate4sd3_1 hold487 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ),
    .X(net517));
 sg13g2_dlygate4sd3_1 hold488 (.A(\spiking_network_top_uut.debug_inst.debug_config[1] ),
    .X(net518));
 sg13g2_dlygate4sd3_1 hold489 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ),
    .X(net519));
 sg13g2_dlygate4sd3_1 hold490 (.A(\spiking_network_top_uut.debug_inst.debug_config[2] ),
    .X(net520));
 sg13g2_dlygate4sd3_1 hold491 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ),
    .X(net521));
 sg13g2_dlygate4sd3_1 hold492 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[0] ),
    .X(net522));
 sg13g2_dlygate4sd3_1 hold493 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ),
    .X(net523));
 sg13g2_dlygate4sd3_1 hold494 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_dout ),
    .X(net524));
 sg13g2_dlygate4sd3_1 hold495 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_dout ),
    .X(net525));
 sg13g2_dlygate4sd3_1 hold496 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ),
    .X(net526));
 sg13g2_dlygate4sd3_1 hold497 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_reg1 ),
    .X(net527));
 sg13g2_dlygate4sd3_1 hold498 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ),
    .X(net528));
 sg13g2_dlygate4sd3_1 hold499 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ),
    .X(net529));
 sg13g2_dlygate4sd3_1 hold500 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ),
    .X(net530));
 sg13g2_dlygate4sd3_1 hold501 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ),
    .X(net531));
 sg13g2_dlygate4sd3_1 hold502 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ),
    .X(net532));
 sg13g2_dlygate4sd3_1 hold503 (.A(\spiking_network_top_uut.debug_inst.debug_config[0] ),
    .X(net533));
 sg13g2_dlygate4sd3_1 hold504 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ),
    .X(net534));
 sg13g2_dlygate4sd3_1 hold505 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ),
    .X(net535));
 sg13g2_dlygate4sd3_1 hold506 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ),
    .X(net536));
 sg13g2_dlygate4sd3_1 hold507 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ),
    .X(net537));
 sg13g2_dlygate4sd3_1 hold508 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ),
    .X(net538));
 sg13g2_dlygate4sd3_1 hold509 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ),
    .X(net539));
 sg13g2_dlygate4sd3_1 hold510 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ),
    .X(net540));
 sg13g2_dlygate4sd3_1 hold511 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ),
    .X(net541));
 sg13g2_dlygate4sd3_1 hold512 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ),
    .X(net542));
 sg13g2_dlygate4sd3_1 hold513 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ),
    .X(net543));
 sg13g2_dlygate4sd3_1 hold514 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ),
    .X(net544));
 sg13g2_dlygate4sd3_1 hold515 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ),
    .X(net545));
 sg13g2_dlygate4sd3_1 hold516 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ),
    .X(net546));
 sg13g2_dlygate4sd3_1 hold517 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ),
    .X(net547));
 sg13g2_dlygate4sd3_1 hold518 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ),
    .X(net548));
 sg13g2_dlygate4sd3_1 hold519 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ),
    .X(net549));
 sg13g2_dlygate4sd3_1 hold520 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[1] ),
    .X(net550));
 sg13g2_dlygate4sd3_1 hold521 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[2] ),
    .X(net551));
 sg13g2_dlygate4sd3_1 hold522 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ),
    .X(net552));
 sg13g2_dlygate4sd3_1 hold523 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.enable_LYR_3 ),
    .X(net553));
 sg13g2_dlygate4sd3_1 hold524 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[1] ),
    .X(net554));
 sg13g2_dlygate4sd3_1 hold525 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer3.neuron_gen[1].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[0] ),
    .X(net555));
 sg13g2_dlygate4sd3_1 hold526 (.A(_05361_),
    .X(net556));
 sg13g2_dlygate4sd3_1 hold527 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.lif_neuron_inst.lif_neuron_inst.refractory_counter[1] ),
    .X(net557));
 sg13g2_antennanp ANTENNA_1 (.A(_00026_));
 sg13g2_antennanp ANTENNA_2 (.A(_00026_));
 sg13g2_antennanp ANTENNA_3 (.A(_00026_));
 sg13g2_antennanp ANTENNA_4 (.A(_00026_));
 sg13g2_antennanp ANTENNA_5 (.A(_00026_));
 sg13g2_antennanp ANTENNA_6 (.A(_00026_));
 sg13g2_antennanp ANTENNA_7 (.A(_00146_));
 sg13g2_antennanp ANTENNA_8 (.A(_00158_));
 sg13g2_antennanp ANTENNA_9 (.A(_00164_));
 sg13g2_antennanp ANTENNA_10 (.A(_00188_));
 sg13g2_antennanp ANTENNA_11 (.A(_00197_));
 sg13g2_antennanp ANTENNA_12 (.A(_00201_));
 sg13g2_antennanp ANTENNA_13 (.A(_00209_));
 sg13g2_antennanp ANTENNA_14 (.A(_00213_));
 sg13g2_antennanp ANTENNA_15 (.A(_00217_));
 sg13g2_antennanp ANTENNA_16 (.A(_00226_));
 sg13g2_antennanp ANTENNA_17 (.A(_00232_));
 sg13g2_antennanp ANTENNA_18 (.A(_00251_));
 sg13g2_antennanp ANTENNA_19 (.A(_00258_));
 sg13g2_antennanp ANTENNA_20 (.A(_00271_));
 sg13g2_antennanp ANTENNA_21 (.A(_00283_));
 sg13g2_antennanp ANTENNA_22 (.A(_00284_));
 sg13g2_antennanp ANTENNA_23 (.A(_00288_));
 sg13g2_antennanp ANTENNA_24 (.A(_00299_));
 sg13g2_antennanp ANTENNA_25 (.A(_00343_));
 sg13g2_antennanp ANTENNA_26 (.A(_00347_));
 sg13g2_antennanp ANTENNA_27 (.A(_00349_));
 sg13g2_antennanp ANTENNA_28 (.A(_00390_));
 sg13g2_antennanp ANTENNA_29 (.A(_00391_));
 sg13g2_antennanp ANTENNA_30 (.A(_00415_));
 sg13g2_antennanp ANTENNA_31 (.A(_00419_));
 sg13g2_antennanp ANTENNA_32 (.A(_02122_));
 sg13g2_antennanp ANTENNA_33 (.A(_02122_));
 sg13g2_antennanp ANTENNA_34 (.A(_02122_));
 sg13g2_antennanp ANTENNA_35 (.A(_02122_));
 sg13g2_antennanp ANTENNA_36 (.A(_02215_));
 sg13g2_antennanp ANTENNA_37 (.A(_02216_));
 sg13g2_antennanp ANTENNA_38 (.A(_02405_));
 sg13g2_antennanp ANTENNA_39 (.A(_02405_));
 sg13g2_antennanp ANTENNA_40 (.A(_02405_));
 sg13g2_antennanp ANTENNA_41 (.A(_02405_));
 sg13g2_antennanp ANTENNA_42 (.A(_02405_));
 sg13g2_antennanp ANTENNA_43 (.A(_02405_));
 sg13g2_antennanp ANTENNA_44 (.A(_02405_));
 sg13g2_antennanp ANTENNA_45 (.A(_02405_));
 sg13g2_antennanp ANTENNA_46 (.A(_02405_));
 sg13g2_antennanp ANTENNA_47 (.A(_02405_));
 sg13g2_antennanp ANTENNA_48 (.A(_02405_));
 sg13g2_antennanp ANTENNA_49 (.A(_02405_));
 sg13g2_antennanp ANTENNA_50 (.A(_02405_));
 sg13g2_antennanp ANTENNA_51 (.A(_02405_));
 sg13g2_antennanp ANTENNA_52 (.A(_02405_));
 sg13g2_antennanp ANTENNA_53 (.A(_02405_));
 sg13g2_antennanp ANTENNA_54 (.A(_02405_));
 sg13g2_antennanp ANTENNA_55 (.A(_02405_));
 sg13g2_antennanp ANTENNA_56 (.A(_02406_));
 sg13g2_antennanp ANTENNA_57 (.A(_02406_));
 sg13g2_antennanp ANTENNA_58 (.A(_02406_));
 sg13g2_antennanp ANTENNA_59 (.A(_02406_));
 sg13g2_antennanp ANTENNA_60 (.A(_02438_));
 sg13g2_antennanp ANTENNA_61 (.A(_02438_));
 sg13g2_antennanp ANTENNA_62 (.A(_02438_));
 sg13g2_antennanp ANTENNA_63 (.A(_02438_));
 sg13g2_antennanp ANTENNA_64 (.A(_02483_));
 sg13g2_antennanp ANTENNA_65 (.A(_02483_));
 sg13g2_antennanp ANTENNA_66 (.A(_02483_));
 sg13g2_antennanp ANTENNA_67 (.A(_02483_));
 sg13g2_antennanp ANTENNA_68 (.A(_02483_));
 sg13g2_antennanp ANTENNA_69 (.A(_02483_));
 sg13g2_antennanp ANTENNA_70 (.A(_02483_));
 sg13g2_antennanp ANTENNA_71 (.A(_02483_));
 sg13g2_antennanp ANTENNA_72 (.A(_02483_));
 sg13g2_antennanp ANTENNA_73 (.A(_02484_));
 sg13g2_antennanp ANTENNA_74 (.A(_02484_));
 sg13g2_antennanp ANTENNA_75 (.A(_02484_));
 sg13g2_antennanp ANTENNA_76 (.A(_02484_));
 sg13g2_antennanp ANTENNA_77 (.A(_02494_));
 sg13g2_antennanp ANTENNA_78 (.A(_02494_));
 sg13g2_antennanp ANTENNA_79 (.A(_02494_));
 sg13g2_antennanp ANTENNA_80 (.A(_02494_));
 sg13g2_antennanp ANTENNA_81 (.A(_02495_));
 sg13g2_antennanp ANTENNA_82 (.A(_02495_));
 sg13g2_antennanp ANTENNA_83 (.A(_02495_));
 sg13g2_antennanp ANTENNA_84 (.A(_02495_));
 sg13g2_antennanp ANTENNA_85 (.A(_02495_));
 sg13g2_antennanp ANTENNA_86 (.A(_02495_));
 sg13g2_antennanp ANTENNA_87 (.A(_02495_));
 sg13g2_antennanp ANTENNA_88 (.A(_02495_));
 sg13g2_antennanp ANTENNA_89 (.A(_02495_));
 sg13g2_antennanp ANTENNA_90 (.A(_02509_));
 sg13g2_antennanp ANTENNA_91 (.A(_02509_));
 sg13g2_antennanp ANTENNA_92 (.A(_02509_));
 sg13g2_antennanp ANTENNA_93 (.A(_02509_));
 sg13g2_antennanp ANTENNA_94 (.A(_02700_));
 sg13g2_antennanp ANTENNA_95 (.A(_02700_));
 sg13g2_antennanp ANTENNA_96 (.A(_02700_));
 sg13g2_antennanp ANTENNA_97 (.A(_02700_));
 sg13g2_antennanp ANTENNA_98 (.A(_02700_));
 sg13g2_antennanp ANTENNA_99 (.A(_02700_));
 sg13g2_antennanp ANTENNA_100 (.A(_02700_));
 sg13g2_antennanp ANTENNA_101 (.A(_02700_));
 sg13g2_antennanp ANTENNA_102 (.A(_02700_));
 sg13g2_antennanp ANTENNA_103 (.A(_02700_));
 sg13g2_antennanp ANTENNA_104 (.A(_02700_));
 sg13g2_antennanp ANTENNA_105 (.A(_02700_));
 sg13g2_antennanp ANTENNA_106 (.A(_02777_));
 sg13g2_antennanp ANTENNA_107 (.A(_02777_));
 sg13g2_antennanp ANTENNA_108 (.A(_02777_));
 sg13g2_antennanp ANTENNA_109 (.A(_02777_));
 sg13g2_antennanp ANTENNA_110 (.A(_02785_));
 sg13g2_antennanp ANTENNA_111 (.A(_02991_));
 sg13g2_antennanp ANTENNA_112 (.A(_02991_));
 sg13g2_antennanp ANTENNA_113 (.A(_02991_));
 sg13g2_antennanp ANTENNA_114 (.A(_02991_));
 sg13g2_antennanp ANTENNA_115 (.A(_02991_));
 sg13g2_antennanp ANTENNA_116 (.A(_02991_));
 sg13g2_antennanp ANTENNA_117 (.A(_02991_));
 sg13g2_antennanp ANTENNA_118 (.A(_02991_));
 sg13g2_antennanp ANTENNA_119 (.A(_02991_));
 sg13g2_antennanp ANTENNA_120 (.A(_03509_));
 sg13g2_antennanp ANTENNA_121 (.A(_03518_));
 sg13g2_antennanp ANTENNA_122 (.A(_03522_));
 sg13g2_antennanp ANTENNA_123 (.A(_03526_));
 sg13g2_antennanp ANTENNA_124 (.A(_03534_));
 sg13g2_antennanp ANTENNA_125 (.A(_03536_));
 sg13g2_antennanp ANTENNA_126 (.A(_03537_));
 sg13g2_antennanp ANTENNA_127 (.A(_03543_));
 sg13g2_antennanp ANTENNA_128 (.A(_03549_));
 sg13g2_antennanp ANTENNA_129 (.A(_03550_));
 sg13g2_antennanp ANTENNA_130 (.A(_03551_));
 sg13g2_antennanp ANTENNA_131 (.A(_03560_));
 sg13g2_antennanp ANTENNA_132 (.A(_03567_));
 sg13g2_antennanp ANTENNA_133 (.A(_03571_));
 sg13g2_antennanp ANTENNA_134 (.A(_03573_));
 sg13g2_antennanp ANTENNA_135 (.A(_03574_));
 sg13g2_antennanp ANTENNA_136 (.A(_03576_));
 sg13g2_antennanp ANTENNA_137 (.A(_03578_));
 sg13g2_antennanp ANTENNA_138 (.A(_03589_));
 sg13g2_antennanp ANTENNA_139 (.A(_03602_));
 sg13g2_antennanp ANTENNA_140 (.A(_03609_));
 sg13g2_antennanp ANTENNA_141 (.A(_03613_));
 sg13g2_antennanp ANTENNA_142 (.A(_03614_));
 sg13g2_antennanp ANTENNA_143 (.A(_03622_));
 sg13g2_antennanp ANTENNA_144 (.A(_03625_));
 sg13g2_antennanp ANTENNA_145 (.A(_03629_));
 sg13g2_antennanp ANTENNA_146 (.A(_03631_));
 sg13g2_antennanp ANTENNA_147 (.A(_03633_));
 sg13g2_antennanp ANTENNA_148 (.A(_03648_));
 sg13g2_antennanp ANTENNA_149 (.A(_03650_));
 sg13g2_antennanp ANTENNA_150 (.A(_03651_));
 sg13g2_antennanp ANTENNA_151 (.A(_03652_));
 sg13g2_antennanp ANTENNA_152 (.A(_03654_));
 sg13g2_antennanp ANTENNA_153 (.A(_03794_));
 sg13g2_antennanp ANTENNA_154 (.A(_03794_));
 sg13g2_antennanp ANTENNA_155 (.A(_03794_));
 sg13g2_antennanp ANTENNA_156 (.A(_03794_));
 sg13g2_antennanp ANTENNA_157 (.A(_03794_));
 sg13g2_antennanp ANTENNA_158 (.A(_03794_));
 sg13g2_antennanp ANTENNA_159 (.A(_03794_));
 sg13g2_antennanp ANTENNA_160 (.A(_03794_));
 sg13g2_antennanp ANTENNA_161 (.A(_03794_));
 sg13g2_antennanp ANTENNA_162 (.A(_03794_));
 sg13g2_antennanp ANTENNA_163 (.A(_03794_));
 sg13g2_antennanp ANTENNA_164 (.A(_03794_));
 sg13g2_antennanp ANTENNA_165 (.A(_03794_));
 sg13g2_antennanp ANTENNA_166 (.A(_03794_));
 sg13g2_antennanp ANTENNA_167 (.A(_03794_));
 sg13g2_antennanp ANTENNA_168 (.A(_03794_));
 sg13g2_antennanp ANTENNA_169 (.A(_03794_));
 sg13g2_antennanp ANTENNA_170 (.A(_03794_));
 sg13g2_antennanp ANTENNA_171 (.A(_03794_));
 sg13g2_antennanp ANTENNA_172 (.A(_03794_));
 sg13g2_antennanp ANTENNA_173 (.A(_03858_));
 sg13g2_antennanp ANTENNA_174 (.A(_03893_));
 sg13g2_antennanp ANTENNA_175 (.A(_03906_));
 sg13g2_antennanp ANTENNA_176 (.A(_03913_));
 sg13g2_antennanp ANTENNA_177 (.A(_03981_));
 sg13g2_antennanp ANTENNA_178 (.A(_03988_));
 sg13g2_antennanp ANTENNA_179 (.A(_03990_));
 sg13g2_antennanp ANTENNA_180 (.A(_03993_));
 sg13g2_antennanp ANTENNA_181 (.A(_03999_));
 sg13g2_antennanp ANTENNA_182 (.A(_04005_));
 sg13g2_antennanp ANTENNA_183 (.A(_04025_));
 sg13g2_antennanp ANTENNA_184 (.A(_04028_));
 sg13g2_antennanp ANTENNA_185 (.A(_04043_));
 sg13g2_antennanp ANTENNA_186 (.A(_04046_));
 sg13g2_antennanp ANTENNA_187 (.A(_04081_));
 sg13g2_antennanp ANTENNA_188 (.A(_04092_));
 sg13g2_antennanp ANTENNA_189 (.A(_04103_));
 sg13g2_antennanp ANTENNA_190 (.A(_04114_));
 sg13g2_antennanp ANTENNA_191 (.A(_04119_));
 sg13g2_antennanp ANTENNA_192 (.A(_04130_));
 sg13g2_antennanp ANTENNA_193 (.A(_04131_));
 sg13g2_antennanp ANTENNA_194 (.A(_04132_));
 sg13g2_antennanp ANTENNA_195 (.A(_04137_));
 sg13g2_antennanp ANTENNA_196 (.A(_04145_));
 sg13g2_antennanp ANTENNA_197 (.A(_04148_));
 sg13g2_antennanp ANTENNA_198 (.A(_04157_));
 sg13g2_antennanp ANTENNA_199 (.A(_04167_));
 sg13g2_antennanp ANTENNA_200 (.A(_04186_));
 sg13g2_antennanp ANTENNA_201 (.A(_04191_));
 sg13g2_antennanp ANTENNA_202 (.A(_04194_));
 sg13g2_antennanp ANTENNA_203 (.A(_04202_));
 sg13g2_antennanp ANTENNA_204 (.A(_04213_));
 sg13g2_antennanp ANTENNA_205 (.A(_04216_));
 sg13g2_antennanp ANTENNA_206 (.A(_04221_));
 sg13g2_antennanp ANTENNA_207 (.A(_04231_));
 sg13g2_antennanp ANTENNA_208 (.A(_04238_));
 sg13g2_antennanp ANTENNA_209 (.A(_04243_));
 sg13g2_antennanp ANTENNA_210 (.A(_04267_));
 sg13g2_antennanp ANTENNA_211 (.A(_04270_));
 sg13g2_antennanp ANTENNA_212 (.A(_04271_));
 sg13g2_antennanp ANTENNA_213 (.A(_04280_));
 sg13g2_antennanp ANTENNA_214 (.A(_04289_));
 sg13g2_antennanp ANTENNA_215 (.A(_04301_));
 sg13g2_antennanp ANTENNA_216 (.A(_04312_));
 sg13g2_antennanp ANTENNA_217 (.A(_04319_));
 sg13g2_antennanp ANTENNA_218 (.A(_04337_));
 sg13g2_antennanp ANTENNA_219 (.A(_04352_));
 sg13g2_antennanp ANTENNA_220 (.A(_04362_));
 sg13g2_antennanp ANTENNA_221 (.A(_04374_));
 sg13g2_antennanp ANTENNA_222 (.A(_04401_));
 sg13g2_antennanp ANTENNA_223 (.A(_04403_));
 sg13g2_antennanp ANTENNA_224 (.A(_04410_));
 sg13g2_antennanp ANTENNA_225 (.A(_04415_));
 sg13g2_antennanp ANTENNA_226 (.A(_04417_));
 sg13g2_antennanp ANTENNA_227 (.A(_04436_));
 sg13g2_antennanp ANTENNA_228 (.A(_04450_));
 sg13g2_antennanp ANTENNA_229 (.A(_04480_));
 sg13g2_antennanp ANTENNA_230 (.A(_04498_));
 sg13g2_antennanp ANTENNA_231 (.A(_04500_));
 sg13g2_antennanp ANTENNA_232 (.A(_04504_));
 sg13g2_antennanp ANTENNA_233 (.A(_04508_));
 sg13g2_antennanp ANTENNA_234 (.A(_04511_));
 sg13g2_antennanp ANTENNA_235 (.A(_04514_));
 sg13g2_antennanp ANTENNA_236 (.A(_04523_));
 sg13g2_antennanp ANTENNA_237 (.A(_04546_));
 sg13g2_antennanp ANTENNA_238 (.A(_04556_));
 sg13g2_antennanp ANTENNA_239 (.A(_04559_));
 sg13g2_antennanp ANTENNA_240 (.A(_04562_));
 sg13g2_antennanp ANTENNA_241 (.A(_04578_));
 sg13g2_antennanp ANTENNA_242 (.A(_04579_));
 sg13g2_antennanp ANTENNA_243 (.A(_04580_));
 sg13g2_antennanp ANTENNA_244 (.A(_04584_));
 sg13g2_antennanp ANTENNA_245 (.A(_05709_));
 sg13g2_antennanp ANTENNA_246 (.A(_05709_));
 sg13g2_antennanp ANTENNA_247 (.A(_05709_));
 sg13g2_antennanp ANTENNA_248 (.A(_05709_));
 sg13g2_antennanp ANTENNA_249 (.A(_05804_));
 sg13g2_antennanp ANTENNA_250 (.A(_05805_));
 sg13g2_antennanp ANTENNA_251 (.A(_05995_));
 sg13g2_antennanp ANTENNA_252 (.A(_05995_));
 sg13g2_antennanp ANTENNA_253 (.A(_05995_));
 sg13g2_antennanp ANTENNA_254 (.A(_05995_));
 sg13g2_antennanp ANTENNA_255 (.A(_06082_));
 sg13g2_antennanp ANTENNA_256 (.A(_06284_));
 sg13g2_antennanp ANTENNA_257 (.A(_06284_));
 sg13g2_antennanp ANTENNA_258 (.A(_06284_));
 sg13g2_antennanp ANTENNA_259 (.A(_06284_));
 sg13g2_antennanp ANTENNA_260 (.A(_06286_));
 sg13g2_antennanp ANTENNA_261 (.A(_06286_));
 sg13g2_antennanp ANTENNA_262 (.A(_06286_));
 sg13g2_antennanp ANTENNA_263 (.A(_06286_));
 sg13g2_antennanp ANTENNA_264 (.A(_06625_));
 sg13g2_antennanp ANTENNA_265 (.A(_06625_));
 sg13g2_antennanp ANTENNA_266 (.A(_06625_));
 sg13g2_antennanp ANTENNA_267 (.A(_06625_));
 sg13g2_antennanp ANTENNA_268 (.A(_06679_));
 sg13g2_antennanp ANTENNA_269 (.A(_06679_));
 sg13g2_antennanp ANTENNA_270 (.A(_06679_));
 sg13g2_antennanp ANTENNA_271 (.A(_06679_));
 sg13g2_antennanp ANTENNA_272 (.A(_07526_));
 sg13g2_antennanp ANTENNA_273 (.A(_07721_));
 sg13g2_antennanp ANTENNA_274 (.A(_07721_));
 sg13g2_antennanp ANTENNA_275 (.A(_07721_));
 sg13g2_antennanp ANTENNA_276 (.A(_07721_));
 sg13g2_antennanp ANTENNA_277 (.A(_08106_));
 sg13g2_antennanp ANTENNA_278 (.A(_08106_));
 sg13g2_antennanp ANTENNA_279 (.A(_08106_));
 sg13g2_antennanp ANTENNA_280 (.A(_08106_));
 sg13g2_antennanp ANTENNA_281 (.A(_08570_));
 sg13g2_antennanp ANTENNA_282 (.A(_08570_));
 sg13g2_antennanp ANTENNA_283 (.A(_08570_));
 sg13g2_antennanp ANTENNA_284 (.A(_08570_));
 sg13g2_antennanp ANTENNA_285 (.A(_08572_));
 sg13g2_antennanp ANTENNA_286 (.A(_08572_));
 sg13g2_antennanp ANTENNA_287 (.A(_08572_));
 sg13g2_antennanp ANTENNA_288 (.A(_08572_));
 sg13g2_antennanp ANTENNA_289 (.A(_08849_));
 sg13g2_antennanp ANTENNA_290 (.A(_08849_));
 sg13g2_antennanp ANTENNA_291 (.A(_08849_));
 sg13g2_antennanp ANTENNA_292 (.A(_08849_));
 sg13g2_antennanp ANTENNA_293 (.A(_08849_));
 sg13g2_antennanp ANTENNA_294 (.A(_08849_));
 sg13g2_antennanp ANTENNA_295 (.A(_08849_));
 sg13g2_antennanp ANTENNA_296 (.A(_08849_));
 sg13g2_antennanp ANTENNA_297 (.A(_08849_));
 sg13g2_antennanp ANTENNA_298 (.A(_08851_));
 sg13g2_antennanp ANTENNA_299 (.A(_08851_));
 sg13g2_antennanp ANTENNA_300 (.A(_08851_));
 sg13g2_antennanp ANTENNA_301 (.A(_08851_));
 sg13g2_antennanp ANTENNA_302 (.A(_08851_));
 sg13g2_antennanp ANTENNA_303 (.A(_08851_));
 sg13g2_antennanp ANTENNA_304 (.A(_08851_));
 sg13g2_antennanp ANTENNA_305 (.A(_08851_));
 sg13g2_antennanp ANTENNA_306 (.A(_08851_));
 sg13g2_antennanp ANTENNA_307 (.A(_08860_));
 sg13g2_antennanp ANTENNA_308 (.A(_08860_));
 sg13g2_antennanp ANTENNA_309 (.A(_08860_));
 sg13g2_antennanp ANTENNA_310 (.A(_08860_));
 sg13g2_antennanp ANTENNA_311 (.A(\spiking_network_top_uut.all_data_out[17] ));
 sg13g2_antennanp ANTENNA_312 (.A(\spiking_network_top_uut.all_data_out[17] ));
 sg13g2_antennanp ANTENNA_313 (.A(\spiking_network_top_uut.all_data_out[17] ));
 sg13g2_antennanp ANTENNA_314 (.A(\spiking_network_top_uut.all_data_out[17] ));
 sg13g2_antennanp ANTENNA_315 (.A(\spiking_network_top_uut.all_data_out[273] ));
 sg13g2_antennanp ANTENNA_316 (.A(\spiking_network_top_uut.all_data_out[273] ));
 sg13g2_antennanp ANTENNA_317 (.A(\spiking_network_top_uut.all_data_out[273] ));
 sg13g2_antennanp ANTENNA_318 (.A(\spiking_network_top_uut.all_data_out[291] ));
 sg13g2_antennanp ANTENNA_319 (.A(\spiking_network_top_uut.all_data_out[291] ));
 sg13g2_antennanp ANTENNA_320 (.A(\spiking_network_top_uut.all_data_out[291] ));
 sg13g2_antennanp ANTENNA_321 (.A(\spiking_network_top_uut.all_data_out[291] ));
 sg13g2_antennanp ANTENNA_322 (.A(\spiking_network_top_uut.all_data_out[291] ));
 sg13g2_antennanp ANTENNA_323 (.A(\spiking_network_top_uut.all_data_out[291] ));
 sg13g2_antennanp ANTENNA_324 (.A(\spiking_network_top_uut.all_data_out[294] ));
 sg13g2_antennanp ANTENNA_325 (.A(\spiking_network_top_uut.all_data_out[294] ));
 sg13g2_antennanp ANTENNA_326 (.A(\spiking_network_top_uut.all_data_out[294] ));
 sg13g2_antennanp ANTENNA_327 (.A(\spiking_network_top_uut.all_data_out[294] ));
 sg13g2_antennanp ANTENNA_328 (.A(\spiking_network_top_uut.all_data_out[294] ));
 sg13g2_antennanp ANTENNA_329 (.A(\spiking_network_top_uut.all_data_out[294] ));
 sg13g2_antennanp ANTENNA_330 (.A(\spiking_network_top_uut.all_data_out[294] ));
 sg13g2_antennanp ANTENNA_331 (.A(\spiking_network_top_uut.all_data_out[294] ));
 sg13g2_antennanp ANTENNA_332 (.A(\spiking_network_top_uut.all_data_out[294] ));
 sg13g2_antennanp ANTENNA_333 (.A(\spiking_network_top_uut.all_data_out[295] ));
 sg13g2_antennanp ANTENNA_334 (.A(\spiking_network_top_uut.all_data_out[295] ));
 sg13g2_antennanp ANTENNA_335 (.A(\spiking_network_top_uut.all_data_out[295] ));
 sg13g2_antennanp ANTENNA_336 (.A(\spiking_network_top_uut.all_data_out[299] ));
 sg13g2_antennanp ANTENNA_337 (.A(\spiking_network_top_uut.all_data_out[299] ));
 sg13g2_antennanp ANTENNA_338 (.A(\spiking_network_top_uut.all_data_out[299] ));
 sg13g2_antennanp ANTENNA_339 (.A(\spiking_network_top_uut.all_data_out[299] ));
 sg13g2_antennanp ANTENNA_340 (.A(\spiking_network_top_uut.all_data_out[299] ));
 sg13g2_antennanp ANTENNA_341 (.A(\spiking_network_top_uut.all_data_out[307] ));
 sg13g2_antennanp ANTENNA_342 (.A(\spiking_network_top_uut.all_data_out[307] ));
 sg13g2_antennanp ANTENNA_343 (.A(\spiking_network_top_uut.all_data_out[307] ));
 sg13g2_antennanp ANTENNA_344 (.A(\spiking_network_top_uut.all_data_out[308] ));
 sg13g2_antennanp ANTENNA_345 (.A(\spiking_network_top_uut.all_data_out[308] ));
 sg13g2_antennanp ANTENNA_346 (.A(\spiking_network_top_uut.all_data_out[308] ));
 sg13g2_antennanp ANTENNA_347 (.A(\spiking_network_top_uut.all_data_out[308] ));
 sg13g2_antennanp ANTENNA_348 (.A(\spiking_network_top_uut.all_data_out[311] ));
 sg13g2_antennanp ANTENNA_349 (.A(\spiking_network_top_uut.all_data_out[311] ));
 sg13g2_antennanp ANTENNA_350 (.A(\spiking_network_top_uut.all_data_out[311] ));
 sg13g2_antennanp ANTENNA_351 (.A(\spiking_network_top_uut.all_data_out[330] ));
 sg13g2_antennanp ANTENNA_352 (.A(\spiking_network_top_uut.all_data_out[330] ));
 sg13g2_antennanp ANTENNA_353 (.A(\spiking_network_top_uut.all_data_out[330] ));
 sg13g2_antennanp ANTENNA_354 (.A(\spiking_network_top_uut.all_data_out[330] ));
 sg13g2_antennanp ANTENNA_355 (.A(\spiking_network_top_uut.all_data_out[392] ));
 sg13g2_antennanp ANTENNA_356 (.A(\spiking_network_top_uut.all_data_out[392] ));
 sg13g2_antennanp ANTENNA_357 (.A(\spiking_network_top_uut.all_data_out[392] ));
 sg13g2_antennanp ANTENNA_358 (.A(\spiking_network_top_uut.all_data_out[392] ));
 sg13g2_antennanp ANTENNA_359 (.A(\spiking_network_top_uut.all_data_out[392] ));
 sg13g2_antennanp ANTENNA_360 (.A(\spiking_network_top_uut.all_data_out[392] ));
 sg13g2_antennanp ANTENNA_361 (.A(\spiking_network_top_uut.all_data_out[392] ));
 sg13g2_antennanp ANTENNA_362 (.A(\spiking_network_top_uut.all_data_out[392] ));
 sg13g2_antennanp ANTENNA_363 (.A(\spiking_network_top_uut.all_data_out[516] ));
 sg13g2_antennanp ANTENNA_364 (.A(\spiking_network_top_uut.all_data_out[516] ));
 sg13g2_antennanp ANTENNA_365 (.A(\spiking_network_top_uut.all_data_out[516] ));
 sg13g2_antennanp ANTENNA_366 (.A(\spiking_network_top_uut.all_data_out[516] ));
 sg13g2_antennanp ANTENNA_367 (.A(\spiking_network_top_uut.all_data_out[516] ));
 sg13g2_antennanp ANTENNA_368 (.A(\spiking_network_top_uut.all_data_out[516] ));
 sg13g2_antennanp ANTENNA_369 (.A(\spiking_network_top_uut.all_data_out[516] ));
 sg13g2_antennanp ANTENNA_370 (.A(\spiking_network_top_uut.all_data_out[516] ));
 sg13g2_antennanp ANTENNA_371 (.A(\spiking_network_top_uut.all_data_out[584] ));
 sg13g2_antennanp ANTENNA_372 (.A(\spiking_network_top_uut.all_data_out[584] ));
 sg13g2_antennanp ANTENNA_373 (.A(\spiking_network_top_uut.all_data_out[584] ));
 sg13g2_antennanp ANTENNA_374 (.A(\spiking_network_top_uut.all_data_out[584] ));
 sg13g2_antennanp ANTENNA_375 (.A(\spiking_network_top_uut.all_data_out[584] ));
 sg13g2_antennanp ANTENNA_376 (.A(\spiking_network_top_uut.all_data_out[584] ));
 sg13g2_antennanp ANTENNA_377 (.A(\spiking_network_top_uut.all_data_out[584] ));
 sg13g2_antennanp ANTENNA_378 (.A(\spiking_network_top_uut.all_data_out[584] ));
 sg13g2_antennanp ANTENNA_379 (.A(\spiking_network_top_uut.all_data_out[587] ));
 sg13g2_antennanp ANTENNA_380 (.A(\spiking_network_top_uut.all_data_out[587] ));
 sg13g2_antennanp ANTENNA_381 (.A(\spiking_network_top_uut.all_data_out[587] ));
 sg13g2_antennanp ANTENNA_382 (.A(\spiking_network_top_uut.all_data_out[587] ));
 sg13g2_antennanp ANTENNA_383 (.A(\spiking_network_top_uut.all_data_out[587] ));
 sg13g2_antennanp ANTENNA_384 (.A(\spiking_network_top_uut.all_data_out[76] ));
 sg13g2_antennanp ANTENNA_385 (.A(\spiking_network_top_uut.all_data_out[76] ));
 sg13g2_antennanp ANTENNA_386 (.A(\spiking_network_top_uut.all_data_out[76] ));
 sg13g2_antennanp ANTENNA_387 (.A(\spiking_network_top_uut.all_data_out[76] ));
 sg13g2_antennanp ANTENNA_388 (.A(\spiking_network_top_uut.all_data_out[79] ));
 sg13g2_antennanp ANTENNA_389 (.A(\spiking_network_top_uut.all_data_out[79] ));
 sg13g2_antennanp ANTENNA_390 (.A(\spiking_network_top_uut.all_data_out[79] ));
 sg13g2_antennanp ANTENNA_391 (.A(\spiking_network_top_uut.all_data_out[79] ));
 sg13g2_antennanp ANTENNA_392 (.A(\spiking_network_top_uut.all_data_out[79] ));
 sg13g2_antennanp ANTENNA_393 (.A(\spiking_network_top_uut.all_data_out[79] ));
 sg13g2_antennanp ANTENNA_394 (.A(\spiking_network_top_uut.all_data_out[79] ));
 sg13g2_antennanp ANTENNA_395 (.A(\spiking_network_top_uut.all_data_out[79] ));
 sg13g2_antennanp ANTENNA_396 (.A(\spiking_network_top_uut.all_data_out[79] ));
 sg13g2_antennanp ANTENNA_397 (.A(\spiking_network_top_uut.all_data_out[79] ));
 sg13g2_antennanp ANTENNA_398 (.A(\spiking_network_top_uut.all_data_out[79] ));
 sg13g2_antennanp ANTENNA_399 (.A(\spiking_network_top_uut.all_data_out[79] ));
 sg13g2_antennanp ANTENNA_400 (.A(\spiking_network_top_uut.all_data_out[79] ));
 sg13g2_antennanp ANTENNA_401 (.A(\spiking_network_top_uut.all_data_out[848] ));
 sg13g2_antennanp ANTENNA_402 (.A(\spiking_network_top_uut.all_data_out[848] ));
 sg13g2_antennanp ANTENNA_403 (.A(\spiking_network_top_uut.all_data_out[848] ));
 sg13g2_antennanp ANTENNA_404 (.A(\spiking_network_top_uut.all_data_out[848] ));
 sg13g2_antennanp ANTENNA_405 (.A(\spiking_network_top_uut.all_data_out[848] ));
 sg13g2_antennanp ANTENNA_406 (.A(\spiking_network_top_uut.all_data_out[848] ));
 sg13g2_antennanp ANTENNA_407 (.A(\spiking_network_top_uut.all_data_out[848] ));
 sg13g2_antennanp ANTENNA_408 (.A(\spiking_network_top_uut.all_data_out[848] ));
 sg13g2_antennanp ANTENNA_409 (.A(\spiking_network_top_uut.all_data_out[848] ));
 sg13g2_antennanp ANTENNA_410 (.A(\spiking_network_top_uut.all_data_out[867] ));
 sg13g2_antennanp ANTENNA_411 (.A(\spiking_network_top_uut.all_data_out[867] ));
 sg13g2_antennanp ANTENNA_412 (.A(\spiking_network_top_uut.all_data_out[867] ));
 sg13g2_antennanp ANTENNA_413 (.A(\spiking_network_top_uut.all_data_out[867] ));
 sg13g2_antennanp ANTENNA_414 (.A(\spiking_network_top_uut.all_data_out[867] ));
 sg13g2_antennanp ANTENNA_415 (.A(\spiking_network_top_uut.all_data_out[867] ));
 sg13g2_antennanp ANTENNA_416 (.A(\spiking_network_top_uut.all_data_out[867] ));
 sg13g2_antennanp ANTENNA_417 (.A(\spiking_network_top_uut.all_data_out[867] ));
 sg13g2_antennanp ANTENNA_418 (.A(\spiking_network_top_uut.all_data_out[867] ));
 sg13g2_antennanp ANTENNA_419 (.A(\spiking_network_top_uut.all_data_out[867] ));
 sg13g2_antennanp ANTENNA_420 (.A(\spiking_network_top_uut.all_data_out[896] ));
 sg13g2_antennanp ANTENNA_421 (.A(\spiking_network_top_uut.all_data_out[896] ));
 sg13g2_antennanp ANTENNA_422 (.A(\spiking_network_top_uut.all_data_out[896] ));
 sg13g2_antennanp ANTENNA_423 (.A(\spiking_network_top_uut.all_data_out[896] ));
 sg13g2_antennanp ANTENNA_424 (.A(\spiking_network_top_uut.all_data_out[896] ));
 sg13g2_antennanp ANTENNA_425 (.A(\spiking_network_top_uut.all_data_out[896] ));
 sg13g2_antennanp ANTENNA_426 (.A(\spiking_network_top_uut.all_data_out[896] ));
 sg13g2_antennanp ANTENNA_427 (.A(\spiking_network_top_uut.all_data_out[896] ));
 sg13g2_antennanp ANTENNA_428 (.A(\spiking_network_top_uut.all_data_out[896] ));
 sg13g2_antennanp ANTENNA_429 (.A(\spiking_network_top_uut.all_data_out[897] ));
 sg13g2_antennanp ANTENNA_430 (.A(\spiking_network_top_uut.all_data_out[897] ));
 sg13g2_antennanp ANTENNA_431 (.A(\spiking_network_top_uut.all_data_out[897] ));
 sg13g2_antennanp ANTENNA_432 (.A(\spiking_network_top_uut.all_data_out[897] ));
 sg13g2_antennanp ANTENNA_433 (.A(\spiking_network_top_uut.all_data_out[897] ));
 sg13g2_antennanp ANTENNA_434 (.A(\spiking_network_top_uut.all_data_out[897] ));
 sg13g2_antennanp ANTENNA_435 (.A(\spiking_network_top_uut.all_data_out[898] ));
 sg13g2_antennanp ANTENNA_436 (.A(\spiking_network_top_uut.all_data_out[898] ));
 sg13g2_antennanp ANTENNA_437 (.A(\spiking_network_top_uut.all_data_out[898] ));
 sg13g2_antennanp ANTENNA_438 (.A(\spiking_network_top_uut.all_data_out[898] ));
 sg13g2_antennanp ANTENNA_439 (.A(\spiking_network_top_uut.all_data_out[898] ));
 sg13g2_antennanp ANTENNA_440 (.A(\spiking_network_top_uut.all_data_out[898] ));
 sg13g2_antennanp ANTENNA_441 (.A(\spiking_network_top_uut.all_data_out[898] ));
 sg13g2_antennanp ANTENNA_442 (.A(\spiking_network_top_uut.all_data_out[898] ));
 sg13g2_antennanp ANTENNA_443 (.A(\spiking_network_top_uut.all_data_out[898] ));
 sg13g2_antennanp ANTENNA_444 (.A(\spiking_network_top_uut.all_data_out[899] ));
 sg13g2_antennanp ANTENNA_445 (.A(\spiking_network_top_uut.all_data_out[899] ));
 sg13g2_antennanp ANTENNA_446 (.A(\spiking_network_top_uut.all_data_out[899] ));
 sg13g2_antennanp ANTENNA_447 (.A(\spiking_network_top_uut.all_data_out[899] ));
 sg13g2_antennanp ANTENNA_448 (.A(\spiking_network_top_uut.all_data_out[899] ));
 sg13g2_antennanp ANTENNA_449 (.A(\spiking_network_top_uut.all_data_out[899] ));
 sg13g2_antennanp ANTENNA_450 (.A(\spiking_network_top_uut.all_data_out[901] ));
 sg13g2_antennanp ANTENNA_451 (.A(\spiking_network_top_uut.all_data_out[901] ));
 sg13g2_antennanp ANTENNA_452 (.A(\spiking_network_top_uut.all_data_out[901] ));
 sg13g2_antennanp ANTENNA_453 (.A(\spiking_network_top_uut.all_data_out[901] ));
 sg13g2_antennanp ANTENNA_454 (.A(\spiking_network_top_uut.all_data_out[901] ));
 sg13g2_antennanp ANTENNA_455 (.A(\spiking_network_top_uut.all_data_out[901] ));
 sg13g2_antennanp ANTENNA_456 (.A(\spiking_network_top_uut.all_data_out[902] ));
 sg13g2_antennanp ANTENNA_457 (.A(\spiking_network_top_uut.all_data_out[902] ));
 sg13g2_antennanp ANTENNA_458 (.A(\spiking_network_top_uut.all_data_out[902] ));
 sg13g2_antennanp ANTENNA_459 (.A(\spiking_network_top_uut.all_data_out[902] ));
 sg13g2_antennanp ANTENNA_460 (.A(\spiking_network_top_uut.all_data_out[902] ));
 sg13g2_antennanp ANTENNA_461 (.A(\spiking_network_top_uut.all_data_out[902] ));
 sg13g2_antennanp ANTENNA_462 (.A(\spiking_network_top_uut.all_data_out[902] ));
 sg13g2_antennanp ANTENNA_463 (.A(\spiking_network_top_uut.all_data_out[902] ));
 sg13g2_antennanp ANTENNA_464 (.A(\spiking_network_top_uut.all_data_out[902] ));
 sg13g2_antennanp ANTENNA_465 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.enable_LYR_2 ));
 sg13g2_antennanp ANTENNA_466 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.enable_LYR_2 ));
 sg13g2_antennanp ANTENNA_467 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.enable_LYR_2 ));
 sg13g2_antennanp ANTENNA_468 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.enable_LYR_2 ));
 sg13g2_antennanp ANTENNA_469 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.enable_LYR_2 ));
 sg13g2_antennanp ANTENNA_470 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.enable_LYR_2 ));
 sg13g2_antennanp ANTENNA_471 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.enable_LYR_2 ));
 sg13g2_antennanp ANTENNA_472 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.enable_LYR_2 ));
 sg13g2_antennanp ANTENNA_473 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.enable_LYR_2 ));
 sg13g2_antennanp ANTENNA_474 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.enable_LYR_2 ));
 sg13g2_antennanp ANTENNA_475 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.enable_LYR_2 ));
 sg13g2_antennanp ANTENNA_476 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.enable_LYR_2 ));
 sg13g2_antennanp ANTENNA_477 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.enable_LYR_2 ));
 sg13g2_antennanp ANTENNA_478 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.enable_LYR_2 ));
 sg13g2_antennanp ANTENNA_479 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ));
 sg13g2_antennanp ANTENNA_480 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ));
 sg13g2_antennanp ANTENNA_481 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ));
 sg13g2_antennanp ANTENNA_482 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ));
 sg13g2_antennanp ANTENNA_483 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ));
 sg13g2_antennanp ANTENNA_484 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ));
 sg13g2_antennanp ANTENNA_485 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[4] ));
 sg13g2_antennanp ANTENNA_486 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_487 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_488 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_489 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_490 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_491 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_492 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_493 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_494 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_495 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_496 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_497 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_498 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_499 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_500 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_501 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_502 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ));
 sg13g2_antennanp ANTENNA_503 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ));
 sg13g2_antennanp ANTENNA_504 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ));
 sg13g2_antennanp ANTENNA_505 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ));
 sg13g2_antennanp ANTENNA_506 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ));
 sg13g2_antennanp ANTENNA_507 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ));
 sg13g2_antennanp ANTENNA_508 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ));
 sg13g2_antennanp ANTENNA_509 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.lif_neuron_inst.lif_neuron_inst.membrane_potential[3] ));
 sg13g2_antennanp ANTENNA_510 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_511 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_512 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_513 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_514 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_515 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_516 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_517 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_518 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_519 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_520 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.spike_out ));
 sg13g2_antennanp ANTENNA_521 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.spike_out ));
 sg13g2_antennanp ANTENNA_522 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.spike_out ));
 sg13g2_antennanp ANTENNA_523 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_524 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_525 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_526 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_527 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_528 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_529 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_530 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_531 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_532 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_533 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_534 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[7].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_535 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_536 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_537 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_538 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_539 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_540 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_541 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_542 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_543 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.neuron_delay_gen[5].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_544 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.spike_out ));
 sg13g2_antennanp ANTENNA_545 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.spike_out ));
 sg13g2_antennanp ANTENNA_546 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.spike_out ));
 sg13g2_antennanp ANTENNA_547 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.spike_out ));
 sg13g2_antennanp ANTENNA_548 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.spike_out ));
 sg13g2_antennanp ANTENNA_549 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.spike_out ));
 sg13g2_antennanp ANTENNA_550 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.spike_out ));
 sg13g2_antennanp ANTENNA_551 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.lif_neuron_inst.lif_neuron_inst.spike_out ));
 sg13g2_antennanp ANTENNA_552 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_reg1 ));
 sg13g2_antennanp ANTENNA_553 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_reg1 ));
 sg13g2_antennanp ANTENNA_554 (.A(net3658));
 sg13g2_antennanp ANTENNA_555 (.A(net3658));
 sg13g2_antennanp ANTENNA_556 (.A(net3658));
 sg13g2_antennanp ANTENNA_557 (.A(net3658));
 sg13g2_antennanp ANTENNA_558 (.A(net3658));
 sg13g2_antennanp ANTENNA_559 (.A(net3658));
 sg13g2_antennanp ANTENNA_560 (.A(net3728));
 sg13g2_antennanp ANTENNA_561 (.A(net3728));
 sg13g2_antennanp ANTENNA_562 (.A(net3728));
 sg13g2_antennanp ANTENNA_563 (.A(net3728));
 sg13g2_antennanp ANTENNA_564 (.A(net3728));
 sg13g2_antennanp ANTENNA_565 (.A(net3728));
 sg13g2_antennanp ANTENNA_566 (.A(net3728));
 sg13g2_antennanp ANTENNA_567 (.A(net3728));
 sg13g2_antennanp ANTENNA_568 (.A(net3965));
 sg13g2_antennanp ANTENNA_569 (.A(net3965));
 sg13g2_antennanp ANTENNA_570 (.A(net3965));
 sg13g2_antennanp ANTENNA_571 (.A(net3965));
 sg13g2_antennanp ANTENNA_572 (.A(net3965));
 sg13g2_antennanp ANTENNA_573 (.A(net3965));
 sg13g2_antennanp ANTENNA_574 (.A(net3965));
 sg13g2_antennanp ANTENNA_575 (.A(net3965));
 sg13g2_antennanp ANTENNA_576 (.A(net3965));
 sg13g2_antennanp ANTENNA_577 (.A(net3965));
 sg13g2_antennanp ANTENNA_578 (.A(net3965));
 sg13g2_antennanp ANTENNA_579 (.A(net3965));
 sg13g2_antennanp ANTENNA_580 (.A(net3965));
 sg13g2_antennanp ANTENNA_581 (.A(net3965));
 sg13g2_antennanp ANTENNA_582 (.A(net3965));
 sg13g2_antennanp ANTENNA_583 (.A(net3965));
 sg13g2_antennanp ANTENNA_584 (.A(net3965));
 sg13g2_antennanp ANTENNA_585 (.A(net3965));
 sg13g2_antennanp ANTENNA_586 (.A(net3965));
 sg13g2_antennanp ANTENNA_587 (.A(net4136));
 sg13g2_antennanp ANTENNA_588 (.A(net4136));
 sg13g2_antennanp ANTENNA_589 (.A(net4136));
 sg13g2_antennanp ANTENNA_590 (.A(net4136));
 sg13g2_antennanp ANTENNA_591 (.A(net4136));
 sg13g2_antennanp ANTENNA_592 (.A(net4162));
 sg13g2_antennanp ANTENNA_593 (.A(net4162));
 sg13g2_antennanp ANTENNA_594 (.A(net4162));
 sg13g2_antennanp ANTENNA_595 (.A(net4162));
 sg13g2_antennanp ANTENNA_596 (.A(net4162));
 sg13g2_antennanp ANTENNA_597 (.A(net4162));
 sg13g2_antennanp ANTENNA_598 (.A(net4162));
 sg13g2_antennanp ANTENNA_599 (.A(net4162));
 sg13g2_antennanp ANTENNA_600 (.A(net4162));
 sg13g2_antennanp ANTENNA_601 (.A(net4162));
 sg13g2_antennanp ANTENNA_602 (.A(net4162));
 sg13g2_antennanp ANTENNA_603 (.A(net4709));
 sg13g2_antennanp ANTENNA_604 (.A(net4709));
 sg13g2_antennanp ANTENNA_605 (.A(net4709));
 sg13g2_antennanp ANTENNA_606 (.A(net4709));
 sg13g2_antennanp ANTENNA_607 (.A(net4709));
 sg13g2_antennanp ANTENNA_608 (.A(net2));
 sg13g2_antennanp ANTENNA_609 (.A(net3));
 sg13g2_antennanp ANTENNA_610 (.A(net4));
 sg13g2_antennanp ANTENNA_611 (.A(net5));
 sg13g2_antennanp ANTENNA_612 (.A(net6));
 sg13g2_antennanp ANTENNA_613 (.A(net8));
 sg13g2_antennanp ANTENNA_614 (.A(net9));
 sg13g2_antennanp ANTENNA_615 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_616 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_617 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_618 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_619 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_620 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_621 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_622 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_623 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_624 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_625 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_626 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_627 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_628 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_629 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_630 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_631 (.A(clknet_4_3__leaf_clk));
 sg13g2_antennanp ANTENNA_632 (.A(clknet_4_3__leaf_clk));
 sg13g2_antennanp ANTENNA_633 (.A(clknet_4_3__leaf_clk));
 sg13g2_antennanp ANTENNA_634 (.A(clknet_4_3__leaf_clk));
 sg13g2_antennanp ANTENNA_635 (.A(clknet_4_3__leaf_clk));
 sg13g2_antennanp ANTENNA_636 (.A(clknet_4_3__leaf_clk));
 sg13g2_antennanp ANTENNA_637 (.A(clknet_4_3__leaf_clk));
 sg13g2_antennanp ANTENNA_638 (.A(clknet_4_3__leaf_clk));
 sg13g2_antennanp ANTENNA_639 (.A(clknet_4_3__leaf_clk));
 sg13g2_antennanp ANTENNA_640 (.A(clknet_4_3__leaf_clk));
 sg13g2_antennanp ANTENNA_641 (.A(clknet_4_3__leaf_clk));
 sg13g2_antennanp ANTENNA_642 (.A(_00026_));
 sg13g2_antennanp ANTENNA_643 (.A(_00026_));
 sg13g2_antennanp ANTENNA_644 (.A(_00026_));
 sg13g2_antennanp ANTENNA_645 (.A(_00026_));
 sg13g2_antennanp ANTENNA_646 (.A(_00146_));
 sg13g2_antennanp ANTENNA_647 (.A(_00148_));
 sg13g2_antennanp ANTENNA_648 (.A(_00158_));
 sg13g2_antennanp ANTENNA_649 (.A(_00188_));
 sg13g2_antennanp ANTENNA_650 (.A(_00197_));
 sg13g2_antennanp ANTENNA_651 (.A(_00199_));
 sg13g2_antennanp ANTENNA_652 (.A(_00201_));
 sg13g2_antennanp ANTENNA_653 (.A(_00208_));
 sg13g2_antennanp ANTENNA_654 (.A(_00209_));
 sg13g2_antennanp ANTENNA_655 (.A(_00213_));
 sg13g2_antennanp ANTENNA_656 (.A(_00217_));
 sg13g2_antennanp ANTENNA_657 (.A(_00226_));
 sg13g2_antennanp ANTENNA_658 (.A(_00251_));
 sg13g2_antennanp ANTENNA_659 (.A(_00258_));
 sg13g2_antennanp ANTENNA_660 (.A(_00259_));
 sg13g2_antennanp ANTENNA_661 (.A(_00271_));
 sg13g2_antennanp ANTENNA_662 (.A(_00283_));
 sg13g2_antennanp ANTENNA_663 (.A(_00284_));
 sg13g2_antennanp ANTENNA_664 (.A(_00288_));
 sg13g2_antennanp ANTENNA_665 (.A(_00299_));
 sg13g2_antennanp ANTENNA_666 (.A(_00328_));
 sg13g2_antennanp ANTENNA_667 (.A(_00329_));
 sg13g2_antennanp ANTENNA_668 (.A(_00347_));
 sg13g2_antennanp ANTENNA_669 (.A(_00390_));
 sg13g2_antennanp ANTENNA_670 (.A(_00391_));
 sg13g2_antennanp ANTENNA_671 (.A(_00411_));
 sg13g2_antennanp ANTENNA_672 (.A(_00415_));
 sg13g2_antennanp ANTENNA_673 (.A(_00419_));
 sg13g2_antennanp ANTENNA_674 (.A(_02216_));
 sg13g2_antennanp ANTENNA_675 (.A(_02406_));
 sg13g2_antennanp ANTENNA_676 (.A(_02406_));
 sg13g2_antennanp ANTENNA_677 (.A(_02406_));
 sg13g2_antennanp ANTENNA_678 (.A(_02406_));
 sg13g2_antennanp ANTENNA_679 (.A(_02483_));
 sg13g2_antennanp ANTENNA_680 (.A(_02483_));
 sg13g2_antennanp ANTENNA_681 (.A(_02483_));
 sg13g2_antennanp ANTENNA_682 (.A(_02483_));
 sg13g2_antennanp ANTENNA_683 (.A(_02483_));
 sg13g2_antennanp ANTENNA_684 (.A(_02483_));
 sg13g2_antennanp ANTENNA_685 (.A(_02483_));
 sg13g2_antennanp ANTENNA_686 (.A(_02483_));
 sg13g2_antennanp ANTENNA_687 (.A(_02483_));
 sg13g2_antennanp ANTENNA_688 (.A(_02484_));
 sg13g2_antennanp ANTENNA_689 (.A(_02484_));
 sg13g2_antennanp ANTENNA_690 (.A(_02484_));
 sg13g2_antennanp ANTENNA_691 (.A(_02484_));
 sg13g2_antennanp ANTENNA_692 (.A(_02494_));
 sg13g2_antennanp ANTENNA_693 (.A(_02494_));
 sg13g2_antennanp ANTENNA_694 (.A(_02494_));
 sg13g2_antennanp ANTENNA_695 (.A(_02494_));
 sg13g2_antennanp ANTENNA_696 (.A(_02495_));
 sg13g2_antennanp ANTENNA_697 (.A(_02495_));
 sg13g2_antennanp ANTENNA_698 (.A(_02495_));
 sg13g2_antennanp ANTENNA_699 (.A(_02495_));
 sg13g2_antennanp ANTENNA_700 (.A(_02495_));
 sg13g2_antennanp ANTENNA_701 (.A(_02495_));
 sg13g2_antennanp ANTENNA_702 (.A(_02495_));
 sg13g2_antennanp ANTENNA_703 (.A(_02495_));
 sg13g2_antennanp ANTENNA_704 (.A(_02495_));
 sg13g2_antennanp ANTENNA_705 (.A(_02509_));
 sg13g2_antennanp ANTENNA_706 (.A(_02509_));
 sg13g2_antennanp ANTENNA_707 (.A(_02509_));
 sg13g2_antennanp ANTENNA_708 (.A(_02509_));
 sg13g2_antennanp ANTENNA_709 (.A(_02777_));
 sg13g2_antennanp ANTENNA_710 (.A(_02777_));
 sg13g2_antennanp ANTENNA_711 (.A(_02777_));
 sg13g2_antennanp ANTENNA_712 (.A(_02777_));
 sg13g2_antennanp ANTENNA_713 (.A(_02785_));
 sg13g2_antennanp ANTENNA_714 (.A(_02991_));
 sg13g2_antennanp ANTENNA_715 (.A(_02991_));
 sg13g2_antennanp ANTENNA_716 (.A(_02991_));
 sg13g2_antennanp ANTENNA_717 (.A(_02991_));
 sg13g2_antennanp ANTENNA_718 (.A(_02991_));
 sg13g2_antennanp ANTENNA_719 (.A(_02991_));
 sg13g2_antennanp ANTENNA_720 (.A(_02991_));
 sg13g2_antennanp ANTENNA_721 (.A(_02991_));
 sg13g2_antennanp ANTENNA_722 (.A(_02991_));
 sg13g2_antennanp ANTENNA_723 (.A(_03215_));
 sg13g2_antennanp ANTENNA_724 (.A(_03215_));
 sg13g2_antennanp ANTENNA_725 (.A(_03215_));
 sg13g2_antennanp ANTENNA_726 (.A(_03215_));
 sg13g2_antennanp ANTENNA_727 (.A(_03215_));
 sg13g2_antennanp ANTENNA_728 (.A(_03215_));
 sg13g2_antennanp ANTENNA_729 (.A(_03215_));
 sg13g2_antennanp ANTENNA_730 (.A(_03215_));
 sg13g2_antennanp ANTENNA_731 (.A(_03215_));
 sg13g2_antennanp ANTENNA_732 (.A(_03215_));
 sg13g2_antennanp ANTENNA_733 (.A(_03215_));
 sg13g2_antennanp ANTENNA_734 (.A(_03215_));
 sg13g2_antennanp ANTENNA_735 (.A(_03215_));
 sg13g2_antennanp ANTENNA_736 (.A(_03215_));
 sg13g2_antennanp ANTENNA_737 (.A(_03215_));
 sg13g2_antennanp ANTENNA_738 (.A(_03215_));
 sg13g2_antennanp ANTENNA_739 (.A(_03215_));
 sg13g2_antennanp ANTENNA_740 (.A(_03509_));
 sg13g2_antennanp ANTENNA_741 (.A(_03518_));
 sg13g2_antennanp ANTENNA_742 (.A(_03522_));
 sg13g2_antennanp ANTENNA_743 (.A(_03534_));
 sg13g2_antennanp ANTENNA_744 (.A(_03543_));
 sg13g2_antennanp ANTENNA_745 (.A(_03549_));
 sg13g2_antennanp ANTENNA_746 (.A(_03550_));
 sg13g2_antennanp ANTENNA_747 (.A(_03551_));
 sg13g2_antennanp ANTENNA_748 (.A(_03567_));
 sg13g2_antennanp ANTENNA_749 (.A(_03571_));
 sg13g2_antennanp ANTENNA_750 (.A(_03573_));
 sg13g2_antennanp ANTENNA_751 (.A(_03574_));
 sg13g2_antennanp ANTENNA_752 (.A(_03576_));
 sg13g2_antennanp ANTENNA_753 (.A(_03578_));
 sg13g2_antennanp ANTENNA_754 (.A(_03589_));
 sg13g2_antennanp ANTENNA_755 (.A(_03609_));
 sg13g2_antennanp ANTENNA_756 (.A(_03613_));
 sg13g2_antennanp ANTENNA_757 (.A(_03614_));
 sg13g2_antennanp ANTENNA_758 (.A(_03622_));
 sg13g2_antennanp ANTENNA_759 (.A(_03625_));
 sg13g2_antennanp ANTENNA_760 (.A(_03648_));
 sg13g2_antennanp ANTENNA_761 (.A(_03650_));
 sg13g2_antennanp ANTENNA_762 (.A(_03651_));
 sg13g2_antennanp ANTENNA_763 (.A(_03652_));
 sg13g2_antennanp ANTENNA_764 (.A(_03654_));
 sg13g2_antennanp ANTENNA_765 (.A(_03794_));
 sg13g2_antennanp ANTENNA_766 (.A(_03794_));
 sg13g2_antennanp ANTENNA_767 (.A(_03794_));
 sg13g2_antennanp ANTENNA_768 (.A(_03794_));
 sg13g2_antennanp ANTENNA_769 (.A(_03794_));
 sg13g2_antennanp ANTENNA_770 (.A(_03794_));
 sg13g2_antennanp ANTENNA_771 (.A(_03794_));
 sg13g2_antennanp ANTENNA_772 (.A(_03794_));
 sg13g2_antennanp ANTENNA_773 (.A(_03794_));
 sg13g2_antennanp ANTENNA_774 (.A(_03794_));
 sg13g2_antennanp ANTENNA_775 (.A(_03794_));
 sg13g2_antennanp ANTENNA_776 (.A(_03794_));
 sg13g2_antennanp ANTENNA_777 (.A(_03794_));
 sg13g2_antennanp ANTENNA_778 (.A(_03794_));
 sg13g2_antennanp ANTENNA_779 (.A(_03794_));
 sg13g2_antennanp ANTENNA_780 (.A(_03794_));
 sg13g2_antennanp ANTENNA_781 (.A(_03794_));
 sg13g2_antennanp ANTENNA_782 (.A(_03794_));
 sg13g2_antennanp ANTENNA_783 (.A(_03794_));
 sg13g2_antennanp ANTENNA_784 (.A(_03794_));
 sg13g2_antennanp ANTENNA_785 (.A(_03893_));
 sg13g2_antennanp ANTENNA_786 (.A(_03906_));
 sg13g2_antennanp ANTENNA_787 (.A(_03913_));
 sg13g2_antennanp ANTENNA_788 (.A(_03988_));
 sg13g2_antennanp ANTENNA_789 (.A(_03990_));
 sg13g2_antennanp ANTENNA_790 (.A(_03993_));
 sg13g2_antennanp ANTENNA_791 (.A(_03999_));
 sg13g2_antennanp ANTENNA_792 (.A(_04005_));
 sg13g2_antennanp ANTENNA_793 (.A(_04025_));
 sg13g2_antennanp ANTENNA_794 (.A(_04028_));
 sg13g2_antennanp ANTENNA_795 (.A(_04043_));
 sg13g2_antennanp ANTENNA_796 (.A(_04046_));
 sg13g2_antennanp ANTENNA_797 (.A(_04081_));
 sg13g2_antennanp ANTENNA_798 (.A(_04092_));
 sg13g2_antennanp ANTENNA_799 (.A(_04114_));
 sg13g2_antennanp ANTENNA_800 (.A(_04130_));
 sg13g2_antennanp ANTENNA_801 (.A(_04131_));
 sg13g2_antennanp ANTENNA_802 (.A(_04132_));
 sg13g2_antennanp ANTENNA_803 (.A(_04137_));
 sg13g2_antennanp ANTENNA_804 (.A(_04148_));
 sg13g2_antennanp ANTENNA_805 (.A(_04167_));
 sg13g2_antennanp ANTENNA_806 (.A(_04180_));
 sg13g2_antennanp ANTENNA_807 (.A(_04191_));
 sg13g2_antennanp ANTENNA_808 (.A(_04194_));
 sg13g2_antennanp ANTENNA_809 (.A(_04202_));
 sg13g2_antennanp ANTENNA_810 (.A(_04213_));
 sg13g2_antennanp ANTENNA_811 (.A(_04216_));
 sg13g2_antennanp ANTENNA_812 (.A(_04221_));
 sg13g2_antennanp ANTENNA_813 (.A(_04231_));
 sg13g2_antennanp ANTENNA_814 (.A(_04238_));
 sg13g2_antennanp ANTENNA_815 (.A(_04243_));
 sg13g2_antennanp ANTENNA_816 (.A(_04270_));
 sg13g2_antennanp ANTENNA_817 (.A(_04271_));
 sg13g2_antennanp ANTENNA_818 (.A(_04280_));
 sg13g2_antennanp ANTENNA_819 (.A(_04289_));
 sg13g2_antennanp ANTENNA_820 (.A(_04312_));
 sg13g2_antennanp ANTENNA_821 (.A(_04319_));
 sg13g2_antennanp ANTENNA_822 (.A(_04352_));
 sg13g2_antennanp ANTENNA_823 (.A(_04362_));
 sg13g2_antennanp ANTENNA_824 (.A(_04374_));
 sg13g2_antennanp ANTENNA_825 (.A(_04401_));
 sg13g2_antennanp ANTENNA_826 (.A(_04410_));
 sg13g2_antennanp ANTENNA_827 (.A(_04415_));
 sg13g2_antennanp ANTENNA_828 (.A(_04417_));
 sg13g2_antennanp ANTENNA_829 (.A(_04436_));
 sg13g2_antennanp ANTENNA_830 (.A(_04450_));
 sg13g2_antennanp ANTENNA_831 (.A(_04480_));
 sg13g2_antennanp ANTENNA_832 (.A(_04498_));
 sg13g2_antennanp ANTENNA_833 (.A(_04500_));
 sg13g2_antennanp ANTENNA_834 (.A(_04504_));
 sg13g2_antennanp ANTENNA_835 (.A(_04508_));
 sg13g2_antennanp ANTENNA_836 (.A(_04511_));
 sg13g2_antennanp ANTENNA_837 (.A(_04523_));
 sg13g2_antennanp ANTENNA_838 (.A(_04556_));
 sg13g2_antennanp ANTENNA_839 (.A(_04559_));
 sg13g2_antennanp ANTENNA_840 (.A(_04562_));
 sg13g2_antennanp ANTENNA_841 (.A(_04578_));
 sg13g2_antennanp ANTENNA_842 (.A(_04579_));
 sg13g2_antennanp ANTENNA_843 (.A(_04580_));
 sg13g2_antennanp ANTENNA_844 (.A(_04584_));
 sg13g2_antennanp ANTENNA_845 (.A(_05709_));
 sg13g2_antennanp ANTENNA_846 (.A(_05709_));
 sg13g2_antennanp ANTENNA_847 (.A(_05709_));
 sg13g2_antennanp ANTENNA_848 (.A(_05709_));
 sg13g2_antennanp ANTENNA_849 (.A(_05805_));
 sg13g2_antennanp ANTENNA_850 (.A(_06082_));
 sg13g2_antennanp ANTENNA_851 (.A(_06284_));
 sg13g2_antennanp ANTENNA_852 (.A(_06284_));
 sg13g2_antennanp ANTENNA_853 (.A(_06284_));
 sg13g2_antennanp ANTENNA_854 (.A(_06284_));
 sg13g2_antennanp ANTENNA_855 (.A(_06286_));
 sg13g2_antennanp ANTENNA_856 (.A(_06286_));
 sg13g2_antennanp ANTENNA_857 (.A(_06286_));
 sg13g2_antennanp ANTENNA_858 (.A(_06286_));
 sg13g2_antennanp ANTENNA_859 (.A(_06625_));
 sg13g2_antennanp ANTENNA_860 (.A(_06625_));
 sg13g2_antennanp ANTENNA_861 (.A(_06625_));
 sg13g2_antennanp ANTENNA_862 (.A(_06625_));
 sg13g2_antennanp ANTENNA_863 (.A(_07721_));
 sg13g2_antennanp ANTENNA_864 (.A(_07721_));
 sg13g2_antennanp ANTENNA_865 (.A(_07721_));
 sg13g2_antennanp ANTENNA_866 (.A(_07721_));
 sg13g2_antennanp ANTENNA_867 (.A(_08106_));
 sg13g2_antennanp ANTENNA_868 (.A(_08106_));
 sg13g2_antennanp ANTENNA_869 (.A(_08106_));
 sg13g2_antennanp ANTENNA_870 (.A(_08106_));
 sg13g2_antennanp ANTENNA_871 (.A(_08570_));
 sg13g2_antennanp ANTENNA_872 (.A(_08570_));
 sg13g2_antennanp ANTENNA_873 (.A(_08570_));
 sg13g2_antennanp ANTENNA_874 (.A(_08570_));
 sg13g2_antennanp ANTENNA_875 (.A(_08849_));
 sg13g2_antennanp ANTENNA_876 (.A(_08849_));
 sg13g2_antennanp ANTENNA_877 (.A(_08849_));
 sg13g2_antennanp ANTENNA_878 (.A(_08849_));
 sg13g2_antennanp ANTENNA_879 (.A(_08849_));
 sg13g2_antennanp ANTENNA_880 (.A(_08849_));
 sg13g2_antennanp ANTENNA_881 (.A(_08849_));
 sg13g2_antennanp ANTENNA_882 (.A(_08849_));
 sg13g2_antennanp ANTENNA_883 (.A(_08849_));
 sg13g2_antennanp ANTENNA_884 (.A(_08860_));
 sg13g2_antennanp ANTENNA_885 (.A(_08860_));
 sg13g2_antennanp ANTENNA_886 (.A(_08860_));
 sg13g2_antennanp ANTENNA_887 (.A(_08860_));
 sg13g2_antennanp ANTENNA_888 (.A(\spiking_network_top_uut.all_data_out[17] ));
 sg13g2_antennanp ANTENNA_889 (.A(\spiking_network_top_uut.all_data_out[17] ));
 sg13g2_antennanp ANTENNA_890 (.A(\spiking_network_top_uut.all_data_out[17] ));
 sg13g2_antennanp ANTENNA_891 (.A(\spiking_network_top_uut.all_data_out[17] ));
 sg13g2_antennanp ANTENNA_892 (.A(\spiking_network_top_uut.all_data_out[273] ));
 sg13g2_antennanp ANTENNA_893 (.A(\spiking_network_top_uut.all_data_out[273] ));
 sg13g2_antennanp ANTENNA_894 (.A(\spiking_network_top_uut.all_data_out[273] ));
 sg13g2_antennanp ANTENNA_895 (.A(\spiking_network_top_uut.all_data_out[294] ));
 sg13g2_antennanp ANTENNA_896 (.A(\spiking_network_top_uut.all_data_out[294] ));
 sg13g2_antennanp ANTENNA_897 (.A(\spiking_network_top_uut.all_data_out[294] ));
 sg13g2_antennanp ANTENNA_898 (.A(\spiking_network_top_uut.all_data_out[294] ));
 sg13g2_antennanp ANTENNA_899 (.A(\spiking_network_top_uut.all_data_out[294] ));
 sg13g2_antennanp ANTENNA_900 (.A(\spiking_network_top_uut.all_data_out[294] ));
 sg13g2_antennanp ANTENNA_901 (.A(\spiking_network_top_uut.all_data_out[294] ));
 sg13g2_antennanp ANTENNA_902 (.A(\spiking_network_top_uut.all_data_out[294] ));
 sg13g2_antennanp ANTENNA_903 (.A(\spiking_network_top_uut.all_data_out[294] ));
 sg13g2_antennanp ANTENNA_904 (.A(\spiking_network_top_uut.all_data_out[295] ));
 sg13g2_antennanp ANTENNA_905 (.A(\spiking_network_top_uut.all_data_out[295] ));
 sg13g2_antennanp ANTENNA_906 (.A(\spiking_network_top_uut.all_data_out[295] ));
 sg13g2_antennanp ANTENNA_907 (.A(\spiking_network_top_uut.all_data_out[295] ));
 sg13g2_antennanp ANTENNA_908 (.A(\spiking_network_top_uut.all_data_out[295] ));
 sg13g2_antennanp ANTENNA_909 (.A(\spiking_network_top_uut.all_data_out[295] ));
 sg13g2_antennanp ANTENNA_910 (.A(\spiking_network_top_uut.all_data_out[295] ));
 sg13g2_antennanp ANTENNA_911 (.A(\spiking_network_top_uut.all_data_out[295] ));
 sg13g2_antennanp ANTENNA_912 (.A(\spiking_network_top_uut.all_data_out[299] ));
 sg13g2_antennanp ANTENNA_913 (.A(\spiking_network_top_uut.all_data_out[299] ));
 sg13g2_antennanp ANTENNA_914 (.A(\spiking_network_top_uut.all_data_out[299] ));
 sg13g2_antennanp ANTENNA_915 (.A(\spiking_network_top_uut.all_data_out[299] ));
 sg13g2_antennanp ANTENNA_916 (.A(\spiking_network_top_uut.all_data_out[299] ));
 sg13g2_antennanp ANTENNA_917 (.A(\spiking_network_top_uut.all_data_out[299] ));
 sg13g2_antennanp ANTENNA_918 (.A(\spiking_network_top_uut.all_data_out[299] ));
 sg13g2_antennanp ANTENNA_919 (.A(\spiking_network_top_uut.all_data_out[299] ));
 sg13g2_antennanp ANTENNA_920 (.A(\spiking_network_top_uut.all_data_out[299] ));
 sg13g2_antennanp ANTENNA_921 (.A(\spiking_network_top_uut.all_data_out[299] ));
 sg13g2_antennanp ANTENNA_922 (.A(\spiking_network_top_uut.all_data_out[299] ));
 sg13g2_antennanp ANTENNA_923 (.A(\spiking_network_top_uut.all_data_out[299] ));
 sg13g2_antennanp ANTENNA_924 (.A(\spiking_network_top_uut.all_data_out[299] ));
 sg13g2_antennanp ANTENNA_925 (.A(\spiking_network_top_uut.all_data_out[307] ));
 sg13g2_antennanp ANTENNA_926 (.A(\spiking_network_top_uut.all_data_out[307] ));
 sg13g2_antennanp ANTENNA_927 (.A(\spiking_network_top_uut.all_data_out[307] ));
 sg13g2_antennanp ANTENNA_928 (.A(\spiking_network_top_uut.all_data_out[308] ));
 sg13g2_antennanp ANTENNA_929 (.A(\spiking_network_top_uut.all_data_out[308] ));
 sg13g2_antennanp ANTENNA_930 (.A(\spiking_network_top_uut.all_data_out[308] ));
 sg13g2_antennanp ANTENNA_931 (.A(\spiking_network_top_uut.all_data_out[311] ));
 sg13g2_antennanp ANTENNA_932 (.A(\spiking_network_top_uut.all_data_out[311] ));
 sg13g2_antennanp ANTENNA_933 (.A(\spiking_network_top_uut.all_data_out[311] ));
 sg13g2_antennanp ANTENNA_934 (.A(\spiking_network_top_uut.all_data_out[311] ));
 sg13g2_antennanp ANTENNA_935 (.A(\spiking_network_top_uut.all_data_out[311] ));
 sg13g2_antennanp ANTENNA_936 (.A(\spiking_network_top_uut.all_data_out[311] ));
 sg13g2_antennanp ANTENNA_937 (.A(\spiking_network_top_uut.all_data_out[330] ));
 sg13g2_antennanp ANTENNA_938 (.A(\spiking_network_top_uut.all_data_out[330] ));
 sg13g2_antennanp ANTENNA_939 (.A(\spiking_network_top_uut.all_data_out[330] ));
 sg13g2_antennanp ANTENNA_940 (.A(\spiking_network_top_uut.all_data_out[330] ));
 sg13g2_antennanp ANTENNA_941 (.A(\spiking_network_top_uut.all_data_out[584] ));
 sg13g2_antennanp ANTENNA_942 (.A(\spiking_network_top_uut.all_data_out[584] ));
 sg13g2_antennanp ANTENNA_943 (.A(\spiking_network_top_uut.all_data_out[584] ));
 sg13g2_antennanp ANTENNA_944 (.A(\spiking_network_top_uut.all_data_out[584] ));
 sg13g2_antennanp ANTENNA_945 (.A(\spiking_network_top_uut.all_data_out[584] ));
 sg13g2_antennanp ANTENNA_946 (.A(\spiking_network_top_uut.all_data_out[584] ));
 sg13g2_antennanp ANTENNA_947 (.A(\spiking_network_top_uut.all_data_out[584] ));
 sg13g2_antennanp ANTENNA_948 (.A(\spiking_network_top_uut.all_data_out[584] ));
 sg13g2_antennanp ANTENNA_949 (.A(\spiking_network_top_uut.all_data_out[584] ));
 sg13g2_antennanp ANTENNA_950 (.A(\spiking_network_top_uut.all_data_out[584] ));
 sg13g2_antennanp ANTENNA_951 (.A(\spiking_network_top_uut.all_data_out[584] ));
 sg13g2_antennanp ANTENNA_952 (.A(\spiking_network_top_uut.all_data_out[584] ));
 sg13g2_antennanp ANTENNA_953 (.A(\spiking_network_top_uut.all_data_out[584] ));
 sg13g2_antennanp ANTENNA_954 (.A(\spiking_network_top_uut.all_data_out[584] ));
 sg13g2_antennanp ANTENNA_955 (.A(\spiking_network_top_uut.all_data_out[584] ));
 sg13g2_antennanp ANTENNA_956 (.A(\spiking_network_top_uut.all_data_out[584] ));
 sg13g2_antennanp ANTENNA_957 (.A(\spiking_network_top_uut.all_data_out[76] ));
 sg13g2_antennanp ANTENNA_958 (.A(\spiking_network_top_uut.all_data_out[76] ));
 sg13g2_antennanp ANTENNA_959 (.A(\spiking_network_top_uut.all_data_out[76] ));
 sg13g2_antennanp ANTENNA_960 (.A(\spiking_network_top_uut.all_data_out[76] ));
 sg13g2_antennanp ANTENNA_961 (.A(\spiking_network_top_uut.all_data_out[79] ));
 sg13g2_antennanp ANTENNA_962 (.A(\spiking_network_top_uut.all_data_out[79] ));
 sg13g2_antennanp ANTENNA_963 (.A(\spiking_network_top_uut.all_data_out[79] ));
 sg13g2_antennanp ANTENNA_964 (.A(\spiking_network_top_uut.all_data_out[79] ));
 sg13g2_antennanp ANTENNA_965 (.A(\spiking_network_top_uut.all_data_out[79] ));
 sg13g2_antennanp ANTENNA_966 (.A(\spiking_network_top_uut.all_data_out[79] ));
 sg13g2_antennanp ANTENNA_967 (.A(\spiking_network_top_uut.all_data_out[79] ));
 sg13g2_antennanp ANTENNA_968 (.A(\spiking_network_top_uut.all_data_out[79] ));
 sg13g2_antennanp ANTENNA_969 (.A(\spiking_network_top_uut.all_data_out[79] ));
 sg13g2_antennanp ANTENNA_970 (.A(\spiking_network_top_uut.all_data_out[79] ));
 sg13g2_antennanp ANTENNA_971 (.A(\spiking_network_top_uut.all_data_out[79] ));
 sg13g2_antennanp ANTENNA_972 (.A(\spiking_network_top_uut.all_data_out[79] ));
 sg13g2_antennanp ANTENNA_973 (.A(\spiking_network_top_uut.all_data_out[79] ));
 sg13g2_antennanp ANTENNA_974 (.A(\spiking_network_top_uut.all_data_out[855] ));
 sg13g2_antennanp ANTENNA_975 (.A(\spiking_network_top_uut.all_data_out[855] ));
 sg13g2_antennanp ANTENNA_976 (.A(\spiking_network_top_uut.all_data_out[855] ));
 sg13g2_antennanp ANTENNA_977 (.A(\spiking_network_top_uut.all_data_out[896] ));
 sg13g2_antennanp ANTENNA_978 (.A(\spiking_network_top_uut.all_data_out[896] ));
 sg13g2_antennanp ANTENNA_979 (.A(\spiking_network_top_uut.all_data_out[896] ));
 sg13g2_antennanp ANTENNA_980 (.A(\spiking_network_top_uut.all_data_out[896] ));
 sg13g2_antennanp ANTENNA_981 (.A(\spiking_network_top_uut.all_data_out[896] ));
 sg13g2_antennanp ANTENNA_982 (.A(\spiking_network_top_uut.all_data_out[896] ));
 sg13g2_antennanp ANTENNA_983 (.A(\spiking_network_top_uut.all_data_out[896] ));
 sg13g2_antennanp ANTENNA_984 (.A(\spiking_network_top_uut.all_data_out[896] ));
 sg13g2_antennanp ANTENNA_985 (.A(\spiking_network_top_uut.all_data_out[896] ));
 sg13g2_antennanp ANTENNA_986 (.A(\spiking_network_top_uut.all_data_out[897] ));
 sg13g2_antennanp ANTENNA_987 (.A(\spiking_network_top_uut.all_data_out[897] ));
 sg13g2_antennanp ANTENNA_988 (.A(\spiking_network_top_uut.all_data_out[897] ));
 sg13g2_antennanp ANTENNA_989 (.A(\spiking_network_top_uut.all_data_out[897] ));
 sg13g2_antennanp ANTENNA_990 (.A(\spiking_network_top_uut.all_data_out[897] ));
 sg13g2_antennanp ANTENNA_991 (.A(\spiking_network_top_uut.all_data_out[897] ));
 sg13g2_antennanp ANTENNA_992 (.A(\spiking_network_top_uut.all_data_out[898] ));
 sg13g2_antennanp ANTENNA_993 (.A(\spiking_network_top_uut.all_data_out[898] ));
 sg13g2_antennanp ANTENNA_994 (.A(\spiking_network_top_uut.all_data_out[898] ));
 sg13g2_antennanp ANTENNA_995 (.A(\spiking_network_top_uut.all_data_out[898] ));
 sg13g2_antennanp ANTENNA_996 (.A(\spiking_network_top_uut.all_data_out[898] ));
 sg13g2_antennanp ANTENNA_997 (.A(\spiking_network_top_uut.all_data_out[898] ));
 sg13g2_antennanp ANTENNA_998 (.A(\spiking_network_top_uut.all_data_out[898] ));
 sg13g2_antennanp ANTENNA_999 (.A(\spiking_network_top_uut.all_data_out[898] ));
 sg13g2_antennanp ANTENNA_1000 (.A(\spiking_network_top_uut.all_data_out[898] ));
 sg13g2_antennanp ANTENNA_1001 (.A(\spiking_network_top_uut.all_data_out[899] ));
 sg13g2_antennanp ANTENNA_1002 (.A(\spiking_network_top_uut.all_data_out[899] ));
 sg13g2_antennanp ANTENNA_1003 (.A(\spiking_network_top_uut.all_data_out[899] ));
 sg13g2_antennanp ANTENNA_1004 (.A(\spiking_network_top_uut.all_data_out[899] ));
 sg13g2_antennanp ANTENNA_1005 (.A(\spiking_network_top_uut.all_data_out[899] ));
 sg13g2_antennanp ANTENNA_1006 (.A(\spiking_network_top_uut.all_data_out[899] ));
 sg13g2_antennanp ANTENNA_1007 (.A(\spiking_network_top_uut.all_data_out[902] ));
 sg13g2_antennanp ANTENNA_1008 (.A(\spiking_network_top_uut.all_data_out[902] ));
 sg13g2_antennanp ANTENNA_1009 (.A(\spiking_network_top_uut.all_data_out[902] ));
 sg13g2_antennanp ANTENNA_1010 (.A(\spiking_network_top_uut.all_data_out[902] ));
 sg13g2_antennanp ANTENNA_1011 (.A(\spiking_network_top_uut.all_data_out[902] ));
 sg13g2_antennanp ANTENNA_1012 (.A(\spiking_network_top_uut.all_data_out[902] ));
 sg13g2_antennanp ANTENNA_1013 (.A(\spiking_network_top_uut.all_data_out[902] ));
 sg13g2_antennanp ANTENNA_1014 (.A(\spiking_network_top_uut.all_data_out[902] ));
 sg13g2_antennanp ANTENNA_1015 (.A(\spiking_network_top_uut.all_data_out[902] ));
 sg13g2_antennanp ANTENNA_1016 (.A(\spiking_network_top_uut.all_data_out[903] ));
 sg13g2_antennanp ANTENNA_1017 (.A(\spiking_network_top_uut.all_data_out[903] ));
 sg13g2_antennanp ANTENNA_1018 (.A(\spiking_network_top_uut.all_data_out[903] ));
 sg13g2_antennanp ANTENNA_1019 (.A(\spiking_network_top_uut.all_data_out[903] ));
 sg13g2_antennanp ANTENNA_1020 (.A(\spiking_network_top_uut.all_data_out[903] ));
 sg13g2_antennanp ANTENNA_1021 (.A(\spiking_network_top_uut.all_data_out[903] ));
 sg13g2_antennanp ANTENNA_1022 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_1023 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_1024 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_1025 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_1026 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_1027 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_1028 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_1029 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.spike_out ));
 sg13g2_antennanp ANTENNA_1030 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.spike_out ));
 sg13g2_antennanp ANTENNA_1031 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.spike_out ));
 sg13g2_antennanp ANTENNA_1032 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_1033 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_1034 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_1035 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_1036 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_1037 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_1038 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_1039 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_1040 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_1041 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_1042 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_1043 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_1044 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_1045 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_1046 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_1047 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_1048 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_1049 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_1050 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_1051 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_1052 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_1053 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_1054 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_1055 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_1056 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_1057 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_1058 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_1059 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_1060 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_1061 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_1062 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_1063 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_1064 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_1065 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_1066 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_1067 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[3].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_1068 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_1069 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_1070 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_1071 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_1072 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_1073 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_1074 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_1075 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_1076 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_1077 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_1078 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_reg1 ));
 sg13g2_antennanp ANTENNA_1079 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_reg1 ));
 sg13g2_antennanp ANTENNA_1080 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_reg1 ));
 sg13g2_antennanp ANTENNA_1081 (.A(net3658));
 sg13g2_antennanp ANTENNA_1082 (.A(net3658));
 sg13g2_antennanp ANTENNA_1083 (.A(net3658));
 sg13g2_antennanp ANTENNA_1084 (.A(net3658));
 sg13g2_antennanp ANTENNA_1085 (.A(net3658));
 sg13g2_antennanp ANTENNA_1086 (.A(net3658));
 sg13g2_antennanp ANTENNA_1087 (.A(net3728));
 sg13g2_antennanp ANTENNA_1088 (.A(net3728));
 sg13g2_antennanp ANTENNA_1089 (.A(net3728));
 sg13g2_antennanp ANTENNA_1090 (.A(net3728));
 sg13g2_antennanp ANTENNA_1091 (.A(net3728));
 sg13g2_antennanp ANTENNA_1092 (.A(net3728));
 sg13g2_antennanp ANTENNA_1093 (.A(net3728));
 sg13g2_antennanp ANTENNA_1094 (.A(net3728));
 sg13g2_antennanp ANTENNA_1095 (.A(net4136));
 sg13g2_antennanp ANTENNA_1096 (.A(net4136));
 sg13g2_antennanp ANTENNA_1097 (.A(net4136));
 sg13g2_antennanp ANTENNA_1098 (.A(net4136));
 sg13g2_antennanp ANTENNA_1099 (.A(net4136));
 sg13g2_antennanp ANTENNA_1100 (.A(net4162));
 sg13g2_antennanp ANTENNA_1101 (.A(net4162));
 sg13g2_antennanp ANTENNA_1102 (.A(net4162));
 sg13g2_antennanp ANTENNA_1103 (.A(net4162));
 sg13g2_antennanp ANTENNA_1104 (.A(net4162));
 sg13g2_antennanp ANTENNA_1105 (.A(net4162));
 sg13g2_antennanp ANTENNA_1106 (.A(net4162));
 sg13g2_antennanp ANTENNA_1107 (.A(net4162));
 sg13g2_antennanp ANTENNA_1108 (.A(net4162));
 sg13g2_antennanp ANTENNA_1109 (.A(net4162));
 sg13g2_antennanp ANTENNA_1110 (.A(net4162));
 sg13g2_antennanp ANTENNA_1111 (.A(net4162));
 sg13g2_antennanp ANTENNA_1112 (.A(net4162));
 sg13g2_antennanp ANTENNA_1113 (.A(net4275));
 sg13g2_antennanp ANTENNA_1114 (.A(net4275));
 sg13g2_antennanp ANTENNA_1115 (.A(net4275));
 sg13g2_antennanp ANTENNA_1116 (.A(net4275));
 sg13g2_antennanp ANTENNA_1117 (.A(net4275));
 sg13g2_antennanp ANTENNA_1118 (.A(net4275));
 sg13g2_antennanp ANTENNA_1119 (.A(net4275));
 sg13g2_antennanp ANTENNA_1120 (.A(net4275));
 sg13g2_antennanp ANTENNA_1121 (.A(net4275));
 sg13g2_antennanp ANTENNA_1122 (.A(net4275));
 sg13g2_antennanp ANTENNA_1123 (.A(net4275));
 sg13g2_antennanp ANTENNA_1124 (.A(net4275));
 sg13g2_antennanp ANTENNA_1125 (.A(net4275));
 sg13g2_antennanp ANTENNA_1126 (.A(net4275));
 sg13g2_antennanp ANTENNA_1127 (.A(net4275));
 sg13g2_antennanp ANTENNA_1128 (.A(net4275));
 sg13g2_antennanp ANTENNA_1129 (.A(net4379));
 sg13g2_antennanp ANTENNA_1130 (.A(net4379));
 sg13g2_antennanp ANTENNA_1131 (.A(net4379));
 sg13g2_antennanp ANTENNA_1132 (.A(net4379));
 sg13g2_antennanp ANTENNA_1133 (.A(net4379));
 sg13g2_antennanp ANTENNA_1134 (.A(net4379));
 sg13g2_antennanp ANTENNA_1135 (.A(net4379));
 sg13g2_antennanp ANTENNA_1136 (.A(net4379));
 sg13g2_antennanp ANTENNA_1137 (.A(net4709));
 sg13g2_antennanp ANTENNA_1138 (.A(net4709));
 sg13g2_antennanp ANTENNA_1139 (.A(net4709));
 sg13g2_antennanp ANTENNA_1140 (.A(net4709));
 sg13g2_antennanp ANTENNA_1141 (.A(net4709));
 sg13g2_antennanp ANTENNA_1142 (.A(net4709));
 sg13g2_antennanp ANTENNA_1143 (.A(net4709));
 sg13g2_antennanp ANTENNA_1144 (.A(net4709));
 sg13g2_antennanp ANTENNA_1145 (.A(net4709));
 sg13g2_antennanp ANTENNA_1146 (.A(net4709));
 sg13g2_antennanp ANTENNA_1147 (.A(net4709));
 sg13g2_antennanp ANTENNA_1148 (.A(net4709));
 sg13g2_antennanp ANTENNA_1149 (.A(net4709));
 sg13g2_antennanp ANTENNA_1150 (.A(net2));
 sg13g2_antennanp ANTENNA_1151 (.A(net4));
 sg13g2_antennanp ANTENNA_1152 (.A(net6));
 sg13g2_antennanp ANTENNA_1153 (.A(net7));
 sg13g2_antennanp ANTENNA_1154 (.A(net8));
 sg13g2_antennanp ANTENNA_1155 (.A(net9));
 sg13g2_antennanp ANTENNA_1156 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_1157 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_1158 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_1159 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_1160 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_1161 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_1162 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_1163 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_1164 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_1165 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_1166 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_1167 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_1168 (.A(_00026_));
 sg13g2_antennanp ANTENNA_1169 (.A(_00026_));
 sg13g2_antennanp ANTENNA_1170 (.A(_00026_));
 sg13g2_antennanp ANTENNA_1171 (.A(_00026_));
 sg13g2_antennanp ANTENNA_1172 (.A(_00146_));
 sg13g2_antennanp ANTENNA_1173 (.A(_00148_));
 sg13g2_antennanp ANTENNA_1174 (.A(_00188_));
 sg13g2_antennanp ANTENNA_1175 (.A(_00197_));
 sg13g2_antennanp ANTENNA_1176 (.A(_00199_));
 sg13g2_antennanp ANTENNA_1177 (.A(_00201_));
 sg13g2_antennanp ANTENNA_1178 (.A(_00209_));
 sg13g2_antennanp ANTENNA_1179 (.A(_00213_));
 sg13g2_antennanp ANTENNA_1180 (.A(_00217_));
 sg13g2_antennanp ANTENNA_1181 (.A(_00226_));
 sg13g2_antennanp ANTENNA_1182 (.A(_00232_));
 sg13g2_antennanp ANTENNA_1183 (.A(_00251_));
 sg13g2_antennanp ANTENNA_1184 (.A(_00258_));
 sg13g2_antennanp ANTENNA_1185 (.A(_00259_));
 sg13g2_antennanp ANTENNA_1186 (.A(_00271_));
 sg13g2_antennanp ANTENNA_1187 (.A(_00283_));
 sg13g2_antennanp ANTENNA_1188 (.A(_00284_));
 sg13g2_antennanp ANTENNA_1189 (.A(_00299_));
 sg13g2_antennanp ANTENNA_1190 (.A(_00328_));
 sg13g2_antennanp ANTENNA_1191 (.A(_00329_));
 sg13g2_antennanp ANTENNA_1192 (.A(_00390_));
 sg13g2_antennanp ANTENNA_1193 (.A(_00391_));
 sg13g2_antennanp ANTENNA_1194 (.A(_00411_));
 sg13g2_antennanp ANTENNA_1195 (.A(_00415_));
 sg13g2_antennanp ANTENNA_1196 (.A(_00419_));
 sg13g2_antennanp ANTENNA_1197 (.A(_02216_));
 sg13g2_antennanp ANTENNA_1198 (.A(_02483_));
 sg13g2_antennanp ANTENNA_1199 (.A(_02483_));
 sg13g2_antennanp ANTENNA_1200 (.A(_02483_));
 sg13g2_antennanp ANTENNA_1201 (.A(_02483_));
 sg13g2_antennanp ANTENNA_1202 (.A(_02483_));
 sg13g2_antennanp ANTENNA_1203 (.A(_02483_));
 sg13g2_antennanp ANTENNA_1204 (.A(_02483_));
 sg13g2_antennanp ANTENNA_1205 (.A(_02483_));
 sg13g2_antennanp ANTENNA_1206 (.A(_02483_));
 sg13g2_antennanp ANTENNA_1207 (.A(_02484_));
 sg13g2_antennanp ANTENNA_1208 (.A(_02484_));
 sg13g2_antennanp ANTENNA_1209 (.A(_02484_));
 sg13g2_antennanp ANTENNA_1210 (.A(_02484_));
 sg13g2_antennanp ANTENNA_1211 (.A(_02494_));
 sg13g2_antennanp ANTENNA_1212 (.A(_02494_));
 sg13g2_antennanp ANTENNA_1213 (.A(_02494_));
 sg13g2_antennanp ANTENNA_1214 (.A(_02494_));
 sg13g2_antennanp ANTENNA_1215 (.A(_02495_));
 sg13g2_antennanp ANTENNA_1216 (.A(_02495_));
 sg13g2_antennanp ANTENNA_1217 (.A(_02495_));
 sg13g2_antennanp ANTENNA_1218 (.A(_02495_));
 sg13g2_antennanp ANTENNA_1219 (.A(_02495_));
 sg13g2_antennanp ANTENNA_1220 (.A(_02495_));
 sg13g2_antennanp ANTENNA_1221 (.A(_02495_));
 sg13g2_antennanp ANTENNA_1222 (.A(_02495_));
 sg13g2_antennanp ANTENNA_1223 (.A(_02495_));
 sg13g2_antennanp ANTENNA_1224 (.A(_02509_));
 sg13g2_antennanp ANTENNA_1225 (.A(_02509_));
 sg13g2_antennanp ANTENNA_1226 (.A(_02509_));
 sg13g2_antennanp ANTENNA_1227 (.A(_02509_));
 sg13g2_antennanp ANTENNA_1228 (.A(_02777_));
 sg13g2_antennanp ANTENNA_1229 (.A(_02777_));
 sg13g2_antennanp ANTENNA_1230 (.A(_02777_));
 sg13g2_antennanp ANTENNA_1231 (.A(_02777_));
 sg13g2_antennanp ANTENNA_1232 (.A(_02991_));
 sg13g2_antennanp ANTENNA_1233 (.A(_02991_));
 sg13g2_antennanp ANTENNA_1234 (.A(_02991_));
 sg13g2_antennanp ANTENNA_1235 (.A(_02991_));
 sg13g2_antennanp ANTENNA_1236 (.A(_02991_));
 sg13g2_antennanp ANTENNA_1237 (.A(_02991_));
 sg13g2_antennanp ANTENNA_1238 (.A(_02991_));
 sg13g2_antennanp ANTENNA_1239 (.A(_02991_));
 sg13g2_antennanp ANTENNA_1240 (.A(_02991_));
 sg13g2_antennanp ANTENNA_1241 (.A(_03215_));
 sg13g2_antennanp ANTENNA_1242 (.A(_03215_));
 sg13g2_antennanp ANTENNA_1243 (.A(_03215_));
 sg13g2_antennanp ANTENNA_1244 (.A(_03215_));
 sg13g2_antennanp ANTENNA_1245 (.A(_03215_));
 sg13g2_antennanp ANTENNA_1246 (.A(_03215_));
 sg13g2_antennanp ANTENNA_1247 (.A(_03215_));
 sg13g2_antennanp ANTENNA_1248 (.A(_03215_));
 sg13g2_antennanp ANTENNA_1249 (.A(_03215_));
 sg13g2_antennanp ANTENNA_1250 (.A(_03215_));
 sg13g2_antennanp ANTENNA_1251 (.A(_03215_));
 sg13g2_antennanp ANTENNA_1252 (.A(_03215_));
 sg13g2_antennanp ANTENNA_1253 (.A(_03215_));
 sg13g2_antennanp ANTENNA_1254 (.A(_03215_));
 sg13g2_antennanp ANTENNA_1255 (.A(_03215_));
 sg13g2_antennanp ANTENNA_1256 (.A(_03215_));
 sg13g2_antennanp ANTENNA_1257 (.A(_03215_));
 sg13g2_antennanp ANTENNA_1258 (.A(_03509_));
 sg13g2_antennanp ANTENNA_1259 (.A(_03518_));
 sg13g2_antennanp ANTENNA_1260 (.A(_03522_));
 sg13g2_antennanp ANTENNA_1261 (.A(_03534_));
 sg13g2_antennanp ANTENNA_1262 (.A(_03543_));
 sg13g2_antennanp ANTENNA_1263 (.A(_03549_));
 sg13g2_antennanp ANTENNA_1264 (.A(_03550_));
 sg13g2_antennanp ANTENNA_1265 (.A(_03551_));
 sg13g2_antennanp ANTENNA_1266 (.A(_03567_));
 sg13g2_antennanp ANTENNA_1267 (.A(_03571_));
 sg13g2_antennanp ANTENNA_1268 (.A(_03573_));
 sg13g2_antennanp ANTENNA_1269 (.A(_03574_));
 sg13g2_antennanp ANTENNA_1270 (.A(_03576_));
 sg13g2_antennanp ANTENNA_1271 (.A(_03578_));
 sg13g2_antennanp ANTENNA_1272 (.A(_03609_));
 sg13g2_antennanp ANTENNA_1273 (.A(_03613_));
 sg13g2_antennanp ANTENNA_1274 (.A(_03614_));
 sg13g2_antennanp ANTENNA_1275 (.A(_03622_));
 sg13g2_antennanp ANTENNA_1276 (.A(_03625_));
 sg13g2_antennanp ANTENNA_1277 (.A(_03648_));
 sg13g2_antennanp ANTENNA_1278 (.A(_03650_));
 sg13g2_antennanp ANTENNA_1279 (.A(_03651_));
 sg13g2_antennanp ANTENNA_1280 (.A(_03652_));
 sg13g2_antennanp ANTENNA_1281 (.A(_03654_));
 sg13g2_antennanp ANTENNA_1282 (.A(_03794_));
 sg13g2_antennanp ANTENNA_1283 (.A(_03794_));
 sg13g2_antennanp ANTENNA_1284 (.A(_03794_));
 sg13g2_antennanp ANTENNA_1285 (.A(_03794_));
 sg13g2_antennanp ANTENNA_1286 (.A(_03794_));
 sg13g2_antennanp ANTENNA_1287 (.A(_03794_));
 sg13g2_antennanp ANTENNA_1288 (.A(_03794_));
 sg13g2_antennanp ANTENNA_1289 (.A(_03794_));
 sg13g2_antennanp ANTENNA_1290 (.A(_03794_));
 sg13g2_antennanp ANTENNA_1291 (.A(_03794_));
 sg13g2_antennanp ANTENNA_1292 (.A(_03794_));
 sg13g2_antennanp ANTENNA_1293 (.A(_03794_));
 sg13g2_antennanp ANTENNA_1294 (.A(_03794_));
 sg13g2_antennanp ANTENNA_1295 (.A(_03794_));
 sg13g2_antennanp ANTENNA_1296 (.A(_03794_));
 sg13g2_antennanp ANTENNA_1297 (.A(_03794_));
 sg13g2_antennanp ANTENNA_1298 (.A(_03794_));
 sg13g2_antennanp ANTENNA_1299 (.A(_03794_));
 sg13g2_antennanp ANTENNA_1300 (.A(_03794_));
 sg13g2_antennanp ANTENNA_1301 (.A(_03794_));
 sg13g2_antennanp ANTENNA_1302 (.A(_03893_));
 sg13g2_antennanp ANTENNA_1303 (.A(_03906_));
 sg13g2_antennanp ANTENNA_1304 (.A(_03913_));
 sg13g2_antennanp ANTENNA_1305 (.A(_03988_));
 sg13g2_antennanp ANTENNA_1306 (.A(_03990_));
 sg13g2_antennanp ANTENNA_1307 (.A(_03993_));
 sg13g2_antennanp ANTENNA_1308 (.A(_03999_));
 sg13g2_antennanp ANTENNA_1309 (.A(_04005_));
 sg13g2_antennanp ANTENNA_1310 (.A(_04025_));
 sg13g2_antennanp ANTENNA_1311 (.A(_04028_));
 sg13g2_antennanp ANTENNA_1312 (.A(_04043_));
 sg13g2_antennanp ANTENNA_1313 (.A(_04046_));
 sg13g2_antennanp ANTENNA_1314 (.A(_04092_));
 sg13g2_antennanp ANTENNA_1315 (.A(_04114_));
 sg13g2_antennanp ANTENNA_1316 (.A(_04130_));
 sg13g2_antennanp ANTENNA_1317 (.A(_04131_));
 sg13g2_antennanp ANTENNA_1318 (.A(_04132_));
 sg13g2_antennanp ANTENNA_1319 (.A(_04148_));
 sg13g2_antennanp ANTENNA_1320 (.A(_04180_));
 sg13g2_antennanp ANTENNA_1321 (.A(_04194_));
 sg13g2_antennanp ANTENNA_1322 (.A(_04202_));
 sg13g2_antennanp ANTENNA_1323 (.A(_04213_));
 sg13g2_antennanp ANTENNA_1324 (.A(_04216_));
 sg13g2_antennanp ANTENNA_1325 (.A(_04221_));
 sg13g2_antennanp ANTENNA_1326 (.A(_04231_));
 sg13g2_antennanp ANTENNA_1327 (.A(_04238_));
 sg13g2_antennanp ANTENNA_1328 (.A(_04270_));
 sg13g2_antennanp ANTENNA_1329 (.A(_04271_));
 sg13g2_antennanp ANTENNA_1330 (.A(_04280_));
 sg13g2_antennanp ANTENNA_1331 (.A(_04289_));
 sg13g2_antennanp ANTENNA_1332 (.A(_04312_));
 sg13g2_antennanp ANTENNA_1333 (.A(_04319_));
 sg13g2_antennanp ANTENNA_1334 (.A(_04352_));
 sg13g2_antennanp ANTENNA_1335 (.A(_04362_));
 sg13g2_antennanp ANTENNA_1336 (.A(_04374_));
 sg13g2_antennanp ANTENNA_1337 (.A(_04401_));
 sg13g2_antennanp ANTENNA_1338 (.A(_04403_));
 sg13g2_antennanp ANTENNA_1339 (.A(_04410_));
 sg13g2_antennanp ANTENNA_1340 (.A(_04415_));
 sg13g2_antennanp ANTENNA_1341 (.A(_04417_));
 sg13g2_antennanp ANTENNA_1342 (.A(_04436_));
 sg13g2_antennanp ANTENNA_1343 (.A(_04450_));
 sg13g2_antennanp ANTENNA_1344 (.A(_04480_));
 sg13g2_antennanp ANTENNA_1345 (.A(_04498_));
 sg13g2_antennanp ANTENNA_1346 (.A(_04500_));
 sg13g2_antennanp ANTENNA_1347 (.A(_04504_));
 sg13g2_antennanp ANTENNA_1348 (.A(_04508_));
 sg13g2_antennanp ANTENNA_1349 (.A(_04511_));
 sg13g2_antennanp ANTENNA_1350 (.A(_04523_));
 sg13g2_antennanp ANTENNA_1351 (.A(_04543_));
 sg13g2_antennanp ANTENNA_1352 (.A(_04559_));
 sg13g2_antennanp ANTENNA_1353 (.A(_04562_));
 sg13g2_antennanp ANTENNA_1354 (.A(_04579_));
 sg13g2_antennanp ANTENNA_1355 (.A(_04580_));
 sg13g2_antennanp ANTENNA_1356 (.A(_04584_));
 sg13g2_antennanp ANTENNA_1357 (.A(_05709_));
 sg13g2_antennanp ANTENNA_1358 (.A(_05709_));
 sg13g2_antennanp ANTENNA_1359 (.A(_05709_));
 sg13g2_antennanp ANTENNA_1360 (.A(_05709_));
 sg13g2_antennanp ANTENNA_1361 (.A(_06082_));
 sg13g2_antennanp ANTENNA_1362 (.A(_06284_));
 sg13g2_antennanp ANTENNA_1363 (.A(_06284_));
 sg13g2_antennanp ANTENNA_1364 (.A(_06284_));
 sg13g2_antennanp ANTENNA_1365 (.A(_06284_));
 sg13g2_antennanp ANTENNA_1366 (.A(_06286_));
 sg13g2_antennanp ANTENNA_1367 (.A(_06286_));
 sg13g2_antennanp ANTENNA_1368 (.A(_06286_));
 sg13g2_antennanp ANTENNA_1369 (.A(_06286_));
 sg13g2_antennanp ANTENNA_1370 (.A(_06625_));
 sg13g2_antennanp ANTENNA_1371 (.A(_06625_));
 sg13g2_antennanp ANTENNA_1372 (.A(_06625_));
 sg13g2_antennanp ANTENNA_1373 (.A(_06625_));
 sg13g2_antennanp ANTENNA_1374 (.A(_07721_));
 sg13g2_antennanp ANTENNA_1375 (.A(_07721_));
 sg13g2_antennanp ANTENNA_1376 (.A(_07721_));
 sg13g2_antennanp ANTENNA_1377 (.A(_07721_));
 sg13g2_antennanp ANTENNA_1378 (.A(_08106_));
 sg13g2_antennanp ANTENNA_1379 (.A(_08106_));
 sg13g2_antennanp ANTENNA_1380 (.A(_08106_));
 sg13g2_antennanp ANTENNA_1381 (.A(_08106_));
 sg13g2_antennanp ANTENNA_1382 (.A(_08570_));
 sg13g2_antennanp ANTENNA_1383 (.A(_08570_));
 sg13g2_antennanp ANTENNA_1384 (.A(_08570_));
 sg13g2_antennanp ANTENNA_1385 (.A(_08570_));
 sg13g2_antennanp ANTENNA_1386 (.A(_08572_));
 sg13g2_antennanp ANTENNA_1387 (.A(_08572_));
 sg13g2_antennanp ANTENNA_1388 (.A(_08572_));
 sg13g2_antennanp ANTENNA_1389 (.A(_08572_));
 sg13g2_antennanp ANTENNA_1390 (.A(_08572_));
 sg13g2_antennanp ANTENNA_1391 (.A(_08572_));
 sg13g2_antennanp ANTENNA_1392 (.A(_08572_));
 sg13g2_antennanp ANTENNA_1393 (.A(_08572_));
 sg13g2_antennanp ANTENNA_1394 (.A(_08572_));
 sg13g2_antennanp ANTENNA_1395 (.A(_08572_));
 sg13g2_antennanp ANTENNA_1396 (.A(_08572_));
 sg13g2_antennanp ANTENNA_1397 (.A(_08572_));
 sg13g2_antennanp ANTENNA_1398 (.A(_08849_));
 sg13g2_antennanp ANTENNA_1399 (.A(_08849_));
 sg13g2_antennanp ANTENNA_1400 (.A(_08849_));
 sg13g2_antennanp ANTENNA_1401 (.A(_08849_));
 sg13g2_antennanp ANTENNA_1402 (.A(_08849_));
 sg13g2_antennanp ANTENNA_1403 (.A(_08849_));
 sg13g2_antennanp ANTENNA_1404 (.A(_08849_));
 sg13g2_antennanp ANTENNA_1405 (.A(_08849_));
 sg13g2_antennanp ANTENNA_1406 (.A(_08849_));
 sg13g2_antennanp ANTENNA_1407 (.A(_08860_));
 sg13g2_antennanp ANTENNA_1408 (.A(_08860_));
 sg13g2_antennanp ANTENNA_1409 (.A(_08860_));
 sg13g2_antennanp ANTENNA_1410 (.A(_08860_));
 sg13g2_antennanp ANTENNA_1411 (.A(\spiking_network_top_uut.all_data_out[273] ));
 sg13g2_antennanp ANTENNA_1412 (.A(\spiking_network_top_uut.all_data_out[273] ));
 sg13g2_antennanp ANTENNA_1413 (.A(\spiking_network_top_uut.all_data_out[273] ));
 sg13g2_antennanp ANTENNA_1414 (.A(\spiking_network_top_uut.all_data_out[294] ));
 sg13g2_antennanp ANTENNA_1415 (.A(\spiking_network_top_uut.all_data_out[294] ));
 sg13g2_antennanp ANTENNA_1416 (.A(\spiking_network_top_uut.all_data_out[294] ));
 sg13g2_antennanp ANTENNA_1417 (.A(\spiking_network_top_uut.all_data_out[294] ));
 sg13g2_antennanp ANTENNA_1418 (.A(\spiking_network_top_uut.all_data_out[294] ));
 sg13g2_antennanp ANTENNA_1419 (.A(\spiking_network_top_uut.all_data_out[294] ));
 sg13g2_antennanp ANTENNA_1420 (.A(\spiking_network_top_uut.all_data_out[294] ));
 sg13g2_antennanp ANTENNA_1421 (.A(\spiking_network_top_uut.all_data_out[294] ));
 sg13g2_antennanp ANTENNA_1422 (.A(\spiking_network_top_uut.all_data_out[294] ));
 sg13g2_antennanp ANTENNA_1423 (.A(\spiking_network_top_uut.all_data_out[307] ));
 sg13g2_antennanp ANTENNA_1424 (.A(\spiking_network_top_uut.all_data_out[307] ));
 sg13g2_antennanp ANTENNA_1425 (.A(\spiking_network_top_uut.all_data_out[307] ));
 sg13g2_antennanp ANTENNA_1426 (.A(\spiking_network_top_uut.all_data_out[308] ));
 sg13g2_antennanp ANTENNA_1427 (.A(\spiking_network_top_uut.all_data_out[308] ));
 sg13g2_antennanp ANTENNA_1428 (.A(\spiking_network_top_uut.all_data_out[308] ));
 sg13g2_antennanp ANTENNA_1429 (.A(\spiking_network_top_uut.all_data_out[308] ));
 sg13g2_antennanp ANTENNA_1430 (.A(\spiking_network_top_uut.all_data_out[311] ));
 sg13g2_antennanp ANTENNA_1431 (.A(\spiking_network_top_uut.all_data_out[311] ));
 sg13g2_antennanp ANTENNA_1432 (.A(\spiking_network_top_uut.all_data_out[311] ));
 sg13g2_antennanp ANTENNA_1433 (.A(\spiking_network_top_uut.all_data_out[311] ));
 sg13g2_antennanp ANTENNA_1434 (.A(\spiking_network_top_uut.all_data_out[311] ));
 sg13g2_antennanp ANTENNA_1435 (.A(\spiking_network_top_uut.all_data_out[311] ));
 sg13g2_antennanp ANTENNA_1436 (.A(\spiking_network_top_uut.all_data_out[311] ));
 sg13g2_antennanp ANTENNA_1437 (.A(\spiking_network_top_uut.all_data_out[311] ));
 sg13g2_antennanp ANTENNA_1438 (.A(\spiking_network_top_uut.all_data_out[311] ));
 sg13g2_antennanp ANTENNA_1439 (.A(\spiking_network_top_uut.all_data_out[330] ));
 sg13g2_antennanp ANTENNA_1440 (.A(\spiking_network_top_uut.all_data_out[330] ));
 sg13g2_antennanp ANTENNA_1441 (.A(\spiking_network_top_uut.all_data_out[330] ));
 sg13g2_antennanp ANTENNA_1442 (.A(\spiking_network_top_uut.all_data_out[330] ));
 sg13g2_antennanp ANTENNA_1443 (.A(\spiking_network_top_uut.all_data_out[584] ));
 sg13g2_antennanp ANTENNA_1444 (.A(\spiking_network_top_uut.all_data_out[584] ));
 sg13g2_antennanp ANTENNA_1445 (.A(\spiking_network_top_uut.all_data_out[584] ));
 sg13g2_antennanp ANTENNA_1446 (.A(\spiking_network_top_uut.all_data_out[584] ));
 sg13g2_antennanp ANTENNA_1447 (.A(\spiking_network_top_uut.all_data_out[584] ));
 sg13g2_antennanp ANTENNA_1448 (.A(\spiking_network_top_uut.all_data_out[584] ));
 sg13g2_antennanp ANTENNA_1449 (.A(\spiking_network_top_uut.all_data_out[584] ));
 sg13g2_antennanp ANTENNA_1450 (.A(\spiking_network_top_uut.all_data_out[584] ));
 sg13g2_antennanp ANTENNA_1451 (.A(\spiking_network_top_uut.all_data_out[584] ));
 sg13g2_antennanp ANTENNA_1452 (.A(\spiking_network_top_uut.all_data_out[584] ));
 sg13g2_antennanp ANTENNA_1453 (.A(\spiking_network_top_uut.all_data_out[584] ));
 sg13g2_antennanp ANTENNA_1454 (.A(\spiking_network_top_uut.all_data_out[584] ));
 sg13g2_antennanp ANTENNA_1455 (.A(\spiking_network_top_uut.all_data_out[584] ));
 sg13g2_antennanp ANTENNA_1456 (.A(\spiking_network_top_uut.all_data_out[584] ));
 sg13g2_antennanp ANTENNA_1457 (.A(\spiking_network_top_uut.all_data_out[584] ));
 sg13g2_antennanp ANTENNA_1458 (.A(\spiking_network_top_uut.all_data_out[584] ));
 sg13g2_antennanp ANTENNA_1459 (.A(\spiking_network_top_uut.all_data_out[76] ));
 sg13g2_antennanp ANTENNA_1460 (.A(\spiking_network_top_uut.all_data_out[76] ));
 sg13g2_antennanp ANTENNA_1461 (.A(\spiking_network_top_uut.all_data_out[76] ));
 sg13g2_antennanp ANTENNA_1462 (.A(\spiking_network_top_uut.all_data_out[76] ));
 sg13g2_antennanp ANTENNA_1463 (.A(\spiking_network_top_uut.all_data_out[855] ));
 sg13g2_antennanp ANTENNA_1464 (.A(\spiking_network_top_uut.all_data_out[855] ));
 sg13g2_antennanp ANTENNA_1465 (.A(\spiking_network_top_uut.all_data_out[855] ));
 sg13g2_antennanp ANTENNA_1466 (.A(\spiking_network_top_uut.all_data_out[896] ));
 sg13g2_antennanp ANTENNA_1467 (.A(\spiking_network_top_uut.all_data_out[896] ));
 sg13g2_antennanp ANTENNA_1468 (.A(\spiking_network_top_uut.all_data_out[896] ));
 sg13g2_antennanp ANTENNA_1469 (.A(\spiking_network_top_uut.all_data_out[896] ));
 sg13g2_antennanp ANTENNA_1470 (.A(\spiking_network_top_uut.all_data_out[896] ));
 sg13g2_antennanp ANTENNA_1471 (.A(\spiking_network_top_uut.all_data_out[896] ));
 sg13g2_antennanp ANTENNA_1472 (.A(\spiking_network_top_uut.all_data_out[896] ));
 sg13g2_antennanp ANTENNA_1473 (.A(\spiking_network_top_uut.all_data_out[896] ));
 sg13g2_antennanp ANTENNA_1474 (.A(\spiking_network_top_uut.all_data_out[896] ));
 sg13g2_antennanp ANTENNA_1475 (.A(\spiking_network_top_uut.all_data_out[897] ));
 sg13g2_antennanp ANTENNA_1476 (.A(\spiking_network_top_uut.all_data_out[897] ));
 sg13g2_antennanp ANTENNA_1477 (.A(\spiking_network_top_uut.all_data_out[897] ));
 sg13g2_antennanp ANTENNA_1478 (.A(\spiking_network_top_uut.all_data_out[897] ));
 sg13g2_antennanp ANTENNA_1479 (.A(\spiking_network_top_uut.all_data_out[897] ));
 sg13g2_antennanp ANTENNA_1480 (.A(\spiking_network_top_uut.all_data_out[897] ));
 sg13g2_antennanp ANTENNA_1481 (.A(\spiking_network_top_uut.all_data_out[897] ));
 sg13g2_antennanp ANTENNA_1482 (.A(\spiking_network_top_uut.all_data_out[897] ));
 sg13g2_antennanp ANTENNA_1483 (.A(\spiking_network_top_uut.all_data_out[897] ));
 sg13g2_antennanp ANTENNA_1484 (.A(\spiking_network_top_uut.all_data_out[898] ));
 sg13g2_antennanp ANTENNA_1485 (.A(\spiking_network_top_uut.all_data_out[898] ));
 sg13g2_antennanp ANTENNA_1486 (.A(\spiking_network_top_uut.all_data_out[898] ));
 sg13g2_antennanp ANTENNA_1487 (.A(\spiking_network_top_uut.all_data_out[898] ));
 sg13g2_antennanp ANTENNA_1488 (.A(\spiking_network_top_uut.all_data_out[898] ));
 sg13g2_antennanp ANTENNA_1489 (.A(\spiking_network_top_uut.all_data_out[898] ));
 sg13g2_antennanp ANTENNA_1490 (.A(\spiking_network_top_uut.all_data_out[898] ));
 sg13g2_antennanp ANTENNA_1491 (.A(\spiking_network_top_uut.all_data_out[898] ));
 sg13g2_antennanp ANTENNA_1492 (.A(\spiking_network_top_uut.all_data_out[898] ));
 sg13g2_antennanp ANTENNA_1493 (.A(\spiking_network_top_uut.all_data_out[899] ));
 sg13g2_antennanp ANTENNA_1494 (.A(\spiking_network_top_uut.all_data_out[899] ));
 sg13g2_antennanp ANTENNA_1495 (.A(\spiking_network_top_uut.all_data_out[899] ));
 sg13g2_antennanp ANTENNA_1496 (.A(\spiking_network_top_uut.all_data_out[899] ));
 sg13g2_antennanp ANTENNA_1497 (.A(\spiking_network_top_uut.all_data_out[899] ));
 sg13g2_antennanp ANTENNA_1498 (.A(\spiking_network_top_uut.all_data_out[899] ));
 sg13g2_antennanp ANTENNA_1499 (.A(\spiking_network_top_uut.all_data_out[902] ));
 sg13g2_antennanp ANTENNA_1500 (.A(\spiking_network_top_uut.all_data_out[902] ));
 sg13g2_antennanp ANTENNA_1501 (.A(\spiking_network_top_uut.all_data_out[902] ));
 sg13g2_antennanp ANTENNA_1502 (.A(\spiking_network_top_uut.all_data_out[902] ));
 sg13g2_antennanp ANTENNA_1503 (.A(\spiking_network_top_uut.all_data_out[902] ));
 sg13g2_antennanp ANTENNA_1504 (.A(\spiking_network_top_uut.all_data_out[902] ));
 sg13g2_antennanp ANTENNA_1505 (.A(\spiking_network_top_uut.all_data_out[902] ));
 sg13g2_antennanp ANTENNA_1506 (.A(\spiking_network_top_uut.all_data_out[902] ));
 sg13g2_antennanp ANTENNA_1507 (.A(\spiking_network_top_uut.all_data_out[902] ));
 sg13g2_antennanp ANTENNA_1508 (.A(\spiking_network_top_uut.all_data_out[902] ));
 sg13g2_antennanp ANTENNA_1509 (.A(\spiking_network_top_uut.all_data_out[903] ));
 sg13g2_antennanp ANTENNA_1510 (.A(\spiking_network_top_uut.all_data_out[903] ));
 sg13g2_antennanp ANTENNA_1511 (.A(\spiking_network_top_uut.all_data_out[903] ));
 sg13g2_antennanp ANTENNA_1512 (.A(\spiking_network_top_uut.all_data_out[903] ));
 sg13g2_antennanp ANTENNA_1513 (.A(\spiking_network_top_uut.all_data_out[903] ));
 sg13g2_antennanp ANTENNA_1514 (.A(\spiking_network_top_uut.all_data_out[903] ));
 sg13g2_antennanp ANTENNA_1515 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_1516 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_1517 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[0].neuron_inst.neuron_delay_gen[6].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_1518 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_1519 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_1520 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_1521 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[1].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_1522 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.spike_out ));
 sg13g2_antennanp ANTENNA_1523 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.spike_out ));
 sg13g2_antennanp ANTENNA_1524 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.lif_neuron_inst.lif_neuron_inst.spike_out ));
 sg13g2_antennanp ANTENNA_1525 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_1526 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_1527 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_1528 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_1529 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_1530 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_1531 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_1532 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[2].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_1533 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_1534 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_1535 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[4].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_1536 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_1537 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_1538 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_1539 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.neuron_delay_gen[1].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_1540 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_1541 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_1542 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_1543 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[5].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_1544 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_1545 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_1546 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_1547 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer1.neuron_gen[6].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_1548 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_1549 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_1550 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[0].neuron_inst.neuron_delay_gen[7].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_1551 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_1552 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[1].neuron_inst.neuron_delay_gen[4].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_1553 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_1554 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_1555 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_1556 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[4].neuron_inst.neuron_delay_gen[3].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_1557 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_1558 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[5].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_1559 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_1560 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[6].neuron_inst.neuron_delay_gen[2].neuron_delay_inst.sync_dout ));
 sg13g2_antennanp ANTENNA_1561 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_reg1 ));
 sg13g2_antennanp ANTENNA_1562 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_reg1 ));
 sg13g2_antennanp ANTENNA_1563 (.A(\spiking_network_top_uut.snn_inst.three_layer_network_inst.layer2.neuron_gen[7].neuron_inst.neuron_delay_gen[0].neuron_delay_inst.sync_reg1 ));
 sg13g2_antennanp ANTENNA_1564 (.A(net3728));
 sg13g2_antennanp ANTENNA_1565 (.A(net3728));
 sg13g2_antennanp ANTENNA_1566 (.A(net3728));
 sg13g2_antennanp ANTENNA_1567 (.A(net3728));
 sg13g2_antennanp ANTENNA_1568 (.A(net3728));
 sg13g2_antennanp ANTENNA_1569 (.A(net3728));
 sg13g2_antennanp ANTENNA_1570 (.A(net3728));
 sg13g2_antennanp ANTENNA_1571 (.A(net3728));
 sg13g2_antennanp ANTENNA_1572 (.A(net4136));
 sg13g2_antennanp ANTENNA_1573 (.A(net4136));
 sg13g2_antennanp ANTENNA_1574 (.A(net4136));
 sg13g2_antennanp ANTENNA_1575 (.A(net4136));
 sg13g2_antennanp ANTENNA_1576 (.A(net4136));
 sg13g2_antennanp ANTENNA_1577 (.A(net4709));
 sg13g2_antennanp ANTENNA_1578 (.A(net4709));
 sg13g2_antennanp ANTENNA_1579 (.A(net4709));
 sg13g2_antennanp ANTENNA_1580 (.A(net4709));
 sg13g2_antennanp ANTENNA_1581 (.A(net4709));
 sg13g2_antennanp ANTENNA_1582 (.A(net4709));
 sg13g2_antennanp ANTENNA_1583 (.A(net4709));
 sg13g2_antennanp ANTENNA_1584 (.A(net4709));
 sg13g2_antennanp ANTENNA_1585 (.A(net4709));
 sg13g2_antennanp ANTENNA_1586 (.A(net4709));
 sg13g2_antennanp ANTENNA_1587 (.A(net4709));
 sg13g2_antennanp ANTENNA_1588 (.A(net4709));
 sg13g2_antennanp ANTENNA_1589 (.A(net4709));
 sg13g2_antennanp ANTENNA_1590 (.A(net2));
 sg13g2_antennanp ANTENNA_1591 (.A(net4));
 sg13g2_antennanp ANTENNA_1592 (.A(net6));
 sg13g2_antennanp ANTENNA_1593 (.A(net7));
 sg13g2_antennanp ANTENNA_1594 (.A(net8));
 sg13g2_antennanp ANTENNA_1595 (.A(net9));
 sg13g2_antennanp ANTENNA_1596 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_1597 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_1598 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_1599 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_1600 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_1601 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_1602 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_1603 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_1604 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_1605 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_1606 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_1607 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_1608 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_1609 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_1610 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_1611 (.A(clknet_0_clk));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_fill_2 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_188 ();
 sg13g2_decap_8 FILLER_0_199 ();
 sg13g2_decap_8 FILLER_0_206 ();
 sg13g2_decap_8 FILLER_0_213 ();
 sg13g2_decap_8 FILLER_0_220 ();
 sg13g2_decap_8 FILLER_0_227 ();
 sg13g2_decap_8 FILLER_0_234 ();
 sg13g2_decap_8 FILLER_0_241 ();
 sg13g2_decap_8 FILLER_0_248 ();
 sg13g2_decap_8 FILLER_0_255 ();
 sg13g2_decap_8 FILLER_0_262 ();
 sg13g2_fill_2 FILLER_0_269 ();
 sg13g2_decap_8 FILLER_0_275 ();
 sg13g2_decap_8 FILLER_0_282 ();
 sg13g2_decap_8 FILLER_0_289 ();
 sg13g2_decap_8 FILLER_0_296 ();
 sg13g2_decap_8 FILLER_0_303 ();
 sg13g2_decap_8 FILLER_0_310 ();
 sg13g2_decap_8 FILLER_0_317 ();
 sg13g2_decap_8 FILLER_0_324 ();
 sg13g2_decap_8 FILLER_0_331 ();
 sg13g2_decap_8 FILLER_0_338 ();
 sg13g2_decap_8 FILLER_0_345 ();
 sg13g2_decap_8 FILLER_0_352 ();
 sg13g2_decap_8 FILLER_0_359 ();
 sg13g2_fill_2 FILLER_0_366 ();
 sg13g2_fill_1 FILLER_0_368 ();
 sg13g2_decap_8 FILLER_0_379 ();
 sg13g2_decap_8 FILLER_0_386 ();
 sg13g2_decap_8 FILLER_0_393 ();
 sg13g2_decap_8 FILLER_0_400 ();
 sg13g2_decap_8 FILLER_0_407 ();
 sg13g2_decap_8 FILLER_0_414 ();
 sg13g2_decap_8 FILLER_0_421 ();
 sg13g2_decap_8 FILLER_0_428 ();
 sg13g2_decap_8 FILLER_0_435 ();
 sg13g2_decap_8 FILLER_0_442 ();
 sg13g2_decap_8 FILLER_0_449 ();
 sg13g2_decap_8 FILLER_0_456 ();
 sg13g2_decap_8 FILLER_0_463 ();
 sg13g2_decap_8 FILLER_0_470 ();
 sg13g2_fill_1 FILLER_0_477 ();
 sg13g2_decap_8 FILLER_0_488 ();
 sg13g2_decap_8 FILLER_0_495 ();
 sg13g2_decap_8 FILLER_0_502 ();
 sg13g2_decap_8 FILLER_0_509 ();
 sg13g2_decap_8 FILLER_0_516 ();
 sg13g2_decap_8 FILLER_0_523 ();
 sg13g2_decap_8 FILLER_0_530 ();
 sg13g2_decap_8 FILLER_0_537 ();
 sg13g2_decap_8 FILLER_0_544 ();
 sg13g2_decap_8 FILLER_0_551 ();
 sg13g2_decap_8 FILLER_0_558 ();
 sg13g2_decap_8 FILLER_0_565 ();
 sg13g2_decap_8 FILLER_0_572 ();
 sg13g2_decap_8 FILLER_0_579 ();
 sg13g2_decap_8 FILLER_0_586 ();
 sg13g2_decap_8 FILLER_0_593 ();
 sg13g2_decap_8 FILLER_0_600 ();
 sg13g2_decap_8 FILLER_0_607 ();
 sg13g2_decap_8 FILLER_0_614 ();
 sg13g2_decap_8 FILLER_0_621 ();
 sg13g2_decap_8 FILLER_0_628 ();
 sg13g2_decap_8 FILLER_0_635 ();
 sg13g2_decap_8 FILLER_0_642 ();
 sg13g2_decap_8 FILLER_0_649 ();
 sg13g2_decap_8 FILLER_0_656 ();
 sg13g2_decap_8 FILLER_0_663 ();
 sg13g2_decap_8 FILLER_0_670 ();
 sg13g2_decap_8 FILLER_0_677 ();
 sg13g2_decap_8 FILLER_0_684 ();
 sg13g2_decap_8 FILLER_0_691 ();
 sg13g2_decap_8 FILLER_0_698 ();
 sg13g2_decap_8 FILLER_0_705 ();
 sg13g2_fill_2 FILLER_0_712 ();
 sg13g2_decap_8 FILLER_0_719 ();
 sg13g2_decap_8 FILLER_0_726 ();
 sg13g2_decap_8 FILLER_0_733 ();
 sg13g2_decap_8 FILLER_0_740 ();
 sg13g2_decap_8 FILLER_0_747 ();
 sg13g2_fill_2 FILLER_0_754 ();
 sg13g2_fill_1 FILLER_0_756 ();
 sg13g2_decap_8 FILLER_0_767 ();
 sg13g2_decap_4 FILLER_0_774 ();
 sg13g2_decap_8 FILLER_0_788 ();
 sg13g2_decap_8 FILLER_0_795 ();
 sg13g2_decap_8 FILLER_0_802 ();
 sg13g2_decap_8 FILLER_0_809 ();
 sg13g2_decap_8 FILLER_0_816 ();
 sg13g2_decap_8 FILLER_0_823 ();
 sg13g2_decap_4 FILLER_0_830 ();
 sg13g2_fill_1 FILLER_0_834 ();
 sg13g2_decap_8 FILLER_0_845 ();
 sg13g2_decap_8 FILLER_0_852 ();
 sg13g2_decap_8 FILLER_0_859 ();
 sg13g2_decap_8 FILLER_0_866 ();
 sg13g2_decap_8 FILLER_0_873 ();
 sg13g2_decap_8 FILLER_0_880 ();
 sg13g2_decap_8 FILLER_0_887 ();
 sg13g2_decap_8 FILLER_0_894 ();
 sg13g2_decap_8 FILLER_0_901 ();
 sg13g2_fill_2 FILLER_0_908 ();
 sg13g2_decap_8 FILLER_0_936 ();
 sg13g2_decap_8 FILLER_0_943 ();
 sg13g2_decap_8 FILLER_0_950 ();
 sg13g2_decap_8 FILLER_0_957 ();
 sg13g2_decap_8 FILLER_0_964 ();
 sg13g2_decap_8 FILLER_0_971 ();
 sg13g2_decap_8 FILLER_0_978 ();
 sg13g2_decap_8 FILLER_0_985 ();
 sg13g2_decap_8 FILLER_0_992 ();
 sg13g2_decap_8 FILLER_0_999 ();
 sg13g2_decap_8 FILLER_0_1006 ();
 sg13g2_decap_8 FILLER_0_1013 ();
 sg13g2_decap_8 FILLER_0_1020 ();
 sg13g2_decap_8 FILLER_0_1027 ();
 sg13g2_decap_8 FILLER_0_1034 ();
 sg13g2_decap_8 FILLER_0_1041 ();
 sg13g2_decap_8 FILLER_0_1048 ();
 sg13g2_decap_8 FILLER_0_1055 ();
 sg13g2_decap_8 FILLER_0_1062 ();
 sg13g2_decap_8 FILLER_0_1069 ();
 sg13g2_decap_8 FILLER_0_1076 ();
 sg13g2_decap_8 FILLER_0_1083 ();
 sg13g2_decap_8 FILLER_0_1090 ();
 sg13g2_decap_8 FILLER_0_1097 ();
 sg13g2_decap_8 FILLER_0_1104 ();
 sg13g2_decap_8 FILLER_0_1111 ();
 sg13g2_decap_8 FILLER_0_1118 ();
 sg13g2_fill_1 FILLER_0_1125 ();
 sg13g2_decap_8 FILLER_0_1161 ();
 sg13g2_decap_8 FILLER_0_1168 ();
 sg13g2_decap_8 FILLER_0_1175 ();
 sg13g2_decap_8 FILLER_0_1182 ();
 sg13g2_decap_8 FILLER_0_1189 ();
 sg13g2_decap_8 FILLER_0_1196 ();
 sg13g2_decap_8 FILLER_0_1203 ();
 sg13g2_decap_8 FILLER_0_1210 ();
 sg13g2_decap_8 FILLER_0_1217 ();
 sg13g2_decap_8 FILLER_0_1224 ();
 sg13g2_decap_8 FILLER_0_1231 ();
 sg13g2_decap_8 FILLER_0_1238 ();
 sg13g2_decap_4 FILLER_0_1245 ();
 sg13g2_decap_8 FILLER_0_1254 ();
 sg13g2_decap_8 FILLER_0_1261 ();
 sg13g2_decap_8 FILLER_0_1268 ();
 sg13g2_decap_8 FILLER_0_1275 ();
 sg13g2_decap_8 FILLER_0_1282 ();
 sg13g2_decap_8 FILLER_0_1289 ();
 sg13g2_decap_8 FILLER_0_1296 ();
 sg13g2_decap_4 FILLER_0_1303 ();
 sg13g2_fill_2 FILLER_0_1307 ();
 sg13g2_decap_8 FILLER_0_1314 ();
 sg13g2_decap_8 FILLER_0_1321 ();
 sg13g2_decap_8 FILLER_0_1328 ();
 sg13g2_decap_8 FILLER_0_1335 ();
 sg13g2_decap_8 FILLER_0_1342 ();
 sg13g2_decap_8 FILLER_0_1349 ();
 sg13g2_decap_8 FILLER_0_1382 ();
 sg13g2_decap_8 FILLER_0_1389 ();
 sg13g2_decap_8 FILLER_0_1396 ();
 sg13g2_decap_8 FILLER_0_1403 ();
 sg13g2_decap_8 FILLER_0_1410 ();
 sg13g2_decap_8 FILLER_0_1417 ();
 sg13g2_decap_8 FILLER_0_1424 ();
 sg13g2_decap_8 FILLER_0_1431 ();
 sg13g2_decap_8 FILLER_0_1438 ();
 sg13g2_decap_8 FILLER_0_1445 ();
 sg13g2_decap_8 FILLER_0_1452 ();
 sg13g2_decap_8 FILLER_0_1459 ();
 sg13g2_decap_8 FILLER_0_1466 ();
 sg13g2_decap_8 FILLER_0_1473 ();
 sg13g2_decap_8 FILLER_0_1480 ();
 sg13g2_decap_8 FILLER_0_1487 ();
 sg13g2_decap_8 FILLER_0_1494 ();
 sg13g2_decap_8 FILLER_0_1501 ();
 sg13g2_decap_8 FILLER_0_1508 ();
 sg13g2_decap_8 FILLER_0_1515 ();
 sg13g2_decap_8 FILLER_0_1522 ();
 sg13g2_decap_8 FILLER_0_1529 ();
 sg13g2_decap_8 FILLER_0_1536 ();
 sg13g2_decap_8 FILLER_0_1543 ();
 sg13g2_decap_8 FILLER_0_1550 ();
 sg13g2_decap_8 FILLER_0_1557 ();
 sg13g2_decap_8 FILLER_0_1564 ();
 sg13g2_decap_8 FILLER_0_1571 ();
 sg13g2_fill_1 FILLER_0_1578 ();
 sg13g2_decap_8 FILLER_0_1605 ();
 sg13g2_decap_8 FILLER_0_1612 ();
 sg13g2_decap_8 FILLER_0_1619 ();
 sg13g2_decap_8 FILLER_0_1626 ();
 sg13g2_decap_8 FILLER_0_1633 ();
 sg13g2_decap_8 FILLER_0_1640 ();
 sg13g2_decap_8 FILLER_0_1647 ();
 sg13g2_decap_8 FILLER_0_1654 ();
 sg13g2_decap_8 FILLER_0_1661 ();
 sg13g2_decap_8 FILLER_0_1668 ();
 sg13g2_decap_8 FILLER_0_1675 ();
 sg13g2_fill_1 FILLER_0_1682 ();
 sg13g2_decap_8 FILLER_0_1709 ();
 sg13g2_decap_8 FILLER_0_1716 ();
 sg13g2_decap_8 FILLER_0_1723 ();
 sg13g2_decap_8 FILLER_0_1730 ();
 sg13g2_decap_8 FILLER_0_1737 ();
 sg13g2_decap_8 FILLER_0_1744 ();
 sg13g2_decap_8 FILLER_0_1751 ();
 sg13g2_decap_8 FILLER_0_1758 ();
 sg13g2_decap_8 FILLER_0_1765 ();
 sg13g2_decap_8 FILLER_0_1772 ();
 sg13g2_decap_8 FILLER_0_1779 ();
 sg13g2_decap_8 FILLER_0_1786 ();
 sg13g2_decap_8 FILLER_0_1793 ();
 sg13g2_decap_8 FILLER_0_1800 ();
 sg13g2_decap_8 FILLER_0_1807 ();
 sg13g2_decap_8 FILLER_0_1814 ();
 sg13g2_decap_8 FILLER_0_1821 ();
 sg13g2_decap_8 FILLER_0_1828 ();
 sg13g2_decap_8 FILLER_0_1835 ();
 sg13g2_decap_8 FILLER_0_1842 ();
 sg13g2_fill_1 FILLER_0_1849 ();
 sg13g2_decap_8 FILLER_0_1876 ();
 sg13g2_decap_8 FILLER_0_1883 ();
 sg13g2_decap_8 FILLER_0_1890 ();
 sg13g2_decap_8 FILLER_0_1897 ();
 sg13g2_fill_2 FILLER_0_1904 ();
 sg13g2_decap_8 FILLER_0_1932 ();
 sg13g2_decap_8 FILLER_0_1939 ();
 sg13g2_decap_8 FILLER_0_1946 ();
 sg13g2_decap_8 FILLER_0_1953 ();
 sg13g2_decap_8 FILLER_0_1960 ();
 sg13g2_decap_8 FILLER_0_1967 ();
 sg13g2_decap_8 FILLER_0_1974 ();
 sg13g2_decap_8 FILLER_0_1981 ();
 sg13g2_decap_8 FILLER_0_1988 ();
 sg13g2_decap_8 FILLER_0_1995 ();
 sg13g2_decap_8 FILLER_0_2002 ();
 sg13g2_decap_8 FILLER_0_2009 ();
 sg13g2_decap_8 FILLER_0_2016 ();
 sg13g2_decap_8 FILLER_0_2023 ();
 sg13g2_decap_8 FILLER_0_2030 ();
 sg13g2_decap_8 FILLER_0_2037 ();
 sg13g2_decap_8 FILLER_0_2044 ();
 sg13g2_decap_8 FILLER_0_2051 ();
 sg13g2_decap_8 FILLER_0_2058 ();
 sg13g2_decap_8 FILLER_0_2065 ();
 sg13g2_decap_8 FILLER_0_2072 ();
 sg13g2_decap_8 FILLER_0_2079 ();
 sg13g2_decap_8 FILLER_0_2086 ();
 sg13g2_decap_8 FILLER_0_2093 ();
 sg13g2_decap_8 FILLER_0_2100 ();
 sg13g2_decap_8 FILLER_0_2107 ();
 sg13g2_decap_8 FILLER_0_2114 ();
 sg13g2_decap_8 FILLER_0_2121 ();
 sg13g2_decap_8 FILLER_0_2128 ();
 sg13g2_decap_8 FILLER_0_2135 ();
 sg13g2_decap_8 FILLER_0_2142 ();
 sg13g2_decap_8 FILLER_0_2149 ();
 sg13g2_decap_8 FILLER_0_2156 ();
 sg13g2_decap_8 FILLER_0_2163 ();
 sg13g2_decap_4 FILLER_0_2170 ();
 sg13g2_fill_2 FILLER_0_2174 ();
 sg13g2_decap_8 FILLER_0_2202 ();
 sg13g2_decap_8 FILLER_0_2209 ();
 sg13g2_decap_8 FILLER_0_2216 ();
 sg13g2_decap_8 FILLER_0_2223 ();
 sg13g2_decap_8 FILLER_0_2230 ();
 sg13g2_decap_8 FILLER_0_2237 ();
 sg13g2_decap_8 FILLER_0_2244 ();
 sg13g2_decap_8 FILLER_0_2251 ();
 sg13g2_decap_8 FILLER_0_2258 ();
 sg13g2_decap_8 FILLER_0_2265 ();
 sg13g2_decap_8 FILLER_0_2272 ();
 sg13g2_decap_8 FILLER_0_2279 ();
 sg13g2_decap_8 FILLER_0_2286 ();
 sg13g2_decap_8 FILLER_0_2293 ();
 sg13g2_decap_8 FILLER_0_2300 ();
 sg13g2_decap_8 FILLER_0_2307 ();
 sg13g2_decap_8 FILLER_0_2314 ();
 sg13g2_decap_8 FILLER_0_2321 ();
 sg13g2_decap_8 FILLER_0_2328 ();
 sg13g2_decap_8 FILLER_0_2335 ();
 sg13g2_decap_8 FILLER_0_2342 ();
 sg13g2_decap_8 FILLER_0_2349 ();
 sg13g2_decap_8 FILLER_0_2356 ();
 sg13g2_decap_8 FILLER_0_2363 ();
 sg13g2_decap_8 FILLER_0_2370 ();
 sg13g2_decap_8 FILLER_0_2377 ();
 sg13g2_decap_8 FILLER_0_2384 ();
 sg13g2_decap_8 FILLER_0_2391 ();
 sg13g2_decap_8 FILLER_0_2398 ();
 sg13g2_decap_8 FILLER_0_2405 ();
 sg13g2_decap_8 FILLER_0_2412 ();
 sg13g2_decap_8 FILLER_0_2419 ();
 sg13g2_decap_8 FILLER_0_2426 ();
 sg13g2_decap_8 FILLER_0_2433 ();
 sg13g2_decap_8 FILLER_0_2440 ();
 sg13g2_decap_8 FILLER_0_2447 ();
 sg13g2_decap_8 FILLER_0_2454 ();
 sg13g2_decap_8 FILLER_0_2461 ();
 sg13g2_decap_8 FILLER_0_2468 ();
 sg13g2_decap_8 FILLER_0_2475 ();
 sg13g2_decap_8 FILLER_0_2482 ();
 sg13g2_decap_8 FILLER_0_2489 ();
 sg13g2_decap_8 FILLER_0_2496 ();
 sg13g2_decap_8 FILLER_0_2503 ();
 sg13g2_decap_8 FILLER_0_2510 ();
 sg13g2_decap_8 FILLER_0_2517 ();
 sg13g2_decap_8 FILLER_0_2524 ();
 sg13g2_decap_8 FILLER_0_2531 ();
 sg13g2_decap_8 FILLER_0_2538 ();
 sg13g2_decap_8 FILLER_0_2545 ();
 sg13g2_decap_8 FILLER_0_2552 ();
 sg13g2_decap_8 FILLER_0_2559 ();
 sg13g2_decap_8 FILLER_0_2566 ();
 sg13g2_decap_8 FILLER_0_2573 ();
 sg13g2_decap_8 FILLER_0_2580 ();
 sg13g2_decap_8 FILLER_0_2587 ();
 sg13g2_decap_8 FILLER_0_2594 ();
 sg13g2_decap_8 FILLER_0_2601 ();
 sg13g2_decap_8 FILLER_0_2608 ();
 sg13g2_decap_8 FILLER_0_2615 ();
 sg13g2_decap_8 FILLER_0_2622 ();
 sg13g2_decap_8 FILLER_0_2629 ();
 sg13g2_decap_8 FILLER_0_2636 ();
 sg13g2_decap_8 FILLER_0_2643 ();
 sg13g2_decap_8 FILLER_0_2650 ();
 sg13g2_decap_8 FILLER_0_2657 ();
 sg13g2_decap_8 FILLER_0_2664 ();
 sg13g2_decap_8 FILLER_0_2671 ();
 sg13g2_decap_8 FILLER_0_2678 ();
 sg13g2_decap_8 FILLER_0_2685 ();
 sg13g2_decap_8 FILLER_0_2692 ();
 sg13g2_decap_8 FILLER_0_2699 ();
 sg13g2_decap_8 FILLER_0_2706 ();
 sg13g2_decap_8 FILLER_0_2713 ();
 sg13g2_decap_8 FILLER_0_2720 ();
 sg13g2_decap_8 FILLER_0_2727 ();
 sg13g2_decap_8 FILLER_0_2734 ();
 sg13g2_decap_8 FILLER_0_2741 ();
 sg13g2_decap_8 FILLER_0_2748 ();
 sg13g2_decap_8 FILLER_0_2755 ();
 sg13g2_decap_8 FILLER_0_2762 ();
 sg13g2_decap_8 FILLER_0_2769 ();
 sg13g2_decap_8 FILLER_0_2776 ();
 sg13g2_decap_8 FILLER_0_2783 ();
 sg13g2_decap_8 FILLER_0_2790 ();
 sg13g2_decap_8 FILLER_0_2797 ();
 sg13g2_decap_8 FILLER_0_2804 ();
 sg13g2_decap_8 FILLER_0_2811 ();
 sg13g2_decap_8 FILLER_0_2818 ();
 sg13g2_decap_8 FILLER_0_2825 ();
 sg13g2_decap_8 FILLER_0_2832 ();
 sg13g2_decap_8 FILLER_0_2839 ();
 sg13g2_decap_8 FILLER_0_2846 ();
 sg13g2_decap_8 FILLER_0_2853 ();
 sg13g2_decap_8 FILLER_0_2860 ();
 sg13g2_decap_8 FILLER_0_2867 ();
 sg13g2_decap_8 FILLER_0_2874 ();
 sg13g2_decap_8 FILLER_0_2881 ();
 sg13g2_decap_8 FILLER_0_2888 ();
 sg13g2_decap_8 FILLER_0_2895 ();
 sg13g2_decap_8 FILLER_0_2902 ();
 sg13g2_decap_8 FILLER_0_2909 ();
 sg13g2_decap_8 FILLER_0_2916 ();
 sg13g2_decap_8 FILLER_0_2923 ();
 sg13g2_decap_8 FILLER_0_2930 ();
 sg13g2_decap_8 FILLER_0_2937 ();
 sg13g2_decap_8 FILLER_0_2944 ();
 sg13g2_decap_8 FILLER_0_2951 ();
 sg13g2_decap_8 FILLER_0_2958 ();
 sg13g2_decap_8 FILLER_0_2965 ();
 sg13g2_decap_8 FILLER_0_2972 ();
 sg13g2_decap_8 FILLER_0_2979 ();
 sg13g2_decap_8 FILLER_0_2986 ();
 sg13g2_decap_8 FILLER_0_2993 ();
 sg13g2_decap_8 FILLER_0_3000 ();
 sg13g2_decap_8 FILLER_0_3007 ();
 sg13g2_decap_8 FILLER_0_3014 ();
 sg13g2_decap_8 FILLER_0_3021 ();
 sg13g2_decap_8 FILLER_0_3028 ();
 sg13g2_decap_8 FILLER_0_3035 ();
 sg13g2_decap_8 FILLER_0_3042 ();
 sg13g2_decap_8 FILLER_0_3049 ();
 sg13g2_decap_8 FILLER_0_3056 ();
 sg13g2_decap_8 FILLER_0_3063 ();
 sg13g2_decap_8 FILLER_0_3070 ();
 sg13g2_decap_8 FILLER_0_3077 ();
 sg13g2_decap_8 FILLER_0_3084 ();
 sg13g2_decap_8 FILLER_0_3091 ();
 sg13g2_decap_8 FILLER_0_3098 ();
 sg13g2_decap_8 FILLER_0_3105 ();
 sg13g2_decap_8 FILLER_0_3112 ();
 sg13g2_decap_8 FILLER_0_3119 ();
 sg13g2_decap_8 FILLER_0_3126 ();
 sg13g2_decap_8 FILLER_0_3133 ();
 sg13g2_decap_8 FILLER_0_3140 ();
 sg13g2_decap_8 FILLER_0_3147 ();
 sg13g2_decap_8 FILLER_0_3154 ();
 sg13g2_decap_8 FILLER_0_3161 ();
 sg13g2_decap_4 FILLER_0_3168 ();
 sg13g2_fill_1 FILLER_0_3172 ();
 sg13g2_decap_8 FILLER_0_3181 ();
 sg13g2_decap_8 FILLER_0_3188 ();
 sg13g2_decap_8 FILLER_0_3195 ();
 sg13g2_decap_8 FILLER_0_3202 ();
 sg13g2_decap_8 FILLER_0_3209 ();
 sg13g2_decap_8 FILLER_0_3224 ();
 sg13g2_decap_8 FILLER_0_3231 ();
 sg13g2_decap_8 FILLER_0_3238 ();
 sg13g2_decap_8 FILLER_0_3245 ();
 sg13g2_decap_8 FILLER_0_3252 ();
 sg13g2_decap_8 FILLER_0_3259 ();
 sg13g2_decap_8 FILLER_0_3266 ();
 sg13g2_decap_8 FILLER_0_3273 ();
 sg13g2_decap_8 FILLER_0_3280 ();
 sg13g2_decap_8 FILLER_0_3287 ();
 sg13g2_decap_8 FILLER_0_3294 ();
 sg13g2_decap_8 FILLER_0_3301 ();
 sg13g2_decap_8 FILLER_0_3308 ();
 sg13g2_decap_8 FILLER_0_3315 ();
 sg13g2_decap_8 FILLER_0_3322 ();
 sg13g2_decap_8 FILLER_0_3329 ();
 sg13g2_decap_8 FILLER_0_3336 ();
 sg13g2_decap_8 FILLER_0_3343 ();
 sg13g2_decap_8 FILLER_0_3350 ();
 sg13g2_decap_8 FILLER_0_3357 ();
 sg13g2_decap_8 FILLER_0_3364 ();
 sg13g2_decap_8 FILLER_0_3371 ();
 sg13g2_decap_8 FILLER_0_3378 ();
 sg13g2_decap_8 FILLER_0_3385 ();
 sg13g2_decap_8 FILLER_0_3392 ();
 sg13g2_decap_8 FILLER_0_3399 ();
 sg13g2_decap_8 FILLER_0_3406 ();
 sg13g2_decap_8 FILLER_0_3413 ();
 sg13g2_decap_8 FILLER_0_3420 ();
 sg13g2_decap_8 FILLER_0_3427 ();
 sg13g2_decap_8 FILLER_0_3434 ();
 sg13g2_decap_8 FILLER_0_3441 ();
 sg13g2_decap_8 FILLER_0_3448 ();
 sg13g2_decap_8 FILLER_0_3455 ();
 sg13g2_decap_8 FILLER_0_3462 ();
 sg13g2_decap_8 FILLER_0_3469 ();
 sg13g2_decap_8 FILLER_0_3476 ();
 sg13g2_decap_8 FILLER_0_3483 ();
 sg13g2_decap_8 FILLER_0_3490 ();
 sg13g2_decap_8 FILLER_0_3497 ();
 sg13g2_decap_8 FILLER_0_3504 ();
 sg13g2_decap_8 FILLER_0_3511 ();
 sg13g2_decap_8 FILLER_0_3518 ();
 sg13g2_decap_8 FILLER_0_3525 ();
 sg13g2_decap_8 FILLER_0_3532 ();
 sg13g2_decap_8 FILLER_0_3539 ();
 sg13g2_decap_8 FILLER_0_3546 ();
 sg13g2_decap_8 FILLER_0_3553 ();
 sg13g2_decap_8 FILLER_0_3560 ();
 sg13g2_decap_8 FILLER_0_3567 ();
 sg13g2_decap_4 FILLER_0_3574 ();
 sg13g2_fill_2 FILLER_0_3578 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_4 FILLER_1_63 ();
 sg13g2_fill_2 FILLER_1_67 ();
 sg13g2_decap_8 FILLER_1_95 ();
 sg13g2_decap_8 FILLER_1_102 ();
 sg13g2_decap_8 FILLER_1_109 ();
 sg13g2_decap_8 FILLER_1_116 ();
 sg13g2_decap_8 FILLER_1_123 ();
 sg13g2_decap_8 FILLER_1_130 ();
 sg13g2_decap_8 FILLER_1_137 ();
 sg13g2_decap_8 FILLER_1_144 ();
 sg13g2_decap_8 FILLER_1_151 ();
 sg13g2_decap_8 FILLER_1_158 ();
 sg13g2_decap_8 FILLER_1_165 ();
 sg13g2_decap_8 FILLER_1_172 ();
 sg13g2_fill_1 FILLER_1_179 ();
 sg13g2_fill_2 FILLER_1_185 ();
 sg13g2_fill_1 FILLER_1_187 ();
 sg13g2_decap_8 FILLER_1_223 ();
 sg13g2_decap_8 FILLER_1_230 ();
 sg13g2_decap_8 FILLER_1_237 ();
 sg13g2_decap_4 FILLER_1_244 ();
 sg13g2_fill_2 FILLER_1_248 ();
 sg13g2_decap_8 FILLER_1_281 ();
 sg13g2_fill_1 FILLER_1_288 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_4 FILLER_1_362 ();
 sg13g2_fill_1 FILLER_1_366 ();
 sg13g2_decap_8 FILLER_1_393 ();
 sg13g2_fill_2 FILLER_1_400 ();
 sg13g2_fill_2 FILLER_1_438 ();
 sg13g2_fill_1 FILLER_1_440 ();
 sg13g2_decap_4 FILLER_1_477 ();
 sg13g2_fill_2 FILLER_1_481 ();
 sg13g2_decap_8 FILLER_1_509 ();
 sg13g2_decap_8 FILLER_1_516 ();
 sg13g2_decap_8 FILLER_1_531 ();
 sg13g2_decap_8 FILLER_1_538 ();
 sg13g2_decap_8 FILLER_1_545 ();
 sg13g2_decap_8 FILLER_1_552 ();
 sg13g2_fill_2 FILLER_1_559 ();
 sg13g2_decap_8 FILLER_1_587 ();
 sg13g2_fill_1 FILLER_1_594 ();
 sg13g2_decap_8 FILLER_1_621 ();
 sg13g2_decap_8 FILLER_1_628 ();
 sg13g2_decap_8 FILLER_1_635 ();
 sg13g2_decap_8 FILLER_1_642 ();
 sg13g2_fill_1 FILLER_1_649 ();
 sg13g2_decap_4 FILLER_1_660 ();
 sg13g2_fill_2 FILLER_1_664 ();
 sg13g2_decap_8 FILLER_1_675 ();
 sg13g2_decap_8 FILLER_1_682 ();
 sg13g2_decap_8 FILLER_1_689 ();
 sg13g2_decap_4 FILLER_1_696 ();
 sg13g2_fill_1 FILLER_1_700 ();
 sg13g2_decap_8 FILLER_1_727 ();
 sg13g2_decap_8 FILLER_1_734 ();
 sg13g2_decap_8 FILLER_1_741 ();
 sg13g2_decap_8 FILLER_1_748 ();
 sg13g2_fill_2 FILLER_1_755 ();
 sg13g2_decap_8 FILLER_1_786 ();
 sg13g2_decap_8 FILLER_1_793 ();
 sg13g2_decap_8 FILLER_1_800 ();
 sg13g2_decap_8 FILLER_1_807 ();
 sg13g2_decap_8 FILLER_1_814 ();
 sg13g2_decap_8 FILLER_1_821 ();
 sg13g2_decap_4 FILLER_1_828 ();
 sg13g2_fill_1 FILLER_1_832 ();
 sg13g2_decap_8 FILLER_1_859 ();
 sg13g2_decap_8 FILLER_1_866 ();
 sg13g2_fill_2 FILLER_1_873 ();
 sg13g2_decap_8 FILLER_1_901 ();
 sg13g2_decap_8 FILLER_1_908 ();
 sg13g2_decap_4 FILLER_1_915 ();
 sg13g2_decap_8 FILLER_1_945 ();
 sg13g2_decap_8 FILLER_1_952 ();
 sg13g2_decap_4 FILLER_1_959 ();
 sg13g2_fill_2 FILLER_1_971 ();
 sg13g2_fill_2 FILLER_1_999 ();
 sg13g2_decap_8 FILLER_1_1053 ();
 sg13g2_decap_8 FILLER_1_1060 ();
 sg13g2_decap_8 FILLER_1_1067 ();
 sg13g2_fill_2 FILLER_1_1074 ();
 sg13g2_fill_1 FILLER_1_1076 ();
 sg13g2_decap_8 FILLER_1_1103 ();
 sg13g2_decap_8 FILLER_1_1110 ();
 sg13g2_decap_8 FILLER_1_1117 ();
 sg13g2_fill_2 FILLER_1_1124 ();
 sg13g2_fill_1 FILLER_1_1126 ();
 sg13g2_decap_8 FILLER_1_1157 ();
 sg13g2_decap_8 FILLER_1_1164 ();
 sg13g2_decap_8 FILLER_1_1171 ();
 sg13g2_fill_2 FILLER_1_1178 ();
 sg13g2_fill_1 FILLER_1_1180 ();
 sg13g2_fill_1 FILLER_1_1189 ();
 sg13g2_decap_8 FILLER_1_1216 ();
 sg13g2_decap_8 FILLER_1_1223 ();
 sg13g2_decap_4 FILLER_1_1230 ();
 sg13g2_fill_2 FILLER_1_1234 ();
 sg13g2_decap_8 FILLER_1_1261 ();
 sg13g2_decap_8 FILLER_1_1268 ();
 sg13g2_fill_2 FILLER_1_1275 ();
 sg13g2_fill_1 FILLER_1_1277 ();
 sg13g2_decap_8 FILLER_1_1288 ();
 sg13g2_decap_8 FILLER_1_1295 ();
 sg13g2_decap_8 FILLER_1_1325 ();
 sg13g2_decap_8 FILLER_1_1332 ();
 sg13g2_decap_8 FILLER_1_1339 ();
 sg13g2_decap_8 FILLER_1_1356 ();
 sg13g2_decap_8 FILLER_1_1389 ();
 sg13g2_decap_8 FILLER_1_1396 ();
 sg13g2_decap_8 FILLER_1_1403 ();
 sg13g2_decap_8 FILLER_1_1410 ();
 sg13g2_decap_8 FILLER_1_1417 ();
 sg13g2_decap_8 FILLER_1_1424 ();
 sg13g2_decap_8 FILLER_1_1431 ();
 sg13g2_decap_8 FILLER_1_1438 ();
 sg13g2_decap_8 FILLER_1_1445 ();
 sg13g2_decap_8 FILLER_1_1452 ();
 sg13g2_decap_8 FILLER_1_1459 ();
 sg13g2_decap_4 FILLER_1_1466 ();
 sg13g2_fill_1 FILLER_1_1470 ();
 sg13g2_decap_8 FILLER_1_1497 ();
 sg13g2_decap_8 FILLER_1_1504 ();
 sg13g2_decap_8 FILLER_1_1511 ();
 sg13g2_decap_4 FILLER_1_1518 ();
 sg13g2_fill_2 FILLER_1_1522 ();
 sg13g2_decap_8 FILLER_1_1550 ();
 sg13g2_decap_8 FILLER_1_1557 ();
 sg13g2_decap_8 FILLER_1_1564 ();
 sg13g2_fill_2 FILLER_1_1571 ();
 sg13g2_fill_1 FILLER_1_1573 ();
 sg13g2_decap_8 FILLER_1_1609 ();
 sg13g2_decap_8 FILLER_1_1616 ();
 sg13g2_decap_4 FILLER_1_1623 ();
 sg13g2_fill_2 FILLER_1_1627 ();
 sg13g2_decap_8 FILLER_1_1655 ();
 sg13g2_decap_8 FILLER_1_1662 ();
 sg13g2_decap_8 FILLER_1_1669 ();
 sg13g2_decap_8 FILLER_1_1676 ();
 sg13g2_decap_4 FILLER_1_1683 ();
 sg13g2_decap_8 FILLER_1_1716 ();
 sg13g2_decap_8 FILLER_1_1723 ();
 sg13g2_decap_8 FILLER_1_1730 ();
 sg13g2_fill_1 FILLER_1_1737 ();
 sg13g2_fill_2 FILLER_1_1781 ();
 sg13g2_fill_1 FILLER_1_1783 ();
 sg13g2_decap_8 FILLER_1_1792 ();
 sg13g2_fill_1 FILLER_1_1799 ();
 sg13g2_decap_8 FILLER_1_1826 ();
 sg13g2_decap_8 FILLER_1_1833 ();
 sg13g2_decap_4 FILLER_1_1840 ();
 sg13g2_decap_8 FILLER_1_1882 ();
 sg13g2_decap_8 FILLER_1_1889 ();
 sg13g2_decap_4 FILLER_1_1922 ();
 sg13g2_decap_8 FILLER_1_1935 ();
 sg13g2_decap_8 FILLER_1_1942 ();
 sg13g2_decap_8 FILLER_1_1949 ();
 sg13g2_decap_8 FILLER_1_1956 ();
 sg13g2_decap_8 FILLER_1_1963 ();
 sg13g2_decap_8 FILLER_1_1996 ();
 sg13g2_decap_8 FILLER_1_2003 ();
 sg13g2_decap_4 FILLER_1_2010 ();
 sg13g2_fill_1 FILLER_1_2014 ();
 sg13g2_decap_8 FILLER_1_2023 ();
 sg13g2_decap_8 FILLER_1_2030 ();
 sg13g2_fill_2 FILLER_1_2037 ();
 sg13g2_decap_8 FILLER_1_2047 ();
 sg13g2_decap_8 FILLER_1_2054 ();
 sg13g2_decap_4 FILLER_1_2061 ();
 sg13g2_decap_8 FILLER_1_2097 ();
 sg13g2_fill_2 FILLER_1_2104 ();
 sg13g2_fill_1 FILLER_1_2106 ();
 sg13g2_decap_8 FILLER_1_2133 ();
 sg13g2_decap_8 FILLER_1_2140 ();
 sg13g2_decap_8 FILLER_1_2147 ();
 sg13g2_decap_8 FILLER_1_2154 ();
 sg13g2_decap_4 FILLER_1_2161 ();
 sg13g2_decap_8 FILLER_1_2191 ();
 sg13g2_decap_8 FILLER_1_2198 ();
 sg13g2_decap_8 FILLER_1_2205 ();
 sg13g2_decap_8 FILLER_1_2212 ();
 sg13g2_decap_8 FILLER_1_2219 ();
 sg13g2_decap_4 FILLER_1_2226 ();
 sg13g2_fill_2 FILLER_1_2230 ();
 sg13g2_fill_2 FILLER_1_2258 ();
 sg13g2_decap_8 FILLER_1_2286 ();
 sg13g2_decap_8 FILLER_1_2293 ();
 sg13g2_decap_8 FILLER_1_2300 ();
 sg13g2_decap_8 FILLER_1_2307 ();
 sg13g2_decap_8 FILLER_1_2314 ();
 sg13g2_fill_1 FILLER_1_2321 ();
 sg13g2_fill_1 FILLER_1_2332 ();
 sg13g2_decap_8 FILLER_1_2359 ();
 sg13g2_decap_8 FILLER_1_2366 ();
 sg13g2_decap_8 FILLER_1_2373 ();
 sg13g2_decap_8 FILLER_1_2380 ();
 sg13g2_decap_8 FILLER_1_2387 ();
 sg13g2_fill_1 FILLER_1_2394 ();
 sg13g2_decap_8 FILLER_1_2405 ();
 sg13g2_decap_8 FILLER_1_2438 ();
 sg13g2_decap_8 FILLER_1_2445 ();
 sg13g2_decap_4 FILLER_1_2452 ();
 sg13g2_fill_2 FILLER_1_2456 ();
 sg13g2_decap_8 FILLER_1_2484 ();
 sg13g2_decap_8 FILLER_1_2491 ();
 sg13g2_decap_8 FILLER_1_2498 ();
 sg13g2_decap_8 FILLER_1_2505 ();
 sg13g2_decap_4 FILLER_1_2512 ();
 sg13g2_decap_8 FILLER_1_2529 ();
 sg13g2_decap_8 FILLER_1_2536 ();
 sg13g2_decap_8 FILLER_1_2543 ();
 sg13g2_decap_4 FILLER_1_2560 ();
 sg13g2_decap_8 FILLER_1_2590 ();
 sg13g2_decap_8 FILLER_1_2597 ();
 sg13g2_decap_8 FILLER_1_2604 ();
 sg13g2_decap_4 FILLER_1_2611 ();
 sg13g2_fill_2 FILLER_1_2615 ();
 sg13g2_decap_8 FILLER_1_2632 ();
 sg13g2_decap_8 FILLER_1_2639 ();
 sg13g2_decap_8 FILLER_1_2646 ();
 sg13g2_decap_8 FILLER_1_2653 ();
 sg13g2_fill_2 FILLER_1_2660 ();
 sg13g2_fill_1 FILLER_1_2662 ();
 sg13g2_decap_8 FILLER_1_2689 ();
 sg13g2_decap_8 FILLER_1_2696 ();
 sg13g2_decap_8 FILLER_1_2703 ();
 sg13g2_decap_8 FILLER_1_2710 ();
 sg13g2_decap_8 FILLER_1_2717 ();
 sg13g2_decap_8 FILLER_1_2724 ();
 sg13g2_decap_4 FILLER_1_2731 ();
 sg13g2_fill_1 FILLER_1_2735 ();
 sg13g2_decap_8 FILLER_1_2762 ();
 sg13g2_decap_8 FILLER_1_2769 ();
 sg13g2_decap_4 FILLER_1_2776 ();
 sg13g2_fill_2 FILLER_1_2806 ();
 sg13g2_fill_1 FILLER_1_2813 ();
 sg13g2_decap_8 FILLER_1_2819 ();
 sg13g2_fill_2 FILLER_1_2826 ();
 sg13g2_fill_1 FILLER_1_2828 ();
 sg13g2_decap_8 FILLER_1_2858 ();
 sg13g2_decap_4 FILLER_1_2865 ();
 sg13g2_decap_8 FILLER_1_2877 ();
 sg13g2_decap_4 FILLER_1_2884 ();
 sg13g2_fill_1 FILLER_1_2888 ();
 sg13g2_decap_8 FILLER_1_2915 ();
 sg13g2_decap_8 FILLER_1_2922 ();
 sg13g2_decap_8 FILLER_1_2929 ();
 sg13g2_fill_1 FILLER_1_2936 ();
 sg13g2_decap_8 FILLER_1_2945 ();
 sg13g2_decap_8 FILLER_1_2952 ();
 sg13g2_decap_8 FILLER_1_2959 ();
 sg13g2_decap_8 FILLER_1_2966 ();
 sg13g2_decap_8 FILLER_1_2973 ();
 sg13g2_fill_2 FILLER_1_2980 ();
 sg13g2_fill_1 FILLER_1_3008 ();
 sg13g2_decap_8 FILLER_1_3012 ();
 sg13g2_decap_8 FILLER_1_3071 ();
 sg13g2_decap_8 FILLER_1_3078 ();
 sg13g2_decap_4 FILLER_1_3085 ();
 sg13g2_decap_8 FILLER_1_3118 ();
 sg13g2_decap_8 FILLER_1_3125 ();
 sg13g2_decap_8 FILLER_1_3132 ();
 sg13g2_decap_8 FILLER_1_3191 ();
 sg13g2_decap_4 FILLER_1_3198 ();
 sg13g2_fill_1 FILLER_1_3202 ();
 sg13g2_decap_8 FILLER_1_3242 ();
 sg13g2_decap_8 FILLER_1_3249 ();
 sg13g2_decap_8 FILLER_1_3256 ();
 sg13g2_decap_8 FILLER_1_3263 ();
 sg13g2_decap_8 FILLER_1_3270 ();
 sg13g2_decap_8 FILLER_1_3277 ();
 sg13g2_decap_8 FILLER_1_3284 ();
 sg13g2_decap_8 FILLER_1_3291 ();
 sg13g2_decap_8 FILLER_1_3298 ();
 sg13g2_decap_8 FILLER_1_3305 ();
 sg13g2_decap_8 FILLER_1_3312 ();
 sg13g2_decap_8 FILLER_1_3319 ();
 sg13g2_decap_8 FILLER_1_3326 ();
 sg13g2_decap_8 FILLER_1_3333 ();
 sg13g2_decap_8 FILLER_1_3340 ();
 sg13g2_decap_8 FILLER_1_3347 ();
 sg13g2_decap_8 FILLER_1_3354 ();
 sg13g2_decap_8 FILLER_1_3361 ();
 sg13g2_decap_8 FILLER_1_3368 ();
 sg13g2_decap_8 FILLER_1_3375 ();
 sg13g2_decap_8 FILLER_1_3382 ();
 sg13g2_decap_8 FILLER_1_3389 ();
 sg13g2_decap_8 FILLER_1_3396 ();
 sg13g2_decap_8 FILLER_1_3403 ();
 sg13g2_decap_8 FILLER_1_3410 ();
 sg13g2_decap_8 FILLER_1_3417 ();
 sg13g2_decap_8 FILLER_1_3424 ();
 sg13g2_decap_8 FILLER_1_3431 ();
 sg13g2_decap_8 FILLER_1_3438 ();
 sg13g2_decap_8 FILLER_1_3445 ();
 sg13g2_decap_8 FILLER_1_3452 ();
 sg13g2_decap_8 FILLER_1_3459 ();
 sg13g2_decap_8 FILLER_1_3466 ();
 sg13g2_decap_8 FILLER_1_3473 ();
 sg13g2_decap_8 FILLER_1_3480 ();
 sg13g2_decap_8 FILLER_1_3487 ();
 sg13g2_decap_8 FILLER_1_3494 ();
 sg13g2_decap_8 FILLER_1_3501 ();
 sg13g2_decap_8 FILLER_1_3508 ();
 sg13g2_decap_8 FILLER_1_3515 ();
 sg13g2_decap_8 FILLER_1_3522 ();
 sg13g2_decap_8 FILLER_1_3529 ();
 sg13g2_decap_8 FILLER_1_3536 ();
 sg13g2_decap_8 FILLER_1_3543 ();
 sg13g2_decap_8 FILLER_1_3550 ();
 sg13g2_decap_8 FILLER_1_3557 ();
 sg13g2_decap_8 FILLER_1_3564 ();
 sg13g2_decap_8 FILLER_1_3571 ();
 sg13g2_fill_2 FILLER_1_3578 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_fill_1 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_97 ();
 sg13g2_decap_8 FILLER_2_104 ();
 sg13g2_decap_8 FILLER_2_111 ();
 sg13g2_decap_8 FILLER_2_118 ();
 sg13g2_decap_8 FILLER_2_125 ();
 sg13g2_decap_8 FILLER_2_132 ();
 sg13g2_decap_8 FILLER_2_139 ();
 sg13g2_decap_8 FILLER_2_146 ();
 sg13g2_decap_8 FILLER_2_153 ();
 sg13g2_decap_8 FILLER_2_160 ();
 sg13g2_fill_1 FILLER_2_167 ();
 sg13g2_decap_8 FILLER_2_225 ();
 sg13g2_decap_8 FILLER_2_232 ();
 sg13g2_decap_8 FILLER_2_239 ();
 sg13g2_decap_8 FILLER_2_246 ();
 sg13g2_fill_2 FILLER_2_253 ();
 sg13g2_fill_1 FILLER_2_255 ();
 sg13g2_fill_2 FILLER_2_261 ();
 sg13g2_fill_2 FILLER_2_271 ();
 sg13g2_fill_1 FILLER_2_273 ();
 sg13g2_fill_1 FILLER_2_283 ();
 sg13g2_fill_1 FILLER_2_302 ();
 sg13g2_decap_8 FILLER_2_312 ();
 sg13g2_decap_8 FILLER_2_319 ();
 sg13g2_decap_8 FILLER_2_326 ();
 sg13g2_fill_2 FILLER_2_333 ();
 sg13g2_decap_8 FILLER_2_361 ();
 sg13g2_decap_8 FILLER_2_368 ();
 sg13g2_decap_8 FILLER_2_375 ();
 sg13g2_decap_8 FILLER_2_382 ();
 sg13g2_decap_8 FILLER_2_389 ();
 sg13g2_decap_4 FILLER_2_396 ();
 sg13g2_fill_1 FILLER_2_400 ();
 sg13g2_decap_4 FILLER_2_411 ();
 sg13g2_fill_1 FILLER_2_415 ();
 sg13g2_decap_8 FILLER_2_426 ();
 sg13g2_decap_8 FILLER_2_433 ();
 sg13g2_decap_8 FILLER_2_440 ();
 sg13g2_decap_4 FILLER_2_447 ();
 sg13g2_decap_8 FILLER_2_461 ();
 sg13g2_decap_4 FILLER_2_468 ();
 sg13g2_fill_2 FILLER_2_472 ();
 sg13g2_decap_8 FILLER_2_484 ();
 sg13g2_decap_8 FILLER_2_491 ();
 sg13g2_decap_8 FILLER_2_498 ();
 sg13g2_decap_8 FILLER_2_505 ();
 sg13g2_fill_2 FILLER_2_512 ();
 sg13g2_decap_8 FILLER_2_548 ();
 sg13g2_fill_2 FILLER_2_555 ();
 sg13g2_fill_1 FILLER_2_557 ();
 sg13g2_decap_4 FILLER_2_584 ();
 sg13g2_fill_2 FILLER_2_588 ();
 sg13g2_fill_1 FILLER_2_626 ();
 sg13g2_decap_8 FILLER_2_679 ();
 sg13g2_decap_8 FILLER_2_686 ();
 sg13g2_decap_4 FILLER_2_745 ();
 sg13g2_decap_8 FILLER_2_795 ();
 sg13g2_decap_8 FILLER_2_802 ();
 sg13g2_decap_8 FILLER_2_809 ();
 sg13g2_fill_2 FILLER_2_816 ();
 sg13g2_fill_1 FILLER_2_818 ();
 sg13g2_decap_8 FILLER_2_855 ();
 sg13g2_decap_8 FILLER_2_862 ();
 sg13g2_decap_8 FILLER_2_869 ();
 sg13g2_decap_8 FILLER_2_886 ();
 sg13g2_decap_8 FILLER_2_893 ();
 sg13g2_fill_1 FILLER_2_900 ();
 sg13g2_decap_8 FILLER_2_921 ();
 sg13g2_decap_8 FILLER_2_928 ();
 sg13g2_decap_8 FILLER_2_935 ();
 sg13g2_decap_8 FILLER_2_942 ();
 sg13g2_decap_8 FILLER_2_949 ();
 sg13g2_decap_8 FILLER_2_956 ();
 sg13g2_decap_8 FILLER_2_963 ();
 sg13g2_decap_8 FILLER_2_970 ();
 sg13g2_decap_8 FILLER_2_977 ();
 sg13g2_decap_8 FILLER_2_984 ();
 sg13g2_decap_8 FILLER_2_991 ();
 sg13g2_fill_2 FILLER_2_998 ();
 sg13g2_decap_8 FILLER_2_1009 ();
 sg13g2_decap_8 FILLER_2_1016 ();
 sg13g2_decap_4 FILLER_2_1023 ();
 sg13g2_fill_2 FILLER_2_1068 ();
 sg13g2_decap_8 FILLER_2_1106 ();
 sg13g2_decap_8 FILLER_2_1113 ();
 sg13g2_decap_8 FILLER_2_1120 ();
 sg13g2_decap_8 FILLER_2_1127 ();
 sg13g2_decap_8 FILLER_2_1134 ();
 sg13g2_fill_2 FILLER_2_1141 ();
 sg13g2_decap_8 FILLER_2_1146 ();
 sg13g2_fill_2 FILLER_2_1153 ();
 sg13g2_fill_1 FILLER_2_1155 ();
 sg13g2_fill_2 FILLER_2_1182 ();
 sg13g2_fill_1 FILLER_2_1184 ();
 sg13g2_decap_8 FILLER_2_1221 ();
 sg13g2_decap_4 FILLER_2_1228 ();
 sg13g2_fill_2 FILLER_2_1232 ();
 sg13g2_decap_8 FILLER_2_1270 ();
 sg13g2_fill_2 FILLER_2_1277 ();
 sg13g2_fill_1 FILLER_2_1279 ();
 sg13g2_decap_8 FILLER_2_1340 ();
 sg13g2_decap_8 FILLER_2_1367 ();
 sg13g2_decap_8 FILLER_2_1374 ();
 sg13g2_decap_8 FILLER_2_1381 ();
 sg13g2_decap_8 FILLER_2_1388 ();
 sg13g2_decap_8 FILLER_2_1395 ();
 sg13g2_decap_4 FILLER_2_1402 ();
 sg13g2_decap_8 FILLER_2_1432 ();
 sg13g2_decap_8 FILLER_2_1439 ();
 sg13g2_decap_8 FILLER_2_1446 ();
 sg13g2_decap_8 FILLER_2_1453 ();
 sg13g2_decap_8 FILLER_2_1460 ();
 sg13g2_decap_4 FILLER_2_1467 ();
 sg13g2_fill_1 FILLER_2_1471 ();
 sg13g2_decap_8 FILLER_2_1498 ();
 sg13g2_decap_4 FILLER_2_1505 ();
 sg13g2_fill_1 FILLER_2_1509 ();
 sg13g2_decap_4 FILLER_2_1520 ();
 sg13g2_decap_8 FILLER_2_1550 ();
 sg13g2_decap_8 FILLER_2_1565 ();
 sg13g2_decap_8 FILLER_2_1572 ();
 sg13g2_decap_4 FILLER_2_1579 ();
 sg13g2_decap_8 FILLER_2_1593 ();
 sg13g2_decap_8 FILLER_2_1600 ();
 sg13g2_decap_8 FILLER_2_1607 ();
 sg13g2_decap_8 FILLER_2_1614 ();
 sg13g2_decap_8 FILLER_2_1621 ();
 sg13g2_decap_8 FILLER_2_1628 ();
 sg13g2_decap_4 FILLER_2_1635 ();
 sg13g2_fill_2 FILLER_2_1639 ();
 sg13g2_decap_8 FILLER_2_1665 ();
 sg13g2_decap_8 FILLER_2_1672 ();
 sg13g2_decap_4 FILLER_2_1679 ();
 sg13g2_fill_1 FILLER_2_1683 ();
 sg13g2_fill_2 FILLER_2_1697 ();
 sg13g2_fill_1 FILLER_2_1699 ();
 sg13g2_fill_1 FILLER_2_1713 ();
 sg13g2_decap_8 FILLER_2_1723 ();
 sg13g2_decap_8 FILLER_2_1730 ();
 sg13g2_decap_8 FILLER_2_1737 ();
 sg13g2_decap_8 FILLER_2_1744 ();
 sg13g2_fill_2 FILLER_2_1751 ();
 sg13g2_fill_1 FILLER_2_1753 ();
 sg13g2_fill_1 FILLER_2_1779 ();
 sg13g2_fill_2 FILLER_2_1806 ();
 sg13g2_decap_8 FILLER_2_1818 ();
 sg13g2_decap_8 FILLER_2_1825 ();
 sg13g2_decap_8 FILLER_2_1832 ();
 sg13g2_fill_2 FILLER_2_1839 ();
 sg13g2_decap_8 FILLER_2_1865 ();
 sg13g2_decap_8 FILLER_2_1872 ();
 sg13g2_decap_8 FILLER_2_1879 ();
 sg13g2_decap_4 FILLER_2_1886 ();
 sg13g2_fill_2 FILLER_2_1890 ();
 sg13g2_fill_1 FILLER_2_1902 ();
 sg13g2_decap_8 FILLER_2_1925 ();
 sg13g2_decap_8 FILLER_2_1932 ();
 sg13g2_decap_8 FILLER_2_1939 ();
 sg13g2_decap_8 FILLER_2_1946 ();
 sg13g2_decap_8 FILLER_2_1953 ();
 sg13g2_decap_8 FILLER_2_1960 ();
 sg13g2_decap_4 FILLER_2_1967 ();
 sg13g2_fill_1 FILLER_2_1971 ();
 sg13g2_decap_4 FILLER_2_1982 ();
 sg13g2_decap_4 FILLER_2_1995 ();
 sg13g2_fill_1 FILLER_2_2025 ();
 sg13g2_fill_2 FILLER_2_2060 ();
 sg13g2_decap_8 FILLER_2_2095 ();
 sg13g2_decap_8 FILLER_2_2102 ();
 sg13g2_fill_2 FILLER_2_2109 ();
 sg13g2_fill_1 FILLER_2_2111 ();
 sg13g2_decap_8 FILLER_2_2138 ();
 sg13g2_fill_2 FILLER_2_2150 ();
 sg13g2_fill_2 FILLER_2_2178 ();
 sg13g2_fill_1 FILLER_2_2180 ();
 sg13g2_decap_8 FILLER_2_2207 ();
 sg13g2_decap_8 FILLER_2_2214 ();
 sg13g2_fill_1 FILLER_2_2221 ();
 sg13g2_decap_8 FILLER_2_2248 ();
 sg13g2_decap_8 FILLER_2_2255 ();
 sg13g2_decap_8 FILLER_2_2262 ();
 sg13g2_decap_8 FILLER_2_2269 ();
 sg13g2_decap_4 FILLER_2_2276 ();
 sg13g2_fill_1 FILLER_2_2280 ();
 sg13g2_fill_2 FILLER_2_2307 ();
 sg13g2_decap_8 FILLER_2_2371 ();
 sg13g2_decap_4 FILLER_2_2378 ();
 sg13g2_fill_1 FILLER_2_2382 ();
 sg13g2_decap_8 FILLER_2_2435 ();
 sg13g2_decap_4 FILLER_2_2442 ();
 sg13g2_fill_1 FILLER_2_2446 ();
 sg13g2_decap_8 FILLER_2_2499 ();
 sg13g2_fill_2 FILLER_2_2506 ();
 sg13g2_decap_8 FILLER_2_2534 ();
 sg13g2_fill_1 FILLER_2_2541 ();
 sg13g2_decap_4 FILLER_2_2594 ();
 sg13g2_fill_2 FILLER_2_2602 ();
 sg13g2_fill_1 FILLER_2_2604 ();
 sg13g2_fill_2 FILLER_2_2657 ();
 sg13g2_fill_1 FILLER_2_2659 ();
 sg13g2_fill_2 FILLER_2_2686 ();
 sg13g2_decap_4 FILLER_2_2698 ();
 sg13g2_fill_1 FILLER_2_2728 ();
 sg13g2_decap_8 FILLER_2_2755 ();
 sg13g2_decap_8 FILLER_2_2762 ();
 sg13g2_decap_8 FILLER_2_2769 ();
 sg13g2_decap_4 FILLER_2_2776 ();
 sg13g2_fill_2 FILLER_2_2806 ();
 sg13g2_fill_1 FILLER_2_2808 ();
 sg13g2_fill_1 FILLER_2_2835 ();
 sg13g2_decap_8 FILLER_2_2862 ();
 sg13g2_decap_4 FILLER_2_2869 ();
 sg13g2_fill_2 FILLER_2_2873 ();
 sg13g2_decap_8 FILLER_2_2927 ();
 sg13g2_decap_8 FILLER_2_2934 ();
 sg13g2_decap_8 FILLER_2_2941 ();
 sg13g2_decap_8 FILLER_2_2948 ();
 sg13g2_decap_8 FILLER_2_2955 ();
 sg13g2_decap_8 FILLER_2_2962 ();
 sg13g2_decap_8 FILLER_2_2969 ();
 sg13g2_decap_4 FILLER_2_2976 ();
 sg13g2_decap_8 FILLER_2_3028 ();
 sg13g2_decap_8 FILLER_2_3035 ();
 sg13g2_decap_4 FILLER_2_3042 ();
 sg13g2_decap_8 FILLER_2_3064 ();
 sg13g2_decap_4 FILLER_2_3071 ();
 sg13g2_fill_1 FILLER_2_3075 ();
 sg13g2_fill_1 FILLER_2_3106 ();
 sg13g2_decap_8 FILLER_2_3143 ();
 sg13g2_decap_4 FILLER_2_3150 ();
 sg13g2_fill_2 FILLER_2_3154 ();
 sg13g2_decap_8 FILLER_2_3174 ();
 sg13g2_decap_8 FILLER_2_3181 ();
 sg13g2_decap_8 FILLER_2_3188 ();
 sg13g2_decap_8 FILLER_2_3195 ();
 sg13g2_fill_2 FILLER_2_3202 ();
 sg13g2_decap_8 FILLER_2_3230 ();
 sg13g2_decap_8 FILLER_2_3237 ();
 sg13g2_decap_8 FILLER_2_3244 ();
 sg13g2_decap_8 FILLER_2_3251 ();
 sg13g2_decap_8 FILLER_2_3258 ();
 sg13g2_decap_8 FILLER_2_3265 ();
 sg13g2_decap_8 FILLER_2_3272 ();
 sg13g2_decap_8 FILLER_2_3279 ();
 sg13g2_decap_8 FILLER_2_3286 ();
 sg13g2_decap_8 FILLER_2_3293 ();
 sg13g2_decap_8 FILLER_2_3300 ();
 sg13g2_decap_8 FILLER_2_3307 ();
 sg13g2_decap_8 FILLER_2_3314 ();
 sg13g2_decap_8 FILLER_2_3321 ();
 sg13g2_decap_8 FILLER_2_3328 ();
 sg13g2_decap_8 FILLER_2_3335 ();
 sg13g2_decap_8 FILLER_2_3342 ();
 sg13g2_decap_8 FILLER_2_3349 ();
 sg13g2_decap_8 FILLER_2_3356 ();
 sg13g2_decap_8 FILLER_2_3363 ();
 sg13g2_decap_8 FILLER_2_3370 ();
 sg13g2_decap_8 FILLER_2_3377 ();
 sg13g2_decap_8 FILLER_2_3384 ();
 sg13g2_decap_8 FILLER_2_3391 ();
 sg13g2_decap_8 FILLER_2_3398 ();
 sg13g2_decap_8 FILLER_2_3405 ();
 sg13g2_decap_8 FILLER_2_3412 ();
 sg13g2_decap_8 FILLER_2_3419 ();
 sg13g2_decap_8 FILLER_2_3426 ();
 sg13g2_decap_8 FILLER_2_3433 ();
 sg13g2_decap_8 FILLER_2_3440 ();
 sg13g2_decap_8 FILLER_2_3447 ();
 sg13g2_decap_8 FILLER_2_3454 ();
 sg13g2_decap_8 FILLER_2_3461 ();
 sg13g2_decap_8 FILLER_2_3468 ();
 sg13g2_decap_8 FILLER_2_3475 ();
 sg13g2_decap_8 FILLER_2_3482 ();
 sg13g2_decap_8 FILLER_2_3489 ();
 sg13g2_decap_8 FILLER_2_3496 ();
 sg13g2_decap_8 FILLER_2_3503 ();
 sg13g2_decap_8 FILLER_2_3510 ();
 sg13g2_decap_8 FILLER_2_3517 ();
 sg13g2_decap_8 FILLER_2_3524 ();
 sg13g2_decap_8 FILLER_2_3531 ();
 sg13g2_decap_8 FILLER_2_3538 ();
 sg13g2_decap_8 FILLER_2_3545 ();
 sg13g2_decap_8 FILLER_2_3552 ();
 sg13g2_decap_8 FILLER_2_3559 ();
 sg13g2_decap_8 FILLER_2_3566 ();
 sg13g2_decap_8 FILLER_2_3573 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_fill_2 FILLER_3_56 ();
 sg13g2_fill_1 FILLER_3_58 ();
 sg13g2_decap_8 FILLER_3_117 ();
 sg13g2_decap_8 FILLER_3_124 ();
 sg13g2_decap_8 FILLER_3_131 ();
 sg13g2_decap_8 FILLER_3_138 ();
 sg13g2_decap_8 FILLER_3_145 ();
 sg13g2_decap_8 FILLER_3_152 ();
 sg13g2_decap_4 FILLER_3_159 ();
 sg13g2_fill_2 FILLER_3_172 ();
 sg13g2_fill_1 FILLER_3_184 ();
 sg13g2_fill_2 FILLER_3_207 ();
 sg13g2_fill_1 FILLER_3_209 ();
 sg13g2_decap_8 FILLER_3_219 ();
 sg13g2_decap_8 FILLER_3_226 ();
 sg13g2_decap_8 FILLER_3_233 ();
 sg13g2_fill_1 FILLER_3_271 ();
 sg13g2_decap_8 FILLER_3_291 ();
 sg13g2_decap_8 FILLER_3_298 ();
 sg13g2_decap_8 FILLER_3_305 ();
 sg13g2_decap_8 FILLER_3_312 ();
 sg13g2_decap_8 FILLER_3_319 ();
 sg13g2_fill_2 FILLER_3_326 ();
 sg13g2_fill_1 FILLER_3_328 ();
 sg13g2_decap_8 FILLER_3_359 ();
 sg13g2_decap_8 FILLER_3_366 ();
 sg13g2_decap_8 FILLER_3_373 ();
 sg13g2_decap_8 FILLER_3_380 ();
 sg13g2_decap_8 FILLER_3_387 ();
 sg13g2_fill_1 FILLER_3_394 ();
 sg13g2_decap_8 FILLER_3_416 ();
 sg13g2_decap_4 FILLER_3_423 ();
 sg13g2_decap_8 FILLER_3_437 ();
 sg13g2_decap_8 FILLER_3_444 ();
 sg13g2_decap_8 FILLER_3_451 ();
 sg13g2_decap_8 FILLER_3_458 ();
 sg13g2_decap_8 FILLER_3_465 ();
 sg13g2_decap_4 FILLER_3_472 ();
 sg13g2_fill_2 FILLER_3_476 ();
 sg13g2_decap_8 FILLER_3_488 ();
 sg13g2_decap_8 FILLER_3_495 ();
 sg13g2_fill_2 FILLER_3_502 ();
 sg13g2_decap_8 FILLER_3_508 ();
 sg13g2_decap_8 FILLER_3_515 ();
 sg13g2_decap_8 FILLER_3_522 ();
 sg13g2_decap_8 FILLER_3_529 ();
 sg13g2_decap_8 FILLER_3_536 ();
 sg13g2_decap_8 FILLER_3_543 ();
 sg13g2_decap_8 FILLER_3_550 ();
 sg13g2_decap_8 FILLER_3_557 ();
 sg13g2_fill_2 FILLER_3_564 ();
 sg13g2_fill_1 FILLER_3_566 ();
 sg13g2_decap_8 FILLER_3_577 ();
 sg13g2_decap_8 FILLER_3_584 ();
 sg13g2_fill_2 FILLER_3_591 ();
 sg13g2_fill_1 FILLER_3_593 ();
 sg13g2_decap_8 FILLER_3_604 ();
 sg13g2_decap_8 FILLER_3_611 ();
 sg13g2_decap_8 FILLER_3_618 ();
 sg13g2_decap_8 FILLER_3_625 ();
 sg13g2_decap_8 FILLER_3_632 ();
 sg13g2_fill_2 FILLER_3_639 ();
 sg13g2_decap_8 FILLER_3_680 ();
 sg13g2_decap_8 FILLER_3_687 ();
 sg13g2_fill_2 FILLER_3_694 ();
 sg13g2_fill_1 FILLER_3_696 ();
 sg13g2_fill_2 FILLER_3_717 ();
 sg13g2_fill_1 FILLER_3_719 ();
 sg13g2_decap_8 FILLER_3_730 ();
 sg13g2_decap_8 FILLER_3_737 ();
 sg13g2_decap_8 FILLER_3_744 ();
 sg13g2_decap_8 FILLER_3_751 ();
 sg13g2_fill_2 FILLER_3_758 ();
 sg13g2_decap_8 FILLER_3_786 ();
 sg13g2_decap_8 FILLER_3_793 ();
 sg13g2_decap_8 FILLER_3_800 ();
 sg13g2_decap_8 FILLER_3_807 ();
 sg13g2_decap_8 FILLER_3_814 ();
 sg13g2_decap_8 FILLER_3_821 ();
 sg13g2_fill_1 FILLER_3_828 ();
 sg13g2_decap_8 FILLER_3_855 ();
 sg13g2_decap_8 FILLER_3_862 ();
 sg13g2_decap_8 FILLER_3_869 ();
 sg13g2_decap_8 FILLER_3_876 ();
 sg13g2_decap_4 FILLER_3_883 ();
 sg13g2_fill_1 FILLER_3_887 ();
 sg13g2_decap_8 FILLER_3_898 ();
 sg13g2_decap_8 FILLER_3_905 ();
 sg13g2_decap_8 FILLER_3_912 ();
 sg13g2_decap_8 FILLER_3_919 ();
 sg13g2_decap_8 FILLER_3_926 ();
 sg13g2_decap_8 FILLER_3_933 ();
 sg13g2_decap_8 FILLER_3_940 ();
 sg13g2_fill_2 FILLER_3_947 ();
 sg13g2_decap_4 FILLER_3_954 ();
 sg13g2_fill_2 FILLER_3_958 ();
 sg13g2_decap_4 FILLER_3_968 ();
 sg13g2_fill_1 FILLER_3_972 ();
 sg13g2_decap_8 FILLER_3_983 ();
 sg13g2_decap_8 FILLER_3_990 ();
 sg13g2_decap_8 FILLER_3_997 ();
 sg13g2_decap_8 FILLER_3_1004 ();
 sg13g2_decap_8 FILLER_3_1011 ();
 sg13g2_decap_8 FILLER_3_1018 ();
 sg13g2_decap_8 FILLER_3_1025 ();
 sg13g2_decap_8 FILLER_3_1032 ();
 sg13g2_decap_4 FILLER_3_1039 ();
 sg13g2_decap_8 FILLER_3_1066 ();
 sg13g2_decap_8 FILLER_3_1073 ();
 sg13g2_fill_1 FILLER_3_1080 ();
 sg13g2_decap_8 FILLER_3_1107 ();
 sg13g2_decap_8 FILLER_3_1114 ();
 sg13g2_decap_8 FILLER_3_1121 ();
 sg13g2_decap_4 FILLER_3_1128 ();
 sg13g2_fill_1 FILLER_3_1132 ();
 sg13g2_decap_8 FILLER_3_1158 ();
 sg13g2_decap_8 FILLER_3_1165 ();
 sg13g2_decap_8 FILLER_3_1172 ();
 sg13g2_decap_4 FILLER_3_1179 ();
 sg13g2_fill_2 FILLER_3_1183 ();
 sg13g2_fill_1 FILLER_3_1193 ();
 sg13g2_decap_8 FILLER_3_1204 ();
 sg13g2_decap_8 FILLER_3_1211 ();
 sg13g2_decap_8 FILLER_3_1218 ();
 sg13g2_decap_8 FILLER_3_1225 ();
 sg13g2_decap_8 FILLER_3_1232 ();
 sg13g2_fill_2 FILLER_3_1239 ();
 sg13g2_fill_2 FILLER_3_1259 ();
 sg13g2_decap_8 FILLER_3_1271 ();
 sg13g2_decap_8 FILLER_3_1278 ();
 sg13g2_decap_8 FILLER_3_1285 ();
 sg13g2_decap_8 FILLER_3_1292 ();
 sg13g2_fill_1 FILLER_3_1299 ();
 sg13g2_fill_1 FILLER_3_1308 ();
 sg13g2_fill_1 FILLER_3_1319 ();
 sg13g2_decap_8 FILLER_3_1325 ();
 sg13g2_decap_8 FILLER_3_1332 ();
 sg13g2_decap_8 FILLER_3_1339 ();
 sg13g2_decap_8 FILLER_3_1346 ();
 sg13g2_fill_2 FILLER_3_1353 ();
 sg13g2_decap_8 FILLER_3_1370 ();
 sg13g2_decap_8 FILLER_3_1377 ();
 sg13g2_decap_8 FILLER_3_1384 ();
 sg13g2_decap_8 FILLER_3_1391 ();
 sg13g2_decap_8 FILLER_3_1398 ();
 sg13g2_decap_8 FILLER_3_1405 ();
 sg13g2_decap_8 FILLER_3_1412 ();
 sg13g2_decap_8 FILLER_3_1445 ();
 sg13g2_decap_8 FILLER_3_1452 ();
 sg13g2_decap_8 FILLER_3_1459 ();
 sg13g2_fill_1 FILLER_3_1466 ();
 sg13g2_decap_8 FILLER_3_1471 ();
 sg13g2_fill_2 FILLER_3_1478 ();
 sg13g2_fill_2 FILLER_3_1506 ();
 sg13g2_decap_8 FILLER_3_1544 ();
 sg13g2_fill_2 FILLER_3_1551 ();
 sg13g2_decap_8 FILLER_3_1561 ();
 sg13g2_decap_4 FILLER_3_1568 ();
 sg13g2_fill_2 FILLER_3_1572 ();
 sg13g2_fill_2 FILLER_3_1584 ();
 sg13g2_decap_8 FILLER_3_1604 ();
 sg13g2_decap_8 FILLER_3_1611 ();
 sg13g2_decap_8 FILLER_3_1618 ();
 sg13g2_decap_8 FILLER_3_1625 ();
 sg13g2_decap_8 FILLER_3_1632 ();
 sg13g2_decap_4 FILLER_3_1639 ();
 sg13g2_fill_1 FILLER_3_1643 ();
 sg13g2_fill_1 FILLER_3_1647 ();
 sg13g2_fill_2 FILLER_3_1657 ();
 sg13g2_fill_1 FILLER_3_1659 ();
 sg13g2_decap_8 FILLER_3_1670 ();
 sg13g2_decap_8 FILLER_3_1677 ();
 sg13g2_decap_8 FILLER_3_1684 ();
 sg13g2_decap_4 FILLER_3_1691 ();
 sg13g2_decap_8 FILLER_3_1705 ();
 sg13g2_decap_8 FILLER_3_1712 ();
 sg13g2_decap_8 FILLER_3_1719 ();
 sg13g2_decap_8 FILLER_3_1726 ();
 sg13g2_decap_8 FILLER_3_1733 ();
 sg13g2_decap_8 FILLER_3_1740 ();
 sg13g2_decap_8 FILLER_3_1747 ();
 sg13g2_fill_1 FILLER_3_1754 ();
 sg13g2_decap_8 FILLER_3_1781 ();
 sg13g2_fill_1 FILLER_3_1788 ();
 sg13g2_decap_4 FILLER_3_1802 ();
 sg13g2_fill_1 FILLER_3_1806 ();
 sg13g2_decap_8 FILLER_3_1816 ();
 sg13g2_decap_8 FILLER_3_1823 ();
 sg13g2_decap_8 FILLER_3_1830 ();
 sg13g2_decap_8 FILLER_3_1837 ();
 sg13g2_decap_8 FILLER_3_1844 ();
 sg13g2_decap_8 FILLER_3_1877 ();
 sg13g2_decap_8 FILLER_3_1884 ();
 sg13g2_decap_8 FILLER_3_1891 ();
 sg13g2_decap_8 FILLER_3_1898 ();
 sg13g2_decap_8 FILLER_3_1905 ();
 sg13g2_fill_2 FILLER_3_1912 ();
 sg13g2_decap_8 FILLER_3_1940 ();
 sg13g2_decap_8 FILLER_3_1947 ();
 sg13g2_decap_8 FILLER_3_1954 ();
 sg13g2_decap_8 FILLER_3_1961 ();
 sg13g2_fill_2 FILLER_3_1968 ();
 sg13g2_decap_8 FILLER_3_1996 ();
 sg13g2_decap_4 FILLER_3_2003 ();
 sg13g2_decap_8 FILLER_3_2017 ();
 sg13g2_decap_8 FILLER_3_2024 ();
 sg13g2_decap_8 FILLER_3_2070 ();
 sg13g2_decap_4 FILLER_3_2077 ();
 sg13g2_decap_8 FILLER_3_2096 ();
 sg13g2_decap_8 FILLER_3_2103 ();
 sg13g2_decap_8 FILLER_3_2110 ();
 sg13g2_fill_1 FILLER_3_2117 ();
 sg13g2_decap_8 FILLER_3_2158 ();
 sg13g2_decap_4 FILLER_3_2165 ();
 sg13g2_decap_8 FILLER_3_2174 ();
 sg13g2_fill_2 FILLER_3_2186 ();
 sg13g2_fill_2 FILLER_3_2210 ();
 sg13g2_fill_2 FILLER_3_2232 ();
 sg13g2_fill_1 FILLER_3_2234 ();
 sg13g2_decap_8 FILLER_3_2240 ();
 sg13g2_decap_4 FILLER_3_2247 ();
 sg13g2_fill_2 FILLER_3_2251 ();
 sg13g2_decap_4 FILLER_3_2258 ();
 sg13g2_decap_4 FILLER_3_2266 ();
 sg13g2_fill_1 FILLER_3_2270 ();
 sg13g2_fill_2 FILLER_3_2275 ();
 sg13g2_fill_1 FILLER_3_2277 ();
 sg13g2_decap_8 FILLER_3_2292 ();
 sg13g2_decap_8 FILLER_3_2299 ();
 sg13g2_decap_4 FILLER_3_2306 ();
 sg13g2_decap_8 FILLER_3_2326 ();
 sg13g2_decap_8 FILLER_3_2343 ();
 sg13g2_decap_4 FILLER_3_2350 ();
 sg13g2_decap_8 FILLER_3_2362 ();
 sg13g2_decap_8 FILLER_3_2369 ();
 sg13g2_decap_8 FILLER_3_2376 ();
 sg13g2_decap_8 FILLER_3_2383 ();
 sg13g2_fill_2 FILLER_3_2390 ();
 sg13g2_fill_2 FILLER_3_2401 ();
 sg13g2_fill_1 FILLER_3_2403 ();
 sg13g2_fill_2 FILLER_3_2412 ();
 sg13g2_decap_8 FILLER_3_2433 ();
 sg13g2_decap_8 FILLER_3_2440 ();
 sg13g2_decap_8 FILLER_3_2447 ();
 sg13g2_decap_8 FILLER_3_2454 ();
 sg13g2_decap_4 FILLER_3_2461 ();
 sg13g2_decap_8 FILLER_3_2502 ();
 sg13g2_decap_8 FILLER_3_2535 ();
 sg13g2_decap_8 FILLER_3_2542 ();
 sg13g2_decap_8 FILLER_3_2549 ();
 sg13g2_decap_4 FILLER_3_2556 ();
 sg13g2_fill_1 FILLER_3_2560 ();
 sg13g2_decap_4 FILLER_3_2578 ();
 sg13g2_decap_8 FILLER_3_2591 ();
 sg13g2_decap_8 FILLER_3_2598 ();
 sg13g2_fill_2 FILLER_3_2605 ();
 sg13g2_fill_1 FILLER_3_2607 ();
 sg13g2_fill_2 FILLER_3_2613 ();
 sg13g2_decap_8 FILLER_3_2630 ();
 sg13g2_decap_8 FILLER_3_2637 ();
 sg13g2_decap_8 FILLER_3_2644 ();
 sg13g2_decap_4 FILLER_3_2690 ();
 sg13g2_decap_8 FILLER_3_2702 ();
 sg13g2_decap_8 FILLER_3_2709 ();
 sg13g2_fill_2 FILLER_3_2716 ();
 sg13g2_fill_1 FILLER_3_2718 ();
 sg13g2_decap_8 FILLER_3_2757 ();
 sg13g2_decap_8 FILLER_3_2764 ();
 sg13g2_decap_8 FILLER_3_2771 ();
 sg13g2_fill_2 FILLER_3_2778 ();
 sg13g2_fill_1 FILLER_3_2780 ();
 sg13g2_decap_8 FILLER_3_2809 ();
 sg13g2_decap_8 FILLER_3_2816 ();
 sg13g2_decap_4 FILLER_3_2823 ();
 sg13g2_fill_1 FILLER_3_2827 ();
 sg13g2_fill_2 FILLER_3_2842 ();
 sg13g2_decap_8 FILLER_3_2862 ();
 sg13g2_decap_8 FILLER_3_2869 ();
 sg13g2_decap_8 FILLER_3_2876 ();
 sg13g2_fill_2 FILLER_3_2883 ();
 sg13g2_decap_8 FILLER_3_2911 ();
 sg13g2_decap_8 FILLER_3_2918 ();
 sg13g2_decap_8 FILLER_3_2925 ();
 sg13g2_fill_2 FILLER_3_2932 ();
 sg13g2_decap_8 FILLER_3_2960 ();
 sg13g2_decap_8 FILLER_3_2967 ();
 sg13g2_decap_8 FILLER_3_2974 ();
 sg13g2_decap_8 FILLER_3_2981 ();
 sg13g2_decap_8 FILLER_3_3007 ();
 sg13g2_decap_8 FILLER_3_3014 ();
 sg13g2_decap_8 FILLER_3_3021 ();
 sg13g2_decap_4 FILLER_3_3028 ();
 sg13g2_fill_2 FILLER_3_3036 ();
 sg13g2_fill_1 FILLER_3_3064 ();
 sg13g2_decap_4 FILLER_3_3092 ();
 sg13g2_fill_2 FILLER_3_3096 ();
 sg13g2_decap_8 FILLER_3_3108 ();
 sg13g2_fill_1 FILLER_3_3115 ();
 sg13g2_decap_8 FILLER_3_3126 ();
 sg13g2_decap_8 FILLER_3_3133 ();
 sg13g2_decap_8 FILLER_3_3140 ();
 sg13g2_decap_8 FILLER_3_3147 ();
 sg13g2_decap_8 FILLER_3_3154 ();
 sg13g2_decap_4 FILLER_3_3161 ();
 sg13g2_fill_2 FILLER_3_3165 ();
 sg13g2_decap_8 FILLER_3_3172 ();
 sg13g2_decap_8 FILLER_3_3179 ();
 sg13g2_decap_8 FILLER_3_3186 ();
 sg13g2_decap_8 FILLER_3_3193 ();
 sg13g2_decap_8 FILLER_3_3200 ();
 sg13g2_decap_8 FILLER_3_3207 ();
 sg13g2_decap_8 FILLER_3_3214 ();
 sg13g2_fill_1 FILLER_3_3221 ();
 sg13g2_decap_8 FILLER_3_3225 ();
 sg13g2_decap_8 FILLER_3_3232 ();
 sg13g2_decap_8 FILLER_3_3239 ();
 sg13g2_decap_8 FILLER_3_3246 ();
 sg13g2_decap_8 FILLER_3_3253 ();
 sg13g2_decap_8 FILLER_3_3260 ();
 sg13g2_decap_8 FILLER_3_3267 ();
 sg13g2_decap_8 FILLER_3_3274 ();
 sg13g2_decap_8 FILLER_3_3281 ();
 sg13g2_decap_8 FILLER_3_3288 ();
 sg13g2_decap_8 FILLER_3_3295 ();
 sg13g2_decap_8 FILLER_3_3302 ();
 sg13g2_decap_8 FILLER_3_3309 ();
 sg13g2_decap_8 FILLER_3_3316 ();
 sg13g2_decap_8 FILLER_3_3323 ();
 sg13g2_decap_8 FILLER_3_3330 ();
 sg13g2_decap_8 FILLER_3_3337 ();
 sg13g2_decap_8 FILLER_3_3344 ();
 sg13g2_decap_8 FILLER_3_3351 ();
 sg13g2_decap_8 FILLER_3_3358 ();
 sg13g2_decap_8 FILLER_3_3365 ();
 sg13g2_decap_8 FILLER_3_3372 ();
 sg13g2_decap_8 FILLER_3_3379 ();
 sg13g2_decap_8 FILLER_3_3386 ();
 sg13g2_decap_8 FILLER_3_3393 ();
 sg13g2_decap_8 FILLER_3_3400 ();
 sg13g2_decap_8 FILLER_3_3407 ();
 sg13g2_decap_8 FILLER_3_3414 ();
 sg13g2_decap_8 FILLER_3_3421 ();
 sg13g2_decap_8 FILLER_3_3428 ();
 sg13g2_decap_8 FILLER_3_3435 ();
 sg13g2_decap_8 FILLER_3_3442 ();
 sg13g2_decap_8 FILLER_3_3449 ();
 sg13g2_decap_8 FILLER_3_3456 ();
 sg13g2_decap_8 FILLER_3_3463 ();
 sg13g2_decap_8 FILLER_3_3470 ();
 sg13g2_decap_8 FILLER_3_3477 ();
 sg13g2_decap_8 FILLER_3_3484 ();
 sg13g2_decap_8 FILLER_3_3491 ();
 sg13g2_decap_8 FILLER_3_3498 ();
 sg13g2_decap_8 FILLER_3_3505 ();
 sg13g2_decap_8 FILLER_3_3512 ();
 sg13g2_decap_8 FILLER_3_3519 ();
 sg13g2_decap_8 FILLER_3_3526 ();
 sg13g2_decap_8 FILLER_3_3533 ();
 sg13g2_decap_8 FILLER_3_3540 ();
 sg13g2_decap_8 FILLER_3_3547 ();
 sg13g2_decap_8 FILLER_3_3554 ();
 sg13g2_decap_8 FILLER_3_3561 ();
 sg13g2_decap_8 FILLER_3_3568 ();
 sg13g2_decap_4 FILLER_3_3575 ();
 sg13g2_fill_1 FILLER_3_3579 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_4 FILLER_4_63 ();
 sg13g2_fill_2 FILLER_4_67 ();
 sg13g2_fill_1 FILLER_4_83 ();
 sg13g2_decap_8 FILLER_4_102 ();
 sg13g2_decap_8 FILLER_4_109 ();
 sg13g2_decap_8 FILLER_4_116 ();
 sg13g2_decap_8 FILLER_4_123 ();
 sg13g2_decap_8 FILLER_4_130 ();
 sg13g2_decap_8 FILLER_4_137 ();
 sg13g2_decap_8 FILLER_4_144 ();
 sg13g2_fill_2 FILLER_4_151 ();
 sg13g2_fill_2 FILLER_4_179 ();
 sg13g2_fill_1 FILLER_4_181 ();
 sg13g2_fill_2 FILLER_4_191 ();
 sg13g2_fill_1 FILLER_4_193 ();
 sg13g2_fill_2 FILLER_4_204 ();
 sg13g2_fill_1 FILLER_4_206 ();
 sg13g2_decap_8 FILLER_4_216 ();
 sg13g2_decap_8 FILLER_4_223 ();
 sg13g2_decap_8 FILLER_4_230 ();
 sg13g2_decap_8 FILLER_4_237 ();
 sg13g2_fill_2 FILLER_4_244 ();
 sg13g2_decap_4 FILLER_4_255 ();
 sg13g2_fill_1 FILLER_4_264 ();
 sg13g2_fill_2 FILLER_4_274 ();
 sg13g2_fill_1 FILLER_4_276 ();
 sg13g2_decap_8 FILLER_4_281 ();
 sg13g2_fill_1 FILLER_4_288 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_4 FILLER_4_329 ();
 sg13g2_fill_1 FILLER_4_333 ();
 sg13g2_decap_8 FILLER_4_386 ();
 sg13g2_decap_4 FILLER_4_393 ();
 sg13g2_fill_1 FILLER_4_397 ();
 sg13g2_fill_1 FILLER_4_403 ();
 sg13g2_decap_8 FILLER_4_409 ();
 sg13g2_decap_4 FILLER_4_416 ();
 sg13g2_fill_2 FILLER_4_430 ();
 sg13g2_fill_1 FILLER_4_432 ();
 sg13g2_decap_8 FILLER_4_438 ();
 sg13g2_decap_8 FILLER_4_455 ();
 sg13g2_fill_2 FILLER_4_462 ();
 sg13g2_decap_8 FILLER_4_474 ();
 sg13g2_fill_1 FILLER_4_481 ();
 sg13g2_fill_1 FILLER_4_535 ();
 sg13g2_decap_8 FILLER_4_572 ();
 sg13g2_decap_8 FILLER_4_579 ();
 sg13g2_decap_8 FILLER_4_586 ();
 sg13g2_decap_8 FILLER_4_593 ();
 sg13g2_decap_4 FILLER_4_600 ();
 sg13g2_fill_2 FILLER_4_604 ();
 sg13g2_decap_8 FILLER_4_627 ();
 sg13g2_fill_1 FILLER_4_634 ();
 sg13g2_decap_8 FILLER_4_640 ();
 sg13g2_decap_4 FILLER_4_647 ();
 sg13g2_fill_1 FILLER_4_651 ();
 sg13g2_decap_4 FILLER_4_662 ();
 sg13g2_fill_2 FILLER_4_666 ();
 sg13g2_decap_8 FILLER_4_677 ();
 sg13g2_decap_8 FILLER_4_684 ();
 sg13g2_decap_8 FILLER_4_691 ();
 sg13g2_decap_8 FILLER_4_698 ();
 sg13g2_decap_8 FILLER_4_705 ();
 sg13g2_decap_8 FILLER_4_712 ();
 sg13g2_decap_8 FILLER_4_719 ();
 sg13g2_decap_8 FILLER_4_747 ();
 sg13g2_decap_8 FILLER_4_754 ();
 sg13g2_decap_8 FILLER_4_761 ();
 sg13g2_decap_8 FILLER_4_768 ();
 sg13g2_decap_8 FILLER_4_775 ();
 sg13g2_decap_8 FILLER_4_782 ();
 sg13g2_decap_8 FILLER_4_789 ();
 sg13g2_decap_4 FILLER_4_796 ();
 sg13g2_decap_8 FILLER_4_805 ();
 sg13g2_decap_8 FILLER_4_812 ();
 sg13g2_decap_8 FILLER_4_819 ();
 sg13g2_decap_4 FILLER_4_826 ();
 sg13g2_decap_8 FILLER_4_840 ();
 sg13g2_decap_8 FILLER_4_847 ();
 sg13g2_decap_8 FILLER_4_854 ();
 sg13g2_decap_8 FILLER_4_861 ();
 sg13g2_decap_8 FILLER_4_868 ();
 sg13g2_decap_8 FILLER_4_875 ();
 sg13g2_fill_1 FILLER_4_882 ();
 sg13g2_decap_8 FILLER_4_903 ();
 sg13g2_decap_8 FILLER_4_930 ();
 sg13g2_decap_8 FILLER_4_937 ();
 sg13g2_decap_8 FILLER_4_944 ();
 sg13g2_decap_8 FILLER_4_951 ();
 sg13g2_decap_4 FILLER_4_958 ();
 sg13g2_decap_8 FILLER_4_993 ();
 sg13g2_decap_4 FILLER_4_1000 ();
 sg13g2_fill_2 FILLER_4_1004 ();
 sg13g2_decap_8 FILLER_4_1032 ();
 sg13g2_decap_8 FILLER_4_1039 ();
 sg13g2_fill_2 FILLER_4_1046 ();
 sg13g2_fill_1 FILLER_4_1048 ();
 sg13g2_decap_8 FILLER_4_1053 ();
 sg13g2_decap_8 FILLER_4_1060 ();
 sg13g2_decap_8 FILLER_4_1067 ();
 sg13g2_decap_4 FILLER_4_1074 ();
 sg13g2_fill_1 FILLER_4_1078 ();
 sg13g2_decap_8 FILLER_4_1089 ();
 sg13g2_decap_8 FILLER_4_1096 ();
 sg13g2_decap_8 FILLER_4_1103 ();
 sg13g2_decap_8 FILLER_4_1110 ();
 sg13g2_decap_8 FILLER_4_1117 ();
 sg13g2_decap_8 FILLER_4_1124 ();
 sg13g2_fill_2 FILLER_4_1131 ();
 sg13g2_decap_8 FILLER_4_1147 ();
 sg13g2_decap_8 FILLER_4_1154 ();
 sg13g2_decap_8 FILLER_4_1161 ();
 sg13g2_decap_8 FILLER_4_1168 ();
 sg13g2_decap_8 FILLER_4_1175 ();
 sg13g2_decap_4 FILLER_4_1182 ();
 sg13g2_fill_2 FILLER_4_1186 ();
 sg13g2_decap_8 FILLER_4_1191 ();
 sg13g2_decap_8 FILLER_4_1198 ();
 sg13g2_decap_8 FILLER_4_1205 ();
 sg13g2_decap_8 FILLER_4_1212 ();
 sg13g2_decap_8 FILLER_4_1219 ();
 sg13g2_decap_8 FILLER_4_1226 ();
 sg13g2_decap_8 FILLER_4_1233 ();
 sg13g2_decap_4 FILLER_4_1240 ();
 sg13g2_fill_1 FILLER_4_1244 ();
 sg13g2_fill_2 FILLER_4_1250 ();
 sg13g2_fill_1 FILLER_4_1252 ();
 sg13g2_decap_8 FILLER_4_1258 ();
 sg13g2_decap_8 FILLER_4_1265 ();
 sg13g2_decap_8 FILLER_4_1272 ();
 sg13g2_decap_8 FILLER_4_1279 ();
 sg13g2_decap_8 FILLER_4_1286 ();
 sg13g2_decap_8 FILLER_4_1293 ();
 sg13g2_decap_4 FILLER_4_1300 ();
 sg13g2_fill_1 FILLER_4_1304 ();
 sg13g2_decap_8 FILLER_4_1310 ();
 sg13g2_decap_8 FILLER_4_1317 ();
 sg13g2_decap_8 FILLER_4_1324 ();
 sg13g2_decap_8 FILLER_4_1331 ();
 sg13g2_decap_8 FILLER_4_1338 ();
 sg13g2_decap_8 FILLER_4_1345 ();
 sg13g2_decap_8 FILLER_4_1352 ();
 sg13g2_decap_8 FILLER_4_1359 ();
 sg13g2_decap_8 FILLER_4_1366 ();
 sg13g2_decap_8 FILLER_4_1373 ();
 sg13g2_decap_8 FILLER_4_1380 ();
 sg13g2_decap_8 FILLER_4_1387 ();
 sg13g2_decap_8 FILLER_4_1394 ();
 sg13g2_decap_8 FILLER_4_1401 ();
 sg13g2_decap_8 FILLER_4_1408 ();
 sg13g2_decap_4 FILLER_4_1415 ();
 sg13g2_decap_8 FILLER_4_1445 ();
 sg13g2_decap_8 FILLER_4_1452 ();
 sg13g2_decap_8 FILLER_4_1459 ();
 sg13g2_decap_8 FILLER_4_1466 ();
 sg13g2_decap_8 FILLER_4_1473 ();
 sg13g2_decap_8 FILLER_4_1480 ();
 sg13g2_fill_2 FILLER_4_1487 ();
 sg13g2_decap_8 FILLER_4_1493 ();
 sg13g2_decap_8 FILLER_4_1500 ();
 sg13g2_fill_2 FILLER_4_1507 ();
 sg13g2_decap_8 FILLER_4_1519 ();
 sg13g2_decap_8 FILLER_4_1526 ();
 sg13g2_decap_4 FILLER_4_1533 ();
 sg13g2_fill_1 FILLER_4_1537 ();
 sg13g2_decap_8 FILLER_4_1546 ();
 sg13g2_decap_8 FILLER_4_1553 ();
 sg13g2_decap_8 FILLER_4_1560 ();
 sg13g2_decap_8 FILLER_4_1567 ();
 sg13g2_decap_4 FILLER_4_1574 ();
 sg13g2_fill_1 FILLER_4_1578 ();
 sg13g2_decap_8 FILLER_4_1604 ();
 sg13g2_decap_8 FILLER_4_1611 ();
 sg13g2_decap_8 FILLER_4_1618 ();
 sg13g2_fill_2 FILLER_4_1625 ();
 sg13g2_decap_8 FILLER_4_1688 ();
 sg13g2_decap_8 FILLER_4_1695 ();
 sg13g2_decap_8 FILLER_4_1702 ();
 sg13g2_decap_8 FILLER_4_1709 ();
 sg13g2_decap_4 FILLER_4_1716 ();
 sg13g2_decap_8 FILLER_4_1746 ();
 sg13g2_decap_8 FILLER_4_1753 ();
 sg13g2_decap_8 FILLER_4_1760 ();
 sg13g2_decap_4 FILLER_4_1767 ();
 sg13g2_decap_8 FILLER_4_1779 ();
 sg13g2_decap_8 FILLER_4_1786 ();
 sg13g2_fill_2 FILLER_4_1793 ();
 sg13g2_fill_1 FILLER_4_1795 ();
 sg13g2_decap_8 FILLER_4_1801 ();
 sg13g2_decap_8 FILLER_4_1808 ();
 sg13g2_decap_8 FILLER_4_1815 ();
 sg13g2_decap_8 FILLER_4_1822 ();
 sg13g2_decap_8 FILLER_4_1829 ();
 sg13g2_decap_8 FILLER_4_1836 ();
 sg13g2_decap_8 FILLER_4_1843 ();
 sg13g2_decap_8 FILLER_4_1876 ();
 sg13g2_decap_8 FILLER_4_1883 ();
 sg13g2_decap_8 FILLER_4_1890 ();
 sg13g2_decap_8 FILLER_4_1897 ();
 sg13g2_decap_8 FILLER_4_1904 ();
 sg13g2_decap_4 FILLER_4_1911 ();
 sg13g2_fill_2 FILLER_4_1951 ();
 sg13g2_fill_1 FILLER_4_1953 ();
 sg13g2_decap_8 FILLER_4_1990 ();
 sg13g2_decap_8 FILLER_4_1997 ();
 sg13g2_fill_2 FILLER_4_2004 ();
 sg13g2_decap_8 FILLER_4_2015 ();
 sg13g2_decap_8 FILLER_4_2022 ();
 sg13g2_fill_1 FILLER_4_2042 ();
 sg13g2_decap_8 FILLER_4_2048 ();
 sg13g2_decap_8 FILLER_4_2055 ();
 sg13g2_decap_8 FILLER_4_2062 ();
 sg13g2_decap_4 FILLER_4_2069 ();
 sg13g2_decap_8 FILLER_4_2078 ();
 sg13g2_fill_2 FILLER_4_2085 ();
 sg13g2_fill_1 FILLER_4_2087 ();
 sg13g2_decap_8 FILLER_4_2098 ();
 sg13g2_decap_8 FILLER_4_2105 ();
 sg13g2_decap_8 FILLER_4_2112 ();
 sg13g2_fill_2 FILLER_4_2119 ();
 sg13g2_fill_1 FILLER_4_2121 ();
 sg13g2_decap_8 FILLER_4_2136 ();
 sg13g2_fill_1 FILLER_4_2143 ();
 sg13g2_decap_8 FILLER_4_2148 ();
 sg13g2_decap_8 FILLER_4_2155 ();
 sg13g2_decap_8 FILLER_4_2162 ();
 sg13g2_decap_8 FILLER_4_2169 ();
 sg13g2_fill_2 FILLER_4_2176 ();
 sg13g2_decap_8 FILLER_4_2187 ();
 sg13g2_decap_8 FILLER_4_2194 ();
 sg13g2_decap_8 FILLER_4_2201 ();
 sg13g2_decap_8 FILLER_4_2208 ();
 sg13g2_decap_8 FILLER_4_2215 ();
 sg13g2_decap_8 FILLER_4_2222 ();
 sg13g2_fill_2 FILLER_4_2229 ();
 sg13g2_fill_1 FILLER_4_2231 ();
 sg13g2_decap_8 FILLER_4_2240 ();
 sg13g2_decap_8 FILLER_4_2247 ();
 sg13g2_decap_8 FILLER_4_2259 ();
 sg13g2_fill_2 FILLER_4_2266 ();
 sg13g2_decap_8 FILLER_4_2304 ();
 sg13g2_decap_8 FILLER_4_2311 ();
 sg13g2_decap_8 FILLER_4_2318 ();
 sg13g2_decap_8 FILLER_4_2325 ();
 sg13g2_decap_8 FILLER_4_2332 ();
 sg13g2_decap_8 FILLER_4_2344 ();
 sg13g2_decap_8 FILLER_4_2351 ();
 sg13g2_decap_8 FILLER_4_2358 ();
 sg13g2_decap_8 FILLER_4_2365 ();
 sg13g2_decap_8 FILLER_4_2372 ();
 sg13g2_decap_4 FILLER_4_2384 ();
 sg13g2_fill_1 FILLER_4_2388 ();
 sg13g2_decap_8 FILLER_4_2428 ();
 sg13g2_decap_8 FILLER_4_2435 ();
 sg13g2_decap_8 FILLER_4_2442 ();
 sg13g2_decap_8 FILLER_4_2449 ();
 sg13g2_decap_8 FILLER_4_2456 ();
 sg13g2_fill_1 FILLER_4_2463 ();
 sg13g2_fill_2 FILLER_4_2473 ();
 sg13g2_fill_1 FILLER_4_2475 ();
 sg13g2_decap_8 FILLER_4_2489 ();
 sg13g2_decap_8 FILLER_4_2496 ();
 sg13g2_decap_8 FILLER_4_2503 ();
 sg13g2_fill_2 FILLER_4_2510 ();
 sg13g2_fill_1 FILLER_4_2512 ();
 sg13g2_decap_8 FILLER_4_2540 ();
 sg13g2_decap_8 FILLER_4_2547 ();
 sg13g2_decap_8 FILLER_4_2554 ();
 sg13g2_decap_8 FILLER_4_2571 ();
 sg13g2_decap_8 FILLER_4_2578 ();
 sg13g2_decap_8 FILLER_4_2585 ();
 sg13g2_fill_2 FILLER_4_2592 ();
 sg13g2_decap_8 FILLER_4_2630 ();
 sg13g2_decap_8 FILLER_4_2637 ();
 sg13g2_decap_8 FILLER_4_2644 ();
 sg13g2_decap_8 FILLER_4_2651 ();
 sg13g2_decap_8 FILLER_4_2658 ();
 sg13g2_decap_8 FILLER_4_2665 ();
 sg13g2_decap_8 FILLER_4_2672 ();
 sg13g2_decap_8 FILLER_4_2679 ();
 sg13g2_fill_2 FILLER_4_2686 ();
 sg13g2_decap_8 FILLER_4_2693 ();
 sg13g2_decap_8 FILLER_4_2700 ();
 sg13g2_decap_8 FILLER_4_2707 ();
 sg13g2_decap_8 FILLER_4_2714 ();
 sg13g2_decap_4 FILLER_4_2721 ();
 sg13g2_fill_2 FILLER_4_2725 ();
 sg13g2_decap_8 FILLER_4_2743 ();
 sg13g2_decap_8 FILLER_4_2750 ();
 sg13g2_decap_8 FILLER_4_2757 ();
 sg13g2_decap_8 FILLER_4_2764 ();
 sg13g2_decap_8 FILLER_4_2771 ();
 sg13g2_decap_8 FILLER_4_2778 ();
 sg13g2_decap_4 FILLER_4_2785 ();
 sg13g2_fill_2 FILLER_4_2793 ();
 sg13g2_decap_8 FILLER_4_2809 ();
 sg13g2_decap_8 FILLER_4_2816 ();
 sg13g2_decap_8 FILLER_4_2823 ();
 sg13g2_decap_4 FILLER_4_2830 ();
 sg13g2_fill_1 FILLER_4_2834 ();
 sg13g2_fill_2 FILLER_4_2840 ();
 sg13g2_decap_8 FILLER_4_2850 ();
 sg13g2_decap_8 FILLER_4_2857 ();
 sg13g2_decap_8 FILLER_4_2864 ();
 sg13g2_fill_1 FILLER_4_2871 ();
 sg13g2_decap_8 FILLER_4_2881 ();
 sg13g2_decap_8 FILLER_4_2888 ();
 sg13g2_decap_8 FILLER_4_2895 ();
 sg13g2_decap_8 FILLER_4_2902 ();
 sg13g2_decap_8 FILLER_4_2909 ();
 sg13g2_decap_4 FILLER_4_2916 ();
 sg13g2_fill_2 FILLER_4_2930 ();
 sg13g2_fill_1 FILLER_4_2932 ();
 sg13g2_decap_8 FILLER_4_2959 ();
 sg13g2_decap_8 FILLER_4_2966 ();
 sg13g2_decap_8 FILLER_4_2973 ();
 sg13g2_decap_4 FILLER_4_2980 ();
 sg13g2_fill_2 FILLER_4_2984 ();
 sg13g2_decap_8 FILLER_4_2991 ();
 sg13g2_decap_4 FILLER_4_2998 ();
 sg13g2_fill_1 FILLER_4_3002 ();
 sg13g2_decap_4 FILLER_4_3016 ();
 sg13g2_fill_2 FILLER_4_3020 ();
 sg13g2_fill_1 FILLER_4_3045 ();
 sg13g2_fill_2 FILLER_4_3057 ();
 sg13g2_decap_8 FILLER_4_3085 ();
 sg13g2_decap_8 FILLER_4_3092 ();
 sg13g2_decap_4 FILLER_4_3099 ();
 sg13g2_decap_8 FILLER_4_3129 ();
 sg13g2_decap_8 FILLER_4_3136 ();
 sg13g2_decap_8 FILLER_4_3143 ();
 sg13g2_decap_4 FILLER_4_3150 ();
 sg13g2_fill_2 FILLER_4_3154 ();
 sg13g2_decap_8 FILLER_4_3192 ();
 sg13g2_decap_8 FILLER_4_3199 ();
 sg13g2_decap_4 FILLER_4_3206 ();
 sg13g2_fill_2 FILLER_4_3210 ();
 sg13g2_decap_8 FILLER_4_3231 ();
 sg13g2_decap_8 FILLER_4_3238 ();
 sg13g2_decap_8 FILLER_4_3245 ();
 sg13g2_decap_8 FILLER_4_3252 ();
 sg13g2_decap_8 FILLER_4_3259 ();
 sg13g2_decap_8 FILLER_4_3266 ();
 sg13g2_decap_8 FILLER_4_3273 ();
 sg13g2_decap_8 FILLER_4_3280 ();
 sg13g2_decap_8 FILLER_4_3287 ();
 sg13g2_decap_8 FILLER_4_3294 ();
 sg13g2_decap_8 FILLER_4_3301 ();
 sg13g2_decap_8 FILLER_4_3308 ();
 sg13g2_decap_8 FILLER_4_3315 ();
 sg13g2_decap_8 FILLER_4_3322 ();
 sg13g2_decap_8 FILLER_4_3329 ();
 sg13g2_decap_8 FILLER_4_3336 ();
 sg13g2_decap_8 FILLER_4_3343 ();
 sg13g2_decap_8 FILLER_4_3350 ();
 sg13g2_decap_8 FILLER_4_3357 ();
 sg13g2_decap_8 FILLER_4_3364 ();
 sg13g2_decap_8 FILLER_4_3371 ();
 sg13g2_decap_8 FILLER_4_3378 ();
 sg13g2_decap_8 FILLER_4_3385 ();
 sg13g2_decap_8 FILLER_4_3392 ();
 sg13g2_decap_8 FILLER_4_3399 ();
 sg13g2_decap_8 FILLER_4_3406 ();
 sg13g2_decap_8 FILLER_4_3413 ();
 sg13g2_decap_8 FILLER_4_3420 ();
 sg13g2_decap_8 FILLER_4_3427 ();
 sg13g2_decap_8 FILLER_4_3434 ();
 sg13g2_decap_8 FILLER_4_3441 ();
 sg13g2_decap_8 FILLER_4_3448 ();
 sg13g2_decap_8 FILLER_4_3455 ();
 sg13g2_decap_8 FILLER_4_3462 ();
 sg13g2_decap_8 FILLER_4_3469 ();
 sg13g2_decap_8 FILLER_4_3476 ();
 sg13g2_decap_8 FILLER_4_3483 ();
 sg13g2_decap_8 FILLER_4_3490 ();
 sg13g2_decap_8 FILLER_4_3497 ();
 sg13g2_decap_8 FILLER_4_3504 ();
 sg13g2_decap_8 FILLER_4_3511 ();
 sg13g2_decap_8 FILLER_4_3518 ();
 sg13g2_decap_8 FILLER_4_3525 ();
 sg13g2_decap_8 FILLER_4_3532 ();
 sg13g2_decap_8 FILLER_4_3539 ();
 sg13g2_decap_8 FILLER_4_3546 ();
 sg13g2_decap_8 FILLER_4_3553 ();
 sg13g2_decap_8 FILLER_4_3560 ();
 sg13g2_decap_8 FILLER_4_3567 ();
 sg13g2_decap_4 FILLER_4_3574 ();
 sg13g2_fill_2 FILLER_4_3578 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_4 FILLER_5_70 ();
 sg13g2_fill_1 FILLER_5_83 ();
 sg13g2_decap_8 FILLER_5_94 ();
 sg13g2_decap_8 FILLER_5_101 ();
 sg13g2_fill_2 FILLER_5_116 ();
 sg13g2_fill_1 FILLER_5_118 ();
 sg13g2_decap_8 FILLER_5_135 ();
 sg13g2_decap_8 FILLER_5_142 ();
 sg13g2_decap_8 FILLER_5_149 ();
 sg13g2_decap_8 FILLER_5_156 ();
 sg13g2_decap_8 FILLER_5_163 ();
 sg13g2_decap_4 FILLER_5_170 ();
 sg13g2_decap_4 FILLER_5_179 ();
 sg13g2_fill_1 FILLER_5_183 ();
 sg13g2_fill_2 FILLER_5_188 ();
 sg13g2_fill_1 FILLER_5_208 ();
 sg13g2_decap_8 FILLER_5_218 ();
 sg13g2_decap_8 FILLER_5_225 ();
 sg13g2_decap_8 FILLER_5_232 ();
 sg13g2_decap_8 FILLER_5_239 ();
 sg13g2_fill_2 FILLER_5_246 ();
 sg13g2_fill_1 FILLER_5_248 ();
 sg13g2_decap_4 FILLER_5_259 ();
 sg13g2_fill_1 FILLER_5_263 ();
 sg13g2_decap_8 FILLER_5_272 ();
 sg13g2_decap_8 FILLER_5_310 ();
 sg13g2_decap_8 FILLER_5_317 ();
 sg13g2_decap_8 FILLER_5_324 ();
 sg13g2_decap_8 FILLER_5_331 ();
 sg13g2_decap_8 FILLER_5_338 ();
 sg13g2_decap_8 FILLER_5_345 ();
 sg13g2_decap_4 FILLER_5_352 ();
 sg13g2_decap_8 FILLER_5_366 ();
 sg13g2_decap_8 FILLER_5_373 ();
 sg13g2_decap_8 FILLER_5_380 ();
 sg13g2_decap_8 FILLER_5_387 ();
 sg13g2_decap_8 FILLER_5_394 ();
 sg13g2_decap_8 FILLER_5_401 ();
 sg13g2_decap_8 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_5_415 ();
 sg13g2_decap_8 FILLER_5_422 ();
 sg13g2_fill_2 FILLER_5_429 ();
 sg13g2_fill_1 FILLER_5_431 ();
 sg13g2_decap_8 FILLER_5_500 ();
 sg13g2_decap_8 FILLER_5_507 ();
 sg13g2_decap_8 FILLER_5_514 ();
 sg13g2_fill_2 FILLER_5_521 ();
 sg13g2_decap_8 FILLER_5_538 ();
 sg13g2_decap_8 FILLER_5_545 ();
 sg13g2_decap_8 FILLER_5_552 ();
 sg13g2_fill_1 FILLER_5_559 ();
 sg13g2_decap_8 FILLER_5_579 ();
 sg13g2_decap_8 FILLER_5_586 ();
 sg13g2_decap_8 FILLER_5_593 ();
 sg13g2_decap_4 FILLER_5_600 ();
 sg13g2_fill_2 FILLER_5_604 ();
 sg13g2_decap_8 FILLER_5_627 ();
 sg13g2_decap_8 FILLER_5_634 ();
 sg13g2_decap_8 FILLER_5_641 ();
 sg13g2_fill_1 FILLER_5_648 ();
 sg13g2_decap_8 FILLER_5_653 ();
 sg13g2_decap_8 FILLER_5_660 ();
 sg13g2_decap_4 FILLER_5_667 ();
 sg13g2_fill_1 FILLER_5_671 ();
 sg13g2_fill_1 FILLER_5_702 ();
 sg13g2_decap_8 FILLER_5_708 ();
 sg13g2_decap_8 FILLER_5_715 ();
 sg13g2_fill_2 FILLER_5_722 ();
 sg13g2_fill_1 FILLER_5_724 ();
 sg13g2_decap_8 FILLER_5_746 ();
 sg13g2_decap_8 FILLER_5_753 ();
 sg13g2_decap_8 FILLER_5_760 ();
 sg13g2_decap_8 FILLER_5_767 ();
 sg13g2_decap_4 FILLER_5_774 ();
 sg13g2_decap_8 FILLER_5_788 ();
 sg13g2_decap_8 FILLER_5_795 ();
 sg13g2_decap_8 FILLER_5_802 ();
 sg13g2_decap_8 FILLER_5_809 ();
 sg13g2_decap_8 FILLER_5_816 ();
 sg13g2_decap_8 FILLER_5_823 ();
 sg13g2_fill_2 FILLER_5_830 ();
 sg13g2_fill_1 FILLER_5_832 ();
 sg13g2_decap_8 FILLER_5_859 ();
 sg13g2_decap_8 FILLER_5_866 ();
 sg13g2_fill_2 FILLER_5_873 ();
 sg13g2_fill_1 FILLER_5_896 ();
 sg13g2_fill_1 FILLER_5_922 ();
 sg13g2_decap_8 FILLER_5_928 ();
 sg13g2_decap_8 FILLER_5_935 ();
 sg13g2_decap_8 FILLER_5_942 ();
 sg13g2_decap_8 FILLER_5_949 ();
 sg13g2_decap_8 FILLER_5_956 ();
 sg13g2_decap_4 FILLER_5_963 ();
 sg13g2_decap_8 FILLER_5_993 ();
 sg13g2_decap_8 FILLER_5_1000 ();
 sg13g2_fill_2 FILLER_5_1007 ();
 sg13g2_decap_8 FILLER_5_1035 ();
 sg13g2_decap_8 FILLER_5_1042 ();
 sg13g2_fill_2 FILLER_5_1049 ();
 sg13g2_decap_8 FILLER_5_1054 ();
 sg13g2_decap_8 FILLER_5_1061 ();
 sg13g2_decap_4 FILLER_5_1068 ();
 sg13g2_fill_1 FILLER_5_1072 ();
 sg13g2_fill_2 FILLER_5_1076 ();
 sg13g2_fill_2 FILLER_5_1081 ();
 sg13g2_decap_8 FILLER_5_1096 ();
 sg13g2_decap_8 FILLER_5_1103 ();
 sg13g2_decap_8 FILLER_5_1110 ();
 sg13g2_decap_8 FILLER_5_1117 ();
 sg13g2_decap_8 FILLER_5_1124 ();
 sg13g2_decap_8 FILLER_5_1131 ();
 sg13g2_decap_8 FILLER_5_1138 ();
 sg13g2_decap_8 FILLER_5_1145 ();
 sg13g2_decap_8 FILLER_5_1152 ();
 sg13g2_decap_8 FILLER_5_1159 ();
 sg13g2_decap_8 FILLER_5_1166 ();
 sg13g2_decap_8 FILLER_5_1173 ();
 sg13g2_decap_4 FILLER_5_1180 ();
 sg13g2_fill_1 FILLER_5_1184 ();
 sg13g2_decap_4 FILLER_5_1193 ();
 sg13g2_fill_2 FILLER_5_1197 ();
 sg13g2_decap_8 FILLER_5_1209 ();
 sg13g2_decap_8 FILLER_5_1216 ();
 sg13g2_decap_8 FILLER_5_1223 ();
 sg13g2_decap_4 FILLER_5_1230 ();
 sg13g2_decap_8 FILLER_5_1239 ();
 sg13g2_decap_8 FILLER_5_1273 ();
 sg13g2_decap_8 FILLER_5_1280 ();
 sg13g2_decap_8 FILLER_5_1287 ();
 sg13g2_decap_8 FILLER_5_1294 ();
 sg13g2_decap_8 FILLER_5_1301 ();
 sg13g2_decap_8 FILLER_5_1308 ();
 sg13g2_decap_8 FILLER_5_1315 ();
 sg13g2_decap_8 FILLER_5_1322 ();
 sg13g2_decap_8 FILLER_5_1329 ();
 sg13g2_fill_2 FILLER_5_1336 ();
 sg13g2_decap_4 FILLER_5_1348 ();
 sg13g2_decap_8 FILLER_5_1378 ();
 sg13g2_decap_8 FILLER_5_1385 ();
 sg13g2_decap_8 FILLER_5_1392 ();
 sg13g2_fill_1 FILLER_5_1399 ();
 sg13g2_fill_2 FILLER_5_1410 ();
 sg13g2_fill_1 FILLER_5_1412 ();
 sg13g2_decap_8 FILLER_5_1423 ();
 sg13g2_decap_8 FILLER_5_1430 ();
 sg13g2_decap_8 FILLER_5_1437 ();
 sg13g2_decap_8 FILLER_5_1444 ();
 sg13g2_decap_8 FILLER_5_1451 ();
 sg13g2_decap_4 FILLER_5_1458 ();
 sg13g2_fill_2 FILLER_5_1462 ();
 sg13g2_decap_8 FILLER_5_1477 ();
 sg13g2_decap_8 FILLER_5_1484 ();
 sg13g2_decap_8 FILLER_5_1491 ();
 sg13g2_decap_4 FILLER_5_1498 ();
 sg13g2_decap_8 FILLER_5_1512 ();
 sg13g2_decap_8 FILLER_5_1519 ();
 sg13g2_decap_8 FILLER_5_1526 ();
 sg13g2_decap_8 FILLER_5_1533 ();
 sg13g2_decap_8 FILLER_5_1540 ();
 sg13g2_decap_8 FILLER_5_1547 ();
 sg13g2_decap_8 FILLER_5_1554 ();
 sg13g2_decap_8 FILLER_5_1561 ();
 sg13g2_decap_4 FILLER_5_1568 ();
 sg13g2_fill_2 FILLER_5_1572 ();
 sg13g2_decap_8 FILLER_5_1595 ();
 sg13g2_decap_8 FILLER_5_1602 ();
 sg13g2_decap_4 FILLER_5_1609 ();
 sg13g2_fill_2 FILLER_5_1621 ();
 sg13g2_fill_1 FILLER_5_1623 ();
 sg13g2_decap_8 FILLER_5_1629 ();
 sg13g2_decap_8 FILLER_5_1636 ();
 sg13g2_decap_8 FILLER_5_1648 ();
 sg13g2_fill_2 FILLER_5_1655 ();
 sg13g2_decap_8 FILLER_5_1666 ();
 sg13g2_decap_8 FILLER_5_1673 ();
 sg13g2_decap_8 FILLER_5_1680 ();
 sg13g2_decap_8 FILLER_5_1687 ();
 sg13g2_decap_4 FILLER_5_1694 ();
 sg13g2_decap_8 FILLER_5_1724 ();
 sg13g2_decap_8 FILLER_5_1731 ();
 sg13g2_decap_8 FILLER_5_1738 ();
 sg13g2_decap_8 FILLER_5_1745 ();
 sg13g2_decap_8 FILLER_5_1752 ();
 sg13g2_decap_8 FILLER_5_1759 ();
 sg13g2_decap_8 FILLER_5_1766 ();
 sg13g2_decap_8 FILLER_5_1773 ();
 sg13g2_decap_8 FILLER_5_1780 ();
 sg13g2_decap_8 FILLER_5_1787 ();
 sg13g2_decap_8 FILLER_5_1794 ();
 sg13g2_decap_8 FILLER_5_1801 ();
 sg13g2_decap_4 FILLER_5_1808 ();
 sg13g2_fill_1 FILLER_5_1812 ();
 sg13g2_decap_8 FILLER_5_1839 ();
 sg13g2_decap_4 FILLER_5_1846 ();
 sg13g2_decap_8 FILLER_5_1860 ();
 sg13g2_decap_8 FILLER_5_1867 ();
 sg13g2_decap_8 FILLER_5_1874 ();
 sg13g2_decap_8 FILLER_5_1881 ();
 sg13g2_decap_8 FILLER_5_1888 ();
 sg13g2_decap_8 FILLER_5_1895 ();
 sg13g2_decap_8 FILLER_5_1902 ();
 sg13g2_fill_1 FILLER_5_1909 ();
 sg13g2_decap_8 FILLER_5_1915 ();
 sg13g2_decap_8 FILLER_5_1922 ();
 sg13g2_decap_8 FILLER_5_1929 ();
 sg13g2_fill_2 FILLER_5_1950 ();
 sg13g2_fill_1 FILLER_5_1952 ();
 sg13g2_fill_1 FILLER_5_1962 ();
 sg13g2_decap_8 FILLER_5_1991 ();
 sg13g2_decap_8 FILLER_5_1998 ();
 sg13g2_decap_8 FILLER_5_2005 ();
 sg13g2_decap_8 FILLER_5_2020 ();
 sg13g2_decap_8 FILLER_5_2027 ();
 sg13g2_decap_8 FILLER_5_2034 ();
 sg13g2_decap_8 FILLER_5_2041 ();
 sg13g2_decap_8 FILLER_5_2048 ();
 sg13g2_decap_8 FILLER_5_2055 ();
 sg13g2_decap_8 FILLER_5_2062 ();
 sg13g2_decap_8 FILLER_5_2069 ();
 sg13g2_fill_2 FILLER_5_2076 ();
 sg13g2_decap_8 FILLER_5_2109 ();
 sg13g2_decap_8 FILLER_5_2116 ();
 sg13g2_decap_8 FILLER_5_2123 ();
 sg13g2_decap_8 FILLER_5_2130 ();
 sg13g2_decap_8 FILLER_5_2137 ();
 sg13g2_decap_8 FILLER_5_2144 ();
 sg13g2_decap_8 FILLER_5_2151 ();
 sg13g2_fill_2 FILLER_5_2158 ();
 sg13g2_fill_1 FILLER_5_2160 ();
 sg13g2_decap_8 FILLER_5_2166 ();
 sg13g2_decap_8 FILLER_5_2173 ();
 sg13g2_decap_8 FILLER_5_2180 ();
 sg13g2_decap_8 FILLER_5_2187 ();
 sg13g2_decap_8 FILLER_5_2194 ();
 sg13g2_fill_1 FILLER_5_2201 ();
 sg13g2_decap_4 FILLER_5_2207 ();
 sg13g2_decap_8 FILLER_5_2219 ();
 sg13g2_decap_8 FILLER_5_2226 ();
 sg13g2_decap_8 FILLER_5_2233 ();
 sg13g2_decap_8 FILLER_5_2240 ();
 sg13g2_decap_8 FILLER_5_2247 ();
 sg13g2_decap_4 FILLER_5_2254 ();
 sg13g2_fill_1 FILLER_5_2258 ();
 sg13g2_decap_8 FILLER_5_2264 ();
 sg13g2_fill_2 FILLER_5_2271 ();
 sg13g2_decap_8 FILLER_5_2293 ();
 sg13g2_decap_8 FILLER_5_2300 ();
 sg13g2_decap_8 FILLER_5_2307 ();
 sg13g2_decap_8 FILLER_5_2314 ();
 sg13g2_decap_8 FILLER_5_2321 ();
 sg13g2_decap_4 FILLER_5_2328 ();
 sg13g2_decap_8 FILLER_5_2346 ();
 sg13g2_decap_8 FILLER_5_2353 ();
 sg13g2_decap_8 FILLER_5_2360 ();
 sg13g2_decap_8 FILLER_5_2367 ();
 sg13g2_decap_8 FILLER_5_2374 ();
 sg13g2_decap_8 FILLER_5_2381 ();
 sg13g2_decap_8 FILLER_5_2398 ();
 sg13g2_fill_2 FILLER_5_2405 ();
 sg13g2_fill_1 FILLER_5_2407 ();
 sg13g2_fill_2 FILLER_5_2417 ();
 sg13g2_fill_1 FILLER_5_2419 ();
 sg13g2_decap_8 FILLER_5_2429 ();
 sg13g2_decap_8 FILLER_5_2436 ();
 sg13g2_decap_8 FILLER_5_2443 ();
 sg13g2_decap_8 FILLER_5_2450 ();
 sg13g2_decap_8 FILLER_5_2457 ();
 sg13g2_decap_8 FILLER_5_2464 ();
 sg13g2_decap_4 FILLER_5_2471 ();
 sg13g2_fill_2 FILLER_5_2475 ();
 sg13g2_decap_8 FILLER_5_2482 ();
 sg13g2_decap_8 FILLER_5_2489 ();
 sg13g2_decap_8 FILLER_5_2496 ();
 sg13g2_decap_8 FILLER_5_2503 ();
 sg13g2_decap_8 FILLER_5_2510 ();
 sg13g2_decap_8 FILLER_5_2526 ();
 sg13g2_decap_8 FILLER_5_2533 ();
 sg13g2_fill_1 FILLER_5_2540 ();
 sg13g2_decap_8 FILLER_5_2546 ();
 sg13g2_decap_8 FILLER_5_2553 ();
 sg13g2_decap_8 FILLER_5_2560 ();
 sg13g2_decap_4 FILLER_5_2567 ();
 sg13g2_fill_1 FILLER_5_2571 ();
 sg13g2_decap_8 FILLER_5_2577 ();
 sg13g2_decap_4 FILLER_5_2584 ();
 sg13g2_fill_1 FILLER_5_2588 ();
 sg13g2_decap_8 FILLER_5_2594 ();
 sg13g2_decap_8 FILLER_5_2601 ();
 sg13g2_decap_8 FILLER_5_2608 ();
 sg13g2_decap_8 FILLER_5_2615 ();
 sg13g2_decap_8 FILLER_5_2622 ();
 sg13g2_decap_8 FILLER_5_2629 ();
 sg13g2_decap_8 FILLER_5_2636 ();
 sg13g2_decap_8 FILLER_5_2643 ();
 sg13g2_decap_8 FILLER_5_2650 ();
 sg13g2_decap_8 FILLER_5_2657 ();
 sg13g2_decap_8 FILLER_5_2664 ();
 sg13g2_decap_8 FILLER_5_2671 ();
 sg13g2_decap_8 FILLER_5_2678 ();
 sg13g2_decap_8 FILLER_5_2685 ();
 sg13g2_decap_4 FILLER_5_2692 ();
 sg13g2_decap_8 FILLER_5_2700 ();
 sg13g2_decap_8 FILLER_5_2707 ();
 sg13g2_fill_2 FILLER_5_2714 ();
 sg13g2_decap_8 FILLER_5_2742 ();
 sg13g2_decap_8 FILLER_5_2749 ();
 sg13g2_decap_8 FILLER_5_2756 ();
 sg13g2_decap_8 FILLER_5_2763 ();
 sg13g2_decap_8 FILLER_5_2770 ();
 sg13g2_fill_2 FILLER_5_2777 ();
 sg13g2_fill_1 FILLER_5_2779 ();
 sg13g2_decap_8 FILLER_5_2805 ();
 sg13g2_decap_8 FILLER_5_2812 ();
 sg13g2_decap_8 FILLER_5_2819 ();
 sg13g2_decap_8 FILLER_5_2826 ();
 sg13g2_fill_2 FILLER_5_2833 ();
 sg13g2_decap_8 FILLER_5_2840 ();
 sg13g2_decap_8 FILLER_5_2847 ();
 sg13g2_decap_8 FILLER_5_2854 ();
 sg13g2_fill_1 FILLER_5_2861 ();
 sg13g2_decap_8 FILLER_5_2887 ();
 sg13g2_decap_8 FILLER_5_2894 ();
 sg13g2_decap_8 FILLER_5_2901 ();
 sg13g2_decap_4 FILLER_5_2908 ();
 sg13g2_fill_1 FILLER_5_2912 ();
 sg13g2_decap_8 FILLER_5_2933 ();
 sg13g2_decap_8 FILLER_5_2966 ();
 sg13g2_decap_4 FILLER_5_2973 ();
 sg13g2_fill_2 FILLER_5_2977 ();
 sg13g2_decap_8 FILLER_5_2987 ();
 sg13g2_fill_2 FILLER_5_2994 ();
 sg13g2_decap_8 FILLER_5_3067 ();
 sg13g2_decap_4 FILLER_5_3074 ();
 sg13g2_fill_2 FILLER_5_3078 ();
 sg13g2_decap_8 FILLER_5_3085 ();
 sg13g2_fill_2 FILLER_5_3092 ();
 sg13g2_fill_1 FILLER_5_3094 ();
 sg13g2_decap_8 FILLER_5_3105 ();
 sg13g2_decap_8 FILLER_5_3112 ();
 sg13g2_decap_8 FILLER_5_3119 ();
 sg13g2_decap_8 FILLER_5_3126 ();
 sg13g2_decap_8 FILLER_5_3133 ();
 sg13g2_decap_8 FILLER_5_3140 ();
 sg13g2_decap_8 FILLER_5_3147 ();
 sg13g2_fill_2 FILLER_5_3154 ();
 sg13g2_decap_8 FILLER_5_3192 ();
 sg13g2_decap_8 FILLER_5_3199 ();
 sg13g2_decap_4 FILLER_5_3206 ();
 sg13g2_decap_8 FILLER_5_3214 ();
 sg13g2_fill_2 FILLER_5_3230 ();
 sg13g2_decap_8 FILLER_5_3242 ();
 sg13g2_decap_8 FILLER_5_3249 ();
 sg13g2_decap_8 FILLER_5_3265 ();
 sg13g2_decap_8 FILLER_5_3272 ();
 sg13g2_decap_8 FILLER_5_3279 ();
 sg13g2_decap_8 FILLER_5_3286 ();
 sg13g2_decap_8 FILLER_5_3293 ();
 sg13g2_decap_8 FILLER_5_3300 ();
 sg13g2_decap_8 FILLER_5_3307 ();
 sg13g2_decap_8 FILLER_5_3314 ();
 sg13g2_decap_8 FILLER_5_3321 ();
 sg13g2_decap_8 FILLER_5_3328 ();
 sg13g2_decap_8 FILLER_5_3335 ();
 sg13g2_decap_8 FILLER_5_3342 ();
 sg13g2_decap_8 FILLER_5_3349 ();
 sg13g2_decap_8 FILLER_5_3356 ();
 sg13g2_decap_8 FILLER_5_3363 ();
 sg13g2_decap_8 FILLER_5_3370 ();
 sg13g2_decap_8 FILLER_5_3377 ();
 sg13g2_decap_8 FILLER_5_3384 ();
 sg13g2_decap_8 FILLER_5_3391 ();
 sg13g2_decap_8 FILLER_5_3398 ();
 sg13g2_decap_8 FILLER_5_3405 ();
 sg13g2_decap_8 FILLER_5_3412 ();
 sg13g2_decap_8 FILLER_5_3419 ();
 sg13g2_decap_8 FILLER_5_3426 ();
 sg13g2_decap_8 FILLER_5_3433 ();
 sg13g2_decap_8 FILLER_5_3440 ();
 sg13g2_decap_8 FILLER_5_3447 ();
 sg13g2_decap_8 FILLER_5_3454 ();
 sg13g2_decap_8 FILLER_5_3461 ();
 sg13g2_decap_8 FILLER_5_3468 ();
 sg13g2_decap_8 FILLER_5_3475 ();
 sg13g2_decap_8 FILLER_5_3482 ();
 sg13g2_decap_8 FILLER_5_3489 ();
 sg13g2_decap_8 FILLER_5_3496 ();
 sg13g2_decap_8 FILLER_5_3503 ();
 sg13g2_decap_8 FILLER_5_3510 ();
 sg13g2_decap_8 FILLER_5_3517 ();
 sg13g2_decap_8 FILLER_5_3524 ();
 sg13g2_decap_8 FILLER_5_3531 ();
 sg13g2_decap_8 FILLER_5_3538 ();
 sg13g2_decap_8 FILLER_5_3545 ();
 sg13g2_decap_8 FILLER_5_3552 ();
 sg13g2_decap_8 FILLER_5_3559 ();
 sg13g2_decap_8 FILLER_5_3566 ();
 sg13g2_decap_8 FILLER_5_3573 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_4 FILLER_6_63 ();
 sg13g2_fill_1 FILLER_6_67 ();
 sg13g2_decap_8 FILLER_6_135 ();
 sg13g2_decap_8 FILLER_6_142 ();
 sg13g2_decap_8 FILLER_6_149 ();
 sg13g2_decap_8 FILLER_6_156 ();
 sg13g2_decap_8 FILLER_6_163 ();
 sg13g2_decap_8 FILLER_6_170 ();
 sg13g2_decap_8 FILLER_6_177 ();
 sg13g2_decap_4 FILLER_6_184 ();
 sg13g2_fill_2 FILLER_6_188 ();
 sg13g2_decap_8 FILLER_6_221 ();
 sg13g2_decap_8 FILLER_6_228 ();
 sg13g2_decap_8 FILLER_6_235 ();
 sg13g2_decap_8 FILLER_6_242 ();
 sg13g2_decap_8 FILLER_6_249 ();
 sg13g2_decap_8 FILLER_6_256 ();
 sg13g2_decap_8 FILLER_6_263 ();
 sg13g2_decap_8 FILLER_6_270 ();
 sg13g2_fill_2 FILLER_6_281 ();
 sg13g2_fill_1 FILLER_6_283 ();
 sg13g2_decap_8 FILLER_6_292 ();
 sg13g2_decap_8 FILLER_6_299 ();
 sg13g2_decap_8 FILLER_6_306 ();
 sg13g2_decap_8 FILLER_6_313 ();
 sg13g2_decap_8 FILLER_6_320 ();
 sg13g2_decap_8 FILLER_6_327 ();
 sg13g2_decap_8 FILLER_6_334 ();
 sg13g2_decap_8 FILLER_6_341 ();
 sg13g2_decap_8 FILLER_6_348 ();
 sg13g2_decap_8 FILLER_6_355 ();
 sg13g2_decap_8 FILLER_6_362 ();
 sg13g2_decap_8 FILLER_6_369 ();
 sg13g2_decap_8 FILLER_6_376 ();
 sg13g2_decap_8 FILLER_6_383 ();
 sg13g2_decap_8 FILLER_6_390 ();
 sg13g2_decap_8 FILLER_6_397 ();
 sg13g2_decap_8 FILLER_6_404 ();
 sg13g2_decap_8 FILLER_6_411 ();
 sg13g2_decap_8 FILLER_6_418 ();
 sg13g2_decap_8 FILLER_6_425 ();
 sg13g2_decap_8 FILLER_6_432 ();
 sg13g2_decap_8 FILLER_6_439 ();
 sg13g2_decap_8 FILLER_6_446 ();
 sg13g2_decap_8 FILLER_6_453 ();
 sg13g2_decap_4 FILLER_6_460 ();
 sg13g2_fill_1 FILLER_6_464 ();
 sg13g2_decap_4 FILLER_6_479 ();
 sg13g2_fill_1 FILLER_6_483 ();
 sg13g2_decap_8 FILLER_6_493 ();
 sg13g2_decap_8 FILLER_6_500 ();
 sg13g2_decap_8 FILLER_6_507 ();
 sg13g2_decap_8 FILLER_6_514 ();
 sg13g2_decap_8 FILLER_6_521 ();
 sg13g2_decap_8 FILLER_6_528 ();
 sg13g2_decap_8 FILLER_6_535 ();
 sg13g2_decap_8 FILLER_6_542 ();
 sg13g2_decap_8 FILLER_6_549 ();
 sg13g2_decap_8 FILLER_6_556 ();
 sg13g2_fill_2 FILLER_6_563 ();
 sg13g2_fill_1 FILLER_6_570 ();
 sg13g2_decap_8 FILLER_6_581 ();
 sg13g2_decap_8 FILLER_6_588 ();
 sg13g2_decap_8 FILLER_6_595 ();
 sg13g2_decap_8 FILLER_6_602 ();
 sg13g2_decap_8 FILLER_6_609 ();
 sg13g2_decap_8 FILLER_6_616 ();
 sg13g2_decap_8 FILLER_6_623 ();
 sg13g2_fill_1 FILLER_6_630 ();
 sg13g2_fill_2 FILLER_6_636 ();
 sg13g2_fill_1 FILLER_6_638 ();
 sg13g2_decap_8 FILLER_6_674 ();
 sg13g2_decap_4 FILLER_6_681 ();
 sg13g2_fill_1 FILLER_6_685 ();
 sg13g2_decap_8 FILLER_6_695 ();
 sg13g2_decap_8 FILLER_6_702 ();
 sg13g2_decap_8 FILLER_6_709 ();
 sg13g2_decap_8 FILLER_6_716 ();
 sg13g2_decap_8 FILLER_6_723 ();
 sg13g2_decap_4 FILLER_6_730 ();
 sg13g2_fill_2 FILLER_6_734 ();
 sg13g2_fill_2 FILLER_6_741 ();
 sg13g2_decap_8 FILLER_6_748 ();
 sg13g2_decap_8 FILLER_6_755 ();
 sg13g2_decap_4 FILLER_6_762 ();
 sg13g2_fill_2 FILLER_6_766 ();
 sg13g2_decap_8 FILLER_6_798 ();
 sg13g2_decap_8 FILLER_6_805 ();
 sg13g2_decap_8 FILLER_6_812 ();
 sg13g2_decap_8 FILLER_6_863 ();
 sg13g2_decap_8 FILLER_6_870 ();
 sg13g2_fill_2 FILLER_6_877 ();
 sg13g2_fill_1 FILLER_6_884 ();
 sg13g2_decap_8 FILLER_6_890 ();
 sg13g2_fill_2 FILLER_6_897 ();
 sg13g2_decap_8 FILLER_6_904 ();
 sg13g2_decap_8 FILLER_6_911 ();
 sg13g2_decap_8 FILLER_6_922 ();
 sg13g2_decap_8 FILLER_6_929 ();
 sg13g2_decap_8 FILLER_6_936 ();
 sg13g2_decap_8 FILLER_6_943 ();
 sg13g2_fill_2 FILLER_6_950 ();
 sg13g2_fill_1 FILLER_6_952 ();
 sg13g2_decap_8 FILLER_6_958 ();
 sg13g2_decap_8 FILLER_6_965 ();
 sg13g2_fill_1 FILLER_6_972 ();
 sg13g2_decap_8 FILLER_6_991 ();
 sg13g2_fill_1 FILLER_6_1001 ();
 sg13g2_decap_8 FILLER_6_1022 ();
 sg13g2_decap_8 FILLER_6_1029 ();
 sg13g2_decap_8 FILLER_6_1036 ();
 sg13g2_fill_1 FILLER_6_1043 ();
 sg13g2_decap_4 FILLER_6_1047 ();
 sg13g2_decap_8 FILLER_6_1061 ();
 sg13g2_decap_4 FILLER_6_1068 ();
 sg13g2_fill_1 FILLER_6_1072 ();
 sg13g2_decap_8 FILLER_6_1103 ();
 sg13g2_decap_8 FILLER_6_1110 ();
 sg13g2_decap_8 FILLER_6_1117 ();
 sg13g2_decap_8 FILLER_6_1124 ();
 sg13g2_decap_4 FILLER_6_1131 ();
 sg13g2_fill_2 FILLER_6_1135 ();
 sg13g2_decap_8 FILLER_6_1163 ();
 sg13g2_decap_8 FILLER_6_1170 ();
 sg13g2_decap_8 FILLER_6_1177 ();
 sg13g2_decap_4 FILLER_6_1184 ();
 sg13g2_decap_8 FILLER_6_1217 ();
 sg13g2_decap_8 FILLER_6_1224 ();
 sg13g2_decap_8 FILLER_6_1231 ();
 sg13g2_decap_8 FILLER_6_1238 ();
 sg13g2_fill_1 FILLER_6_1245 ();
 sg13g2_fill_1 FILLER_6_1272 ();
 sg13g2_decap_8 FILLER_6_1281 ();
 sg13g2_decap_8 FILLER_6_1288 ();
 sg13g2_decap_8 FILLER_6_1295 ();
 sg13g2_decap_4 FILLER_6_1302 ();
 sg13g2_fill_2 FILLER_6_1306 ();
 sg13g2_decap_8 FILLER_6_1313 ();
 sg13g2_decap_8 FILLER_6_1320 ();
 sg13g2_decap_8 FILLER_6_1327 ();
 sg13g2_decap_4 FILLER_6_1334 ();
 sg13g2_fill_1 FILLER_6_1338 ();
 sg13g2_fill_1 FILLER_6_1349 ();
 sg13g2_decap_8 FILLER_6_1376 ();
 sg13g2_decap_8 FILLER_6_1383 ();
 sg13g2_decap_8 FILLER_6_1390 ();
 sg13g2_decap_8 FILLER_6_1397 ();
 sg13g2_decap_8 FILLER_6_1404 ();
 sg13g2_fill_1 FILLER_6_1411 ();
 sg13g2_decap_8 FILLER_6_1422 ();
 sg13g2_decap_8 FILLER_6_1429 ();
 sg13g2_decap_8 FILLER_6_1436 ();
 sg13g2_decap_8 FILLER_6_1443 ();
 sg13g2_decap_8 FILLER_6_1450 ();
 sg13g2_decap_8 FILLER_6_1457 ();
 sg13g2_decap_8 FILLER_6_1464 ();
 sg13g2_decap_8 FILLER_6_1471 ();
 sg13g2_decap_8 FILLER_6_1478 ();
 sg13g2_decap_8 FILLER_6_1485 ();
 sg13g2_decap_4 FILLER_6_1492 ();
 sg13g2_fill_2 FILLER_6_1496 ();
 sg13g2_decap_8 FILLER_6_1534 ();
 sg13g2_decap_8 FILLER_6_1541 ();
 sg13g2_decap_8 FILLER_6_1548 ();
 sg13g2_decap_4 FILLER_6_1555 ();
 sg13g2_fill_2 FILLER_6_1559 ();
 sg13g2_decap_8 FILLER_6_1587 ();
 sg13g2_decap_8 FILLER_6_1594 ();
 sg13g2_decap_8 FILLER_6_1601 ();
 sg13g2_decap_8 FILLER_6_1608 ();
 sg13g2_decap_8 FILLER_6_1615 ();
 sg13g2_decap_8 FILLER_6_1638 ();
 sg13g2_decap_8 FILLER_6_1645 ();
 sg13g2_fill_2 FILLER_6_1652 ();
 sg13g2_decap_8 FILLER_6_1680 ();
 sg13g2_decap_8 FILLER_6_1687 ();
 sg13g2_decap_8 FILLER_6_1694 ();
 sg13g2_decap_8 FILLER_6_1701 ();
 sg13g2_decap_8 FILLER_6_1708 ();
 sg13g2_fill_1 FILLER_6_1715 ();
 sg13g2_fill_2 FILLER_6_1731 ();
 sg13g2_fill_1 FILLER_6_1733 ();
 sg13g2_fill_1 FILLER_6_1750 ();
 sg13g2_decap_4 FILLER_6_1761 ();
 sg13g2_fill_1 FILLER_6_1765 ();
 sg13g2_decap_8 FILLER_6_1771 ();
 sg13g2_decap_8 FILLER_6_1778 ();
 sg13g2_decap_4 FILLER_6_1795 ();
 sg13g2_fill_1 FILLER_6_1799 ();
 sg13g2_decap_4 FILLER_6_1810 ();
 sg13g2_fill_2 FILLER_6_1814 ();
 sg13g2_decap_8 FILLER_6_1826 ();
 sg13g2_decap_8 FILLER_6_1833 ();
 sg13g2_decap_8 FILLER_6_1840 ();
 sg13g2_fill_2 FILLER_6_1847 ();
 sg13g2_fill_1 FILLER_6_1849 ();
 sg13g2_fill_2 FILLER_6_1860 ();
 sg13g2_fill_1 FILLER_6_1862 ();
 sg13g2_decap_8 FILLER_6_1871 ();
 sg13g2_decap_4 FILLER_6_1878 ();
 sg13g2_fill_2 FILLER_6_1882 ();
 sg13g2_decap_8 FILLER_6_1894 ();
 sg13g2_decap_8 FILLER_6_1916 ();
 sg13g2_decap_8 FILLER_6_1923 ();
 sg13g2_decap_8 FILLER_6_1930 ();
 sg13g2_decap_4 FILLER_6_1937 ();
 sg13g2_decap_8 FILLER_6_1945 ();
 sg13g2_decap_8 FILLER_6_1952 ();
 sg13g2_decap_8 FILLER_6_1959 ();
 sg13g2_decap_8 FILLER_6_1966 ();
 sg13g2_decap_8 FILLER_6_1973 ();
 sg13g2_decap_8 FILLER_6_1980 ();
 sg13g2_decap_8 FILLER_6_1987 ();
 sg13g2_decap_8 FILLER_6_1994 ();
 sg13g2_decap_8 FILLER_6_2001 ();
 sg13g2_decap_8 FILLER_6_2008 ();
 sg13g2_decap_8 FILLER_6_2015 ();
 sg13g2_decap_8 FILLER_6_2022 ();
 sg13g2_decap_8 FILLER_6_2029 ();
 sg13g2_decap_8 FILLER_6_2036 ();
 sg13g2_decap_8 FILLER_6_2043 ();
 sg13g2_decap_8 FILLER_6_2050 ();
 sg13g2_decap_8 FILLER_6_2057 ();
 sg13g2_decap_8 FILLER_6_2064 ();
 sg13g2_decap_8 FILLER_6_2071 ();
 sg13g2_decap_8 FILLER_6_2078 ();
 sg13g2_fill_1 FILLER_6_2085 ();
 sg13g2_decap_4 FILLER_6_2104 ();
 sg13g2_decap_8 FILLER_6_2118 ();
 sg13g2_fill_2 FILLER_6_2125 ();
 sg13g2_fill_1 FILLER_6_2127 ();
 sg13g2_fill_1 FILLER_6_2143 ();
 sg13g2_decap_8 FILLER_6_2149 ();
 sg13g2_decap_8 FILLER_6_2156 ();
 sg13g2_fill_1 FILLER_6_2163 ();
 sg13g2_decap_8 FILLER_6_2179 ();
 sg13g2_decap_8 FILLER_6_2186 ();
 sg13g2_decap_8 FILLER_6_2193 ();
 sg13g2_decap_4 FILLER_6_2200 ();
 sg13g2_fill_2 FILLER_6_2204 ();
 sg13g2_decap_8 FILLER_6_2221 ();
 sg13g2_decap_8 FILLER_6_2228 ();
 sg13g2_decap_8 FILLER_6_2235 ();
 sg13g2_fill_1 FILLER_6_2242 ();
 sg13g2_fill_2 FILLER_6_2248 ();
 sg13g2_fill_1 FILLER_6_2250 ();
 sg13g2_decap_8 FILLER_6_2261 ();
 sg13g2_decap_8 FILLER_6_2268 ();
 sg13g2_decap_8 FILLER_6_2275 ();
 sg13g2_decap_8 FILLER_6_2287 ();
 sg13g2_decap_8 FILLER_6_2294 ();
 sg13g2_decap_4 FILLER_6_2301 ();
 sg13g2_fill_1 FILLER_6_2305 ();
 sg13g2_decap_8 FILLER_6_2311 ();
 sg13g2_decap_8 FILLER_6_2318 ();
 sg13g2_fill_2 FILLER_6_2325 ();
 sg13g2_decap_8 FILLER_6_2358 ();
 sg13g2_decap_8 FILLER_6_2365 ();
 sg13g2_decap_8 FILLER_6_2398 ();
 sg13g2_decap_8 FILLER_6_2405 ();
 sg13g2_decap_4 FILLER_6_2412 ();
 sg13g2_fill_2 FILLER_6_2416 ();
 sg13g2_fill_2 FILLER_6_2423 ();
 sg13g2_decap_8 FILLER_6_2440 ();
 sg13g2_decap_8 FILLER_6_2447 ();
 sg13g2_fill_1 FILLER_6_2454 ();
 sg13g2_decap_4 FILLER_6_2476 ();
 sg13g2_decap_8 FILLER_6_2495 ();
 sg13g2_decap_8 FILLER_6_2502 ();
 sg13g2_decap_4 FILLER_6_2509 ();
 sg13g2_fill_2 FILLER_6_2513 ();
 sg13g2_decap_8 FILLER_6_2530 ();
 sg13g2_decap_8 FILLER_6_2537 ();
 sg13g2_fill_2 FILLER_6_2544 ();
 sg13g2_fill_2 FILLER_6_2561 ();
 sg13g2_decap_8 FILLER_6_2604 ();
 sg13g2_decap_8 FILLER_6_2611 ();
 sg13g2_decap_4 FILLER_6_2618 ();
 sg13g2_decap_8 FILLER_6_2627 ();
 sg13g2_decap_8 FILLER_6_2634 ();
 sg13g2_fill_2 FILLER_6_2641 ();
 sg13g2_fill_2 FILLER_6_2647 ();
 sg13g2_fill_1 FILLER_6_2649 ();
 sg13g2_decap_8 FILLER_6_2669 ();
 sg13g2_decap_4 FILLER_6_2676 ();
 sg13g2_fill_2 FILLER_6_2684 ();
 sg13g2_fill_1 FILLER_6_2686 ();
 sg13g2_fill_1 FILLER_6_2727 ();
 sg13g2_decap_8 FILLER_6_2737 ();
 sg13g2_decap_8 FILLER_6_2744 ();
 sg13g2_decap_8 FILLER_6_2751 ();
 sg13g2_decap_8 FILLER_6_2758 ();
 sg13g2_decap_8 FILLER_6_2765 ();
 sg13g2_decap_8 FILLER_6_2812 ();
 sg13g2_decap_8 FILLER_6_2819 ();
 sg13g2_decap_8 FILLER_6_2826 ();
 sg13g2_decap_4 FILLER_6_2843 ();
 sg13g2_decap_8 FILLER_6_2852 ();
 sg13g2_decap_8 FILLER_6_2859 ();
 sg13g2_fill_2 FILLER_6_2866 ();
 sg13g2_fill_2 FILLER_6_2872 ();
 sg13g2_fill_1 FILLER_6_2874 ();
 sg13g2_decap_8 FILLER_6_2884 ();
 sg13g2_decap_8 FILLER_6_2891 ();
 sg13g2_decap_4 FILLER_6_2898 ();
 sg13g2_fill_1 FILLER_6_2902 ();
 sg13g2_decap_8 FILLER_6_2911 ();
 sg13g2_decap_8 FILLER_6_2918 ();
 sg13g2_decap_8 FILLER_6_2930 ();
 sg13g2_decap_8 FILLER_6_2937 ();
 sg13g2_decap_8 FILLER_6_2944 ();
 sg13g2_decap_8 FILLER_6_2951 ();
 sg13g2_decap_8 FILLER_6_2958 ();
 sg13g2_decap_8 FILLER_6_2965 ();
 sg13g2_decap_8 FILLER_6_2972 ();
 sg13g2_decap_8 FILLER_6_2979 ();
 sg13g2_decap_8 FILLER_6_2986 ();
 sg13g2_decap_8 FILLER_6_2993 ();
 sg13g2_decap_8 FILLER_6_3000 ();
 sg13g2_decap_8 FILLER_6_3007 ();
 sg13g2_decap_8 FILLER_6_3014 ();
 sg13g2_decap_4 FILLER_6_3021 ();
 sg13g2_decap_4 FILLER_6_3031 ();
 sg13g2_fill_1 FILLER_6_3035 ();
 sg13g2_decap_8 FILLER_6_3052 ();
 sg13g2_decap_8 FILLER_6_3059 ();
 sg13g2_decap_8 FILLER_6_3066 ();
 sg13g2_decap_8 FILLER_6_3073 ();
 sg13g2_decap_8 FILLER_6_3080 ();
 sg13g2_decap_8 FILLER_6_3087 ();
 sg13g2_decap_8 FILLER_6_3094 ();
 sg13g2_decap_4 FILLER_6_3101 ();
 sg13g2_fill_1 FILLER_6_3105 ();
 sg13g2_decap_8 FILLER_6_3132 ();
 sg13g2_decap_4 FILLER_6_3139 ();
 sg13g2_decap_8 FILLER_6_3153 ();
 sg13g2_decap_8 FILLER_6_3160 ();
 sg13g2_decap_8 FILLER_6_3172 ();
 sg13g2_decap_8 FILLER_6_3179 ();
 sg13g2_decap_8 FILLER_6_3186 ();
 sg13g2_decap_8 FILLER_6_3193 ();
 sg13g2_decap_8 FILLER_6_3200 ();
 sg13g2_decap_4 FILLER_6_3207 ();
 sg13g2_fill_2 FILLER_6_3216 ();
 sg13g2_fill_2 FILLER_6_3222 ();
 sg13g2_decap_4 FILLER_6_3276 ();
 sg13g2_decap_8 FILLER_6_3306 ();
 sg13g2_decap_8 FILLER_6_3313 ();
 sg13g2_decap_8 FILLER_6_3320 ();
 sg13g2_decap_8 FILLER_6_3327 ();
 sg13g2_decap_8 FILLER_6_3334 ();
 sg13g2_decap_8 FILLER_6_3341 ();
 sg13g2_decap_8 FILLER_6_3348 ();
 sg13g2_decap_8 FILLER_6_3355 ();
 sg13g2_decap_8 FILLER_6_3362 ();
 sg13g2_decap_8 FILLER_6_3369 ();
 sg13g2_decap_8 FILLER_6_3376 ();
 sg13g2_decap_8 FILLER_6_3383 ();
 sg13g2_decap_8 FILLER_6_3390 ();
 sg13g2_decap_8 FILLER_6_3397 ();
 sg13g2_decap_8 FILLER_6_3404 ();
 sg13g2_decap_8 FILLER_6_3411 ();
 sg13g2_decap_8 FILLER_6_3418 ();
 sg13g2_decap_8 FILLER_6_3425 ();
 sg13g2_decap_8 FILLER_6_3432 ();
 sg13g2_decap_8 FILLER_6_3439 ();
 sg13g2_decap_8 FILLER_6_3446 ();
 sg13g2_decap_8 FILLER_6_3453 ();
 sg13g2_decap_8 FILLER_6_3460 ();
 sg13g2_decap_8 FILLER_6_3467 ();
 sg13g2_decap_8 FILLER_6_3474 ();
 sg13g2_decap_8 FILLER_6_3481 ();
 sg13g2_decap_8 FILLER_6_3488 ();
 sg13g2_decap_8 FILLER_6_3495 ();
 sg13g2_decap_8 FILLER_6_3502 ();
 sg13g2_decap_8 FILLER_6_3509 ();
 sg13g2_decap_8 FILLER_6_3516 ();
 sg13g2_decap_8 FILLER_6_3523 ();
 sg13g2_decap_8 FILLER_6_3530 ();
 sg13g2_decap_8 FILLER_6_3537 ();
 sg13g2_decap_8 FILLER_6_3544 ();
 sg13g2_decap_8 FILLER_6_3551 ();
 sg13g2_decap_8 FILLER_6_3558 ();
 sg13g2_decap_8 FILLER_6_3565 ();
 sg13g2_decap_8 FILLER_6_3572 ();
 sg13g2_fill_1 FILLER_6_3579 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_fill_2 FILLER_7_77 ();
 sg13g2_fill_1 FILLER_7_79 ();
 sg13g2_fill_2 FILLER_7_88 ();
 sg13g2_fill_1 FILLER_7_90 ();
 sg13g2_decap_8 FILLER_7_100 ();
 sg13g2_fill_1 FILLER_7_107 ();
 sg13g2_fill_1 FILLER_7_117 ();
 sg13g2_decap_8 FILLER_7_123 ();
 sg13g2_fill_2 FILLER_7_130 ();
 sg13g2_decap_4 FILLER_7_137 ();
 sg13g2_decap_8 FILLER_7_149 ();
 sg13g2_decap_8 FILLER_7_156 ();
 sg13g2_decap_8 FILLER_7_163 ();
 sg13g2_decap_8 FILLER_7_170 ();
 sg13g2_decap_8 FILLER_7_177 ();
 sg13g2_fill_1 FILLER_7_184 ();
 sg13g2_decap_8 FILLER_7_190 ();
 sg13g2_fill_1 FILLER_7_197 ();
 sg13g2_decap_8 FILLER_7_213 ();
 sg13g2_decap_8 FILLER_7_220 ();
 sg13g2_fill_2 FILLER_7_227 ();
 sg13g2_fill_1 FILLER_7_229 ();
 sg13g2_decap_8 FILLER_7_256 ();
 sg13g2_decap_8 FILLER_7_263 ();
 sg13g2_decap_8 FILLER_7_270 ();
 sg13g2_decap_4 FILLER_7_277 ();
 sg13g2_fill_1 FILLER_7_281 ();
 sg13g2_decap_4 FILLER_7_287 ();
 sg13g2_fill_2 FILLER_7_291 ();
 sg13g2_decap_8 FILLER_7_298 ();
 sg13g2_decap_8 FILLER_7_305 ();
 sg13g2_decap_8 FILLER_7_312 ();
 sg13g2_decap_8 FILLER_7_319 ();
 sg13g2_decap_8 FILLER_7_326 ();
 sg13g2_decap_4 FILLER_7_333 ();
 sg13g2_fill_1 FILLER_7_337 ();
 sg13g2_decap_4 FILLER_7_342 ();
 sg13g2_decap_8 FILLER_7_351 ();
 sg13g2_decap_8 FILLER_7_358 ();
 sg13g2_decap_8 FILLER_7_365 ();
 sg13g2_decap_8 FILLER_7_372 ();
 sg13g2_decap_4 FILLER_7_379 ();
 sg13g2_fill_2 FILLER_7_383 ();
 sg13g2_fill_1 FILLER_7_390 ();
 sg13g2_decap_8 FILLER_7_407 ();
 sg13g2_decap_8 FILLER_7_414 ();
 sg13g2_fill_1 FILLER_7_421 ();
 sg13g2_decap_8 FILLER_7_426 ();
 sg13g2_decap_8 FILLER_7_433 ();
 sg13g2_fill_2 FILLER_7_440 ();
 sg13g2_decap_8 FILLER_7_455 ();
 sg13g2_decap_8 FILLER_7_462 ();
 sg13g2_decap_8 FILLER_7_469 ();
 sg13g2_decap_8 FILLER_7_476 ();
 sg13g2_decap_8 FILLER_7_483 ();
 sg13g2_decap_8 FILLER_7_490 ();
 sg13g2_decap_8 FILLER_7_497 ();
 sg13g2_decap_8 FILLER_7_504 ();
 sg13g2_decap_4 FILLER_7_511 ();
 sg13g2_decap_8 FILLER_7_530 ();
 sg13g2_decap_8 FILLER_7_537 ();
 sg13g2_decap_8 FILLER_7_544 ();
 sg13g2_decap_8 FILLER_7_551 ();
 sg13g2_decap_4 FILLER_7_558 ();
 sg13g2_fill_1 FILLER_7_562 ();
 sg13g2_decap_8 FILLER_7_589 ();
 sg13g2_decap_8 FILLER_7_596 ();
 sg13g2_decap_8 FILLER_7_603 ();
 sg13g2_decap_8 FILLER_7_610 ();
 sg13g2_decap_8 FILLER_7_617 ();
 sg13g2_fill_2 FILLER_7_629 ();
 sg13g2_fill_2 FILLER_7_636 ();
 sg13g2_decap_8 FILLER_7_643 ();
 sg13g2_decap_8 FILLER_7_650 ();
 sg13g2_decap_8 FILLER_7_657 ();
 sg13g2_decap_8 FILLER_7_664 ();
 sg13g2_fill_2 FILLER_7_697 ();
 sg13g2_decap_8 FILLER_7_704 ();
 sg13g2_decap_8 FILLER_7_711 ();
 sg13g2_decap_8 FILLER_7_718 ();
 sg13g2_decap_8 FILLER_7_725 ();
 sg13g2_decap_8 FILLER_7_732 ();
 sg13g2_decap_4 FILLER_7_739 ();
 sg13g2_decap_8 FILLER_7_748 ();
 sg13g2_decap_8 FILLER_7_755 ();
 sg13g2_fill_2 FILLER_7_762 ();
 sg13g2_fill_1 FILLER_7_764 ();
 sg13g2_decap_8 FILLER_7_798 ();
 sg13g2_decap_8 FILLER_7_805 ();
 sg13g2_decap_8 FILLER_7_812 ();
 sg13g2_decap_8 FILLER_7_819 ();
 sg13g2_decap_4 FILLER_7_826 ();
 sg13g2_decap_8 FILLER_7_840 ();
 sg13g2_decap_8 FILLER_7_847 ();
 sg13g2_decap_8 FILLER_7_854 ();
 sg13g2_decap_8 FILLER_7_861 ();
 sg13g2_decap_8 FILLER_7_868 ();
 sg13g2_decap_8 FILLER_7_875 ();
 sg13g2_decap_8 FILLER_7_882 ();
 sg13g2_decap_8 FILLER_7_889 ();
 sg13g2_fill_2 FILLER_7_896 ();
 sg13g2_fill_1 FILLER_7_898 ();
 sg13g2_decap_8 FILLER_7_908 ();
 sg13g2_decap_8 FILLER_7_915 ();
 sg13g2_fill_2 FILLER_7_922 ();
 sg13g2_decap_8 FILLER_7_929 ();
 sg13g2_fill_2 FILLER_7_936 ();
 sg13g2_decap_4 FILLER_7_942 ();
 sg13g2_fill_1 FILLER_7_946 ();
 sg13g2_decap_8 FILLER_7_956 ();
 sg13g2_decap_8 FILLER_7_963 ();
 sg13g2_decap_8 FILLER_7_970 ();
 sg13g2_decap_8 FILLER_7_977 ();
 sg13g2_decap_8 FILLER_7_984 ();
 sg13g2_decap_4 FILLER_7_991 ();
 sg13g2_decap_8 FILLER_7_1007 ();
 sg13g2_decap_8 FILLER_7_1014 ();
 sg13g2_decap_8 FILLER_7_1021 ();
 sg13g2_decap_8 FILLER_7_1028 ();
 sg13g2_decap_8 FILLER_7_1035 ();
 sg13g2_fill_2 FILLER_7_1042 ();
 sg13g2_decap_4 FILLER_7_1075 ();
 sg13g2_decap_4 FILLER_7_1084 ();
 sg13g2_fill_2 FILLER_7_1088 ();
 sg13g2_fill_1 FILLER_7_1094 ();
 sg13g2_decap_8 FILLER_7_1112 ();
 sg13g2_decap_8 FILLER_7_1119 ();
 sg13g2_decap_4 FILLER_7_1126 ();
 sg13g2_decap_4 FILLER_7_1166 ();
 sg13g2_fill_2 FILLER_7_1170 ();
 sg13g2_decap_4 FILLER_7_1192 ();
 sg13g2_decap_8 FILLER_7_1222 ();
 sg13g2_decap_4 FILLER_7_1229 ();
 sg13g2_fill_2 FILLER_7_1233 ();
 sg13g2_decap_8 FILLER_7_1243 ();
 sg13g2_fill_2 FILLER_7_1250 ();
 sg13g2_fill_1 FILLER_7_1252 ();
 sg13g2_decap_8 FILLER_7_1279 ();
 sg13g2_decap_4 FILLER_7_1286 ();
 sg13g2_fill_2 FILLER_7_1290 ();
 sg13g2_fill_1 FILLER_7_1297 ();
 sg13g2_decap_8 FILLER_7_1324 ();
 sg13g2_decap_8 FILLER_7_1331 ();
 sg13g2_decap_8 FILLER_7_1338 ();
 sg13g2_decap_8 FILLER_7_1345 ();
 sg13g2_decap_8 FILLER_7_1352 ();
 sg13g2_decap_8 FILLER_7_1359 ();
 sg13g2_decap_8 FILLER_7_1366 ();
 sg13g2_decap_8 FILLER_7_1373 ();
 sg13g2_fill_2 FILLER_7_1380 ();
 sg13g2_decap_8 FILLER_7_1387 ();
 sg13g2_decap_8 FILLER_7_1394 ();
 sg13g2_decap_8 FILLER_7_1401 ();
 sg13g2_decap_8 FILLER_7_1408 ();
 sg13g2_decap_8 FILLER_7_1415 ();
 sg13g2_decap_4 FILLER_7_1422 ();
 sg13g2_decap_8 FILLER_7_1434 ();
 sg13g2_decap_8 FILLER_7_1441 ();
 sg13g2_decap_8 FILLER_7_1448 ();
 sg13g2_decap_8 FILLER_7_1455 ();
 sg13g2_decap_8 FILLER_7_1462 ();
 sg13g2_decap_8 FILLER_7_1469 ();
 sg13g2_decap_8 FILLER_7_1476 ();
 sg13g2_decap_4 FILLER_7_1483 ();
 sg13g2_decap_8 FILLER_7_1496 ();
 sg13g2_fill_2 FILLER_7_1503 ();
 sg13g2_fill_1 FILLER_7_1505 ();
 sg13g2_decap_8 FILLER_7_1532 ();
 sg13g2_decap_8 FILLER_7_1539 ();
 sg13g2_fill_1 FILLER_7_1546 ();
 sg13g2_fill_1 FILLER_7_1552 ();
 sg13g2_decap_8 FILLER_7_1563 ();
 sg13g2_decap_8 FILLER_7_1570 ();
 sg13g2_fill_2 FILLER_7_1577 ();
 sg13g2_decap_8 FILLER_7_1589 ();
 sg13g2_decap_8 FILLER_7_1596 ();
 sg13g2_decap_8 FILLER_7_1603 ();
 sg13g2_decap_8 FILLER_7_1610 ();
 sg13g2_decap_8 FILLER_7_1617 ();
 sg13g2_decap_8 FILLER_7_1624 ();
 sg13g2_decap_8 FILLER_7_1636 ();
 sg13g2_decap_8 FILLER_7_1643 ();
 sg13g2_decap_8 FILLER_7_1650 ();
 sg13g2_fill_2 FILLER_7_1657 ();
 sg13g2_fill_1 FILLER_7_1659 ();
 sg13g2_fill_2 FILLER_7_1670 ();
 sg13g2_decap_8 FILLER_7_1681 ();
 sg13g2_decap_8 FILLER_7_1688 ();
 sg13g2_decap_8 FILLER_7_1695 ();
 sg13g2_decap_8 FILLER_7_1702 ();
 sg13g2_decap_8 FILLER_7_1709 ();
 sg13g2_fill_2 FILLER_7_1716 ();
 sg13g2_decap_8 FILLER_7_1749 ();
 sg13g2_fill_1 FILLER_7_1756 ();
 sg13g2_decap_4 FILLER_7_1804 ();
 sg13g2_fill_2 FILLER_7_1808 ();
 sg13g2_decap_8 FILLER_7_1815 ();
 sg13g2_decap_4 FILLER_7_1822 ();
 sg13g2_decap_4 FILLER_7_1836 ();
 sg13g2_decap_8 FILLER_7_1845 ();
 sg13g2_decap_4 FILLER_7_1852 ();
 sg13g2_decap_8 FILLER_7_1861 ();
 sg13g2_decap_4 FILLER_7_1868 ();
 sg13g2_fill_2 FILLER_7_1872 ();
 sg13g2_decap_8 FILLER_7_1905 ();
 sg13g2_decap_8 FILLER_7_1912 ();
 sg13g2_decap_8 FILLER_7_1919 ();
 sg13g2_decap_8 FILLER_7_1926 ();
 sg13g2_decap_8 FILLER_7_1933 ();
 sg13g2_decap_8 FILLER_7_1940 ();
 sg13g2_decap_8 FILLER_7_1947 ();
 sg13g2_decap_8 FILLER_7_1954 ();
 sg13g2_decap_8 FILLER_7_1961 ();
 sg13g2_decap_8 FILLER_7_1968 ();
 sg13g2_decap_8 FILLER_7_1975 ();
 sg13g2_decap_8 FILLER_7_1982 ();
 sg13g2_fill_2 FILLER_7_1989 ();
 sg13g2_fill_1 FILLER_7_1991 ();
 sg13g2_fill_2 FILLER_7_2018 ();
 sg13g2_decap_8 FILLER_7_2046 ();
 sg13g2_decap_8 FILLER_7_2053 ();
 sg13g2_decap_8 FILLER_7_2060 ();
 sg13g2_decap_8 FILLER_7_2067 ();
 sg13g2_fill_2 FILLER_7_2074 ();
 sg13g2_decap_8 FILLER_7_2107 ();
 sg13g2_decap_4 FILLER_7_2114 ();
 sg13g2_fill_2 FILLER_7_2118 ();
 sg13g2_decap_4 FILLER_7_2151 ();
 sg13g2_fill_1 FILLER_7_2155 ();
 sg13g2_decap_8 FILLER_7_2186 ();
 sg13g2_fill_1 FILLER_7_2193 ();
 sg13g2_decap_8 FILLER_7_2227 ();
 sg13g2_fill_2 FILLER_7_2234 ();
 sg13g2_fill_1 FILLER_7_2236 ();
 sg13g2_decap_8 FILLER_7_2273 ();
 sg13g2_fill_1 FILLER_7_2280 ();
 sg13g2_decap_4 FILLER_7_2291 ();
 sg13g2_fill_1 FILLER_7_2295 ();
 sg13g2_decap_8 FILLER_7_2316 ();
 sg13g2_decap_8 FILLER_7_2323 ();
 sg13g2_fill_2 FILLER_7_2330 ();
 sg13g2_fill_2 FILLER_7_2336 ();
 sg13g2_decap_8 FILLER_7_2364 ();
 sg13g2_decap_8 FILLER_7_2371 ();
 sg13g2_decap_4 FILLER_7_2378 ();
 sg13g2_fill_1 FILLER_7_2382 ();
 sg13g2_decap_8 FILLER_7_2392 ();
 sg13g2_decap_8 FILLER_7_2399 ();
 sg13g2_decap_8 FILLER_7_2406 ();
 sg13g2_fill_1 FILLER_7_2413 ();
 sg13g2_fill_2 FILLER_7_2424 ();
 sg13g2_decap_8 FILLER_7_2446 ();
 sg13g2_fill_1 FILLER_7_2453 ();
 sg13g2_decap_8 FILLER_7_2501 ();
 sg13g2_decap_4 FILLER_7_2534 ();
 sg13g2_fill_1 FILLER_7_2538 ();
 sg13g2_decap_8 FILLER_7_2570 ();
 sg13g2_decap_8 FILLER_7_2577 ();
 sg13g2_decap_8 FILLER_7_2584 ();
 sg13g2_decap_4 FILLER_7_2591 ();
 sg13g2_fill_1 FILLER_7_2616 ();
 sg13g2_decap_8 FILLER_7_2694 ();
 sg13g2_decap_8 FILLER_7_2701 ();
 sg13g2_fill_2 FILLER_7_2708 ();
 sg13g2_fill_1 FILLER_7_2710 ();
 sg13g2_decap_4 FILLER_7_2730 ();
 sg13g2_fill_2 FILLER_7_2734 ();
 sg13g2_decap_8 FILLER_7_2749 ();
 sg13g2_decap_8 FILLER_7_2756 ();
 sg13g2_decap_8 FILLER_7_2763 ();
 sg13g2_decap_8 FILLER_7_2770 ();
 sg13g2_fill_2 FILLER_7_2777 ();
 sg13g2_decap_8 FILLER_7_2809 ();
 sg13g2_decap_4 FILLER_7_2816 ();
 sg13g2_fill_2 FILLER_7_2820 ();
 sg13g2_decap_8 FILLER_7_2853 ();
 sg13g2_decap_8 FILLER_7_2860 ();
 sg13g2_decap_8 FILLER_7_2867 ();
 sg13g2_decap_8 FILLER_7_2874 ();
 sg13g2_decap_8 FILLER_7_2881 ();
 sg13g2_decap_4 FILLER_7_2901 ();
 sg13g2_decap_8 FILLER_7_2920 ();
 sg13g2_decap_8 FILLER_7_2927 ();
 sg13g2_decap_8 FILLER_7_2934 ();
 sg13g2_decap_8 FILLER_7_2941 ();
 sg13g2_decap_8 FILLER_7_2948 ();
 sg13g2_decap_8 FILLER_7_2955 ();
 sg13g2_decap_8 FILLER_7_2962 ();
 sg13g2_decap_8 FILLER_7_2969 ();
 sg13g2_decap_8 FILLER_7_2976 ();
 sg13g2_decap_8 FILLER_7_2983 ();
 sg13g2_decap_8 FILLER_7_2990 ();
 sg13g2_decap_8 FILLER_7_3002 ();
 sg13g2_decap_8 FILLER_7_3014 ();
 sg13g2_decap_8 FILLER_7_3021 ();
 sg13g2_decap_8 FILLER_7_3028 ();
 sg13g2_decap_8 FILLER_7_3035 ();
 sg13g2_decap_8 FILLER_7_3051 ();
 sg13g2_decap_8 FILLER_7_3058 ();
 sg13g2_decap_8 FILLER_7_3065 ();
 sg13g2_decap_8 FILLER_7_3072 ();
 sg13g2_decap_8 FILLER_7_3079 ();
 sg13g2_decap_8 FILLER_7_3086 ();
 sg13g2_decap_8 FILLER_7_3093 ();
 sg13g2_decap_8 FILLER_7_3100 ();
 sg13g2_decap_8 FILLER_7_3107 ();
 sg13g2_decap_8 FILLER_7_3114 ();
 sg13g2_decap_8 FILLER_7_3121 ();
 sg13g2_decap_8 FILLER_7_3128 ();
 sg13g2_fill_2 FILLER_7_3135 ();
 sg13g2_fill_1 FILLER_7_3137 ();
 sg13g2_decap_8 FILLER_7_3158 ();
 sg13g2_decap_8 FILLER_7_3165 ();
 sg13g2_fill_1 FILLER_7_3172 ();
 sg13g2_decap_4 FILLER_7_3189 ();
 sg13g2_fill_2 FILLER_7_3193 ();
 sg13g2_decap_8 FILLER_7_3200 ();
 sg13g2_fill_1 FILLER_7_3207 ();
 sg13g2_decap_8 FILLER_7_3212 ();
 sg13g2_decap_8 FILLER_7_3219 ();
 sg13g2_decap_8 FILLER_7_3226 ();
 sg13g2_fill_2 FILLER_7_3233 ();
 sg13g2_decap_8 FILLER_7_3244 ();
 sg13g2_decap_8 FILLER_7_3251 ();
 sg13g2_decap_8 FILLER_7_3258 ();
 sg13g2_fill_1 FILLER_7_3265 ();
 sg13g2_decap_4 FILLER_7_3292 ();
 sg13g2_fill_2 FILLER_7_3296 ();
 sg13g2_decap_8 FILLER_7_3303 ();
 sg13g2_decap_8 FILLER_7_3310 ();
 sg13g2_decap_8 FILLER_7_3317 ();
 sg13g2_decap_8 FILLER_7_3324 ();
 sg13g2_decap_8 FILLER_7_3331 ();
 sg13g2_decap_8 FILLER_7_3338 ();
 sg13g2_decap_8 FILLER_7_3345 ();
 sg13g2_decap_8 FILLER_7_3352 ();
 sg13g2_decap_4 FILLER_7_3359 ();
 sg13g2_fill_1 FILLER_7_3363 ();
 sg13g2_decap_8 FILLER_7_3372 ();
 sg13g2_decap_8 FILLER_7_3379 ();
 sg13g2_decap_8 FILLER_7_3386 ();
 sg13g2_decap_8 FILLER_7_3393 ();
 sg13g2_decap_8 FILLER_7_3400 ();
 sg13g2_decap_4 FILLER_7_3407 ();
 sg13g2_fill_1 FILLER_7_3411 ();
 sg13g2_decap_8 FILLER_7_3422 ();
 sg13g2_fill_2 FILLER_7_3429 ();
 sg13g2_fill_1 FILLER_7_3431 ();
 sg13g2_decap_8 FILLER_7_3441 ();
 sg13g2_decap_8 FILLER_7_3448 ();
 sg13g2_decap_8 FILLER_7_3455 ();
 sg13g2_decap_8 FILLER_7_3462 ();
 sg13g2_decap_8 FILLER_7_3469 ();
 sg13g2_decap_8 FILLER_7_3476 ();
 sg13g2_decap_8 FILLER_7_3483 ();
 sg13g2_decap_8 FILLER_7_3490 ();
 sg13g2_decap_8 FILLER_7_3497 ();
 sg13g2_decap_8 FILLER_7_3504 ();
 sg13g2_decap_8 FILLER_7_3511 ();
 sg13g2_decap_8 FILLER_7_3518 ();
 sg13g2_decap_8 FILLER_7_3525 ();
 sg13g2_decap_8 FILLER_7_3532 ();
 sg13g2_decap_8 FILLER_7_3539 ();
 sg13g2_decap_8 FILLER_7_3546 ();
 sg13g2_decap_8 FILLER_7_3553 ();
 sg13g2_decap_8 FILLER_7_3560 ();
 sg13g2_decap_8 FILLER_7_3567 ();
 sg13g2_decap_4 FILLER_7_3574 ();
 sg13g2_fill_2 FILLER_7_3578 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_4 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_92 ();
 sg13g2_decap_8 FILLER_8_99 ();
 sg13g2_decap_8 FILLER_8_106 ();
 sg13g2_decap_8 FILLER_8_113 ();
 sg13g2_decap_8 FILLER_8_120 ();
 sg13g2_fill_2 FILLER_8_127 ();
 sg13g2_decap_8 FILLER_8_160 ();
 sg13g2_decap_8 FILLER_8_167 ();
 sg13g2_fill_1 FILLER_8_174 ();
 sg13g2_decap_4 FILLER_8_190 ();
 sg13g2_decap_8 FILLER_8_204 ();
 sg13g2_decap_8 FILLER_8_211 ();
 sg13g2_decap_8 FILLER_8_218 ();
 sg13g2_decap_8 FILLER_8_225 ();
 sg13g2_fill_1 FILLER_8_232 ();
 sg13g2_decap_4 FILLER_8_268 ();
 sg13g2_fill_2 FILLER_8_272 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_4 FILLER_8_322 ();
 sg13g2_fill_2 FILLER_8_326 ();
 sg13g2_decap_8 FILLER_8_360 ();
 sg13g2_decap_8 FILLER_8_367 ();
 sg13g2_decap_4 FILLER_8_374 ();
 sg13g2_fill_2 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_403 ();
 sg13g2_decap_8 FILLER_8_410 ();
 sg13g2_decap_4 FILLER_8_417 ();
 sg13g2_fill_1 FILLER_8_421 ();
 sg13g2_decap_4 FILLER_8_427 ();
 sg13g2_fill_1 FILLER_8_431 ();
 sg13g2_decap_8 FILLER_8_440 ();
 sg13g2_fill_2 FILLER_8_447 ();
 sg13g2_fill_1 FILLER_8_449 ();
 sg13g2_decap_8 FILLER_8_455 ();
 sg13g2_decap_8 FILLER_8_462 ();
 sg13g2_decap_8 FILLER_8_469 ();
 sg13g2_decap_8 FILLER_8_476 ();
 sg13g2_decap_8 FILLER_8_483 ();
 sg13g2_fill_2 FILLER_8_490 ();
 sg13g2_fill_1 FILLER_8_492 ();
 sg13g2_decap_8 FILLER_8_501 ();
 sg13g2_fill_2 FILLER_8_508 ();
 sg13g2_decap_8 FILLER_8_545 ();
 sg13g2_fill_1 FILLER_8_552 ();
 sg13g2_decap_8 FILLER_8_589 ();
 sg13g2_decap_8 FILLER_8_596 ();
 sg13g2_decap_8 FILLER_8_603 ();
 sg13g2_decap_4 FILLER_8_610 ();
 sg13g2_decap_8 FILLER_8_644 ();
 sg13g2_decap_8 FILLER_8_651 ();
 sg13g2_decap_8 FILLER_8_658 ();
 sg13g2_decap_8 FILLER_8_665 ();
 sg13g2_fill_1 FILLER_8_672 ();
 sg13g2_decap_8 FILLER_8_678 ();
 sg13g2_decap_8 FILLER_8_685 ();
 sg13g2_decap_4 FILLER_8_692 ();
 sg13g2_fill_1 FILLER_8_696 ();
 sg13g2_fill_2 FILLER_8_711 ();
 sg13g2_fill_1 FILLER_8_713 ();
 sg13g2_decap_8 FILLER_8_726 ();
 sg13g2_decap_8 FILLER_8_733 ();
 sg13g2_decap_8 FILLER_8_740 ();
 sg13g2_decap_8 FILLER_8_747 ();
 sg13g2_decap_8 FILLER_8_754 ();
 sg13g2_decap_4 FILLER_8_761 ();
 sg13g2_fill_1 FILLER_8_765 ();
 sg13g2_decap_8 FILLER_8_797 ();
 sg13g2_decap_8 FILLER_8_804 ();
 sg13g2_decap_8 FILLER_8_811 ();
 sg13g2_decap_8 FILLER_8_818 ();
 sg13g2_decap_8 FILLER_8_825 ();
 sg13g2_decap_8 FILLER_8_832 ();
 sg13g2_decap_8 FILLER_8_839 ();
 sg13g2_decap_8 FILLER_8_846 ();
 sg13g2_decap_8 FILLER_8_853 ();
 sg13g2_decap_8 FILLER_8_860 ();
 sg13g2_decap_8 FILLER_8_867 ();
 sg13g2_decap_8 FILLER_8_874 ();
 sg13g2_decap_4 FILLER_8_881 ();
 sg13g2_fill_2 FILLER_8_885 ();
 sg13g2_decap_4 FILLER_8_922 ();
 sg13g2_fill_1 FILLER_8_926 ();
 sg13g2_decap_8 FILLER_8_963 ();
 sg13g2_decap_8 FILLER_8_970 ();
 sg13g2_decap_8 FILLER_8_977 ();
 sg13g2_decap_8 FILLER_8_984 ();
 sg13g2_decap_8 FILLER_8_991 ();
 sg13g2_decap_8 FILLER_8_1001 ();
 sg13g2_fill_1 FILLER_8_1008 ();
 sg13g2_decap_4 FILLER_8_1035 ();
 sg13g2_fill_1 FILLER_8_1039 ();
 sg13g2_fill_2 FILLER_8_1044 ();
 sg13g2_fill_1 FILLER_8_1046 ();
 sg13g2_fill_2 FILLER_8_1052 ();
 sg13g2_fill_1 FILLER_8_1054 ();
 sg13g2_decap_8 FILLER_8_1064 ();
 sg13g2_decap_8 FILLER_8_1071 ();
 sg13g2_fill_1 FILLER_8_1078 ();
 sg13g2_fill_2 FILLER_8_1084 ();
 sg13g2_fill_1 FILLER_8_1086 ();
 sg13g2_decap_4 FILLER_8_1092 ();
 sg13g2_fill_2 FILLER_8_1096 ();
 sg13g2_decap_8 FILLER_8_1107 ();
 sg13g2_decap_8 FILLER_8_1114 ();
 sg13g2_decap_8 FILLER_8_1121 ();
 sg13g2_decap_8 FILLER_8_1128 ();
 sg13g2_decap_8 FILLER_8_1135 ();
 sg13g2_fill_1 FILLER_8_1142 ();
 sg13g2_decap_8 FILLER_8_1153 ();
 sg13g2_decap_8 FILLER_8_1160 ();
 sg13g2_decap_4 FILLER_8_1173 ();
 sg13g2_fill_1 FILLER_8_1177 ();
 sg13g2_decap_8 FILLER_8_1204 ();
 sg13g2_decap_8 FILLER_8_1211 ();
 sg13g2_decap_8 FILLER_8_1218 ();
 sg13g2_decap_8 FILLER_8_1225 ();
 sg13g2_decap_8 FILLER_8_1232 ();
 sg13g2_decap_8 FILLER_8_1239 ();
 sg13g2_decap_8 FILLER_8_1246 ();
 sg13g2_fill_1 FILLER_8_1253 ();
 sg13g2_fill_1 FILLER_8_1272 ();
 sg13g2_fill_1 FILLER_8_1282 ();
 sg13g2_decap_8 FILLER_8_1323 ();
 sg13g2_decap_8 FILLER_8_1330 ();
 sg13g2_decap_8 FILLER_8_1337 ();
 sg13g2_decap_8 FILLER_8_1344 ();
 sg13g2_decap_8 FILLER_8_1351 ();
 sg13g2_fill_2 FILLER_8_1358 ();
 sg13g2_fill_1 FILLER_8_1360 ();
 sg13g2_decap_8 FILLER_8_1387 ();
 sg13g2_decap_4 FILLER_8_1394 ();
 sg13g2_decap_8 FILLER_8_1424 ();
 sg13g2_decap_8 FILLER_8_1431 ();
 sg13g2_fill_2 FILLER_8_1438 ();
 sg13g2_fill_1 FILLER_8_1440 ();
 sg13g2_decap_4 FILLER_8_1467 ();
 sg13g2_decap_8 FILLER_8_1507 ();
 sg13g2_decap_8 FILLER_8_1514 ();
 sg13g2_fill_2 FILLER_8_1521 ();
 sg13g2_fill_1 FILLER_8_1523 ();
 sg13g2_fill_2 FILLER_8_1529 ();
 sg13g2_decap_8 FILLER_8_1539 ();
 sg13g2_decap_8 FILLER_8_1546 ();
 sg13g2_decap_8 FILLER_8_1553 ();
 sg13g2_decap_8 FILLER_8_1560 ();
 sg13g2_decap_4 FILLER_8_1567 ();
 sg13g2_fill_2 FILLER_8_1571 ();
 sg13g2_decap_8 FILLER_8_1604 ();
 sg13g2_decap_8 FILLER_8_1611 ();
 sg13g2_decap_4 FILLER_8_1618 ();
 sg13g2_fill_2 FILLER_8_1622 ();
 sg13g2_decap_8 FILLER_8_1632 ();
 sg13g2_decap_8 FILLER_8_1639 ();
 sg13g2_fill_2 FILLER_8_1646 ();
 sg13g2_decap_8 FILLER_8_1674 ();
 sg13g2_decap_8 FILLER_8_1707 ();
 sg13g2_decap_8 FILLER_8_1714 ();
 sg13g2_decap_8 FILLER_8_1721 ();
 sg13g2_decap_8 FILLER_8_1736 ();
 sg13g2_decap_8 FILLER_8_1743 ();
 sg13g2_decap_8 FILLER_8_1750 ();
 sg13g2_decap_4 FILLER_8_1757 ();
 sg13g2_fill_2 FILLER_8_1761 ();
 sg13g2_decap_8 FILLER_8_1767 ();
 sg13g2_decap_8 FILLER_8_1774 ();
 sg13g2_decap_4 FILLER_8_1781 ();
 sg13g2_fill_2 FILLER_8_1785 ();
 sg13g2_decap_8 FILLER_8_1792 ();
 sg13g2_decap_4 FILLER_8_1799 ();
 sg13g2_fill_1 FILLER_8_1803 ();
 sg13g2_fill_2 FILLER_8_1809 ();
 sg13g2_fill_1 FILLER_8_1811 ();
 sg13g2_fill_2 FILLER_8_1822 ();
 sg13g2_fill_1 FILLER_8_1824 ();
 sg13g2_decap_8 FILLER_8_1835 ();
 sg13g2_decap_8 FILLER_8_1842 ();
 sg13g2_decap_8 FILLER_8_1849 ();
 sg13g2_decap_8 FILLER_8_1856 ();
 sg13g2_decap_8 FILLER_8_1863 ();
 sg13g2_fill_2 FILLER_8_1870 ();
 sg13g2_decap_8 FILLER_8_1892 ();
 sg13g2_decap_8 FILLER_8_1904 ();
 sg13g2_decap_8 FILLER_8_1911 ();
 sg13g2_decap_8 FILLER_8_1918 ();
 sg13g2_fill_1 FILLER_8_1925 ();
 sg13g2_decap_8 FILLER_8_1936 ();
 sg13g2_decap_4 FILLER_8_1943 ();
 sg13g2_fill_1 FILLER_8_1947 ();
 sg13g2_decap_8 FILLER_8_1974 ();
 sg13g2_fill_2 FILLER_8_1981 ();
 sg13g2_decap_8 FILLER_8_1993 ();
 sg13g2_decap_8 FILLER_8_2000 ();
 sg13g2_decap_4 FILLER_8_2007 ();
 sg13g2_fill_2 FILLER_8_2011 ();
 sg13g2_decap_8 FILLER_8_2023 ();
 sg13g2_fill_2 FILLER_8_2030 ();
 sg13g2_decap_8 FILLER_8_2058 ();
 sg13g2_decap_8 FILLER_8_2065 ();
 sg13g2_decap_8 FILLER_8_2072 ();
 sg13g2_decap_8 FILLER_8_2079 ();
 sg13g2_decap_4 FILLER_8_2086 ();
 sg13g2_decap_8 FILLER_8_2102 ();
 sg13g2_decap_8 FILLER_8_2109 ();
 sg13g2_decap_8 FILLER_8_2116 ();
 sg13g2_decap_8 FILLER_8_2123 ();
 sg13g2_fill_1 FILLER_8_2130 ();
 sg13g2_decap_8 FILLER_8_2136 ();
 sg13g2_decap_8 FILLER_8_2143 ();
 sg13g2_decap_8 FILLER_8_2150 ();
 sg13g2_decap_8 FILLER_8_2157 ();
 sg13g2_fill_2 FILLER_8_2164 ();
 sg13g2_decap_8 FILLER_8_2180 ();
 sg13g2_decap_8 FILLER_8_2187 ();
 sg13g2_decap_8 FILLER_8_2194 ();
 sg13g2_decap_8 FILLER_8_2201 ();
 sg13g2_fill_1 FILLER_8_2208 ();
 sg13g2_decap_8 FILLER_8_2220 ();
 sg13g2_decap_8 FILLER_8_2227 ();
 sg13g2_decap_8 FILLER_8_2234 ();
 sg13g2_decap_4 FILLER_8_2241 ();
 sg13g2_fill_1 FILLER_8_2245 ();
 sg13g2_decap_8 FILLER_8_2256 ();
 sg13g2_decap_8 FILLER_8_2263 ();
 sg13g2_decap_8 FILLER_8_2270 ();
 sg13g2_decap_8 FILLER_8_2277 ();
 sg13g2_decap_8 FILLER_8_2284 ();
 sg13g2_decap_4 FILLER_8_2291 ();
 sg13g2_fill_2 FILLER_8_2295 ();
 sg13g2_fill_2 FILLER_8_2306 ();
 sg13g2_fill_1 FILLER_8_2308 ();
 sg13g2_decap_8 FILLER_8_2319 ();
 sg13g2_decap_8 FILLER_8_2326 ();
 sg13g2_decap_8 FILLER_8_2333 ();
 sg13g2_decap_8 FILLER_8_2340 ();
 sg13g2_fill_2 FILLER_8_2347 ();
 sg13g2_decap_8 FILLER_8_2374 ();
 sg13g2_decap_8 FILLER_8_2381 ();
 sg13g2_decap_4 FILLER_8_2388 ();
 sg13g2_decap_8 FILLER_8_2400 ();
 sg13g2_decap_8 FILLER_8_2407 ();
 sg13g2_decap_8 FILLER_8_2414 ();
 sg13g2_fill_1 FILLER_8_2421 ();
 sg13g2_decap_8 FILLER_8_2444 ();
 sg13g2_decap_8 FILLER_8_2451 ();
 sg13g2_decap_8 FILLER_8_2458 ();
 sg13g2_decap_8 FILLER_8_2465 ();
 sg13g2_decap_8 FILLER_8_2472 ();
 sg13g2_fill_1 FILLER_8_2479 ();
 sg13g2_decap_8 FILLER_8_2495 ();
 sg13g2_decap_8 FILLER_8_2502 ();
 sg13g2_decap_4 FILLER_8_2509 ();
 sg13g2_fill_1 FILLER_8_2513 ();
 sg13g2_decap_8 FILLER_8_2529 ();
 sg13g2_decap_8 FILLER_8_2536 ();
 sg13g2_decap_8 FILLER_8_2543 ();
 sg13g2_decap_8 FILLER_8_2560 ();
 sg13g2_decap_8 FILLER_8_2567 ();
 sg13g2_decap_8 FILLER_8_2574 ();
 sg13g2_decap_8 FILLER_8_2581 ();
 sg13g2_decap_8 FILLER_8_2588 ();
 sg13g2_decap_4 FILLER_8_2595 ();
 sg13g2_fill_2 FILLER_8_2599 ();
 sg13g2_fill_1 FILLER_8_2606 ();
 sg13g2_fill_2 FILLER_8_2627 ();
 sg13g2_fill_1 FILLER_8_2629 ();
 sg13g2_decap_8 FILLER_8_2635 ();
 sg13g2_decap_8 FILLER_8_2642 ();
 sg13g2_fill_2 FILLER_8_2649 ();
 sg13g2_fill_1 FILLER_8_2651 ();
 sg13g2_fill_2 FILLER_8_2661 ();
 sg13g2_fill_1 FILLER_8_2663 ();
 sg13g2_fill_2 FILLER_8_2674 ();
 sg13g2_fill_1 FILLER_8_2676 ();
 sg13g2_decap_8 FILLER_8_2692 ();
 sg13g2_decap_8 FILLER_8_2699 ();
 sg13g2_decap_8 FILLER_8_2706 ();
 sg13g2_decap_8 FILLER_8_2713 ();
 sg13g2_decap_8 FILLER_8_2720 ();
 sg13g2_decap_8 FILLER_8_2727 ();
 sg13g2_decap_8 FILLER_8_2734 ();
 sg13g2_decap_8 FILLER_8_2741 ();
 sg13g2_decap_8 FILLER_8_2748 ();
 sg13g2_decap_8 FILLER_8_2755 ();
 sg13g2_decap_8 FILLER_8_2762 ();
 sg13g2_decap_8 FILLER_8_2769 ();
 sg13g2_decap_8 FILLER_8_2776 ();
 sg13g2_fill_2 FILLER_8_2783 ();
 sg13g2_fill_1 FILLER_8_2785 ();
 sg13g2_decap_8 FILLER_8_2802 ();
 sg13g2_decap_8 FILLER_8_2809 ();
 sg13g2_decap_8 FILLER_8_2816 ();
 sg13g2_decap_8 FILLER_8_2823 ();
 sg13g2_fill_1 FILLER_8_2830 ();
 sg13g2_fill_1 FILLER_8_2836 ();
 sg13g2_decap_8 FILLER_8_2842 ();
 sg13g2_decap_8 FILLER_8_2849 ();
 sg13g2_decap_8 FILLER_8_2856 ();
 sg13g2_fill_1 FILLER_8_2863 ();
 sg13g2_decap_8 FILLER_8_2868 ();
 sg13g2_decap_8 FILLER_8_2875 ();
 sg13g2_decap_8 FILLER_8_2882 ();
 sg13g2_decap_8 FILLER_8_2889 ();
 sg13g2_fill_1 FILLER_8_2896 ();
 sg13g2_fill_2 FILLER_8_2902 ();
 sg13g2_fill_1 FILLER_8_2904 ();
 sg13g2_decap_8 FILLER_8_2915 ();
 sg13g2_decap_8 FILLER_8_2922 ();
 sg13g2_decap_8 FILLER_8_2929 ();
 sg13g2_decap_8 FILLER_8_2936 ();
 sg13g2_decap_4 FILLER_8_2943 ();
 sg13g2_fill_1 FILLER_8_2947 ();
 sg13g2_decap_8 FILLER_8_2964 ();
 sg13g2_decap_8 FILLER_8_2979 ();
 sg13g2_fill_2 FILLER_8_2986 ();
 sg13g2_decap_8 FILLER_8_2996 ();
 sg13g2_decap_8 FILLER_8_3003 ();
 sg13g2_decap_4 FILLER_8_3010 ();
 sg13g2_fill_1 FILLER_8_3019 ();
 sg13g2_fill_1 FILLER_8_3025 ();
 sg13g2_decap_8 FILLER_8_3057 ();
 sg13g2_decap_8 FILLER_8_3064 ();
 sg13g2_decap_8 FILLER_8_3071 ();
 sg13g2_fill_2 FILLER_8_3078 ();
 sg13g2_fill_1 FILLER_8_3080 ();
 sg13g2_fill_1 FILLER_8_3091 ();
 sg13g2_decap_8 FILLER_8_3118 ();
 sg13g2_decap_8 FILLER_8_3125 ();
 sg13g2_decap_8 FILLER_8_3132 ();
 sg13g2_decap_8 FILLER_8_3139 ();
 sg13g2_fill_1 FILLER_8_3146 ();
 sg13g2_decap_8 FILLER_8_3152 ();
 sg13g2_decap_8 FILLER_8_3159 ();
 sg13g2_decap_4 FILLER_8_3166 ();
 sg13g2_fill_2 FILLER_8_3170 ();
 sg13g2_decap_8 FILLER_8_3176 ();
 sg13g2_decap_8 FILLER_8_3183 ();
 sg13g2_decap_8 FILLER_8_3190 ();
 sg13g2_decap_4 FILLER_8_3197 ();
 sg13g2_fill_1 FILLER_8_3201 ();
 sg13g2_decap_8 FILLER_8_3237 ();
 sg13g2_decap_8 FILLER_8_3244 ();
 sg13g2_decap_8 FILLER_8_3251 ();
 sg13g2_decap_8 FILLER_8_3258 ();
 sg13g2_decap_8 FILLER_8_3265 ();
 sg13g2_fill_1 FILLER_8_3272 ();
 sg13g2_decap_8 FILLER_8_3308 ();
 sg13g2_fill_1 FILLER_8_3356 ();
 sg13g2_decap_8 FILLER_8_3383 ();
 sg13g2_fill_2 FILLER_8_3390 ();
 sg13g2_decap_4 FILLER_8_3418 ();
 sg13g2_decap_8 FILLER_8_3456 ();
 sg13g2_decap_8 FILLER_8_3463 ();
 sg13g2_decap_8 FILLER_8_3470 ();
 sg13g2_decap_8 FILLER_8_3477 ();
 sg13g2_decap_8 FILLER_8_3484 ();
 sg13g2_decap_8 FILLER_8_3491 ();
 sg13g2_decap_8 FILLER_8_3498 ();
 sg13g2_decap_8 FILLER_8_3505 ();
 sg13g2_decap_8 FILLER_8_3512 ();
 sg13g2_decap_8 FILLER_8_3519 ();
 sg13g2_decap_8 FILLER_8_3526 ();
 sg13g2_decap_8 FILLER_8_3533 ();
 sg13g2_decap_8 FILLER_8_3540 ();
 sg13g2_decap_8 FILLER_8_3547 ();
 sg13g2_decap_8 FILLER_8_3554 ();
 sg13g2_decap_8 FILLER_8_3561 ();
 sg13g2_decap_8 FILLER_8_3568 ();
 sg13g2_decap_4 FILLER_8_3575 ();
 sg13g2_fill_1 FILLER_8_3579 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_4 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_96 ();
 sg13g2_decap_8 FILLER_9_103 ();
 sg13g2_decap_8 FILLER_9_110 ();
 sg13g2_decap_8 FILLER_9_117 ();
 sg13g2_decap_4 FILLER_9_124 ();
 sg13g2_decap_8 FILLER_9_159 ();
 sg13g2_decap_8 FILLER_9_166 ();
 sg13g2_fill_2 FILLER_9_173 ();
 sg13g2_fill_1 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_4 FILLER_9_273 ();
 sg13g2_fill_2 FILLER_9_277 ();
 sg13g2_decap_8 FILLER_9_313 ();
 sg13g2_decap_4 FILLER_9_320 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_408 ();
 sg13g2_decap_4 FILLER_9_415 ();
 sg13g2_fill_1 FILLER_9_419 ();
 sg13g2_decap_4 FILLER_9_428 ();
 sg13g2_fill_2 FILLER_9_432 ();
 sg13g2_decap_4 FILLER_9_439 ();
 sg13g2_fill_2 FILLER_9_443 ();
 sg13g2_decap_8 FILLER_9_461 ();
 sg13g2_decap_8 FILLER_9_468 ();
 sg13g2_decap_8 FILLER_9_475 ();
 sg13g2_fill_1 FILLER_9_482 ();
 sg13g2_fill_2 FILLER_9_488 ();
 sg13g2_fill_2 FILLER_9_515 ();
 sg13g2_fill_2 FILLER_9_522 ();
 sg13g2_decap_8 FILLER_9_534 ();
 sg13g2_decap_8 FILLER_9_541 ();
 sg13g2_decap_8 FILLER_9_548 ();
 sg13g2_decap_4 FILLER_9_555 ();
 sg13g2_fill_2 FILLER_9_559 ();
 sg13g2_decap_8 FILLER_9_587 ();
 sg13g2_decap_8 FILLER_9_594 ();
 sg13g2_fill_2 FILLER_9_601 ();
 sg13g2_fill_1 FILLER_9_603 ();
 sg13g2_fill_1 FILLER_9_614 ();
 sg13g2_fill_2 FILLER_9_629 ();
 sg13g2_decap_8 FILLER_9_643 ();
 sg13g2_decap_8 FILLER_9_650 ();
 sg13g2_decap_4 FILLER_9_657 ();
 sg13g2_fill_2 FILLER_9_661 ();
 sg13g2_decap_8 FILLER_9_671 ();
 sg13g2_decap_8 FILLER_9_678 ();
 sg13g2_decap_8 FILLER_9_685 ();
 sg13g2_fill_2 FILLER_9_692 ();
 sg13g2_decap_8 FILLER_9_746 ();
 sg13g2_decap_8 FILLER_9_753 ();
 sg13g2_decap_8 FILLER_9_760 ();
 sg13g2_decap_8 FILLER_9_767 ();
 sg13g2_fill_1 FILLER_9_774 ();
 sg13g2_decap_8 FILLER_9_780 ();
 sg13g2_decap_8 FILLER_9_787 ();
 sg13g2_decap_8 FILLER_9_794 ();
 sg13g2_decap_8 FILLER_9_801 ();
 sg13g2_decap_8 FILLER_9_808 ();
 sg13g2_decap_8 FILLER_9_815 ();
 sg13g2_decap_4 FILLER_9_822 ();
 sg13g2_fill_2 FILLER_9_826 ();
 sg13g2_decap_8 FILLER_9_854 ();
 sg13g2_decap_8 FILLER_9_861 ();
 sg13g2_decap_8 FILLER_9_868 ();
 sg13g2_decap_8 FILLER_9_875 ();
 sg13g2_decap_8 FILLER_9_882 ();
 sg13g2_fill_1 FILLER_9_889 ();
 sg13g2_decap_8 FILLER_9_916 ();
 sg13g2_decap_8 FILLER_9_923 ();
 sg13g2_decap_8 FILLER_9_930 ();
 sg13g2_decap_8 FILLER_9_937 ();
 sg13g2_decap_4 FILLER_9_944 ();
 sg13g2_fill_1 FILLER_9_948 ();
 sg13g2_fill_2 FILLER_9_984 ();
 sg13g2_fill_1 FILLER_9_986 ();
 sg13g2_decap_8 FILLER_9_997 ();
 sg13g2_decap_8 FILLER_9_1004 ();
 sg13g2_decap_8 FILLER_9_1011 ();
 sg13g2_decap_8 FILLER_9_1018 ();
 sg13g2_decap_8 FILLER_9_1025 ();
 sg13g2_decap_4 FILLER_9_1032 ();
 sg13g2_fill_2 FILLER_9_1036 ();
 sg13g2_decap_8 FILLER_9_1055 ();
 sg13g2_decap_8 FILLER_9_1062 ();
 sg13g2_decap_8 FILLER_9_1069 ();
 sg13g2_decap_8 FILLER_9_1076 ();
 sg13g2_decap_8 FILLER_9_1083 ();
 sg13g2_decap_8 FILLER_9_1090 ();
 sg13g2_fill_1 FILLER_9_1097 ();
 sg13g2_decap_8 FILLER_9_1133 ();
 sg13g2_decap_8 FILLER_9_1140 ();
 sg13g2_decap_8 FILLER_9_1147 ();
 sg13g2_decap_8 FILLER_9_1154 ();
 sg13g2_decap_8 FILLER_9_1161 ();
 sg13g2_decap_8 FILLER_9_1168 ();
 sg13g2_decap_8 FILLER_9_1175 ();
 sg13g2_decap_8 FILLER_9_1182 ();
 sg13g2_decap_8 FILLER_9_1189 ();
 sg13g2_decap_8 FILLER_9_1196 ();
 sg13g2_decap_8 FILLER_9_1203 ();
 sg13g2_decap_8 FILLER_9_1210 ();
 sg13g2_decap_8 FILLER_9_1217 ();
 sg13g2_decap_8 FILLER_9_1224 ();
 sg13g2_decap_8 FILLER_9_1231 ();
 sg13g2_decap_8 FILLER_9_1238 ();
 sg13g2_decap_8 FILLER_9_1245 ();
 sg13g2_decap_8 FILLER_9_1252 ();
 sg13g2_fill_1 FILLER_9_1263 ();
 sg13g2_decap_8 FILLER_9_1273 ();
 sg13g2_decap_8 FILLER_9_1280 ();
 sg13g2_fill_2 FILLER_9_1287 ();
 sg13g2_fill_1 FILLER_9_1289 ();
 sg13g2_fill_1 FILLER_9_1304 ();
 sg13g2_decap_8 FILLER_9_1328 ();
 sg13g2_fill_1 FILLER_9_1335 ();
 sg13g2_decap_8 FILLER_9_1372 ();
 sg13g2_decap_8 FILLER_9_1379 ();
 sg13g2_decap_8 FILLER_9_1386 ();
 sg13g2_decap_8 FILLER_9_1393 ();
 sg13g2_decap_4 FILLER_9_1400 ();
 sg13g2_fill_2 FILLER_9_1404 ();
 sg13g2_decap_4 FILLER_9_1409 ();
 sg13g2_fill_1 FILLER_9_1413 ();
 sg13g2_fill_2 FILLER_9_1435 ();
 sg13g2_decap_8 FILLER_9_1466 ();
 sg13g2_decap_8 FILLER_9_1473 ();
 sg13g2_decap_8 FILLER_9_1480 ();
 sg13g2_decap_8 FILLER_9_1487 ();
 sg13g2_decap_8 FILLER_9_1494 ();
 sg13g2_decap_8 FILLER_9_1501 ();
 sg13g2_decap_8 FILLER_9_1508 ();
 sg13g2_decap_8 FILLER_9_1515 ();
 sg13g2_decap_4 FILLER_9_1522 ();
 sg13g2_fill_2 FILLER_9_1526 ();
 sg13g2_decap_8 FILLER_9_1559 ();
 sg13g2_decap_8 FILLER_9_1571 ();
 sg13g2_fill_2 FILLER_9_1578 ();
 sg13g2_fill_1 FILLER_9_1580 ();
 sg13g2_fill_2 FILLER_9_1590 ();
 sg13g2_decap_8 FILLER_9_1606 ();
 sg13g2_decap_8 FILLER_9_1613 ();
 sg13g2_fill_1 FILLER_9_1620 ();
 sg13g2_decap_8 FILLER_9_1626 ();
 sg13g2_fill_1 FILLER_9_1633 ();
 sg13g2_decap_8 FILLER_9_1642 ();
 sg13g2_decap_8 FILLER_9_1649 ();
 sg13g2_fill_1 FILLER_9_1656 ();
 sg13g2_fill_2 FILLER_9_1702 ();
 sg13g2_fill_1 FILLER_9_1704 ();
 sg13g2_decap_8 FILLER_9_1710 ();
 sg13g2_decap_8 FILLER_9_1717 ();
 sg13g2_decap_8 FILLER_9_1724 ();
 sg13g2_decap_8 FILLER_9_1731 ();
 sg13g2_fill_1 FILLER_9_1738 ();
 sg13g2_decap_8 FILLER_9_1754 ();
 sg13g2_decap_8 FILLER_9_1761 ();
 sg13g2_decap_8 FILLER_9_1768 ();
 sg13g2_decap_8 FILLER_9_1775 ();
 sg13g2_decap_8 FILLER_9_1782 ();
 sg13g2_decap_8 FILLER_9_1789 ();
 sg13g2_decap_8 FILLER_9_1796 ();
 sg13g2_decap_8 FILLER_9_1803 ();
 sg13g2_decap_4 FILLER_9_1810 ();
 sg13g2_fill_2 FILLER_9_1814 ();
 sg13g2_fill_2 FILLER_9_1821 ();
 sg13g2_decap_8 FILLER_9_1838 ();
 sg13g2_decap_8 FILLER_9_1845 ();
 sg13g2_decap_8 FILLER_9_1852 ();
 sg13g2_decap_8 FILLER_9_1859 ();
 sg13g2_decap_4 FILLER_9_1866 ();
 sg13g2_fill_2 FILLER_9_1870 ();
 sg13g2_fill_1 FILLER_9_1893 ();
 sg13g2_decap_8 FILLER_9_1904 ();
 sg13g2_decap_8 FILLER_9_1911 ();
 sg13g2_decap_4 FILLER_9_1918 ();
 sg13g2_decap_8 FILLER_9_1948 ();
 sg13g2_fill_2 FILLER_9_1955 ();
 sg13g2_decap_8 FILLER_9_1983 ();
 sg13g2_decap_8 FILLER_9_1990 ();
 sg13g2_decap_8 FILLER_9_1997 ();
 sg13g2_decap_8 FILLER_9_2004 ();
 sg13g2_decap_8 FILLER_9_2011 ();
 sg13g2_decap_8 FILLER_9_2018 ();
 sg13g2_decap_8 FILLER_9_2035 ();
 sg13g2_decap_8 FILLER_9_2042 ();
 sg13g2_decap_8 FILLER_9_2049 ();
 sg13g2_decap_8 FILLER_9_2056 ();
 sg13g2_decap_8 FILLER_9_2063 ();
 sg13g2_decap_8 FILLER_9_2070 ();
 sg13g2_decap_8 FILLER_9_2077 ();
 sg13g2_decap_4 FILLER_9_2084 ();
 sg13g2_decap_8 FILLER_9_2091 ();
 sg13g2_decap_8 FILLER_9_2098 ();
 sg13g2_decap_8 FILLER_9_2105 ();
 sg13g2_decap_8 FILLER_9_2112 ();
 sg13g2_decap_8 FILLER_9_2119 ();
 sg13g2_decap_8 FILLER_9_2126 ();
 sg13g2_decap_8 FILLER_9_2133 ();
 sg13g2_decap_8 FILLER_9_2140 ();
 sg13g2_decap_8 FILLER_9_2147 ();
 sg13g2_decap_8 FILLER_9_2154 ();
 sg13g2_decap_8 FILLER_9_2161 ();
 sg13g2_decap_8 FILLER_9_2168 ();
 sg13g2_decap_8 FILLER_9_2175 ();
 sg13g2_decap_8 FILLER_9_2182 ();
 sg13g2_decap_8 FILLER_9_2189 ();
 sg13g2_decap_4 FILLER_9_2196 ();
 sg13g2_fill_2 FILLER_9_2200 ();
 sg13g2_decap_8 FILLER_9_2207 ();
 sg13g2_decap_8 FILLER_9_2214 ();
 sg13g2_decap_8 FILLER_9_2221 ();
 sg13g2_decap_8 FILLER_9_2228 ();
 sg13g2_decap_8 FILLER_9_2235 ();
 sg13g2_decap_8 FILLER_9_2242 ();
 sg13g2_decap_8 FILLER_9_2249 ();
 sg13g2_decap_8 FILLER_9_2256 ();
 sg13g2_fill_2 FILLER_9_2263 ();
 sg13g2_decap_8 FILLER_9_2268 ();
 sg13g2_decap_8 FILLER_9_2275 ();
 sg13g2_decap_8 FILLER_9_2282 ();
 sg13g2_decap_8 FILLER_9_2289 ();
 sg13g2_decap_8 FILLER_9_2296 ();
 sg13g2_decap_8 FILLER_9_2303 ();
 sg13g2_decap_8 FILLER_9_2310 ();
 sg13g2_decap_8 FILLER_9_2317 ();
 sg13g2_decap_8 FILLER_9_2324 ();
 sg13g2_decap_8 FILLER_9_2331 ();
 sg13g2_decap_8 FILLER_9_2338 ();
 sg13g2_decap_8 FILLER_9_2345 ();
 sg13g2_decap_8 FILLER_9_2352 ();
 sg13g2_decap_8 FILLER_9_2359 ();
 sg13g2_decap_8 FILLER_9_2366 ();
 sg13g2_decap_8 FILLER_9_2373 ();
 sg13g2_decap_8 FILLER_9_2380 ();
 sg13g2_decap_8 FILLER_9_2387 ();
 sg13g2_decap_8 FILLER_9_2394 ();
 sg13g2_decap_8 FILLER_9_2401 ();
 sg13g2_fill_2 FILLER_9_2408 ();
 sg13g2_fill_1 FILLER_9_2410 ();
 sg13g2_decap_8 FILLER_9_2414 ();
 sg13g2_decap_8 FILLER_9_2421 ();
 sg13g2_decap_8 FILLER_9_2432 ();
 sg13g2_decap_8 FILLER_9_2439 ();
 sg13g2_decap_8 FILLER_9_2446 ();
 sg13g2_decap_8 FILLER_9_2453 ();
 sg13g2_decap_8 FILLER_9_2460 ();
 sg13g2_decap_8 FILLER_9_2467 ();
 sg13g2_decap_8 FILLER_9_2474 ();
 sg13g2_decap_8 FILLER_9_2481 ();
 sg13g2_decap_8 FILLER_9_2488 ();
 sg13g2_decap_8 FILLER_9_2495 ();
 sg13g2_decap_8 FILLER_9_2502 ();
 sg13g2_decap_8 FILLER_9_2509 ();
 sg13g2_decap_8 FILLER_9_2516 ();
 sg13g2_decap_8 FILLER_9_2523 ();
 sg13g2_decap_8 FILLER_9_2530 ();
 sg13g2_decap_8 FILLER_9_2537 ();
 sg13g2_decap_8 FILLER_9_2544 ();
 sg13g2_decap_8 FILLER_9_2551 ();
 sg13g2_decap_8 FILLER_9_2558 ();
 sg13g2_decap_8 FILLER_9_2565 ();
 sg13g2_decap_8 FILLER_9_2572 ();
 sg13g2_decap_8 FILLER_9_2579 ();
 sg13g2_decap_8 FILLER_9_2586 ();
 sg13g2_decap_8 FILLER_9_2593 ();
 sg13g2_decap_8 FILLER_9_2600 ();
 sg13g2_decap_8 FILLER_9_2607 ();
 sg13g2_decap_4 FILLER_9_2614 ();
 sg13g2_fill_1 FILLER_9_2618 ();
 sg13g2_decap_8 FILLER_9_2624 ();
 sg13g2_decap_8 FILLER_9_2631 ();
 sg13g2_decap_8 FILLER_9_2638 ();
 sg13g2_decap_8 FILLER_9_2645 ();
 sg13g2_decap_8 FILLER_9_2652 ();
 sg13g2_decap_8 FILLER_9_2659 ();
 sg13g2_decap_8 FILLER_9_2666 ();
 sg13g2_fill_2 FILLER_9_2673 ();
 sg13g2_decap_8 FILLER_9_2685 ();
 sg13g2_decap_8 FILLER_9_2692 ();
 sg13g2_decap_8 FILLER_9_2699 ();
 sg13g2_decap_8 FILLER_9_2706 ();
 sg13g2_decap_8 FILLER_9_2713 ();
 sg13g2_decap_8 FILLER_9_2720 ();
 sg13g2_decap_8 FILLER_9_2727 ();
 sg13g2_decap_8 FILLER_9_2744 ();
 sg13g2_decap_8 FILLER_9_2751 ();
 sg13g2_decap_8 FILLER_9_2758 ();
 sg13g2_decap_8 FILLER_9_2765 ();
 sg13g2_fill_1 FILLER_9_2772 ();
 sg13g2_decap_8 FILLER_9_2778 ();
 sg13g2_decap_8 FILLER_9_2785 ();
 sg13g2_decap_8 FILLER_9_2792 ();
 sg13g2_decap_8 FILLER_9_2799 ();
 sg13g2_decap_8 FILLER_9_2806 ();
 sg13g2_decap_8 FILLER_9_2813 ();
 sg13g2_decap_8 FILLER_9_2820 ();
 sg13g2_decap_8 FILLER_9_2827 ();
 sg13g2_decap_8 FILLER_9_2834 ();
 sg13g2_decap_8 FILLER_9_2841 ();
 sg13g2_decap_8 FILLER_9_2848 ();
 sg13g2_decap_8 FILLER_9_2855 ();
 sg13g2_decap_8 FILLER_9_2862 ();
 sg13g2_decap_8 FILLER_9_2869 ();
 sg13g2_decap_8 FILLER_9_2876 ();
 sg13g2_decap_8 FILLER_9_2883 ();
 sg13g2_fill_2 FILLER_9_2890 ();
 sg13g2_fill_1 FILLER_9_2892 ();
 sg13g2_fill_2 FILLER_9_2898 ();
 sg13g2_fill_1 FILLER_9_2900 ();
 sg13g2_decap_8 FILLER_9_2927 ();
 sg13g2_fill_1 FILLER_9_2934 ();
 sg13g2_decap_4 FILLER_9_2940 ();
 sg13g2_decap_8 FILLER_9_2996 ();
 sg13g2_decap_8 FILLER_9_3003 ();
 sg13g2_fill_2 FILLER_9_3010 ();
 sg13g2_decap_8 FILLER_9_3058 ();
 sg13g2_decap_4 FILLER_9_3065 ();
 sg13g2_fill_2 FILLER_9_3069 ();
 sg13g2_fill_2 FILLER_9_3092 ();
 sg13g2_decap_8 FILLER_9_3104 ();
 sg13g2_decap_4 FILLER_9_3111 ();
 sg13g2_decap_8 FILLER_9_3136 ();
 sg13g2_decap_8 FILLER_9_3143 ();
 sg13g2_decap_8 FILLER_9_3150 ();
 sg13g2_decap_4 FILLER_9_3157 ();
 sg13g2_fill_1 FILLER_9_3161 ();
 sg13g2_fill_2 FILLER_9_3167 ();
 sg13g2_fill_1 FILLER_9_3173 ();
 sg13g2_decap_8 FILLER_9_3184 ();
 sg13g2_fill_2 FILLER_9_3191 ();
 sg13g2_fill_1 FILLER_9_3193 ();
 sg13g2_fill_2 FILLER_9_3199 ();
 sg13g2_fill_1 FILLER_9_3201 ();
 sg13g2_decap_8 FILLER_9_3238 ();
 sg13g2_decap_8 FILLER_9_3245 ();
 sg13g2_decap_8 FILLER_9_3252 ();
 sg13g2_fill_2 FILLER_9_3259 ();
 sg13g2_fill_1 FILLER_9_3261 ();
 sg13g2_fill_1 FILLER_9_3267 ();
 sg13g2_decap_8 FILLER_9_3297 ();
 sg13g2_decap_8 FILLER_9_3304 ();
 sg13g2_decap_8 FILLER_9_3311 ();
 sg13g2_fill_2 FILLER_9_3344 ();
 sg13g2_decap_4 FILLER_9_3356 ();
 sg13g2_fill_2 FILLER_9_3360 ();
 sg13g2_decap_8 FILLER_9_3367 ();
 sg13g2_decap_8 FILLER_9_3374 ();
 sg13g2_decap_8 FILLER_9_3381 ();
 sg13g2_decap_8 FILLER_9_3388 ();
 sg13g2_decap_8 FILLER_9_3395 ();
 sg13g2_fill_2 FILLER_9_3402 ();
 sg13g2_fill_1 FILLER_9_3404 ();
 sg13g2_decap_4 FILLER_9_3409 ();
 sg13g2_decap_8 FILLER_9_3435 ();
 sg13g2_decap_8 FILLER_9_3442 ();
 sg13g2_decap_8 FILLER_9_3449 ();
 sg13g2_decap_8 FILLER_9_3456 ();
 sg13g2_decap_8 FILLER_9_3463 ();
 sg13g2_decap_8 FILLER_9_3470 ();
 sg13g2_decap_8 FILLER_9_3477 ();
 sg13g2_decap_8 FILLER_9_3484 ();
 sg13g2_decap_8 FILLER_9_3491 ();
 sg13g2_decap_8 FILLER_9_3498 ();
 sg13g2_decap_8 FILLER_9_3505 ();
 sg13g2_decap_8 FILLER_9_3512 ();
 sg13g2_decap_8 FILLER_9_3519 ();
 sg13g2_decap_8 FILLER_9_3526 ();
 sg13g2_decap_8 FILLER_9_3533 ();
 sg13g2_decap_8 FILLER_9_3540 ();
 sg13g2_decap_8 FILLER_9_3547 ();
 sg13g2_decap_8 FILLER_9_3554 ();
 sg13g2_decap_8 FILLER_9_3561 ();
 sg13g2_decap_8 FILLER_9_3568 ();
 sg13g2_decap_4 FILLER_9_3575 ();
 sg13g2_fill_1 FILLER_9_3579 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_4 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_29 ();
 sg13g2_decap_8 FILLER_10_36 ();
 sg13g2_decap_8 FILLER_10_43 ();
 sg13g2_decap_8 FILLER_10_50 ();
 sg13g2_fill_2 FILLER_10_57 ();
 sg13g2_decap_8 FILLER_10_85 ();
 sg13g2_decap_8 FILLER_10_92 ();
 sg13g2_decap_8 FILLER_10_99 ();
 sg13g2_decap_8 FILLER_10_106 ();
 sg13g2_decap_8 FILLER_10_113 ();
 sg13g2_decap_8 FILLER_10_120 ();
 sg13g2_decap_8 FILLER_10_127 ();
 sg13g2_decap_8 FILLER_10_134 ();
 sg13g2_fill_2 FILLER_10_141 ();
 sg13g2_fill_2 FILLER_10_147 ();
 sg13g2_fill_1 FILLER_10_149 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_fill_1 FILLER_10_182 ();
 sg13g2_fill_2 FILLER_10_187 ();
 sg13g2_decap_4 FILLER_10_210 ();
 sg13g2_fill_2 FILLER_10_214 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_fill_2 FILLER_10_287 ();
 sg13g2_fill_1 FILLER_10_289 ();
 sg13g2_decap_8 FILLER_10_299 ();
 sg13g2_decap_8 FILLER_10_306 ();
 sg13g2_decap_8 FILLER_10_313 ();
 sg13g2_decap_8 FILLER_10_320 ();
 sg13g2_fill_1 FILLER_10_335 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_fill_2 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_397 ();
 sg13g2_decap_4 FILLER_10_404 ();
 sg13g2_fill_2 FILLER_10_408 ();
 sg13g2_fill_1 FILLER_10_415 ();
 sg13g2_decap_8 FILLER_10_428 ();
 sg13g2_decap_8 FILLER_10_435 ();
 sg13g2_decap_4 FILLER_10_442 ();
 sg13g2_fill_1 FILLER_10_446 ();
 sg13g2_fill_2 FILLER_10_480 ();
 sg13g2_fill_1 FILLER_10_482 ();
 sg13g2_decap_4 FILLER_10_509 ();
 sg13g2_fill_2 FILLER_10_513 ();
 sg13g2_decap_8 FILLER_10_524 ();
 sg13g2_decap_8 FILLER_10_531 ();
 sg13g2_decap_8 FILLER_10_538 ();
 sg13g2_decap_8 FILLER_10_545 ();
 sg13g2_decap_8 FILLER_10_552 ();
 sg13g2_decap_8 FILLER_10_559 ();
 sg13g2_fill_1 FILLER_10_566 ();
 sg13g2_decap_8 FILLER_10_577 ();
 sg13g2_decap_8 FILLER_10_584 ();
 sg13g2_decap_8 FILLER_10_591 ();
 sg13g2_fill_2 FILLER_10_598 ();
 sg13g2_fill_1 FILLER_10_600 ();
 sg13g2_decap_8 FILLER_10_635 ();
 sg13g2_decap_8 FILLER_10_642 ();
 sg13g2_decap_8 FILLER_10_649 ();
 sg13g2_decap_8 FILLER_10_656 ();
 sg13g2_decap_8 FILLER_10_663 ();
 sg13g2_decap_4 FILLER_10_670 ();
 sg13g2_fill_2 FILLER_10_674 ();
 sg13g2_decap_4 FILLER_10_680 ();
 sg13g2_fill_2 FILLER_10_694 ();
 sg13g2_fill_1 FILLER_10_696 ();
 sg13g2_decap_8 FILLER_10_707 ();
 sg13g2_fill_2 FILLER_10_714 ();
 sg13g2_decap_8 FILLER_10_726 ();
 sg13g2_decap_8 FILLER_10_733 ();
 sg13g2_decap_8 FILLER_10_740 ();
 sg13g2_decap_8 FILLER_10_747 ();
 sg13g2_decap_8 FILLER_10_754 ();
 sg13g2_decap_8 FILLER_10_761 ();
 sg13g2_decap_8 FILLER_10_768 ();
 sg13g2_decap_8 FILLER_10_775 ();
 sg13g2_decap_8 FILLER_10_782 ();
 sg13g2_decap_8 FILLER_10_789 ();
 sg13g2_decap_8 FILLER_10_796 ();
 sg13g2_decap_8 FILLER_10_803 ();
 sg13g2_decap_8 FILLER_10_810 ();
 sg13g2_decap_8 FILLER_10_817 ();
 sg13g2_fill_1 FILLER_10_824 ();
 sg13g2_decap_8 FILLER_10_869 ();
 sg13g2_decap_8 FILLER_10_876 ();
 sg13g2_decap_8 FILLER_10_883 ();
 sg13g2_decap_8 FILLER_10_890 ();
 sg13g2_fill_2 FILLER_10_897 ();
 sg13g2_fill_1 FILLER_10_909 ();
 sg13g2_decap_8 FILLER_10_919 ();
 sg13g2_decap_8 FILLER_10_926 ();
 sg13g2_decap_8 FILLER_10_933 ();
 sg13g2_decap_8 FILLER_10_940 ();
 sg13g2_decap_8 FILLER_10_947 ();
 sg13g2_decap_8 FILLER_10_954 ();
 sg13g2_decap_8 FILLER_10_961 ();
 sg13g2_fill_2 FILLER_10_968 ();
 sg13g2_fill_1 FILLER_10_970 ();
 sg13g2_decap_8 FILLER_10_997 ();
 sg13g2_decap_8 FILLER_10_1004 ();
 sg13g2_decap_8 FILLER_10_1047 ();
 sg13g2_decap_8 FILLER_10_1054 ();
 sg13g2_decap_8 FILLER_10_1061 ();
 sg13g2_decap_4 FILLER_10_1068 ();
 sg13g2_fill_2 FILLER_10_1072 ();
 sg13g2_decap_8 FILLER_10_1084 ();
 sg13g2_decap_8 FILLER_10_1091 ();
 sg13g2_decap_4 FILLER_10_1098 ();
 sg13g2_fill_2 FILLER_10_1102 ();
 sg13g2_decap_8 FILLER_10_1107 ();
 sg13g2_fill_2 FILLER_10_1114 ();
 sg13g2_fill_1 FILLER_10_1116 ();
 sg13g2_decap_8 FILLER_10_1125 ();
 sg13g2_decap_8 FILLER_10_1132 ();
 sg13g2_fill_2 FILLER_10_1139 ();
 sg13g2_fill_1 FILLER_10_1141 ();
 sg13g2_fill_2 FILLER_10_1168 ();
 sg13g2_fill_1 FILLER_10_1170 ();
 sg13g2_decap_8 FILLER_10_1181 ();
 sg13g2_decap_8 FILLER_10_1188 ();
 sg13g2_decap_8 FILLER_10_1195 ();
 sg13g2_decap_8 FILLER_10_1202 ();
 sg13g2_decap_8 FILLER_10_1209 ();
 sg13g2_decap_8 FILLER_10_1216 ();
 sg13g2_decap_8 FILLER_10_1223 ();
 sg13g2_decap_8 FILLER_10_1230 ();
 sg13g2_decap_8 FILLER_10_1237 ();
 sg13g2_decap_8 FILLER_10_1244 ();
 sg13g2_fill_2 FILLER_10_1251 ();
 sg13g2_fill_1 FILLER_10_1253 ();
 sg13g2_decap_8 FILLER_10_1258 ();
 sg13g2_decap_8 FILLER_10_1265 ();
 sg13g2_decap_8 FILLER_10_1272 ();
 sg13g2_decap_8 FILLER_10_1279 ();
 sg13g2_decap_8 FILLER_10_1286 ();
 sg13g2_decap_8 FILLER_10_1293 ();
 sg13g2_decap_8 FILLER_10_1323 ();
 sg13g2_decap_8 FILLER_10_1330 ();
 sg13g2_decap_8 FILLER_10_1337 ();
 sg13g2_decap_8 FILLER_10_1344 ();
 sg13g2_decap_8 FILLER_10_1351 ();
 sg13g2_decap_8 FILLER_10_1358 ();
 sg13g2_decap_8 FILLER_10_1365 ();
 sg13g2_decap_8 FILLER_10_1372 ();
 sg13g2_decap_4 FILLER_10_1379 ();
 sg13g2_fill_2 FILLER_10_1383 ();
 sg13g2_decap_8 FILLER_10_1395 ();
 sg13g2_decap_4 FILLER_10_1402 ();
 sg13g2_fill_2 FILLER_10_1406 ();
 sg13g2_decap_8 FILLER_10_1443 ();
 sg13g2_decap_8 FILLER_10_1450 ();
 sg13g2_decap_8 FILLER_10_1457 ();
 sg13g2_decap_8 FILLER_10_1464 ();
 sg13g2_decap_8 FILLER_10_1471 ();
 sg13g2_decap_8 FILLER_10_1478 ();
 sg13g2_decap_8 FILLER_10_1485 ();
 sg13g2_decap_8 FILLER_10_1492 ();
 sg13g2_decap_8 FILLER_10_1499 ();
 sg13g2_decap_4 FILLER_10_1506 ();
 sg13g2_fill_2 FILLER_10_1510 ();
 sg13g2_decap_8 FILLER_10_1527 ();
 sg13g2_decap_8 FILLER_10_1534 ();
 sg13g2_decap_8 FILLER_10_1541 ();
 sg13g2_fill_1 FILLER_10_1548 ();
 sg13g2_fill_2 FILLER_10_1564 ();
 sg13g2_decap_8 FILLER_10_1576 ();
 sg13g2_decap_8 FILLER_10_1583 ();
 sg13g2_decap_8 FILLER_10_1590 ();
 sg13g2_fill_2 FILLER_10_1597 ();
 sg13g2_fill_1 FILLER_10_1599 ();
 sg13g2_decap_8 FILLER_10_1619 ();
 sg13g2_fill_2 FILLER_10_1626 ();
 sg13g2_decap_8 FILLER_10_1637 ();
 sg13g2_decap_8 FILLER_10_1644 ();
 sg13g2_decap_8 FILLER_10_1651 ();
 sg13g2_decap_4 FILLER_10_1658 ();
 sg13g2_fill_1 FILLER_10_1662 ();
 sg13g2_decap_4 FILLER_10_1672 ();
 sg13g2_fill_1 FILLER_10_1676 ();
 sg13g2_decap_4 FILLER_10_1681 ();
 sg13g2_decap_8 FILLER_10_1703 ();
 sg13g2_decap_8 FILLER_10_1710 ();
 sg13g2_decap_8 FILLER_10_1717 ();
 sg13g2_decap_8 FILLER_10_1724 ();
 sg13g2_fill_2 FILLER_10_1731 ();
 sg13g2_fill_1 FILLER_10_1733 ();
 sg13g2_decap_8 FILLER_10_1765 ();
 sg13g2_decap_8 FILLER_10_1772 ();
 sg13g2_decap_4 FILLER_10_1779 ();
 sg13g2_fill_2 FILLER_10_1783 ();
 sg13g2_decap_8 FILLER_10_1800 ();
 sg13g2_decap_8 FILLER_10_1807 ();
 sg13g2_decap_4 FILLER_10_1814 ();
 sg13g2_fill_2 FILLER_10_1837 ();
 sg13g2_fill_1 FILLER_10_1839 ();
 sg13g2_decap_8 FILLER_10_1855 ();
 sg13g2_decap_8 FILLER_10_1862 ();
 sg13g2_decap_8 FILLER_10_1869 ();
 sg13g2_decap_8 FILLER_10_1876 ();
 sg13g2_decap_8 FILLER_10_1888 ();
 sg13g2_decap_8 FILLER_10_1895 ();
 sg13g2_decap_8 FILLER_10_1902 ();
 sg13g2_decap_8 FILLER_10_1909 ();
 sg13g2_fill_2 FILLER_10_1942 ();
 sg13g2_fill_1 FILLER_10_1944 ();
 sg13g2_decap_4 FILLER_10_1948 ();
 sg13g2_fill_1 FILLER_10_1952 ();
 sg13g2_fill_1 FILLER_10_1963 ();
 sg13g2_decap_8 FILLER_10_1974 ();
 sg13g2_decap_4 FILLER_10_1981 ();
 sg13g2_fill_2 FILLER_10_1985 ();
 sg13g2_decap_8 FILLER_10_2023 ();
 sg13g2_decap_8 FILLER_10_2030 ();
 sg13g2_decap_8 FILLER_10_2037 ();
 sg13g2_fill_2 FILLER_10_2044 ();
 sg13g2_fill_1 FILLER_10_2046 ();
 sg13g2_decap_8 FILLER_10_2073 ();
 sg13g2_decap_8 FILLER_10_2080 ();
 sg13g2_decap_8 FILLER_10_2087 ();
 sg13g2_fill_1 FILLER_10_2094 ();
 sg13g2_decap_8 FILLER_10_2121 ();
 sg13g2_decap_8 FILLER_10_2128 ();
 sg13g2_decap_8 FILLER_10_2135 ();
 sg13g2_decap_4 FILLER_10_2142 ();
 sg13g2_decap_8 FILLER_10_2172 ();
 sg13g2_decap_8 FILLER_10_2179 ();
 sg13g2_decap_8 FILLER_10_2186 ();
 sg13g2_fill_1 FILLER_10_2193 ();
 sg13g2_decap_8 FILLER_10_2220 ();
 sg13g2_decap_8 FILLER_10_2227 ();
 sg13g2_decap_4 FILLER_10_2234 ();
 sg13g2_fill_2 FILLER_10_2238 ();
 sg13g2_decap_8 FILLER_10_2276 ();
 sg13g2_decap_8 FILLER_10_2283 ();
 sg13g2_fill_2 FILLER_10_2290 ();
 sg13g2_fill_1 FILLER_10_2292 ();
 sg13g2_decap_8 FILLER_10_2303 ();
 sg13g2_decap_8 FILLER_10_2310 ();
 sg13g2_decap_8 FILLER_10_2317 ();
 sg13g2_decap_8 FILLER_10_2324 ();
 sg13g2_decap_8 FILLER_10_2331 ();
 sg13g2_decap_8 FILLER_10_2338 ();
 sg13g2_decap_4 FILLER_10_2345 ();
 sg13g2_decap_8 FILLER_10_2359 ();
 sg13g2_decap_8 FILLER_10_2366 ();
 sg13g2_decap_8 FILLER_10_2373 ();
 sg13g2_fill_2 FILLER_10_2380 ();
 sg13g2_fill_1 FILLER_10_2382 ();
 sg13g2_decap_8 FILLER_10_2414 ();
 sg13g2_decap_8 FILLER_10_2421 ();
 sg13g2_decap_8 FILLER_10_2428 ();
 sg13g2_decap_8 FILLER_10_2435 ();
 sg13g2_decap_8 FILLER_10_2442 ();
 sg13g2_decap_8 FILLER_10_2449 ();
 sg13g2_decap_8 FILLER_10_2456 ();
 sg13g2_decap_8 FILLER_10_2463 ();
 sg13g2_decap_8 FILLER_10_2470 ();
 sg13g2_decap_8 FILLER_10_2477 ();
 sg13g2_decap_8 FILLER_10_2484 ();
 sg13g2_decap_8 FILLER_10_2491 ();
 sg13g2_decap_8 FILLER_10_2498 ();
 sg13g2_fill_1 FILLER_10_2505 ();
 sg13g2_decap_8 FILLER_10_2516 ();
 sg13g2_decap_8 FILLER_10_2523 ();
 sg13g2_decap_8 FILLER_10_2530 ();
 sg13g2_decap_4 FILLER_10_2537 ();
 sg13g2_fill_2 FILLER_10_2541 ();
 sg13g2_decap_8 FILLER_10_2553 ();
 sg13g2_decap_8 FILLER_10_2560 ();
 sg13g2_decap_8 FILLER_10_2567 ();
 sg13g2_decap_8 FILLER_10_2574 ();
 sg13g2_decap_8 FILLER_10_2581 ();
 sg13g2_decap_8 FILLER_10_2588 ();
 sg13g2_decap_8 FILLER_10_2595 ();
 sg13g2_decap_8 FILLER_10_2602 ();
 sg13g2_fill_2 FILLER_10_2609 ();
 sg13g2_fill_1 FILLER_10_2611 ();
 sg13g2_decap_8 FILLER_10_2622 ();
 sg13g2_decap_8 FILLER_10_2629 ();
 sg13g2_decap_8 FILLER_10_2636 ();
 sg13g2_decap_8 FILLER_10_2643 ();
 sg13g2_decap_8 FILLER_10_2650 ();
 sg13g2_decap_8 FILLER_10_2657 ();
 sg13g2_decap_8 FILLER_10_2664 ();
 sg13g2_decap_8 FILLER_10_2671 ();
 sg13g2_decap_8 FILLER_10_2678 ();
 sg13g2_decap_8 FILLER_10_2685 ();
 sg13g2_decap_4 FILLER_10_2692 ();
 sg13g2_fill_2 FILLER_10_2696 ();
 sg13g2_decap_8 FILLER_10_2708 ();
 sg13g2_decap_8 FILLER_10_2715 ();
 sg13g2_decap_8 FILLER_10_2722 ();
 sg13g2_decap_8 FILLER_10_2729 ();
 sg13g2_decap_8 FILLER_10_2736 ();
 sg13g2_decap_4 FILLER_10_2743 ();
 sg13g2_decap_8 FILLER_10_2773 ();
 sg13g2_decap_8 FILLER_10_2780 ();
 sg13g2_decap_8 FILLER_10_2802 ();
 sg13g2_decap_8 FILLER_10_2809 ();
 sg13g2_decap_8 FILLER_10_2816 ();
 sg13g2_decap_8 FILLER_10_2833 ();
 sg13g2_decap_8 FILLER_10_2840 ();
 sg13g2_decap_8 FILLER_10_2847 ();
 sg13g2_decap_8 FILLER_10_2880 ();
 sg13g2_decap_8 FILLER_10_2887 ();
 sg13g2_fill_2 FILLER_10_2894 ();
 sg13g2_fill_1 FILLER_10_2896 ();
 sg13g2_decap_8 FILLER_10_2928 ();
 sg13g2_decap_8 FILLER_10_2935 ();
 sg13g2_decap_8 FILLER_10_2942 ();
 sg13g2_fill_2 FILLER_10_2949 ();
 sg13g2_fill_1 FILLER_10_2951 ();
 sg13g2_fill_2 FILLER_10_2975 ();
 sg13g2_fill_1 FILLER_10_2977 ();
 sg13g2_decap_8 FILLER_10_2987 ();
 sg13g2_decap_8 FILLER_10_2994 ();
 sg13g2_decap_8 FILLER_10_3001 ();
 sg13g2_decap_8 FILLER_10_3008 ();
 sg13g2_decap_8 FILLER_10_3015 ();
 sg13g2_decap_8 FILLER_10_3022 ();
 sg13g2_fill_2 FILLER_10_3029 ();
 sg13g2_decap_8 FILLER_10_3051 ();
 sg13g2_decap_8 FILLER_10_3058 ();
 sg13g2_decap_8 FILLER_10_3065 ();
 sg13g2_decap_8 FILLER_10_3093 ();
 sg13g2_fill_1 FILLER_10_3100 ();
 sg13g2_fill_2 FILLER_10_3106 ();
 sg13g2_decap_8 FILLER_10_3129 ();
 sg13g2_decap_8 FILLER_10_3136 ();
 sg13g2_decap_8 FILLER_10_3143 ();
 sg13g2_fill_2 FILLER_10_3150 ();
 sg13g2_fill_1 FILLER_10_3152 ();
 sg13g2_decap_8 FILLER_10_3195 ();
 sg13g2_decap_8 FILLER_10_3202 ();
 sg13g2_fill_1 FILLER_10_3209 ();
 sg13g2_decap_8 FILLER_10_3219 ();
 sg13g2_decap_8 FILLER_10_3226 ();
 sg13g2_decap_8 FILLER_10_3233 ();
 sg13g2_decap_4 FILLER_10_3240 ();
 sg13g2_fill_2 FILLER_10_3244 ();
 sg13g2_decap_4 FILLER_10_3256 ();
 sg13g2_decap_8 FILLER_10_3264 ();
 sg13g2_fill_2 FILLER_10_3271 ();
 sg13g2_decap_8 FILLER_10_3292 ();
 sg13g2_decap_8 FILLER_10_3299 ();
 sg13g2_decap_4 FILLER_10_3306 ();
 sg13g2_fill_1 FILLER_10_3310 ();
 sg13g2_decap_8 FILLER_10_3321 ();
 sg13g2_decap_8 FILLER_10_3328 ();
 sg13g2_decap_4 FILLER_10_3335 ();
 sg13g2_fill_2 FILLER_10_3339 ();
 sg13g2_decap_8 FILLER_10_3346 ();
 sg13g2_decap_8 FILLER_10_3353 ();
 sg13g2_decap_8 FILLER_10_3360 ();
 sg13g2_decap_8 FILLER_10_3367 ();
 sg13g2_decap_8 FILLER_10_3374 ();
 sg13g2_decap_4 FILLER_10_3381 ();
 sg13g2_fill_1 FILLER_10_3390 ();
 sg13g2_decap_8 FILLER_10_3396 ();
 sg13g2_decap_8 FILLER_10_3403 ();
 sg13g2_decap_8 FILLER_10_3410 ();
 sg13g2_decap_8 FILLER_10_3417 ();
 sg13g2_decap_8 FILLER_10_3424 ();
 sg13g2_decap_8 FILLER_10_3431 ();
 sg13g2_fill_2 FILLER_10_3438 ();
 sg13g2_decap_8 FILLER_10_3466 ();
 sg13g2_decap_8 FILLER_10_3473 ();
 sg13g2_decap_8 FILLER_10_3480 ();
 sg13g2_decap_8 FILLER_10_3487 ();
 sg13g2_decap_8 FILLER_10_3494 ();
 sg13g2_decap_8 FILLER_10_3501 ();
 sg13g2_decap_8 FILLER_10_3508 ();
 sg13g2_decap_8 FILLER_10_3515 ();
 sg13g2_decap_8 FILLER_10_3522 ();
 sg13g2_decap_8 FILLER_10_3529 ();
 sg13g2_decap_8 FILLER_10_3536 ();
 sg13g2_decap_8 FILLER_10_3543 ();
 sg13g2_decap_8 FILLER_10_3550 ();
 sg13g2_decap_8 FILLER_10_3557 ();
 sg13g2_decap_8 FILLER_10_3564 ();
 sg13g2_decap_8 FILLER_10_3571 ();
 sg13g2_fill_2 FILLER_10_3578 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_4 FILLER_11_7 ();
 sg13g2_fill_2 FILLER_11_11 ();
 sg13g2_decap_8 FILLER_11_52 ();
 sg13g2_fill_2 FILLER_11_59 ();
 sg13g2_fill_1 FILLER_11_95 ();
 sg13g2_decap_8 FILLER_11_101 ();
 sg13g2_decap_8 FILLER_11_108 ();
 sg13g2_fill_2 FILLER_11_115 ();
 sg13g2_decap_8 FILLER_11_125 ();
 sg13g2_decap_8 FILLER_11_132 ();
 sg13g2_decap_8 FILLER_11_139 ();
 sg13g2_decap_4 FILLER_11_146 ();
 sg13g2_fill_2 FILLER_11_155 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_fill_2 FILLER_11_203 ();
 sg13g2_fill_1 FILLER_11_205 ();
 sg13g2_fill_2 FILLER_11_222 ();
 sg13g2_fill_2 FILLER_11_237 ();
 sg13g2_decap_8 FILLER_11_243 ();
 sg13g2_decap_8 FILLER_11_250 ();
 sg13g2_decap_8 FILLER_11_257 ();
 sg13g2_decap_8 FILLER_11_264 ();
 sg13g2_decap_8 FILLER_11_271 ();
 sg13g2_decap_8 FILLER_11_278 ();
 sg13g2_decap_8 FILLER_11_285 ();
 sg13g2_decap_8 FILLER_11_292 ();
 sg13g2_fill_1 FILLER_11_299 ();
 sg13g2_decap_8 FILLER_11_304 ();
 sg13g2_decap_8 FILLER_11_311 ();
 sg13g2_fill_1 FILLER_11_318 ();
 sg13g2_fill_1 FILLER_11_324 ();
 sg13g2_fill_2 FILLER_11_338 ();
 sg13g2_fill_1 FILLER_11_340 ();
 sg13g2_decap_8 FILLER_11_348 ();
 sg13g2_decap_8 FILLER_11_355 ();
 sg13g2_decap_8 FILLER_11_362 ();
 sg13g2_decap_8 FILLER_11_369 ();
 sg13g2_decap_4 FILLER_11_376 ();
 sg13g2_fill_2 FILLER_11_380 ();
 sg13g2_decap_8 FILLER_11_389 ();
 sg13g2_decap_8 FILLER_11_396 ();
 sg13g2_decap_4 FILLER_11_403 ();
 sg13g2_fill_2 FILLER_11_407 ();
 sg13g2_decap_8 FILLER_11_417 ();
 sg13g2_decap_8 FILLER_11_424 ();
 sg13g2_decap_8 FILLER_11_431 ();
 sg13g2_decap_8 FILLER_11_438 ();
 sg13g2_decap_8 FILLER_11_445 ();
 sg13g2_fill_2 FILLER_11_452 ();
 sg13g2_fill_1 FILLER_11_454 ();
 sg13g2_decap_8 FILLER_11_459 ();
 sg13g2_decap_8 FILLER_11_466 ();
 sg13g2_decap_8 FILLER_11_473 ();
 sg13g2_decap_4 FILLER_11_480 ();
 sg13g2_fill_2 FILLER_11_484 ();
 sg13g2_decap_8 FILLER_11_497 ();
 sg13g2_decap_8 FILLER_11_504 ();
 sg13g2_decap_8 FILLER_11_511 ();
 sg13g2_decap_8 FILLER_11_518 ();
 sg13g2_decap_8 FILLER_11_525 ();
 sg13g2_decap_8 FILLER_11_532 ();
 sg13g2_decap_8 FILLER_11_539 ();
 sg13g2_decap_8 FILLER_11_546 ();
 sg13g2_decap_8 FILLER_11_553 ();
 sg13g2_decap_8 FILLER_11_560 ();
 sg13g2_decap_8 FILLER_11_567 ();
 sg13g2_fill_2 FILLER_11_574 ();
 sg13g2_decap_8 FILLER_11_586 ();
 sg13g2_decap_8 FILLER_11_593 ();
 sg13g2_decap_8 FILLER_11_600 ();
 sg13g2_decap_8 FILLER_11_607 ();
 sg13g2_decap_8 FILLER_11_614 ();
 sg13g2_decap_8 FILLER_11_621 ();
 sg13g2_decap_4 FILLER_11_628 ();
 sg13g2_fill_1 FILLER_11_632 ();
 sg13g2_decap_8 FILLER_11_646 ();
 sg13g2_decap_8 FILLER_11_653 ();
 sg13g2_decap_8 FILLER_11_660 ();
 sg13g2_fill_2 FILLER_11_667 ();
 sg13g2_decap_8 FILLER_11_695 ();
 sg13g2_decap_8 FILLER_11_702 ();
 sg13g2_fill_1 FILLER_11_709 ();
 sg13g2_decap_4 FILLER_11_736 ();
 sg13g2_fill_2 FILLER_11_740 ();
 sg13g2_decap_8 FILLER_11_747 ();
 sg13g2_decap_8 FILLER_11_754 ();
 sg13g2_decap_8 FILLER_11_761 ();
 sg13g2_decap_8 FILLER_11_789 ();
 sg13g2_decap_8 FILLER_11_796 ();
 sg13g2_decap_8 FILLER_11_803 ();
 sg13g2_decap_8 FILLER_11_810 ();
 sg13g2_decap_4 FILLER_11_817 ();
 sg13g2_fill_2 FILLER_11_821 ();
 sg13g2_decap_8 FILLER_11_849 ();
 sg13g2_decap_8 FILLER_11_856 ();
 sg13g2_decap_8 FILLER_11_863 ();
 sg13g2_decap_8 FILLER_11_870 ();
 sg13g2_decap_4 FILLER_11_877 ();
 sg13g2_decap_8 FILLER_11_907 ();
 sg13g2_decap_8 FILLER_11_914 ();
 sg13g2_decap_8 FILLER_11_921 ();
 sg13g2_decap_8 FILLER_11_928 ();
 sg13g2_decap_8 FILLER_11_935 ();
 sg13g2_decap_8 FILLER_11_942 ();
 sg13g2_decap_8 FILLER_11_949 ();
 sg13g2_decap_8 FILLER_11_956 ();
 sg13g2_decap_8 FILLER_11_963 ();
 sg13g2_decap_8 FILLER_11_970 ();
 sg13g2_fill_2 FILLER_11_977 ();
 sg13g2_fill_1 FILLER_11_979 ();
 sg13g2_decap_8 FILLER_11_1016 ();
 sg13g2_decap_8 FILLER_11_1023 ();
 sg13g2_fill_2 FILLER_11_1030 ();
 sg13g2_decap_8 FILLER_11_1058 ();
 sg13g2_fill_1 FILLER_11_1065 ();
 sg13g2_decap_8 FILLER_11_1092 ();
 sg13g2_decap_8 FILLER_11_1099 ();
 sg13g2_decap_8 FILLER_11_1106 ();
 sg13g2_decap_8 FILLER_11_1113 ();
 sg13g2_decap_8 FILLER_11_1120 ();
 sg13g2_decap_8 FILLER_11_1127 ();
 sg13g2_decap_8 FILLER_11_1134 ();
 sg13g2_decap_4 FILLER_11_1141 ();
 sg13g2_fill_2 FILLER_11_1153 ();
 sg13g2_decap_8 FILLER_11_1181 ();
 sg13g2_decap_8 FILLER_11_1188 ();
 sg13g2_decap_8 FILLER_11_1195 ();
 sg13g2_fill_2 FILLER_11_1202 ();
 sg13g2_fill_1 FILLER_11_1204 ();
 sg13g2_fill_1 FILLER_11_1211 ();
 sg13g2_decap_8 FILLER_11_1224 ();
 sg13g2_decap_8 FILLER_11_1231 ();
 sg13g2_fill_2 FILLER_11_1238 ();
 sg13g2_decap_8 FILLER_11_1279 ();
 sg13g2_decap_8 FILLER_11_1286 ();
 sg13g2_decap_4 FILLER_11_1293 ();
 sg13g2_fill_2 FILLER_11_1297 ();
 sg13g2_decap_8 FILLER_11_1304 ();
 sg13g2_fill_1 FILLER_11_1311 ();
 sg13g2_decap_8 FILLER_11_1315 ();
 sg13g2_decap_8 FILLER_11_1322 ();
 sg13g2_decap_8 FILLER_11_1329 ();
 sg13g2_decap_8 FILLER_11_1336 ();
 sg13g2_decap_8 FILLER_11_1343 ();
 sg13g2_fill_1 FILLER_11_1350 ();
 sg13g2_decap_4 FILLER_11_1380 ();
 sg13g2_fill_1 FILLER_11_1384 ();
 sg13g2_fill_2 FILLER_11_1403 ();
 sg13g2_decap_8 FILLER_11_1435 ();
 sg13g2_decap_8 FILLER_11_1442 ();
 sg13g2_decap_8 FILLER_11_1449 ();
 sg13g2_decap_8 FILLER_11_1456 ();
 sg13g2_decap_8 FILLER_11_1463 ();
 sg13g2_decap_8 FILLER_11_1470 ();
 sg13g2_decap_8 FILLER_11_1477 ();
 sg13g2_decap_8 FILLER_11_1484 ();
 sg13g2_decap_8 FILLER_11_1491 ();
 sg13g2_decap_8 FILLER_11_1498 ();
 sg13g2_decap_4 FILLER_11_1505 ();
 sg13g2_fill_1 FILLER_11_1509 ();
 sg13g2_fill_2 FILLER_11_1525 ();
 sg13g2_decap_8 FILLER_11_1532 ();
 sg13g2_decap_8 FILLER_11_1539 ();
 sg13g2_decap_8 FILLER_11_1546 ();
 sg13g2_decap_4 FILLER_11_1553 ();
 sg13g2_decap_8 FILLER_11_1562 ();
 sg13g2_decap_8 FILLER_11_1569 ();
 sg13g2_fill_2 FILLER_11_1576 ();
 sg13g2_fill_1 FILLER_11_1578 ();
 sg13g2_decap_8 FILLER_11_1600 ();
 sg13g2_fill_1 FILLER_11_1607 ();
 sg13g2_decap_8 FILLER_11_1639 ();
 sg13g2_decap_8 FILLER_11_1646 ();
 sg13g2_decap_8 FILLER_11_1653 ();
 sg13g2_decap_8 FILLER_11_1660 ();
 sg13g2_decap_8 FILLER_11_1667 ();
 sg13g2_decap_4 FILLER_11_1674 ();
 sg13g2_fill_2 FILLER_11_1678 ();
 sg13g2_decap_8 FILLER_11_1688 ();
 sg13g2_decap_8 FILLER_11_1695 ();
 sg13g2_decap_8 FILLER_11_1702 ();
 sg13g2_decap_4 FILLER_11_1709 ();
 sg13g2_fill_2 FILLER_11_1713 ();
 sg13g2_decap_4 FILLER_11_1720 ();
 sg13g2_fill_1 FILLER_11_1724 ();
 sg13g2_fill_2 FILLER_11_1746 ();
 sg13g2_fill_1 FILLER_11_1748 ();
 sg13g2_decap_8 FILLER_11_1754 ();
 sg13g2_decap_8 FILLER_11_1761 ();
 sg13g2_decap_8 FILLER_11_1768 ();
 sg13g2_decap_8 FILLER_11_1810 ();
 sg13g2_decap_8 FILLER_11_1817 ();
 sg13g2_decap_4 FILLER_11_1824 ();
 sg13g2_fill_2 FILLER_11_1828 ();
 sg13g2_decap_8 FILLER_11_1860 ();
 sg13g2_decap_8 FILLER_11_1867 ();
 sg13g2_decap_8 FILLER_11_1874 ();
 sg13g2_decap_8 FILLER_11_1881 ();
 sg13g2_decap_8 FILLER_11_1888 ();
 sg13g2_decap_8 FILLER_11_1895 ();
 sg13g2_decap_8 FILLER_11_1902 ();
 sg13g2_decap_8 FILLER_11_1909 ();
 sg13g2_decap_8 FILLER_11_1926 ();
 sg13g2_decap_8 FILLER_11_1933 ();
 sg13g2_decap_8 FILLER_11_1940 ();
 sg13g2_decap_8 FILLER_11_1947 ();
 sg13g2_decap_8 FILLER_11_1954 ();
 sg13g2_decap_8 FILLER_11_1961 ();
 sg13g2_decap_8 FILLER_11_1968 ();
 sg13g2_decap_8 FILLER_11_1975 ();
 sg13g2_fill_2 FILLER_11_1982 ();
 sg13g2_fill_1 FILLER_11_1984 ();
 sg13g2_decap_4 FILLER_11_1995 ();
 sg13g2_decap_8 FILLER_11_2009 ();
 sg13g2_decap_8 FILLER_11_2016 ();
 sg13g2_decap_8 FILLER_11_2023 ();
 sg13g2_decap_8 FILLER_11_2030 ();
 sg13g2_decap_8 FILLER_11_2037 ();
 sg13g2_decap_8 FILLER_11_2044 ();
 sg13g2_decap_4 FILLER_11_2051 ();
 sg13g2_decap_8 FILLER_11_2065 ();
 sg13g2_decap_8 FILLER_11_2072 ();
 sg13g2_decap_8 FILLER_11_2114 ();
 sg13g2_decap_8 FILLER_11_2121 ();
 sg13g2_decap_4 FILLER_11_2128 ();
 sg13g2_decap_8 FILLER_11_2168 ();
 sg13g2_decap_8 FILLER_11_2175 ();
 sg13g2_decap_8 FILLER_11_2182 ();
 sg13g2_decap_4 FILLER_11_2189 ();
 sg13g2_fill_1 FILLER_11_2193 ();
 sg13g2_decap_8 FILLER_11_2208 ();
 sg13g2_decap_4 FILLER_11_2215 ();
 sg13g2_fill_1 FILLER_11_2219 ();
 sg13g2_decap_8 FILLER_11_2230 ();
 sg13g2_decap_8 FILLER_11_2263 ();
 sg13g2_decap_4 FILLER_11_2296 ();
 sg13g2_decap_8 FILLER_11_2334 ();
 sg13g2_fill_2 FILLER_11_2341 ();
 sg13g2_fill_1 FILLER_11_2343 ();
 sg13g2_decap_8 FILLER_11_2370 ();
 sg13g2_decap_8 FILLER_11_2377 ();
 sg13g2_decap_8 FILLER_11_2384 ();
 sg13g2_decap_8 FILLER_11_2391 ();
 sg13g2_decap_4 FILLER_11_2398 ();
 sg13g2_decap_8 FILLER_11_2416 ();
 sg13g2_decap_8 FILLER_11_2423 ();
 sg13g2_fill_2 FILLER_11_2430 ();
 sg13g2_fill_1 FILLER_11_2432 ();
 sg13g2_fill_2 FILLER_11_2459 ();
 sg13g2_fill_1 FILLER_11_2461 ();
 sg13g2_decap_4 FILLER_11_2472 ();
 sg13g2_fill_1 FILLER_11_2476 ();
 sg13g2_decap_8 FILLER_11_2487 ();
 sg13g2_fill_2 FILLER_11_2494 ();
 sg13g2_fill_1 FILLER_11_2496 ();
 sg13g2_decap_8 FILLER_11_2523 ();
 sg13g2_decap_8 FILLER_11_2530 ();
 sg13g2_fill_2 FILLER_11_2537 ();
 sg13g2_fill_1 FILLER_11_2539 ();
 sg13g2_decap_8 FILLER_11_2576 ();
 sg13g2_decap_8 FILLER_11_2583 ();
 sg13g2_fill_1 FILLER_11_2590 ();
 sg13g2_decap_8 FILLER_11_2627 ();
 sg13g2_decap_8 FILLER_11_2634 ();
 sg13g2_decap_8 FILLER_11_2641 ();
 sg13g2_decap_8 FILLER_11_2648 ();
 sg13g2_decap_8 FILLER_11_2681 ();
 sg13g2_decap_8 FILLER_11_2688 ();
 sg13g2_fill_2 FILLER_11_2695 ();
 sg13g2_fill_1 FILLER_11_2697 ();
 sg13g2_decap_8 FILLER_11_2750 ();
 sg13g2_decap_8 FILLER_11_2757 ();
 sg13g2_decap_8 FILLER_11_2764 ();
 sg13g2_decap_8 FILLER_11_2771 ();
 sg13g2_decap_4 FILLER_11_2778 ();
 sg13g2_fill_2 FILLER_11_2811 ();
 sg13g2_fill_1 FILLER_11_2813 ();
 sg13g2_fill_2 FILLER_11_2845 ();
 sg13g2_fill_1 FILLER_11_2847 ();
 sg13g2_decap_8 FILLER_11_2853 ();
 sg13g2_fill_2 FILLER_11_2860 ();
 sg13g2_fill_1 FILLER_11_2862 ();
 sg13g2_decap_8 FILLER_11_2878 ();
 sg13g2_fill_1 FILLER_11_2895 ();
 sg13g2_decap_8 FILLER_11_2911 ();
 sg13g2_decap_8 FILLER_11_2918 ();
 sg13g2_decap_8 FILLER_11_2925 ();
 sg13g2_decap_8 FILLER_11_2932 ();
 sg13g2_decap_8 FILLER_11_2939 ();
 sg13g2_decap_8 FILLER_11_2946 ();
 sg13g2_decap_8 FILLER_11_2953 ();
 sg13g2_decap_8 FILLER_11_2960 ();
 sg13g2_decap_8 FILLER_11_2967 ();
 sg13g2_decap_8 FILLER_11_2974 ();
 sg13g2_decap_8 FILLER_11_2981 ();
 sg13g2_decap_8 FILLER_11_2988 ();
 sg13g2_decap_8 FILLER_11_2995 ();
 sg13g2_decap_8 FILLER_11_3002 ();
 sg13g2_decap_8 FILLER_11_3009 ();
 sg13g2_decap_8 FILLER_11_3016 ();
 sg13g2_decap_8 FILLER_11_3023 ();
 sg13g2_decap_8 FILLER_11_3030 ();
 sg13g2_fill_2 FILLER_11_3037 ();
 sg13g2_decap_8 FILLER_11_3044 ();
 sg13g2_decap_8 FILLER_11_3051 ();
 sg13g2_decap_8 FILLER_11_3058 ();
 sg13g2_decap_8 FILLER_11_3065 ();
 sg13g2_decap_8 FILLER_11_3072 ();
 sg13g2_decap_8 FILLER_11_3079 ();
 sg13g2_decap_8 FILLER_11_3086 ();
 sg13g2_decap_8 FILLER_11_3093 ();
 sg13g2_decap_8 FILLER_11_3100 ();
 sg13g2_fill_1 FILLER_11_3107 ();
 sg13g2_decap_8 FILLER_11_3128 ();
 sg13g2_decap_8 FILLER_11_3135 ();
 sg13g2_decap_4 FILLER_11_3142 ();
 sg13g2_decap_8 FILLER_11_3151 ();
 sg13g2_decap_4 FILLER_11_3158 ();
 sg13g2_fill_1 FILLER_11_3167 ();
 sg13g2_decap_8 FILLER_11_3188 ();
 sg13g2_decap_8 FILLER_11_3195 ();
 sg13g2_decap_8 FILLER_11_3202 ();
 sg13g2_decap_8 FILLER_11_3209 ();
 sg13g2_decap_8 FILLER_11_3216 ();
 sg13g2_decap_8 FILLER_11_3223 ();
 sg13g2_decap_8 FILLER_11_3230 ();
 sg13g2_decap_4 FILLER_11_3237 ();
 sg13g2_decap_4 FILLER_11_3266 ();
 sg13g2_fill_2 FILLER_11_3270 ();
 sg13g2_decap_8 FILLER_11_3281 ();
 sg13g2_fill_2 FILLER_11_3288 ();
 sg13g2_decap_8 FILLER_11_3300 ();
 sg13g2_decap_8 FILLER_11_3307 ();
 sg13g2_decap_8 FILLER_11_3314 ();
 sg13g2_decap_8 FILLER_11_3321 ();
 sg13g2_decap_8 FILLER_11_3328 ();
 sg13g2_decap_8 FILLER_11_3335 ();
 sg13g2_fill_2 FILLER_11_3342 ();
 sg13g2_decap_8 FILLER_11_3347 ();
 sg13g2_decap_8 FILLER_11_3354 ();
 sg13g2_decap_4 FILLER_11_3361 ();
 sg13g2_fill_1 FILLER_11_3365 ();
 sg13g2_fill_2 FILLER_11_3376 ();
 sg13g2_decap_8 FILLER_11_3412 ();
 sg13g2_decap_8 FILLER_11_3419 ();
 sg13g2_decap_8 FILLER_11_3426 ();
 sg13g2_decap_8 FILLER_11_3459 ();
 sg13g2_decap_8 FILLER_11_3466 ();
 sg13g2_decap_8 FILLER_11_3473 ();
 sg13g2_decap_8 FILLER_11_3480 ();
 sg13g2_decap_8 FILLER_11_3487 ();
 sg13g2_decap_8 FILLER_11_3494 ();
 sg13g2_decap_8 FILLER_11_3501 ();
 sg13g2_decap_8 FILLER_11_3508 ();
 sg13g2_decap_8 FILLER_11_3515 ();
 sg13g2_decap_8 FILLER_11_3522 ();
 sg13g2_decap_8 FILLER_11_3529 ();
 sg13g2_decap_8 FILLER_11_3536 ();
 sg13g2_decap_8 FILLER_11_3543 ();
 sg13g2_decap_8 FILLER_11_3550 ();
 sg13g2_decap_8 FILLER_11_3557 ();
 sg13g2_decap_8 FILLER_11_3564 ();
 sg13g2_decap_8 FILLER_11_3571 ();
 sg13g2_fill_2 FILLER_11_3578 ();
 sg13g2_fill_2 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_47 ();
 sg13g2_fill_2 FILLER_12_54 ();
 sg13g2_fill_1 FILLER_12_56 ();
 sg13g2_fill_2 FILLER_12_76 ();
 sg13g2_fill_1 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_132 ();
 sg13g2_decap_8 FILLER_12_139 ();
 sg13g2_fill_1 FILLER_12_146 ();
 sg13g2_decap_8 FILLER_12_186 ();
 sg13g2_decap_8 FILLER_12_193 ();
 sg13g2_fill_2 FILLER_12_226 ();
 sg13g2_decap_8 FILLER_12_250 ();
 sg13g2_decap_8 FILLER_12_257 ();
 sg13g2_decap_4 FILLER_12_264 ();
 sg13g2_decap_4 FILLER_12_271 ();
 sg13g2_fill_2 FILLER_12_275 ();
 sg13g2_decap_8 FILLER_12_282 ();
 sg13g2_decap_8 FILLER_12_289 ();
 sg13g2_decap_8 FILLER_12_296 ();
 sg13g2_decap_8 FILLER_12_303 ();
 sg13g2_decap_8 FILLER_12_310 ();
 sg13g2_decap_8 FILLER_12_317 ();
 sg13g2_decap_4 FILLER_12_324 ();
 sg13g2_fill_1 FILLER_12_332 ();
 sg13g2_fill_1 FILLER_12_337 ();
 sg13g2_decap_8 FILLER_12_342 ();
 sg13g2_decap_8 FILLER_12_349 ();
 sg13g2_decap_8 FILLER_12_356 ();
 sg13g2_decap_8 FILLER_12_363 ();
 sg13g2_decap_4 FILLER_12_370 ();
 sg13g2_fill_2 FILLER_12_374 ();
 sg13g2_decap_8 FILLER_12_381 ();
 sg13g2_decap_8 FILLER_12_388 ();
 sg13g2_decap_4 FILLER_12_395 ();
 sg13g2_decap_8 FILLER_12_422 ();
 sg13g2_decap_8 FILLER_12_429 ();
 sg13g2_decap_4 FILLER_12_436 ();
 sg13g2_decap_8 FILLER_12_445 ();
 sg13g2_decap_8 FILLER_12_452 ();
 sg13g2_decap_8 FILLER_12_459 ();
 sg13g2_decap_8 FILLER_12_466 ();
 sg13g2_decap_8 FILLER_12_473 ();
 sg13g2_decap_4 FILLER_12_480 ();
 sg13g2_fill_2 FILLER_12_484 ();
 sg13g2_decap_8 FILLER_12_512 ();
 sg13g2_decap_8 FILLER_12_519 ();
 sg13g2_decap_8 FILLER_12_526 ();
 sg13g2_decap_8 FILLER_12_533 ();
 sg13g2_fill_2 FILLER_12_540 ();
 sg13g2_decap_8 FILLER_12_547 ();
 sg13g2_decap_8 FILLER_12_554 ();
 sg13g2_decap_8 FILLER_12_561 ();
 sg13g2_decap_8 FILLER_12_568 ();
 sg13g2_decap_8 FILLER_12_575 ();
 sg13g2_decap_8 FILLER_12_582 ();
 sg13g2_decap_8 FILLER_12_589 ();
 sg13g2_decap_8 FILLER_12_596 ();
 sg13g2_decap_8 FILLER_12_603 ();
 sg13g2_decap_8 FILLER_12_610 ();
 sg13g2_decap_8 FILLER_12_617 ();
 sg13g2_decap_4 FILLER_12_624 ();
 sg13g2_decap_8 FILLER_12_654 ();
 sg13g2_decap_8 FILLER_12_661 ();
 sg13g2_decap_8 FILLER_12_668 ();
 sg13g2_decap_8 FILLER_12_675 ();
 sg13g2_decap_8 FILLER_12_682 ();
 sg13g2_decap_8 FILLER_12_689 ();
 sg13g2_decap_8 FILLER_12_696 ();
 sg13g2_decap_8 FILLER_12_703 ();
 sg13g2_decap_4 FILLER_12_710 ();
 sg13g2_fill_2 FILLER_12_714 ();
 sg13g2_decap_8 FILLER_12_726 ();
 sg13g2_decap_8 FILLER_12_754 ();
 sg13g2_fill_1 FILLER_12_761 ();
 sg13g2_decap_8 FILLER_12_798 ();
 sg13g2_decap_8 FILLER_12_805 ();
 sg13g2_decap_8 FILLER_12_812 ();
 sg13g2_decap_4 FILLER_12_824 ();
 sg13g2_fill_2 FILLER_12_828 ();
 sg13g2_decap_8 FILLER_12_835 ();
 sg13g2_decap_8 FILLER_12_842 ();
 sg13g2_decap_8 FILLER_12_849 ();
 sg13g2_decap_8 FILLER_12_856 ();
 sg13g2_decap_8 FILLER_12_863 ();
 sg13g2_decap_8 FILLER_12_870 ();
 sg13g2_decap_8 FILLER_12_877 ();
 sg13g2_decap_8 FILLER_12_910 ();
 sg13g2_fill_1 FILLER_12_917 ();
 sg13g2_decap_8 FILLER_12_944 ();
 sg13g2_decap_8 FILLER_12_951 ();
 sg13g2_decap_8 FILLER_12_958 ();
 sg13g2_fill_2 FILLER_12_965 ();
 sg13g2_decap_8 FILLER_12_998 ();
 sg13g2_decap_8 FILLER_12_1005 ();
 sg13g2_decap_8 FILLER_12_1012 ();
 sg13g2_decap_8 FILLER_12_1019 ();
 sg13g2_decap_8 FILLER_12_1026 ();
 sg13g2_decap_8 FILLER_12_1033 ();
 sg13g2_decap_8 FILLER_12_1057 ();
 sg13g2_fill_1 FILLER_12_1064 ();
 sg13g2_decap_8 FILLER_12_1082 ();
 sg13g2_decap_8 FILLER_12_1089 ();
 sg13g2_decap_8 FILLER_12_1096 ();
 sg13g2_fill_1 FILLER_12_1103 ();
 sg13g2_decap_4 FILLER_12_1112 ();
 sg13g2_fill_2 FILLER_12_1116 ();
 sg13g2_decap_8 FILLER_12_1126 ();
 sg13g2_decap_8 FILLER_12_1133 ();
 sg13g2_decap_4 FILLER_12_1140 ();
 sg13g2_fill_1 FILLER_12_1144 ();
 sg13g2_decap_8 FILLER_12_1155 ();
 sg13g2_decap_8 FILLER_12_1162 ();
 sg13g2_decap_8 FILLER_12_1169 ();
 sg13g2_fill_1 FILLER_12_1176 ();
 sg13g2_decap_8 FILLER_12_1182 ();
 sg13g2_fill_2 FILLER_12_1189 ();
 sg13g2_fill_1 FILLER_12_1191 ();
 sg13g2_fill_2 FILLER_12_1218 ();
 sg13g2_fill_1 FILLER_12_1220 ();
 sg13g2_decap_8 FILLER_12_1230 ();
 sg13g2_decap_4 FILLER_12_1237 ();
 sg13g2_fill_2 FILLER_12_1288 ();
 sg13g2_fill_1 FILLER_12_1290 ();
 sg13g2_decap_8 FILLER_12_1327 ();
 sg13g2_fill_2 FILLER_12_1334 ();
 sg13g2_decap_8 FILLER_12_1346 ();
 sg13g2_decap_8 FILLER_12_1353 ();
 sg13g2_decap_8 FILLER_12_1360 ();
 sg13g2_decap_8 FILLER_12_1367 ();
 sg13g2_decap_8 FILLER_12_1374 ();
 sg13g2_decap_4 FILLER_12_1381 ();
 sg13g2_decap_8 FILLER_12_1394 ();
 sg13g2_fill_2 FILLER_12_1410 ();
 sg13g2_fill_1 FILLER_12_1412 ();
 sg13g2_decap_8 FILLER_12_1417 ();
 sg13g2_decap_8 FILLER_12_1424 ();
 sg13g2_fill_2 FILLER_12_1444 ();
 sg13g2_fill_1 FILLER_12_1446 ();
 sg13g2_decap_8 FILLER_12_1457 ();
 sg13g2_decap_8 FILLER_12_1464 ();
 sg13g2_decap_8 FILLER_12_1471 ();
 sg13g2_decap_8 FILLER_12_1478 ();
 sg13g2_decap_8 FILLER_12_1485 ();
 sg13g2_fill_2 FILLER_12_1492 ();
 sg13g2_decap_4 FILLER_12_1504 ();
 sg13g2_fill_1 FILLER_12_1508 ();
 sg13g2_decap_8 FILLER_12_1528 ();
 sg13g2_decap_8 FILLER_12_1535 ();
 sg13g2_decap_8 FILLER_12_1542 ();
 sg13g2_decap_8 FILLER_12_1549 ();
 sg13g2_decap_8 FILLER_12_1556 ();
 sg13g2_decap_8 FILLER_12_1563 ();
 sg13g2_fill_1 FILLER_12_1570 ();
 sg13g2_decap_8 FILLER_12_1609 ();
 sg13g2_decap_8 FILLER_12_1616 ();
 sg13g2_decap_8 FILLER_12_1623 ();
 sg13g2_decap_8 FILLER_12_1630 ();
 sg13g2_decap_8 FILLER_12_1637 ();
 sg13g2_decap_8 FILLER_12_1644 ();
 sg13g2_decap_8 FILLER_12_1651 ();
 sg13g2_decap_8 FILLER_12_1658 ();
 sg13g2_decap_8 FILLER_12_1665 ();
 sg13g2_decap_8 FILLER_12_1672 ();
 sg13g2_decap_8 FILLER_12_1679 ();
 sg13g2_decap_8 FILLER_12_1686 ();
 sg13g2_decap_8 FILLER_12_1693 ();
 sg13g2_decap_8 FILLER_12_1700 ();
 sg13g2_decap_4 FILLER_12_1707 ();
 sg13g2_fill_2 FILLER_12_1711 ();
 sg13g2_decap_4 FILLER_12_1739 ();
 sg13g2_fill_1 FILLER_12_1743 ();
 sg13g2_decap_8 FILLER_12_1749 ();
 sg13g2_decap_8 FILLER_12_1756 ();
 sg13g2_decap_8 FILLER_12_1763 ();
 sg13g2_decap_8 FILLER_12_1770 ();
 sg13g2_decap_4 FILLER_12_1777 ();
 sg13g2_fill_1 FILLER_12_1781 ();
 sg13g2_decap_4 FILLER_12_1785 ();
 sg13g2_fill_1 FILLER_12_1789 ();
 sg13g2_decap_8 FILLER_12_1804 ();
 sg13g2_decap_8 FILLER_12_1811 ();
 sg13g2_decap_8 FILLER_12_1818 ();
 sg13g2_decap_4 FILLER_12_1825 ();
 sg13g2_fill_1 FILLER_12_1829 ();
 sg13g2_fill_2 FILLER_12_1835 ();
 sg13g2_decap_8 FILLER_12_1851 ();
 sg13g2_decap_8 FILLER_12_1858 ();
 sg13g2_decap_8 FILLER_12_1865 ();
 sg13g2_fill_2 FILLER_12_1872 ();
 sg13g2_fill_1 FILLER_12_1874 ();
 sg13g2_decap_8 FILLER_12_1885 ();
 sg13g2_decap_8 FILLER_12_1892 ();
 sg13g2_decap_8 FILLER_12_1899 ();
 sg13g2_decap_8 FILLER_12_1906 ();
 sg13g2_decap_8 FILLER_12_1913 ();
 sg13g2_decap_8 FILLER_12_1920 ();
 sg13g2_decap_8 FILLER_12_1927 ();
 sg13g2_decap_8 FILLER_12_1934 ();
 sg13g2_decap_8 FILLER_12_1941 ();
 sg13g2_decap_8 FILLER_12_1951 ();
 sg13g2_decap_8 FILLER_12_1958 ();
 sg13g2_decap_8 FILLER_12_1965 ();
 sg13g2_decap_8 FILLER_12_1972 ();
 sg13g2_decap_8 FILLER_12_1979 ();
 sg13g2_decap_4 FILLER_12_1986 ();
 sg13g2_fill_2 FILLER_12_1990 ();
 sg13g2_decap_8 FILLER_12_2044 ();
 sg13g2_fill_2 FILLER_12_2051 ();
 sg13g2_decap_8 FILLER_12_2063 ();
 sg13g2_decap_8 FILLER_12_2070 ();
 sg13g2_decap_8 FILLER_12_2077 ();
 sg13g2_decap_8 FILLER_12_2094 ();
 sg13g2_decap_8 FILLER_12_2101 ();
 sg13g2_decap_4 FILLER_12_2108 ();
 sg13g2_fill_1 FILLER_12_2112 ();
 sg13g2_decap_8 FILLER_12_2116 ();
 sg13g2_decap_8 FILLER_12_2123 ();
 sg13g2_decap_8 FILLER_12_2130 ();
 sg13g2_decap_8 FILLER_12_2147 ();
 sg13g2_decap_8 FILLER_12_2154 ();
 sg13g2_decap_8 FILLER_12_2161 ();
 sg13g2_decap_8 FILLER_12_2168 ();
 sg13g2_fill_1 FILLER_12_2175 ();
 sg13g2_decap_8 FILLER_12_2181 ();
 sg13g2_fill_1 FILLER_12_2188 ();
 sg13g2_decap_4 FILLER_12_2215 ();
 sg13g2_fill_2 FILLER_12_2219 ();
 sg13g2_decap_8 FILLER_12_2225 ();
 sg13g2_decap_8 FILLER_12_2232 ();
 sg13g2_decap_8 FILLER_12_2239 ();
 sg13g2_fill_1 FILLER_12_2246 ();
 sg13g2_decap_8 FILLER_12_2257 ();
 sg13g2_decap_8 FILLER_12_2264 ();
 sg13g2_decap_8 FILLER_12_2271 ();
 sg13g2_decap_8 FILLER_12_2278 ();
 sg13g2_decap_4 FILLER_12_2285 ();
 sg13g2_fill_2 FILLER_12_2289 ();
 sg13g2_decap_8 FILLER_12_2296 ();
 sg13g2_fill_2 FILLER_12_2303 ();
 sg13g2_fill_1 FILLER_12_2305 ();
 sg13g2_decap_4 FILLER_12_2316 ();
 sg13g2_decap_8 FILLER_12_2346 ();
 sg13g2_fill_2 FILLER_12_2353 ();
 sg13g2_fill_1 FILLER_12_2355 ();
 sg13g2_decap_8 FILLER_12_2360 ();
 sg13g2_decap_8 FILLER_12_2367 ();
 sg13g2_fill_2 FILLER_12_2374 ();
 sg13g2_fill_1 FILLER_12_2376 ();
 sg13g2_fill_1 FILLER_12_2382 ();
 sg13g2_decap_8 FILLER_12_2413 ();
 sg13g2_fill_1 FILLER_12_2420 ();
 sg13g2_decap_8 FILLER_12_2509 ();
 sg13g2_decap_8 FILLER_12_2516 ();
 sg13g2_decap_8 FILLER_12_2523 ();
 sg13g2_decap_4 FILLER_12_2530 ();
 sg13g2_decap_8 FILLER_12_2570 ();
 sg13g2_decap_8 FILLER_12_2577 ();
 sg13g2_decap_4 FILLER_12_2584 ();
 sg13g2_decap_8 FILLER_12_2624 ();
 sg13g2_decap_8 FILLER_12_2631 ();
 sg13g2_decap_8 FILLER_12_2638 ();
 sg13g2_decap_8 FILLER_12_2645 ();
 sg13g2_fill_1 FILLER_12_2652 ();
 sg13g2_decap_8 FILLER_12_2679 ();
 sg13g2_decap_8 FILLER_12_2686 ();
 sg13g2_decap_4 FILLER_12_2693 ();
 sg13g2_fill_2 FILLER_12_2697 ();
 sg13g2_decap_8 FILLER_12_2709 ();
 sg13g2_decap_4 FILLER_12_2716 ();
 sg13g2_fill_1 FILLER_12_2720 ();
 sg13g2_decap_8 FILLER_12_2747 ();
 sg13g2_decap_8 FILLER_12_2754 ();
 sg13g2_decap_8 FILLER_12_2761 ();
 sg13g2_decap_8 FILLER_12_2768 ();
 sg13g2_decap_8 FILLER_12_2775 ();
 sg13g2_decap_4 FILLER_12_2782 ();
 sg13g2_fill_1 FILLER_12_2789 ();
 sg13g2_decap_8 FILLER_12_2805 ();
 sg13g2_decap_8 FILLER_12_2812 ();
 sg13g2_fill_1 FILLER_12_2819 ();
 sg13g2_decap_8 FILLER_12_2835 ();
 sg13g2_decap_8 FILLER_12_2842 ();
 sg13g2_decap_8 FILLER_12_2849 ();
 sg13g2_decap_8 FILLER_12_2856 ();
 sg13g2_decap_8 FILLER_12_2878 ();
 sg13g2_decap_8 FILLER_12_2885 ();
 sg13g2_decap_4 FILLER_12_2892 ();
 sg13g2_fill_2 FILLER_12_2896 ();
 sg13g2_decap_8 FILLER_12_2903 ();
 sg13g2_fill_1 FILLER_12_2910 ();
 sg13g2_decap_4 FILLER_12_2921 ();
 sg13g2_fill_1 FILLER_12_2925 ();
 sg13g2_decap_8 FILLER_12_2930 ();
 sg13g2_decap_8 FILLER_12_2937 ();
 sg13g2_decap_8 FILLER_12_2944 ();
 sg13g2_decap_8 FILLER_12_2951 ();
 sg13g2_decap_8 FILLER_12_2958 ();
 sg13g2_decap_8 FILLER_12_2965 ();
 sg13g2_decap_8 FILLER_12_2972 ();
 sg13g2_decap_4 FILLER_12_2979 ();
 sg13g2_fill_2 FILLER_12_2983 ();
 sg13g2_decap_8 FILLER_12_3011 ();
 sg13g2_decap_8 FILLER_12_3018 ();
 sg13g2_decap_8 FILLER_12_3025 ();
 sg13g2_decap_8 FILLER_12_3032 ();
 sg13g2_decap_8 FILLER_12_3039 ();
 sg13g2_decap_8 FILLER_12_3046 ();
 sg13g2_decap_8 FILLER_12_3053 ();
 sg13g2_decap_8 FILLER_12_3060 ();
 sg13g2_decap_8 FILLER_12_3067 ();
 sg13g2_decap_8 FILLER_12_3074 ();
 sg13g2_decap_8 FILLER_12_3081 ();
 sg13g2_decap_8 FILLER_12_3088 ();
 sg13g2_decap_4 FILLER_12_3095 ();
 sg13g2_fill_2 FILLER_12_3099 ();
 sg13g2_decap_8 FILLER_12_3104 ();
 sg13g2_decap_8 FILLER_12_3111 ();
 sg13g2_fill_1 FILLER_12_3123 ();
 sg13g2_fill_2 FILLER_12_3134 ();
 sg13g2_fill_1 FILLER_12_3136 ();
 sg13g2_decap_8 FILLER_12_3142 ();
 sg13g2_decap_8 FILLER_12_3154 ();
 sg13g2_decap_8 FILLER_12_3161 ();
 sg13g2_decap_8 FILLER_12_3168 ();
 sg13g2_decap_8 FILLER_12_3175 ();
 sg13g2_decap_8 FILLER_12_3182 ();
 sg13g2_decap_8 FILLER_12_3189 ();
 sg13g2_decap_8 FILLER_12_3196 ();
 sg13g2_decap_8 FILLER_12_3203 ();
 sg13g2_decap_8 FILLER_12_3210 ();
 sg13g2_decap_8 FILLER_12_3217 ();
 sg13g2_decap_8 FILLER_12_3224 ();
 sg13g2_decap_8 FILLER_12_3231 ();
 sg13g2_decap_8 FILLER_12_3258 ();
 sg13g2_fill_2 FILLER_12_3265 ();
 sg13g2_fill_1 FILLER_12_3267 ();
 sg13g2_decap_8 FILLER_12_3298 ();
 sg13g2_fill_2 FILLER_12_3305 ();
 sg13g2_decap_4 FILLER_12_3338 ();
 sg13g2_fill_2 FILLER_12_3342 ();
 sg13g2_decap_8 FILLER_12_3365 ();
 sg13g2_fill_2 FILLER_12_3380 ();
 sg13g2_fill_1 FILLER_12_3382 ();
 sg13g2_decap_8 FILLER_12_3393 ();
 sg13g2_decap_8 FILLER_12_3400 ();
 sg13g2_decap_8 FILLER_12_3407 ();
 sg13g2_decap_4 FILLER_12_3414 ();
 sg13g2_fill_2 FILLER_12_3418 ();
 sg13g2_decap_8 FILLER_12_3440 ();
 sg13g2_decap_8 FILLER_12_3447 ();
 sg13g2_decap_8 FILLER_12_3454 ();
 sg13g2_decap_4 FILLER_12_3461 ();
 sg13g2_decap_8 FILLER_12_3470 ();
 sg13g2_decap_8 FILLER_12_3477 ();
 sg13g2_decap_8 FILLER_12_3484 ();
 sg13g2_decap_8 FILLER_12_3491 ();
 sg13g2_decap_8 FILLER_12_3498 ();
 sg13g2_decap_8 FILLER_12_3505 ();
 sg13g2_decap_8 FILLER_12_3512 ();
 sg13g2_decap_8 FILLER_12_3519 ();
 sg13g2_decap_8 FILLER_12_3526 ();
 sg13g2_decap_8 FILLER_12_3533 ();
 sg13g2_decap_8 FILLER_12_3540 ();
 sg13g2_decap_8 FILLER_12_3547 ();
 sg13g2_decap_8 FILLER_12_3554 ();
 sg13g2_decap_8 FILLER_12_3561 ();
 sg13g2_decap_8 FILLER_12_3568 ();
 sg13g2_decap_4 FILLER_12_3575 ();
 sg13g2_fill_1 FILLER_12_3579 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_4 FILLER_13_7 ();
 sg13g2_fill_2 FILLER_13_11 ();
 sg13g2_decap_8 FILLER_13_46 ();
 sg13g2_decap_8 FILLER_13_53 ();
 sg13g2_decap_4 FILLER_13_60 ();
 sg13g2_fill_2 FILLER_13_110 ();
 sg13g2_fill_1 FILLER_13_112 ();
 sg13g2_fill_2 FILLER_13_123 ();
 sg13g2_decap_4 FILLER_13_141 ();
 sg13g2_fill_2 FILLER_13_145 ();
 sg13g2_decap_8 FILLER_13_165 ();
 sg13g2_decap_8 FILLER_13_172 ();
 sg13g2_decap_8 FILLER_13_179 ();
 sg13g2_decap_8 FILLER_13_186 ();
 sg13g2_decap_8 FILLER_13_193 ();
 sg13g2_decap_4 FILLER_13_200 ();
 sg13g2_fill_1 FILLER_13_204 ();
 sg13g2_decap_8 FILLER_13_236 ();
 sg13g2_decap_8 FILLER_13_243 ();
 sg13g2_decap_8 FILLER_13_250 ();
 sg13g2_decap_4 FILLER_13_257 ();
 sg13g2_fill_1 FILLER_13_261 ();
 sg13g2_decap_8 FILLER_13_296 ();
 sg13g2_decap_8 FILLER_13_303 ();
 sg13g2_decap_8 FILLER_13_310 ();
 sg13g2_decap_8 FILLER_13_317 ();
 sg13g2_decap_8 FILLER_13_324 ();
 sg13g2_decap_4 FILLER_13_331 ();
 sg13g2_fill_2 FILLER_13_335 ();
 sg13g2_decap_8 FILLER_13_351 ();
 sg13g2_decap_8 FILLER_13_358 ();
 sg13g2_decap_8 FILLER_13_365 ();
 sg13g2_decap_8 FILLER_13_372 ();
 sg13g2_decap_8 FILLER_13_379 ();
 sg13g2_decap_8 FILLER_13_386 ();
 sg13g2_decap_4 FILLER_13_393 ();
 sg13g2_fill_1 FILLER_13_397 ();
 sg13g2_fill_2 FILLER_13_416 ();
 sg13g2_decap_8 FILLER_13_463 ();
 sg13g2_decap_8 FILLER_13_470 ();
 sg13g2_decap_8 FILLER_13_477 ();
 sg13g2_decap_8 FILLER_13_484 ();
 sg13g2_decap_8 FILLER_13_491 ();
 sg13g2_decap_4 FILLER_13_498 ();
 sg13g2_fill_2 FILLER_13_502 ();
 sg13g2_decap_8 FILLER_13_530 ();
 sg13g2_decap_8 FILLER_13_589 ();
 sg13g2_decap_8 FILLER_13_596 ();
 sg13g2_decap_8 FILLER_13_603 ();
 sg13g2_decap_8 FILLER_13_610 ();
 sg13g2_decap_8 FILLER_13_617 ();
 sg13g2_decap_8 FILLER_13_624 ();
 sg13g2_decap_4 FILLER_13_631 ();
 sg13g2_decap_8 FILLER_13_661 ();
 sg13g2_decap_8 FILLER_13_668 ();
 sg13g2_decap_8 FILLER_13_675 ();
 sg13g2_decap_8 FILLER_13_682 ();
 sg13g2_decap_8 FILLER_13_689 ();
 sg13g2_decap_8 FILLER_13_696 ();
 sg13g2_decap_8 FILLER_13_703 ();
 sg13g2_decap_8 FILLER_13_710 ();
 sg13g2_decap_8 FILLER_13_717 ();
 sg13g2_decap_8 FILLER_13_724 ();
 sg13g2_decap_8 FILLER_13_731 ();
 sg13g2_fill_2 FILLER_13_738 ();
 sg13g2_decap_4 FILLER_13_766 ();
 sg13g2_fill_2 FILLER_13_770 ();
 sg13g2_fill_1 FILLER_13_808 ();
 sg13g2_decap_8 FILLER_13_822 ();
 sg13g2_decap_8 FILLER_13_829 ();
 sg13g2_decap_4 FILLER_13_836 ();
 sg13g2_decap_8 FILLER_13_845 ();
 sg13g2_decap_8 FILLER_13_852 ();
 sg13g2_decap_8 FILLER_13_859 ();
 sg13g2_fill_1 FILLER_13_866 ();
 sg13g2_decap_8 FILLER_13_887 ();
 sg13g2_decap_8 FILLER_13_894 ();
 sg13g2_decap_8 FILLER_13_901 ();
 sg13g2_fill_1 FILLER_13_908 ();
 sg13g2_decap_8 FILLER_13_919 ();
 sg13g2_decap_8 FILLER_13_926 ();
 sg13g2_decap_8 FILLER_13_933 ();
 sg13g2_decap_8 FILLER_13_940 ();
 sg13g2_decap_8 FILLER_13_947 ();
 sg13g2_decap_8 FILLER_13_954 ();
 sg13g2_decap_4 FILLER_13_961 ();
 sg13g2_decap_8 FILLER_13_973 ();
 sg13g2_decap_8 FILLER_13_980 ();
 sg13g2_decap_8 FILLER_13_987 ();
 sg13g2_decap_8 FILLER_13_994 ();
 sg13g2_decap_8 FILLER_13_1001 ();
 sg13g2_decap_8 FILLER_13_1008 ();
 sg13g2_fill_2 FILLER_13_1015 ();
 sg13g2_decap_4 FILLER_13_1022 ();
 sg13g2_fill_2 FILLER_13_1034 ();
 sg13g2_fill_1 FILLER_13_1036 ();
 sg13g2_decap_8 FILLER_13_1048 ();
 sg13g2_decap_8 FILLER_13_1055 ();
 sg13g2_decap_8 FILLER_13_1062 ();
 sg13g2_fill_2 FILLER_13_1069 ();
 sg13g2_fill_1 FILLER_13_1071 ();
 sg13g2_fill_1 FILLER_13_1081 ();
 sg13g2_decap_8 FILLER_13_1085 ();
 sg13g2_decap_8 FILLER_13_1092 ();
 sg13g2_fill_2 FILLER_13_1099 ();
 sg13g2_fill_1 FILLER_13_1101 ();
 sg13g2_decap_8 FILLER_13_1110 ();
 sg13g2_fill_1 FILLER_13_1117 ();
 sg13g2_decap_8 FILLER_13_1133 ();
 sg13g2_decap_4 FILLER_13_1140 ();
 sg13g2_fill_2 FILLER_13_1144 ();
 sg13g2_decap_8 FILLER_13_1151 ();
 sg13g2_decap_8 FILLER_13_1158 ();
 sg13g2_decap_8 FILLER_13_1165 ();
 sg13g2_decap_8 FILLER_13_1172 ();
 sg13g2_decap_8 FILLER_13_1179 ();
 sg13g2_fill_1 FILLER_13_1186 ();
 sg13g2_decap_8 FILLER_13_1208 ();
 sg13g2_decap_8 FILLER_13_1215 ();
 sg13g2_decap_8 FILLER_13_1222 ();
 sg13g2_decap_8 FILLER_13_1229 ();
 sg13g2_decap_8 FILLER_13_1236 ();
 sg13g2_decap_4 FILLER_13_1243 ();
 sg13g2_decap_8 FILLER_13_1291 ();
 sg13g2_decap_8 FILLER_13_1356 ();
 sg13g2_decap_8 FILLER_13_1363 ();
 sg13g2_decap_8 FILLER_13_1370 ();
 sg13g2_decap_4 FILLER_13_1377 ();
 sg13g2_fill_1 FILLER_13_1381 ();
 sg13g2_decap_8 FILLER_13_1411 ();
 sg13g2_fill_2 FILLER_13_1418 ();
 sg13g2_fill_1 FILLER_13_1420 ();
 sg13g2_decap_8 FILLER_13_1425 ();
 sg13g2_decap_8 FILLER_13_1432 ();
 sg13g2_decap_8 FILLER_13_1439 ();
 sg13g2_fill_1 FILLER_13_1446 ();
 sg13g2_decap_8 FILLER_13_1473 ();
 sg13g2_fill_2 FILLER_13_1480 ();
 sg13g2_fill_1 FILLER_13_1482 ();
 sg13g2_decap_8 FILLER_13_1519 ();
 sg13g2_decap_8 FILLER_13_1526 ();
 sg13g2_decap_8 FILLER_13_1533 ();
 sg13g2_decap_8 FILLER_13_1540 ();
 sg13g2_decap_4 FILLER_13_1547 ();
 sg13g2_fill_2 FILLER_13_1551 ();
 sg13g2_fill_2 FILLER_13_1563 ();
 sg13g2_fill_2 FILLER_13_1575 ();
 sg13g2_decap_8 FILLER_13_1593 ();
 sg13g2_decap_8 FILLER_13_1600 ();
 sg13g2_decap_8 FILLER_13_1607 ();
 sg13g2_decap_8 FILLER_13_1614 ();
 sg13g2_fill_1 FILLER_13_1621 ();
 sg13g2_decap_8 FILLER_13_1648 ();
 sg13g2_fill_2 FILLER_13_1655 ();
 sg13g2_fill_1 FILLER_13_1657 ();
 sg13g2_decap_8 FILLER_13_1684 ();
 sg13g2_decap_8 FILLER_13_1691 ();
 sg13g2_decap_8 FILLER_13_1698 ();
 sg13g2_decap_8 FILLER_13_1705 ();
 sg13g2_fill_1 FILLER_13_1712 ();
 sg13g2_decap_8 FILLER_13_1716 ();
 sg13g2_decap_8 FILLER_13_1727 ();
 sg13g2_decap_8 FILLER_13_1734 ();
 sg13g2_decap_8 FILLER_13_1741 ();
 sg13g2_decap_8 FILLER_13_1748 ();
 sg13g2_decap_8 FILLER_13_1755 ();
 sg13g2_decap_8 FILLER_13_1762 ();
 sg13g2_decap_8 FILLER_13_1769 ();
 sg13g2_decap_4 FILLER_13_1776 ();
 sg13g2_fill_2 FILLER_13_1780 ();
 sg13g2_decap_8 FILLER_13_1785 ();
 sg13g2_decap_8 FILLER_13_1792 ();
 sg13g2_decap_8 FILLER_13_1799 ();
 sg13g2_decap_8 FILLER_13_1806 ();
 sg13g2_decap_8 FILLER_13_1813 ();
 sg13g2_decap_8 FILLER_13_1820 ();
 sg13g2_decap_8 FILLER_13_1827 ();
 sg13g2_decap_8 FILLER_13_1834 ();
 sg13g2_decap_8 FILLER_13_1841 ();
 sg13g2_decap_8 FILLER_13_1848 ();
 sg13g2_decap_8 FILLER_13_1855 ();
 sg13g2_decap_4 FILLER_13_1862 ();
 sg13g2_decap_8 FILLER_13_1905 ();
 sg13g2_decap_8 FILLER_13_1912 ();
 sg13g2_decap_8 FILLER_13_1919 ();
 sg13g2_fill_1 FILLER_13_1948 ();
 sg13g2_decap_8 FILLER_13_1956 ();
 sg13g2_decap_8 FILLER_13_1963 ();
 sg13g2_decap_8 FILLER_13_1970 ();
 sg13g2_decap_8 FILLER_13_1977 ();
 sg13g2_decap_8 FILLER_13_1984 ();
 sg13g2_decap_8 FILLER_13_1991 ();
 sg13g2_decap_4 FILLER_13_1998 ();
 sg13g2_fill_1 FILLER_13_2002 ();
 sg13g2_decap_8 FILLER_13_2008 ();
 sg13g2_decap_8 FILLER_13_2015 ();
 sg13g2_decap_8 FILLER_13_2038 ();
 sg13g2_decap_8 FILLER_13_2071 ();
 sg13g2_decap_8 FILLER_13_2078 ();
 sg13g2_fill_2 FILLER_13_2085 ();
 sg13g2_fill_1 FILLER_13_2087 ();
 sg13g2_fill_1 FILLER_13_2098 ();
 sg13g2_decap_8 FILLER_13_2125 ();
 sg13g2_decap_8 FILLER_13_2132 ();
 sg13g2_decap_8 FILLER_13_2139 ();
 sg13g2_decap_8 FILLER_13_2156 ();
 sg13g2_decap_8 FILLER_13_2163 ();
 sg13g2_decap_4 FILLER_13_2170 ();
 sg13g2_decap_8 FILLER_13_2177 ();
 sg13g2_decap_8 FILLER_13_2184 ();
 sg13g2_decap_8 FILLER_13_2191 ();
 sg13g2_decap_8 FILLER_13_2198 ();
 sg13g2_decap_8 FILLER_13_2205 ();
 sg13g2_decap_8 FILLER_13_2212 ();
 sg13g2_decap_8 FILLER_13_2219 ();
 sg13g2_decap_8 FILLER_13_2226 ();
 sg13g2_decap_8 FILLER_13_2233 ();
 sg13g2_decap_8 FILLER_13_2240 ();
 sg13g2_decap_8 FILLER_13_2247 ();
 sg13g2_decap_8 FILLER_13_2254 ();
 sg13g2_decap_8 FILLER_13_2261 ();
 sg13g2_decap_8 FILLER_13_2268 ();
 sg13g2_decap_8 FILLER_13_2275 ();
 sg13g2_decap_8 FILLER_13_2282 ();
 sg13g2_fill_2 FILLER_13_2289 ();
 sg13g2_fill_1 FILLER_13_2291 ();
 sg13g2_decap_8 FILLER_13_2295 ();
 sg13g2_decap_8 FILLER_13_2302 ();
 sg13g2_decap_8 FILLER_13_2309 ();
 sg13g2_decap_8 FILLER_13_2316 ();
 sg13g2_decap_8 FILLER_13_2323 ();
 sg13g2_decap_8 FILLER_13_2330 ();
 sg13g2_fill_2 FILLER_13_2337 ();
 sg13g2_decap_8 FILLER_13_2355 ();
 sg13g2_decap_8 FILLER_13_2362 ();
 sg13g2_decap_8 FILLER_13_2369 ();
 sg13g2_decap_8 FILLER_13_2376 ();
 sg13g2_decap_8 FILLER_13_2383 ();
 sg13g2_fill_2 FILLER_13_2390 ();
 sg13g2_fill_1 FILLER_13_2392 ();
 sg13g2_decap_8 FILLER_13_2397 ();
 sg13g2_decap_8 FILLER_13_2404 ();
 sg13g2_decap_8 FILLER_13_2411 ();
 sg13g2_decap_4 FILLER_13_2418 ();
 sg13g2_fill_2 FILLER_13_2422 ();
 sg13g2_decap_8 FILLER_13_2434 ();
 sg13g2_decap_8 FILLER_13_2441 ();
 sg13g2_decap_8 FILLER_13_2448 ();
 sg13g2_decap_8 FILLER_13_2455 ();
 sg13g2_fill_1 FILLER_13_2462 ();
 sg13g2_decap_8 FILLER_13_2467 ();
 sg13g2_decap_8 FILLER_13_2474 ();
 sg13g2_decap_8 FILLER_13_2481 ();
 sg13g2_decap_8 FILLER_13_2488 ();
 sg13g2_decap_8 FILLER_13_2495 ();
 sg13g2_decap_8 FILLER_13_2512 ();
 sg13g2_decap_8 FILLER_13_2519 ();
 sg13g2_decap_8 FILLER_13_2526 ();
 sg13g2_decap_8 FILLER_13_2533 ();
 sg13g2_decap_8 FILLER_13_2540 ();
 sg13g2_fill_2 FILLER_13_2547 ();
 sg13g2_fill_1 FILLER_13_2549 ();
 sg13g2_decap_8 FILLER_13_2579 ();
 sg13g2_decap_8 FILLER_13_2586 ();
 sg13g2_decap_8 FILLER_13_2593 ();
 sg13g2_decap_8 FILLER_13_2600 ();
 sg13g2_fill_1 FILLER_13_2607 ();
 sg13g2_fill_2 FILLER_13_2638 ();
 sg13g2_fill_1 FILLER_13_2650 ();
 sg13g2_decap_8 FILLER_13_2661 ();
 sg13g2_decap_8 FILLER_13_2668 ();
 sg13g2_decap_8 FILLER_13_2675 ();
 sg13g2_decap_8 FILLER_13_2682 ();
 sg13g2_decap_8 FILLER_13_2699 ();
 sg13g2_fill_1 FILLER_13_2706 ();
 sg13g2_decap_4 FILLER_13_2733 ();
 sg13g2_decap_8 FILLER_13_2747 ();
 sg13g2_decap_8 FILLER_13_2754 ();
 sg13g2_decap_8 FILLER_13_2761 ();
 sg13g2_decap_4 FILLER_13_2768 ();
 sg13g2_fill_1 FILLER_13_2772 ();
 sg13g2_decap_8 FILLER_13_2778 ();
 sg13g2_decap_8 FILLER_13_2785 ();
 sg13g2_decap_8 FILLER_13_2792 ();
 sg13g2_decap_8 FILLER_13_2799 ();
 sg13g2_decap_4 FILLER_13_2806 ();
 sg13g2_fill_1 FILLER_13_2810 ();
 sg13g2_decap_8 FILLER_13_2816 ();
 sg13g2_decap_8 FILLER_13_2823 ();
 sg13g2_fill_2 FILLER_13_2830 ();
 sg13g2_fill_1 FILLER_13_2832 ();
 sg13g2_fill_2 FILLER_13_2838 ();
 sg13g2_fill_1 FILLER_13_2840 ();
 sg13g2_decap_8 FILLER_13_2845 ();
 sg13g2_decap_8 FILLER_13_2852 ();
 sg13g2_decap_8 FILLER_13_2859 ();
 sg13g2_decap_8 FILLER_13_2866 ();
 sg13g2_fill_2 FILLER_13_2873 ();
 sg13g2_fill_1 FILLER_13_2875 ();
 sg13g2_decap_8 FILLER_13_2881 ();
 sg13g2_decap_8 FILLER_13_2888 ();
 sg13g2_decap_8 FILLER_13_2895 ();
 sg13g2_decap_8 FILLER_13_2902 ();
 sg13g2_decap_8 FILLER_13_2909 ();
 sg13g2_fill_2 FILLER_13_2916 ();
 sg13g2_decap_8 FILLER_13_2953 ();
 sg13g2_decap_8 FILLER_13_2960 ();
 sg13g2_decap_8 FILLER_13_2967 ();
 sg13g2_decap_4 FILLER_13_2974 ();
 sg13g2_fill_2 FILLER_13_2978 ();
 sg13g2_decap_8 FILLER_13_3016 ();
 sg13g2_decap_8 FILLER_13_3023 ();
 sg13g2_fill_2 FILLER_13_3030 ();
 sg13g2_decap_8 FILLER_13_3058 ();
 sg13g2_decap_8 FILLER_13_3065 ();
 sg13g2_decap_8 FILLER_13_3072 ();
 sg13g2_decap_4 FILLER_13_3079 ();
 sg13g2_decap_8 FILLER_13_3087 ();
 sg13g2_decap_8 FILLER_13_3094 ();
 sg13g2_fill_1 FILLER_13_3101 ();
 sg13g2_decap_8 FILLER_13_3105 ();
 sg13g2_decap_8 FILLER_13_3112 ();
 sg13g2_decap_8 FILLER_13_3119 ();
 sg13g2_decap_4 FILLER_13_3126 ();
 sg13g2_fill_2 FILLER_13_3130 ();
 sg13g2_decap_4 FILLER_13_3137 ();
 sg13g2_fill_2 FILLER_13_3141 ();
 sg13g2_decap_8 FILLER_13_3152 ();
 sg13g2_decap_8 FILLER_13_3159 ();
 sg13g2_decap_8 FILLER_13_3166 ();
 sg13g2_decap_8 FILLER_13_3173 ();
 sg13g2_decap_8 FILLER_13_3180 ();
 sg13g2_decap_8 FILLER_13_3187 ();
 sg13g2_decap_8 FILLER_13_3194 ();
 sg13g2_decap_4 FILLER_13_3201 ();
 sg13g2_decap_8 FILLER_13_3218 ();
 sg13g2_decap_8 FILLER_13_3225 ();
 sg13g2_fill_2 FILLER_13_3232 ();
 sg13g2_decap_4 FILLER_13_3242 ();
 sg13g2_decap_8 FILLER_13_3251 ();
 sg13g2_decap_8 FILLER_13_3258 ();
 sg13g2_decap_8 FILLER_13_3270 ();
 sg13g2_decap_8 FILLER_13_3277 ();
 sg13g2_decap_8 FILLER_13_3284 ();
 sg13g2_decap_8 FILLER_13_3291 ();
 sg13g2_decap_8 FILLER_13_3298 ();
 sg13g2_decap_8 FILLER_13_3305 ();
 sg13g2_decap_8 FILLER_13_3312 ();
 sg13g2_decap_8 FILLER_13_3319 ();
 sg13g2_decap_8 FILLER_13_3326 ();
 sg13g2_decap_8 FILLER_13_3333 ();
 sg13g2_decap_4 FILLER_13_3340 ();
 sg13g2_decap_8 FILLER_13_3365 ();
 sg13g2_decap_4 FILLER_13_3372 ();
 sg13g2_fill_1 FILLER_13_3376 ();
 sg13g2_decap_8 FILLER_13_3387 ();
 sg13g2_decap_8 FILLER_13_3394 ();
 sg13g2_decap_8 FILLER_13_3406 ();
 sg13g2_decap_4 FILLER_13_3413 ();
 sg13g2_fill_2 FILLER_13_3417 ();
 sg13g2_fill_2 FILLER_13_3424 ();
 sg13g2_fill_2 FILLER_13_3431 ();
 sg13g2_fill_2 FILLER_13_3451 ();
 sg13g2_decap_8 FILLER_13_3479 ();
 sg13g2_decap_8 FILLER_13_3486 ();
 sg13g2_decap_8 FILLER_13_3493 ();
 sg13g2_decap_8 FILLER_13_3500 ();
 sg13g2_decap_8 FILLER_13_3507 ();
 sg13g2_decap_8 FILLER_13_3514 ();
 sg13g2_decap_8 FILLER_13_3521 ();
 sg13g2_decap_8 FILLER_13_3528 ();
 sg13g2_decap_8 FILLER_13_3535 ();
 sg13g2_decap_8 FILLER_13_3542 ();
 sg13g2_decap_8 FILLER_13_3549 ();
 sg13g2_decap_8 FILLER_13_3556 ();
 sg13g2_decap_8 FILLER_13_3563 ();
 sg13g2_decap_8 FILLER_13_3570 ();
 sg13g2_fill_2 FILLER_13_3577 ();
 sg13g2_fill_1 FILLER_13_3579 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_fill_2 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_40 ();
 sg13g2_decap_8 FILLER_14_47 ();
 sg13g2_decap_8 FILLER_14_54 ();
 sg13g2_fill_2 FILLER_14_61 ();
 sg13g2_fill_2 FILLER_14_85 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_4 FILLER_14_112 ();
 sg13g2_fill_2 FILLER_14_116 ();
 sg13g2_fill_1 FILLER_14_122 ();
 sg13g2_fill_1 FILLER_14_128 ();
 sg13g2_decap_8 FILLER_14_134 ();
 sg13g2_decap_4 FILLER_14_141 ();
 sg13g2_fill_1 FILLER_14_145 ();
 sg13g2_decap_8 FILLER_14_163 ();
 sg13g2_decap_8 FILLER_14_170 ();
 sg13g2_decap_8 FILLER_14_177 ();
 sg13g2_decap_8 FILLER_14_184 ();
 sg13g2_decap_8 FILLER_14_191 ();
 sg13g2_decap_8 FILLER_14_198 ();
 sg13g2_decap_8 FILLER_14_205 ();
 sg13g2_fill_2 FILLER_14_212 ();
 sg13g2_fill_1 FILLER_14_214 ();
 sg13g2_decap_8 FILLER_14_228 ();
 sg13g2_decap_8 FILLER_14_235 ();
 sg13g2_decap_8 FILLER_14_242 ();
 sg13g2_decap_8 FILLER_14_249 ();
 sg13g2_decap_4 FILLER_14_256 ();
 sg13g2_fill_2 FILLER_14_260 ();
 sg13g2_decap_4 FILLER_14_282 ();
 sg13g2_decap_8 FILLER_14_297 ();
 sg13g2_decap_8 FILLER_14_304 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_fill_2 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_353 ();
 sg13g2_fill_1 FILLER_14_360 ();
 sg13g2_fill_2 FILLER_14_369 ();
 sg13g2_decap_8 FILLER_14_379 ();
 sg13g2_decap_8 FILLER_14_386 ();
 sg13g2_decap_8 FILLER_14_393 ();
 sg13g2_decap_8 FILLER_14_400 ();
 sg13g2_fill_2 FILLER_14_415 ();
 sg13g2_fill_1 FILLER_14_417 ();
 sg13g2_fill_2 FILLER_14_426 ();
 sg13g2_decap_4 FILLER_14_433 ();
 sg13g2_fill_1 FILLER_14_437 ();
 sg13g2_fill_2 FILLER_14_446 ();
 sg13g2_decap_8 FILLER_14_456 ();
 sg13g2_decap_8 FILLER_14_463 ();
 sg13g2_decap_8 FILLER_14_470 ();
 sg13g2_decap_8 FILLER_14_477 ();
 sg13g2_fill_2 FILLER_14_484 ();
 sg13g2_decap_8 FILLER_14_496 ();
 sg13g2_decap_8 FILLER_14_503 ();
 sg13g2_fill_2 FILLER_14_510 ();
 sg13g2_decap_8 FILLER_14_522 ();
 sg13g2_decap_8 FILLER_14_529 ();
 sg13g2_fill_1 FILLER_14_536 ();
 sg13g2_decap_8 FILLER_14_547 ();
 sg13g2_decap_4 FILLER_14_554 ();
 sg13g2_fill_1 FILLER_14_558 ();
 sg13g2_decap_8 FILLER_14_569 ();
 sg13g2_fill_2 FILLER_14_576 ();
 sg13g2_fill_1 FILLER_14_578 ();
 sg13g2_decap_8 FILLER_14_605 ();
 sg13g2_decap_8 FILLER_14_612 ();
 sg13g2_decap_8 FILLER_14_619 ();
 sg13g2_decap_8 FILLER_14_626 ();
 sg13g2_decap_8 FILLER_14_633 ();
 sg13g2_decap_4 FILLER_14_640 ();
 sg13g2_decap_8 FILLER_14_670 ();
 sg13g2_decap_8 FILLER_14_697 ();
 sg13g2_fill_1 FILLER_14_704 ();
 sg13g2_decap_4 FILLER_14_715 ();
 sg13g2_fill_2 FILLER_14_719 ();
 sg13g2_decap_8 FILLER_14_726 ();
 sg13g2_decap_8 FILLER_14_733 ();
 sg13g2_decap_8 FILLER_14_740 ();
 sg13g2_decap_8 FILLER_14_747 ();
 sg13g2_decap_4 FILLER_14_754 ();
 sg13g2_decap_8 FILLER_14_768 ();
 sg13g2_decap_4 FILLER_14_775 ();
 sg13g2_fill_1 FILLER_14_779 ();
 sg13g2_decap_8 FILLER_14_789 ();
 sg13g2_decap_8 FILLER_14_796 ();
 sg13g2_decap_8 FILLER_14_803 ();
 sg13g2_decap_8 FILLER_14_810 ();
 sg13g2_decap_8 FILLER_14_817 ();
 sg13g2_fill_2 FILLER_14_824 ();
 sg13g2_decap_8 FILLER_14_855 ();
 sg13g2_decap_8 FILLER_14_862 ();
 sg13g2_decap_8 FILLER_14_905 ();
 sg13g2_decap_8 FILLER_14_912 ();
 sg13g2_decap_4 FILLER_14_919 ();
 sg13g2_decap_8 FILLER_14_933 ();
 sg13g2_fill_2 FILLER_14_940 ();
 sg13g2_decap_8 FILLER_14_978 ();
 sg13g2_decap_8 FILLER_14_985 ();
 sg13g2_decap_8 FILLER_14_992 ();
 sg13g2_decap_8 FILLER_14_999 ();
 sg13g2_fill_2 FILLER_14_1006 ();
 sg13g2_decap_4 FILLER_14_1034 ();
 sg13g2_fill_2 FILLER_14_1038 ();
 sg13g2_decap_8 FILLER_14_1043 ();
 sg13g2_decap_8 FILLER_14_1050 ();
 sg13g2_decap_4 FILLER_14_1057 ();
 sg13g2_decap_8 FILLER_14_1092 ();
 sg13g2_decap_4 FILLER_14_1099 ();
 sg13g2_fill_2 FILLER_14_1103 ();
 sg13g2_decap_4 FILLER_14_1110 ();
 sg13g2_fill_1 FILLER_14_1114 ();
 sg13g2_fill_2 FILLER_14_1126 ();
 sg13g2_fill_1 FILLER_14_1128 ();
 sg13g2_decap_8 FILLER_14_1143 ();
 sg13g2_decap_8 FILLER_14_1150 ();
 sg13g2_decap_8 FILLER_14_1157 ();
 sg13g2_decap_8 FILLER_14_1164 ();
 sg13g2_decap_8 FILLER_14_1171 ();
 sg13g2_fill_1 FILLER_14_1178 ();
 sg13g2_decap_8 FILLER_14_1215 ();
 sg13g2_decap_8 FILLER_14_1222 ();
 sg13g2_decap_8 FILLER_14_1229 ();
 sg13g2_decap_8 FILLER_14_1236 ();
 sg13g2_decap_8 FILLER_14_1243 ();
 sg13g2_decap_4 FILLER_14_1250 ();
 sg13g2_fill_2 FILLER_14_1254 ();
 sg13g2_fill_1 FILLER_14_1268 ();
 sg13g2_decap_8 FILLER_14_1274 ();
 sg13g2_decap_8 FILLER_14_1281 ();
 sg13g2_decap_8 FILLER_14_1288 ();
 sg13g2_decap_8 FILLER_14_1295 ();
 sg13g2_decap_4 FILLER_14_1302 ();
 sg13g2_decap_4 FILLER_14_1325 ();
 sg13g2_decap_4 FILLER_14_1338 ();
 sg13g2_fill_1 FILLER_14_1342 ();
 sg13g2_decap_8 FILLER_14_1352 ();
 sg13g2_decap_8 FILLER_14_1359 ();
 sg13g2_decap_8 FILLER_14_1366 ();
 sg13g2_decap_8 FILLER_14_1373 ();
 sg13g2_decap_4 FILLER_14_1380 ();
 sg13g2_fill_1 FILLER_14_1384 ();
 sg13g2_decap_8 FILLER_14_1388 ();
 sg13g2_decap_8 FILLER_14_1395 ();
 sg13g2_decap_8 FILLER_14_1402 ();
 sg13g2_decap_8 FILLER_14_1409 ();
 sg13g2_fill_1 FILLER_14_1416 ();
 sg13g2_decap_8 FILLER_14_1423 ();
 sg13g2_decap_8 FILLER_14_1430 ();
 sg13g2_decap_8 FILLER_14_1437 ();
 sg13g2_decap_8 FILLER_14_1444 ();
 sg13g2_decap_8 FILLER_14_1451 ();
 sg13g2_decap_8 FILLER_14_1458 ();
 sg13g2_decap_8 FILLER_14_1465 ();
 sg13g2_decap_8 FILLER_14_1472 ();
 sg13g2_decap_4 FILLER_14_1479 ();
 sg13g2_fill_2 FILLER_14_1501 ();
 sg13g2_fill_1 FILLER_14_1503 ();
 sg13g2_decap_8 FILLER_14_1514 ();
 sg13g2_decap_8 FILLER_14_1521 ();
 sg13g2_decap_8 FILLER_14_1528 ();
 sg13g2_decap_8 FILLER_14_1535 ();
 sg13g2_decap_8 FILLER_14_1542 ();
 sg13g2_decap_8 FILLER_14_1585 ();
 sg13g2_decap_8 FILLER_14_1592 ();
 sg13g2_decap_8 FILLER_14_1599 ();
 sg13g2_decap_8 FILLER_14_1606 ();
 sg13g2_decap_8 FILLER_14_1613 ();
 sg13g2_decap_4 FILLER_14_1620 ();
 sg13g2_fill_2 FILLER_14_1624 ();
 sg13g2_decap_8 FILLER_14_1652 ();
 sg13g2_fill_2 FILLER_14_1659 ();
 sg13g2_fill_1 FILLER_14_1661 ();
 sg13g2_decap_8 FILLER_14_1688 ();
 sg13g2_decap_8 FILLER_14_1695 ();
 sg13g2_decap_4 FILLER_14_1702 ();
 sg13g2_fill_1 FILLER_14_1706 ();
 sg13g2_decap_8 FILLER_14_1712 ();
 sg13g2_fill_2 FILLER_14_1719 ();
 sg13g2_fill_1 FILLER_14_1721 ();
 sg13g2_decap_8 FILLER_14_1748 ();
 sg13g2_fill_1 FILLER_14_1755 ();
 sg13g2_decap_8 FILLER_14_1766 ();
 sg13g2_decap_4 FILLER_14_1773 ();
 sg13g2_fill_2 FILLER_14_1777 ();
 sg13g2_decap_8 FILLER_14_1798 ();
 sg13g2_decap_8 FILLER_14_1805 ();
 sg13g2_decap_8 FILLER_14_1812 ();
 sg13g2_decap_8 FILLER_14_1819 ();
 sg13g2_decap_8 FILLER_14_1826 ();
 sg13g2_decap_8 FILLER_14_1833 ();
 sg13g2_decap_8 FILLER_14_1840 ();
 sg13g2_decap_8 FILLER_14_1847 ();
 sg13g2_decap_8 FILLER_14_1854 ();
 sg13g2_decap_8 FILLER_14_1861 ();
 sg13g2_fill_2 FILLER_14_1868 ();
 sg13g2_decap_8 FILLER_14_1886 ();
 sg13g2_decap_8 FILLER_14_1893 ();
 sg13g2_decap_8 FILLER_14_1900 ();
 sg13g2_decap_8 FILLER_14_1907 ();
 sg13g2_decap_8 FILLER_14_1914 ();
 sg13g2_decap_4 FILLER_14_1921 ();
 sg13g2_fill_2 FILLER_14_1925 ();
 sg13g2_decap_8 FILLER_14_1968 ();
 sg13g2_decap_8 FILLER_14_1975 ();
 sg13g2_decap_8 FILLER_14_1982 ();
 sg13g2_decap_8 FILLER_14_1989 ();
 sg13g2_decap_8 FILLER_14_1996 ();
 sg13g2_decap_8 FILLER_14_2003 ();
 sg13g2_decap_8 FILLER_14_2010 ();
 sg13g2_decap_8 FILLER_14_2017 ();
 sg13g2_decap_8 FILLER_14_2024 ();
 sg13g2_decap_8 FILLER_14_2031 ();
 sg13g2_fill_2 FILLER_14_2038 ();
 sg13g2_fill_1 FILLER_14_2040 ();
 sg13g2_fill_2 FILLER_14_2045 ();
 sg13g2_fill_1 FILLER_14_2047 ();
 sg13g2_decap_8 FILLER_14_2056 ();
 sg13g2_decap_8 FILLER_14_2063 ();
 sg13g2_decap_8 FILLER_14_2070 ();
 sg13g2_decap_8 FILLER_14_2077 ();
 sg13g2_decap_8 FILLER_14_2084 ();
 sg13g2_fill_2 FILLER_14_2091 ();
 sg13g2_decap_8 FILLER_14_2106 ();
 sg13g2_decap_8 FILLER_14_2113 ();
 sg13g2_fill_2 FILLER_14_2120 ();
 sg13g2_decap_8 FILLER_14_2127 ();
 sg13g2_decap_8 FILLER_14_2134 ();
 sg13g2_fill_2 FILLER_14_2141 ();
 sg13g2_decap_8 FILLER_14_2169 ();
 sg13g2_decap_8 FILLER_14_2176 ();
 sg13g2_fill_1 FILLER_14_2183 ();
 sg13g2_decap_8 FILLER_14_2213 ();
 sg13g2_decap_8 FILLER_14_2220 ();
 sg13g2_decap_8 FILLER_14_2227 ();
 sg13g2_decap_8 FILLER_14_2234 ();
 sg13g2_decap_8 FILLER_14_2241 ();
 sg13g2_fill_1 FILLER_14_2248 ();
 sg13g2_fill_1 FILLER_14_2267 ();
 sg13g2_decap_8 FILLER_14_2304 ();
 sg13g2_decap_8 FILLER_14_2311 ();
 sg13g2_decap_8 FILLER_14_2318 ();
 sg13g2_decap_8 FILLER_14_2325 ();
 sg13g2_decap_8 FILLER_14_2332 ();
 sg13g2_decap_8 FILLER_14_2339 ();
 sg13g2_decap_8 FILLER_14_2346 ();
 sg13g2_decap_8 FILLER_14_2353 ();
 sg13g2_decap_8 FILLER_14_2360 ();
 sg13g2_decap_8 FILLER_14_2367 ();
 sg13g2_decap_8 FILLER_14_2374 ();
 sg13g2_fill_2 FILLER_14_2381 ();
 sg13g2_decap_8 FILLER_14_2393 ();
 sg13g2_decap_8 FILLER_14_2400 ();
 sg13g2_decap_8 FILLER_14_2407 ();
 sg13g2_decap_8 FILLER_14_2414 ();
 sg13g2_decap_8 FILLER_14_2421 ();
 sg13g2_decap_8 FILLER_14_2428 ();
 sg13g2_decap_8 FILLER_14_2441 ();
 sg13g2_decap_8 FILLER_14_2448 ();
 sg13g2_decap_8 FILLER_14_2455 ();
 sg13g2_decap_8 FILLER_14_2462 ();
 sg13g2_decap_8 FILLER_14_2469 ();
 sg13g2_decap_8 FILLER_14_2476 ();
 sg13g2_decap_8 FILLER_14_2483 ();
 sg13g2_decap_8 FILLER_14_2490 ();
 sg13g2_decap_4 FILLER_14_2497 ();
 sg13g2_decap_8 FILLER_14_2527 ();
 sg13g2_decap_8 FILLER_14_2534 ();
 sg13g2_decap_8 FILLER_14_2541 ();
 sg13g2_decap_8 FILLER_14_2548 ();
 sg13g2_decap_8 FILLER_14_2555 ();
 sg13g2_decap_8 FILLER_14_2562 ();
 sg13g2_decap_8 FILLER_14_2569 ();
 sg13g2_decap_8 FILLER_14_2576 ();
 sg13g2_decap_8 FILLER_14_2583 ();
 sg13g2_decap_8 FILLER_14_2590 ();
 sg13g2_decap_8 FILLER_14_2597 ();
 sg13g2_decap_8 FILLER_14_2604 ();
 sg13g2_decap_8 FILLER_14_2611 ();
 sg13g2_decap_8 FILLER_14_2618 ();
 sg13g2_decap_8 FILLER_14_2625 ();
 sg13g2_decap_8 FILLER_14_2632 ();
 sg13g2_decap_8 FILLER_14_2639 ();
 sg13g2_decap_8 FILLER_14_2646 ();
 sg13g2_decap_8 FILLER_14_2653 ();
 sg13g2_decap_8 FILLER_14_2660 ();
 sg13g2_decap_8 FILLER_14_2667 ();
 sg13g2_decap_8 FILLER_14_2674 ();
 sg13g2_decap_4 FILLER_14_2681 ();
 sg13g2_fill_1 FILLER_14_2695 ();
 sg13g2_decap_8 FILLER_14_2722 ();
 sg13g2_decap_8 FILLER_14_2729 ();
 sg13g2_decap_8 FILLER_14_2736 ();
 sg13g2_decap_8 FILLER_14_2743 ();
 sg13g2_decap_8 FILLER_14_2750 ();
 sg13g2_decap_8 FILLER_14_2793 ();
 sg13g2_decap_8 FILLER_14_2800 ();
 sg13g2_decap_8 FILLER_14_2807 ();
 sg13g2_decap_8 FILLER_14_2814 ();
 sg13g2_decap_8 FILLER_14_2821 ();
 sg13g2_decap_4 FILLER_14_2863 ();
 sg13g2_fill_2 FILLER_14_2867 ();
 sg13g2_decap_8 FILLER_14_2895 ();
 sg13g2_decap_8 FILLER_14_2902 ();
 sg13g2_decap_8 FILLER_14_2909 ();
 sg13g2_decap_4 FILLER_14_2916 ();
 sg13g2_fill_1 FILLER_14_2920 ();
 sg13g2_decap_8 FILLER_14_2955 ();
 sg13g2_decap_8 FILLER_14_2962 ();
 sg13g2_decap_8 FILLER_14_2969 ();
 sg13g2_fill_2 FILLER_14_2976 ();
 sg13g2_fill_1 FILLER_14_2978 ();
 sg13g2_decap_8 FILLER_14_3007 ();
 sg13g2_decap_8 FILLER_14_3014 ();
 sg13g2_decap_8 FILLER_14_3021 ();
 sg13g2_decap_4 FILLER_14_3038 ();
 sg13g2_decap_8 FILLER_14_3068 ();
 sg13g2_fill_2 FILLER_14_3075 ();
 sg13g2_fill_1 FILLER_14_3077 ();
 sg13g2_decap_8 FILLER_14_3109 ();
 sg13g2_decap_8 FILLER_14_3116 ();
 sg13g2_decap_8 FILLER_14_3123 ();
 sg13g2_decap_4 FILLER_14_3130 ();
 sg13g2_decap_8 FILLER_14_3173 ();
 sg13g2_decap_8 FILLER_14_3180 ();
 sg13g2_decap_4 FILLER_14_3187 ();
 sg13g2_decap_8 FILLER_14_3204 ();
 sg13g2_decap_8 FILLER_14_3211 ();
 sg13g2_decap_8 FILLER_14_3218 ();
 sg13g2_decap_8 FILLER_14_3225 ();
 sg13g2_decap_8 FILLER_14_3232 ();
 sg13g2_fill_2 FILLER_14_3239 ();
 sg13g2_fill_1 FILLER_14_3259 ();
 sg13g2_decap_8 FILLER_14_3265 ();
 sg13g2_decap_8 FILLER_14_3272 ();
 sg13g2_decap_8 FILLER_14_3279 ();
 sg13g2_decap_8 FILLER_14_3286 ();
 sg13g2_decap_8 FILLER_14_3293 ();
 sg13g2_decap_8 FILLER_14_3300 ();
 sg13g2_decap_8 FILLER_14_3307 ();
 sg13g2_decap_8 FILLER_14_3314 ();
 sg13g2_decap_8 FILLER_14_3321 ();
 sg13g2_decap_4 FILLER_14_3328 ();
 sg13g2_fill_1 FILLER_14_3332 ();
 sg13g2_decap_8 FILLER_14_3353 ();
 sg13g2_decap_8 FILLER_14_3360 ();
 sg13g2_decap_8 FILLER_14_3367 ();
 sg13g2_decap_8 FILLER_14_3374 ();
 sg13g2_fill_1 FILLER_14_3381 ();
 sg13g2_decap_8 FILLER_14_3400 ();
 sg13g2_decap_8 FILLER_14_3407 ();
 sg13g2_decap_8 FILLER_14_3414 ();
 sg13g2_decap_4 FILLER_14_3421 ();
 sg13g2_decap_4 FILLER_14_3429 ();
 sg13g2_fill_2 FILLER_14_3433 ();
 sg13g2_decap_8 FILLER_14_3443 ();
 sg13g2_fill_2 FILLER_14_3450 ();
 sg13g2_decap_8 FILLER_14_3478 ();
 sg13g2_decap_8 FILLER_14_3485 ();
 sg13g2_decap_8 FILLER_14_3492 ();
 sg13g2_decap_8 FILLER_14_3499 ();
 sg13g2_decap_8 FILLER_14_3506 ();
 sg13g2_decap_8 FILLER_14_3513 ();
 sg13g2_decap_8 FILLER_14_3520 ();
 sg13g2_decap_8 FILLER_14_3527 ();
 sg13g2_decap_8 FILLER_14_3534 ();
 sg13g2_decap_8 FILLER_14_3541 ();
 sg13g2_decap_8 FILLER_14_3548 ();
 sg13g2_decap_8 FILLER_14_3555 ();
 sg13g2_decap_8 FILLER_14_3562 ();
 sg13g2_decap_8 FILLER_14_3569 ();
 sg13g2_decap_4 FILLER_14_3576 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_fill_2 FILLER_15_21 ();
 sg13g2_fill_2 FILLER_15_41 ();
 sg13g2_decap_8 FILLER_15_52 ();
 sg13g2_decap_8 FILLER_15_59 ();
 sg13g2_decap_4 FILLER_15_66 ();
 sg13g2_fill_1 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_97 ();
 sg13g2_decap_8 FILLER_15_104 ();
 sg13g2_decap_8 FILLER_15_111 ();
 sg13g2_decap_8 FILLER_15_118 ();
 sg13g2_decap_8 FILLER_15_125 ();
 sg13g2_decap_8 FILLER_15_132 ();
 sg13g2_decap_8 FILLER_15_139 ();
 sg13g2_decap_8 FILLER_15_146 ();
 sg13g2_decap_8 FILLER_15_153 ();
 sg13g2_decap_8 FILLER_15_160 ();
 sg13g2_decap_8 FILLER_15_167 ();
 sg13g2_decap_8 FILLER_15_174 ();
 sg13g2_decap_8 FILLER_15_181 ();
 sg13g2_decap_8 FILLER_15_188 ();
 sg13g2_decap_8 FILLER_15_195 ();
 sg13g2_decap_8 FILLER_15_202 ();
 sg13g2_decap_8 FILLER_15_209 ();
 sg13g2_decap_8 FILLER_15_230 ();
 sg13g2_fill_2 FILLER_15_237 ();
 sg13g2_decap_8 FILLER_15_243 ();
 sg13g2_decap_8 FILLER_15_250 ();
 sg13g2_decap_8 FILLER_15_257 ();
 sg13g2_fill_1 FILLER_15_264 ();
 sg13g2_decap_8 FILLER_15_270 ();
 sg13g2_decap_8 FILLER_15_277 ();
 sg13g2_decap_8 FILLER_15_284 ();
 sg13g2_decap_8 FILLER_15_291 ();
 sg13g2_decap_8 FILLER_15_298 ();
 sg13g2_decap_8 FILLER_15_305 ();
 sg13g2_fill_1 FILLER_15_312 ();
 sg13g2_decap_8 FILLER_15_376 ();
 sg13g2_decap_4 FILLER_15_383 ();
 sg13g2_fill_2 FILLER_15_387 ();
 sg13g2_decap_4 FILLER_15_393 ();
 sg13g2_decap_8 FILLER_15_401 ();
 sg13g2_decap_8 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_15_415 ();
 sg13g2_decap_8 FILLER_15_422 ();
 sg13g2_decap_8 FILLER_15_429 ();
 sg13g2_decap_8 FILLER_15_436 ();
 sg13g2_decap_8 FILLER_15_443 ();
 sg13g2_decap_8 FILLER_15_450 ();
 sg13g2_decap_8 FILLER_15_457 ();
 sg13g2_decap_8 FILLER_15_464 ();
 sg13g2_decap_8 FILLER_15_471 ();
 sg13g2_decap_4 FILLER_15_478 ();
 sg13g2_decap_8 FILLER_15_492 ();
 sg13g2_decap_8 FILLER_15_499 ();
 sg13g2_decap_8 FILLER_15_506 ();
 sg13g2_fill_2 FILLER_15_513 ();
 sg13g2_fill_1 FILLER_15_515 ();
 sg13g2_decap_8 FILLER_15_531 ();
 sg13g2_decap_4 FILLER_15_538 ();
 sg13g2_fill_2 FILLER_15_542 ();
 sg13g2_decap_8 FILLER_15_549 ();
 sg13g2_decap_8 FILLER_15_556 ();
 sg13g2_decap_8 FILLER_15_563 ();
 sg13g2_decap_8 FILLER_15_570 ();
 sg13g2_fill_1 FILLER_15_577 ();
 sg13g2_decap_8 FILLER_15_588 ();
 sg13g2_decap_8 FILLER_15_595 ();
 sg13g2_decap_8 FILLER_15_602 ();
 sg13g2_decap_8 FILLER_15_609 ();
 sg13g2_decap_8 FILLER_15_616 ();
 sg13g2_decap_8 FILLER_15_623 ();
 sg13g2_decap_8 FILLER_15_630 ();
 sg13g2_decap_8 FILLER_15_637 ();
 sg13g2_decap_8 FILLER_15_644 ();
 sg13g2_fill_1 FILLER_15_670 ();
 sg13g2_fill_1 FILLER_15_675 ();
 sg13g2_fill_2 FILLER_15_679 ();
 sg13g2_fill_2 FILLER_15_691 ();
 sg13g2_fill_1 FILLER_15_693 ();
 sg13g2_fill_2 FILLER_15_704 ();
 sg13g2_fill_2 FILLER_15_716 ();
 sg13g2_fill_1 FILLER_15_718 ();
 sg13g2_decap_8 FILLER_15_724 ();
 sg13g2_fill_2 FILLER_15_731 ();
 sg13g2_decap_8 FILLER_15_743 ();
 sg13g2_decap_8 FILLER_15_750 ();
 sg13g2_decap_8 FILLER_15_757 ();
 sg13g2_decap_8 FILLER_15_764 ();
 sg13g2_decap_8 FILLER_15_771 ();
 sg13g2_decap_8 FILLER_15_778 ();
 sg13g2_decap_8 FILLER_15_785 ();
 sg13g2_decap_8 FILLER_15_792 ();
 sg13g2_decap_8 FILLER_15_799 ();
 sg13g2_decap_8 FILLER_15_806 ();
 sg13g2_decap_8 FILLER_15_813 ();
 sg13g2_decap_8 FILLER_15_820 ();
 sg13g2_decap_4 FILLER_15_827 ();
 sg13g2_fill_2 FILLER_15_841 ();
 sg13g2_decap_8 FILLER_15_869 ();
 sg13g2_decap_8 FILLER_15_876 ();
 sg13g2_decap_8 FILLER_15_883 ();
 sg13g2_decap_8 FILLER_15_890 ();
 sg13g2_decap_8 FILLER_15_897 ();
 sg13g2_decap_8 FILLER_15_904 ();
 sg13g2_decap_8 FILLER_15_911 ();
 sg13g2_decap_8 FILLER_15_918 ();
 sg13g2_decap_8 FILLER_15_925 ();
 sg13g2_decap_8 FILLER_15_932 ();
 sg13g2_fill_1 FILLER_15_939 ();
 sg13g2_decap_8 FILLER_15_976 ();
 sg13g2_decap_8 FILLER_15_983 ();
 sg13g2_decap_8 FILLER_15_990 ();
 sg13g2_decap_8 FILLER_15_997 ();
 sg13g2_fill_2 FILLER_15_1014 ();
 sg13g2_decap_8 FILLER_15_1042 ();
 sg13g2_decap_8 FILLER_15_1049 ();
 sg13g2_decap_8 FILLER_15_1056 ();
 sg13g2_decap_8 FILLER_15_1063 ();
 sg13g2_decap_8 FILLER_15_1070 ();
 sg13g2_decap_8 FILLER_15_1077 ();
 sg13g2_decap_8 FILLER_15_1084 ();
 sg13g2_decap_8 FILLER_15_1091 ();
 sg13g2_decap_4 FILLER_15_1098 ();
 sg13g2_fill_1 FILLER_15_1121 ();
 sg13g2_decap_8 FILLER_15_1151 ();
 sg13g2_decap_8 FILLER_15_1158 ();
 sg13g2_decap_8 FILLER_15_1165 ();
 sg13g2_decap_8 FILLER_15_1172 ();
 sg13g2_decap_4 FILLER_15_1179 ();
 sg13g2_fill_2 FILLER_15_1183 ();
 sg13g2_fill_2 FILLER_15_1190 ();
 sg13g2_fill_1 FILLER_15_1192 ();
 sg13g2_decap_8 FILLER_15_1201 ();
 sg13g2_decap_8 FILLER_15_1208 ();
 sg13g2_decap_8 FILLER_15_1215 ();
 sg13g2_fill_1 FILLER_15_1222 ();
 sg13g2_decap_8 FILLER_15_1236 ();
 sg13g2_decap_8 FILLER_15_1243 ();
 sg13g2_decap_8 FILLER_15_1250 ();
 sg13g2_decap_4 FILLER_15_1257 ();
 sg13g2_decap_8 FILLER_15_1266 ();
 sg13g2_decap_4 FILLER_15_1273 ();
 sg13g2_decap_4 FILLER_15_1282 ();
 sg13g2_fill_1 FILLER_15_1286 ();
 sg13g2_decap_8 FILLER_15_1290 ();
 sg13g2_fill_1 FILLER_15_1297 ();
 sg13g2_decap_4 FILLER_15_1304 ();
 sg13g2_fill_1 FILLER_15_1308 ();
 sg13g2_decap_8 FILLER_15_1314 ();
 sg13g2_decap_8 FILLER_15_1321 ();
 sg13g2_decap_4 FILLER_15_1328 ();
 sg13g2_fill_1 FILLER_15_1332 ();
 sg13g2_decap_8 FILLER_15_1338 ();
 sg13g2_decap_8 FILLER_15_1345 ();
 sg13g2_decap_8 FILLER_15_1352 ();
 sg13g2_decap_8 FILLER_15_1359 ();
 sg13g2_decap_8 FILLER_15_1366 ();
 sg13g2_decap_8 FILLER_15_1373 ();
 sg13g2_decap_8 FILLER_15_1380 ();
 sg13g2_decap_8 FILLER_15_1387 ();
 sg13g2_decap_8 FILLER_15_1394 ();
 sg13g2_decap_8 FILLER_15_1401 ();
 sg13g2_decap_8 FILLER_15_1408 ();
 sg13g2_decap_8 FILLER_15_1415 ();
 sg13g2_decap_4 FILLER_15_1422 ();
 sg13g2_fill_1 FILLER_15_1426 ();
 sg13g2_decap_8 FILLER_15_1453 ();
 sg13g2_fill_2 FILLER_15_1460 ();
 sg13g2_decap_8 FILLER_15_1467 ();
 sg13g2_decap_8 FILLER_15_1474 ();
 sg13g2_decap_8 FILLER_15_1481 ();
 sg13g2_decap_8 FILLER_15_1488 ();
 sg13g2_fill_2 FILLER_15_1495 ();
 sg13g2_decap_8 FILLER_15_1517 ();
 sg13g2_decap_8 FILLER_15_1524 ();
 sg13g2_decap_8 FILLER_15_1531 ();
 sg13g2_decap_8 FILLER_15_1538 ();
 sg13g2_fill_2 FILLER_15_1545 ();
 sg13g2_fill_2 FILLER_15_1569 ();
 sg13g2_decap_8 FILLER_15_1586 ();
 sg13g2_decap_8 FILLER_15_1593 ();
 sg13g2_decap_8 FILLER_15_1600 ();
 sg13g2_decap_8 FILLER_15_1607 ();
 sg13g2_fill_2 FILLER_15_1614 ();
 sg13g2_fill_1 FILLER_15_1616 ();
 sg13g2_decap_8 FILLER_15_1627 ();
 sg13g2_decap_8 FILLER_15_1634 ();
 sg13g2_decap_8 FILLER_15_1641 ();
 sg13g2_decap_8 FILLER_15_1648 ();
 sg13g2_decap_8 FILLER_15_1655 ();
 sg13g2_decap_8 FILLER_15_1662 ();
 sg13g2_decap_8 FILLER_15_1669 ();
 sg13g2_decap_8 FILLER_15_1676 ();
 sg13g2_fill_2 FILLER_15_1683 ();
 sg13g2_fill_1 FILLER_15_1685 ();
 sg13g2_decap_8 FILLER_15_1785 ();
 sg13g2_decap_8 FILLER_15_1792 ();
 sg13g2_decap_8 FILLER_15_1799 ();
 sg13g2_decap_8 FILLER_15_1806 ();
 sg13g2_decap_8 FILLER_15_1849 ();
 sg13g2_decap_8 FILLER_15_1856 ();
 sg13g2_decap_8 FILLER_15_1863 ();
 sg13g2_decap_8 FILLER_15_1870 ();
 sg13g2_fill_2 FILLER_15_1877 ();
 sg13g2_decap_8 FILLER_15_1892 ();
 sg13g2_decap_8 FILLER_15_1899 ();
 sg13g2_decap_8 FILLER_15_1906 ();
 sg13g2_decap_8 FILLER_15_1913 ();
 sg13g2_decap_8 FILLER_15_1920 ();
 sg13g2_fill_2 FILLER_15_1927 ();
 sg13g2_fill_1 FILLER_15_1929 ();
 sg13g2_decap_4 FILLER_15_1944 ();
 sg13g2_fill_2 FILLER_15_1955 ();
 sg13g2_fill_1 FILLER_15_1957 ();
 sg13g2_decap_8 FILLER_15_1975 ();
 sg13g2_decap_8 FILLER_15_1982 ();
 sg13g2_decap_8 FILLER_15_1989 ();
 sg13g2_decap_8 FILLER_15_1996 ();
 sg13g2_decap_8 FILLER_15_2003 ();
 sg13g2_decap_8 FILLER_15_2010 ();
 sg13g2_decap_8 FILLER_15_2017 ();
 sg13g2_decap_8 FILLER_15_2024 ();
 sg13g2_decap_8 FILLER_15_2031 ();
 sg13g2_decap_8 FILLER_15_2038 ();
 sg13g2_decap_8 FILLER_15_2045 ();
 sg13g2_decap_8 FILLER_15_2052 ();
 sg13g2_decap_8 FILLER_15_2059 ();
 sg13g2_decap_8 FILLER_15_2066 ();
 sg13g2_decap_8 FILLER_15_2073 ();
 sg13g2_decap_8 FILLER_15_2080 ();
 sg13g2_decap_8 FILLER_15_2087 ();
 sg13g2_fill_1 FILLER_15_2094 ();
 sg13g2_decap_8 FILLER_15_2103 ();
 sg13g2_decap_8 FILLER_15_2110 ();
 sg13g2_decap_8 FILLER_15_2117 ();
 sg13g2_decap_8 FILLER_15_2124 ();
 sg13g2_decap_8 FILLER_15_2131 ();
 sg13g2_decap_8 FILLER_15_2138 ();
 sg13g2_decap_8 FILLER_15_2153 ();
 sg13g2_decap_8 FILLER_15_2160 ();
 sg13g2_decap_8 FILLER_15_2167 ();
 sg13g2_decap_8 FILLER_15_2174 ();
 sg13g2_fill_1 FILLER_15_2191 ();
 sg13g2_decap_8 FILLER_15_2218 ();
 sg13g2_decap_8 FILLER_15_2225 ();
 sg13g2_decap_4 FILLER_15_2232 ();
 sg13g2_fill_2 FILLER_15_2236 ();
 sg13g2_decap_8 FILLER_15_2264 ();
 sg13g2_decap_8 FILLER_15_2271 ();
 sg13g2_fill_1 FILLER_15_2278 ();
 sg13g2_decap_8 FILLER_15_2305 ();
 sg13g2_decap_8 FILLER_15_2312 ();
 sg13g2_decap_8 FILLER_15_2319 ();
 sg13g2_decap_8 FILLER_15_2326 ();
 sg13g2_decap_8 FILLER_15_2333 ();
 sg13g2_decap_8 FILLER_15_2340 ();
 sg13g2_decap_8 FILLER_15_2347 ();
 sg13g2_decap_8 FILLER_15_2354 ();
 sg13g2_decap_4 FILLER_15_2361 ();
 sg13g2_fill_1 FILLER_15_2365 ();
 sg13g2_decap_8 FILLER_15_2371 ();
 sg13g2_decap_8 FILLER_15_2404 ();
 sg13g2_decap_8 FILLER_15_2411 ();
 sg13g2_decap_8 FILLER_15_2418 ();
 sg13g2_decap_8 FILLER_15_2425 ();
 sg13g2_decap_8 FILLER_15_2432 ();
 sg13g2_decap_8 FILLER_15_2439 ();
 sg13g2_decap_8 FILLER_15_2446 ();
 sg13g2_decap_8 FILLER_15_2453 ();
 sg13g2_decap_4 FILLER_15_2460 ();
 sg13g2_fill_2 FILLER_15_2464 ();
 sg13g2_decap_8 FILLER_15_2492 ();
 sg13g2_decap_8 FILLER_15_2499 ();
 sg13g2_decap_8 FILLER_15_2506 ();
 sg13g2_decap_8 FILLER_15_2513 ();
 sg13g2_decap_8 FILLER_15_2520 ();
 sg13g2_fill_2 FILLER_15_2527 ();
 sg13g2_decap_8 FILLER_15_2539 ();
 sg13g2_decap_8 FILLER_15_2546 ();
 sg13g2_decap_8 FILLER_15_2553 ();
 sg13g2_decap_8 FILLER_15_2560 ();
 sg13g2_decap_8 FILLER_15_2567 ();
 sg13g2_decap_8 FILLER_15_2574 ();
 sg13g2_decap_8 FILLER_15_2581 ();
 sg13g2_decap_8 FILLER_15_2588 ();
 sg13g2_decap_8 FILLER_15_2595 ();
 sg13g2_decap_8 FILLER_15_2602 ();
 sg13g2_decap_8 FILLER_15_2609 ();
 sg13g2_decap_4 FILLER_15_2616 ();
 sg13g2_fill_2 FILLER_15_2620 ();
 sg13g2_decap_8 FILLER_15_2633 ();
 sg13g2_decap_8 FILLER_15_2640 ();
 sg13g2_decap_8 FILLER_15_2647 ();
 sg13g2_decap_8 FILLER_15_2654 ();
 sg13g2_decap_8 FILLER_15_2661 ();
 sg13g2_decap_8 FILLER_15_2668 ();
 sg13g2_decap_8 FILLER_15_2675 ();
 sg13g2_decap_8 FILLER_15_2682 ();
 sg13g2_decap_8 FILLER_15_2689 ();
 sg13g2_decap_8 FILLER_15_2696 ();
 sg13g2_decap_8 FILLER_15_2703 ();
 sg13g2_decap_8 FILLER_15_2710 ();
 sg13g2_decap_8 FILLER_15_2717 ();
 sg13g2_decap_8 FILLER_15_2724 ();
 sg13g2_decap_8 FILLER_15_2731 ();
 sg13g2_decap_8 FILLER_15_2738 ();
 sg13g2_decap_8 FILLER_15_2745 ();
 sg13g2_decap_8 FILLER_15_2752 ();
 sg13g2_fill_2 FILLER_15_2759 ();
 sg13g2_decap_8 FILLER_15_2791 ();
 sg13g2_decap_8 FILLER_15_2798 ();
 sg13g2_decap_8 FILLER_15_2805 ();
 sg13g2_decap_8 FILLER_15_2812 ();
 sg13g2_decap_8 FILLER_15_2819 ();
 sg13g2_fill_1 FILLER_15_2826 ();
 sg13g2_decap_4 FILLER_15_2832 ();
 sg13g2_decap_8 FILLER_15_2839 ();
 sg13g2_decap_4 FILLER_15_2846 ();
 sg13g2_decap_8 FILLER_15_2860 ();
 sg13g2_decap_8 FILLER_15_2867 ();
 sg13g2_fill_2 FILLER_15_2874 ();
 sg13g2_decap_8 FILLER_15_2889 ();
 sg13g2_decap_8 FILLER_15_2896 ();
 sg13g2_decap_8 FILLER_15_2903 ();
 sg13g2_decap_8 FILLER_15_2910 ();
 sg13g2_decap_4 FILLER_15_2917 ();
 sg13g2_fill_1 FILLER_15_2921 ();
 sg13g2_decap_8 FILLER_15_2947 ();
 sg13g2_decap_8 FILLER_15_2954 ();
 sg13g2_decap_8 FILLER_15_2961 ();
 sg13g2_decap_8 FILLER_15_2968 ();
 sg13g2_fill_2 FILLER_15_2975 ();
 sg13g2_fill_1 FILLER_15_2977 ();
 sg13g2_decap_8 FILLER_15_3004 ();
 sg13g2_decap_8 FILLER_15_3011 ();
 sg13g2_decap_8 FILLER_15_3018 ();
 sg13g2_decap_8 FILLER_15_3025 ();
 sg13g2_decap_8 FILLER_15_3032 ();
 sg13g2_fill_2 FILLER_15_3039 ();
 sg13g2_fill_1 FILLER_15_3041 ();
 sg13g2_decap_8 FILLER_15_3060 ();
 sg13g2_decap_8 FILLER_15_3067 ();
 sg13g2_fill_2 FILLER_15_3074 ();
 sg13g2_fill_1 FILLER_15_3076 ();
 sg13g2_decap_8 FILLER_15_3107 ();
 sg13g2_decap_8 FILLER_15_3114 ();
 sg13g2_decap_8 FILLER_15_3121 ();
 sg13g2_decap_8 FILLER_15_3128 ();
 sg13g2_decap_8 FILLER_15_3135 ();
 sg13g2_fill_2 FILLER_15_3142 ();
 sg13g2_fill_1 FILLER_15_3144 ();
 sg13g2_decap_8 FILLER_15_3171 ();
 sg13g2_decap_8 FILLER_15_3204 ();
 sg13g2_decap_8 FILLER_15_3211 ();
 sg13g2_decap_8 FILLER_15_3218 ();
 sg13g2_decap_8 FILLER_15_3225 ();
 sg13g2_decap_4 FILLER_15_3232 ();
 sg13g2_decap_8 FILLER_15_3270 ();
 sg13g2_decap_8 FILLER_15_3277 ();
 sg13g2_decap_8 FILLER_15_3284 ();
 sg13g2_decap_4 FILLER_15_3291 ();
 sg13g2_decap_8 FILLER_15_3305 ();
 sg13g2_decap_8 FILLER_15_3312 ();
 sg13g2_decap_4 FILLER_15_3319 ();
 sg13g2_decap_8 FILLER_15_3364 ();
 sg13g2_decap_8 FILLER_15_3371 ();
 sg13g2_decap_8 FILLER_15_3378 ();
 sg13g2_decap_8 FILLER_15_3385 ();
 sg13g2_decap_8 FILLER_15_3397 ();
 sg13g2_fill_2 FILLER_15_3404 ();
 sg13g2_decap_8 FILLER_15_3426 ();
 sg13g2_fill_2 FILLER_15_3433 ();
 sg13g2_fill_1 FILLER_15_3435 ();
 sg13g2_fill_2 FILLER_15_3441 ();
 sg13g2_decap_8 FILLER_15_3447 ();
 sg13g2_decap_4 FILLER_15_3454 ();
 sg13g2_fill_2 FILLER_15_3467 ();
 sg13g2_fill_1 FILLER_15_3469 ();
 sg13g2_decap_8 FILLER_15_3483 ();
 sg13g2_decap_8 FILLER_15_3490 ();
 sg13g2_decap_8 FILLER_15_3497 ();
 sg13g2_decap_8 FILLER_15_3504 ();
 sg13g2_decap_8 FILLER_15_3511 ();
 sg13g2_decap_8 FILLER_15_3518 ();
 sg13g2_decap_8 FILLER_15_3525 ();
 sg13g2_decap_8 FILLER_15_3532 ();
 sg13g2_decap_8 FILLER_15_3539 ();
 sg13g2_decap_8 FILLER_15_3546 ();
 sg13g2_decap_8 FILLER_15_3553 ();
 sg13g2_decap_8 FILLER_15_3560 ();
 sg13g2_decap_8 FILLER_15_3567 ();
 sg13g2_decap_4 FILLER_15_3574 ();
 sg13g2_fill_2 FILLER_15_3578 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_4 FILLER_16_7 ();
 sg13g2_fill_1 FILLER_16_11 ();
 sg13g2_fill_1 FILLER_16_47 ();
 sg13g2_decap_8 FILLER_16_58 ();
 sg13g2_decap_8 FILLER_16_65 ();
 sg13g2_decap_8 FILLER_16_72 ();
 sg13g2_decap_4 FILLER_16_79 ();
 sg13g2_fill_2 FILLER_16_83 ();
 sg13g2_decap_4 FILLER_16_90 ();
 sg13g2_fill_2 FILLER_16_94 ();
 sg13g2_decap_8 FILLER_16_104 ();
 sg13g2_decap_8 FILLER_16_111 ();
 sg13g2_decap_8 FILLER_16_118 ();
 sg13g2_decap_8 FILLER_16_125 ();
 sg13g2_decap_8 FILLER_16_132 ();
 sg13g2_decap_4 FILLER_16_139 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_fill_2 FILLER_16_161 ();
 sg13g2_fill_2 FILLER_16_169 ();
 sg13g2_fill_1 FILLER_16_171 ();
 sg13g2_decap_8 FILLER_16_180 ();
 sg13g2_decap_8 FILLER_16_187 ();
 sg13g2_decap_8 FILLER_16_194 ();
 sg13g2_decap_8 FILLER_16_201 ();
 sg13g2_decap_8 FILLER_16_216 ();
 sg13g2_decap_8 FILLER_16_223 ();
 sg13g2_decap_8 FILLER_16_235 ();
 sg13g2_decap_8 FILLER_16_242 ();
 sg13g2_decap_8 FILLER_16_249 ();
 sg13g2_decap_8 FILLER_16_256 ();
 sg13g2_decap_8 FILLER_16_263 ();
 sg13g2_decap_8 FILLER_16_270 ();
 sg13g2_decap_8 FILLER_16_277 ();
 sg13g2_decap_8 FILLER_16_284 ();
 sg13g2_decap_8 FILLER_16_291 ();
 sg13g2_decap_8 FILLER_16_298 ();
 sg13g2_decap_8 FILLER_16_305 ();
 sg13g2_fill_2 FILLER_16_312 ();
 sg13g2_fill_1 FILLER_16_314 ();
 sg13g2_decap_4 FILLER_16_321 ();
 sg13g2_decap_4 FILLER_16_328 ();
 sg13g2_fill_1 FILLER_16_332 ();
 sg13g2_decap_8 FILLER_16_342 ();
 sg13g2_decap_8 FILLER_16_349 ();
 sg13g2_decap_4 FILLER_16_356 ();
 sg13g2_fill_1 FILLER_16_360 ();
 sg13g2_decap_8 FILLER_16_378 ();
 sg13g2_decap_8 FILLER_16_385 ();
 sg13g2_decap_8 FILLER_16_392 ();
 sg13g2_decap_8 FILLER_16_399 ();
 sg13g2_decap_8 FILLER_16_406 ();
 sg13g2_decap_4 FILLER_16_413 ();
 sg13g2_fill_1 FILLER_16_417 ();
 sg13g2_decap_8 FILLER_16_434 ();
 sg13g2_decap_8 FILLER_16_441 ();
 sg13g2_decap_8 FILLER_16_448 ();
 sg13g2_decap_8 FILLER_16_455 ();
 sg13g2_decap_8 FILLER_16_462 ();
 sg13g2_decap_8 FILLER_16_513 ();
 sg13g2_decap_8 FILLER_16_520 ();
 sg13g2_decap_8 FILLER_16_527 ();
 sg13g2_fill_2 FILLER_16_534 ();
 sg13g2_fill_1 FILLER_16_536 ();
 sg13g2_fill_2 FILLER_16_552 ();
 sg13g2_fill_1 FILLER_16_554 ();
 sg13g2_decap_8 FILLER_16_560 ();
 sg13g2_decap_4 FILLER_16_567 ();
 sg13g2_fill_2 FILLER_16_571 ();
 sg13g2_decap_8 FILLER_16_593 ();
 sg13g2_decap_8 FILLER_16_600 ();
 sg13g2_decap_8 FILLER_16_607 ();
 sg13g2_decap_8 FILLER_16_614 ();
 sg13g2_decap_8 FILLER_16_621 ();
 sg13g2_decap_8 FILLER_16_628 ();
 sg13g2_decap_4 FILLER_16_635 ();
 sg13g2_fill_2 FILLER_16_639 ();
 sg13g2_decap_8 FILLER_16_644 ();
 sg13g2_decap_4 FILLER_16_651 ();
 sg13g2_decap_8 FILLER_16_660 ();
 sg13g2_decap_8 FILLER_16_667 ();
 sg13g2_decap_8 FILLER_16_674 ();
 sg13g2_decap_4 FILLER_16_681 ();
 sg13g2_fill_1 FILLER_16_685 ();
 sg13g2_decap_4 FILLER_16_700 ();
 sg13g2_fill_1 FILLER_16_704 ();
 sg13g2_decap_4 FILLER_16_710 ();
 sg13g2_fill_1 FILLER_16_714 ();
 sg13g2_decap_8 FILLER_16_718 ();
 sg13g2_decap_8 FILLER_16_725 ();
 sg13g2_decap_8 FILLER_16_732 ();
 sg13g2_decap_8 FILLER_16_739 ();
 sg13g2_decap_8 FILLER_16_746 ();
 sg13g2_decap_8 FILLER_16_753 ();
 sg13g2_fill_2 FILLER_16_760 ();
 sg13g2_fill_1 FILLER_16_766 ();
 sg13g2_decap_8 FILLER_16_803 ();
 sg13g2_decap_8 FILLER_16_810 ();
 sg13g2_decap_8 FILLER_16_817 ();
 sg13g2_decap_8 FILLER_16_824 ();
 sg13g2_decap_8 FILLER_16_831 ();
 sg13g2_decap_8 FILLER_16_838 ();
 sg13g2_fill_2 FILLER_16_845 ();
 sg13g2_decap_8 FILLER_16_857 ();
 sg13g2_decap_8 FILLER_16_864 ();
 sg13g2_decap_8 FILLER_16_871 ();
 sg13g2_decap_8 FILLER_16_878 ();
 sg13g2_decap_8 FILLER_16_885 ();
 sg13g2_decap_8 FILLER_16_892 ();
 sg13g2_decap_8 FILLER_16_899 ();
 sg13g2_decap_8 FILLER_16_906 ();
 sg13g2_decap_8 FILLER_16_913 ();
 sg13g2_decap_8 FILLER_16_920 ();
 sg13g2_decap_8 FILLER_16_927 ();
 sg13g2_decap_8 FILLER_16_934 ();
 sg13g2_decap_8 FILLER_16_941 ();
 sg13g2_decap_8 FILLER_16_948 ();
 sg13g2_decap_8 FILLER_16_955 ();
 sg13g2_fill_1 FILLER_16_962 ();
 sg13g2_decap_8 FILLER_16_976 ();
 sg13g2_decap_8 FILLER_16_983 ();
 sg13g2_decap_8 FILLER_16_990 ();
 sg13g2_decap_8 FILLER_16_997 ();
 sg13g2_decap_8 FILLER_16_1004 ();
 sg13g2_decap_8 FILLER_16_1011 ();
 sg13g2_fill_2 FILLER_16_1018 ();
 sg13g2_fill_1 FILLER_16_1020 ();
 sg13g2_decap_8 FILLER_16_1057 ();
 sg13g2_decap_8 FILLER_16_1064 ();
 sg13g2_decap_4 FILLER_16_1071 ();
 sg13g2_fill_1 FILLER_16_1075 ();
 sg13g2_decap_8 FILLER_16_1086 ();
 sg13g2_decap_8 FILLER_16_1093 ();
 sg13g2_decap_8 FILLER_16_1100 ();
 sg13g2_decap_8 FILLER_16_1107 ();
 sg13g2_decap_4 FILLER_16_1114 ();
 sg13g2_fill_2 FILLER_16_1121 ();
 sg13g2_fill_1 FILLER_16_1123 ();
 sg13g2_decap_8 FILLER_16_1150 ();
 sg13g2_decap_4 FILLER_16_1157 ();
 sg13g2_fill_1 FILLER_16_1161 ();
 sg13g2_decap_4 FILLER_16_1180 ();
 sg13g2_fill_1 FILLER_16_1184 ();
 sg13g2_decap_8 FILLER_16_1189 ();
 sg13g2_decap_8 FILLER_16_1196 ();
 sg13g2_decap_8 FILLER_16_1203 ();
 sg13g2_decap_8 FILLER_16_1210 ();
 sg13g2_decap_8 FILLER_16_1217 ();
 sg13g2_decap_8 FILLER_16_1224 ();
 sg13g2_decap_8 FILLER_16_1231 ();
 sg13g2_decap_8 FILLER_16_1238 ();
 sg13g2_decap_8 FILLER_16_1245 ();
 sg13g2_fill_2 FILLER_16_1252 ();
 sg13g2_fill_1 FILLER_16_1258 ();
 sg13g2_fill_2 FILLER_16_1267 ();
 sg13g2_fill_2 FILLER_16_1272 ();
 sg13g2_decap_8 FILLER_16_1291 ();
 sg13g2_decap_4 FILLER_16_1298 ();
 sg13g2_fill_1 FILLER_16_1302 ();
 sg13g2_decap_8 FILLER_16_1308 ();
 sg13g2_decap_4 FILLER_16_1315 ();
 sg13g2_fill_1 FILLER_16_1319 ();
 sg13g2_decap_8 FILLER_16_1333 ();
 sg13g2_decap_8 FILLER_16_1340 ();
 sg13g2_fill_2 FILLER_16_1347 ();
 sg13g2_fill_1 FILLER_16_1349 ();
 sg13g2_decap_4 FILLER_16_1386 ();
 sg13g2_decap_8 FILLER_16_1398 ();
 sg13g2_decap_8 FILLER_16_1405 ();
 sg13g2_decap_4 FILLER_16_1412 ();
 sg13g2_fill_1 FILLER_16_1416 ();
 sg13g2_decap_8 FILLER_16_1422 ();
 sg13g2_decap_8 FILLER_16_1429 ();
 sg13g2_decap_8 FILLER_16_1436 ();
 sg13g2_fill_2 FILLER_16_1443 ();
 sg13g2_decap_8 FILLER_16_1453 ();
 sg13g2_decap_8 FILLER_16_1460 ();
 sg13g2_decap_8 FILLER_16_1467 ();
 sg13g2_decap_8 FILLER_16_1474 ();
 sg13g2_decap_8 FILLER_16_1481 ();
 sg13g2_decap_4 FILLER_16_1488 ();
 sg13g2_fill_2 FILLER_16_1492 ();
 sg13g2_fill_1 FILLER_16_1509 ();
 sg13g2_decap_8 FILLER_16_1519 ();
 sg13g2_decap_8 FILLER_16_1526 ();
 sg13g2_decap_8 FILLER_16_1533 ();
 sg13g2_decap_8 FILLER_16_1540 ();
 sg13g2_decap_8 FILLER_16_1547 ();
 sg13g2_fill_1 FILLER_16_1573 ();
 sg13g2_decap_8 FILLER_16_1579 ();
 sg13g2_decap_8 FILLER_16_1586 ();
 sg13g2_decap_8 FILLER_16_1593 ();
 sg13g2_decap_8 FILLER_16_1600 ();
 sg13g2_decap_8 FILLER_16_1607 ();
 sg13g2_decap_8 FILLER_16_1624 ();
 sg13g2_decap_8 FILLER_16_1631 ();
 sg13g2_decap_8 FILLER_16_1638 ();
 sg13g2_decap_8 FILLER_16_1645 ();
 sg13g2_decap_8 FILLER_16_1652 ();
 sg13g2_decap_8 FILLER_16_1659 ();
 sg13g2_decap_8 FILLER_16_1666 ();
 sg13g2_decap_8 FILLER_16_1673 ();
 sg13g2_fill_1 FILLER_16_1680 ();
 sg13g2_decap_8 FILLER_16_1686 ();
 sg13g2_decap_8 FILLER_16_1693 ();
 sg13g2_decap_8 FILLER_16_1700 ();
 sg13g2_fill_2 FILLER_16_1707 ();
 sg13g2_fill_2 FILLER_16_1713 ();
 sg13g2_fill_1 FILLER_16_1715 ();
 sg13g2_decap_8 FILLER_16_1719 ();
 sg13g2_decap_8 FILLER_16_1726 ();
 sg13g2_decap_4 FILLER_16_1733 ();
 sg13g2_fill_2 FILLER_16_1737 ();
 sg13g2_decap_8 FILLER_16_1749 ();
 sg13g2_decap_8 FILLER_16_1756 ();
 sg13g2_fill_2 FILLER_16_1763 ();
 sg13g2_fill_1 FILLER_16_1765 ();
 sg13g2_decap_8 FILLER_16_1769 ();
 sg13g2_decap_4 FILLER_16_1776 ();
 sg13g2_fill_2 FILLER_16_1780 ();
 sg13g2_decap_4 FILLER_16_1785 ();
 sg13g2_decap_8 FILLER_16_1792 ();
 sg13g2_decap_8 FILLER_16_1799 ();
 sg13g2_decap_4 FILLER_16_1806 ();
 sg13g2_decap_8 FILLER_16_1846 ();
 sg13g2_decap_8 FILLER_16_1853 ();
 sg13g2_decap_8 FILLER_16_1860 ();
 sg13g2_decap_8 FILLER_16_1867 ();
 sg13g2_decap_8 FILLER_16_1874 ();
 sg13g2_decap_8 FILLER_16_1881 ();
 sg13g2_decap_8 FILLER_16_1888 ();
 sg13g2_fill_2 FILLER_16_1895 ();
 sg13g2_fill_1 FILLER_16_1897 ();
 sg13g2_decap_4 FILLER_16_1902 ();
 sg13g2_fill_2 FILLER_16_1906 ();
 sg13g2_decap_4 FILLER_16_1913 ();
 sg13g2_decap_8 FILLER_16_1930 ();
 sg13g2_decap_8 FILLER_16_1937 ();
 sg13g2_decap_8 FILLER_16_1944 ();
 sg13g2_fill_2 FILLER_16_1991 ();
 sg13g2_decap_8 FILLER_16_2014 ();
 sg13g2_decap_8 FILLER_16_2021 ();
 sg13g2_fill_2 FILLER_16_2028 ();
 sg13g2_decap_4 FILLER_16_2040 ();
 sg13g2_decap_8 FILLER_16_2075 ();
 sg13g2_fill_1 FILLER_16_2082 ();
 sg13g2_decap_4 FILLER_16_2119 ();
 sg13g2_fill_2 FILLER_16_2123 ();
 sg13g2_decap_8 FILLER_16_2161 ();
 sg13g2_decap_8 FILLER_16_2168 ();
 sg13g2_decap_8 FILLER_16_2175 ();
 sg13g2_decap_8 FILLER_16_2182 ();
 sg13g2_decap_8 FILLER_16_2189 ();
 sg13g2_decap_8 FILLER_16_2196 ();
 sg13g2_decap_8 FILLER_16_2203 ();
 sg13g2_decap_8 FILLER_16_2210 ();
 sg13g2_decap_8 FILLER_16_2220 ();
 sg13g2_decap_8 FILLER_16_2227 ();
 sg13g2_decap_8 FILLER_16_2234 ();
 sg13g2_decap_8 FILLER_16_2241 ();
 sg13g2_decap_8 FILLER_16_2248 ();
 sg13g2_decap_8 FILLER_16_2255 ();
 sg13g2_fill_1 FILLER_16_2262 ();
 sg13g2_fill_2 FILLER_16_2268 ();
 sg13g2_fill_1 FILLER_16_2270 ();
 sg13g2_decap_8 FILLER_16_2297 ();
 sg13g2_decap_8 FILLER_16_2304 ();
 sg13g2_decap_8 FILLER_16_2311 ();
 sg13g2_decap_8 FILLER_16_2318 ();
 sg13g2_decap_8 FILLER_16_2325 ();
 sg13g2_fill_2 FILLER_16_2332 ();
 sg13g2_decap_8 FILLER_16_2378 ();
 sg13g2_decap_8 FILLER_16_2385 ();
 sg13g2_decap_8 FILLER_16_2392 ();
 sg13g2_decap_8 FILLER_16_2399 ();
 sg13g2_fill_2 FILLER_16_2406 ();
 sg13g2_decap_8 FILLER_16_2434 ();
 sg13g2_decap_8 FILLER_16_2441 ();
 sg13g2_decap_4 FILLER_16_2448 ();
 sg13g2_decap_8 FILLER_16_2488 ();
 sg13g2_decap_8 FILLER_16_2495 ();
 sg13g2_fill_2 FILLER_16_2502 ();
 sg13g2_fill_1 FILLER_16_2504 ();
 sg13g2_decap_8 FILLER_16_2513 ();
 sg13g2_decap_4 FILLER_16_2520 ();
 sg13g2_fill_1 FILLER_16_2524 ();
 sg13g2_decap_8 FILLER_16_2575 ();
 sg13g2_decap_8 FILLER_16_2582 ();
 sg13g2_decap_8 FILLER_16_2589 ();
 sg13g2_fill_2 FILLER_16_2596 ();
 sg13g2_fill_1 FILLER_16_2608 ();
 sg13g2_decap_8 FILLER_16_2635 ();
 sg13g2_decap_8 FILLER_16_2642 ();
 sg13g2_decap_8 FILLER_16_2649 ();
 sg13g2_decap_8 FILLER_16_2656 ();
 sg13g2_decap_8 FILLER_16_2663 ();
 sg13g2_decap_4 FILLER_16_2670 ();
 sg13g2_fill_2 FILLER_16_2674 ();
 sg13g2_decap_8 FILLER_16_2712 ();
 sg13g2_decap_8 FILLER_16_2719 ();
 sg13g2_decap_8 FILLER_16_2726 ();
 sg13g2_decap_8 FILLER_16_2733 ();
 sg13g2_decap_8 FILLER_16_2740 ();
 sg13g2_decap_8 FILLER_16_2747 ();
 sg13g2_decap_8 FILLER_16_2754 ();
 sg13g2_decap_4 FILLER_16_2761 ();
 sg13g2_fill_2 FILLER_16_2765 ();
 sg13g2_decap_8 FILLER_16_2803 ();
 sg13g2_decap_8 FILLER_16_2810 ();
 sg13g2_decap_4 FILLER_16_2817 ();
 sg13g2_fill_2 FILLER_16_2821 ();
 sg13g2_fill_2 FILLER_16_2858 ();
 sg13g2_fill_1 FILLER_16_2860 ();
 sg13g2_decap_8 FILLER_16_2887 ();
 sg13g2_decap_8 FILLER_16_2894 ();
 sg13g2_decap_8 FILLER_16_2901 ();
 sg13g2_decap_8 FILLER_16_2908 ();
 sg13g2_decap_8 FILLER_16_2915 ();
 sg13g2_fill_2 FILLER_16_2922 ();
 sg13g2_decap_8 FILLER_16_2942 ();
 sg13g2_fill_2 FILLER_16_2949 ();
 sg13g2_fill_1 FILLER_16_2951 ();
 sg13g2_decap_8 FILLER_16_2961 ();
 sg13g2_decap_8 FILLER_16_2968 ();
 sg13g2_decap_8 FILLER_16_2975 ();
 sg13g2_decap_8 FILLER_16_2982 ();
 sg13g2_decap_8 FILLER_16_2989 ();
 sg13g2_decap_8 FILLER_16_2996 ();
 sg13g2_decap_8 FILLER_16_3003 ();
 sg13g2_fill_2 FILLER_16_3010 ();
 sg13g2_fill_2 FILLER_16_3038 ();
 sg13g2_fill_1 FILLER_16_3040 ();
 sg13g2_decap_8 FILLER_16_3061 ();
 sg13g2_decap_8 FILLER_16_3068 ();
 sg13g2_decap_8 FILLER_16_3075 ();
 sg13g2_fill_2 FILLER_16_3082 ();
 sg13g2_fill_1 FILLER_16_3084 ();
 sg13g2_decap_4 FILLER_16_3090 ();
 sg13g2_fill_1 FILLER_16_3094 ();
 sg13g2_decap_8 FILLER_16_3101 ();
 sg13g2_decap_8 FILLER_16_3108 ();
 sg13g2_decap_8 FILLER_16_3115 ();
 sg13g2_decap_8 FILLER_16_3122 ();
 sg13g2_decap_8 FILLER_16_3129 ();
 sg13g2_decap_8 FILLER_16_3136 ();
 sg13g2_decap_8 FILLER_16_3143 ();
 sg13g2_decap_8 FILLER_16_3150 ();
 sg13g2_decap_4 FILLER_16_3157 ();
 sg13g2_fill_1 FILLER_16_3171 ();
 sg13g2_decap_8 FILLER_16_3181 ();
 sg13g2_decap_8 FILLER_16_3188 ();
 sg13g2_fill_2 FILLER_16_3195 ();
 sg13g2_decap_8 FILLER_16_3215 ();
 sg13g2_decap_8 FILLER_16_3222 ();
 sg13g2_decap_8 FILLER_16_3229 ();
 sg13g2_decap_8 FILLER_16_3271 ();
 sg13g2_decap_4 FILLER_16_3278 ();
 sg13g2_fill_1 FILLER_16_3282 ();
 sg13g2_decap_8 FILLER_16_3314 ();
 sg13g2_decap_8 FILLER_16_3321 ();
 sg13g2_fill_1 FILLER_16_3328 ();
 sg13g2_decap_8 FILLER_16_3349 ();
 sg13g2_decap_8 FILLER_16_3356 ();
 sg13g2_decap_8 FILLER_16_3363 ();
 sg13g2_decap_4 FILLER_16_3370 ();
 sg13g2_fill_2 FILLER_16_3374 ();
 sg13g2_decap_4 FILLER_16_3386 ();
 sg13g2_fill_2 FILLER_16_3390 ();
 sg13g2_decap_8 FILLER_16_3425 ();
 sg13g2_decap_8 FILLER_16_3432 ();
 sg13g2_decap_8 FILLER_16_3439 ();
 sg13g2_decap_4 FILLER_16_3446 ();
 sg13g2_fill_2 FILLER_16_3461 ();
 sg13g2_fill_1 FILLER_16_3463 ();
 sg13g2_decap_8 FILLER_16_3508 ();
 sg13g2_decap_8 FILLER_16_3515 ();
 sg13g2_decap_8 FILLER_16_3522 ();
 sg13g2_decap_8 FILLER_16_3529 ();
 sg13g2_decap_8 FILLER_16_3536 ();
 sg13g2_decap_8 FILLER_16_3543 ();
 sg13g2_decap_8 FILLER_16_3550 ();
 sg13g2_decap_8 FILLER_16_3557 ();
 sg13g2_decap_8 FILLER_16_3564 ();
 sg13g2_decap_8 FILLER_16_3571 ();
 sg13g2_fill_2 FILLER_16_3578 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_4 FILLER_17_21 ();
 sg13g2_fill_1 FILLER_17_25 ();
 sg13g2_decap_8 FILLER_17_60 ();
 sg13g2_decap_8 FILLER_17_67 ();
 sg13g2_decap_8 FILLER_17_74 ();
 sg13g2_decap_8 FILLER_17_81 ();
 sg13g2_decap_8 FILLER_17_88 ();
 sg13g2_fill_1 FILLER_17_95 ();
 sg13g2_decap_8 FILLER_17_122 ();
 sg13g2_decap_8 FILLER_17_129 ();
 sg13g2_decap_8 FILLER_17_136 ();
 sg13g2_decap_8 FILLER_17_143 ();
 sg13g2_decap_4 FILLER_17_150 ();
 sg13g2_fill_1 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_189 ();
 sg13g2_fill_1 FILLER_17_196 ();
 sg13g2_fill_2 FILLER_17_219 ();
 sg13g2_fill_1 FILLER_17_224 ();
 sg13g2_decap_8 FILLER_17_230 ();
 sg13g2_decap_4 FILLER_17_237 ();
 sg13g2_fill_1 FILLER_17_241 ();
 sg13g2_decap_8 FILLER_17_247 ();
 sg13g2_fill_1 FILLER_17_254 ();
 sg13g2_fill_1 FILLER_17_259 ();
 sg13g2_fill_1 FILLER_17_268 ();
 sg13g2_fill_1 FILLER_17_274 ();
 sg13g2_decap_8 FILLER_17_288 ();
 sg13g2_decap_8 FILLER_17_295 ();
 sg13g2_decap_8 FILLER_17_302 ();
 sg13g2_fill_1 FILLER_17_309 ();
 sg13g2_decap_8 FILLER_17_330 ();
 sg13g2_decap_8 FILLER_17_337 ();
 sg13g2_decap_8 FILLER_17_344 ();
 sg13g2_decap_4 FILLER_17_351 ();
 sg13g2_decap_8 FILLER_17_381 ();
 sg13g2_decap_8 FILLER_17_388 ();
 sg13g2_decap_8 FILLER_17_395 ();
 sg13g2_decap_8 FILLER_17_402 ();
 sg13g2_decap_4 FILLER_17_409 ();
 sg13g2_fill_2 FILLER_17_413 ();
 sg13g2_decap_8 FILLER_17_436 ();
 sg13g2_decap_8 FILLER_17_443 ();
 sg13g2_decap_8 FILLER_17_450 ();
 sg13g2_decap_8 FILLER_17_457 ();
 sg13g2_decap_8 FILLER_17_464 ();
 sg13g2_decap_8 FILLER_17_471 ();
 sg13g2_decap_4 FILLER_17_478 ();
 sg13g2_decap_8 FILLER_17_518 ();
 sg13g2_fill_2 FILLER_17_525 ();
 sg13g2_fill_1 FILLER_17_527 ();
 sg13g2_fill_2 FILLER_17_554 ();
 sg13g2_fill_2 FILLER_17_561 ();
 sg13g2_decap_8 FILLER_17_573 ();
 sg13g2_fill_2 FILLER_17_599 ();
 sg13g2_fill_1 FILLER_17_601 ();
 sg13g2_decap_8 FILLER_17_628 ();
 sg13g2_decap_4 FILLER_17_635 ();
 sg13g2_fill_1 FILLER_17_639 ();
 sg13g2_decap_8 FILLER_17_649 ();
 sg13g2_decap_8 FILLER_17_656 ();
 sg13g2_decap_8 FILLER_17_663 ();
 sg13g2_decap_8 FILLER_17_670 ();
 sg13g2_decap_8 FILLER_17_677 ();
 sg13g2_decap_8 FILLER_17_684 ();
 sg13g2_decap_4 FILLER_17_691 ();
 sg13g2_fill_1 FILLER_17_695 ();
 sg13g2_decap_8 FILLER_17_736 ();
 sg13g2_decap_8 FILLER_17_743 ();
 sg13g2_decap_4 FILLER_17_750 ();
 sg13g2_decap_8 FILLER_17_811 ();
 sg13g2_decap_8 FILLER_17_818 ();
 sg13g2_decap_8 FILLER_17_825 ();
 sg13g2_decap_8 FILLER_17_832 ();
 sg13g2_decap_8 FILLER_17_839 ();
 sg13g2_decap_8 FILLER_17_846 ();
 sg13g2_decap_8 FILLER_17_853 ();
 sg13g2_decap_8 FILLER_17_860 ();
 sg13g2_decap_8 FILLER_17_867 ();
 sg13g2_decap_8 FILLER_17_874 ();
 sg13g2_fill_2 FILLER_17_881 ();
 sg13g2_decap_4 FILLER_17_893 ();
 sg13g2_fill_1 FILLER_17_897 ();
 sg13g2_decap_8 FILLER_17_934 ();
 sg13g2_decap_8 FILLER_17_941 ();
 sg13g2_decap_8 FILLER_17_948 ();
 sg13g2_decap_8 FILLER_17_955 ();
 sg13g2_decap_8 FILLER_17_962 ();
 sg13g2_decap_8 FILLER_17_969 ();
 sg13g2_decap_8 FILLER_17_976 ();
 sg13g2_decap_8 FILLER_17_983 ();
 sg13g2_fill_2 FILLER_17_990 ();
 sg13g2_fill_1 FILLER_17_992 ();
 sg13g2_decap_8 FILLER_17_1003 ();
 sg13g2_decap_8 FILLER_17_1010 ();
 sg13g2_decap_8 FILLER_17_1017 ();
 sg13g2_decap_8 FILLER_17_1024 ();
 sg13g2_decap_8 FILLER_17_1031 ();
 sg13g2_decap_8 FILLER_17_1038 ();
 sg13g2_decap_4 FILLER_17_1045 ();
 sg13g2_fill_2 FILLER_17_1049 ();
 sg13g2_decap_4 FILLER_17_1057 ();
 sg13g2_fill_2 FILLER_17_1061 ();
 sg13g2_decap_8 FILLER_17_1089 ();
 sg13g2_decap_8 FILLER_17_1096 ();
 sg13g2_fill_2 FILLER_17_1103 ();
 sg13g2_decap_8 FILLER_17_1115 ();
 sg13g2_decap_8 FILLER_17_1122 ();
 sg13g2_decap_4 FILLER_17_1129 ();
 sg13g2_fill_1 FILLER_17_1133 ();
 sg13g2_decap_8 FILLER_17_1186 ();
 sg13g2_decap_8 FILLER_17_1193 ();
 sg13g2_decap_8 FILLER_17_1200 ();
 sg13g2_decap_8 FILLER_17_1207 ();
 sg13g2_decap_8 FILLER_17_1214 ();
 sg13g2_fill_2 FILLER_17_1221 ();
 sg13g2_fill_1 FILLER_17_1223 ();
 sg13g2_decap_8 FILLER_17_1232 ();
 sg13g2_decap_8 FILLER_17_1239 ();
 sg13g2_fill_2 FILLER_17_1246 ();
 sg13g2_decap_8 FILLER_17_1292 ();
 sg13g2_decap_8 FILLER_17_1299 ();
 sg13g2_decap_4 FILLER_17_1306 ();
 sg13g2_fill_1 FILLER_17_1310 ();
 sg13g2_decap_8 FILLER_17_1337 ();
 sg13g2_decap_8 FILLER_17_1344 ();
 sg13g2_fill_2 FILLER_17_1351 ();
 sg13g2_decap_8 FILLER_17_1394 ();
 sg13g2_fill_2 FILLER_17_1401 ();
 sg13g2_decap_8 FILLER_17_1408 ();
 sg13g2_decap_8 FILLER_17_1415 ();
 sg13g2_decap_8 FILLER_17_1422 ();
 sg13g2_decap_8 FILLER_17_1429 ();
 sg13g2_decap_4 FILLER_17_1467 ();
 sg13g2_fill_1 FILLER_17_1471 ();
 sg13g2_decap_8 FILLER_17_1482 ();
 sg13g2_decap_4 FILLER_17_1489 ();
 sg13g2_fill_1 FILLER_17_1493 ();
 sg13g2_decap_4 FILLER_17_1499 ();
 sg13g2_fill_1 FILLER_17_1503 ();
 sg13g2_decap_8 FILLER_17_1517 ();
 sg13g2_decap_8 FILLER_17_1524 ();
 sg13g2_decap_8 FILLER_17_1531 ();
 sg13g2_decap_8 FILLER_17_1538 ();
 sg13g2_decap_8 FILLER_17_1545 ();
 sg13g2_decap_4 FILLER_17_1552 ();
 sg13g2_fill_1 FILLER_17_1556 ();
 sg13g2_decap_8 FILLER_17_1568 ();
 sg13g2_decap_8 FILLER_17_1575 ();
 sg13g2_decap_8 FILLER_17_1582 ();
 sg13g2_decap_8 FILLER_17_1589 ();
 sg13g2_decap_8 FILLER_17_1596 ();
 sg13g2_decap_8 FILLER_17_1603 ();
 sg13g2_decap_4 FILLER_17_1610 ();
 sg13g2_fill_1 FILLER_17_1614 ();
 sg13g2_decap_8 FILLER_17_1651 ();
 sg13g2_decap_8 FILLER_17_1658 ();
 sg13g2_decap_8 FILLER_17_1665 ();
 sg13g2_decap_8 FILLER_17_1672 ();
 sg13g2_decap_8 FILLER_17_1679 ();
 sg13g2_decap_8 FILLER_17_1686 ();
 sg13g2_decap_8 FILLER_17_1693 ();
 sg13g2_decap_8 FILLER_17_1700 ();
 sg13g2_decap_8 FILLER_17_1707 ();
 sg13g2_decap_8 FILLER_17_1714 ();
 sg13g2_decap_8 FILLER_17_1721 ();
 sg13g2_decap_8 FILLER_17_1728 ();
 sg13g2_decap_8 FILLER_17_1735 ();
 sg13g2_decap_8 FILLER_17_1742 ();
 sg13g2_decap_8 FILLER_17_1749 ();
 sg13g2_fill_1 FILLER_17_1756 ();
 sg13g2_decap_8 FILLER_17_1760 ();
 sg13g2_decap_8 FILLER_17_1767 ();
 sg13g2_decap_8 FILLER_17_1774 ();
 sg13g2_decap_8 FILLER_17_1781 ();
 sg13g2_fill_2 FILLER_17_1788 ();
 sg13g2_fill_1 FILLER_17_1790 ();
 sg13g2_decap_8 FILLER_17_1794 ();
 sg13g2_decap_4 FILLER_17_1801 ();
 sg13g2_fill_1 FILLER_17_1805 ();
 sg13g2_fill_2 FILLER_17_1847 ();
 sg13g2_decap_8 FILLER_17_1857 ();
 sg13g2_decap_8 FILLER_17_1864 ();
 sg13g2_decap_8 FILLER_17_1871 ();
 sg13g2_fill_2 FILLER_17_1878 ();
 sg13g2_decap_4 FILLER_17_1893 ();
 sg13g2_fill_1 FILLER_17_1897 ();
 sg13g2_fill_2 FILLER_17_1912 ();
 sg13g2_fill_1 FILLER_17_1914 ();
 sg13g2_decap_8 FILLER_17_1929 ();
 sg13g2_decap_8 FILLER_17_1936 ();
 sg13g2_decap_8 FILLER_17_1943 ();
 sg13g2_decap_4 FILLER_17_1950 ();
 sg13g2_decap_8 FILLER_17_1964 ();
 sg13g2_decap_8 FILLER_17_1971 ();
 sg13g2_decap_8 FILLER_17_1978 ();
 sg13g2_decap_8 FILLER_17_1985 ();
 sg13g2_decap_4 FILLER_17_1992 ();
 sg13g2_fill_1 FILLER_17_1996 ();
 sg13g2_decap_4 FILLER_17_2054 ();
 sg13g2_decap_8 FILLER_17_2068 ();
 sg13g2_decap_8 FILLER_17_2075 ();
 sg13g2_decap_8 FILLER_17_2082 ();
 sg13g2_decap_8 FILLER_17_2089 ();
 sg13g2_decap_8 FILLER_17_2096 ();
 sg13g2_decap_8 FILLER_17_2103 ();
 sg13g2_decap_8 FILLER_17_2110 ();
 sg13g2_decap_8 FILLER_17_2117 ();
 sg13g2_decap_8 FILLER_17_2124 ();
 sg13g2_decap_8 FILLER_17_2131 ();
 sg13g2_decap_8 FILLER_17_2138 ();
 sg13g2_decap_4 FILLER_17_2145 ();
 sg13g2_fill_2 FILLER_17_2149 ();
 sg13g2_decap_8 FILLER_17_2161 ();
 sg13g2_decap_8 FILLER_17_2168 ();
 sg13g2_decap_8 FILLER_17_2175 ();
 sg13g2_decap_8 FILLER_17_2182 ();
 sg13g2_decap_8 FILLER_17_2189 ();
 sg13g2_fill_2 FILLER_17_2196 ();
 sg13g2_fill_1 FILLER_17_2198 ();
 sg13g2_decap_8 FILLER_17_2209 ();
 sg13g2_fill_1 FILLER_17_2216 ();
 sg13g2_decap_8 FILLER_17_2246 ();
 sg13g2_decap_8 FILLER_17_2253 ();
 sg13g2_fill_1 FILLER_17_2260 ();
 sg13g2_decap_8 FILLER_17_2274 ();
 sg13g2_decap_8 FILLER_17_2281 ();
 sg13g2_decap_8 FILLER_17_2288 ();
 sg13g2_decap_4 FILLER_17_2295 ();
 sg13g2_fill_2 FILLER_17_2299 ();
 sg13g2_decap_8 FILLER_17_2344 ();
 sg13g2_decap_8 FILLER_17_2351 ();
 sg13g2_decap_8 FILLER_17_2358 ();
 sg13g2_fill_2 FILLER_17_2365 ();
 sg13g2_fill_1 FILLER_17_2367 ();
 sg13g2_decap_8 FILLER_17_2384 ();
 sg13g2_decap_8 FILLER_17_2391 ();
 sg13g2_decap_8 FILLER_17_2398 ();
 sg13g2_fill_2 FILLER_17_2405 ();
 sg13g2_decap_8 FILLER_17_2443 ();
 sg13g2_decap_8 FILLER_17_2450 ();
 sg13g2_decap_8 FILLER_17_2457 ();
 sg13g2_decap_8 FILLER_17_2479 ();
 sg13g2_decap_8 FILLER_17_2486 ();
 sg13g2_decap_8 FILLER_17_2493 ();
 sg13g2_decap_8 FILLER_17_2500 ();
 sg13g2_decap_8 FILLER_17_2507 ();
 sg13g2_decap_8 FILLER_17_2514 ();
 sg13g2_decap_8 FILLER_17_2521 ();
 sg13g2_decap_8 FILLER_17_2528 ();
 sg13g2_decap_8 FILLER_17_2535 ();
 sg13g2_decap_4 FILLER_17_2542 ();
 sg13g2_fill_1 FILLER_17_2546 ();
 sg13g2_decap_4 FILLER_17_2552 ();
 sg13g2_fill_2 FILLER_17_2556 ();
 sg13g2_decap_8 FILLER_17_2584 ();
 sg13g2_fill_1 FILLER_17_2591 ();
 sg13g2_decap_4 FILLER_17_2618 ();
 sg13g2_fill_2 FILLER_17_2622 ();
 sg13g2_decap_8 FILLER_17_2632 ();
 sg13g2_decap_4 FILLER_17_2639 ();
 sg13g2_decap_4 FILLER_17_2651 ();
 sg13g2_fill_1 FILLER_17_2655 ();
 sg13g2_decap_8 FILLER_17_2682 ();
 sg13g2_decap_8 FILLER_17_2689 ();
 sg13g2_decap_8 FILLER_17_2696 ();
 sg13g2_decap_8 FILLER_17_2703 ();
 sg13g2_decap_8 FILLER_17_2710 ();
 sg13g2_decap_8 FILLER_17_2717 ();
 sg13g2_decap_8 FILLER_17_2724 ();
 sg13g2_decap_8 FILLER_17_2731 ();
 sg13g2_decap_8 FILLER_17_2738 ();
 sg13g2_decap_8 FILLER_17_2745 ();
 sg13g2_decap_8 FILLER_17_2752 ();
 sg13g2_decap_8 FILLER_17_2759 ();
 sg13g2_fill_2 FILLER_17_2766 ();
 sg13g2_decap_8 FILLER_17_2773 ();
 sg13g2_decap_8 FILLER_17_2780 ();
 sg13g2_decap_8 FILLER_17_2787 ();
 sg13g2_decap_8 FILLER_17_2794 ();
 sg13g2_decap_8 FILLER_17_2801 ();
 sg13g2_decap_8 FILLER_17_2808 ();
 sg13g2_decap_8 FILLER_17_2815 ();
 sg13g2_fill_1 FILLER_17_2822 ();
 sg13g2_decap_8 FILLER_17_2833 ();
 sg13g2_decap_8 FILLER_17_2840 ();
 sg13g2_decap_8 FILLER_17_2847 ();
 sg13g2_decap_4 FILLER_17_2854 ();
 sg13g2_fill_2 FILLER_17_2867 ();
 sg13g2_fill_1 FILLER_17_2869 ();
 sg13g2_decap_8 FILLER_17_2906 ();
 sg13g2_decap_8 FILLER_17_2913 ();
 sg13g2_decap_4 FILLER_17_2920 ();
 sg13g2_fill_1 FILLER_17_2924 ();
 sg13g2_fill_2 FILLER_17_2935 ();
 sg13g2_decap_8 FILLER_17_2963 ();
 sg13g2_decap_8 FILLER_17_2970 ();
 sg13g2_fill_2 FILLER_17_2977 ();
 sg13g2_fill_2 FILLER_17_2992 ();
 sg13g2_decap_8 FILLER_17_3004 ();
 sg13g2_decap_8 FILLER_17_3011 ();
 sg13g2_decap_8 FILLER_17_3018 ();
 sg13g2_decap_8 FILLER_17_3025 ();
 sg13g2_decap_8 FILLER_17_3035 ();
 sg13g2_decap_8 FILLER_17_3042 ();
 sg13g2_decap_8 FILLER_17_3049 ();
 sg13g2_decap_8 FILLER_17_3056 ();
 sg13g2_decap_8 FILLER_17_3063 ();
 sg13g2_decap_8 FILLER_17_3070 ();
 sg13g2_decap_8 FILLER_17_3077 ();
 sg13g2_decap_8 FILLER_17_3084 ();
 sg13g2_decap_8 FILLER_17_3091 ();
 sg13g2_decap_8 FILLER_17_3098 ();
 sg13g2_fill_2 FILLER_17_3105 ();
 sg13g2_decap_8 FILLER_17_3133 ();
 sg13g2_decap_8 FILLER_17_3140 ();
 sg13g2_decap_8 FILLER_17_3147 ();
 sg13g2_decap_8 FILLER_17_3154 ();
 sg13g2_decap_8 FILLER_17_3161 ();
 sg13g2_decap_8 FILLER_17_3168 ();
 sg13g2_decap_8 FILLER_17_3175 ();
 sg13g2_decap_8 FILLER_17_3182 ();
 sg13g2_decap_8 FILLER_17_3189 ();
 sg13g2_decap_8 FILLER_17_3196 ();
 sg13g2_decap_8 FILLER_17_3203 ();
 sg13g2_decap_8 FILLER_17_3210 ();
 sg13g2_decap_8 FILLER_17_3217 ();
 sg13g2_decap_8 FILLER_17_3224 ();
 sg13g2_decap_8 FILLER_17_3231 ();
 sg13g2_fill_1 FILLER_17_3238 ();
 sg13g2_decap_8 FILLER_17_3264 ();
 sg13g2_decap_8 FILLER_17_3271 ();
 sg13g2_decap_8 FILLER_17_3278 ();
 sg13g2_decap_8 FILLER_17_3285 ();
 sg13g2_decap_4 FILLER_17_3292 ();
 sg13g2_fill_1 FILLER_17_3306 ();
 sg13g2_decap_4 FILLER_17_3317 ();
 sg13g2_decap_8 FILLER_17_3325 ();
 sg13g2_decap_8 FILLER_17_3332 ();
 sg13g2_decap_8 FILLER_17_3339 ();
 sg13g2_decap_8 FILLER_17_3346 ();
 sg13g2_decap_8 FILLER_17_3353 ();
 sg13g2_decap_8 FILLER_17_3360 ();
 sg13g2_decap_4 FILLER_17_3372 ();
 sg13g2_fill_1 FILLER_17_3376 ();
 sg13g2_fill_1 FILLER_17_3382 ();
 sg13g2_decap_8 FILLER_17_3387 ();
 sg13g2_decap_8 FILLER_17_3394 ();
 sg13g2_decap_8 FILLER_17_3401 ();
 sg13g2_decap_8 FILLER_17_3408 ();
 sg13g2_decap_4 FILLER_17_3415 ();
 sg13g2_decap_8 FILLER_17_3424 ();
 sg13g2_fill_1 FILLER_17_3431 ();
 sg13g2_decap_8 FILLER_17_3440 ();
 sg13g2_decap_8 FILLER_17_3447 ();
 sg13g2_decap_8 FILLER_17_3454 ();
 sg13g2_decap_8 FILLER_17_3461 ();
 sg13g2_decap_4 FILLER_17_3468 ();
 sg13g2_decap_8 FILLER_17_3480 ();
 sg13g2_decap_8 FILLER_17_3487 ();
 sg13g2_decap_8 FILLER_17_3494 ();
 sg13g2_decap_8 FILLER_17_3501 ();
 sg13g2_decap_8 FILLER_17_3508 ();
 sg13g2_decap_8 FILLER_17_3515 ();
 sg13g2_decap_8 FILLER_17_3522 ();
 sg13g2_decap_8 FILLER_17_3529 ();
 sg13g2_decap_8 FILLER_17_3536 ();
 sg13g2_decap_8 FILLER_17_3543 ();
 sg13g2_decap_8 FILLER_17_3550 ();
 sg13g2_decap_8 FILLER_17_3557 ();
 sg13g2_decap_8 FILLER_17_3564 ();
 sg13g2_decap_8 FILLER_17_3571 ();
 sg13g2_fill_2 FILLER_17_3578 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_4 FILLER_18_21 ();
 sg13g2_fill_2 FILLER_18_25 ();
 sg13g2_decap_8 FILLER_18_53 ();
 sg13g2_decap_8 FILLER_18_60 ();
 sg13g2_decap_8 FILLER_18_67 ();
 sg13g2_decap_8 FILLER_18_74 ();
 sg13g2_decap_8 FILLER_18_81 ();
 sg13g2_decap_8 FILLER_18_88 ();
 sg13g2_fill_1 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_129 ();
 sg13g2_decap_8 FILLER_18_136 ();
 sg13g2_decap_8 FILLER_18_143 ();
 sg13g2_fill_2 FILLER_18_150 ();
 sg13g2_decap_4 FILLER_18_188 ();
 sg13g2_fill_2 FILLER_18_192 ();
 sg13g2_decap_4 FILLER_18_210 ();
 sg13g2_decap_4 FILLER_18_261 ();
 sg13g2_fill_2 FILLER_18_265 ();
 sg13g2_decap_8 FILLER_18_271 ();
 sg13g2_decap_8 FILLER_18_291 ();
 sg13g2_decap_8 FILLER_18_298 ();
 sg13g2_decap_8 FILLER_18_305 ();
 sg13g2_decap_4 FILLER_18_312 ();
 sg13g2_fill_2 FILLER_18_316 ();
 sg13g2_decap_8 FILLER_18_323 ();
 sg13g2_decap_8 FILLER_18_330 ();
 sg13g2_decap_8 FILLER_18_337 ();
 sg13g2_decap_8 FILLER_18_344 ();
 sg13g2_decap_8 FILLER_18_360 ();
 sg13g2_fill_2 FILLER_18_367 ();
 sg13g2_fill_1 FILLER_18_369 ();
 sg13g2_decap_8 FILLER_18_383 ();
 sg13g2_fill_1 FILLER_18_395 ();
 sg13g2_decap_8 FILLER_18_443 ();
 sg13g2_decap_8 FILLER_18_450 ();
 sg13g2_decap_8 FILLER_18_457 ();
 sg13g2_decap_8 FILLER_18_464 ();
 sg13g2_decap_8 FILLER_18_471 ();
 sg13g2_decap_4 FILLER_18_478 ();
 sg13g2_decap_8 FILLER_18_508 ();
 sg13g2_decap_8 FILLER_18_515 ();
 sg13g2_decap_8 FILLER_18_522 ();
 sg13g2_decap_8 FILLER_18_529 ();
 sg13g2_decap_4 FILLER_18_536 ();
 sg13g2_fill_1 FILLER_18_540 ();
 sg13g2_decap_8 FILLER_18_546 ();
 sg13g2_fill_1 FILLER_18_558 ();
 sg13g2_fill_2 FILLER_18_573 ();
 sg13g2_fill_1 FILLER_18_575 ();
 sg13g2_decap_4 FILLER_18_586 ();
 sg13g2_fill_2 FILLER_18_590 ();
 sg13g2_decap_8 FILLER_18_596 ();
 sg13g2_decap_8 FILLER_18_603 ();
 sg13g2_fill_2 FILLER_18_610 ();
 sg13g2_fill_1 FILLER_18_612 ();
 sg13g2_fill_2 FILLER_18_617 ();
 sg13g2_fill_1 FILLER_18_619 ();
 sg13g2_decap_8 FILLER_18_656 ();
 sg13g2_decap_8 FILLER_18_663 ();
 sg13g2_decap_8 FILLER_18_670 ();
 sg13g2_decap_8 FILLER_18_677 ();
 sg13g2_decap_8 FILLER_18_684 ();
 sg13g2_decap_8 FILLER_18_691 ();
 sg13g2_decap_8 FILLER_18_729 ();
 sg13g2_decap_8 FILLER_18_736 ();
 sg13g2_decap_8 FILLER_18_743 ();
 sg13g2_decap_8 FILLER_18_750 ();
 sg13g2_decap_8 FILLER_18_757 ();
 sg13g2_decap_8 FILLER_18_764 ();
 sg13g2_decap_4 FILLER_18_771 ();
 sg13g2_decap_8 FILLER_18_785 ();
 sg13g2_decap_4 FILLER_18_792 ();
 sg13g2_fill_1 FILLER_18_796 ();
 sg13g2_decap_8 FILLER_18_803 ();
 sg13g2_decap_4 FILLER_18_810 ();
 sg13g2_fill_2 FILLER_18_814 ();
 sg13g2_decap_4 FILLER_18_822 ();
 sg13g2_decap_8 FILLER_18_852 ();
 sg13g2_decap_8 FILLER_18_859 ();
 sg13g2_decap_8 FILLER_18_866 ();
 sg13g2_decap_8 FILLER_18_873 ();
 sg13g2_fill_2 FILLER_18_880 ();
 sg13g2_fill_1 FILLER_18_882 ();
 sg13g2_fill_1 FILLER_18_893 ();
 sg13g2_decap_8 FILLER_18_920 ();
 sg13g2_decap_8 FILLER_18_927 ();
 sg13g2_decap_8 FILLER_18_934 ();
 sg13g2_decap_8 FILLER_18_941 ();
 sg13g2_decap_8 FILLER_18_948 ();
 sg13g2_fill_2 FILLER_18_955 ();
 sg13g2_fill_1 FILLER_18_957 ();
 sg13g2_decap_8 FILLER_18_974 ();
 sg13g2_fill_1 FILLER_18_981 ();
 sg13g2_fill_2 FILLER_18_992 ();
 sg13g2_fill_1 FILLER_18_994 ();
 sg13g2_decap_8 FILLER_18_1021 ();
 sg13g2_decap_8 FILLER_18_1028 ();
 sg13g2_decap_8 FILLER_18_1035 ();
 sg13g2_decap_8 FILLER_18_1042 ();
 sg13g2_decap_8 FILLER_18_1059 ();
 sg13g2_decap_4 FILLER_18_1066 ();
 sg13g2_fill_2 FILLER_18_1070 ();
 sg13g2_decap_8 FILLER_18_1081 ();
 sg13g2_decap_8 FILLER_18_1088 ();
 sg13g2_decap_8 FILLER_18_1095 ();
 sg13g2_decap_8 FILLER_18_1102 ();
 sg13g2_decap_8 FILLER_18_1109 ();
 sg13g2_decap_8 FILLER_18_1116 ();
 sg13g2_decap_8 FILLER_18_1123 ();
 sg13g2_decap_4 FILLER_18_1130 ();
 sg13g2_decap_8 FILLER_18_1154 ();
 sg13g2_decap_8 FILLER_18_1161 ();
 sg13g2_decap_8 FILLER_18_1168 ();
 sg13g2_fill_1 FILLER_18_1175 ();
 sg13g2_decap_8 FILLER_18_1212 ();
 sg13g2_decap_8 FILLER_18_1219 ();
 sg13g2_decap_8 FILLER_18_1226 ();
 sg13g2_decap_8 FILLER_18_1233 ();
 sg13g2_decap_8 FILLER_18_1240 ();
 sg13g2_decap_8 FILLER_18_1247 ();
 sg13g2_decap_8 FILLER_18_1254 ();
 sg13g2_decap_8 FILLER_18_1261 ();
 sg13g2_decap_8 FILLER_18_1268 ();
 sg13g2_decap_4 FILLER_18_1280 ();
 sg13g2_decap_8 FILLER_18_1287 ();
 sg13g2_decap_8 FILLER_18_1294 ();
 sg13g2_decap_4 FILLER_18_1301 ();
 sg13g2_fill_1 FILLER_18_1305 ();
 sg13g2_decap_8 FILLER_18_1311 ();
 sg13g2_decap_8 FILLER_18_1318 ();
 sg13g2_decap_8 FILLER_18_1325 ();
 sg13g2_decap_4 FILLER_18_1332 ();
 sg13g2_fill_2 FILLER_18_1336 ();
 sg13g2_decap_8 FILLER_18_1346 ();
 sg13g2_decap_8 FILLER_18_1353 ();
 sg13g2_decap_8 FILLER_18_1360 ();
 sg13g2_decap_8 FILLER_18_1367 ();
 sg13g2_decap_8 FILLER_18_1374 ();
 sg13g2_decap_4 FILLER_18_1381 ();
 sg13g2_fill_2 FILLER_18_1385 ();
 sg13g2_decap_8 FILLER_18_1419 ();
 sg13g2_fill_2 FILLER_18_1426 ();
 sg13g2_decap_8 FILLER_18_1436 ();
 sg13g2_decap_8 FILLER_18_1443 ();
 sg13g2_decap_8 FILLER_18_1450 ();
 sg13g2_decap_4 FILLER_18_1457 ();
 sg13g2_fill_1 FILLER_18_1461 ();
 sg13g2_decap_8 FILLER_18_1493 ();
 sg13g2_decap_8 FILLER_18_1500 ();
 sg13g2_decap_8 FILLER_18_1507 ();
 sg13g2_decap_8 FILLER_18_1514 ();
 sg13g2_decap_8 FILLER_18_1521 ();
 sg13g2_decap_8 FILLER_18_1528 ();
 sg13g2_decap_8 FILLER_18_1535 ();
 sg13g2_decap_8 FILLER_18_1551 ();
 sg13g2_decap_8 FILLER_18_1558 ();
 sg13g2_decap_8 FILLER_18_1565 ();
 sg13g2_decap_8 FILLER_18_1572 ();
 sg13g2_decap_8 FILLER_18_1579 ();
 sg13g2_fill_2 FILLER_18_1586 ();
 sg13g2_fill_1 FILLER_18_1588 ();
 sg13g2_decap_8 FILLER_18_1599 ();
 sg13g2_decap_8 FILLER_18_1632 ();
 sg13g2_decap_8 FILLER_18_1639 ();
 sg13g2_decap_8 FILLER_18_1646 ();
 sg13g2_fill_1 FILLER_18_1653 ();
 sg13g2_fill_1 FILLER_18_1664 ();
 sg13g2_decap_8 FILLER_18_1691 ();
 sg13g2_decap_8 FILLER_18_1698 ();
 sg13g2_decap_4 FILLER_18_1705 ();
 sg13g2_decap_8 FILLER_18_1719 ();
 sg13g2_decap_8 FILLER_18_1726 ();
 sg13g2_decap_8 FILLER_18_1733 ();
 sg13g2_decap_8 FILLER_18_1740 ();
 sg13g2_decap_8 FILLER_18_1747 ();
 sg13g2_decap_8 FILLER_18_1754 ();
 sg13g2_decap_8 FILLER_18_1761 ();
 sg13g2_fill_2 FILLER_18_1768 ();
 sg13g2_decap_8 FILLER_18_1776 ();
 sg13g2_decap_8 FILLER_18_1783 ();
 sg13g2_decap_8 FILLER_18_1790 ();
 sg13g2_fill_2 FILLER_18_1797 ();
 sg13g2_fill_1 FILLER_18_1799 ();
 sg13g2_decap_8 FILLER_18_1806 ();
 sg13g2_decap_8 FILLER_18_1813 ();
 sg13g2_decap_8 FILLER_18_1820 ();
 sg13g2_decap_8 FILLER_18_1827 ();
 sg13g2_decap_8 FILLER_18_1834 ();
 sg13g2_fill_1 FILLER_18_1841 ();
 sg13g2_decap_8 FILLER_18_1847 ();
 sg13g2_decap_8 FILLER_18_1862 ();
 sg13g2_decap_8 FILLER_18_1869 ();
 sg13g2_fill_2 FILLER_18_1876 ();
 sg13g2_fill_1 FILLER_18_1878 ();
 sg13g2_decap_8 FILLER_18_1905 ();
 sg13g2_decap_8 FILLER_18_1918 ();
 sg13g2_decap_8 FILLER_18_1925 ();
 sg13g2_decap_8 FILLER_18_1932 ();
 sg13g2_decap_8 FILLER_18_1939 ();
 sg13g2_decap_8 FILLER_18_1946 ();
 sg13g2_fill_2 FILLER_18_1953 ();
 sg13g2_decap_8 FILLER_18_1981 ();
 sg13g2_decap_8 FILLER_18_1988 ();
 sg13g2_decap_8 FILLER_18_1995 ();
 sg13g2_decap_8 FILLER_18_2002 ();
 sg13g2_decap_8 FILLER_18_2009 ();
 sg13g2_decap_8 FILLER_18_2016 ();
 sg13g2_decap_8 FILLER_18_2023 ();
 sg13g2_decap_4 FILLER_18_2030 ();
 sg13g2_fill_1 FILLER_18_2034 ();
 sg13g2_decap_4 FILLER_18_2038 ();
 sg13g2_fill_1 FILLER_18_2042 ();
 sg13g2_decap_8 FILLER_18_2051 ();
 sg13g2_decap_8 FILLER_18_2063 ();
 sg13g2_decap_8 FILLER_18_2070 ();
 sg13g2_decap_8 FILLER_18_2077 ();
 sg13g2_decap_4 FILLER_18_2084 ();
 sg13g2_fill_1 FILLER_18_2088 ();
 sg13g2_decap_8 FILLER_18_2115 ();
 sg13g2_decap_8 FILLER_18_2122 ();
 sg13g2_decap_8 FILLER_18_2129 ();
 sg13g2_decap_8 FILLER_18_2136 ();
 sg13g2_decap_4 FILLER_18_2143 ();
 sg13g2_fill_1 FILLER_18_2147 ();
 sg13g2_decap_8 FILLER_18_2174 ();
 sg13g2_decap_8 FILLER_18_2181 ();
 sg13g2_decap_8 FILLER_18_2188 ();
 sg13g2_decap_4 FILLER_18_2195 ();
 sg13g2_fill_1 FILLER_18_2199 ();
 sg13g2_fill_2 FILLER_18_2209 ();
 sg13g2_decap_8 FILLER_18_2221 ();
 sg13g2_fill_2 FILLER_18_2228 ();
 sg13g2_fill_1 FILLER_18_2230 ();
 sg13g2_decap_8 FILLER_18_2237 ();
 sg13g2_decap_8 FILLER_18_2244 ();
 sg13g2_decap_8 FILLER_18_2251 ();
 sg13g2_decap_4 FILLER_18_2258 ();
 sg13g2_decap_8 FILLER_18_2272 ();
 sg13g2_decap_8 FILLER_18_2279 ();
 sg13g2_decap_8 FILLER_18_2286 ();
 sg13g2_decap_8 FILLER_18_2293 ();
 sg13g2_decap_8 FILLER_18_2300 ();
 sg13g2_decap_4 FILLER_18_2307 ();
 sg13g2_fill_1 FILLER_18_2311 ();
 sg13g2_decap_8 FILLER_18_2322 ();
 sg13g2_decap_8 FILLER_18_2329 ();
 sg13g2_decap_8 FILLER_18_2336 ();
 sg13g2_fill_2 FILLER_18_2343 ();
 sg13g2_fill_1 FILLER_18_2345 ();
 sg13g2_decap_8 FILLER_18_2383 ();
 sg13g2_decap_8 FILLER_18_2390 ();
 sg13g2_decap_8 FILLER_18_2397 ();
 sg13g2_decap_8 FILLER_18_2404 ();
 sg13g2_decap_8 FILLER_18_2411 ();
 sg13g2_fill_2 FILLER_18_2418 ();
 sg13g2_decap_8 FILLER_18_2434 ();
 sg13g2_decap_8 FILLER_18_2441 ();
 sg13g2_decap_8 FILLER_18_2448 ();
 sg13g2_decap_8 FILLER_18_2455 ();
 sg13g2_decap_4 FILLER_18_2462 ();
 sg13g2_fill_2 FILLER_18_2466 ();
 sg13g2_decap_8 FILLER_18_2482 ();
 sg13g2_decap_8 FILLER_18_2489 ();
 sg13g2_fill_2 FILLER_18_2496 ();
 sg13g2_fill_1 FILLER_18_2498 ();
 sg13g2_decap_8 FILLER_18_2525 ();
 sg13g2_fill_2 FILLER_18_2532 ();
 sg13g2_fill_1 FILLER_18_2534 ();
 sg13g2_decap_4 FILLER_18_2539 ();
 sg13g2_fill_1 FILLER_18_2543 ();
 sg13g2_decap_8 FILLER_18_2552 ();
 sg13g2_decap_8 FILLER_18_2559 ();
 sg13g2_fill_1 FILLER_18_2566 ();
 sg13g2_decap_8 FILLER_18_2577 ();
 sg13g2_decap_8 FILLER_18_2584 ();
 sg13g2_decap_8 FILLER_18_2591 ();
 sg13g2_decap_4 FILLER_18_2598 ();
 sg13g2_fill_1 FILLER_18_2602 ();
 sg13g2_decap_4 FILLER_18_2613 ();
 sg13g2_fill_1 FILLER_18_2617 ();
 sg13g2_fill_2 FILLER_18_2624 ();
 sg13g2_fill_1 FILLER_18_2626 ();
 sg13g2_decap_8 FILLER_18_2632 ();
 sg13g2_decap_8 FILLER_18_2642 ();
 sg13g2_decap_4 FILLER_18_2649 ();
 sg13g2_decap_4 FILLER_18_2656 ();
 sg13g2_fill_2 FILLER_18_2660 ();
 sg13g2_decap_8 FILLER_18_2672 ();
 sg13g2_decap_8 FILLER_18_2679 ();
 sg13g2_decap_8 FILLER_18_2686 ();
 sg13g2_fill_2 FILLER_18_2693 ();
 sg13g2_fill_1 FILLER_18_2695 ();
 sg13g2_decap_4 FILLER_18_2706 ();
 sg13g2_fill_2 FILLER_18_2710 ();
 sg13g2_decap_8 FILLER_18_2743 ();
 sg13g2_decap_8 FILLER_18_2750 ();
 sg13g2_decap_8 FILLER_18_2757 ();
 sg13g2_decap_8 FILLER_18_2774 ();
 sg13g2_decap_4 FILLER_18_2781 ();
 sg13g2_decap_8 FILLER_18_2793 ();
 sg13g2_decap_8 FILLER_18_2800 ();
 sg13g2_decap_4 FILLER_18_2807 ();
 sg13g2_fill_2 FILLER_18_2811 ();
 sg13g2_decap_8 FILLER_18_2839 ();
 sg13g2_decap_8 FILLER_18_2846 ();
 sg13g2_decap_8 FILLER_18_2853 ();
 sg13g2_decap_8 FILLER_18_2860 ();
 sg13g2_fill_2 FILLER_18_2867 ();
 sg13g2_decap_4 FILLER_18_2874 ();
 sg13g2_decap_8 FILLER_18_2887 ();
 sg13g2_decap_8 FILLER_18_2894 ();
 sg13g2_decap_8 FILLER_18_2901 ();
 sg13g2_decap_8 FILLER_18_2908 ();
 sg13g2_decap_4 FILLER_18_2915 ();
 sg13g2_fill_1 FILLER_18_2919 ();
 sg13g2_decap_8 FILLER_18_2946 ();
 sg13g2_decap_8 FILLER_18_2958 ();
 sg13g2_decap_8 FILLER_18_2965 ();
 sg13g2_decap_8 FILLER_18_3008 ();
 sg13g2_decap_8 FILLER_18_3015 ();
 sg13g2_fill_2 FILLER_18_3022 ();
 sg13g2_fill_1 FILLER_18_3024 ();
 sg13g2_decap_8 FILLER_18_3061 ();
 sg13g2_decap_8 FILLER_18_3068 ();
 sg13g2_decap_8 FILLER_18_3075 ();
 sg13g2_decap_8 FILLER_18_3082 ();
 sg13g2_decap_4 FILLER_18_3089 ();
 sg13g2_fill_2 FILLER_18_3093 ();
 sg13g2_decap_8 FILLER_18_3136 ();
 sg13g2_decap_8 FILLER_18_3143 ();
 sg13g2_decap_8 FILLER_18_3150 ();
 sg13g2_fill_2 FILLER_18_3157 ();
 sg13g2_decap_8 FILLER_18_3185 ();
 sg13g2_decap_8 FILLER_18_3192 ();
 sg13g2_decap_8 FILLER_18_3199 ();
 sg13g2_decap_8 FILLER_18_3216 ();
 sg13g2_decap_8 FILLER_18_3223 ();
 sg13g2_decap_8 FILLER_18_3230 ();
 sg13g2_decap_8 FILLER_18_3237 ();
 sg13g2_fill_2 FILLER_18_3244 ();
 sg13g2_decap_8 FILLER_18_3249 ();
 sg13g2_fill_1 FILLER_18_3256 ();
 sg13g2_decap_8 FILLER_18_3261 ();
 sg13g2_fill_2 FILLER_18_3268 ();
 sg13g2_fill_1 FILLER_18_3270 ();
 sg13g2_decap_8 FILLER_18_3275 ();
 sg13g2_decap_8 FILLER_18_3282 ();
 sg13g2_decap_8 FILLER_18_3289 ();
 sg13g2_fill_2 FILLER_18_3296 ();
 sg13g2_decap_8 FILLER_18_3346 ();
 sg13g2_decap_8 FILLER_18_3353 ();
 sg13g2_decap_8 FILLER_18_3360 ();
 sg13g2_decap_4 FILLER_18_3367 ();
 sg13g2_fill_2 FILLER_18_3371 ();
 sg13g2_decap_8 FILLER_18_3408 ();
 sg13g2_decap_8 FILLER_18_3415 ();
 sg13g2_fill_2 FILLER_18_3422 ();
 sg13g2_decap_8 FILLER_18_3450 ();
 sg13g2_decap_8 FILLER_18_3457 ();
 sg13g2_decap_8 FILLER_18_3464 ();
 sg13g2_decap_8 FILLER_18_3471 ();
 sg13g2_decap_8 FILLER_18_3478 ();
 sg13g2_decap_8 FILLER_18_3485 ();
 sg13g2_decap_8 FILLER_18_3492 ();
 sg13g2_decap_8 FILLER_18_3499 ();
 sg13g2_decap_8 FILLER_18_3532 ();
 sg13g2_decap_8 FILLER_18_3539 ();
 sg13g2_decap_4 FILLER_18_3546 ();
 sg13g2_fill_2 FILLER_18_3550 ();
 sg13g2_decap_8 FILLER_18_3560 ();
 sg13g2_decap_8 FILLER_18_3567 ();
 sg13g2_decap_4 FILLER_18_3574 ();
 sg13g2_fill_2 FILLER_18_3578 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_fill_2 FILLER_19_28 ();
 sg13g2_fill_1 FILLER_19_30 ();
 sg13g2_decap_8 FILLER_19_40 ();
 sg13g2_decap_8 FILLER_19_47 ();
 sg13g2_decap_8 FILLER_19_54 ();
 sg13g2_decap_8 FILLER_19_61 ();
 sg13g2_decap_8 FILLER_19_68 ();
 sg13g2_decap_8 FILLER_19_75 ();
 sg13g2_decap_8 FILLER_19_82 ();
 sg13g2_fill_2 FILLER_19_89 ();
 sg13g2_decap_8 FILLER_19_96 ();
 sg13g2_decap_4 FILLER_19_103 ();
 sg13g2_fill_1 FILLER_19_107 ();
 sg13g2_decap_4 FILLER_19_113 ();
 sg13g2_decap_8 FILLER_19_138 ();
 sg13g2_decap_8 FILLER_19_145 ();
 sg13g2_fill_2 FILLER_19_152 ();
 sg13g2_fill_1 FILLER_19_154 ();
 sg13g2_fill_1 FILLER_19_176 ();
 sg13g2_decap_8 FILLER_19_180 ();
 sg13g2_decap_8 FILLER_19_187 ();
 sg13g2_decap_8 FILLER_19_194 ();
 sg13g2_decap_8 FILLER_19_201 ();
 sg13g2_fill_2 FILLER_19_208 ();
 sg13g2_decap_8 FILLER_19_215 ();
 sg13g2_decap_8 FILLER_19_222 ();
 sg13g2_decap_8 FILLER_19_229 ();
 sg13g2_decap_8 FILLER_19_236 ();
 sg13g2_decap_8 FILLER_19_243 ();
 sg13g2_decap_4 FILLER_19_250 ();
 sg13g2_fill_2 FILLER_19_254 ();
 sg13g2_fill_2 FILLER_19_265 ();
 sg13g2_decap_4 FILLER_19_294 ();
 sg13g2_fill_1 FILLER_19_298 ();
 sg13g2_decap_8 FILLER_19_311 ();
 sg13g2_decap_8 FILLER_19_318 ();
 sg13g2_decap_8 FILLER_19_325 ();
 sg13g2_fill_2 FILLER_19_332 ();
 sg13g2_decap_8 FILLER_19_339 ();
 sg13g2_decap_4 FILLER_19_346 ();
 sg13g2_decap_4 FILLER_19_355 ();
 sg13g2_decap_8 FILLER_19_365 ();
 sg13g2_decap_8 FILLER_19_372 ();
 sg13g2_decap_8 FILLER_19_379 ();
 sg13g2_decap_8 FILLER_19_386 ();
 sg13g2_decap_8 FILLER_19_393 ();
 sg13g2_decap_8 FILLER_19_400 ();
 sg13g2_decap_8 FILLER_19_407 ();
 sg13g2_fill_2 FILLER_19_414 ();
 sg13g2_decap_8 FILLER_19_446 ();
 sg13g2_decap_8 FILLER_19_453 ();
 sg13g2_fill_2 FILLER_19_460 ();
 sg13g2_fill_1 FILLER_19_462 ();
 sg13g2_decap_8 FILLER_19_469 ();
 sg13g2_decap_8 FILLER_19_476 ();
 sg13g2_decap_8 FILLER_19_483 ();
 sg13g2_decap_8 FILLER_19_490 ();
 sg13g2_decap_8 FILLER_19_497 ();
 sg13g2_decap_8 FILLER_19_504 ();
 sg13g2_decap_8 FILLER_19_511 ();
 sg13g2_decap_8 FILLER_19_518 ();
 sg13g2_decap_8 FILLER_19_525 ();
 sg13g2_decap_8 FILLER_19_532 ();
 sg13g2_decap_8 FILLER_19_539 ();
 sg13g2_decap_8 FILLER_19_546 ();
 sg13g2_decap_8 FILLER_19_553 ();
 sg13g2_decap_8 FILLER_19_560 ();
 sg13g2_decap_8 FILLER_19_567 ();
 sg13g2_decap_4 FILLER_19_574 ();
 sg13g2_decap_8 FILLER_19_613 ();
 sg13g2_fill_2 FILLER_19_620 ();
 sg13g2_decap_8 FILLER_19_631 ();
 sg13g2_decap_8 FILLER_19_638 ();
 sg13g2_decap_8 FILLER_19_671 ();
 sg13g2_decap_8 FILLER_19_678 ();
 sg13g2_decap_8 FILLER_19_685 ();
 sg13g2_decap_8 FILLER_19_692 ();
 sg13g2_decap_8 FILLER_19_699 ();
 sg13g2_fill_2 FILLER_19_706 ();
 sg13g2_decap_8 FILLER_19_712 ();
 sg13g2_decap_8 FILLER_19_728 ();
 sg13g2_decap_8 FILLER_19_735 ();
 sg13g2_decap_8 FILLER_19_742 ();
 sg13g2_decap_8 FILLER_19_749 ();
 sg13g2_decap_8 FILLER_19_756 ();
 sg13g2_decap_8 FILLER_19_763 ();
 sg13g2_decap_8 FILLER_19_770 ();
 sg13g2_decap_8 FILLER_19_777 ();
 sg13g2_decap_8 FILLER_19_784 ();
 sg13g2_decap_8 FILLER_19_791 ();
 sg13g2_decap_8 FILLER_19_798 ();
 sg13g2_decap_8 FILLER_19_805 ();
 sg13g2_decap_4 FILLER_19_812 ();
 sg13g2_fill_1 FILLER_19_816 ();
 sg13g2_decap_8 FILLER_19_863 ();
 sg13g2_decap_8 FILLER_19_870 ();
 sg13g2_decap_8 FILLER_19_877 ();
 sg13g2_decap_8 FILLER_19_884 ();
 sg13g2_fill_2 FILLER_19_891 ();
 sg13g2_fill_1 FILLER_19_893 ();
 sg13g2_decap_8 FILLER_19_920 ();
 sg13g2_decap_8 FILLER_19_979 ();
 sg13g2_decap_8 FILLER_19_986 ();
 sg13g2_decap_4 FILLER_19_993 ();
 sg13g2_fill_2 FILLER_19_997 ();
 sg13g2_decap_8 FILLER_19_1025 ();
 sg13g2_decap_8 FILLER_19_1032 ();
 sg13g2_decap_8 FILLER_19_1039 ();
 sg13g2_decap_8 FILLER_19_1046 ();
 sg13g2_fill_2 FILLER_19_1053 ();
 sg13g2_fill_1 FILLER_19_1055 ();
 sg13g2_decap_8 FILLER_19_1092 ();
 sg13g2_decap_8 FILLER_19_1099 ();
 sg13g2_decap_8 FILLER_19_1106 ();
 sg13g2_decap_8 FILLER_19_1113 ();
 sg13g2_fill_2 FILLER_19_1120 ();
 sg13g2_decap_8 FILLER_19_1126 ();
 sg13g2_decap_8 FILLER_19_1133 ();
 sg13g2_decap_8 FILLER_19_1140 ();
 sg13g2_decap_8 FILLER_19_1147 ();
 sg13g2_decap_8 FILLER_19_1154 ();
 sg13g2_decap_8 FILLER_19_1161 ();
 sg13g2_decap_8 FILLER_19_1168 ();
 sg13g2_decap_8 FILLER_19_1175 ();
 sg13g2_decap_8 FILLER_19_1182 ();
 sg13g2_decap_8 FILLER_19_1189 ();
 sg13g2_decap_8 FILLER_19_1196 ();
 sg13g2_fill_2 FILLER_19_1203 ();
 sg13g2_fill_1 FILLER_19_1205 ();
 sg13g2_decap_8 FILLER_19_1216 ();
 sg13g2_decap_8 FILLER_19_1223 ();
 sg13g2_decap_8 FILLER_19_1230 ();
 sg13g2_decap_8 FILLER_19_1237 ();
 sg13g2_decap_8 FILLER_19_1244 ();
 sg13g2_decap_8 FILLER_19_1251 ();
 sg13g2_decap_8 FILLER_19_1258 ();
 sg13g2_fill_1 FILLER_19_1265 ();
 sg13g2_decap_8 FILLER_19_1275 ();
 sg13g2_decap_4 FILLER_19_1282 ();
 sg13g2_fill_2 FILLER_19_1286 ();
 sg13g2_decap_8 FILLER_19_1293 ();
 sg13g2_fill_1 FILLER_19_1300 ();
 sg13g2_decap_8 FILLER_19_1305 ();
 sg13g2_decap_8 FILLER_19_1312 ();
 sg13g2_decap_8 FILLER_19_1319 ();
 sg13g2_fill_2 FILLER_19_1326 ();
 sg13g2_fill_1 FILLER_19_1328 ();
 sg13g2_decap_8 FILLER_19_1345 ();
 sg13g2_decap_8 FILLER_19_1352 ();
 sg13g2_decap_8 FILLER_19_1359 ();
 sg13g2_decap_8 FILLER_19_1366 ();
 sg13g2_decap_8 FILLER_19_1373 ();
 sg13g2_decap_8 FILLER_19_1380 ();
 sg13g2_decap_8 FILLER_19_1387 ();
 sg13g2_decap_8 FILLER_19_1394 ();
 sg13g2_fill_2 FILLER_19_1401 ();
 sg13g2_fill_1 FILLER_19_1403 ();
 sg13g2_decap_4 FILLER_19_1408 ();
 sg13g2_decap_8 FILLER_19_1421 ();
 sg13g2_decap_4 FILLER_19_1428 ();
 sg13g2_fill_2 FILLER_19_1432 ();
 sg13g2_decap_8 FILLER_19_1444 ();
 sg13g2_decap_8 FILLER_19_1451 ();
 sg13g2_decap_8 FILLER_19_1458 ();
 sg13g2_decap_8 FILLER_19_1465 ();
 sg13g2_decap_4 FILLER_19_1472 ();
 sg13g2_fill_1 FILLER_19_1476 ();
 sg13g2_fill_2 FILLER_19_1480 ();
 sg13g2_fill_1 FILLER_19_1482 ();
 sg13g2_decap_8 FILLER_19_1492 ();
 sg13g2_fill_1 FILLER_19_1499 ();
 sg13g2_decap_8 FILLER_19_1510 ();
 sg13g2_decap_8 FILLER_19_1517 ();
 sg13g2_decap_8 FILLER_19_1524 ();
 sg13g2_fill_2 FILLER_19_1531 ();
 sg13g2_fill_1 FILLER_19_1533 ();
 sg13g2_decap_8 FILLER_19_1560 ();
 sg13g2_decap_8 FILLER_19_1567 ();
 sg13g2_fill_2 FILLER_19_1574 ();
 sg13g2_fill_1 FILLER_19_1576 ();
 sg13g2_decap_8 FILLER_19_1587 ();
 sg13g2_decap_8 FILLER_19_1604 ();
 sg13g2_decap_8 FILLER_19_1611 ();
 sg13g2_decap_8 FILLER_19_1618 ();
 sg13g2_decap_8 FILLER_19_1625 ();
 sg13g2_decap_8 FILLER_19_1632 ();
 sg13g2_decap_8 FILLER_19_1639 ();
 sg13g2_decap_8 FILLER_19_1646 ();
 sg13g2_fill_2 FILLER_19_1653 ();
 sg13g2_fill_1 FILLER_19_1665 ();
 sg13g2_decap_8 FILLER_19_1692 ();
 sg13g2_decap_8 FILLER_19_1699 ();
 sg13g2_fill_2 FILLER_19_1706 ();
 sg13g2_decap_8 FILLER_19_1734 ();
 sg13g2_decap_4 FILLER_19_1741 ();
 sg13g2_decap_8 FILLER_19_1797 ();
 sg13g2_decap_8 FILLER_19_1804 ();
 sg13g2_decap_8 FILLER_19_1811 ();
 sg13g2_decap_8 FILLER_19_1818 ();
 sg13g2_decap_8 FILLER_19_1825 ();
 sg13g2_decap_8 FILLER_19_1832 ();
 sg13g2_decap_8 FILLER_19_1842 ();
 sg13g2_decap_8 FILLER_19_1849 ();
 sg13g2_decap_8 FILLER_19_1856 ();
 sg13g2_decap_8 FILLER_19_1863 ();
 sg13g2_decap_8 FILLER_19_1870 ();
 sg13g2_decap_4 FILLER_19_1877 ();
 sg13g2_fill_1 FILLER_19_1881 ();
 sg13g2_decap_8 FILLER_19_1892 ();
 sg13g2_decap_4 FILLER_19_1899 ();
 sg13g2_fill_1 FILLER_19_1903 ();
 sg13g2_decap_8 FILLER_19_1910 ();
 sg13g2_fill_2 FILLER_19_1917 ();
 sg13g2_fill_1 FILLER_19_1919 ();
 sg13g2_decap_8 FILLER_19_1940 ();
 sg13g2_decap_8 FILLER_19_1947 ();
 sg13g2_decap_8 FILLER_19_1954 ();
 sg13g2_decap_8 FILLER_19_1961 ();
 sg13g2_decap_8 FILLER_19_1968 ();
 sg13g2_decap_8 FILLER_19_1975 ();
 sg13g2_decap_8 FILLER_19_1982 ();
 sg13g2_decap_8 FILLER_19_1989 ();
 sg13g2_decap_8 FILLER_19_1996 ();
 sg13g2_decap_8 FILLER_19_2003 ();
 sg13g2_decap_8 FILLER_19_2010 ();
 sg13g2_decap_8 FILLER_19_2017 ();
 sg13g2_decap_8 FILLER_19_2024 ();
 sg13g2_fill_2 FILLER_19_2031 ();
 sg13g2_fill_1 FILLER_19_2033 ();
 sg13g2_decap_8 FILLER_19_2039 ();
 sg13g2_decap_8 FILLER_19_2046 ();
 sg13g2_decap_8 FILLER_19_2053 ();
 sg13g2_decap_8 FILLER_19_2060 ();
 sg13g2_decap_8 FILLER_19_2067 ();
 sg13g2_decap_8 FILLER_19_2074 ();
 sg13g2_decap_4 FILLER_19_2081 ();
 sg13g2_fill_1 FILLER_19_2096 ();
 sg13g2_decap_8 FILLER_19_2114 ();
 sg13g2_decap_8 FILLER_19_2121 ();
 sg13g2_decap_8 FILLER_19_2128 ();
 sg13g2_decap_8 FILLER_19_2135 ();
 sg13g2_decap_4 FILLER_19_2142 ();
 sg13g2_decap_8 FILLER_19_2170 ();
 sg13g2_decap_8 FILLER_19_2177 ();
 sg13g2_decap_8 FILLER_19_2184 ();
 sg13g2_decap_4 FILLER_19_2191 ();
 sg13g2_fill_2 FILLER_19_2195 ();
 sg13g2_fill_2 FILLER_19_2214 ();
 sg13g2_decap_8 FILLER_19_2224 ();
 sg13g2_decap_8 FILLER_19_2231 ();
 sg13g2_decap_8 FILLER_19_2238 ();
 sg13g2_decap_8 FILLER_19_2245 ();
 sg13g2_decap_8 FILLER_19_2252 ();
 sg13g2_fill_2 FILLER_19_2259 ();
 sg13g2_decap_8 FILLER_19_2282 ();
 sg13g2_decap_8 FILLER_19_2289 ();
 sg13g2_decap_8 FILLER_19_2296 ();
 sg13g2_decap_8 FILLER_19_2303 ();
 sg13g2_fill_1 FILLER_19_2310 ();
 sg13g2_decap_8 FILLER_19_2322 ();
 sg13g2_decap_8 FILLER_19_2329 ();
 sg13g2_decap_8 FILLER_19_2346 ();
 sg13g2_decap_8 FILLER_19_2353 ();
 sg13g2_decap_8 FILLER_19_2360 ();
 sg13g2_fill_2 FILLER_19_2367 ();
 sg13g2_fill_1 FILLER_19_2369 ();
 sg13g2_decap_8 FILLER_19_2375 ();
 sg13g2_decap_8 FILLER_19_2382 ();
 sg13g2_fill_2 FILLER_19_2389 ();
 sg13g2_fill_1 FILLER_19_2391 ();
 sg13g2_decap_8 FILLER_19_2403 ();
 sg13g2_decap_8 FILLER_19_2410 ();
 sg13g2_decap_8 FILLER_19_2417 ();
 sg13g2_fill_1 FILLER_19_2424 ();
 sg13g2_decap_8 FILLER_19_2430 ();
 sg13g2_decap_8 FILLER_19_2437 ();
 sg13g2_decap_8 FILLER_19_2444 ();
 sg13g2_decap_8 FILLER_19_2451 ();
 sg13g2_decap_8 FILLER_19_2458 ();
 sg13g2_fill_2 FILLER_19_2465 ();
 sg13g2_fill_1 FILLER_19_2467 ();
 sg13g2_decap_8 FILLER_19_2476 ();
 sg13g2_decap_4 FILLER_19_2486 ();
 sg13g2_fill_1 FILLER_19_2490 ();
 sg13g2_decap_8 FILLER_19_2527 ();
 sg13g2_decap_8 FILLER_19_2534 ();
 sg13g2_decap_8 FILLER_19_2541 ();
 sg13g2_decap_8 FILLER_19_2548 ();
 sg13g2_decap_8 FILLER_19_2555 ();
 sg13g2_decap_8 FILLER_19_2562 ();
 sg13g2_fill_2 FILLER_19_2569 ();
 sg13g2_decap_8 FILLER_19_2574 ();
 sg13g2_decap_8 FILLER_19_2581 ();
 sg13g2_decap_8 FILLER_19_2596 ();
 sg13g2_decap_8 FILLER_19_2603 ();
 sg13g2_fill_2 FILLER_19_2610 ();
 sg13g2_fill_1 FILLER_19_2612 ();
 sg13g2_decap_8 FILLER_19_2639 ();
 sg13g2_decap_8 FILLER_19_2646 ();
 sg13g2_decap_4 FILLER_19_2653 ();
 sg13g2_decap_8 FILLER_19_2683 ();
 sg13g2_decap_4 FILLER_19_2690 ();
 sg13g2_fill_1 FILLER_19_2694 ();
 sg13g2_decap_8 FILLER_19_2742 ();
 sg13g2_decap_8 FILLER_19_2749 ();
 sg13g2_decap_4 FILLER_19_2756 ();
 sg13g2_fill_2 FILLER_19_2760 ();
 sg13g2_decap_8 FILLER_19_2788 ();
 sg13g2_decap_8 FILLER_19_2795 ();
 sg13g2_decap_8 FILLER_19_2802 ();
 sg13g2_decap_8 FILLER_19_2809 ();
 sg13g2_decap_8 FILLER_19_2816 ();
 sg13g2_decap_8 FILLER_19_2823 ();
 sg13g2_decap_8 FILLER_19_2830 ();
 sg13g2_decap_8 FILLER_19_2837 ();
 sg13g2_decap_8 FILLER_19_2844 ();
 sg13g2_decap_8 FILLER_19_2877 ();
 sg13g2_decap_8 FILLER_19_2884 ();
 sg13g2_decap_8 FILLER_19_2891 ();
 sg13g2_decap_8 FILLER_19_2898 ();
 sg13g2_decap_8 FILLER_19_2905 ();
 sg13g2_decap_8 FILLER_19_2912 ();
 sg13g2_decap_8 FILLER_19_2919 ();
 sg13g2_decap_8 FILLER_19_2926 ();
 sg13g2_decap_8 FILLER_19_2933 ();
 sg13g2_decap_8 FILLER_19_2940 ();
 sg13g2_decap_8 FILLER_19_2947 ();
 sg13g2_decap_8 FILLER_19_2954 ();
 sg13g2_decap_8 FILLER_19_2961 ();
 sg13g2_decap_8 FILLER_19_2968 ();
 sg13g2_decap_8 FILLER_19_2975 ();
 sg13g2_decap_8 FILLER_19_2982 ();
 sg13g2_decap_4 FILLER_19_2989 ();
 sg13g2_fill_2 FILLER_19_2993 ();
 sg13g2_decap_8 FILLER_19_3005 ();
 sg13g2_decap_8 FILLER_19_3012 ();
 sg13g2_decap_8 FILLER_19_3061 ();
 sg13g2_decap_8 FILLER_19_3068 ();
 sg13g2_decap_8 FILLER_19_3075 ();
 sg13g2_fill_1 FILLER_19_3082 ();
 sg13g2_fill_1 FILLER_19_3093 ();
 sg13g2_decap_8 FILLER_19_3120 ();
 sg13g2_decap_8 FILLER_19_3127 ();
 sg13g2_decap_8 FILLER_19_3134 ();
 sg13g2_decap_8 FILLER_19_3141 ();
 sg13g2_decap_8 FILLER_19_3148 ();
 sg13g2_decap_8 FILLER_19_3191 ();
 sg13g2_decap_8 FILLER_19_3224 ();
 sg13g2_decap_8 FILLER_19_3231 ();
 sg13g2_decap_8 FILLER_19_3238 ();
 sg13g2_decap_8 FILLER_19_3245 ();
 sg13g2_fill_2 FILLER_19_3252 ();
 sg13g2_fill_1 FILLER_19_3254 ();
 sg13g2_decap_8 FILLER_19_3295 ();
 sg13g2_decap_8 FILLER_19_3302 ();
 sg13g2_decap_8 FILLER_19_3309 ();
 sg13g2_decap_8 FILLER_19_3316 ();
 sg13g2_decap_8 FILLER_19_3323 ();
 sg13g2_decap_4 FILLER_19_3330 ();
 sg13g2_decap_8 FILLER_19_3348 ();
 sg13g2_decap_8 FILLER_19_3355 ();
 sg13g2_decap_8 FILLER_19_3362 ();
 sg13g2_decap_8 FILLER_19_3369 ();
 sg13g2_decap_4 FILLER_19_3376 ();
 sg13g2_fill_2 FILLER_19_3380 ();
 sg13g2_decap_8 FILLER_19_3408 ();
 sg13g2_decap_8 FILLER_19_3415 ();
 sg13g2_decap_4 FILLER_19_3422 ();
 sg13g2_fill_1 FILLER_19_3426 ();
 sg13g2_decap_8 FILLER_19_3462 ();
 sg13g2_fill_2 FILLER_19_3495 ();
 sg13g2_decap_8 FILLER_19_3507 ();
 sg13g2_fill_2 FILLER_19_3514 ();
 sg13g2_decap_8 FILLER_19_3525 ();
 sg13g2_decap_8 FILLER_19_3532 ();
 sg13g2_decap_4 FILLER_19_3552 ();
 sg13g2_decap_8 FILLER_19_3565 ();
 sg13g2_decap_8 FILLER_19_3572 ();
 sg13g2_fill_1 FILLER_19_3579 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_fill_1 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_33 ();
 sg13g2_decap_8 FILLER_20_40 ();
 sg13g2_decap_4 FILLER_20_47 ();
 sg13g2_fill_1 FILLER_20_51 ();
 sg13g2_decap_8 FILLER_20_78 ();
 sg13g2_fill_1 FILLER_20_85 ();
 sg13g2_decap_8 FILLER_20_96 ();
 sg13g2_decap_8 FILLER_20_103 ();
 sg13g2_decap_8 FILLER_20_110 ();
 sg13g2_decap_8 FILLER_20_127 ();
 sg13g2_decap_8 FILLER_20_134 ();
 sg13g2_decap_8 FILLER_20_141 ();
 sg13g2_decap_8 FILLER_20_148 ();
 sg13g2_fill_2 FILLER_20_155 ();
 sg13g2_fill_1 FILLER_20_157 ();
 sg13g2_decap_8 FILLER_20_171 ();
 sg13g2_decap_8 FILLER_20_178 ();
 sg13g2_decap_8 FILLER_20_185 ();
 sg13g2_decap_8 FILLER_20_192 ();
 sg13g2_decap_8 FILLER_20_199 ();
 sg13g2_decap_8 FILLER_20_206 ();
 sg13g2_fill_1 FILLER_20_213 ();
 sg13g2_decap_8 FILLER_20_219 ();
 sg13g2_decap_8 FILLER_20_226 ();
 sg13g2_decap_8 FILLER_20_233 ();
 sg13g2_decap_8 FILLER_20_240 ();
 sg13g2_decap_8 FILLER_20_247 ();
 sg13g2_decap_8 FILLER_20_254 ();
 sg13g2_decap_8 FILLER_20_261 ();
 sg13g2_decap_8 FILLER_20_268 ();
 sg13g2_decap_8 FILLER_20_275 ();
 sg13g2_fill_1 FILLER_20_282 ();
 sg13g2_decap_8 FILLER_20_288 ();
 sg13g2_fill_2 FILLER_20_295 ();
 sg13g2_fill_1 FILLER_20_297 ();
 sg13g2_fill_2 FILLER_20_310 ();
 sg13g2_fill_1 FILLER_20_312 ();
 sg13g2_decap_8 FILLER_20_318 ();
 sg13g2_decap_8 FILLER_20_325 ();
 sg13g2_decap_8 FILLER_20_332 ();
 sg13g2_decap_8 FILLER_20_339 ();
 sg13g2_decap_8 FILLER_20_346 ();
 sg13g2_fill_2 FILLER_20_353 ();
 sg13g2_fill_1 FILLER_20_355 ();
 sg13g2_decap_4 FILLER_20_388 ();
 sg13g2_fill_2 FILLER_20_397 ();
 sg13g2_fill_1 FILLER_20_399 ();
 sg13g2_decap_8 FILLER_20_409 ();
 sg13g2_fill_2 FILLER_20_416 ();
 sg13g2_decap_4 FILLER_20_423 ();
 sg13g2_decap_8 FILLER_20_439 ();
 sg13g2_decap_8 FILLER_20_446 ();
 sg13g2_fill_1 FILLER_20_453 ();
 sg13g2_decap_8 FILLER_20_480 ();
 sg13g2_decap_8 FILLER_20_487 ();
 sg13g2_decap_8 FILLER_20_494 ();
 sg13g2_decap_8 FILLER_20_501 ();
 sg13g2_decap_8 FILLER_20_508 ();
 sg13g2_fill_1 FILLER_20_515 ();
 sg13g2_decap_8 FILLER_20_534 ();
 sg13g2_decap_8 FILLER_20_541 ();
 sg13g2_decap_8 FILLER_20_548 ();
 sg13g2_decap_8 FILLER_20_555 ();
 sg13g2_decap_8 FILLER_20_562 ();
 sg13g2_decap_8 FILLER_20_569 ();
 sg13g2_decap_8 FILLER_20_576 ();
 sg13g2_decap_8 FILLER_20_583 ();
 sg13g2_decap_8 FILLER_20_590 ();
 sg13g2_decap_8 FILLER_20_597 ();
 sg13g2_fill_1 FILLER_20_604 ();
 sg13g2_decap_4 FILLER_20_615 ();
 sg13g2_fill_2 FILLER_20_619 ();
 sg13g2_decap_8 FILLER_20_630 ();
 sg13g2_fill_1 FILLER_20_637 ();
 sg13g2_decap_8 FILLER_20_643 ();
 sg13g2_decap_8 FILLER_20_650 ();
 sg13g2_decap_8 FILLER_20_657 ();
 sg13g2_decap_8 FILLER_20_664 ();
 sg13g2_decap_8 FILLER_20_671 ();
 sg13g2_decap_8 FILLER_20_678 ();
 sg13g2_decap_8 FILLER_20_685 ();
 sg13g2_decap_8 FILLER_20_692 ();
 sg13g2_decap_8 FILLER_20_699 ();
 sg13g2_fill_2 FILLER_20_706 ();
 sg13g2_fill_2 FILLER_20_713 ();
 sg13g2_fill_1 FILLER_20_715 ();
 sg13g2_decap_8 FILLER_20_733 ();
 sg13g2_decap_8 FILLER_20_740 ();
 sg13g2_fill_2 FILLER_20_747 ();
 sg13g2_fill_1 FILLER_20_749 ();
 sg13g2_fill_1 FILLER_20_760 ();
 sg13g2_decap_8 FILLER_20_771 ();
 sg13g2_decap_8 FILLER_20_778 ();
 sg13g2_decap_8 FILLER_20_785 ();
 sg13g2_decap_8 FILLER_20_792 ();
 sg13g2_decap_8 FILLER_20_799 ();
 sg13g2_decap_8 FILLER_20_806 ();
 sg13g2_decap_8 FILLER_20_813 ();
 sg13g2_decap_8 FILLER_20_820 ();
 sg13g2_decap_8 FILLER_20_827 ();
 sg13g2_decap_8 FILLER_20_834 ();
 sg13g2_decap_8 FILLER_20_841 ();
 sg13g2_fill_2 FILLER_20_848 ();
 sg13g2_decap_8 FILLER_20_886 ();
 sg13g2_decap_8 FILLER_20_893 ();
 sg13g2_decap_8 FILLER_20_900 ();
 sg13g2_decap_8 FILLER_20_907 ();
 sg13g2_decap_4 FILLER_20_914 ();
 sg13g2_fill_2 FILLER_20_918 ();
 sg13g2_decap_8 FILLER_20_948 ();
 sg13g2_decap_8 FILLER_20_955 ();
 sg13g2_decap_8 FILLER_20_962 ();
 sg13g2_decap_8 FILLER_20_969 ();
 sg13g2_fill_2 FILLER_20_984 ();
 sg13g2_fill_1 FILLER_20_986 ();
 sg13g2_decap_8 FILLER_20_1000 ();
 sg13g2_decap_8 FILLER_20_1007 ();
 sg13g2_decap_8 FILLER_20_1014 ();
 sg13g2_decap_8 FILLER_20_1021 ();
 sg13g2_decap_8 FILLER_20_1028 ();
 sg13g2_decap_8 FILLER_20_1035 ();
 sg13g2_decap_8 FILLER_20_1042 ();
 sg13g2_decap_8 FILLER_20_1049 ();
 sg13g2_decap_8 FILLER_20_1056 ();
 sg13g2_fill_2 FILLER_20_1063 ();
 sg13g2_decap_8 FILLER_20_1078 ();
 sg13g2_decap_8 FILLER_20_1085 ();
 sg13g2_decap_8 FILLER_20_1092 ();
 sg13g2_decap_4 FILLER_20_1099 ();
 sg13g2_fill_1 FILLER_20_1103 ();
 sg13g2_decap_8 FILLER_20_1138 ();
 sg13g2_decap_8 FILLER_20_1145 ();
 sg13g2_decap_8 FILLER_20_1152 ();
 sg13g2_decap_8 FILLER_20_1159 ();
 sg13g2_decap_8 FILLER_20_1166 ();
 sg13g2_decap_8 FILLER_20_1173 ();
 sg13g2_decap_8 FILLER_20_1180 ();
 sg13g2_decap_8 FILLER_20_1187 ();
 sg13g2_decap_4 FILLER_20_1194 ();
 sg13g2_decap_4 FILLER_20_1206 ();
 sg13g2_fill_2 FILLER_20_1210 ();
 sg13g2_decap_8 FILLER_20_1238 ();
 sg13g2_fill_2 FILLER_20_1245 ();
 sg13g2_decap_8 FILLER_20_1277 ();
 sg13g2_fill_2 FILLER_20_1284 ();
 sg13g2_fill_1 FILLER_20_1286 ();
 sg13g2_fill_2 FILLER_20_1313 ();
 sg13g2_decap_8 FILLER_20_1323 ();
 sg13g2_fill_2 FILLER_20_1330 ();
 sg13g2_decap_8 FILLER_20_1369 ();
 sg13g2_decap_8 FILLER_20_1376 ();
 sg13g2_decap_8 FILLER_20_1383 ();
 sg13g2_decap_8 FILLER_20_1390 ();
 sg13g2_decap_8 FILLER_20_1397 ();
 sg13g2_decap_8 FILLER_20_1404 ();
 sg13g2_decap_8 FILLER_20_1411 ();
 sg13g2_decap_8 FILLER_20_1418 ();
 sg13g2_decap_4 FILLER_20_1425 ();
 sg13g2_fill_1 FILLER_20_1429 ();
 sg13g2_decap_8 FILLER_20_1441 ();
 sg13g2_decap_4 FILLER_20_1448 ();
 sg13g2_fill_1 FILLER_20_1452 ();
 sg13g2_decap_8 FILLER_20_1459 ();
 sg13g2_decap_8 FILLER_20_1466 ();
 sg13g2_decap_8 FILLER_20_1473 ();
 sg13g2_decap_4 FILLER_20_1480 ();
 sg13g2_fill_1 FILLER_20_1484 ();
 sg13g2_decap_8 FILLER_20_1490 ();
 sg13g2_decap_8 FILLER_20_1497 ();
 sg13g2_fill_2 FILLER_20_1504 ();
 sg13g2_fill_1 FILLER_20_1506 ();
 sg13g2_decap_8 FILLER_20_1533 ();
 sg13g2_decap_8 FILLER_20_1540 ();
 sg13g2_decap_8 FILLER_20_1547 ();
 sg13g2_decap_4 FILLER_20_1554 ();
 sg13g2_decap_8 FILLER_20_1610 ();
 sg13g2_decap_8 FILLER_20_1617 ();
 sg13g2_decap_8 FILLER_20_1624 ();
 sg13g2_decap_8 FILLER_20_1631 ();
 sg13g2_decap_8 FILLER_20_1638 ();
 sg13g2_decap_8 FILLER_20_1645 ();
 sg13g2_decap_8 FILLER_20_1652 ();
 sg13g2_decap_8 FILLER_20_1680 ();
 sg13g2_decap_8 FILLER_20_1687 ();
 sg13g2_decap_4 FILLER_20_1694 ();
 sg13g2_decap_4 FILLER_20_1709 ();
 sg13g2_fill_2 FILLER_20_1713 ();
 sg13g2_decap_8 FILLER_20_1721 ();
 sg13g2_decap_8 FILLER_20_1728 ();
 sg13g2_fill_1 FILLER_20_1735 ();
 sg13g2_fill_2 FILLER_20_1773 ();
 sg13g2_fill_1 FILLER_20_1775 ();
 sg13g2_decap_8 FILLER_20_1786 ();
 sg13g2_decap_8 FILLER_20_1793 ();
 sg13g2_decap_8 FILLER_20_1800 ();
 sg13g2_decap_8 FILLER_20_1807 ();
 sg13g2_decap_8 FILLER_20_1814 ();
 sg13g2_fill_1 FILLER_20_1821 ();
 sg13g2_decap_8 FILLER_20_1848 ();
 sg13g2_decap_8 FILLER_20_1855 ();
 sg13g2_decap_8 FILLER_20_1862 ();
 sg13g2_decap_8 FILLER_20_1869 ();
 sg13g2_fill_2 FILLER_20_1876 ();
 sg13g2_decap_8 FILLER_20_1904 ();
 sg13g2_decap_8 FILLER_20_1911 ();
 sg13g2_decap_8 FILLER_20_1918 ();
 sg13g2_decap_8 FILLER_20_1925 ();
 sg13g2_decap_4 FILLER_20_1932 ();
 sg13g2_fill_2 FILLER_20_1952 ();
 sg13g2_decap_8 FILLER_20_1962 ();
 sg13g2_decap_8 FILLER_20_1969 ();
 sg13g2_decap_8 FILLER_20_1976 ();
 sg13g2_fill_2 FILLER_20_1983 ();
 sg13g2_fill_1 FILLER_20_1985 ();
 sg13g2_decap_4 FILLER_20_2016 ();
 sg13g2_decap_8 FILLER_20_2056 ();
 sg13g2_decap_8 FILLER_20_2063 ();
 sg13g2_decap_8 FILLER_20_2070 ();
 sg13g2_fill_2 FILLER_20_2077 ();
 sg13g2_decap_8 FILLER_20_2082 ();
 sg13g2_decap_8 FILLER_20_2089 ();
 sg13g2_decap_8 FILLER_20_2122 ();
 sg13g2_decap_8 FILLER_20_2129 ();
 sg13g2_decap_8 FILLER_20_2136 ();
 sg13g2_decap_8 FILLER_20_2143 ();
 sg13g2_decap_4 FILLER_20_2150 ();
 sg13g2_decap_4 FILLER_20_2180 ();
 sg13g2_fill_2 FILLER_20_2184 ();
 sg13g2_decap_8 FILLER_20_2198 ();
 sg13g2_decap_8 FILLER_20_2208 ();
 sg13g2_decap_8 FILLER_20_2215 ();
 sg13g2_decap_8 FILLER_20_2222 ();
 sg13g2_decap_8 FILLER_20_2229 ();
 sg13g2_decap_8 FILLER_20_2236 ();
 sg13g2_decap_8 FILLER_20_2243 ();
 sg13g2_decap_8 FILLER_20_2250 ();
 sg13g2_decap_8 FILLER_20_2257 ();
 sg13g2_decap_4 FILLER_20_2264 ();
 sg13g2_fill_1 FILLER_20_2268 ();
 sg13g2_decap_4 FILLER_20_2275 ();
 sg13g2_decap_8 FILLER_20_2305 ();
 sg13g2_decap_8 FILLER_20_2312 ();
 sg13g2_decap_8 FILLER_20_2319 ();
 sg13g2_decap_8 FILLER_20_2326 ();
 sg13g2_decap_8 FILLER_20_2333 ();
 sg13g2_decap_8 FILLER_20_2346 ();
 sg13g2_decap_8 FILLER_20_2353 ();
 sg13g2_decap_8 FILLER_20_2360 ();
 sg13g2_decap_8 FILLER_20_2367 ();
 sg13g2_fill_1 FILLER_20_2374 ();
 sg13g2_decap_8 FILLER_20_2385 ();
 sg13g2_decap_8 FILLER_20_2392 ();
 sg13g2_decap_8 FILLER_20_2399 ();
 sg13g2_decap_8 FILLER_20_2406 ();
 sg13g2_decap_8 FILLER_20_2413 ();
 sg13g2_fill_2 FILLER_20_2420 ();
 sg13g2_decap_8 FILLER_20_2453 ();
 sg13g2_decap_8 FILLER_20_2460 ();
 sg13g2_decap_8 FILLER_20_2467 ();
 sg13g2_decap_8 FILLER_20_2474 ();
 sg13g2_decap_8 FILLER_20_2481 ();
 sg13g2_decap_8 FILLER_20_2488 ();
 sg13g2_decap_8 FILLER_20_2500 ();
 sg13g2_decap_8 FILLER_20_2507 ();
 sg13g2_decap_8 FILLER_20_2514 ();
 sg13g2_decap_8 FILLER_20_2521 ();
 sg13g2_decap_8 FILLER_20_2528 ();
 sg13g2_decap_8 FILLER_20_2535 ();
 sg13g2_decap_8 FILLER_20_2542 ();
 sg13g2_decap_8 FILLER_20_2549 ();
 sg13g2_decap_8 FILLER_20_2556 ();
 sg13g2_decap_8 FILLER_20_2563 ();
 sg13g2_decap_8 FILLER_20_2570 ();
 sg13g2_decap_8 FILLER_20_2577 ();
 sg13g2_fill_2 FILLER_20_2584 ();
 sg13g2_fill_1 FILLER_20_2586 ();
 sg13g2_decap_8 FILLER_20_2601 ();
 sg13g2_decap_8 FILLER_20_2608 ();
 sg13g2_decap_8 FILLER_20_2615 ();
 sg13g2_decap_8 FILLER_20_2622 ();
 sg13g2_decap_8 FILLER_20_2629 ();
 sg13g2_decap_8 FILLER_20_2636 ();
 sg13g2_decap_8 FILLER_20_2643 ();
 sg13g2_decap_8 FILLER_20_2650 ();
 sg13g2_decap_4 FILLER_20_2657 ();
 sg13g2_fill_1 FILLER_20_2661 ();
 sg13g2_decap_4 FILLER_20_2672 ();
 sg13g2_decap_8 FILLER_20_2681 ();
 sg13g2_decap_8 FILLER_20_2688 ();
 sg13g2_decap_8 FILLER_20_2695 ();
 sg13g2_decap_8 FILLER_20_2702 ();
 sg13g2_decap_8 FILLER_20_2709 ();
 sg13g2_decap_8 FILLER_20_2716 ();
 sg13g2_decap_8 FILLER_20_2723 ();
 sg13g2_decap_8 FILLER_20_2730 ();
 sg13g2_decap_8 FILLER_20_2737 ();
 sg13g2_decap_8 FILLER_20_2744 ();
 sg13g2_decap_8 FILLER_20_2751 ();
 sg13g2_decap_8 FILLER_20_2794 ();
 sg13g2_decap_8 FILLER_20_2801 ();
 sg13g2_fill_2 FILLER_20_2808 ();
 sg13g2_fill_1 FILLER_20_2810 ();
 sg13g2_decap_4 FILLER_20_2819 ();
 sg13g2_fill_1 FILLER_20_2823 ();
 sg13g2_decap_4 FILLER_20_2836 ();
 sg13g2_fill_2 FILLER_20_2840 ();
 sg13g2_decap_4 FILLER_20_2852 ();
 sg13g2_fill_1 FILLER_20_2856 ();
 sg13g2_decap_4 FILLER_20_2867 ();
 sg13g2_fill_2 FILLER_20_2871 ();
 sg13g2_decap_8 FILLER_20_2912 ();
 sg13g2_fill_1 FILLER_20_2919 ();
 sg13g2_decap_8 FILLER_20_2925 ();
 sg13g2_decap_8 FILLER_20_2932 ();
 sg13g2_fill_2 FILLER_20_2939 ();
 sg13g2_decap_8 FILLER_20_2967 ();
 sg13g2_decap_4 FILLER_20_2974 ();
 sg13g2_fill_1 FILLER_20_2978 ();
 sg13g2_decap_8 FILLER_20_3005 ();
 sg13g2_decap_8 FILLER_20_3012 ();
 sg13g2_decap_4 FILLER_20_3019 ();
 sg13g2_decap_8 FILLER_20_3068 ();
 sg13g2_decap_4 FILLER_20_3075 ();
 sg13g2_decap_8 FILLER_20_3089 ();
 sg13g2_decap_8 FILLER_20_3096 ();
 sg13g2_decap_8 FILLER_20_3103 ();
 sg13g2_decap_8 FILLER_20_3110 ();
 sg13g2_decap_8 FILLER_20_3117 ();
 sg13g2_decap_8 FILLER_20_3124 ();
 sg13g2_decap_8 FILLER_20_3131 ();
 sg13g2_decap_8 FILLER_20_3138 ();
 sg13g2_decap_8 FILLER_20_3145 ();
 sg13g2_fill_2 FILLER_20_3152 ();
 sg13g2_fill_1 FILLER_20_3154 ();
 sg13g2_decap_8 FILLER_20_3181 ();
 sg13g2_decap_8 FILLER_20_3188 ();
 sg13g2_decap_8 FILLER_20_3195 ();
 sg13g2_decap_4 FILLER_20_3202 ();
 sg13g2_decap_8 FILLER_20_3216 ();
 sg13g2_decap_8 FILLER_20_3223 ();
 sg13g2_decap_4 FILLER_20_3230 ();
 sg13g2_decap_8 FILLER_20_3239 ();
 sg13g2_decap_8 FILLER_20_3246 ();
 sg13g2_decap_8 FILLER_20_3253 ();
 sg13g2_decap_8 FILLER_20_3260 ();
 sg13g2_decap_4 FILLER_20_3267 ();
 sg13g2_fill_2 FILLER_20_3271 ();
 sg13g2_decap_8 FILLER_20_3292 ();
 sg13g2_decap_8 FILLER_20_3299 ();
 sg13g2_decap_8 FILLER_20_3306 ();
 sg13g2_decap_8 FILLER_20_3313 ();
 sg13g2_decap_4 FILLER_20_3320 ();
 sg13g2_fill_2 FILLER_20_3324 ();
 sg13g2_decap_8 FILLER_20_3362 ();
 sg13g2_fill_2 FILLER_20_3369 ();
 sg13g2_fill_1 FILLER_20_3371 ();
 sg13g2_decap_8 FILLER_20_3400 ();
 sg13g2_decap_8 FILLER_20_3407 ();
 sg13g2_decap_8 FILLER_20_3414 ();
 sg13g2_decap_8 FILLER_20_3421 ();
 sg13g2_fill_1 FILLER_20_3428 ();
 sg13g2_decap_8 FILLER_20_3452 ();
 sg13g2_decap_8 FILLER_20_3459 ();
 sg13g2_decap_8 FILLER_20_3466 ();
 sg13g2_decap_4 FILLER_20_3473 ();
 sg13g2_fill_2 FILLER_20_3477 ();
 sg13g2_fill_2 FILLER_20_3505 ();
 sg13g2_fill_2 FILLER_20_3533 ();
 sg13g2_fill_1 FILLER_20_3535 ();
 sg13g2_decap_8 FILLER_20_3572 ();
 sg13g2_fill_1 FILLER_20_3579 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_4 FILLER_21_7 ();
 sg13g2_fill_1 FILLER_21_11 ();
 sg13g2_decap_8 FILLER_21_58 ();
 sg13g2_decap_8 FILLER_21_74 ();
 sg13g2_decap_4 FILLER_21_81 ();
 sg13g2_decap_4 FILLER_21_111 ();
 sg13g2_fill_2 FILLER_21_115 ();
 sg13g2_fill_1 FILLER_21_123 ();
 sg13g2_decap_8 FILLER_21_132 ();
 sg13g2_decap_8 FILLER_21_139 ();
 sg13g2_decap_4 FILLER_21_146 ();
 sg13g2_fill_2 FILLER_21_150 ();
 sg13g2_decap_8 FILLER_21_174 ();
 sg13g2_decap_4 FILLER_21_181 ();
 sg13g2_decap_8 FILLER_21_190 ();
 sg13g2_decap_8 FILLER_21_197 ();
 sg13g2_decap_4 FILLER_21_204 ();
 sg13g2_decap_4 FILLER_21_215 ();
 sg13g2_fill_2 FILLER_21_235 ();
 sg13g2_fill_1 FILLER_21_237 ();
 sg13g2_decap_8 FILLER_21_246 ();
 sg13g2_decap_8 FILLER_21_253 ();
 sg13g2_decap_8 FILLER_21_260 ();
 sg13g2_decap_8 FILLER_21_267 ();
 sg13g2_decap_8 FILLER_21_274 ();
 sg13g2_decap_8 FILLER_21_281 ();
 sg13g2_decap_8 FILLER_21_288 ();
 sg13g2_decap_8 FILLER_21_295 ();
 sg13g2_fill_2 FILLER_21_302 ();
 sg13g2_fill_1 FILLER_21_304 ();
 sg13g2_decap_8 FILLER_21_310 ();
 sg13g2_decap_8 FILLER_21_317 ();
 sg13g2_decap_8 FILLER_21_324 ();
 sg13g2_decap_8 FILLER_21_331 ();
 sg13g2_decap_8 FILLER_21_338 ();
 sg13g2_decap_4 FILLER_21_345 ();
 sg13g2_fill_2 FILLER_21_359 ();
 sg13g2_decap_4 FILLER_21_366 ();
 sg13g2_fill_1 FILLER_21_370 ();
 sg13g2_fill_2 FILLER_21_374 ();
 sg13g2_fill_1 FILLER_21_376 ();
 sg13g2_decap_8 FILLER_21_392 ();
 sg13g2_decap_4 FILLER_21_399 ();
 sg13g2_decap_8 FILLER_21_409 ();
 sg13g2_decap_4 FILLER_21_416 ();
 sg13g2_fill_1 FILLER_21_420 ();
 sg13g2_decap_8 FILLER_21_431 ();
 sg13g2_decap_8 FILLER_21_438 ();
 sg13g2_decap_4 FILLER_21_445 ();
 sg13g2_fill_1 FILLER_21_449 ();
 sg13g2_decap_8 FILLER_21_473 ();
 sg13g2_decap_8 FILLER_21_480 ();
 sg13g2_decap_8 FILLER_21_487 ();
 sg13g2_decap_8 FILLER_21_494 ();
 sg13g2_decap_8 FILLER_21_501 ();
 sg13g2_decap_4 FILLER_21_508 ();
 sg13g2_fill_1 FILLER_21_528 ();
 sg13g2_decap_8 FILLER_21_544 ();
 sg13g2_decap_8 FILLER_21_551 ();
 sg13g2_decap_8 FILLER_21_558 ();
 sg13g2_decap_8 FILLER_21_565 ();
 sg13g2_decap_8 FILLER_21_572 ();
 sg13g2_fill_2 FILLER_21_605 ();
 sg13g2_decap_8 FILLER_21_633 ();
 sg13g2_decap_8 FILLER_21_640 ();
 sg13g2_decap_8 FILLER_21_647 ();
 sg13g2_decap_8 FILLER_21_654 ();
 sg13g2_decap_4 FILLER_21_661 ();
 sg13g2_fill_1 FILLER_21_665 ();
 sg13g2_decap_8 FILLER_21_674 ();
 sg13g2_decap_4 FILLER_21_681 ();
 sg13g2_fill_1 FILLER_21_685 ();
 sg13g2_decap_8 FILLER_21_694 ();
 sg13g2_fill_2 FILLER_21_708 ();
 sg13g2_decap_8 FILLER_21_726 ();
 sg13g2_decap_8 FILLER_21_733 ();
 sg13g2_decap_8 FILLER_21_740 ();
 sg13g2_fill_2 FILLER_21_747 ();
 sg13g2_decap_8 FILLER_21_775 ();
 sg13g2_decap_8 FILLER_21_782 ();
 sg13g2_decap_8 FILLER_21_815 ();
 sg13g2_decap_8 FILLER_21_822 ();
 sg13g2_decap_8 FILLER_21_829 ();
 sg13g2_decap_8 FILLER_21_836 ();
 sg13g2_decap_8 FILLER_21_843 ();
 sg13g2_decap_8 FILLER_21_850 ();
 sg13g2_fill_2 FILLER_21_857 ();
 sg13g2_fill_1 FILLER_21_859 ();
 sg13g2_decap_8 FILLER_21_868 ();
 sg13g2_decap_8 FILLER_21_875 ();
 sg13g2_decap_8 FILLER_21_882 ();
 sg13g2_decap_8 FILLER_21_889 ();
 sg13g2_decap_8 FILLER_21_896 ();
 sg13g2_decap_8 FILLER_21_903 ();
 sg13g2_decap_8 FILLER_21_910 ();
 sg13g2_decap_8 FILLER_21_917 ();
 sg13g2_fill_1 FILLER_21_924 ();
 sg13g2_decap_8 FILLER_21_929 ();
 sg13g2_decap_8 FILLER_21_936 ();
 sg13g2_decap_8 FILLER_21_943 ();
 sg13g2_decap_8 FILLER_21_950 ();
 sg13g2_decap_8 FILLER_21_957 ();
 sg13g2_decap_8 FILLER_21_964 ();
 sg13g2_decap_8 FILLER_21_971 ();
 sg13g2_decap_8 FILLER_21_978 ();
 sg13g2_decap_8 FILLER_21_985 ();
 sg13g2_decap_8 FILLER_21_992 ();
 sg13g2_decap_8 FILLER_21_999 ();
 sg13g2_decap_8 FILLER_21_1006 ();
 sg13g2_decap_8 FILLER_21_1019 ();
 sg13g2_decap_8 FILLER_21_1026 ();
 sg13g2_decap_8 FILLER_21_1033 ();
 sg13g2_fill_2 FILLER_21_1040 ();
 sg13g2_decap_4 FILLER_21_1045 ();
 sg13g2_fill_1 FILLER_21_1049 ();
 sg13g2_decap_8 FILLER_21_1069 ();
 sg13g2_decap_8 FILLER_21_1076 ();
 sg13g2_decap_8 FILLER_21_1083 ();
 sg13g2_decap_8 FILLER_21_1090 ();
 sg13g2_decap_4 FILLER_21_1097 ();
 sg13g2_decap_8 FILLER_21_1140 ();
 sg13g2_decap_8 FILLER_21_1147 ();
 sg13g2_decap_8 FILLER_21_1154 ();
 sg13g2_decap_4 FILLER_21_1161 ();
 sg13g2_fill_1 FILLER_21_1191 ();
 sg13g2_decap_8 FILLER_21_1197 ();
 sg13g2_decap_8 FILLER_21_1204 ();
 sg13g2_decap_4 FILLER_21_1211 ();
 sg13g2_decap_4 FILLER_21_1223 ();
 sg13g2_decap_8 FILLER_21_1235 ();
 sg13g2_decap_8 FILLER_21_1242 ();
 sg13g2_decap_4 FILLER_21_1249 ();
 sg13g2_fill_1 FILLER_21_1253 ();
 sg13g2_decap_8 FILLER_21_1291 ();
 sg13g2_decap_8 FILLER_21_1298 ();
 sg13g2_decap_8 FILLER_21_1305 ();
 sg13g2_decap_8 FILLER_21_1312 ();
 sg13g2_decap_8 FILLER_21_1319 ();
 sg13g2_decap_8 FILLER_21_1326 ();
 sg13g2_decap_8 FILLER_21_1333 ();
 sg13g2_decap_8 FILLER_21_1340 ();
 sg13g2_decap_8 FILLER_21_1347 ();
 sg13g2_decap_8 FILLER_21_1354 ();
 sg13g2_decap_8 FILLER_21_1361 ();
 sg13g2_fill_2 FILLER_21_1368 ();
 sg13g2_fill_1 FILLER_21_1370 ();
 sg13g2_decap_8 FILLER_21_1381 ();
 sg13g2_fill_1 FILLER_21_1388 ();
 sg13g2_fill_2 FILLER_21_1420 ();
 sg13g2_fill_1 FILLER_21_1422 ();
 sg13g2_fill_1 FILLER_21_1433 ();
 sg13g2_decap_8 FILLER_21_1442 ();
 sg13g2_decap_4 FILLER_21_1449 ();
 sg13g2_decap_8 FILLER_21_1462 ();
 sg13g2_decap_8 FILLER_21_1469 ();
 sg13g2_decap_8 FILLER_21_1476 ();
 sg13g2_decap_8 FILLER_21_1483 ();
 sg13g2_decap_8 FILLER_21_1490 ();
 sg13g2_decap_8 FILLER_21_1497 ();
 sg13g2_decap_4 FILLER_21_1504 ();
 sg13g2_fill_2 FILLER_21_1508 ();
 sg13g2_decap_8 FILLER_21_1515 ();
 sg13g2_decap_8 FILLER_21_1522 ();
 sg13g2_decap_8 FILLER_21_1529 ();
 sg13g2_decap_8 FILLER_21_1536 ();
 sg13g2_decap_8 FILLER_21_1546 ();
 sg13g2_decap_4 FILLER_21_1553 ();
 sg13g2_decap_8 FILLER_21_1567 ();
 sg13g2_decap_8 FILLER_21_1574 ();
 sg13g2_decap_8 FILLER_21_1581 ();
 sg13g2_decap_8 FILLER_21_1588 ();
 sg13g2_decap_8 FILLER_21_1595 ();
 sg13g2_decap_8 FILLER_21_1628 ();
 sg13g2_decap_8 FILLER_21_1635 ();
 sg13g2_decap_8 FILLER_21_1642 ();
 sg13g2_decap_8 FILLER_21_1649 ();
 sg13g2_decap_8 FILLER_21_1656 ();
 sg13g2_decap_8 FILLER_21_1663 ();
 sg13g2_decap_8 FILLER_21_1670 ();
 sg13g2_decap_8 FILLER_21_1677 ();
 sg13g2_decap_8 FILLER_21_1684 ();
 sg13g2_decap_8 FILLER_21_1691 ();
 sg13g2_decap_8 FILLER_21_1698 ();
 sg13g2_decap_8 FILLER_21_1705 ();
 sg13g2_fill_2 FILLER_21_1712 ();
 sg13g2_fill_1 FILLER_21_1714 ();
 sg13g2_decap_8 FILLER_21_1726 ();
 sg13g2_decap_8 FILLER_21_1753 ();
 sg13g2_decap_4 FILLER_21_1760 ();
 sg13g2_fill_2 FILLER_21_1764 ();
 sg13g2_decap_8 FILLER_21_1772 ();
 sg13g2_decap_8 FILLER_21_1779 ();
 sg13g2_decap_8 FILLER_21_1786 ();
 sg13g2_decap_8 FILLER_21_1793 ();
 sg13g2_decap_8 FILLER_21_1800 ();
 sg13g2_fill_2 FILLER_21_1807 ();
 sg13g2_fill_1 FILLER_21_1809 ();
 sg13g2_decap_8 FILLER_21_1846 ();
 sg13g2_decap_8 FILLER_21_1853 ();
 sg13g2_decap_8 FILLER_21_1860 ();
 sg13g2_fill_2 FILLER_21_1873 ();
 sg13g2_decap_8 FILLER_21_1885 ();
 sg13g2_fill_2 FILLER_21_1912 ();
 sg13g2_decap_8 FILLER_21_1925 ();
 sg13g2_decap_4 FILLER_21_1932 ();
 sg13g2_fill_2 FILLER_21_1936 ();
 sg13g2_decap_8 FILLER_21_1946 ();
 sg13g2_decap_4 FILLER_21_1953 ();
 sg13g2_decap_8 FILLER_21_1965 ();
 sg13g2_decap_8 FILLER_21_1972 ();
 sg13g2_decap_4 FILLER_21_1979 ();
 sg13g2_fill_1 FILLER_21_1983 ();
 sg13g2_decap_8 FILLER_21_2021 ();
 sg13g2_decap_8 FILLER_21_2028 ();
 sg13g2_decap_8 FILLER_21_2035 ();
 sg13g2_decap_8 FILLER_21_2042 ();
 sg13g2_decap_8 FILLER_21_2049 ();
 sg13g2_decap_4 FILLER_21_2056 ();
 sg13g2_fill_2 FILLER_21_2060 ();
 sg13g2_decap_8 FILLER_21_2068 ();
 sg13g2_decap_8 FILLER_21_2075 ();
 sg13g2_decap_8 FILLER_21_2082 ();
 sg13g2_decap_8 FILLER_21_2089 ();
 sg13g2_decap_8 FILLER_21_2096 ();
 sg13g2_decap_8 FILLER_21_2103 ();
 sg13g2_fill_2 FILLER_21_2110 ();
 sg13g2_decap_8 FILLER_21_2138 ();
 sg13g2_decap_8 FILLER_21_2145 ();
 sg13g2_decap_8 FILLER_21_2152 ();
 sg13g2_decap_8 FILLER_21_2159 ();
 sg13g2_decap_8 FILLER_21_2166 ();
 sg13g2_decap_8 FILLER_21_2173 ();
 sg13g2_fill_1 FILLER_21_2180 ();
 sg13g2_decap_8 FILLER_21_2187 ();
 sg13g2_decap_4 FILLER_21_2194 ();
 sg13g2_fill_2 FILLER_21_2198 ();
 sg13g2_fill_1 FILLER_21_2204 ();
 sg13g2_decap_8 FILLER_21_2241 ();
 sg13g2_decap_8 FILLER_21_2248 ();
 sg13g2_fill_2 FILLER_21_2255 ();
 sg13g2_fill_1 FILLER_21_2269 ();
 sg13g2_decap_8 FILLER_21_2291 ();
 sg13g2_decap_8 FILLER_21_2298 ();
 sg13g2_decap_8 FILLER_21_2305 ();
 sg13g2_decap_8 FILLER_21_2312 ();
 sg13g2_fill_2 FILLER_21_2319 ();
 sg13g2_fill_1 FILLER_21_2321 ();
 sg13g2_decap_4 FILLER_21_2337 ();
 sg13g2_fill_2 FILLER_21_2341 ();
 sg13g2_decap_8 FILLER_21_2355 ();
 sg13g2_fill_2 FILLER_21_2362 ();
 sg13g2_fill_1 FILLER_21_2369 ();
 sg13g2_decap_8 FILLER_21_2396 ();
 sg13g2_decap_8 FILLER_21_2403 ();
 sg13g2_decap_8 FILLER_21_2410 ();
 sg13g2_decap_8 FILLER_21_2417 ();
 sg13g2_decap_8 FILLER_21_2424 ();
 sg13g2_fill_2 FILLER_21_2431 ();
 sg13g2_decap_4 FILLER_21_2436 ();
 sg13g2_decap_8 FILLER_21_2449 ();
 sg13g2_decap_4 FILLER_21_2456 ();
 sg13g2_decap_8 FILLER_21_2468 ();
 sg13g2_decap_8 FILLER_21_2475 ();
 sg13g2_decap_8 FILLER_21_2482 ();
 sg13g2_decap_8 FILLER_21_2510 ();
 sg13g2_decap_8 FILLER_21_2517 ();
 sg13g2_decap_8 FILLER_21_2524 ();
 sg13g2_fill_1 FILLER_21_2531 ();
 sg13g2_decap_8 FILLER_21_2542 ();
 sg13g2_decap_8 FILLER_21_2565 ();
 sg13g2_decap_4 FILLER_21_2572 ();
 sg13g2_fill_1 FILLER_21_2576 ();
 sg13g2_decap_8 FILLER_21_2583 ();
 sg13g2_decap_8 FILLER_21_2590 ();
 sg13g2_decap_8 FILLER_21_2597 ();
 sg13g2_fill_2 FILLER_21_2604 ();
 sg13g2_decap_8 FILLER_21_2616 ();
 sg13g2_decap_8 FILLER_21_2623 ();
 sg13g2_fill_1 FILLER_21_2630 ();
 sg13g2_decap_8 FILLER_21_2637 ();
 sg13g2_decap_8 FILLER_21_2644 ();
 sg13g2_decap_8 FILLER_21_2651 ();
 sg13g2_decap_8 FILLER_21_2658 ();
 sg13g2_decap_8 FILLER_21_2665 ();
 sg13g2_fill_2 FILLER_21_2672 ();
 sg13g2_fill_1 FILLER_21_2674 ();
 sg13g2_decap_8 FILLER_21_2680 ();
 sg13g2_decap_8 FILLER_21_2687 ();
 sg13g2_decap_8 FILLER_21_2694 ();
 sg13g2_decap_8 FILLER_21_2701 ();
 sg13g2_decap_8 FILLER_21_2708 ();
 sg13g2_decap_8 FILLER_21_2715 ();
 sg13g2_decap_8 FILLER_21_2722 ();
 sg13g2_decap_8 FILLER_21_2729 ();
 sg13g2_decap_8 FILLER_21_2736 ();
 sg13g2_decap_8 FILLER_21_2743 ();
 sg13g2_decap_8 FILLER_21_2750 ();
 sg13g2_decap_8 FILLER_21_2757 ();
 sg13g2_decap_4 FILLER_21_2764 ();
 sg13g2_decap_8 FILLER_21_2804 ();
 sg13g2_decap_8 FILLER_21_2811 ();
 sg13g2_decap_8 FILLER_21_2818 ();
 sg13g2_decap_8 FILLER_21_2825 ();
 sg13g2_decap_8 FILLER_21_2832 ();
 sg13g2_decap_8 FILLER_21_2839 ();
 sg13g2_decap_8 FILLER_21_2861 ();
 sg13g2_decap_8 FILLER_21_2868 ();
 sg13g2_decap_8 FILLER_21_2875 ();
 sg13g2_decap_8 FILLER_21_2882 ();
 sg13g2_decap_8 FILLER_21_2889 ();
 sg13g2_decap_4 FILLER_21_2896 ();
 sg13g2_fill_1 FILLER_21_2900 ();
 sg13g2_decap_8 FILLER_21_2909 ();
 sg13g2_fill_2 FILLER_21_2916 ();
 sg13g2_fill_1 FILLER_21_2918 ();
 sg13g2_decap_8 FILLER_21_2927 ();
 sg13g2_decap_4 FILLER_21_2934 ();
 sg13g2_fill_2 FILLER_21_2938 ();
 sg13g2_fill_2 FILLER_21_2966 ();
 sg13g2_fill_1 FILLER_21_2968 ();
 sg13g2_decap_8 FILLER_21_2979 ();
 sg13g2_decap_8 FILLER_21_2986 ();
 sg13g2_decap_8 FILLER_21_2993 ();
 sg13g2_decap_8 FILLER_21_3000 ();
 sg13g2_decap_8 FILLER_21_3007 ();
 sg13g2_decap_8 FILLER_21_3014 ();
 sg13g2_decap_8 FILLER_21_3021 ();
 sg13g2_decap_4 FILLER_21_3028 ();
 sg13g2_decap_8 FILLER_21_3041 ();
 sg13g2_decap_8 FILLER_21_3048 ();
 sg13g2_decap_8 FILLER_21_3055 ();
 sg13g2_decap_8 FILLER_21_3062 ();
 sg13g2_fill_2 FILLER_21_3069 ();
 sg13g2_decap_8 FILLER_21_3097 ();
 sg13g2_decap_8 FILLER_21_3104 ();
 sg13g2_decap_8 FILLER_21_3111 ();
 sg13g2_decap_8 FILLER_21_3118 ();
 sg13g2_decap_8 FILLER_21_3125 ();
 sg13g2_decap_8 FILLER_21_3132 ();
 sg13g2_fill_1 FILLER_21_3139 ();
 sg13g2_decap_8 FILLER_21_3150 ();
 sg13g2_decap_8 FILLER_21_3157 ();
 sg13g2_decap_8 FILLER_21_3164 ();
 sg13g2_decap_8 FILLER_21_3171 ();
 sg13g2_decap_8 FILLER_21_3178 ();
 sg13g2_decap_8 FILLER_21_3185 ();
 sg13g2_decap_8 FILLER_21_3192 ();
 sg13g2_decap_8 FILLER_21_3251 ();
 sg13g2_decap_8 FILLER_21_3258 ();
 sg13g2_fill_2 FILLER_21_3265 ();
 sg13g2_decap_8 FILLER_21_3303 ();
 sg13g2_decap_8 FILLER_21_3310 ();
 sg13g2_decap_4 FILLER_21_3317 ();
 sg13g2_fill_1 FILLER_21_3321 ();
 sg13g2_decap_8 FILLER_21_3348 ();
 sg13g2_decap_8 FILLER_21_3355 ();
 sg13g2_decap_8 FILLER_21_3362 ();
 sg13g2_decap_8 FILLER_21_3369 ();
 sg13g2_decap_8 FILLER_21_3376 ();
 sg13g2_decap_8 FILLER_21_3383 ();
 sg13g2_decap_8 FILLER_21_3390 ();
 sg13g2_decap_8 FILLER_21_3397 ();
 sg13g2_decap_8 FILLER_21_3404 ();
 sg13g2_decap_8 FILLER_21_3411 ();
 sg13g2_decap_8 FILLER_21_3418 ();
 sg13g2_decap_8 FILLER_21_3425 ();
 sg13g2_decap_8 FILLER_21_3432 ();
 sg13g2_decap_4 FILLER_21_3439 ();
 sg13g2_fill_2 FILLER_21_3443 ();
 sg13g2_decap_4 FILLER_21_3454 ();
 sg13g2_fill_1 FILLER_21_3462 ();
 sg13g2_decap_4 FILLER_21_3482 ();
 sg13g2_fill_2 FILLER_21_3486 ();
 sg13g2_decap_4 FILLER_21_3492 ();
 sg13g2_fill_2 FILLER_21_3496 ();
 sg13g2_decap_8 FILLER_21_3507 ();
 sg13g2_fill_2 FILLER_21_3514 ();
 sg13g2_fill_1 FILLER_21_3516 ();
 sg13g2_decap_4 FILLER_21_3521 ();
 sg13g2_fill_1 FILLER_21_3525 ();
 sg13g2_decap_4 FILLER_21_3535 ();
 sg13g2_fill_2 FILLER_21_3539 ();
 sg13g2_decap_8 FILLER_21_3549 ();
 sg13g2_decap_8 FILLER_21_3556 ();
 sg13g2_decap_8 FILLER_21_3563 ();
 sg13g2_decap_8 FILLER_21_3570 ();
 sg13g2_fill_2 FILLER_21_3577 ();
 sg13g2_fill_1 FILLER_21_3579 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_4 FILLER_22_7 ();
 sg13g2_fill_2 FILLER_22_45 ();
 sg13g2_decap_8 FILLER_22_65 ();
 sg13g2_fill_2 FILLER_22_72 ();
 sg13g2_fill_1 FILLER_22_74 ();
 sg13g2_decap_8 FILLER_22_104 ();
 sg13g2_decap_8 FILLER_22_111 ();
 sg13g2_decap_8 FILLER_22_118 ();
 sg13g2_decap_8 FILLER_22_125 ();
 sg13g2_decap_8 FILLER_22_132 ();
 sg13g2_decap_8 FILLER_22_139 ();
 sg13g2_fill_1 FILLER_22_164 ();
 sg13g2_decap_8 FILLER_22_179 ();
 sg13g2_decap_8 FILLER_22_186 ();
 sg13g2_decap_8 FILLER_22_193 ();
 sg13g2_fill_1 FILLER_22_200 ();
 sg13g2_decap_4 FILLER_22_216 ();
 sg13g2_decap_4 FILLER_22_243 ();
 sg13g2_fill_1 FILLER_22_247 ();
 sg13g2_decap_8 FILLER_22_254 ();
 sg13g2_fill_2 FILLER_22_266 ();
 sg13g2_decap_8 FILLER_22_276 ();
 sg13g2_fill_1 FILLER_22_283 ();
 sg13g2_fill_1 FILLER_22_288 ();
 sg13g2_decap_4 FILLER_22_295 ();
 sg13g2_fill_1 FILLER_22_299 ();
 sg13g2_decap_8 FILLER_22_313 ();
 sg13g2_fill_2 FILLER_22_320 ();
 sg13g2_fill_1 FILLER_22_322 ();
 sg13g2_decap_8 FILLER_22_329 ();
 sg13g2_decap_8 FILLER_22_336 ();
 sg13g2_decap_8 FILLER_22_343 ();
 sg13g2_decap_8 FILLER_22_350 ();
 sg13g2_fill_1 FILLER_22_357 ();
 sg13g2_decap_8 FILLER_22_383 ();
 sg13g2_decap_8 FILLER_22_390 ();
 sg13g2_decap_8 FILLER_22_440 ();
 sg13g2_decap_8 FILLER_22_447 ();
 sg13g2_decap_8 FILLER_22_463 ();
 sg13g2_decap_8 FILLER_22_470 ();
 sg13g2_decap_8 FILLER_22_477 ();
 sg13g2_decap_8 FILLER_22_484 ();
 sg13g2_decap_8 FILLER_22_491 ();
 sg13g2_decap_8 FILLER_22_498 ();
 sg13g2_decap_8 FILLER_22_505 ();
 sg13g2_decap_8 FILLER_22_512 ();
 sg13g2_fill_2 FILLER_22_519 ();
 sg13g2_fill_1 FILLER_22_521 ();
 sg13g2_decap_8 FILLER_22_552 ();
 sg13g2_decap_8 FILLER_22_559 ();
 sg13g2_decap_8 FILLER_22_566 ();
 sg13g2_decap_4 FILLER_22_573 ();
 sg13g2_fill_2 FILLER_22_577 ();
 sg13g2_decap_8 FILLER_22_589 ();
 sg13g2_decap_8 FILLER_22_596 ();
 sg13g2_decap_8 FILLER_22_603 ();
 sg13g2_decap_8 FILLER_22_610 ();
 sg13g2_decap_8 FILLER_22_617 ();
 sg13g2_decap_8 FILLER_22_624 ();
 sg13g2_decap_8 FILLER_22_631 ();
 sg13g2_decap_8 FILLER_22_638 ();
 sg13g2_fill_2 FILLER_22_645 ();
 sg13g2_fill_1 FILLER_22_647 ();
 sg13g2_fill_2 FILLER_22_656 ();
 sg13g2_fill_1 FILLER_22_658 ();
 sg13g2_decap_8 FILLER_22_668 ();
 sg13g2_fill_2 FILLER_22_675 ();
 sg13g2_fill_2 FILLER_22_700 ();
 sg13g2_decap_4 FILLER_22_710 ();
 sg13g2_decap_8 FILLER_22_729 ();
 sg13g2_decap_8 FILLER_22_736 ();
 sg13g2_decap_8 FILLER_22_743 ();
 sg13g2_decap_8 FILLER_22_750 ();
 sg13g2_decap_8 FILLER_22_757 ();
 sg13g2_fill_2 FILLER_22_764 ();
 sg13g2_fill_1 FILLER_22_766 ();
 sg13g2_decap_8 FILLER_22_803 ();
 sg13g2_decap_8 FILLER_22_810 ();
 sg13g2_decap_4 FILLER_22_817 ();
 sg13g2_fill_1 FILLER_22_821 ();
 sg13g2_decap_8 FILLER_22_848 ();
 sg13g2_decap_8 FILLER_22_855 ();
 sg13g2_decap_8 FILLER_22_862 ();
 sg13g2_decap_8 FILLER_22_869 ();
 sg13g2_decap_8 FILLER_22_876 ();
 sg13g2_decap_8 FILLER_22_883 ();
 sg13g2_decap_8 FILLER_22_890 ();
 sg13g2_decap_4 FILLER_22_897 ();
 sg13g2_fill_2 FILLER_22_901 ();
 sg13g2_decap_8 FILLER_22_929 ();
 sg13g2_decap_8 FILLER_22_936 ();
 sg13g2_decap_8 FILLER_22_943 ();
 sg13g2_decap_8 FILLER_22_950 ();
 sg13g2_decap_8 FILLER_22_957 ();
 sg13g2_decap_8 FILLER_22_964 ();
 sg13g2_decap_8 FILLER_22_971 ();
 sg13g2_fill_1 FILLER_22_978 ();
 sg13g2_decap_4 FILLER_22_987 ();
 sg13g2_decap_4 FILLER_22_1002 ();
 sg13g2_fill_2 FILLER_22_1006 ();
 sg13g2_decap_8 FILLER_22_1030 ();
 sg13g2_fill_2 FILLER_22_1037 ();
 sg13g2_decap_4 FILLER_22_1053 ();
 sg13g2_fill_2 FILLER_22_1057 ();
 sg13g2_decap_8 FILLER_22_1069 ();
 sg13g2_decap_8 FILLER_22_1076 ();
 sg13g2_decap_8 FILLER_22_1083 ();
 sg13g2_decap_8 FILLER_22_1090 ();
 sg13g2_decap_8 FILLER_22_1097 ();
 sg13g2_decap_8 FILLER_22_1104 ();
 sg13g2_decap_8 FILLER_22_1111 ();
 sg13g2_decap_8 FILLER_22_1118 ();
 sg13g2_decap_8 FILLER_22_1125 ();
 sg13g2_decap_8 FILLER_22_1132 ();
 sg13g2_decap_8 FILLER_22_1139 ();
 sg13g2_decap_8 FILLER_22_1146 ();
 sg13g2_decap_8 FILLER_22_1153 ();
 sg13g2_fill_1 FILLER_22_1160 ();
 sg13g2_decap_8 FILLER_22_1197 ();
 sg13g2_decap_8 FILLER_22_1204 ();
 sg13g2_decap_8 FILLER_22_1211 ();
 sg13g2_decap_4 FILLER_22_1218 ();
 sg13g2_fill_2 FILLER_22_1222 ();
 sg13g2_decap_8 FILLER_22_1229 ();
 sg13g2_decap_8 FILLER_22_1236 ();
 sg13g2_decap_8 FILLER_22_1243 ();
 sg13g2_decap_8 FILLER_22_1250 ();
 sg13g2_decap_8 FILLER_22_1257 ();
 sg13g2_decap_4 FILLER_22_1264 ();
 sg13g2_fill_1 FILLER_22_1268 ();
 sg13g2_decap_8 FILLER_22_1274 ();
 sg13g2_decap_8 FILLER_22_1281 ();
 sg13g2_decap_8 FILLER_22_1288 ();
 sg13g2_decap_4 FILLER_22_1295 ();
 sg13g2_fill_1 FILLER_22_1299 ();
 sg13g2_fill_2 FILLER_22_1346 ();
 sg13g2_fill_1 FILLER_22_1348 ();
 sg13g2_decap_8 FILLER_22_1375 ();
 sg13g2_decap_8 FILLER_22_1382 ();
 sg13g2_decap_8 FILLER_22_1389 ();
 sg13g2_decap_8 FILLER_22_1396 ();
 sg13g2_decap_8 FILLER_22_1403 ();
 sg13g2_decap_8 FILLER_22_1410 ();
 sg13g2_decap_4 FILLER_22_1417 ();
 sg13g2_fill_1 FILLER_22_1421 ();
 sg13g2_fill_1 FILLER_22_1437 ();
 sg13g2_decap_8 FILLER_22_1461 ();
 sg13g2_fill_2 FILLER_22_1483 ();
 sg13g2_fill_1 FILLER_22_1485 ();
 sg13g2_decap_8 FILLER_22_1527 ();
 sg13g2_decap_4 FILLER_22_1534 ();
 sg13g2_fill_2 FILLER_22_1538 ();
 sg13g2_decap_8 FILLER_22_1550 ();
 sg13g2_decap_8 FILLER_22_1557 ();
 sg13g2_decap_8 FILLER_22_1564 ();
 sg13g2_decap_4 FILLER_22_1571 ();
 sg13g2_fill_2 FILLER_22_1575 ();
 sg13g2_decap_8 FILLER_22_1595 ();
 sg13g2_decap_8 FILLER_22_1602 ();
 sg13g2_decap_8 FILLER_22_1609 ();
 sg13g2_decap_4 FILLER_22_1616 ();
 sg13g2_fill_2 FILLER_22_1620 ();
 sg13g2_fill_1 FILLER_22_1632 ();
 sg13g2_decap_8 FILLER_22_1637 ();
 sg13g2_decap_8 FILLER_22_1644 ();
 sg13g2_decap_8 FILLER_22_1651 ();
 sg13g2_fill_2 FILLER_22_1658 ();
 sg13g2_fill_1 FILLER_22_1660 ();
 sg13g2_decap_8 FILLER_22_1671 ();
 sg13g2_decap_8 FILLER_22_1678 ();
 sg13g2_decap_8 FILLER_22_1685 ();
 sg13g2_decap_8 FILLER_22_1692 ();
 sg13g2_decap_8 FILLER_22_1699 ();
 sg13g2_decap_8 FILLER_22_1706 ();
 sg13g2_decap_8 FILLER_22_1713 ();
 sg13g2_decap_8 FILLER_22_1720 ();
 sg13g2_decap_8 FILLER_22_1727 ();
 sg13g2_decap_8 FILLER_22_1734 ();
 sg13g2_decap_8 FILLER_22_1741 ();
 sg13g2_decap_8 FILLER_22_1748 ();
 sg13g2_decap_8 FILLER_22_1755 ();
 sg13g2_decap_8 FILLER_22_1762 ();
 sg13g2_decap_8 FILLER_22_1769 ();
 sg13g2_decap_8 FILLER_22_1776 ();
 sg13g2_decap_4 FILLER_22_1783 ();
 sg13g2_fill_1 FILLER_22_1787 ();
 sg13g2_decap_8 FILLER_22_1794 ();
 sg13g2_decap_8 FILLER_22_1801 ();
 sg13g2_decap_8 FILLER_22_1808 ();
 sg13g2_fill_2 FILLER_22_1815 ();
 sg13g2_decap_8 FILLER_22_1827 ();
 sg13g2_decap_8 FILLER_22_1834 ();
 sg13g2_decap_8 FILLER_22_1841 ();
 sg13g2_decap_8 FILLER_22_1848 ();
 sg13g2_decap_8 FILLER_22_1855 ();
 sg13g2_decap_8 FILLER_22_1862 ();
 sg13g2_decap_8 FILLER_22_1869 ();
 sg13g2_decap_4 FILLER_22_1876 ();
 sg13g2_fill_1 FILLER_22_1880 ();
 sg13g2_fill_2 FILLER_22_1891 ();
 sg13g2_fill_1 FILLER_22_1893 ();
 sg13g2_decap_8 FILLER_22_1905 ();
 sg13g2_decap_8 FILLER_22_1912 ();
 sg13g2_decap_8 FILLER_22_1919 ();
 sg13g2_decap_8 FILLER_22_1926 ();
 sg13g2_decap_4 FILLER_22_1933 ();
 sg13g2_fill_1 FILLER_22_1937 ();
 sg13g2_decap_8 FILLER_22_1964 ();
 sg13g2_decap_8 FILLER_22_1971 ();
 sg13g2_decap_8 FILLER_22_1978 ();
 sg13g2_decap_8 FILLER_22_1985 ();
 sg13g2_fill_2 FILLER_22_1992 ();
 sg13g2_fill_1 FILLER_22_1994 ();
 sg13g2_decap_8 FILLER_22_2021 ();
 sg13g2_decap_8 FILLER_22_2028 ();
 sg13g2_decap_8 FILLER_22_2035 ();
 sg13g2_decap_8 FILLER_22_2042 ();
 sg13g2_decap_4 FILLER_22_2049 ();
 sg13g2_fill_2 FILLER_22_2053 ();
 sg13g2_decap_8 FILLER_22_2077 ();
 sg13g2_decap_8 FILLER_22_2084 ();
 sg13g2_decap_8 FILLER_22_2091 ();
 sg13g2_decap_8 FILLER_22_2098 ();
 sg13g2_decap_8 FILLER_22_2105 ();
 sg13g2_decap_8 FILLER_22_2112 ();
 sg13g2_decap_8 FILLER_22_2119 ();
 sg13g2_decap_8 FILLER_22_2132 ();
 sg13g2_decap_8 FILLER_22_2139 ();
 sg13g2_fill_2 FILLER_22_2146 ();
 sg13g2_decap_8 FILLER_22_2184 ();
 sg13g2_decap_8 FILLER_22_2191 ();
 sg13g2_decap_4 FILLER_22_2198 ();
 sg13g2_fill_1 FILLER_22_2202 ();
 sg13g2_fill_2 FILLER_22_2211 ();
 sg13g2_decap_8 FILLER_22_2218 ();
 sg13g2_decap_8 FILLER_22_2225 ();
 sg13g2_decap_8 FILLER_22_2232 ();
 sg13g2_decap_8 FILLER_22_2239 ();
 sg13g2_decap_8 FILLER_22_2246 ();
 sg13g2_decap_8 FILLER_22_2253 ();
 sg13g2_decap_8 FILLER_22_2260 ();
 sg13g2_decap_8 FILLER_22_2267 ();
 sg13g2_decap_8 FILLER_22_2274 ();
 sg13g2_decap_8 FILLER_22_2281 ();
 sg13g2_decap_8 FILLER_22_2288 ();
 sg13g2_decap_8 FILLER_22_2295 ();
 sg13g2_decap_8 FILLER_22_2302 ();
 sg13g2_fill_2 FILLER_22_2309 ();
 sg13g2_decap_8 FILLER_22_2376 ();
 sg13g2_decap_8 FILLER_22_2383 ();
 sg13g2_decap_8 FILLER_22_2390 ();
 sg13g2_decap_8 FILLER_22_2397 ();
 sg13g2_decap_8 FILLER_22_2404 ();
 sg13g2_fill_2 FILLER_22_2411 ();
 sg13g2_decap_4 FILLER_22_2418 ();
 sg13g2_fill_1 FILLER_22_2422 ();
 sg13g2_decap_4 FILLER_22_2447 ();
 sg13g2_fill_2 FILLER_22_2451 ();
 sg13g2_decap_8 FILLER_22_2458 ();
 sg13g2_decap_8 FILLER_22_2465 ();
 sg13g2_decap_8 FILLER_22_2472 ();
 sg13g2_decap_8 FILLER_22_2479 ();
 sg13g2_decap_8 FILLER_22_2486 ();
 sg13g2_decap_8 FILLER_22_2493 ();
 sg13g2_decap_8 FILLER_22_2500 ();
 sg13g2_decap_8 FILLER_22_2507 ();
 sg13g2_decap_8 FILLER_22_2514 ();
 sg13g2_decap_8 FILLER_22_2521 ();
 sg13g2_decap_4 FILLER_22_2528 ();
 sg13g2_fill_1 FILLER_22_2566 ();
 sg13g2_fill_2 FILLER_22_2593 ();
 sg13g2_decap_4 FILLER_22_2601 ();
 sg13g2_decap_8 FILLER_22_2645 ();
 sg13g2_decap_8 FILLER_22_2652 ();
 sg13g2_fill_1 FILLER_22_2667 ();
 sg13g2_decap_4 FILLER_22_2674 ();
 sg13g2_fill_2 FILLER_22_2678 ();
 sg13g2_decap_8 FILLER_22_2724 ();
 sg13g2_decap_8 FILLER_22_2731 ();
 sg13g2_decap_4 FILLER_22_2738 ();
 sg13g2_decap_8 FILLER_22_2757 ();
 sg13g2_decap_8 FILLER_22_2764 ();
 sg13g2_decap_8 FILLER_22_2771 ();
 sg13g2_decap_8 FILLER_22_2778 ();
 sg13g2_decap_8 FILLER_22_2785 ();
 sg13g2_decap_8 FILLER_22_2792 ();
 sg13g2_decap_8 FILLER_22_2799 ();
 sg13g2_decap_8 FILLER_22_2806 ();
 sg13g2_decap_4 FILLER_22_2813 ();
 sg13g2_decap_8 FILLER_22_2846 ();
 sg13g2_decap_4 FILLER_22_2853 ();
 sg13g2_fill_1 FILLER_22_2857 ();
 sg13g2_decap_4 FILLER_22_2863 ();
 sg13g2_fill_1 FILLER_22_2867 ();
 sg13g2_decap_8 FILLER_22_2886 ();
 sg13g2_decap_8 FILLER_22_2893 ();
 sg13g2_decap_8 FILLER_22_2900 ();
 sg13g2_decap_4 FILLER_22_2907 ();
 sg13g2_fill_2 FILLER_22_2911 ();
 sg13g2_decap_8 FILLER_22_2918 ();
 sg13g2_fill_2 FILLER_22_2925 ();
 sg13g2_decap_8 FILLER_22_2932 ();
 sg13g2_fill_2 FILLER_22_2939 ();
 sg13g2_decap_8 FILLER_22_2960 ();
 sg13g2_decap_8 FILLER_22_2967 ();
 sg13g2_decap_8 FILLER_22_2974 ();
 sg13g2_decap_8 FILLER_22_2981 ();
 sg13g2_decap_8 FILLER_22_2988 ();
 sg13g2_fill_2 FILLER_22_2995 ();
 sg13g2_fill_1 FILLER_22_2997 ();
 sg13g2_decap_8 FILLER_22_3011 ();
 sg13g2_decap_8 FILLER_22_3018 ();
 sg13g2_decap_8 FILLER_22_3025 ();
 sg13g2_decap_8 FILLER_22_3032 ();
 sg13g2_decap_8 FILLER_22_3039 ();
 sg13g2_decap_8 FILLER_22_3046 ();
 sg13g2_decap_8 FILLER_22_3053 ();
 sg13g2_decap_8 FILLER_22_3060 ();
 sg13g2_decap_8 FILLER_22_3067 ();
 sg13g2_decap_4 FILLER_22_3074 ();
 sg13g2_fill_1 FILLER_22_3078 ();
 sg13g2_decap_8 FILLER_22_3089 ();
 sg13g2_fill_2 FILLER_22_3096 ();
 sg13g2_fill_1 FILLER_22_3124 ();
 sg13g2_decap_4 FILLER_22_3133 ();
 sg13g2_decap_8 FILLER_22_3160 ();
 sg13g2_decap_8 FILLER_22_3167 ();
 sg13g2_decap_8 FILLER_22_3174 ();
 sg13g2_decap_8 FILLER_22_3181 ();
 sg13g2_decap_8 FILLER_22_3188 ();
 sg13g2_decap_4 FILLER_22_3195 ();
 sg13g2_fill_1 FILLER_22_3199 ();
 sg13g2_decap_8 FILLER_22_3208 ();
 sg13g2_decap_4 FILLER_22_3215 ();
 sg13g2_decap_8 FILLER_22_3224 ();
 sg13g2_decap_4 FILLER_22_3231 ();
 sg13g2_decap_8 FILLER_22_3239 ();
 sg13g2_decap_8 FILLER_22_3246 ();
 sg13g2_decap_8 FILLER_22_3253 ();
 sg13g2_decap_8 FILLER_22_3286 ();
 sg13g2_decap_8 FILLER_22_3293 ();
 sg13g2_decap_8 FILLER_22_3300 ();
 sg13g2_decap_8 FILLER_22_3307 ();
 sg13g2_fill_2 FILLER_22_3314 ();
 sg13g2_fill_1 FILLER_22_3316 ();
 sg13g2_decap_8 FILLER_22_3343 ();
 sg13g2_decap_8 FILLER_22_3350 ();
 sg13g2_decap_8 FILLER_22_3357 ();
 sg13g2_decap_8 FILLER_22_3364 ();
 sg13g2_decap_8 FILLER_22_3371 ();
 sg13g2_fill_2 FILLER_22_3378 ();
 sg13g2_fill_1 FILLER_22_3380 ();
 sg13g2_fill_1 FILLER_22_3391 ();
 sg13g2_decap_8 FILLER_22_3418 ();
 sg13g2_decap_8 FILLER_22_3425 ();
 sg13g2_decap_8 FILLER_22_3432 ();
 sg13g2_decap_8 FILLER_22_3439 ();
 sg13g2_fill_2 FILLER_22_3446 ();
 sg13g2_decap_8 FILLER_22_3488 ();
 sg13g2_decap_8 FILLER_22_3495 ();
 sg13g2_decap_8 FILLER_22_3502 ();
 sg13g2_decap_8 FILLER_22_3509 ();
 sg13g2_decap_8 FILLER_22_3516 ();
 sg13g2_decap_8 FILLER_22_3523 ();
 sg13g2_decap_8 FILLER_22_3530 ();
 sg13g2_decap_8 FILLER_22_3537 ();
 sg13g2_decap_8 FILLER_22_3544 ();
 sg13g2_decap_8 FILLER_22_3551 ();
 sg13g2_decap_8 FILLER_22_3558 ();
 sg13g2_decap_8 FILLER_22_3565 ();
 sg13g2_decap_8 FILLER_22_3572 ();
 sg13g2_fill_1 FILLER_22_3579 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_fill_2 FILLER_23_28 ();
 sg13g2_fill_1 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_55 ();
 sg13g2_decap_8 FILLER_23_62 ();
 sg13g2_decap_8 FILLER_23_69 ();
 sg13g2_decap_8 FILLER_23_76 ();
 sg13g2_fill_2 FILLER_23_83 ();
 sg13g2_fill_1 FILLER_23_85 ();
 sg13g2_decap_8 FILLER_23_90 ();
 sg13g2_decap_4 FILLER_23_97 ();
 sg13g2_fill_1 FILLER_23_101 ();
 sg13g2_decap_8 FILLER_23_108 ();
 sg13g2_decap_8 FILLER_23_115 ();
 sg13g2_decap_8 FILLER_23_122 ();
 sg13g2_decap_8 FILLER_23_129 ();
 sg13g2_decap_8 FILLER_23_136 ();
 sg13g2_decap_8 FILLER_23_143 ();
 sg13g2_decap_8 FILLER_23_150 ();
 sg13g2_decap_8 FILLER_23_195 ();
 sg13g2_decap_4 FILLER_23_202 ();
 sg13g2_decap_4 FILLER_23_225 ();
 sg13g2_decap_8 FILLER_23_235 ();
 sg13g2_fill_2 FILLER_23_242 ();
 sg13g2_fill_1 FILLER_23_281 ();
 sg13g2_fill_2 FILLER_23_287 ();
 sg13g2_fill_2 FILLER_23_315 ();
 sg13g2_decap_8 FILLER_23_331 ();
 sg13g2_fill_1 FILLER_23_338 ();
 sg13g2_fill_1 FILLER_23_347 ();
 sg13g2_fill_2 FILLER_23_360 ();
 sg13g2_decap_8 FILLER_23_380 ();
 sg13g2_decap_8 FILLER_23_387 ();
 sg13g2_decap_8 FILLER_23_394 ();
 sg13g2_decap_8 FILLER_23_401 ();
 sg13g2_fill_1 FILLER_23_408 ();
 sg13g2_fill_2 FILLER_23_422 ();
 sg13g2_decap_8 FILLER_23_429 ();
 sg13g2_decap_8 FILLER_23_436 ();
 sg13g2_decap_8 FILLER_23_443 ();
 sg13g2_decap_8 FILLER_23_450 ();
 sg13g2_decap_8 FILLER_23_457 ();
 sg13g2_decap_8 FILLER_23_464 ();
 sg13g2_decap_8 FILLER_23_471 ();
 sg13g2_fill_1 FILLER_23_478 ();
 sg13g2_decap_8 FILLER_23_490 ();
 sg13g2_decap_8 FILLER_23_497 ();
 sg13g2_decap_8 FILLER_23_504 ();
 sg13g2_decap_8 FILLER_23_511 ();
 sg13g2_decap_8 FILLER_23_518 ();
 sg13g2_decap_8 FILLER_23_525 ();
 sg13g2_fill_2 FILLER_23_532 ();
 sg13g2_decap_4 FILLER_23_564 ();
 sg13g2_fill_2 FILLER_23_594 ();
 sg13g2_decap_8 FILLER_23_604 ();
 sg13g2_decap_8 FILLER_23_611 ();
 sg13g2_decap_8 FILLER_23_618 ();
 sg13g2_decap_8 FILLER_23_625 ();
 sg13g2_decap_4 FILLER_23_632 ();
 sg13g2_decap_4 FILLER_23_668 ();
 sg13g2_fill_2 FILLER_23_685 ();
 sg13g2_decap_8 FILLER_23_731 ();
 sg13g2_decap_8 FILLER_23_738 ();
 sg13g2_decap_8 FILLER_23_745 ();
 sg13g2_decap_8 FILLER_23_778 ();
 sg13g2_decap_8 FILLER_23_785 ();
 sg13g2_decap_8 FILLER_23_792 ();
 sg13g2_decap_8 FILLER_23_799 ();
 sg13g2_fill_2 FILLER_23_806 ();
 sg13g2_decap_8 FILLER_23_818 ();
 sg13g2_fill_1 FILLER_23_825 ();
 sg13g2_decap_8 FILLER_23_852 ();
 sg13g2_decap_8 FILLER_23_859 ();
 sg13g2_decap_8 FILLER_23_866 ();
 sg13g2_decap_8 FILLER_23_873 ();
 sg13g2_decap_8 FILLER_23_880 ();
 sg13g2_decap_8 FILLER_23_887 ();
 sg13g2_decap_8 FILLER_23_894 ();
 sg13g2_decap_8 FILLER_23_901 ();
 sg13g2_decap_8 FILLER_23_908 ();
 sg13g2_decap_8 FILLER_23_921 ();
 sg13g2_decap_8 FILLER_23_928 ();
 sg13g2_decap_4 FILLER_23_935 ();
 sg13g2_fill_1 FILLER_23_939 ();
 sg13g2_decap_8 FILLER_23_976 ();
 sg13g2_decap_8 FILLER_23_983 ();
 sg13g2_decap_8 FILLER_23_990 ();
 sg13g2_decap_8 FILLER_23_997 ();
 sg13g2_fill_1 FILLER_23_1004 ();
 sg13g2_fill_2 FILLER_23_1040 ();
 sg13g2_decap_8 FILLER_23_1045 ();
 sg13g2_decap_8 FILLER_23_1052 ();
 sg13g2_decap_8 FILLER_23_1059 ();
 sg13g2_decap_8 FILLER_23_1092 ();
 sg13g2_decap_8 FILLER_23_1099 ();
 sg13g2_fill_2 FILLER_23_1106 ();
 sg13g2_decap_8 FILLER_23_1150 ();
 sg13g2_decap_8 FILLER_23_1157 ();
 sg13g2_decap_4 FILLER_23_1164 ();
 sg13g2_fill_2 FILLER_23_1171 ();
 sg13g2_fill_1 FILLER_23_1173 ();
 sg13g2_decap_8 FILLER_23_1199 ();
 sg13g2_decap_8 FILLER_23_1206 ();
 sg13g2_decap_8 FILLER_23_1213 ();
 sg13g2_decap_8 FILLER_23_1220 ();
 sg13g2_decap_8 FILLER_23_1227 ();
 sg13g2_decap_4 FILLER_23_1234 ();
 sg13g2_fill_2 FILLER_23_1238 ();
 sg13g2_decap_8 FILLER_23_1266 ();
 sg13g2_decap_8 FILLER_23_1273 ();
 sg13g2_decap_8 FILLER_23_1280 ();
 sg13g2_decap_8 FILLER_23_1287 ();
 sg13g2_decap_4 FILLER_23_1294 ();
 sg13g2_fill_1 FILLER_23_1298 ();
 sg13g2_decap_8 FILLER_23_1335 ();
 sg13g2_decap_8 FILLER_23_1342 ();
 sg13g2_decap_8 FILLER_23_1349 ();
 sg13g2_decap_8 FILLER_23_1356 ();
 sg13g2_decap_8 FILLER_23_1363 ();
 sg13g2_decap_8 FILLER_23_1414 ();
 sg13g2_decap_8 FILLER_23_1421 ();
 sg13g2_decap_4 FILLER_23_1428 ();
 sg13g2_fill_2 FILLER_23_1432 ();
 sg13g2_fill_1 FILLER_23_1446 ();
 sg13g2_fill_2 FILLER_23_1461 ();
 sg13g2_decap_8 FILLER_23_1489 ();
 sg13g2_decap_8 FILLER_23_1496 ();
 sg13g2_decap_8 FILLER_23_1503 ();
 sg13g2_decap_8 FILLER_23_1510 ();
 sg13g2_decap_8 FILLER_23_1517 ();
 sg13g2_decap_8 FILLER_23_1524 ();
 sg13g2_decap_8 FILLER_23_1557 ();
 sg13g2_decap_8 FILLER_23_1564 ();
 sg13g2_decap_8 FILLER_23_1571 ();
 sg13g2_fill_2 FILLER_23_1578 ();
 sg13g2_decap_8 FILLER_23_1595 ();
 sg13g2_decap_8 FILLER_23_1602 ();
 sg13g2_decap_4 FILLER_23_1617 ();
 sg13g2_fill_1 FILLER_23_1621 ();
 sg13g2_decap_8 FILLER_23_1632 ();
 sg13g2_fill_2 FILLER_23_1639 ();
 sg13g2_fill_1 FILLER_23_1672 ();
 sg13g2_decap_8 FILLER_23_1699 ();
 sg13g2_decap_8 FILLER_23_1706 ();
 sg13g2_decap_8 FILLER_23_1713 ();
 sg13g2_fill_1 FILLER_23_1720 ();
 sg13g2_decap_8 FILLER_23_1747 ();
 sg13g2_decap_8 FILLER_23_1754 ();
 sg13g2_decap_8 FILLER_23_1761 ();
 sg13g2_fill_2 FILLER_23_1768 ();
 sg13g2_fill_1 FILLER_23_1770 ();
 sg13g2_fill_1 FILLER_23_1780 ();
 sg13g2_decap_8 FILLER_23_1789 ();
 sg13g2_decap_8 FILLER_23_1796 ();
 sg13g2_decap_8 FILLER_23_1803 ();
 sg13g2_decap_8 FILLER_23_1810 ();
 sg13g2_decap_8 FILLER_23_1817 ();
 sg13g2_decap_8 FILLER_23_1824 ();
 sg13g2_decap_8 FILLER_23_1831 ();
 sg13g2_decap_8 FILLER_23_1838 ();
 sg13g2_decap_8 FILLER_23_1860 ();
 sg13g2_decap_8 FILLER_23_1867 ();
 sg13g2_decap_8 FILLER_23_1874 ();
 sg13g2_fill_1 FILLER_23_1881 ();
 sg13g2_decap_8 FILLER_23_1908 ();
 sg13g2_decap_8 FILLER_23_1915 ();
 sg13g2_decap_8 FILLER_23_1922 ();
 sg13g2_decap_8 FILLER_23_1929 ();
 sg13g2_decap_8 FILLER_23_1936 ();
 sg13g2_decap_8 FILLER_23_1943 ();
 sg13g2_fill_2 FILLER_23_1950 ();
 sg13g2_decap_8 FILLER_23_1956 ();
 sg13g2_fill_1 FILLER_23_1963 ();
 sg13g2_decap_8 FILLER_23_1968 ();
 sg13g2_decap_4 FILLER_23_1975 ();
 sg13g2_fill_2 FILLER_23_1979 ();
 sg13g2_decap_8 FILLER_23_1991 ();
 sg13g2_decap_8 FILLER_23_1998 ();
 sg13g2_decap_8 FILLER_23_2005 ();
 sg13g2_decap_8 FILLER_23_2012 ();
 sg13g2_decap_8 FILLER_23_2019 ();
 sg13g2_fill_2 FILLER_23_2026 ();
 sg13g2_decap_8 FILLER_23_2033 ();
 sg13g2_decap_8 FILLER_23_2040 ();
 sg13g2_fill_1 FILLER_23_2047 ();
 sg13g2_decap_8 FILLER_23_2071 ();
 sg13g2_decap_8 FILLER_23_2078 ();
 sg13g2_decap_8 FILLER_23_2085 ();
 sg13g2_decap_8 FILLER_23_2092 ();
 sg13g2_fill_2 FILLER_23_2111 ();
 sg13g2_decap_8 FILLER_23_2123 ();
 sg13g2_decap_8 FILLER_23_2130 ();
 sg13g2_decap_4 FILLER_23_2137 ();
 sg13g2_decap_8 FILLER_23_2151 ();
 sg13g2_decap_8 FILLER_23_2158 ();
 sg13g2_decap_8 FILLER_23_2165 ();
 sg13g2_decap_8 FILLER_23_2172 ();
 sg13g2_decap_8 FILLER_23_2179 ();
 sg13g2_decap_8 FILLER_23_2186 ();
 sg13g2_decap_4 FILLER_23_2193 ();
 sg13g2_fill_2 FILLER_23_2197 ();
 sg13g2_decap_8 FILLER_23_2241 ();
 sg13g2_decap_4 FILLER_23_2248 ();
 sg13g2_fill_1 FILLER_23_2252 ();
 sg13g2_decap_8 FILLER_23_2283 ();
 sg13g2_decap_8 FILLER_23_2290 ();
 sg13g2_decap_8 FILLER_23_2297 ();
 sg13g2_fill_1 FILLER_23_2304 ();
 sg13g2_decap_8 FILLER_23_2315 ();
 sg13g2_decap_8 FILLER_23_2322 ();
 sg13g2_decap_8 FILLER_23_2329 ();
 sg13g2_decap_8 FILLER_23_2336 ();
 sg13g2_decap_8 FILLER_23_2343 ();
 sg13g2_fill_1 FILLER_23_2350 ();
 sg13g2_decap_8 FILLER_23_2356 ();
 sg13g2_decap_8 FILLER_23_2363 ();
 sg13g2_decap_8 FILLER_23_2370 ();
 sg13g2_decap_8 FILLER_23_2377 ();
 sg13g2_decap_8 FILLER_23_2384 ();
 sg13g2_decap_8 FILLER_23_2391 ();
 sg13g2_decap_8 FILLER_23_2398 ();
 sg13g2_fill_1 FILLER_23_2405 ();
 sg13g2_decap_4 FILLER_23_2428 ();
 sg13g2_fill_1 FILLER_23_2438 ();
 sg13g2_decap_4 FILLER_23_2445 ();
 sg13g2_decap_8 FILLER_23_2483 ();
 sg13g2_fill_2 FILLER_23_2490 ();
 sg13g2_fill_1 FILLER_23_2492 ();
 sg13g2_decap_8 FILLER_23_2519 ();
 sg13g2_decap_8 FILLER_23_2526 ();
 sg13g2_decap_4 FILLER_23_2533 ();
 sg13g2_fill_2 FILLER_23_2537 ();
 sg13g2_decap_8 FILLER_23_2544 ();
 sg13g2_fill_1 FILLER_23_2551 ();
 sg13g2_decap_8 FILLER_23_2557 ();
 sg13g2_decap_8 FILLER_23_2574 ();
 sg13g2_decap_8 FILLER_23_2581 ();
 sg13g2_decap_8 FILLER_23_2588 ();
 sg13g2_decap_8 FILLER_23_2595 ();
 sg13g2_decap_4 FILLER_23_2602 ();
 sg13g2_fill_2 FILLER_23_2606 ();
 sg13g2_decap_8 FILLER_23_2637 ();
 sg13g2_fill_2 FILLER_23_2644 ();
 sg13g2_fill_1 FILLER_23_2646 ();
 sg13g2_decap_8 FILLER_23_2652 ();
 sg13g2_fill_2 FILLER_23_2659 ();
 sg13g2_decap_8 FILLER_23_2665 ();
 sg13g2_decap_8 FILLER_23_2672 ();
 sg13g2_decap_4 FILLER_23_2679 ();
 sg13g2_decap_8 FILLER_23_2701 ();
 sg13g2_decap_8 FILLER_23_2708 ();
 sg13g2_decap_8 FILLER_23_2715 ();
 sg13g2_fill_1 FILLER_23_2722 ();
 sg13g2_fill_2 FILLER_23_2731 ();
 sg13g2_fill_2 FILLER_23_2754 ();
 sg13g2_fill_2 FILLER_23_2766 ();
 sg13g2_decap_8 FILLER_23_2794 ();
 sg13g2_decap_8 FILLER_23_2801 ();
 sg13g2_fill_2 FILLER_23_2808 ();
 sg13g2_fill_1 FILLER_23_2824 ();
 sg13g2_decap_8 FILLER_23_2844 ();
 sg13g2_decap_8 FILLER_23_2851 ();
 sg13g2_decap_4 FILLER_23_2858 ();
 sg13g2_decap_8 FILLER_23_2892 ();
 sg13g2_decap_8 FILLER_23_2899 ();
 sg13g2_decap_8 FILLER_23_2906 ();
 sg13g2_decap_8 FILLER_23_2913 ();
 sg13g2_decap_8 FILLER_23_2920 ();
 sg13g2_decap_8 FILLER_23_2927 ();
 sg13g2_decap_8 FILLER_23_2934 ();
 sg13g2_decap_4 FILLER_23_2941 ();
 sg13g2_decap_8 FILLER_23_2958 ();
 sg13g2_decap_8 FILLER_23_2965 ();
 sg13g2_decap_8 FILLER_23_2972 ();
 sg13g2_decap_8 FILLER_23_2979 ();
 sg13g2_decap_8 FILLER_23_2986 ();
 sg13g2_decap_8 FILLER_23_2993 ();
 sg13g2_decap_8 FILLER_23_3000 ();
 sg13g2_decap_8 FILLER_23_3007 ();
 sg13g2_decap_8 FILLER_23_3014 ();
 sg13g2_decap_8 FILLER_23_3021 ();
 sg13g2_fill_2 FILLER_23_3028 ();
 sg13g2_fill_1 FILLER_23_3030 ();
 sg13g2_decap_8 FILLER_23_3057 ();
 sg13g2_decap_8 FILLER_23_3064 ();
 sg13g2_fill_1 FILLER_23_3071 ();
 sg13g2_decap_8 FILLER_23_3082 ();
 sg13g2_decap_8 FILLER_23_3089 ();
 sg13g2_decap_8 FILLER_23_3096 ();
 sg13g2_decap_8 FILLER_23_3103 ();
 sg13g2_decap_8 FILLER_23_3110 ();
 sg13g2_decap_8 FILLER_23_3117 ();
 sg13g2_decap_8 FILLER_23_3124 ();
 sg13g2_decap_8 FILLER_23_3131 ();
 sg13g2_decap_8 FILLER_23_3138 ();
 sg13g2_decap_8 FILLER_23_3145 ();
 sg13g2_decap_8 FILLER_23_3152 ();
 sg13g2_decap_8 FILLER_23_3159 ();
 sg13g2_decap_8 FILLER_23_3166 ();
 sg13g2_decap_8 FILLER_23_3173 ();
 sg13g2_decap_8 FILLER_23_3180 ();
 sg13g2_decap_8 FILLER_23_3187 ();
 sg13g2_decap_8 FILLER_23_3194 ();
 sg13g2_decap_4 FILLER_23_3201 ();
 sg13g2_fill_1 FILLER_23_3205 ();
 sg13g2_fill_2 FILLER_23_3232 ();
 sg13g2_fill_1 FILLER_23_3234 ();
 sg13g2_decap_8 FILLER_23_3241 ();
 sg13g2_decap_8 FILLER_23_3248 ();
 sg13g2_decap_8 FILLER_23_3255 ();
 sg13g2_decap_8 FILLER_23_3272 ();
 sg13g2_decap_8 FILLER_23_3279 ();
 sg13g2_decap_8 FILLER_23_3286 ();
 sg13g2_decap_4 FILLER_23_3293 ();
 sg13g2_fill_1 FILLER_23_3307 ();
 sg13g2_decap_8 FILLER_23_3318 ();
 sg13g2_decap_8 FILLER_23_3325 ();
 sg13g2_decap_8 FILLER_23_3332 ();
 sg13g2_decap_8 FILLER_23_3339 ();
 sg13g2_decap_8 FILLER_23_3346 ();
 sg13g2_fill_1 FILLER_23_3353 ();
 sg13g2_fill_1 FILLER_23_3364 ();
 sg13g2_decap_8 FILLER_23_3417 ();
 sg13g2_decap_8 FILLER_23_3424 ();
 sg13g2_decap_8 FILLER_23_3431 ();
 sg13g2_decap_8 FILLER_23_3438 ();
 sg13g2_decap_8 FILLER_23_3445 ();
 sg13g2_fill_1 FILLER_23_3452 ();
 sg13g2_decap_8 FILLER_23_3458 ();
 sg13g2_decap_8 FILLER_23_3465 ();
 sg13g2_decap_8 FILLER_23_3472 ();
 sg13g2_decap_8 FILLER_23_3479 ();
 sg13g2_decap_8 FILLER_23_3486 ();
 sg13g2_decap_8 FILLER_23_3493 ();
 sg13g2_fill_1 FILLER_23_3500 ();
 sg13g2_decap_8 FILLER_23_3506 ();
 sg13g2_decap_8 FILLER_23_3513 ();
 sg13g2_decap_8 FILLER_23_3520 ();
 sg13g2_decap_4 FILLER_23_3527 ();
 sg13g2_fill_1 FILLER_23_3535 ();
 sg13g2_decap_8 FILLER_23_3562 ();
 sg13g2_decap_8 FILLER_23_3569 ();
 sg13g2_decap_4 FILLER_23_3576 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_fill_2 FILLER_24_21 ();
 sg13g2_fill_1 FILLER_24_23 ();
 sg13g2_fill_1 FILLER_24_29 ();
 sg13g2_decap_8 FILLER_24_47 ();
 sg13g2_decap_8 FILLER_24_54 ();
 sg13g2_decap_8 FILLER_24_61 ();
 sg13g2_decap_8 FILLER_24_68 ();
 sg13g2_fill_2 FILLER_24_75 ();
 sg13g2_decap_8 FILLER_24_110 ();
 sg13g2_decap_8 FILLER_24_117 ();
 sg13g2_decap_8 FILLER_24_124 ();
 sg13g2_decap_8 FILLER_24_131 ();
 sg13g2_decap_8 FILLER_24_138 ();
 sg13g2_decap_8 FILLER_24_145 ();
 sg13g2_decap_8 FILLER_24_152 ();
 sg13g2_decap_4 FILLER_24_159 ();
 sg13g2_fill_2 FILLER_24_163 ();
 sg13g2_decap_8 FILLER_24_168 ();
 sg13g2_decap_4 FILLER_24_175 ();
 sg13g2_fill_1 FILLER_24_179 ();
 sg13g2_decap_8 FILLER_24_189 ();
 sg13g2_decap_8 FILLER_24_196 ();
 sg13g2_decap_8 FILLER_24_203 ();
 sg13g2_fill_2 FILLER_24_210 ();
 sg13g2_decap_8 FILLER_24_227 ();
 sg13g2_decap_8 FILLER_24_234 ();
 sg13g2_decap_8 FILLER_24_241 ();
 sg13g2_decap_8 FILLER_24_248 ();
 sg13g2_decap_4 FILLER_24_255 ();
 sg13g2_fill_2 FILLER_24_259 ();
 sg13g2_fill_1 FILLER_24_273 ();
 sg13g2_decap_8 FILLER_24_286 ();
 sg13g2_decap_8 FILLER_24_293 ();
 sg13g2_decap_4 FILLER_24_300 ();
 sg13g2_fill_2 FILLER_24_307 ();
 sg13g2_fill_1 FILLER_24_309 ();
 sg13g2_decap_4 FILLER_24_319 ();
 sg13g2_decap_8 FILLER_24_334 ();
 sg13g2_decap_4 FILLER_24_341 ();
 sg13g2_decap_8 FILLER_24_350 ();
 sg13g2_decap_8 FILLER_24_357 ();
 sg13g2_decap_4 FILLER_24_364 ();
 sg13g2_decap_8 FILLER_24_376 ();
 sg13g2_decap_8 FILLER_24_383 ();
 sg13g2_decap_8 FILLER_24_390 ();
 sg13g2_decap_8 FILLER_24_397 ();
 sg13g2_decap_8 FILLER_24_404 ();
 sg13g2_decap_8 FILLER_24_411 ();
 sg13g2_decap_8 FILLER_24_418 ();
 sg13g2_decap_8 FILLER_24_425 ();
 sg13g2_decap_8 FILLER_24_432 ();
 sg13g2_decap_8 FILLER_24_439 ();
 sg13g2_decap_8 FILLER_24_446 ();
 sg13g2_decap_8 FILLER_24_453 ();
 sg13g2_decap_8 FILLER_24_460 ();
 sg13g2_fill_2 FILLER_24_467 ();
 sg13g2_decap_8 FILLER_24_495 ();
 sg13g2_decap_8 FILLER_24_502 ();
 sg13g2_decap_8 FILLER_24_509 ();
 sg13g2_decap_8 FILLER_24_516 ();
 sg13g2_decap_8 FILLER_24_523 ();
 sg13g2_decap_8 FILLER_24_530 ();
 sg13g2_fill_2 FILLER_24_537 ();
 sg13g2_fill_2 FILLER_24_543 ();
 sg13g2_fill_1 FILLER_24_545 ();
 sg13g2_fill_2 FILLER_24_556 ();
 sg13g2_decap_8 FILLER_24_562 ();
 sg13g2_decap_8 FILLER_24_569 ();
 sg13g2_fill_1 FILLER_24_576 ();
 sg13g2_decap_8 FILLER_24_580 ();
 sg13g2_fill_1 FILLER_24_587 ();
 sg13g2_decap_8 FILLER_24_596 ();
 sg13g2_decap_8 FILLER_24_603 ();
 sg13g2_decap_8 FILLER_24_610 ();
 sg13g2_decap_8 FILLER_24_617 ();
 sg13g2_decap_8 FILLER_24_624 ();
 sg13g2_decap_8 FILLER_24_631 ();
 sg13g2_fill_2 FILLER_24_638 ();
 sg13g2_fill_1 FILLER_24_640 ();
 sg13g2_decap_4 FILLER_24_657 ();
 sg13g2_fill_1 FILLER_24_661 ();
 sg13g2_decap_8 FILLER_24_676 ();
 sg13g2_decap_8 FILLER_24_683 ();
 sg13g2_decap_8 FILLER_24_690 ();
 sg13g2_decap_4 FILLER_24_697 ();
 sg13g2_fill_2 FILLER_24_701 ();
 sg13g2_decap_4 FILLER_24_708 ();
 sg13g2_decap_8 FILLER_24_727 ();
 sg13g2_decap_8 FILLER_24_734 ();
 sg13g2_decap_4 FILLER_24_741 ();
 sg13g2_fill_2 FILLER_24_745 ();
 sg13g2_decap_8 FILLER_24_757 ();
 sg13g2_decap_8 FILLER_24_764 ();
 sg13g2_decap_8 FILLER_24_771 ();
 sg13g2_decap_8 FILLER_24_778 ();
 sg13g2_decap_8 FILLER_24_785 ();
 sg13g2_decap_8 FILLER_24_792 ();
 sg13g2_decap_8 FILLER_24_799 ();
 sg13g2_decap_8 FILLER_24_806 ();
 sg13g2_decap_8 FILLER_24_813 ();
 sg13g2_decap_8 FILLER_24_820 ();
 sg13g2_fill_2 FILLER_24_827 ();
 sg13g2_decap_8 FILLER_24_865 ();
 sg13g2_decap_4 FILLER_24_872 ();
 sg13g2_decap_8 FILLER_24_925 ();
 sg13g2_decap_8 FILLER_24_932 ();
 sg13g2_decap_8 FILLER_24_975 ();
 sg13g2_decap_8 FILLER_24_982 ();
 sg13g2_decap_8 FILLER_24_989 ();
 sg13g2_decap_8 FILLER_24_996 ();
 sg13g2_decap_8 FILLER_24_1003 ();
 sg13g2_fill_1 FILLER_24_1019 ();
 sg13g2_decap_8 FILLER_24_1040 ();
 sg13g2_decap_8 FILLER_24_1047 ();
 sg13g2_decap_8 FILLER_24_1054 ();
 sg13g2_decap_8 FILLER_24_1061 ();
 sg13g2_decap_8 FILLER_24_1068 ();
 sg13g2_decap_8 FILLER_24_1075 ();
 sg13g2_decap_8 FILLER_24_1082 ();
 sg13g2_decap_8 FILLER_24_1089 ();
 sg13g2_decap_8 FILLER_24_1096 ();
 sg13g2_decap_8 FILLER_24_1103 ();
 sg13g2_decap_8 FILLER_24_1110 ();
 sg13g2_decap_8 FILLER_24_1117 ();
 sg13g2_decap_8 FILLER_24_1124 ();
 sg13g2_decap_8 FILLER_24_1131 ();
 sg13g2_decap_8 FILLER_24_1138 ();
 sg13g2_decap_8 FILLER_24_1145 ();
 sg13g2_decap_8 FILLER_24_1152 ();
 sg13g2_decap_4 FILLER_24_1159 ();
 sg13g2_fill_2 FILLER_24_1163 ();
 sg13g2_decap_8 FILLER_24_1178 ();
 sg13g2_decap_8 FILLER_24_1185 ();
 sg13g2_decap_8 FILLER_24_1192 ();
 sg13g2_decap_8 FILLER_24_1199 ();
 sg13g2_decap_8 FILLER_24_1206 ();
 sg13g2_decap_8 FILLER_24_1213 ();
 sg13g2_decap_8 FILLER_24_1220 ();
 sg13g2_decap_8 FILLER_24_1227 ();
 sg13g2_decap_8 FILLER_24_1234 ();
 sg13g2_decap_8 FILLER_24_1241 ();
 sg13g2_decap_8 FILLER_24_1248 ();
 sg13g2_fill_2 FILLER_24_1255 ();
 sg13g2_decap_8 FILLER_24_1283 ();
 sg13g2_decap_8 FILLER_24_1290 ();
 sg13g2_decap_8 FILLER_24_1297 ();
 sg13g2_decap_8 FILLER_24_1304 ();
 sg13g2_decap_8 FILLER_24_1311 ();
 sg13g2_decap_8 FILLER_24_1318 ();
 sg13g2_decap_8 FILLER_24_1325 ();
 sg13g2_decap_8 FILLER_24_1332 ();
 sg13g2_decap_8 FILLER_24_1339 ();
 sg13g2_decap_8 FILLER_24_1346 ();
 sg13g2_decap_8 FILLER_24_1353 ();
 sg13g2_decap_8 FILLER_24_1360 ();
 sg13g2_decap_8 FILLER_24_1367 ();
 sg13g2_decap_8 FILLER_24_1374 ();
 sg13g2_decap_8 FILLER_24_1381 ();
 sg13g2_decap_8 FILLER_24_1388 ();
 sg13g2_decap_8 FILLER_24_1395 ();
 sg13g2_decap_8 FILLER_24_1402 ();
 sg13g2_decap_8 FILLER_24_1409 ();
 sg13g2_decap_8 FILLER_24_1416 ();
 sg13g2_decap_8 FILLER_24_1423 ();
 sg13g2_fill_1 FILLER_24_1430 ();
 sg13g2_decap_4 FILLER_24_1443 ();
 sg13g2_decap_8 FILLER_24_1450 ();
 sg13g2_decap_8 FILLER_24_1457 ();
 sg13g2_fill_2 FILLER_24_1472 ();
 sg13g2_decap_8 FILLER_24_1480 ();
 sg13g2_fill_1 FILLER_24_1487 ();
 sg13g2_decap_8 FILLER_24_1501 ();
 sg13g2_decap_8 FILLER_24_1508 ();
 sg13g2_decap_8 FILLER_24_1515 ();
 sg13g2_decap_8 FILLER_24_1522 ();
 sg13g2_decap_8 FILLER_24_1529 ();
 sg13g2_decap_8 FILLER_24_1536 ();
 sg13g2_decap_8 FILLER_24_1543 ();
 sg13g2_decap_8 FILLER_24_1550 ();
 sg13g2_decap_8 FILLER_24_1557 ();
 sg13g2_fill_1 FILLER_24_1564 ();
 sg13g2_decap_8 FILLER_24_1575 ();
 sg13g2_decap_8 FILLER_24_1582 ();
 sg13g2_decap_8 FILLER_24_1589 ();
 sg13g2_decap_8 FILLER_24_1596 ();
 sg13g2_decap_8 FILLER_24_1603 ();
 sg13g2_fill_2 FILLER_24_1610 ();
 sg13g2_decap_8 FILLER_24_1618 ();
 sg13g2_decap_8 FILLER_24_1625 ();
 sg13g2_decap_8 FILLER_24_1632 ();
 sg13g2_fill_2 FILLER_24_1665 ();
 sg13g2_fill_1 FILLER_24_1667 ();
 sg13g2_decap_8 FILLER_24_1676 ();
 sg13g2_decap_8 FILLER_24_1683 ();
 sg13g2_decap_8 FILLER_24_1690 ();
 sg13g2_decap_8 FILLER_24_1697 ();
 sg13g2_decap_8 FILLER_24_1704 ();
 sg13g2_decap_8 FILLER_24_1711 ();
 sg13g2_decap_4 FILLER_24_1718 ();
 sg13g2_fill_2 FILLER_24_1758 ();
 sg13g2_decap_4 FILLER_24_1766 ();
 sg13g2_fill_2 FILLER_24_1770 ();
 sg13g2_decap_8 FILLER_24_1812 ();
 sg13g2_fill_2 FILLER_24_1819 ();
 sg13g2_decap_8 FILLER_24_1831 ();
 sg13g2_decap_4 FILLER_24_1838 ();
 sg13g2_fill_1 FILLER_24_1842 ();
 sg13g2_decap_8 FILLER_24_1869 ();
 sg13g2_decap_8 FILLER_24_1876 ();
 sg13g2_decap_8 FILLER_24_1883 ();
 sg13g2_fill_2 FILLER_24_1890 ();
 sg13g2_fill_1 FILLER_24_1892 ();
 sg13g2_decap_8 FILLER_24_1919 ();
 sg13g2_decap_8 FILLER_24_1926 ();
 sg13g2_decap_4 FILLER_24_1933 ();
 sg13g2_fill_1 FILLER_24_1937 ();
 sg13g2_decap_8 FILLER_24_1948 ();
 sg13g2_decap_8 FILLER_24_1955 ();
 sg13g2_decap_8 FILLER_24_1962 ();
 sg13g2_decap_8 FILLER_24_1969 ();
 sg13g2_decap_8 FILLER_24_1976 ();
 sg13g2_decap_8 FILLER_24_1983 ();
 sg13g2_decap_8 FILLER_24_1990 ();
 sg13g2_decap_8 FILLER_24_1997 ();
 sg13g2_decap_8 FILLER_24_2004 ();
 sg13g2_decap_8 FILLER_24_2011 ();
 sg13g2_decap_8 FILLER_24_2018 ();
 sg13g2_decap_8 FILLER_24_2025 ();
 sg13g2_decap_8 FILLER_24_2032 ();
 sg13g2_decap_8 FILLER_24_2039 ();
 sg13g2_decap_8 FILLER_24_2046 ();
 sg13g2_fill_2 FILLER_24_2053 ();
 sg13g2_decap_8 FILLER_24_2066 ();
 sg13g2_decap_8 FILLER_24_2073 ();
 sg13g2_fill_2 FILLER_24_2080 ();
 sg13g2_fill_1 FILLER_24_2092 ();
 sg13g2_decap_4 FILLER_24_2116 ();
 sg13g2_fill_2 FILLER_24_2120 ();
 sg13g2_decap_8 FILLER_24_2174 ();
 sg13g2_fill_1 FILLER_24_2181 ();
 sg13g2_decap_8 FILLER_24_2190 ();
 sg13g2_decap_8 FILLER_24_2197 ();
 sg13g2_decap_4 FILLER_24_2204 ();
 sg13g2_fill_1 FILLER_24_2208 ();
 sg13g2_decap_8 FILLER_24_2212 ();
 sg13g2_decap_8 FILLER_24_2219 ();
 sg13g2_fill_1 FILLER_24_2226 ();
 sg13g2_decap_8 FILLER_24_2233 ();
 sg13g2_decap_8 FILLER_24_2240 ();
 sg13g2_fill_2 FILLER_24_2247 ();
 sg13g2_fill_1 FILLER_24_2249 ();
 sg13g2_decap_8 FILLER_24_2258 ();
 sg13g2_fill_2 FILLER_24_2265 ();
 sg13g2_decap_8 FILLER_24_2293 ();
 sg13g2_decap_8 FILLER_24_2300 ();
 sg13g2_decap_8 FILLER_24_2307 ();
 sg13g2_fill_2 FILLER_24_2314 ();
 sg13g2_decap_8 FILLER_24_2335 ();
 sg13g2_decap_8 FILLER_24_2342 ();
 sg13g2_decap_8 FILLER_24_2349 ();
 sg13g2_decap_8 FILLER_24_2356 ();
 sg13g2_decap_8 FILLER_24_2363 ();
 sg13g2_decap_8 FILLER_24_2370 ();
 sg13g2_decap_8 FILLER_24_2377 ();
 sg13g2_decap_8 FILLER_24_2384 ();
 sg13g2_decap_8 FILLER_24_2391 ();
 sg13g2_decap_4 FILLER_24_2398 ();
 sg13g2_fill_2 FILLER_24_2402 ();
 sg13g2_decap_4 FILLER_24_2450 ();
 sg13g2_fill_2 FILLER_24_2454 ();
 sg13g2_decap_8 FILLER_24_2460 ();
 sg13g2_decap_8 FILLER_24_2467 ();
 sg13g2_decap_8 FILLER_24_2474 ();
 sg13g2_decap_8 FILLER_24_2481 ();
 sg13g2_decap_8 FILLER_24_2498 ();
 sg13g2_decap_4 FILLER_24_2505 ();
 sg13g2_decap_8 FILLER_24_2515 ();
 sg13g2_fill_2 FILLER_24_2522 ();
 sg13g2_fill_1 FILLER_24_2524 ();
 sg13g2_decap_8 FILLER_24_2542 ();
 sg13g2_decap_8 FILLER_24_2549 ();
 sg13g2_decap_8 FILLER_24_2556 ();
 sg13g2_decap_8 FILLER_24_2563 ();
 sg13g2_decap_8 FILLER_24_2570 ();
 sg13g2_decap_8 FILLER_24_2577 ();
 sg13g2_decap_8 FILLER_24_2584 ();
 sg13g2_decap_8 FILLER_24_2591 ();
 sg13g2_decap_8 FILLER_24_2598 ();
 sg13g2_decap_8 FILLER_24_2605 ();
 sg13g2_fill_1 FILLER_24_2612 ();
 sg13g2_decap_8 FILLER_24_2623 ();
 sg13g2_decap_8 FILLER_24_2630 ();
 sg13g2_decap_8 FILLER_24_2637 ();
 sg13g2_decap_8 FILLER_24_2644 ();
 sg13g2_decap_8 FILLER_24_2651 ();
 sg13g2_fill_2 FILLER_24_2658 ();
 sg13g2_decap_4 FILLER_24_2666 ();
 sg13g2_fill_1 FILLER_24_2670 ();
 sg13g2_decap_8 FILLER_24_2677 ();
 sg13g2_decap_8 FILLER_24_2684 ();
 sg13g2_decap_8 FILLER_24_2717 ();
 sg13g2_decap_8 FILLER_24_2724 ();
 sg13g2_decap_8 FILLER_24_2731 ();
 sg13g2_decap_8 FILLER_24_2738 ();
 sg13g2_decap_4 FILLER_24_2745 ();
 sg13g2_decap_8 FILLER_24_2752 ();
 sg13g2_decap_8 FILLER_24_2759 ();
 sg13g2_decap_8 FILLER_24_2766 ();
 sg13g2_fill_1 FILLER_24_2773 ();
 sg13g2_decap_8 FILLER_24_2800 ();
 sg13g2_decap_4 FILLER_24_2807 ();
 sg13g2_fill_1 FILLER_24_2811 ();
 sg13g2_decap_8 FILLER_24_2841 ();
 sg13g2_decap_8 FILLER_24_2848 ();
 sg13g2_fill_2 FILLER_24_2855 ();
 sg13g2_fill_2 FILLER_24_2880 ();
 sg13g2_decap_8 FILLER_24_2918 ();
 sg13g2_decap_8 FILLER_24_2925 ();
 sg13g2_decap_8 FILLER_24_2932 ();
 sg13g2_decap_4 FILLER_24_2939 ();
 sg13g2_decap_8 FILLER_24_2961 ();
 sg13g2_decap_4 FILLER_24_2968 ();
 sg13g2_fill_2 FILLER_24_2972 ();
 sg13g2_decap_8 FILLER_24_3010 ();
 sg13g2_decap_8 FILLER_24_3017 ();
 sg13g2_decap_8 FILLER_24_3024 ();
 sg13g2_decap_4 FILLER_24_3031 ();
 sg13g2_decap_8 FILLER_24_3045 ();
 sg13g2_decap_8 FILLER_24_3052 ();
 sg13g2_decap_8 FILLER_24_3059 ();
 sg13g2_decap_8 FILLER_24_3092 ();
 sg13g2_decap_8 FILLER_24_3099 ();
 sg13g2_decap_8 FILLER_24_3106 ();
 sg13g2_fill_2 FILLER_24_3113 ();
 sg13g2_decap_8 FILLER_24_3151 ();
 sg13g2_decap_8 FILLER_24_3158 ();
 sg13g2_decap_8 FILLER_24_3165 ();
 sg13g2_decap_8 FILLER_24_3172 ();
 sg13g2_fill_2 FILLER_24_3179 ();
 sg13g2_fill_1 FILLER_24_3181 ();
 sg13g2_decap_8 FILLER_24_3228 ();
 sg13g2_decap_8 FILLER_24_3235 ();
 sg13g2_decap_8 FILLER_24_3242 ();
 sg13g2_decap_8 FILLER_24_3249 ();
 sg13g2_decap_8 FILLER_24_3282 ();
 sg13g2_decap_8 FILLER_24_3289 ();
 sg13g2_decap_8 FILLER_24_3296 ();
 sg13g2_decap_8 FILLER_24_3303 ();
 sg13g2_decap_8 FILLER_24_3310 ();
 sg13g2_decap_8 FILLER_24_3317 ();
 sg13g2_decap_8 FILLER_24_3324 ();
 sg13g2_decap_8 FILLER_24_3331 ();
 sg13g2_decap_8 FILLER_24_3338 ();
 sg13g2_decap_8 FILLER_24_3345 ();
 sg13g2_decap_8 FILLER_24_3352 ();
 sg13g2_decap_8 FILLER_24_3359 ();
 sg13g2_decap_8 FILLER_24_3366 ();
 sg13g2_decap_8 FILLER_24_3373 ();
 sg13g2_fill_2 FILLER_24_3380 ();
 sg13g2_decap_8 FILLER_24_3392 ();
 sg13g2_decap_8 FILLER_24_3399 ();
 sg13g2_decap_8 FILLER_24_3406 ();
 sg13g2_decap_8 FILLER_24_3413 ();
 sg13g2_decap_8 FILLER_24_3420 ();
 sg13g2_decap_8 FILLER_24_3427 ();
 sg13g2_decap_8 FILLER_24_3434 ();
 sg13g2_decap_8 FILLER_24_3456 ();
 sg13g2_decap_8 FILLER_24_3463 ();
 sg13g2_decap_4 FILLER_24_3470 ();
 sg13g2_fill_2 FILLER_24_3474 ();
 sg13g2_decap_8 FILLER_24_3507 ();
 sg13g2_decap_8 FILLER_24_3514 ();
 sg13g2_fill_2 FILLER_24_3521 ();
 sg13g2_fill_1 FILLER_24_3523 ();
 sg13g2_decap_8 FILLER_24_3560 ();
 sg13g2_decap_8 FILLER_24_3567 ();
 sg13g2_decap_4 FILLER_24_3574 ();
 sg13g2_fill_2 FILLER_24_3578 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_43 ();
 sg13g2_fill_2 FILLER_25_50 ();
 sg13g2_fill_1 FILLER_25_52 ();
 sg13g2_fill_1 FILLER_25_101 ();
 sg13g2_decap_8 FILLER_25_113 ();
 sg13g2_decap_8 FILLER_25_120 ();
 sg13g2_decap_8 FILLER_25_127 ();
 sg13g2_decap_8 FILLER_25_155 ();
 sg13g2_decap_8 FILLER_25_162 ();
 sg13g2_decap_8 FILLER_25_169 ();
 sg13g2_decap_8 FILLER_25_176 ();
 sg13g2_decap_8 FILLER_25_183 ();
 sg13g2_decap_8 FILLER_25_190 ();
 sg13g2_decap_8 FILLER_25_197 ();
 sg13g2_decap_8 FILLER_25_204 ();
 sg13g2_fill_2 FILLER_25_211 ();
 sg13g2_fill_1 FILLER_25_213 ();
 sg13g2_decap_8 FILLER_25_219 ();
 sg13g2_decap_8 FILLER_25_226 ();
 sg13g2_decap_8 FILLER_25_233 ();
 sg13g2_decap_8 FILLER_25_240 ();
 sg13g2_decap_8 FILLER_25_247 ();
 sg13g2_decap_8 FILLER_25_254 ();
 sg13g2_decap_8 FILLER_25_261 ();
 sg13g2_decap_4 FILLER_25_268 ();
 sg13g2_fill_1 FILLER_25_272 ();
 sg13g2_decap_8 FILLER_25_276 ();
 sg13g2_decap_8 FILLER_25_283 ();
 sg13g2_decap_8 FILLER_25_290 ();
 sg13g2_decap_8 FILLER_25_297 ();
 sg13g2_decap_8 FILLER_25_304 ();
 sg13g2_decap_8 FILLER_25_311 ();
 sg13g2_fill_2 FILLER_25_318 ();
 sg13g2_fill_1 FILLER_25_320 ();
 sg13g2_decap_8 FILLER_25_326 ();
 sg13g2_decap_8 FILLER_25_333 ();
 sg13g2_decap_8 FILLER_25_340 ();
 sg13g2_decap_8 FILLER_25_347 ();
 sg13g2_fill_1 FILLER_25_354 ();
 sg13g2_decap_8 FILLER_25_363 ();
 sg13g2_decap_8 FILLER_25_370 ();
 sg13g2_decap_8 FILLER_25_377 ();
 sg13g2_decap_8 FILLER_25_384 ();
 sg13g2_decap_8 FILLER_25_391 ();
 sg13g2_decap_8 FILLER_25_398 ();
 sg13g2_decap_8 FILLER_25_405 ();
 sg13g2_decap_8 FILLER_25_412 ();
 sg13g2_decap_8 FILLER_25_419 ();
 sg13g2_decap_8 FILLER_25_426 ();
 sg13g2_decap_8 FILLER_25_433 ();
 sg13g2_decap_4 FILLER_25_440 ();
 sg13g2_decap_4 FILLER_25_454 ();
 sg13g2_fill_2 FILLER_25_485 ();
 sg13g2_fill_1 FILLER_25_487 ();
 sg13g2_decap_8 FILLER_25_501 ();
 sg13g2_decap_8 FILLER_25_508 ();
 sg13g2_decap_8 FILLER_25_515 ();
 sg13g2_decap_8 FILLER_25_522 ();
 sg13g2_fill_2 FILLER_25_529 ();
 sg13g2_decap_8 FILLER_25_536 ();
 sg13g2_decap_8 FILLER_25_543 ();
 sg13g2_decap_8 FILLER_25_550 ();
 sg13g2_decap_8 FILLER_25_557 ();
 sg13g2_decap_8 FILLER_25_564 ();
 sg13g2_fill_2 FILLER_25_571 ();
 sg13g2_fill_1 FILLER_25_573 ();
 sg13g2_decap_8 FILLER_25_590 ();
 sg13g2_decap_8 FILLER_25_597 ();
 sg13g2_decap_8 FILLER_25_604 ();
 sg13g2_decap_8 FILLER_25_611 ();
 sg13g2_decap_8 FILLER_25_618 ();
 sg13g2_decap_8 FILLER_25_625 ();
 sg13g2_fill_2 FILLER_25_632 ();
 sg13g2_fill_1 FILLER_25_644 ();
 sg13g2_fill_1 FILLER_25_649 ();
 sg13g2_decap_8 FILLER_25_659 ();
 sg13g2_decap_8 FILLER_25_670 ();
 sg13g2_decap_8 FILLER_25_677 ();
 sg13g2_decap_8 FILLER_25_684 ();
 sg13g2_decap_8 FILLER_25_691 ();
 sg13g2_decap_8 FILLER_25_698 ();
 sg13g2_decap_8 FILLER_25_705 ();
 sg13g2_decap_8 FILLER_25_712 ();
 sg13g2_fill_2 FILLER_25_719 ();
 sg13g2_decap_8 FILLER_25_727 ();
 sg13g2_decap_8 FILLER_25_734 ();
 sg13g2_decap_8 FILLER_25_770 ();
 sg13g2_decap_8 FILLER_25_777 ();
 sg13g2_decap_8 FILLER_25_784 ();
 sg13g2_decap_8 FILLER_25_791 ();
 sg13g2_decap_8 FILLER_25_798 ();
 sg13g2_decap_4 FILLER_25_805 ();
 sg13g2_decap_4 FILLER_25_825 ();
 sg13g2_decap_8 FILLER_25_834 ();
 sg13g2_fill_1 FILLER_25_841 ();
 sg13g2_decap_8 FILLER_25_847 ();
 sg13g2_decap_8 FILLER_25_854 ();
 sg13g2_decap_8 FILLER_25_861 ();
 sg13g2_decap_8 FILLER_25_868 ();
 sg13g2_decap_8 FILLER_25_875 ();
 sg13g2_decap_8 FILLER_25_882 ();
 sg13g2_decap_8 FILLER_25_926 ();
 sg13g2_decap_8 FILLER_25_933 ();
 sg13g2_decap_8 FILLER_25_976 ();
 sg13g2_decap_8 FILLER_25_983 ();
 sg13g2_decap_8 FILLER_25_990 ();
 sg13g2_fill_1 FILLER_25_997 ();
 sg13g2_decap_8 FILLER_25_1004 ();
 sg13g2_decap_8 FILLER_25_1011 ();
 sg13g2_decap_8 FILLER_25_1018 ();
 sg13g2_decap_8 FILLER_25_1025 ();
 sg13g2_decap_8 FILLER_25_1032 ();
 sg13g2_decap_8 FILLER_25_1039 ();
 sg13g2_decap_8 FILLER_25_1046 ();
 sg13g2_decap_8 FILLER_25_1053 ();
 sg13g2_decap_4 FILLER_25_1060 ();
 sg13g2_fill_1 FILLER_25_1064 ();
 sg13g2_fill_1 FILLER_25_1075 ();
 sg13g2_decap_8 FILLER_25_1112 ();
 sg13g2_decap_8 FILLER_25_1119 ();
 sg13g2_decap_8 FILLER_25_1126 ();
 sg13g2_fill_1 FILLER_25_1133 ();
 sg13g2_decap_8 FILLER_25_1145 ();
 sg13g2_decap_8 FILLER_25_1152 ();
 sg13g2_decap_8 FILLER_25_1159 ();
 sg13g2_fill_2 FILLER_25_1166 ();
 sg13g2_decap_8 FILLER_25_1171 ();
 sg13g2_decap_8 FILLER_25_1178 ();
 sg13g2_decap_4 FILLER_25_1185 ();
 sg13g2_fill_1 FILLER_25_1189 ();
 sg13g2_decap_4 FILLER_25_1242 ();
 sg13g2_decap_8 FILLER_25_1256 ();
 sg13g2_decap_8 FILLER_25_1263 ();
 sg13g2_decap_8 FILLER_25_1270 ();
 sg13g2_decap_8 FILLER_25_1277 ();
 sg13g2_decap_8 FILLER_25_1284 ();
 sg13g2_decap_8 FILLER_25_1291 ();
 sg13g2_decap_8 FILLER_25_1298 ();
 sg13g2_decap_8 FILLER_25_1305 ();
 sg13g2_decap_8 FILLER_25_1312 ();
 sg13g2_decap_8 FILLER_25_1319 ();
 sg13g2_decap_8 FILLER_25_1326 ();
 sg13g2_decap_8 FILLER_25_1333 ();
 sg13g2_decap_8 FILLER_25_1340 ();
 sg13g2_decap_8 FILLER_25_1347 ();
 sg13g2_fill_2 FILLER_25_1354 ();
 sg13g2_fill_1 FILLER_25_1356 ();
 sg13g2_fill_2 FILLER_25_1367 ();
 sg13g2_decap_8 FILLER_25_1401 ();
 sg13g2_decap_8 FILLER_25_1408 ();
 sg13g2_decap_8 FILLER_25_1415 ();
 sg13g2_decap_8 FILLER_25_1422 ();
 sg13g2_decap_8 FILLER_25_1429 ();
 sg13g2_decap_8 FILLER_25_1436 ();
 sg13g2_decap_8 FILLER_25_1443 ();
 sg13g2_decap_8 FILLER_25_1450 ();
 sg13g2_decap_8 FILLER_25_1457 ();
 sg13g2_decap_8 FILLER_25_1464 ();
 sg13g2_decap_8 FILLER_25_1471 ();
 sg13g2_decap_8 FILLER_25_1478 ();
 sg13g2_decap_8 FILLER_25_1485 ();
 sg13g2_decap_8 FILLER_25_1492 ();
 sg13g2_decap_8 FILLER_25_1499 ();
 sg13g2_decap_8 FILLER_25_1506 ();
 sg13g2_decap_8 FILLER_25_1513 ();
 sg13g2_fill_1 FILLER_25_1520 ();
 sg13g2_decap_8 FILLER_25_1537 ();
 sg13g2_decap_8 FILLER_25_1544 ();
 sg13g2_fill_1 FILLER_25_1551 ();
 sg13g2_decap_8 FILLER_25_1558 ();
 sg13g2_decap_4 FILLER_25_1565 ();
 sg13g2_fill_2 FILLER_25_1569 ();
 sg13g2_decap_4 FILLER_25_1597 ();
 sg13g2_fill_1 FILLER_25_1605 ();
 sg13g2_decap_8 FILLER_25_1610 ();
 sg13g2_decap_8 FILLER_25_1617 ();
 sg13g2_decap_8 FILLER_25_1624 ();
 sg13g2_decap_8 FILLER_25_1631 ();
 sg13g2_decap_8 FILLER_25_1638 ();
 sg13g2_decap_8 FILLER_25_1645 ();
 sg13g2_decap_8 FILLER_25_1652 ();
 sg13g2_decap_8 FILLER_25_1659 ();
 sg13g2_fill_2 FILLER_25_1666 ();
 sg13g2_fill_1 FILLER_25_1668 ();
 sg13g2_decap_8 FILLER_25_1687 ();
 sg13g2_decap_8 FILLER_25_1694 ();
 sg13g2_fill_2 FILLER_25_1701 ();
 sg13g2_decap_8 FILLER_25_1707 ();
 sg13g2_decap_8 FILLER_25_1714 ();
 sg13g2_decap_8 FILLER_25_1721 ();
 sg13g2_decap_4 FILLER_25_1728 ();
 sg13g2_fill_1 FILLER_25_1732 ();
 sg13g2_decap_8 FILLER_25_1743 ();
 sg13g2_decap_8 FILLER_25_1750 ();
 sg13g2_decap_8 FILLER_25_1757 ();
 sg13g2_decap_8 FILLER_25_1764 ();
 sg13g2_decap_8 FILLER_25_1771 ();
 sg13g2_fill_2 FILLER_25_1778 ();
 sg13g2_decap_4 FILLER_25_1790 ();
 sg13g2_decap_8 FILLER_25_1856 ();
 sg13g2_decap_8 FILLER_25_1863 ();
 sg13g2_decap_8 FILLER_25_1870 ();
 sg13g2_decap_4 FILLER_25_1877 ();
 sg13g2_decap_8 FILLER_25_1912 ();
 sg13g2_decap_8 FILLER_25_1919 ();
 sg13g2_fill_2 FILLER_25_1926 ();
 sg13g2_fill_1 FILLER_25_1928 ();
 sg13g2_decap_8 FILLER_25_1965 ();
 sg13g2_decap_8 FILLER_25_1972 ();
 sg13g2_decap_4 FILLER_25_1979 ();
 sg13g2_fill_2 FILLER_25_1993 ();
 sg13g2_fill_1 FILLER_25_1995 ();
 sg13g2_decap_8 FILLER_25_2009 ();
 sg13g2_decap_8 FILLER_25_2016 ();
 sg13g2_decap_8 FILLER_25_2023 ();
 sg13g2_decap_8 FILLER_25_2030 ();
 sg13g2_decap_8 FILLER_25_2037 ();
 sg13g2_decap_4 FILLER_25_2044 ();
 sg13g2_decap_4 FILLER_25_2070 ();
 sg13g2_fill_1 FILLER_25_2074 ();
 sg13g2_fill_2 FILLER_25_2097 ();
 sg13g2_decap_8 FILLER_25_2105 ();
 sg13g2_decap_8 FILLER_25_2112 ();
 sg13g2_decap_8 FILLER_25_2119 ();
 sg13g2_decap_8 FILLER_25_2126 ();
 sg13g2_decap_8 FILLER_25_2133 ();
 sg13g2_decap_8 FILLER_25_2140 ();
 sg13g2_decap_8 FILLER_25_2147 ();
 sg13g2_decap_4 FILLER_25_2154 ();
 sg13g2_fill_1 FILLER_25_2158 ();
 sg13g2_decap_8 FILLER_25_2165 ();
 sg13g2_decap_8 FILLER_25_2172 ();
 sg13g2_decap_4 FILLER_25_2179 ();
 sg13g2_decap_8 FILLER_25_2188 ();
 sg13g2_decap_4 FILLER_25_2195 ();
 sg13g2_fill_1 FILLER_25_2205 ();
 sg13g2_fill_1 FILLER_25_2216 ();
 sg13g2_decap_8 FILLER_25_2223 ();
 sg13g2_decap_4 FILLER_25_2230 ();
 sg13g2_decap_8 FILLER_25_2240 ();
 sg13g2_fill_2 FILLER_25_2247 ();
 sg13g2_fill_1 FILLER_25_2249 ();
 sg13g2_decap_8 FILLER_25_2256 ();
 sg13g2_decap_8 FILLER_25_2263 ();
 sg13g2_fill_2 FILLER_25_2270 ();
 sg13g2_fill_1 FILLER_25_2272 ();
 sg13g2_decap_8 FILLER_25_2279 ();
 sg13g2_decap_8 FILLER_25_2286 ();
 sg13g2_fill_1 FILLER_25_2293 ();
 sg13g2_decap_4 FILLER_25_2305 ();
 sg13g2_fill_1 FILLER_25_2309 ();
 sg13g2_decap_8 FILLER_25_2325 ();
 sg13g2_decap_8 FILLER_25_2332 ();
 sg13g2_decap_8 FILLER_25_2339 ();
 sg13g2_decap_8 FILLER_25_2346 ();
 sg13g2_fill_2 FILLER_25_2353 ();
 sg13g2_fill_1 FILLER_25_2355 ();
 sg13g2_decap_8 FILLER_25_2382 ();
 sg13g2_decap_8 FILLER_25_2389 ();
 sg13g2_decap_8 FILLER_25_2396 ();
 sg13g2_decap_8 FILLER_25_2403 ();
 sg13g2_fill_1 FILLER_25_2410 ();
 sg13g2_fill_2 FILLER_25_2442 ();
 sg13g2_fill_1 FILLER_25_2444 ();
 sg13g2_decap_8 FILLER_25_2470 ();
 sg13g2_decap_8 FILLER_25_2477 ();
 sg13g2_decap_8 FILLER_25_2484 ();
 sg13g2_decap_8 FILLER_25_2491 ();
 sg13g2_decap_8 FILLER_25_2498 ();
 sg13g2_decap_8 FILLER_25_2523 ();
 sg13g2_decap_8 FILLER_25_2530 ();
 sg13g2_decap_8 FILLER_25_2537 ();
 sg13g2_decap_8 FILLER_25_2544 ();
 sg13g2_fill_2 FILLER_25_2551 ();
 sg13g2_fill_1 FILLER_25_2553 ();
 sg13g2_decap_8 FILLER_25_2580 ();
 sg13g2_decap_8 FILLER_25_2587 ();
 sg13g2_decap_8 FILLER_25_2594 ();
 sg13g2_fill_2 FILLER_25_2601 ();
 sg13g2_decap_8 FILLER_25_2609 ();
 sg13g2_decap_8 FILLER_25_2616 ();
 sg13g2_decap_8 FILLER_25_2623 ();
 sg13g2_decap_8 FILLER_25_2630 ();
 sg13g2_decap_8 FILLER_25_2648 ();
 sg13g2_decap_8 FILLER_25_2655 ();
 sg13g2_decap_8 FILLER_25_2662 ();
 sg13g2_decap_8 FILLER_25_2669 ();
 sg13g2_decap_8 FILLER_25_2676 ();
 sg13g2_decap_4 FILLER_25_2683 ();
 sg13g2_fill_1 FILLER_25_2687 ();
 sg13g2_decap_8 FILLER_25_2703 ();
 sg13g2_decap_8 FILLER_25_2710 ();
 sg13g2_decap_4 FILLER_25_2717 ();
 sg13g2_decap_8 FILLER_25_2727 ();
 sg13g2_fill_1 FILLER_25_2734 ();
 sg13g2_fill_2 FILLER_25_2763 ();
 sg13g2_decap_8 FILLER_25_2785 ();
 sg13g2_decap_8 FILLER_25_2792 ();
 sg13g2_decap_8 FILLER_25_2799 ();
 sg13g2_decap_8 FILLER_25_2806 ();
 sg13g2_decap_8 FILLER_25_2813 ();
 sg13g2_decap_8 FILLER_25_2820 ();
 sg13g2_decap_4 FILLER_25_2827 ();
 sg13g2_fill_2 FILLER_25_2831 ();
 sg13g2_fill_1 FILLER_25_2841 ();
 sg13g2_decap_8 FILLER_25_2852 ();
 sg13g2_decap_8 FILLER_25_2859 ();
 sg13g2_decap_4 FILLER_25_2866 ();
 sg13g2_fill_2 FILLER_25_2870 ();
 sg13g2_decap_4 FILLER_25_2885 ();
 sg13g2_fill_2 FILLER_25_2889 ();
 sg13g2_decap_8 FILLER_25_2917 ();
 sg13g2_decap_8 FILLER_25_2924 ();
 sg13g2_decap_8 FILLER_25_2931 ();
 sg13g2_fill_2 FILLER_25_2938 ();
 sg13g2_decap_8 FILLER_25_2976 ();
 sg13g2_decap_4 FILLER_25_2983 ();
 sg13g2_fill_1 FILLER_25_2987 ();
 sg13g2_decap_8 FILLER_25_3014 ();
 sg13g2_decap_8 FILLER_25_3021 ();
 sg13g2_decap_8 FILLER_25_3028 ();
 sg13g2_fill_1 FILLER_25_3035 ();
 sg13g2_decap_8 FILLER_25_3062 ();
 sg13g2_decap_8 FILLER_25_3069 ();
 sg13g2_decap_8 FILLER_25_3076 ();
 sg13g2_decap_8 FILLER_25_3083 ();
 sg13g2_decap_8 FILLER_25_3090 ();
 sg13g2_decap_8 FILLER_25_3097 ();
 sg13g2_decap_8 FILLER_25_3104 ();
 sg13g2_decap_8 FILLER_25_3111 ();
 sg13g2_decap_8 FILLER_25_3118 ();
 sg13g2_fill_2 FILLER_25_3125 ();
 sg13g2_fill_1 FILLER_25_3127 ();
 sg13g2_decap_8 FILLER_25_3190 ();
 sg13g2_decap_8 FILLER_25_3197 ();
 sg13g2_decap_8 FILLER_25_3204 ();
 sg13g2_fill_2 FILLER_25_3211 ();
 sg13g2_fill_1 FILLER_25_3213 ();
 sg13g2_decap_8 FILLER_25_3220 ();
 sg13g2_decap_8 FILLER_25_3227 ();
 sg13g2_decap_8 FILLER_25_3234 ();
 sg13g2_decap_8 FILLER_25_3241 ();
 sg13g2_decap_8 FILLER_25_3248 ();
 sg13g2_decap_8 FILLER_25_3255 ();
 sg13g2_decap_4 FILLER_25_3262 ();
 sg13g2_fill_1 FILLER_25_3266 ();
 sg13g2_decap_8 FILLER_25_3273 ();
 sg13g2_decap_8 FILLER_25_3280 ();
 sg13g2_decap_8 FILLER_25_3287 ();
 sg13g2_decap_8 FILLER_25_3294 ();
 sg13g2_decap_8 FILLER_25_3301 ();
 sg13g2_decap_8 FILLER_25_3308 ();
 sg13g2_decap_8 FILLER_25_3315 ();
 sg13g2_decap_8 FILLER_25_3322 ();
 sg13g2_decap_8 FILLER_25_3329 ();
 sg13g2_decap_8 FILLER_25_3336 ();
 sg13g2_decap_8 FILLER_25_3343 ();
 sg13g2_decap_8 FILLER_25_3350 ();
 sg13g2_fill_2 FILLER_25_3357 ();
 sg13g2_fill_1 FILLER_25_3359 ();
 sg13g2_decap_8 FILLER_25_3386 ();
 sg13g2_decap_8 FILLER_25_3393 ();
 sg13g2_decap_8 FILLER_25_3400 ();
 sg13g2_decap_8 FILLER_25_3407 ();
 sg13g2_decap_8 FILLER_25_3414 ();
 sg13g2_decap_8 FILLER_25_3421 ();
 sg13g2_fill_2 FILLER_25_3428 ();
 sg13g2_fill_1 FILLER_25_3430 ();
 sg13g2_decap_8 FILLER_25_3466 ();
 sg13g2_fill_1 FILLER_25_3473 ();
 sg13g2_fill_2 FILLER_25_3484 ();
 sg13g2_decap_8 FILLER_25_3508 ();
 sg13g2_decap_8 FILLER_25_3515 ();
 sg13g2_fill_2 FILLER_25_3522 ();
 sg13g2_fill_1 FILLER_25_3524 ();
 sg13g2_fill_2 FILLER_25_3535 ();
 sg13g2_decap_8 FILLER_25_3568 ();
 sg13g2_decap_4 FILLER_25_3575 ();
 sg13g2_fill_1 FILLER_25_3579 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_fill_2 FILLER_26_7 ();
 sg13g2_fill_1 FILLER_26_9 ();
 sg13g2_decap_8 FILLER_26_41 ();
 sg13g2_decap_8 FILLER_26_48 ();
 sg13g2_decap_8 FILLER_26_55 ();
 sg13g2_decap_8 FILLER_26_62 ();
 sg13g2_decap_8 FILLER_26_69 ();
 sg13g2_fill_2 FILLER_26_76 ();
 sg13g2_fill_1 FILLER_26_78 ();
 sg13g2_fill_2 FILLER_26_88 ();
 sg13g2_decap_8 FILLER_26_94 ();
 sg13g2_fill_1 FILLER_26_101 ();
 sg13g2_decap_8 FILLER_26_105 ();
 sg13g2_decap_8 FILLER_26_112 ();
 sg13g2_decap_8 FILLER_26_119 ();
 sg13g2_fill_1 FILLER_26_126 ();
 sg13g2_decap_8 FILLER_26_159 ();
 sg13g2_decap_8 FILLER_26_166 ();
 sg13g2_decap_8 FILLER_26_173 ();
 sg13g2_decap_8 FILLER_26_180 ();
 sg13g2_fill_2 FILLER_26_187 ();
 sg13g2_decap_8 FILLER_26_201 ();
 sg13g2_decap_8 FILLER_26_208 ();
 sg13g2_decap_8 FILLER_26_215 ();
 sg13g2_decap_4 FILLER_26_222 ();
 sg13g2_decap_8 FILLER_26_231 ();
 sg13g2_decap_8 FILLER_26_238 ();
 sg13g2_decap_8 FILLER_26_245 ();
 sg13g2_decap_8 FILLER_26_252 ();
 sg13g2_decap_8 FILLER_26_259 ();
 sg13g2_fill_2 FILLER_26_266 ();
 sg13g2_decap_8 FILLER_26_272 ();
 sg13g2_decap_8 FILLER_26_279 ();
 sg13g2_decap_8 FILLER_26_286 ();
 sg13g2_decap_8 FILLER_26_293 ();
 sg13g2_fill_2 FILLER_26_300 ();
 sg13g2_fill_1 FILLER_26_302 ();
 sg13g2_decap_8 FILLER_26_313 ();
 sg13g2_decap_8 FILLER_26_320 ();
 sg13g2_decap_8 FILLER_26_327 ();
 sg13g2_decap_8 FILLER_26_334 ();
 sg13g2_decap_8 FILLER_26_341 ();
 sg13g2_decap_8 FILLER_26_348 ();
 sg13g2_fill_2 FILLER_26_355 ();
 sg13g2_fill_2 FILLER_26_369 ();
 sg13g2_fill_1 FILLER_26_371 ();
 sg13g2_fill_2 FILLER_26_377 ();
 sg13g2_fill_1 FILLER_26_384 ();
 sg13g2_fill_1 FILLER_26_398 ();
 sg13g2_decap_4 FILLER_26_431 ();
 sg13g2_fill_2 FILLER_26_441 ();
 sg13g2_decap_8 FILLER_26_448 ();
 sg13g2_decap_4 FILLER_26_455 ();
 sg13g2_fill_1 FILLER_26_459 ();
 sg13g2_fill_2 FILLER_26_465 ();
 sg13g2_fill_2 FILLER_26_484 ();
 sg13g2_fill_1 FILLER_26_486 ();
 sg13g2_decap_8 FILLER_26_500 ();
 sg13g2_decap_4 FILLER_26_507 ();
 sg13g2_fill_1 FILLER_26_511 ();
 sg13g2_decap_8 FILLER_26_518 ();
 sg13g2_fill_1 FILLER_26_525 ();
 sg13g2_fill_1 FILLER_26_531 ();
 sg13g2_decap_8 FILLER_26_553 ();
 sg13g2_decap_8 FILLER_26_560 ();
 sg13g2_decap_8 FILLER_26_567 ();
 sg13g2_fill_2 FILLER_26_574 ();
 sg13g2_fill_1 FILLER_26_576 ();
 sg13g2_decap_8 FILLER_26_580 ();
 sg13g2_decap_8 FILLER_26_587 ();
 sg13g2_decap_8 FILLER_26_594 ();
 sg13g2_decap_8 FILLER_26_601 ();
 sg13g2_decap_8 FILLER_26_608 ();
 sg13g2_decap_8 FILLER_26_615 ();
 sg13g2_decap_8 FILLER_26_622 ();
 sg13g2_decap_4 FILLER_26_629 ();
 sg13g2_fill_1 FILLER_26_633 ();
 sg13g2_decap_8 FILLER_26_672 ();
 sg13g2_decap_8 FILLER_26_679 ();
 sg13g2_decap_8 FILLER_26_686 ();
 sg13g2_decap_8 FILLER_26_693 ();
 sg13g2_decap_8 FILLER_26_700 ();
 sg13g2_decap_8 FILLER_26_707 ();
 sg13g2_decap_8 FILLER_26_714 ();
 sg13g2_decap_4 FILLER_26_724 ();
 sg13g2_decap_8 FILLER_26_780 ();
 sg13g2_decap_8 FILLER_26_787 ();
 sg13g2_decap_8 FILLER_26_794 ();
 sg13g2_fill_1 FILLER_26_801 ();
 sg13g2_decap_8 FILLER_26_807 ();
 sg13g2_decap_8 FILLER_26_814 ();
 sg13g2_decap_8 FILLER_26_821 ();
 sg13g2_decap_8 FILLER_26_828 ();
 sg13g2_decap_8 FILLER_26_835 ();
 sg13g2_decap_8 FILLER_26_842 ();
 sg13g2_decap_8 FILLER_26_849 ();
 sg13g2_decap_8 FILLER_26_856 ();
 sg13g2_decap_8 FILLER_26_863 ();
 sg13g2_decap_4 FILLER_26_870 ();
 sg13g2_decap_8 FILLER_26_890 ();
 sg13g2_decap_8 FILLER_26_897 ();
 sg13g2_decap_4 FILLER_26_904 ();
 sg13g2_decap_8 FILLER_26_913 ();
 sg13g2_decap_8 FILLER_26_920 ();
 sg13g2_decap_8 FILLER_26_927 ();
 sg13g2_decap_8 FILLER_26_934 ();
 sg13g2_decap_8 FILLER_26_941 ();
 sg13g2_decap_8 FILLER_26_948 ();
 sg13g2_decap_8 FILLER_26_955 ();
 sg13g2_decap_8 FILLER_26_962 ();
 sg13g2_decap_8 FILLER_26_969 ();
 sg13g2_decap_8 FILLER_26_976 ();
 sg13g2_decap_8 FILLER_26_983 ();
 sg13g2_fill_2 FILLER_26_1006 ();
 sg13g2_fill_1 FILLER_26_1026 ();
 sg13g2_decap_8 FILLER_26_1053 ();
 sg13g2_fill_2 FILLER_26_1071 ();
 sg13g2_fill_1 FILLER_26_1073 ();
 sg13g2_decap_8 FILLER_26_1100 ();
 sg13g2_decap_8 FILLER_26_1107 ();
 sg13g2_fill_2 FILLER_26_1114 ();
 sg13g2_decap_8 FILLER_26_1121 ();
 sg13g2_fill_2 FILLER_26_1128 ();
 sg13g2_fill_1 FILLER_26_1130 ();
 sg13g2_decap_8 FILLER_26_1145 ();
 sg13g2_decap_8 FILLER_26_1162 ();
 sg13g2_decap_8 FILLER_26_1169 ();
 sg13g2_fill_2 FILLER_26_1176 ();
 sg13g2_decap_8 FILLER_26_1188 ();
 sg13g2_decap_4 FILLER_26_1195 ();
 sg13g2_fill_1 FILLER_26_1199 ();
 sg13g2_decap_8 FILLER_26_1231 ();
 sg13g2_fill_2 FILLER_26_1238 ();
 sg13g2_fill_1 FILLER_26_1240 ();
 sg13g2_decap_8 FILLER_26_1289 ();
 sg13g2_decap_8 FILLER_26_1296 ();
 sg13g2_decap_8 FILLER_26_1303 ();
 sg13g2_decap_8 FILLER_26_1310 ();
 sg13g2_decap_8 FILLER_26_1317 ();
 sg13g2_decap_8 FILLER_26_1324 ();
 sg13g2_fill_2 FILLER_26_1331 ();
 sg13g2_fill_2 FILLER_26_1343 ();
 sg13g2_decap_8 FILLER_26_1371 ();
 sg13g2_decap_8 FILLER_26_1378 ();
 sg13g2_decap_8 FILLER_26_1385 ();
 sg13g2_decap_8 FILLER_26_1392 ();
 sg13g2_decap_8 FILLER_26_1412 ();
 sg13g2_fill_1 FILLER_26_1419 ();
 sg13g2_decap_4 FILLER_26_1456 ();
 sg13g2_fill_1 FILLER_26_1460 ();
 sg13g2_decap_8 FILLER_26_1465 ();
 sg13g2_decap_8 FILLER_26_1472 ();
 sg13g2_decap_8 FILLER_26_1479 ();
 sg13g2_decap_8 FILLER_26_1486 ();
 sg13g2_decap_8 FILLER_26_1493 ();
 sg13g2_decap_8 FILLER_26_1500 ();
 sg13g2_decap_8 FILLER_26_1507 ();
 sg13g2_fill_2 FILLER_26_1514 ();
 sg13g2_fill_1 FILLER_26_1516 ();
 sg13g2_decap_8 FILLER_26_1543 ();
 sg13g2_decap_8 FILLER_26_1550 ();
 sg13g2_decap_8 FILLER_26_1557 ();
 sg13g2_decap_8 FILLER_26_1564 ();
 sg13g2_decap_8 FILLER_26_1571 ();
 sg13g2_decap_4 FILLER_26_1586 ();
 sg13g2_decap_8 FILLER_26_1626 ();
 sg13g2_decap_8 FILLER_26_1633 ();
 sg13g2_decap_8 FILLER_26_1640 ();
 sg13g2_decap_8 FILLER_26_1647 ();
 sg13g2_decap_8 FILLER_26_1654 ();
 sg13g2_decap_8 FILLER_26_1661 ();
 sg13g2_decap_8 FILLER_26_1668 ();
 sg13g2_decap_8 FILLER_26_1675 ();
 sg13g2_decap_8 FILLER_26_1682 ();
 sg13g2_decap_8 FILLER_26_1689 ();
 sg13g2_decap_8 FILLER_26_1696 ();
 sg13g2_decap_8 FILLER_26_1703 ();
 sg13g2_decap_8 FILLER_26_1710 ();
 sg13g2_decap_8 FILLER_26_1717 ();
 sg13g2_decap_8 FILLER_26_1724 ();
 sg13g2_decap_8 FILLER_26_1731 ();
 sg13g2_decap_8 FILLER_26_1738 ();
 sg13g2_decap_8 FILLER_26_1745 ();
 sg13g2_decap_8 FILLER_26_1752 ();
 sg13g2_decap_8 FILLER_26_1759 ();
 sg13g2_decap_8 FILLER_26_1766 ();
 sg13g2_decap_8 FILLER_26_1773 ();
 sg13g2_decap_8 FILLER_26_1780 ();
 sg13g2_decap_8 FILLER_26_1787 ();
 sg13g2_decap_8 FILLER_26_1794 ();
 sg13g2_decap_8 FILLER_26_1801 ();
 sg13g2_decap_8 FILLER_26_1808 ();
 sg13g2_decap_8 FILLER_26_1815 ();
 sg13g2_decap_8 FILLER_26_1822 ();
 sg13g2_decap_8 FILLER_26_1829 ();
 sg13g2_decap_8 FILLER_26_1836 ();
 sg13g2_fill_1 FILLER_26_1843 ();
 sg13g2_decap_8 FILLER_26_1854 ();
 sg13g2_decap_8 FILLER_26_1861 ();
 sg13g2_decap_8 FILLER_26_1868 ();
 sg13g2_decap_8 FILLER_26_1875 ();
 sg13g2_decap_4 FILLER_26_1882 ();
 sg13g2_fill_2 FILLER_26_1886 ();
 sg13g2_decap_8 FILLER_26_1908 ();
 sg13g2_decap_8 FILLER_26_1915 ();
 sg13g2_decap_8 FILLER_26_1922 ();
 sg13g2_decap_8 FILLER_26_1929 ();
 sg13g2_decap_4 FILLER_26_1936 ();
 sg13g2_decap_8 FILLER_26_1966 ();
 sg13g2_decap_8 FILLER_26_1973 ();
 sg13g2_fill_1 FILLER_26_1980 ();
 sg13g2_decap_8 FILLER_26_2011 ();
 sg13g2_decap_8 FILLER_26_2018 ();
 sg13g2_decap_8 FILLER_26_2025 ();
 sg13g2_decap_4 FILLER_26_2032 ();
 sg13g2_fill_1 FILLER_26_2036 ();
 sg13g2_fill_1 FILLER_26_2050 ();
 sg13g2_decap_8 FILLER_26_2066 ();
 sg13g2_decap_8 FILLER_26_2073 ();
 sg13g2_decap_8 FILLER_26_2080 ();
 sg13g2_decap_4 FILLER_26_2087 ();
 sg13g2_fill_1 FILLER_26_2091 ();
 sg13g2_decap_8 FILLER_26_2096 ();
 sg13g2_decap_8 FILLER_26_2103 ();
 sg13g2_decap_8 FILLER_26_2110 ();
 sg13g2_decap_8 FILLER_26_2117 ();
 sg13g2_decap_8 FILLER_26_2124 ();
 sg13g2_decap_8 FILLER_26_2131 ();
 sg13g2_decap_8 FILLER_26_2138 ();
 sg13g2_decap_8 FILLER_26_2145 ();
 sg13g2_decap_8 FILLER_26_2152 ();
 sg13g2_decap_8 FILLER_26_2159 ();
 sg13g2_decap_8 FILLER_26_2166 ();
 sg13g2_decap_8 FILLER_26_2173 ();
 sg13g2_decap_8 FILLER_26_2180 ();
 sg13g2_fill_1 FILLER_26_2187 ();
 sg13g2_fill_2 FILLER_26_2216 ();
 sg13g2_fill_1 FILLER_26_2218 ();
 sg13g2_fill_2 FILLER_26_2237 ();
 sg13g2_decap_8 FILLER_26_2249 ();
 sg13g2_decap_8 FILLER_26_2256 ();
 sg13g2_decap_8 FILLER_26_2263 ();
 sg13g2_decap_8 FILLER_26_2270 ();
 sg13g2_fill_1 FILLER_26_2277 ();
 sg13g2_decap_8 FILLER_26_2284 ();
 sg13g2_fill_2 FILLER_26_2291 ();
 sg13g2_fill_1 FILLER_26_2293 ();
 sg13g2_decap_4 FILLER_26_2300 ();
 sg13g2_decap_4 FILLER_26_2313 ();
 sg13g2_decap_8 FILLER_26_2330 ();
 sg13g2_decap_8 FILLER_26_2337 ();
 sg13g2_fill_2 FILLER_26_2344 ();
 sg13g2_fill_1 FILLER_26_2346 ();
 sg13g2_decap_8 FILLER_26_2383 ();
 sg13g2_decap_8 FILLER_26_2390 ();
 sg13g2_decap_8 FILLER_26_2397 ();
 sg13g2_fill_1 FILLER_26_2404 ();
 sg13g2_decap_8 FILLER_26_2438 ();
 sg13g2_decap_8 FILLER_26_2445 ();
 sg13g2_decap_8 FILLER_26_2452 ();
 sg13g2_decap_8 FILLER_26_2459 ();
 sg13g2_decap_8 FILLER_26_2466 ();
 sg13g2_decap_8 FILLER_26_2473 ();
 sg13g2_decap_8 FILLER_26_2480 ();
 sg13g2_fill_1 FILLER_26_2487 ();
 sg13g2_decap_8 FILLER_26_2514 ();
 sg13g2_decap_8 FILLER_26_2521 ();
 sg13g2_decap_8 FILLER_26_2528 ();
 sg13g2_decap_8 FILLER_26_2535 ();
 sg13g2_decap_8 FILLER_26_2542 ();
 sg13g2_decap_4 FILLER_26_2549 ();
 sg13g2_fill_2 FILLER_26_2553 ();
 sg13g2_decap_8 FILLER_26_2565 ();
 sg13g2_decap_8 FILLER_26_2572 ();
 sg13g2_decap_8 FILLER_26_2579 ();
 sg13g2_decap_8 FILLER_26_2586 ();
 sg13g2_decap_8 FILLER_26_2593 ();
 sg13g2_fill_1 FILLER_26_2600 ();
 sg13g2_decap_8 FILLER_26_2637 ();
 sg13g2_decap_8 FILLER_26_2644 ();
 sg13g2_decap_8 FILLER_26_2651 ();
 sg13g2_decap_8 FILLER_26_2661 ();
 sg13g2_decap_8 FILLER_26_2668 ();
 sg13g2_decap_8 FILLER_26_2675 ();
 sg13g2_decap_4 FILLER_26_2682 ();
 sg13g2_fill_2 FILLER_26_2686 ();
 sg13g2_decap_8 FILLER_26_2714 ();
 sg13g2_decap_8 FILLER_26_2721 ();
 sg13g2_decap_8 FILLER_26_2728 ();
 sg13g2_decap_8 FILLER_26_2735 ();
 sg13g2_fill_2 FILLER_26_2742 ();
 sg13g2_decap_8 FILLER_26_2755 ();
 sg13g2_decap_8 FILLER_26_2762 ();
 sg13g2_decap_8 FILLER_26_2769 ();
 sg13g2_decap_8 FILLER_26_2776 ();
 sg13g2_decap_8 FILLER_26_2783 ();
 sg13g2_decap_4 FILLER_26_2790 ();
 sg13g2_fill_2 FILLER_26_2794 ();
 sg13g2_decap_8 FILLER_26_2802 ();
 sg13g2_decap_8 FILLER_26_2834 ();
 sg13g2_decap_4 FILLER_26_2841 ();
 sg13g2_fill_1 FILLER_26_2845 ();
 sg13g2_decap_8 FILLER_26_2852 ();
 sg13g2_decap_8 FILLER_26_2885 ();
 sg13g2_decap_8 FILLER_26_2892 ();
 sg13g2_fill_2 FILLER_26_2899 ();
 sg13g2_decap_8 FILLER_26_2912 ();
 sg13g2_decap_4 FILLER_26_2919 ();
 sg13g2_fill_2 FILLER_26_2923 ();
 sg13g2_fill_2 FILLER_26_2933 ();
 sg13g2_decap_8 FILLER_26_2940 ();
 sg13g2_decap_8 FILLER_26_2947 ();
 sg13g2_decap_8 FILLER_26_2954 ();
 sg13g2_decap_8 FILLER_26_2961 ();
 sg13g2_decap_8 FILLER_26_2968 ();
 sg13g2_decap_8 FILLER_26_2975 ();
 sg13g2_fill_1 FILLER_26_2992 ();
 sg13g2_decap_8 FILLER_26_3001 ();
 sg13g2_decap_8 FILLER_26_3008 ();
 sg13g2_decap_8 FILLER_26_3015 ();
 sg13g2_decap_8 FILLER_26_3022 ();
 sg13g2_decap_8 FILLER_26_3029 ();
 sg13g2_decap_8 FILLER_26_3068 ();
 sg13g2_decap_8 FILLER_26_3075 ();
 sg13g2_decap_4 FILLER_26_3082 ();
 sg13g2_fill_2 FILLER_26_3086 ();
 sg13g2_decap_8 FILLER_26_3099 ();
 sg13g2_decap_8 FILLER_26_3106 ();
 sg13g2_decap_8 FILLER_26_3113 ();
 sg13g2_decap_8 FILLER_26_3120 ();
 sg13g2_decap_8 FILLER_26_3127 ();
 sg13g2_decap_8 FILLER_26_3134 ();
 sg13g2_fill_2 FILLER_26_3141 ();
 sg13g2_fill_1 FILLER_26_3143 ();
 sg13g2_decap_8 FILLER_26_3147 ();
 sg13g2_decap_8 FILLER_26_3154 ();
 sg13g2_decap_8 FILLER_26_3161 ();
 sg13g2_decap_8 FILLER_26_3168 ();
 sg13g2_decap_8 FILLER_26_3175 ();
 sg13g2_decap_8 FILLER_26_3182 ();
 sg13g2_decap_8 FILLER_26_3189 ();
 sg13g2_decap_4 FILLER_26_3196 ();
 sg13g2_fill_2 FILLER_26_3200 ();
 sg13g2_decap_8 FILLER_26_3208 ();
 sg13g2_decap_8 FILLER_26_3215 ();
 sg13g2_decap_8 FILLER_26_3222 ();
 sg13g2_fill_2 FILLER_26_3229 ();
 sg13g2_fill_1 FILLER_26_3231 ();
 sg13g2_decap_8 FILLER_26_3242 ();
 sg13g2_decap_8 FILLER_26_3249 ();
 sg13g2_decap_8 FILLER_26_3256 ();
 sg13g2_decap_8 FILLER_26_3263 ();
 sg13g2_decap_8 FILLER_26_3270 ();
 sg13g2_decap_8 FILLER_26_3277 ();
 sg13g2_decap_8 FILLER_26_3284 ();
 sg13g2_decap_4 FILLER_26_3291 ();
 sg13g2_fill_1 FILLER_26_3295 ();
 sg13g2_fill_2 FILLER_26_3322 ();
 sg13g2_decap_8 FILLER_26_3334 ();
 sg13g2_fill_2 FILLER_26_3341 ();
 sg13g2_decap_8 FILLER_26_3353 ();
 sg13g2_decap_8 FILLER_26_3360 ();
 sg13g2_decap_8 FILLER_26_3367 ();
 sg13g2_decap_8 FILLER_26_3374 ();
 sg13g2_decap_4 FILLER_26_3381 ();
 sg13g2_decap_8 FILLER_26_3398 ();
 sg13g2_decap_8 FILLER_26_3405 ();
 sg13g2_decap_8 FILLER_26_3412 ();
 sg13g2_decap_8 FILLER_26_3422 ();
 sg13g2_fill_2 FILLER_26_3429 ();
 sg13g2_decap_8 FILLER_26_3462 ();
 sg13g2_decap_8 FILLER_26_3469 ();
 sg13g2_decap_8 FILLER_26_3476 ();
 sg13g2_decap_8 FILLER_26_3483 ();
 sg13g2_decap_8 FILLER_26_3503 ();
 sg13g2_decap_8 FILLER_26_3510 ();
 sg13g2_decap_8 FILLER_26_3517 ();
 sg13g2_decap_8 FILLER_26_3524 ();
 sg13g2_decap_4 FILLER_26_3531 ();
 sg13g2_decap_4 FILLER_26_3539 ();
 sg13g2_fill_2 FILLER_26_3543 ();
 sg13g2_decap_8 FILLER_26_3553 ();
 sg13g2_decap_8 FILLER_26_3560 ();
 sg13g2_decap_8 FILLER_26_3567 ();
 sg13g2_decap_4 FILLER_26_3574 ();
 sg13g2_fill_2 FILLER_26_3578 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_4 FILLER_27_7 ();
 sg13g2_fill_2 FILLER_27_11 ();
 sg13g2_fill_1 FILLER_27_32 ();
 sg13g2_decap_8 FILLER_27_51 ();
 sg13g2_decap_8 FILLER_27_58 ();
 sg13g2_decap_8 FILLER_27_65 ();
 sg13g2_decap_8 FILLER_27_72 ();
 sg13g2_decap_8 FILLER_27_79 ();
 sg13g2_decap_8 FILLER_27_86 ();
 sg13g2_decap_4 FILLER_27_93 ();
 sg13g2_decap_8 FILLER_27_101 ();
 sg13g2_decap_8 FILLER_27_108 ();
 sg13g2_decap_4 FILLER_27_115 ();
 sg13g2_fill_2 FILLER_27_119 ();
 sg13g2_decap_8 FILLER_27_169 ();
 sg13g2_fill_2 FILLER_27_176 ();
 sg13g2_decap_4 FILLER_27_209 ();
 sg13g2_fill_1 FILLER_27_213 ();
 sg13g2_decap_8 FILLER_27_243 ();
 sg13g2_decap_8 FILLER_27_250 ();
 sg13g2_fill_2 FILLER_27_261 ();
 sg13g2_fill_2 FILLER_27_268 ();
 sg13g2_decap_8 FILLER_27_287 ();
 sg13g2_fill_2 FILLER_27_294 ();
 sg13g2_fill_1 FILLER_27_296 ();
 sg13g2_fill_2 FILLER_27_313 ();
 sg13g2_fill_1 FILLER_27_315 ();
 sg13g2_fill_1 FILLER_27_321 ();
 sg13g2_decap_8 FILLER_27_335 ();
 sg13g2_decap_8 FILLER_27_342 ();
 sg13g2_decap_8 FILLER_27_349 ();
 sg13g2_decap_8 FILLER_27_356 ();
 sg13g2_decap_4 FILLER_27_363 ();
 sg13g2_fill_2 FILLER_27_367 ();
 sg13g2_decap_8 FILLER_27_383 ();
 sg13g2_decap_8 FILLER_27_390 ();
 sg13g2_decap_8 FILLER_27_397 ();
 sg13g2_decap_8 FILLER_27_404 ();
 sg13g2_decap_4 FILLER_27_411 ();
 sg13g2_fill_1 FILLER_27_415 ();
 sg13g2_decap_8 FILLER_27_449 ();
 sg13g2_decap_8 FILLER_27_456 ();
 sg13g2_decap_8 FILLER_27_463 ();
 sg13g2_decap_8 FILLER_27_470 ();
 sg13g2_fill_2 FILLER_27_477 ();
 sg13g2_fill_1 FILLER_27_479 ();
 sg13g2_decap_8 FILLER_27_485 ();
 sg13g2_decap_8 FILLER_27_492 ();
 sg13g2_decap_8 FILLER_27_499 ();
 sg13g2_decap_4 FILLER_27_506 ();
 sg13g2_decap_4 FILLER_27_518 ();
 sg13g2_fill_1 FILLER_27_522 ();
 sg13g2_decap_8 FILLER_27_543 ();
 sg13g2_decap_8 FILLER_27_550 ();
 sg13g2_decap_8 FILLER_27_557 ();
 sg13g2_decap_8 FILLER_27_564 ();
 sg13g2_fill_2 FILLER_27_571 ();
 sg13g2_fill_1 FILLER_27_573 ();
 sg13g2_fill_1 FILLER_27_582 ();
 sg13g2_decap_4 FILLER_27_597 ();
 sg13g2_fill_1 FILLER_27_601 ();
 sg13g2_decap_8 FILLER_27_610 ();
 sg13g2_decap_4 FILLER_27_617 ();
 sg13g2_fill_1 FILLER_27_621 ();
 sg13g2_decap_4 FILLER_27_627 ();
 sg13g2_decap_8 FILLER_27_639 ();
 sg13g2_decap_8 FILLER_27_646 ();
 sg13g2_fill_2 FILLER_27_653 ();
 sg13g2_fill_1 FILLER_27_655 ();
 sg13g2_decap_8 FILLER_27_659 ();
 sg13g2_decap_8 FILLER_27_666 ();
 sg13g2_decap_4 FILLER_27_673 ();
 sg13g2_fill_1 FILLER_27_677 ();
 sg13g2_decap_4 FILLER_27_686 ();
 sg13g2_fill_1 FILLER_27_690 ();
 sg13g2_decap_4 FILLER_27_699 ();
 sg13g2_decap_8 FILLER_27_709 ();
 sg13g2_decap_8 FILLER_27_716 ();
 sg13g2_decap_8 FILLER_27_723 ();
 sg13g2_fill_1 FILLER_27_730 ();
 sg13g2_fill_1 FILLER_27_744 ();
 sg13g2_decap_8 FILLER_27_771 ();
 sg13g2_decap_8 FILLER_27_778 ();
 sg13g2_decap_4 FILLER_27_785 ();
 sg13g2_fill_1 FILLER_27_789 ();
 sg13g2_fill_2 FILLER_27_816 ();
 sg13g2_decap_8 FILLER_27_826 ();
 sg13g2_decap_8 FILLER_27_833 ();
 sg13g2_decap_8 FILLER_27_840 ();
 sg13g2_decap_8 FILLER_27_847 ();
 sg13g2_decap_8 FILLER_27_854 ();
 sg13g2_fill_2 FILLER_27_861 ();
 sg13g2_fill_1 FILLER_27_863 ();
 sg13g2_decap_8 FILLER_27_874 ();
 sg13g2_decap_8 FILLER_27_881 ();
 sg13g2_decap_8 FILLER_27_888 ();
 sg13g2_decap_8 FILLER_27_895 ();
 sg13g2_decap_8 FILLER_27_902 ();
 sg13g2_decap_4 FILLER_27_909 ();
 sg13g2_decap_8 FILLER_27_918 ();
 sg13g2_decap_4 FILLER_27_925 ();
 sg13g2_decap_8 FILLER_27_934 ();
 sg13g2_decap_8 FILLER_27_941 ();
 sg13g2_decap_8 FILLER_27_948 ();
 sg13g2_decap_8 FILLER_27_955 ();
 sg13g2_decap_8 FILLER_27_962 ();
 sg13g2_decap_8 FILLER_27_969 ();
 sg13g2_decap_8 FILLER_27_976 ();
 sg13g2_decap_8 FILLER_27_993 ();
 sg13g2_decap_8 FILLER_27_1000 ();
 sg13g2_decap_8 FILLER_27_1007 ();
 sg13g2_decap_8 FILLER_27_1014 ();
 sg13g2_decap_8 FILLER_27_1021 ();
 sg13g2_decap_8 FILLER_27_1028 ();
 sg13g2_decap_8 FILLER_27_1035 ();
 sg13g2_decap_8 FILLER_27_1042 ();
 sg13g2_decap_8 FILLER_27_1049 ();
 sg13g2_decap_8 FILLER_27_1056 ();
 sg13g2_decap_8 FILLER_27_1063 ();
 sg13g2_decap_8 FILLER_27_1070 ();
 sg13g2_decap_8 FILLER_27_1077 ();
 sg13g2_decap_8 FILLER_27_1084 ();
 sg13g2_decap_8 FILLER_27_1091 ();
 sg13g2_decap_8 FILLER_27_1098 ();
 sg13g2_decap_8 FILLER_27_1110 ();
 sg13g2_decap_8 FILLER_27_1117 ();
 sg13g2_decap_8 FILLER_27_1124 ();
 sg13g2_fill_2 FILLER_27_1131 ();
 sg13g2_fill_1 FILLER_27_1133 ();
 sg13g2_fill_2 FILLER_27_1137 ();
 sg13g2_fill_1 FILLER_27_1151 ();
 sg13g2_decap_8 FILLER_27_1178 ();
 sg13g2_decap_4 FILLER_27_1185 ();
 sg13g2_fill_2 FILLER_27_1189 ();
 sg13g2_decap_4 FILLER_27_1199 ();
 sg13g2_fill_2 FILLER_27_1203 ();
 sg13g2_decap_8 FILLER_27_1210 ();
 sg13g2_decap_8 FILLER_27_1217 ();
 sg13g2_decap_8 FILLER_27_1224 ();
 sg13g2_decap_8 FILLER_27_1231 ();
 sg13g2_decap_8 FILLER_27_1238 ();
 sg13g2_decap_8 FILLER_27_1245 ();
 sg13g2_decap_8 FILLER_27_1252 ();
 sg13g2_decap_8 FILLER_27_1259 ();
 sg13g2_decap_8 FILLER_27_1266 ();
 sg13g2_fill_1 FILLER_27_1273 ();
 sg13g2_fill_2 FILLER_27_1288 ();
 sg13g2_decap_8 FILLER_27_1326 ();
 sg13g2_decap_8 FILLER_27_1333 ();
 sg13g2_decap_8 FILLER_27_1340 ();
 sg13g2_decap_4 FILLER_27_1347 ();
 sg13g2_fill_1 FILLER_27_1351 ();
 sg13g2_decap_8 FILLER_27_1377 ();
 sg13g2_decap_8 FILLER_27_1384 ();
 sg13g2_decap_8 FILLER_27_1391 ();
 sg13g2_decap_8 FILLER_27_1398 ();
 sg13g2_fill_2 FILLER_27_1405 ();
 sg13g2_decap_8 FILLER_27_1427 ();
 sg13g2_decap_4 FILLER_27_1434 ();
 sg13g2_fill_1 FILLER_27_1438 ();
 sg13g2_fill_2 FILLER_27_1476 ();
 sg13g2_decap_8 FILLER_27_1491 ();
 sg13g2_decap_8 FILLER_27_1498 ();
 sg13g2_fill_2 FILLER_27_1505 ();
 sg13g2_decap_8 FILLER_27_1515 ();
 sg13g2_decap_8 FILLER_27_1522 ();
 sg13g2_decap_8 FILLER_27_1529 ();
 sg13g2_decap_4 FILLER_27_1536 ();
 sg13g2_decap_8 FILLER_27_1589 ();
 sg13g2_decap_8 FILLER_27_1596 ();
 sg13g2_decap_8 FILLER_27_1603 ();
 sg13g2_decap_8 FILLER_27_1610 ();
 sg13g2_decap_4 FILLER_27_1617 ();
 sg13g2_fill_1 FILLER_27_1621 ();
 sg13g2_decap_8 FILLER_27_1630 ();
 sg13g2_decap_8 FILLER_27_1637 ();
 sg13g2_fill_2 FILLER_27_1644 ();
 sg13g2_fill_1 FILLER_27_1646 ();
 sg13g2_decap_8 FILLER_27_1665 ();
 sg13g2_decap_8 FILLER_27_1672 ();
 sg13g2_decap_8 FILLER_27_1679 ();
 sg13g2_decap_8 FILLER_27_1686 ();
 sg13g2_decap_8 FILLER_27_1693 ();
 sg13g2_decap_8 FILLER_27_1726 ();
 sg13g2_decap_8 FILLER_27_1733 ();
 sg13g2_decap_4 FILLER_27_1740 ();
 sg13g2_decap_8 FILLER_27_1764 ();
 sg13g2_decap_8 FILLER_27_1792 ();
 sg13g2_decap_8 FILLER_27_1799 ();
 sg13g2_decap_8 FILLER_27_1806 ();
 sg13g2_decap_8 FILLER_27_1813 ();
 sg13g2_decap_8 FILLER_27_1820 ();
 sg13g2_decap_8 FILLER_27_1827 ();
 sg13g2_decap_8 FILLER_27_1834 ();
 sg13g2_fill_2 FILLER_27_1841 ();
 sg13g2_decap_8 FILLER_27_1848 ();
 sg13g2_decap_8 FILLER_27_1855 ();
 sg13g2_decap_8 FILLER_27_1862 ();
 sg13g2_decap_8 FILLER_27_1869 ();
 sg13g2_decap_8 FILLER_27_1876 ();
 sg13g2_decap_4 FILLER_27_1883 ();
 sg13g2_decap_4 FILLER_27_1892 ();
 sg13g2_decap_8 FILLER_27_1904 ();
 sg13g2_decap_8 FILLER_27_1911 ();
 sg13g2_decap_8 FILLER_27_1918 ();
 sg13g2_decap_8 FILLER_27_1925 ();
 sg13g2_decap_8 FILLER_27_1932 ();
 sg13g2_decap_8 FILLER_27_1939 ();
 sg13g2_fill_2 FILLER_27_1946 ();
 sg13g2_decap_8 FILLER_27_1954 ();
 sg13g2_decap_8 FILLER_27_1961 ();
 sg13g2_decap_8 FILLER_27_1968 ();
 sg13g2_decap_8 FILLER_27_1975 ();
 sg13g2_decap_8 FILLER_27_1982 ();
 sg13g2_decap_8 FILLER_27_1999 ();
 sg13g2_decap_8 FILLER_27_2006 ();
 sg13g2_decap_8 FILLER_27_2013 ();
 sg13g2_decap_8 FILLER_27_2020 ();
 sg13g2_decap_8 FILLER_27_2027 ();
 sg13g2_decap_8 FILLER_27_2034 ();
 sg13g2_decap_8 FILLER_27_2058 ();
 sg13g2_decap_8 FILLER_27_2065 ();
 sg13g2_decap_8 FILLER_27_2072 ();
 sg13g2_decap_8 FILLER_27_2079 ();
 sg13g2_fill_1 FILLER_27_2086 ();
 sg13g2_decap_4 FILLER_27_2097 ();
 sg13g2_decap_8 FILLER_27_2110 ();
 sg13g2_fill_1 FILLER_27_2117 ();
 sg13g2_decap_8 FILLER_27_2126 ();
 sg13g2_decap_8 FILLER_27_2133 ();
 sg13g2_decap_8 FILLER_27_2140 ();
 sg13g2_fill_1 FILLER_27_2147 ();
 sg13g2_decap_8 FILLER_27_2158 ();
 sg13g2_decap_8 FILLER_27_2165 ();
 sg13g2_decap_8 FILLER_27_2172 ();
 sg13g2_decap_8 FILLER_27_2179 ();
 sg13g2_decap_8 FILLER_27_2186 ();
 sg13g2_decap_8 FILLER_27_2193 ();
 sg13g2_decap_4 FILLER_27_2200 ();
 sg13g2_fill_2 FILLER_27_2204 ();
 sg13g2_decap_4 FILLER_27_2211 ();
 sg13g2_decap_8 FILLER_27_2227 ();
 sg13g2_fill_2 FILLER_27_2234 ();
 sg13g2_decap_8 FILLER_27_2262 ();
 sg13g2_decap_8 FILLER_27_2269 ();
 sg13g2_fill_2 FILLER_27_2276 ();
 sg13g2_decap_8 FILLER_27_2284 ();
 sg13g2_decap_4 FILLER_27_2297 ();
 sg13g2_decap_8 FILLER_27_2306 ();
 sg13g2_decap_8 FILLER_27_2313 ();
 sg13g2_fill_2 FILLER_27_2320 ();
 sg13g2_decap_8 FILLER_27_2330 ();
 sg13g2_decap_8 FILLER_27_2337 ();
 sg13g2_decap_8 FILLER_27_2344 ();
 sg13g2_decap_4 FILLER_27_2351 ();
 sg13g2_decap_8 FILLER_27_2365 ();
 sg13g2_decap_8 FILLER_27_2372 ();
 sg13g2_decap_8 FILLER_27_2379 ();
 sg13g2_decap_8 FILLER_27_2386 ();
 sg13g2_decap_8 FILLER_27_2393 ();
 sg13g2_decap_8 FILLER_27_2400 ();
 sg13g2_decap_8 FILLER_27_2438 ();
 sg13g2_fill_2 FILLER_27_2445 ();
 sg13g2_decap_4 FILLER_27_2452 ();
 sg13g2_fill_2 FILLER_27_2476 ();
 sg13g2_fill_1 FILLER_27_2478 ();
 sg13g2_decap_8 FILLER_27_2531 ();
 sg13g2_decap_8 FILLER_27_2538 ();
 sg13g2_decap_8 FILLER_27_2545 ();
 sg13g2_decap_8 FILLER_27_2552 ();
 sg13g2_decap_4 FILLER_27_2559 ();
 sg13g2_fill_2 FILLER_27_2563 ();
 sg13g2_fill_1 FILLER_27_2591 ();
 sg13g2_fill_2 FILLER_27_2607 ();
 sg13g2_decap_8 FILLER_27_2619 ();
 sg13g2_decap_8 FILLER_27_2626 ();
 sg13g2_decap_8 FILLER_27_2633 ();
 sg13g2_fill_2 FILLER_27_2640 ();
 sg13g2_fill_1 FILLER_27_2642 ();
 sg13g2_fill_2 FILLER_27_2653 ();
 sg13g2_decap_8 FILLER_27_2669 ();
 sg13g2_decap_8 FILLER_27_2676 ();
 sg13g2_decap_8 FILLER_27_2683 ();
 sg13g2_fill_1 FILLER_27_2690 ();
 sg13g2_fill_2 FILLER_27_2696 ();
 sg13g2_fill_1 FILLER_27_2698 ();
 sg13g2_decap_4 FILLER_27_2703 ();
 sg13g2_decap_8 FILLER_27_2712 ();
 sg13g2_decap_8 FILLER_27_2719 ();
 sg13g2_decap_8 FILLER_27_2726 ();
 sg13g2_fill_2 FILLER_27_2733 ();
 sg13g2_fill_2 FILLER_27_2741 ();
 sg13g2_fill_1 FILLER_27_2743 ();
 sg13g2_decap_8 FILLER_27_2755 ();
 sg13g2_decap_4 FILLER_27_2762 ();
 sg13g2_fill_1 FILLER_27_2766 ();
 sg13g2_fill_2 FILLER_27_2811 ();
 sg13g2_decap_8 FILLER_27_2819 ();
 sg13g2_decap_8 FILLER_27_2826 ();
 sg13g2_decap_8 FILLER_27_2833 ();
 sg13g2_fill_1 FILLER_27_2840 ();
 sg13g2_decap_8 FILLER_27_2857 ();
 sg13g2_decap_8 FILLER_27_2864 ();
 sg13g2_decap_8 FILLER_27_2871 ();
 sg13g2_decap_8 FILLER_27_2878 ();
 sg13g2_decap_8 FILLER_27_2885 ();
 sg13g2_decap_8 FILLER_27_2892 ();
 sg13g2_decap_8 FILLER_27_2899 ();
 sg13g2_decap_8 FILLER_27_2906 ();
 sg13g2_decap_8 FILLER_27_2913 ();
 sg13g2_decap_4 FILLER_27_2920 ();
 sg13g2_decap_8 FILLER_27_2932 ();
 sg13g2_decap_4 FILLER_27_2939 ();
 sg13g2_fill_2 FILLER_27_2943 ();
 sg13g2_decap_8 FILLER_27_2953 ();
 sg13g2_decap_8 FILLER_27_2960 ();
 sg13g2_decap_8 FILLER_27_2967 ();
 sg13g2_decap_8 FILLER_27_2974 ();
 sg13g2_decap_8 FILLER_27_2981 ();
 sg13g2_decap_8 FILLER_27_2988 ();
 sg13g2_decap_8 FILLER_27_2995 ();
 sg13g2_decap_8 FILLER_27_3002 ();
 sg13g2_decap_8 FILLER_27_3009 ();
 sg13g2_decap_8 FILLER_27_3016 ();
 sg13g2_decap_8 FILLER_27_3023 ();
 sg13g2_decap_4 FILLER_27_3030 ();
 sg13g2_fill_1 FILLER_27_3034 ();
 sg13g2_decap_8 FILLER_27_3055 ();
 sg13g2_decap_4 FILLER_27_3062 ();
 sg13g2_fill_2 FILLER_27_3066 ();
 sg13g2_decap_8 FILLER_27_3094 ();
 sg13g2_fill_1 FILLER_27_3101 ();
 sg13g2_decap_4 FILLER_27_3128 ();
 sg13g2_fill_1 FILLER_27_3132 ();
 sg13g2_decap_8 FILLER_27_3154 ();
 sg13g2_decap_8 FILLER_27_3161 ();
 sg13g2_fill_2 FILLER_27_3168 ();
 sg13g2_fill_1 FILLER_27_3170 ();
 sg13g2_decap_8 FILLER_27_3190 ();
 sg13g2_decap_8 FILLER_27_3197 ();
 sg13g2_decap_8 FILLER_27_3204 ();
 sg13g2_decap_8 FILLER_27_3211 ();
 sg13g2_decap_4 FILLER_27_3218 ();
 sg13g2_fill_1 FILLER_27_3222 ();
 sg13g2_decap_8 FILLER_27_3249 ();
 sg13g2_decap_8 FILLER_27_3256 ();
 sg13g2_decap_8 FILLER_27_3263 ();
 sg13g2_fill_1 FILLER_27_3270 ();
 sg13g2_decap_8 FILLER_27_3307 ();
 sg13g2_fill_2 FILLER_27_3314 ();
 sg13g2_fill_2 FILLER_27_3326 ();
 sg13g2_decap_8 FILLER_27_3354 ();
 sg13g2_decap_8 FILLER_27_3361 ();
 sg13g2_decap_8 FILLER_27_3368 ();
 sg13g2_decap_4 FILLER_27_3375 ();
 sg13g2_fill_2 FILLER_27_3379 ();
 sg13g2_decap_8 FILLER_27_3411 ();
 sg13g2_decap_8 FILLER_27_3418 ();
 sg13g2_decap_4 FILLER_27_3425 ();
 sg13g2_fill_1 FILLER_27_3429 ();
 sg13g2_decap_8 FILLER_27_3456 ();
 sg13g2_decap_8 FILLER_27_3463 ();
 sg13g2_decap_4 FILLER_27_3470 ();
 sg13g2_fill_2 FILLER_27_3474 ();
 sg13g2_decap_8 FILLER_27_3497 ();
 sg13g2_decap_8 FILLER_27_3504 ();
 sg13g2_decap_8 FILLER_27_3511 ();
 sg13g2_decap_8 FILLER_27_3518 ();
 sg13g2_decap_8 FILLER_27_3525 ();
 sg13g2_decap_8 FILLER_27_3532 ();
 sg13g2_decap_8 FILLER_27_3539 ();
 sg13g2_decap_8 FILLER_27_3546 ();
 sg13g2_decap_8 FILLER_27_3553 ();
 sg13g2_decap_8 FILLER_27_3560 ();
 sg13g2_decap_8 FILLER_27_3567 ();
 sg13g2_decap_4 FILLER_27_3574 ();
 sg13g2_fill_2 FILLER_27_3578 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_4 FILLER_28_14 ();
 sg13g2_fill_1 FILLER_28_18 ();
 sg13g2_decap_8 FILLER_28_71 ();
 sg13g2_decap_8 FILLER_28_78 ();
 sg13g2_decap_8 FILLER_28_85 ();
 sg13g2_decap_4 FILLER_28_92 ();
 sg13g2_decap_8 FILLER_28_102 ();
 sg13g2_fill_2 FILLER_28_109 ();
 sg13g2_fill_1 FILLER_28_111 ();
 sg13g2_decap_8 FILLER_28_115 ();
 sg13g2_decap_8 FILLER_28_122 ();
 sg13g2_decap_4 FILLER_28_129 ();
 sg13g2_decap_8 FILLER_28_159 ();
 sg13g2_decap_8 FILLER_28_166 ();
 sg13g2_decap_8 FILLER_28_173 ();
 sg13g2_decap_4 FILLER_28_180 ();
 sg13g2_decap_8 FILLER_28_205 ();
 sg13g2_decap_8 FILLER_28_212 ();
 sg13g2_decap_8 FILLER_28_219 ();
 sg13g2_decap_8 FILLER_28_241 ();
 sg13g2_decap_4 FILLER_28_248 ();
 sg13g2_fill_1 FILLER_28_303 ();
 sg13g2_fill_2 FILLER_28_312 ();
 sg13g2_decap_8 FILLER_28_343 ();
 sg13g2_decap_8 FILLER_28_350 ();
 sg13g2_fill_2 FILLER_28_363 ();
 sg13g2_fill_1 FILLER_28_365 ();
 sg13g2_decap_8 FILLER_28_389 ();
 sg13g2_decap_8 FILLER_28_396 ();
 sg13g2_decap_8 FILLER_28_403 ();
 sg13g2_decap_8 FILLER_28_410 ();
 sg13g2_decap_8 FILLER_28_417 ();
 sg13g2_fill_2 FILLER_28_424 ();
 sg13g2_fill_1 FILLER_28_426 ();
 sg13g2_fill_2 FILLER_28_442 ();
 sg13g2_decap_8 FILLER_28_457 ();
 sg13g2_decap_8 FILLER_28_469 ();
 sg13g2_decap_8 FILLER_28_476 ();
 sg13g2_decap_8 FILLER_28_483 ();
 sg13g2_decap_8 FILLER_28_490 ();
 sg13g2_decap_8 FILLER_28_510 ();
 sg13g2_decap_8 FILLER_28_517 ();
 sg13g2_decap_8 FILLER_28_524 ();
 sg13g2_decap_8 FILLER_28_531 ();
 sg13g2_decap_4 FILLER_28_538 ();
 sg13g2_decap_8 FILLER_28_557 ();
 sg13g2_decap_4 FILLER_28_564 ();
 sg13g2_fill_2 FILLER_28_585 ();
 sg13g2_fill_1 FILLER_28_599 ();
 sg13g2_fill_1 FILLER_28_613 ();
 sg13g2_decap_8 FILLER_28_650 ();
 sg13g2_decap_8 FILLER_28_657 ();
 sg13g2_decap_8 FILLER_28_664 ();
 sg13g2_decap_8 FILLER_28_671 ();
 sg13g2_fill_2 FILLER_28_686 ();
 sg13g2_decap_8 FILLER_28_720 ();
 sg13g2_decap_8 FILLER_28_727 ();
 sg13g2_decap_8 FILLER_28_734 ();
 sg13g2_decap_8 FILLER_28_741 ();
 sg13g2_decap_8 FILLER_28_748 ();
 sg13g2_decap_8 FILLER_28_755 ();
 sg13g2_decap_8 FILLER_28_762 ();
 sg13g2_decap_8 FILLER_28_769 ();
 sg13g2_decap_8 FILLER_28_776 ();
 sg13g2_decap_8 FILLER_28_783 ();
 sg13g2_decap_4 FILLER_28_790 ();
 sg13g2_decap_8 FILLER_28_804 ();
 sg13g2_decap_4 FILLER_28_811 ();
 sg13g2_fill_2 FILLER_28_815 ();
 sg13g2_decap_8 FILLER_28_822 ();
 sg13g2_decap_4 FILLER_28_829 ();
 sg13g2_fill_2 FILLER_28_833 ();
 sg13g2_decap_8 FILLER_28_843 ();
 sg13g2_decap_8 FILLER_28_850 ();
 sg13g2_fill_2 FILLER_28_857 ();
 sg13g2_fill_1 FILLER_28_859 ();
 sg13g2_fill_1 FILLER_28_872 ();
 sg13g2_decap_8 FILLER_28_899 ();
 sg13g2_decap_8 FILLER_28_906 ();
 sg13g2_decap_8 FILLER_28_913 ();
 sg13g2_fill_2 FILLER_28_920 ();
 sg13g2_fill_1 FILLER_28_922 ();
 sg13g2_fill_1 FILLER_28_928 ();
 sg13g2_decap_8 FILLER_28_955 ();
 sg13g2_decap_8 FILLER_28_962 ();
 sg13g2_decap_8 FILLER_28_969 ();
 sg13g2_decap_8 FILLER_28_976 ();
 sg13g2_decap_8 FILLER_28_1000 ();
 sg13g2_decap_8 FILLER_28_1007 ();
 sg13g2_decap_8 FILLER_28_1014 ();
 sg13g2_fill_2 FILLER_28_1021 ();
 sg13g2_fill_1 FILLER_28_1023 ();
 sg13g2_decap_8 FILLER_28_1050 ();
 sg13g2_decap_8 FILLER_28_1057 ();
 sg13g2_decap_8 FILLER_28_1064 ();
 sg13g2_decap_8 FILLER_28_1071 ();
 sg13g2_decap_8 FILLER_28_1078 ();
 sg13g2_decap_8 FILLER_28_1085 ();
 sg13g2_fill_2 FILLER_28_1092 ();
 sg13g2_fill_1 FILLER_28_1094 ();
 sg13g2_decap_8 FILLER_28_1100 ();
 sg13g2_decap_8 FILLER_28_1107 ();
 sg13g2_decap_8 FILLER_28_1114 ();
 sg13g2_decap_8 FILLER_28_1121 ();
 sg13g2_decap_8 FILLER_28_1128 ();
 sg13g2_decap_8 FILLER_28_1135 ();
 sg13g2_decap_4 FILLER_28_1142 ();
 sg13g2_decap_8 FILLER_28_1154 ();
 sg13g2_decap_8 FILLER_28_1161 ();
 sg13g2_decap_8 FILLER_28_1168 ();
 sg13g2_decap_8 FILLER_28_1175 ();
 sg13g2_decap_8 FILLER_28_1182 ();
 sg13g2_decap_8 FILLER_28_1189 ();
 sg13g2_decap_8 FILLER_28_1196 ();
 sg13g2_decap_8 FILLER_28_1203 ();
 sg13g2_decap_8 FILLER_28_1210 ();
 sg13g2_decap_8 FILLER_28_1217 ();
 sg13g2_decap_8 FILLER_28_1224 ();
 sg13g2_decap_8 FILLER_28_1231 ();
 sg13g2_decap_8 FILLER_28_1238 ();
 sg13g2_decap_8 FILLER_28_1245 ();
 sg13g2_decap_8 FILLER_28_1252 ();
 sg13g2_decap_8 FILLER_28_1259 ();
 sg13g2_decap_8 FILLER_28_1266 ();
 sg13g2_decap_8 FILLER_28_1273 ();
 sg13g2_decap_8 FILLER_28_1286 ();
 sg13g2_fill_2 FILLER_28_1293 ();
 sg13g2_fill_1 FILLER_28_1295 ();
 sg13g2_decap_8 FILLER_28_1332 ();
 sg13g2_decap_8 FILLER_28_1339 ();
 sg13g2_decap_8 FILLER_28_1346 ();
 sg13g2_decap_8 FILLER_28_1353 ();
 sg13g2_fill_1 FILLER_28_1360 ();
 sg13g2_decap_8 FILLER_28_1397 ();
 sg13g2_decap_8 FILLER_28_1404 ();
 sg13g2_decap_8 FILLER_28_1411 ();
 sg13g2_decap_8 FILLER_28_1418 ();
 sg13g2_decap_8 FILLER_28_1425 ();
 sg13g2_decap_8 FILLER_28_1432 ();
 sg13g2_fill_1 FILLER_28_1439 ();
 sg13g2_decap_8 FILLER_28_1476 ();
 sg13g2_decap_8 FILLER_28_1483 ();
 sg13g2_decap_8 FILLER_28_1526 ();
 sg13g2_decap_8 FILLER_28_1533 ();
 sg13g2_decap_8 FILLER_28_1540 ();
 sg13g2_decap_8 FILLER_28_1547 ();
 sg13g2_decap_8 FILLER_28_1554 ();
 sg13g2_decap_8 FILLER_28_1561 ();
 sg13g2_decap_8 FILLER_28_1568 ();
 sg13g2_decap_8 FILLER_28_1575 ();
 sg13g2_decap_8 FILLER_28_1582 ();
 sg13g2_decap_8 FILLER_28_1589 ();
 sg13g2_decap_8 FILLER_28_1596 ();
 sg13g2_decap_8 FILLER_28_1603 ();
 sg13g2_decap_8 FILLER_28_1610 ();
 sg13g2_decap_8 FILLER_28_1617 ();
 sg13g2_decap_4 FILLER_28_1624 ();
 sg13g2_fill_2 FILLER_28_1628 ();
 sg13g2_decap_8 FILLER_28_1638 ();
 sg13g2_fill_1 FILLER_28_1645 ();
 sg13g2_decap_8 FILLER_28_1672 ();
 sg13g2_decap_8 FILLER_28_1679 ();
 sg13g2_decap_4 FILLER_28_1686 ();
 sg13g2_fill_1 FILLER_28_1690 ();
 sg13g2_fill_1 FILLER_28_1701 ();
 sg13g2_decap_8 FILLER_28_1728 ();
 sg13g2_decap_4 FILLER_28_1735 ();
 sg13g2_fill_2 FILLER_28_1739 ();
 sg13g2_fill_2 FILLER_28_1773 ();
 sg13g2_decap_8 FILLER_28_1779 ();
 sg13g2_decap_8 FILLER_28_1786 ();
 sg13g2_decap_8 FILLER_28_1793 ();
 sg13g2_decap_8 FILLER_28_1800 ();
 sg13g2_decap_8 FILLER_28_1807 ();
 sg13g2_decap_8 FILLER_28_1814 ();
 sg13g2_decap_8 FILLER_28_1821 ();
 sg13g2_decap_8 FILLER_28_1828 ();
 sg13g2_fill_2 FILLER_28_1835 ();
 sg13g2_decap_8 FILLER_28_1869 ();
 sg13g2_decap_8 FILLER_28_1876 ();
 sg13g2_decap_8 FILLER_28_1883 ();
 sg13g2_decap_8 FILLER_28_1890 ();
 sg13g2_decap_8 FILLER_28_1897 ();
 sg13g2_decap_8 FILLER_28_1904 ();
 sg13g2_decap_8 FILLER_28_1911 ();
 sg13g2_decap_8 FILLER_28_1918 ();
 sg13g2_decap_8 FILLER_28_1925 ();
 sg13g2_decap_8 FILLER_28_1932 ();
 sg13g2_fill_1 FILLER_28_1939 ();
 sg13g2_decap_8 FILLER_28_1950 ();
 sg13g2_decap_8 FILLER_28_1957 ();
 sg13g2_decap_8 FILLER_28_1964 ();
 sg13g2_decap_8 FILLER_28_1971 ();
 sg13g2_decap_8 FILLER_28_1978 ();
 sg13g2_decap_4 FILLER_28_1985 ();
 sg13g2_decap_4 FILLER_28_2015 ();
 sg13g2_fill_2 FILLER_28_2019 ();
 sg13g2_fill_2 FILLER_28_2036 ();
 sg13g2_fill_1 FILLER_28_2038 ();
 sg13g2_fill_2 FILLER_28_2047 ();
 sg13g2_decap_8 FILLER_28_2065 ();
 sg13g2_decap_8 FILLER_28_2072 ();
 sg13g2_decap_8 FILLER_28_2079 ();
 sg13g2_decap_4 FILLER_28_2117 ();
 sg13g2_fill_1 FILLER_28_2131 ();
 sg13g2_decap_8 FILLER_28_2184 ();
 sg13g2_decap_8 FILLER_28_2191 ();
 sg13g2_fill_2 FILLER_28_2198 ();
 sg13g2_fill_2 FILLER_28_2212 ();
 sg13g2_fill_1 FILLER_28_2214 ();
 sg13g2_decap_8 FILLER_28_2221 ();
 sg13g2_decap_8 FILLER_28_2228 ();
 sg13g2_decap_4 FILLER_28_2235 ();
 sg13g2_fill_1 FILLER_28_2239 ();
 sg13g2_decap_4 FILLER_28_2261 ();
 sg13g2_fill_1 FILLER_28_2265 ();
 sg13g2_decap_8 FILLER_28_2277 ();
 sg13g2_decap_4 FILLER_28_2284 ();
 sg13g2_decap_8 FILLER_28_2291 ();
 sg13g2_decap_4 FILLER_28_2298 ();
 sg13g2_fill_2 FILLER_28_2302 ();
 sg13g2_decap_4 FILLER_28_2310 ();
 sg13g2_decap_4 FILLER_28_2322 ();
 sg13g2_fill_2 FILLER_28_2326 ();
 sg13g2_decap_4 FILLER_28_2338 ();
 sg13g2_fill_2 FILLER_28_2342 ();
 sg13g2_decap_8 FILLER_28_2370 ();
 sg13g2_decap_8 FILLER_28_2377 ();
 sg13g2_decap_8 FILLER_28_2384 ();
 sg13g2_decap_8 FILLER_28_2391 ();
 sg13g2_decap_8 FILLER_28_2398 ();
 sg13g2_decap_4 FILLER_28_2405 ();
 sg13g2_fill_1 FILLER_28_2409 ();
 sg13g2_decap_8 FILLER_28_2416 ();
 sg13g2_decap_8 FILLER_28_2423 ();
 sg13g2_decap_8 FILLER_28_2430 ();
 sg13g2_decap_8 FILLER_28_2437 ();
 sg13g2_fill_2 FILLER_28_2444 ();
 sg13g2_decap_8 FILLER_28_2472 ();
 sg13g2_decap_8 FILLER_28_2479 ();
 sg13g2_fill_2 FILLER_28_2486 ();
 sg13g2_decap_8 FILLER_28_2492 ();
 sg13g2_fill_2 FILLER_28_2499 ();
 sg13g2_decap_8 FILLER_28_2516 ();
 sg13g2_decap_8 FILLER_28_2523 ();
 sg13g2_decap_8 FILLER_28_2530 ();
 sg13g2_decap_4 FILLER_28_2537 ();
 sg13g2_decap_4 FILLER_28_2549 ();
 sg13g2_decap_8 FILLER_28_2589 ();
 sg13g2_fill_2 FILLER_28_2596 ();
 sg13g2_decap_8 FILLER_28_2624 ();
 sg13g2_decap_8 FILLER_28_2631 ();
 sg13g2_decap_8 FILLER_28_2638 ();
 sg13g2_decap_8 FILLER_28_2679 ();
 sg13g2_decap_4 FILLER_28_2686 ();
 sg13g2_fill_1 FILLER_28_2690 ();
 sg13g2_decap_8 FILLER_28_2697 ();
 sg13g2_decap_8 FILLER_28_2704 ();
 sg13g2_decap_8 FILLER_28_2711 ();
 sg13g2_decap_8 FILLER_28_2729 ();
 sg13g2_decap_8 FILLER_28_2736 ();
 sg13g2_decap_8 FILLER_28_2743 ();
 sg13g2_decap_8 FILLER_28_2750 ();
 sg13g2_decap_8 FILLER_28_2757 ();
 sg13g2_decap_8 FILLER_28_2764 ();
 sg13g2_decap_8 FILLER_28_2771 ();
 sg13g2_decap_8 FILLER_28_2778 ();
 sg13g2_decap_8 FILLER_28_2785 ();
 sg13g2_decap_4 FILLER_28_2792 ();
 sg13g2_decap_8 FILLER_28_2807 ();
 sg13g2_decap_8 FILLER_28_2814 ();
 sg13g2_decap_8 FILLER_28_2821 ();
 sg13g2_decap_8 FILLER_28_2828 ();
 sg13g2_decap_8 FILLER_28_2835 ();
 sg13g2_fill_2 FILLER_28_2842 ();
 sg13g2_fill_1 FILLER_28_2844 ();
 sg13g2_decap_8 FILLER_28_2856 ();
 sg13g2_fill_2 FILLER_28_2863 ();
 sg13g2_fill_1 FILLER_28_2865 ();
 sg13g2_decap_8 FILLER_28_2871 ();
 sg13g2_fill_2 FILLER_28_2878 ();
 sg13g2_fill_1 FILLER_28_2880 ();
 sg13g2_decap_8 FILLER_28_2891 ();
 sg13g2_decap_8 FILLER_28_2898 ();
 sg13g2_decap_8 FILLER_28_2905 ();
 sg13g2_decap_8 FILLER_28_2912 ();
 sg13g2_decap_8 FILLER_28_2919 ();
 sg13g2_decap_8 FILLER_28_2926 ();
 sg13g2_decap_8 FILLER_28_2933 ();
 sg13g2_decap_4 FILLER_28_2940 ();
 sg13g2_fill_2 FILLER_28_2944 ();
 sg13g2_decap_4 FILLER_28_2972 ();
 sg13g2_fill_1 FILLER_28_2976 ();
 sg13g2_decap_8 FILLER_28_3014 ();
 sg13g2_decap_8 FILLER_28_3021 ();
 sg13g2_decap_8 FILLER_28_3028 ();
 sg13g2_decap_8 FILLER_28_3035 ();
 sg13g2_decap_8 FILLER_28_3042 ();
 sg13g2_decap_8 FILLER_28_3049 ();
 sg13g2_decap_8 FILLER_28_3056 ();
 sg13g2_fill_2 FILLER_28_3063 ();
 sg13g2_decap_8 FILLER_28_3075 ();
 sg13g2_decap_8 FILLER_28_3082 ();
 sg13g2_decap_8 FILLER_28_3089 ();
 sg13g2_fill_1 FILLER_28_3096 ();
 sg13g2_decap_4 FILLER_28_3107 ();
 sg13g2_fill_1 FILLER_28_3111 ();
 sg13g2_decap_8 FILLER_28_3123 ();
 sg13g2_decap_8 FILLER_28_3130 ();
 sg13g2_decap_8 FILLER_28_3137 ();
 sg13g2_decap_8 FILLER_28_3147 ();
 sg13g2_decap_8 FILLER_28_3154 ();
 sg13g2_decap_4 FILLER_28_3161 ();
 sg13g2_fill_2 FILLER_28_3165 ();
 sg13g2_decap_8 FILLER_28_3175 ();
 sg13g2_decap_4 FILLER_28_3182 ();
 sg13g2_decap_8 FILLER_28_3212 ();
 sg13g2_fill_2 FILLER_28_3219 ();
 sg13g2_fill_1 FILLER_28_3221 ();
 sg13g2_decap_8 FILLER_28_3248 ();
 sg13g2_decap_8 FILLER_28_3255 ();
 sg13g2_decap_8 FILLER_28_3262 ();
 sg13g2_decap_8 FILLER_28_3277 ();
 sg13g2_decap_8 FILLER_28_3284 ();
 sg13g2_fill_2 FILLER_28_3291 ();
 sg13g2_decap_8 FILLER_28_3298 ();
 sg13g2_fill_2 FILLER_28_3305 ();
 sg13g2_fill_2 FILLER_28_3312 ();
 sg13g2_decap_8 FILLER_28_3350 ();
 sg13g2_fill_2 FILLER_28_3357 ();
 sg13g2_decap_8 FILLER_28_3369 ();
 sg13g2_fill_2 FILLER_28_3376 ();
 sg13g2_fill_1 FILLER_28_3378 ();
 sg13g2_decap_8 FILLER_28_3415 ();
 sg13g2_decap_8 FILLER_28_3422 ();
 sg13g2_decap_8 FILLER_28_3429 ();
 sg13g2_fill_2 FILLER_28_3436 ();
 sg13g2_decap_8 FILLER_28_3443 ();
 sg13g2_decap_8 FILLER_28_3450 ();
 sg13g2_decap_8 FILLER_28_3457 ();
 sg13g2_decap_8 FILLER_28_3464 ();
 sg13g2_decap_8 FILLER_28_3471 ();
 sg13g2_decap_8 FILLER_28_3478 ();
 sg13g2_fill_2 FILLER_28_3485 ();
 sg13g2_decap_8 FILLER_28_3497 ();
 sg13g2_fill_2 FILLER_28_3504 ();
 sg13g2_decap_4 FILLER_28_3516 ();
 sg13g2_fill_1 FILLER_28_3520 ();
 sg13g2_decap_4 FILLER_28_3531 ();
 sg13g2_decap_8 FILLER_28_3561 ();
 sg13g2_decap_8 FILLER_28_3568 ();
 sg13g2_decap_4 FILLER_28_3575 ();
 sg13g2_fill_1 FILLER_28_3579 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_fill_2 FILLER_29_7 ();
 sg13g2_fill_1 FILLER_29_9 ();
 sg13g2_fill_1 FILLER_29_45 ();
 sg13g2_decap_8 FILLER_29_73 ();
 sg13g2_fill_2 FILLER_29_80 ();
 sg13g2_fill_1 FILLER_29_82 ();
 sg13g2_decap_8 FILLER_29_127 ();
 sg13g2_decap_4 FILLER_29_134 ();
 sg13g2_fill_2 FILLER_29_138 ();
 sg13g2_decap_8 FILLER_29_159 ();
 sg13g2_decap_8 FILLER_29_166 ();
 sg13g2_decap_8 FILLER_29_173 ();
 sg13g2_decap_8 FILLER_29_180 ();
 sg13g2_decap_8 FILLER_29_187 ();
 sg13g2_decap_8 FILLER_29_194 ();
 sg13g2_decap_4 FILLER_29_201 ();
 sg13g2_decap_8 FILLER_29_210 ();
 sg13g2_decap_8 FILLER_29_217 ();
 sg13g2_decap_8 FILLER_29_224 ();
 sg13g2_fill_2 FILLER_29_231 ();
 sg13g2_fill_1 FILLER_29_233 ();
 sg13g2_decap_8 FILLER_29_239 ();
 sg13g2_decap_8 FILLER_29_246 ();
 sg13g2_decap_4 FILLER_29_253 ();
 sg13g2_fill_1 FILLER_29_257 ();
 sg13g2_fill_1 FILLER_29_263 ();
 sg13g2_decap_8 FILLER_29_283 ();
 sg13g2_decap_8 FILLER_29_290 ();
 sg13g2_decap_8 FILLER_29_297 ();
 sg13g2_decap_8 FILLER_29_304 ();
 sg13g2_decap_8 FILLER_29_311 ();
 sg13g2_decap_4 FILLER_29_318 ();
 sg13g2_decap_8 FILLER_29_331 ();
 sg13g2_decap_8 FILLER_29_338 ();
 sg13g2_decap_8 FILLER_29_345 ();
 sg13g2_decap_8 FILLER_29_352 ();
 sg13g2_decap_8 FILLER_29_359 ();
 sg13g2_fill_1 FILLER_29_387 ();
 sg13g2_decap_4 FILLER_29_402 ();
 sg13g2_fill_1 FILLER_29_406 ();
 sg13g2_decap_8 FILLER_29_416 ();
 sg13g2_decap_8 FILLER_29_423 ();
 sg13g2_fill_2 FILLER_29_430 ();
 sg13g2_decap_8 FILLER_29_437 ();
 sg13g2_decap_8 FILLER_29_444 ();
 sg13g2_decap_8 FILLER_29_451 ();
 sg13g2_decap_8 FILLER_29_458 ();
 sg13g2_decap_8 FILLER_29_465 ();
 sg13g2_decap_8 FILLER_29_472 ();
 sg13g2_fill_1 FILLER_29_484 ();
 sg13g2_decap_8 FILLER_29_505 ();
 sg13g2_decap_8 FILLER_29_512 ();
 sg13g2_decap_8 FILLER_29_519 ();
 sg13g2_decap_8 FILLER_29_526 ();
 sg13g2_decap_8 FILLER_29_533 ();
 sg13g2_decap_4 FILLER_29_540 ();
 sg13g2_fill_2 FILLER_29_548 ();
 sg13g2_decap_8 FILLER_29_566 ();
 sg13g2_decap_4 FILLER_29_573 ();
 sg13g2_decap_8 FILLER_29_602 ();
 sg13g2_decap_8 FILLER_29_609 ();
 sg13g2_decap_8 FILLER_29_616 ();
 sg13g2_decap_4 FILLER_29_623 ();
 sg13g2_fill_1 FILLER_29_627 ();
 sg13g2_fill_2 FILLER_29_634 ();
 sg13g2_fill_1 FILLER_29_636 ();
 sg13g2_decap_8 FILLER_29_658 ();
 sg13g2_decap_4 FILLER_29_665 ();
 sg13g2_fill_1 FILLER_29_669 ();
 sg13g2_decap_8 FILLER_29_678 ();
 sg13g2_decap_8 FILLER_29_685 ();
 sg13g2_decap_8 FILLER_29_692 ();
 sg13g2_decap_4 FILLER_29_699 ();
 sg13g2_fill_2 FILLER_29_703 ();
 sg13g2_decap_8 FILLER_29_730 ();
 sg13g2_decap_8 FILLER_29_737 ();
 sg13g2_decap_8 FILLER_29_744 ();
 sg13g2_decap_8 FILLER_29_751 ();
 sg13g2_decap_8 FILLER_29_758 ();
 sg13g2_decap_8 FILLER_29_765 ();
 sg13g2_decap_8 FILLER_29_772 ();
 sg13g2_decap_8 FILLER_29_779 ();
 sg13g2_decap_8 FILLER_29_786 ();
 sg13g2_fill_2 FILLER_29_793 ();
 sg13g2_fill_1 FILLER_29_795 ();
 sg13g2_decap_8 FILLER_29_806 ();
 sg13g2_decap_8 FILLER_29_813 ();
 sg13g2_fill_2 FILLER_29_820 ();
 sg13g2_fill_2 FILLER_29_858 ();
 sg13g2_decap_8 FILLER_29_905 ();
 sg13g2_decap_8 FILLER_29_912 ();
 sg13g2_fill_1 FILLER_29_919 ();
 sg13g2_fill_2 FILLER_29_930 ();
 sg13g2_fill_1 FILLER_29_932 ();
 sg13g2_decap_8 FILLER_29_967 ();
 sg13g2_decap_8 FILLER_29_974 ();
 sg13g2_fill_1 FILLER_29_1011 ();
 sg13g2_decap_8 FILLER_29_1022 ();
 sg13g2_decap_8 FILLER_29_1029 ();
 sg13g2_decap_8 FILLER_29_1036 ();
 sg13g2_decap_8 FILLER_29_1043 ();
 sg13g2_decap_8 FILLER_29_1050 ();
 sg13g2_decap_4 FILLER_29_1057 ();
 sg13g2_fill_2 FILLER_29_1061 ();
 sg13g2_fill_2 FILLER_29_1099 ();
 sg13g2_decap_8 FILLER_29_1135 ();
 sg13g2_decap_8 FILLER_29_1142 ();
 sg13g2_fill_1 FILLER_29_1149 ();
 sg13g2_decap_8 FILLER_29_1170 ();
 sg13g2_decap_8 FILLER_29_1177 ();
 sg13g2_decap_8 FILLER_29_1184 ();
 sg13g2_decap_8 FILLER_29_1191 ();
 sg13g2_decap_8 FILLER_29_1198 ();
 sg13g2_decap_8 FILLER_29_1205 ();
 sg13g2_fill_1 FILLER_29_1212 ();
 sg13g2_decap_4 FILLER_29_1249 ();
 sg13g2_decap_8 FILLER_29_1263 ();
 sg13g2_decap_8 FILLER_29_1270 ();
 sg13g2_decap_8 FILLER_29_1277 ();
 sg13g2_decap_8 FILLER_29_1284 ();
 sg13g2_decap_8 FILLER_29_1291 ();
 sg13g2_decap_8 FILLER_29_1298 ();
 sg13g2_decap_8 FILLER_29_1305 ();
 sg13g2_decap_8 FILLER_29_1312 ();
 sg13g2_decap_8 FILLER_29_1319 ();
 sg13g2_decap_8 FILLER_29_1326 ();
 sg13g2_decap_8 FILLER_29_1333 ();
 sg13g2_decap_8 FILLER_29_1340 ();
 sg13g2_decap_8 FILLER_29_1347 ();
 sg13g2_decap_8 FILLER_29_1354 ();
 sg13g2_decap_8 FILLER_29_1361 ();
 sg13g2_decap_8 FILLER_29_1368 ();
 sg13g2_decap_8 FILLER_29_1392 ();
 sg13g2_decap_8 FILLER_29_1399 ();
 sg13g2_decap_8 FILLER_29_1406 ();
 sg13g2_decap_8 FILLER_29_1413 ();
 sg13g2_decap_8 FILLER_29_1420 ();
 sg13g2_decap_8 FILLER_29_1427 ();
 sg13g2_decap_8 FILLER_29_1434 ();
 sg13g2_decap_8 FILLER_29_1441 ();
 sg13g2_decap_8 FILLER_29_1448 ();
 sg13g2_decap_8 FILLER_29_1455 ();
 sg13g2_decap_8 FILLER_29_1462 ();
 sg13g2_decap_8 FILLER_29_1469 ();
 sg13g2_decap_8 FILLER_29_1476 ();
 sg13g2_decap_8 FILLER_29_1483 ();
 sg13g2_decap_8 FILLER_29_1490 ();
 sg13g2_decap_4 FILLER_29_1497 ();
 sg13g2_fill_2 FILLER_29_1501 ();
 sg13g2_decap_8 FILLER_29_1539 ();
 sg13g2_decap_8 FILLER_29_1546 ();
 sg13g2_decap_8 FILLER_29_1559 ();
 sg13g2_fill_1 FILLER_29_1566 ();
 sg13g2_decap_8 FILLER_29_1575 ();
 sg13g2_fill_2 FILLER_29_1582 ();
 sg13g2_fill_1 FILLER_29_1584 ();
 sg13g2_decap_8 FILLER_29_1611 ();
 sg13g2_decap_8 FILLER_29_1618 ();
 sg13g2_decap_4 FILLER_29_1625 ();
 sg13g2_decap_8 FILLER_29_1635 ();
 sg13g2_decap_4 FILLER_29_1642 ();
 sg13g2_decap_4 FILLER_29_1652 ();
 sg13g2_fill_2 FILLER_29_1656 ();
 sg13g2_decap_8 FILLER_29_1694 ();
 sg13g2_decap_4 FILLER_29_1701 ();
 sg13g2_fill_1 FILLER_29_1705 ();
 sg13g2_decap_8 FILLER_29_1716 ();
 sg13g2_decap_8 FILLER_29_1723 ();
 sg13g2_decap_8 FILLER_29_1730 ();
 sg13g2_decap_8 FILLER_29_1737 ();
 sg13g2_fill_2 FILLER_29_1744 ();
 sg13g2_decap_8 FILLER_29_1761 ();
 sg13g2_decap_8 FILLER_29_1768 ();
 sg13g2_decap_8 FILLER_29_1775 ();
 sg13g2_decap_4 FILLER_29_1782 ();
 sg13g2_decap_8 FILLER_29_1794 ();
 sg13g2_decap_8 FILLER_29_1801 ();
 sg13g2_decap_8 FILLER_29_1808 ();
 sg13g2_decap_4 FILLER_29_1815 ();
 sg13g2_fill_2 FILLER_29_1829 ();
 sg13g2_decap_8 FILLER_29_1857 ();
 sg13g2_decap_8 FILLER_29_1864 ();
 sg13g2_decap_8 FILLER_29_1871 ();
 sg13g2_decap_4 FILLER_29_1878 ();
 sg13g2_fill_1 FILLER_29_1882 ();
 sg13g2_decap_8 FILLER_29_1888 ();
 sg13g2_decap_4 FILLER_29_1895 ();
 sg13g2_fill_2 FILLER_29_1899 ();
 sg13g2_decap_8 FILLER_29_1906 ();
 sg13g2_decap_8 FILLER_29_1913 ();
 sg13g2_fill_1 FILLER_29_1920 ();
 sg13g2_decap_8 FILLER_29_1973 ();
 sg13g2_decap_8 FILLER_29_1980 ();
 sg13g2_decap_8 FILLER_29_1987 ();
 sg13g2_fill_2 FILLER_29_1994 ();
 sg13g2_fill_1 FILLER_29_1996 ();
 sg13g2_decap_4 FILLER_29_2005 ();
 sg13g2_fill_2 FILLER_29_2009 ();
 sg13g2_decap_8 FILLER_29_2021 ();
 sg13g2_decap_8 FILLER_29_2028 ();
 sg13g2_decap_8 FILLER_29_2035 ();
 sg13g2_decap_8 FILLER_29_2042 ();
 sg13g2_fill_1 FILLER_29_2049 ();
 sg13g2_decap_8 FILLER_29_2058 ();
 sg13g2_decap_8 FILLER_29_2077 ();
 sg13g2_decap_8 FILLER_29_2084 ();
 sg13g2_decap_8 FILLER_29_2091 ();
 sg13g2_decap_8 FILLER_29_2098 ();
 sg13g2_decap_8 FILLER_29_2105 ();
 sg13g2_decap_8 FILLER_29_2112 ();
 sg13g2_decap_8 FILLER_29_2119 ();
 sg13g2_decap_8 FILLER_29_2126 ();
 sg13g2_decap_8 FILLER_29_2133 ();
 sg13g2_decap_8 FILLER_29_2140 ();
 sg13g2_decap_8 FILLER_29_2147 ();
 sg13g2_decap_8 FILLER_29_2154 ();
 sg13g2_decap_8 FILLER_29_2161 ();
 sg13g2_decap_8 FILLER_29_2168 ();
 sg13g2_decap_8 FILLER_29_2175 ();
 sg13g2_decap_8 FILLER_29_2182 ();
 sg13g2_decap_8 FILLER_29_2189 ();
 sg13g2_decap_4 FILLER_29_2196 ();
 sg13g2_fill_1 FILLER_29_2200 ();
 sg13g2_decap_8 FILLER_29_2213 ();
 sg13g2_decap_8 FILLER_29_2220 ();
 sg13g2_decap_8 FILLER_29_2227 ();
 sg13g2_decap_8 FILLER_29_2234 ();
 sg13g2_fill_2 FILLER_29_2241 ();
 sg13g2_fill_1 FILLER_29_2243 ();
 sg13g2_decap_8 FILLER_29_2250 ();
 sg13g2_decap_8 FILLER_29_2257 ();
 sg13g2_decap_4 FILLER_29_2264 ();
 sg13g2_decap_8 FILLER_29_2276 ();
 sg13g2_decap_8 FILLER_29_2283 ();
 sg13g2_decap_8 FILLER_29_2290 ();
 sg13g2_decap_8 FILLER_29_2297 ();
 sg13g2_decap_8 FILLER_29_2315 ();
 sg13g2_decap_8 FILLER_29_2322 ();
 sg13g2_decap_8 FILLER_29_2329 ();
 sg13g2_decap_8 FILLER_29_2336 ();
 sg13g2_decap_8 FILLER_29_2343 ();
 sg13g2_decap_4 FILLER_29_2350 ();
 sg13g2_fill_2 FILLER_29_2354 ();
 sg13g2_decap_8 FILLER_29_2385 ();
 sg13g2_decap_8 FILLER_29_2392 ();
 sg13g2_decap_8 FILLER_29_2399 ();
 sg13g2_decap_8 FILLER_29_2406 ();
 sg13g2_decap_4 FILLER_29_2413 ();
 sg13g2_decap_8 FILLER_29_2423 ();
 sg13g2_decap_8 FILLER_29_2430 ();
 sg13g2_decap_8 FILLER_29_2437 ();
 sg13g2_decap_8 FILLER_29_2444 ();
 sg13g2_decap_4 FILLER_29_2451 ();
 sg13g2_fill_2 FILLER_29_2455 ();
 sg13g2_decap_8 FILLER_29_2460 ();
 sg13g2_decap_8 FILLER_29_2467 ();
 sg13g2_decap_8 FILLER_29_2474 ();
 sg13g2_decap_8 FILLER_29_2481 ();
 sg13g2_decap_8 FILLER_29_2488 ();
 sg13g2_decap_8 FILLER_29_2495 ();
 sg13g2_decap_4 FILLER_29_2502 ();
 sg13g2_decap_8 FILLER_29_2510 ();
 sg13g2_decap_8 FILLER_29_2517 ();
 sg13g2_decap_8 FILLER_29_2524 ();
 sg13g2_decap_4 FILLER_29_2537 ();
 sg13g2_decap_8 FILLER_29_2552 ();
 sg13g2_fill_2 FILLER_29_2569 ();
 sg13g2_fill_1 FILLER_29_2571 ();
 sg13g2_decap_8 FILLER_29_2580 ();
 sg13g2_decap_8 FILLER_29_2587 ();
 sg13g2_decap_8 FILLER_29_2594 ();
 sg13g2_decap_8 FILLER_29_2601 ();
 sg13g2_decap_8 FILLER_29_2608 ();
 sg13g2_decap_8 FILLER_29_2615 ();
 sg13g2_fill_2 FILLER_29_2622 ();
 sg13g2_decap_4 FILLER_29_2639 ();
 sg13g2_fill_2 FILLER_29_2643 ();
 sg13g2_decap_8 FILLER_29_2659 ();
 sg13g2_decap_4 FILLER_29_2666 ();
 sg13g2_fill_1 FILLER_29_2670 ();
 sg13g2_decap_8 FILLER_29_2684 ();
 sg13g2_decap_8 FILLER_29_2691 ();
 sg13g2_decap_8 FILLER_29_2698 ();
 sg13g2_fill_1 FILLER_29_2705 ();
 sg13g2_decap_8 FILLER_29_2711 ();
 sg13g2_decap_8 FILLER_29_2718 ();
 sg13g2_decap_8 FILLER_29_2725 ();
 sg13g2_fill_2 FILLER_29_2732 ();
 sg13g2_decap_8 FILLER_29_2745 ();
 sg13g2_decap_8 FILLER_29_2752 ();
 sg13g2_decap_8 FILLER_29_2759 ();
 sg13g2_decap_8 FILLER_29_2766 ();
 sg13g2_decap_8 FILLER_29_2799 ();
 sg13g2_decap_8 FILLER_29_2806 ();
 sg13g2_decap_8 FILLER_29_2813 ();
 sg13g2_decap_4 FILLER_29_2820 ();
 sg13g2_decap_8 FILLER_29_2856 ();
 sg13g2_decap_8 FILLER_29_2863 ();
 sg13g2_decap_8 FILLER_29_2870 ();
 sg13g2_decap_4 FILLER_29_2877 ();
 sg13g2_fill_1 FILLER_29_2881 ();
 sg13g2_decap_8 FILLER_29_2918 ();
 sg13g2_decap_8 FILLER_29_2925 ();
 sg13g2_decap_8 FILLER_29_2932 ();
 sg13g2_fill_2 FILLER_29_2939 ();
 sg13g2_fill_1 FILLER_29_2941 ();
 sg13g2_decap_8 FILLER_29_2952 ();
 sg13g2_decap_8 FILLER_29_2959 ();
 sg13g2_decap_4 FILLER_29_2966 ();
 sg13g2_fill_1 FILLER_29_2970 ();
 sg13g2_decap_8 FILLER_29_2981 ();
 sg13g2_decap_8 FILLER_29_2988 ();
 sg13g2_decap_8 FILLER_29_2995 ();
 sg13g2_decap_8 FILLER_29_3002 ();
 sg13g2_decap_8 FILLER_29_3009 ();
 sg13g2_decap_8 FILLER_29_3016 ();
 sg13g2_decap_4 FILLER_29_3023 ();
 sg13g2_decap_8 FILLER_29_3048 ();
 sg13g2_decap_8 FILLER_29_3055 ();
 sg13g2_decap_8 FILLER_29_3062 ();
 sg13g2_decap_8 FILLER_29_3069 ();
 sg13g2_decap_8 FILLER_29_3076 ();
 sg13g2_decap_8 FILLER_29_3083 ();
 sg13g2_decap_8 FILLER_29_3090 ();
 sg13g2_decap_8 FILLER_29_3097 ();
 sg13g2_decap_4 FILLER_29_3104 ();
 sg13g2_fill_1 FILLER_29_3108 ();
 sg13g2_decap_8 FILLER_29_3119 ();
 sg13g2_decap_8 FILLER_29_3126 ();
 sg13g2_decap_8 FILLER_29_3133 ();
 sg13g2_decap_8 FILLER_29_3140 ();
 sg13g2_decap_4 FILLER_29_3147 ();
 sg13g2_fill_1 FILLER_29_3151 ();
 sg13g2_decap_8 FILLER_29_3160 ();
 sg13g2_fill_1 FILLER_29_3167 ();
 sg13g2_fill_2 FILLER_29_3176 ();
 sg13g2_fill_1 FILLER_29_3178 ();
 sg13g2_decap_8 FILLER_29_3184 ();
 sg13g2_decap_8 FILLER_29_3191 ();
 sg13g2_decap_8 FILLER_29_3198 ();
 sg13g2_decap_8 FILLER_29_3205 ();
 sg13g2_decap_8 FILLER_29_3212 ();
 sg13g2_decap_8 FILLER_29_3219 ();
 sg13g2_decap_4 FILLER_29_3226 ();
 sg13g2_fill_1 FILLER_29_3230 ();
 sg13g2_decap_8 FILLER_29_3241 ();
 sg13g2_decap_8 FILLER_29_3248 ();
 sg13g2_decap_8 FILLER_29_3255 ();
 sg13g2_decap_8 FILLER_29_3262 ();
 sg13g2_decap_8 FILLER_29_3269 ();
 sg13g2_decap_8 FILLER_29_3276 ();
 sg13g2_decap_8 FILLER_29_3283 ();
 sg13g2_decap_8 FILLER_29_3290 ();
 sg13g2_decap_8 FILLER_29_3297 ();
 sg13g2_decap_8 FILLER_29_3304 ();
 sg13g2_decap_8 FILLER_29_3311 ();
 sg13g2_decap_8 FILLER_29_3318 ();
 sg13g2_decap_8 FILLER_29_3325 ();
 sg13g2_decap_8 FILLER_29_3332 ();
 sg13g2_decap_8 FILLER_29_3339 ();
 sg13g2_decap_8 FILLER_29_3346 ();
 sg13g2_decap_8 FILLER_29_3353 ();
 sg13g2_fill_2 FILLER_29_3360 ();
 sg13g2_fill_1 FILLER_29_3362 ();
 sg13g2_decap_8 FILLER_29_3389 ();
 sg13g2_decap_8 FILLER_29_3396 ();
 sg13g2_decap_8 FILLER_29_3403 ();
 sg13g2_decap_8 FILLER_29_3410 ();
 sg13g2_decap_8 FILLER_29_3417 ();
 sg13g2_decap_8 FILLER_29_3424 ();
 sg13g2_decap_8 FILLER_29_3431 ();
 sg13g2_decap_8 FILLER_29_3438 ();
 sg13g2_decap_8 FILLER_29_3445 ();
 sg13g2_decap_8 FILLER_29_3452 ();
 sg13g2_decap_8 FILLER_29_3459 ();
 sg13g2_decap_8 FILLER_29_3466 ();
 sg13g2_decap_8 FILLER_29_3473 ();
 sg13g2_fill_2 FILLER_29_3480 ();
 sg13g2_decap_8 FILLER_29_3513 ();
 sg13g2_decap_4 FILLER_29_3520 ();
 sg13g2_fill_1 FILLER_29_3524 ();
 sg13g2_fill_2 FILLER_29_3577 ();
 sg13g2_fill_1 FILLER_29_3579 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_fill_2 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_51 ();
 sg13g2_decap_8 FILLER_30_58 ();
 sg13g2_decap_8 FILLER_30_65 ();
 sg13g2_decap_8 FILLER_30_72 ();
 sg13g2_decap_4 FILLER_30_79 ();
 sg13g2_fill_1 FILLER_30_83 ();
 sg13g2_fill_2 FILLER_30_92 ();
 sg13g2_decap_8 FILLER_30_111 ();
 sg13g2_decap_8 FILLER_30_118 ();
 sg13g2_decap_8 FILLER_30_125 ();
 sg13g2_decap_8 FILLER_30_132 ();
 sg13g2_decap_4 FILLER_30_139 ();
 sg13g2_fill_2 FILLER_30_143 ();
 sg13g2_fill_2 FILLER_30_150 ();
 sg13g2_decap_8 FILLER_30_160 ();
 sg13g2_decap_8 FILLER_30_167 ();
 sg13g2_decap_8 FILLER_30_174 ();
 sg13g2_decap_8 FILLER_30_181 ();
 sg13g2_decap_8 FILLER_30_188 ();
 sg13g2_decap_8 FILLER_30_195 ();
 sg13g2_decap_8 FILLER_30_202 ();
 sg13g2_decap_8 FILLER_30_209 ();
 sg13g2_decap_8 FILLER_30_216 ();
 sg13g2_decap_8 FILLER_30_223 ();
 sg13g2_decap_8 FILLER_30_230 ();
 sg13g2_decap_8 FILLER_30_237 ();
 sg13g2_decap_8 FILLER_30_244 ();
 sg13g2_decap_8 FILLER_30_251 ();
 sg13g2_decap_8 FILLER_30_258 ();
 sg13g2_decap_8 FILLER_30_265 ();
 sg13g2_decap_8 FILLER_30_272 ();
 sg13g2_decap_8 FILLER_30_279 ();
 sg13g2_decap_8 FILLER_30_286 ();
 sg13g2_decap_8 FILLER_30_293 ();
 sg13g2_decap_8 FILLER_30_300 ();
 sg13g2_decap_8 FILLER_30_307 ();
 sg13g2_decap_8 FILLER_30_314 ();
 sg13g2_decap_8 FILLER_30_321 ();
 sg13g2_decap_8 FILLER_30_328 ();
 sg13g2_decap_8 FILLER_30_335 ();
 sg13g2_decap_8 FILLER_30_342 ();
 sg13g2_decap_8 FILLER_30_349 ();
 sg13g2_decap_4 FILLER_30_356 ();
 sg13g2_fill_2 FILLER_30_360 ();
 sg13g2_decap_8 FILLER_30_381 ();
 sg13g2_decap_4 FILLER_30_388 ();
 sg13g2_decap_4 FILLER_30_397 ();
 sg13g2_decap_8 FILLER_30_427 ();
 sg13g2_decap_8 FILLER_30_434 ();
 sg13g2_decap_8 FILLER_30_441 ();
 sg13g2_fill_1 FILLER_30_448 ();
 sg13g2_decap_8 FILLER_30_454 ();
 sg13g2_decap_8 FILLER_30_461 ();
 sg13g2_decap_8 FILLER_30_468 ();
 sg13g2_decap_8 FILLER_30_475 ();
 sg13g2_decap_8 FILLER_30_482 ();
 sg13g2_decap_8 FILLER_30_489 ();
 sg13g2_decap_8 FILLER_30_496 ();
 sg13g2_fill_2 FILLER_30_507 ();
 sg13g2_decap_8 FILLER_30_514 ();
 sg13g2_decap_8 FILLER_30_521 ();
 sg13g2_fill_2 FILLER_30_528 ();
 sg13g2_fill_1 FILLER_30_530 ();
 sg13g2_decap_8 FILLER_30_535 ();
 sg13g2_fill_2 FILLER_30_542 ();
 sg13g2_decap_8 FILLER_30_562 ();
 sg13g2_decap_8 FILLER_30_569 ();
 sg13g2_decap_8 FILLER_30_576 ();
 sg13g2_decap_4 FILLER_30_583 ();
 sg13g2_fill_2 FILLER_30_587 ();
 sg13g2_decap_8 FILLER_30_595 ();
 sg13g2_decap_8 FILLER_30_602 ();
 sg13g2_decap_8 FILLER_30_609 ();
 sg13g2_decap_8 FILLER_30_616 ();
 sg13g2_decap_8 FILLER_30_623 ();
 sg13g2_decap_8 FILLER_30_630 ();
 sg13g2_decap_8 FILLER_30_637 ();
 sg13g2_decap_8 FILLER_30_644 ();
 sg13g2_decap_8 FILLER_30_651 ();
 sg13g2_decap_4 FILLER_30_658 ();
 sg13g2_decap_4 FILLER_30_670 ();
 sg13g2_fill_1 FILLER_30_674 ();
 sg13g2_decap_8 FILLER_30_698 ();
 sg13g2_fill_2 FILLER_30_705 ();
 sg13g2_fill_2 FILLER_30_713 ();
 sg13g2_fill_2 FILLER_30_729 ();
 sg13g2_decap_4 FILLER_30_737 ();
 sg13g2_decap_8 FILLER_30_752 ();
 sg13g2_decap_8 FILLER_30_759 ();
 sg13g2_decap_8 FILLER_30_766 ();
 sg13g2_decap_8 FILLER_30_773 ();
 sg13g2_decap_8 FILLER_30_780 ();
 sg13g2_decap_4 FILLER_30_787 ();
 sg13g2_decap_8 FILLER_30_817 ();
 sg13g2_decap_8 FILLER_30_824 ();
 sg13g2_decap_8 FILLER_30_831 ();
 sg13g2_decap_8 FILLER_30_838 ();
 sg13g2_decap_8 FILLER_30_845 ();
 sg13g2_decap_8 FILLER_30_852 ();
 sg13g2_decap_8 FILLER_30_859 ();
 sg13g2_decap_8 FILLER_30_866 ();
 sg13g2_fill_2 FILLER_30_873 ();
 sg13g2_fill_1 FILLER_30_875 ();
 sg13g2_decap_8 FILLER_30_882 ();
 sg13g2_decap_8 FILLER_30_889 ();
 sg13g2_decap_8 FILLER_30_896 ();
 sg13g2_decap_8 FILLER_30_903 ();
 sg13g2_decap_8 FILLER_30_910 ();
 sg13g2_decap_8 FILLER_30_917 ();
 sg13g2_fill_2 FILLER_30_924 ();
 sg13g2_fill_1 FILLER_30_926 ();
 sg13g2_decap_8 FILLER_30_937 ();
 sg13g2_decap_8 FILLER_30_944 ();
 sg13g2_decap_8 FILLER_30_951 ();
 sg13g2_decap_8 FILLER_30_958 ();
 sg13g2_decap_8 FILLER_30_965 ();
 sg13g2_decap_8 FILLER_30_972 ();
 sg13g2_decap_8 FILLER_30_979 ();
 sg13g2_fill_1 FILLER_30_991 ();
 sg13g2_decap_8 FILLER_30_998 ();
 sg13g2_decap_8 FILLER_30_1005 ();
 sg13g2_decap_8 FILLER_30_1012 ();
 sg13g2_decap_8 FILLER_30_1019 ();
 sg13g2_decap_8 FILLER_30_1036 ();
 sg13g2_fill_2 FILLER_30_1043 ();
 sg13g2_fill_1 FILLER_30_1045 ();
 sg13g2_fill_2 FILLER_30_1072 ();
 sg13g2_fill_1 FILLER_30_1100 ();
 sg13g2_decap_8 FILLER_30_1111 ();
 sg13g2_decap_8 FILLER_30_1118 ();
 sg13g2_decap_8 FILLER_30_1125 ();
 sg13g2_decap_8 FILLER_30_1132 ();
 sg13g2_decap_8 FILLER_30_1139 ();
 sg13g2_decap_8 FILLER_30_1146 ();
 sg13g2_decap_8 FILLER_30_1153 ();
 sg13g2_fill_1 FILLER_30_1160 ();
 sg13g2_decap_8 FILLER_30_1197 ();
 sg13g2_decap_8 FILLER_30_1204 ();
 sg13g2_fill_2 FILLER_30_1211 ();
 sg13g2_decap_8 FILLER_30_1247 ();
 sg13g2_decap_4 FILLER_30_1254 ();
 sg13g2_fill_1 FILLER_30_1258 ();
 sg13g2_decap_8 FILLER_30_1285 ();
 sg13g2_decap_4 FILLER_30_1292 ();
 sg13g2_decap_8 FILLER_30_1306 ();
 sg13g2_decap_8 FILLER_30_1313 ();
 sg13g2_decap_8 FILLER_30_1320 ();
 sg13g2_decap_8 FILLER_30_1327 ();
 sg13g2_decap_8 FILLER_30_1334 ();
 sg13g2_decap_8 FILLER_30_1341 ();
 sg13g2_fill_2 FILLER_30_1348 ();
 sg13g2_fill_1 FILLER_30_1350 ();
 sg13g2_decap_8 FILLER_30_1357 ();
 sg13g2_decap_4 FILLER_30_1364 ();
 sg13g2_fill_2 FILLER_30_1368 ();
 sg13g2_decap_8 FILLER_30_1378 ();
 sg13g2_decap_8 FILLER_30_1385 ();
 sg13g2_decap_8 FILLER_30_1392 ();
 sg13g2_decap_8 FILLER_30_1399 ();
 sg13g2_decap_4 FILLER_30_1406 ();
 sg13g2_fill_1 FILLER_30_1410 ();
 sg13g2_decap_4 FILLER_30_1415 ();
 sg13g2_fill_1 FILLER_30_1419 ();
 sg13g2_decap_8 FILLER_30_1424 ();
 sg13g2_decap_8 FILLER_30_1431 ();
 sg13g2_decap_8 FILLER_30_1438 ();
 sg13g2_fill_2 FILLER_30_1445 ();
 sg13g2_fill_1 FILLER_30_1447 ();
 sg13g2_decap_8 FILLER_30_1474 ();
 sg13g2_decap_8 FILLER_30_1481 ();
 sg13g2_decap_8 FILLER_30_1488 ();
 sg13g2_decap_8 FILLER_30_1495 ();
 sg13g2_decap_8 FILLER_30_1502 ();
 sg13g2_decap_8 FILLER_30_1509 ();
 sg13g2_decap_8 FILLER_30_1516 ();
 sg13g2_decap_8 FILLER_30_1523 ();
 sg13g2_decap_8 FILLER_30_1535 ();
 sg13g2_decap_8 FILLER_30_1542 ();
 sg13g2_decap_8 FILLER_30_1549 ();
 sg13g2_decap_8 FILLER_30_1556 ();
 sg13g2_decap_8 FILLER_30_1563 ();
 sg13g2_decap_4 FILLER_30_1570 ();
 sg13g2_decap_8 FILLER_30_1584 ();
 sg13g2_decap_8 FILLER_30_1591 ();
 sg13g2_decap_8 FILLER_30_1598 ();
 sg13g2_decap_8 FILLER_30_1605 ();
 sg13g2_decap_8 FILLER_30_1612 ();
 sg13g2_decap_8 FILLER_30_1619 ();
 sg13g2_decap_8 FILLER_30_1626 ();
 sg13g2_decap_8 FILLER_30_1633 ();
 sg13g2_decap_8 FILLER_30_1640 ();
 sg13g2_decap_8 FILLER_30_1647 ();
 sg13g2_decap_8 FILLER_30_1654 ();
 sg13g2_fill_2 FILLER_30_1661 ();
 sg13g2_fill_1 FILLER_30_1663 ();
 sg13g2_decap_8 FILLER_30_1672 ();
 sg13g2_decap_8 FILLER_30_1679 ();
 sg13g2_decap_8 FILLER_30_1686 ();
 sg13g2_decap_8 FILLER_30_1693 ();
 sg13g2_decap_8 FILLER_30_1700 ();
 sg13g2_decap_8 FILLER_30_1707 ();
 sg13g2_decap_8 FILLER_30_1714 ();
 sg13g2_decap_8 FILLER_30_1721 ();
 sg13g2_decap_8 FILLER_30_1728 ();
 sg13g2_decap_4 FILLER_30_1735 ();
 sg13g2_decap_8 FILLER_30_1770 ();
 sg13g2_decap_4 FILLER_30_1777 ();
 sg13g2_fill_2 FILLER_30_1781 ();
 sg13g2_fill_2 FILLER_30_1799 ();
 sg13g2_fill_1 FILLER_30_1801 ();
 sg13g2_decap_8 FILLER_30_1807 ();
 sg13g2_decap_8 FILLER_30_1814 ();
 sg13g2_decap_8 FILLER_30_1821 ();
 sg13g2_decap_8 FILLER_30_1828 ();
 sg13g2_fill_1 FILLER_30_1835 ();
 sg13g2_fill_2 FILLER_30_1846 ();
 sg13g2_fill_1 FILLER_30_1848 ();
 sg13g2_decap_8 FILLER_30_1857 ();
 sg13g2_decap_8 FILLER_30_1864 ();
 sg13g2_decap_8 FILLER_30_1871 ();
 sg13g2_decap_4 FILLER_30_1878 ();
 sg13g2_fill_1 FILLER_30_1882 ();
 sg13g2_fill_2 FILLER_30_1901 ();
 sg13g2_fill_1 FILLER_30_1903 ();
 sg13g2_decap_4 FILLER_30_1919 ();
 sg13g2_decap_8 FILLER_30_1933 ();
 sg13g2_decap_8 FILLER_30_1940 ();
 sg13g2_fill_1 FILLER_30_1947 ();
 sg13g2_decap_8 FILLER_30_1952 ();
 sg13g2_fill_2 FILLER_30_1959 ();
 sg13g2_fill_1 FILLER_30_1961 ();
 sg13g2_decap_8 FILLER_30_1966 ();
 sg13g2_decap_8 FILLER_30_1973 ();
 sg13g2_decap_8 FILLER_30_1980 ();
 sg13g2_decap_8 FILLER_30_1987 ();
 sg13g2_decap_8 FILLER_30_1994 ();
 sg13g2_decap_8 FILLER_30_2001 ();
 sg13g2_fill_2 FILLER_30_2008 ();
 sg13g2_fill_1 FILLER_30_2036 ();
 sg13g2_fill_2 FILLER_30_2045 ();
 sg13g2_fill_1 FILLER_30_2047 ();
 sg13g2_fill_1 FILLER_30_2056 ();
 sg13g2_decap_8 FILLER_30_2073 ();
 sg13g2_decap_8 FILLER_30_2080 ();
 sg13g2_decap_8 FILLER_30_2087 ();
 sg13g2_decap_8 FILLER_30_2094 ();
 sg13g2_decap_8 FILLER_30_2101 ();
 sg13g2_decap_4 FILLER_30_2108 ();
 sg13g2_decap_8 FILLER_30_2124 ();
 sg13g2_fill_2 FILLER_30_2131 ();
 sg13g2_fill_1 FILLER_30_2133 ();
 sg13g2_decap_8 FILLER_30_2187 ();
 sg13g2_decap_8 FILLER_30_2194 ();
 sg13g2_fill_1 FILLER_30_2201 ();
 sg13g2_decap_8 FILLER_30_2208 ();
 sg13g2_decap_8 FILLER_30_2215 ();
 sg13g2_decap_8 FILLER_30_2222 ();
 sg13g2_decap_8 FILLER_30_2229 ();
 sg13g2_decap_8 FILLER_30_2236 ();
 sg13g2_fill_2 FILLER_30_2243 ();
 sg13g2_decap_8 FILLER_30_2262 ();
 sg13g2_decap_8 FILLER_30_2269 ();
 sg13g2_decap_8 FILLER_30_2284 ();
 sg13g2_decap_8 FILLER_30_2291 ();
 sg13g2_fill_1 FILLER_30_2298 ();
 sg13g2_fill_1 FILLER_30_2304 ();
 sg13g2_decap_8 FILLER_30_2313 ();
 sg13g2_decap_8 FILLER_30_2320 ();
 sg13g2_decap_8 FILLER_30_2327 ();
 sg13g2_decap_8 FILLER_30_2334 ();
 sg13g2_decap_8 FILLER_30_2341 ();
 sg13g2_decap_8 FILLER_30_2348 ();
 sg13g2_decap_8 FILLER_30_2355 ();
 sg13g2_decap_4 FILLER_30_2362 ();
 sg13g2_fill_1 FILLER_30_2366 ();
 sg13g2_decap_8 FILLER_30_2376 ();
 sg13g2_fill_1 FILLER_30_2383 ();
 sg13g2_decap_4 FILLER_30_2396 ();
 sg13g2_fill_1 FILLER_30_2400 ();
 sg13g2_decap_8 FILLER_30_2404 ();
 sg13g2_decap_4 FILLER_30_2411 ();
 sg13g2_fill_2 FILLER_30_2415 ();
 sg13g2_fill_2 FILLER_30_2430 ();
 sg13g2_decap_8 FILLER_30_2435 ();
 sg13g2_decap_8 FILLER_30_2442 ();
 sg13g2_decap_4 FILLER_30_2449 ();
 sg13g2_decap_8 FILLER_30_2470 ();
 sg13g2_decap_8 FILLER_30_2477 ();
 sg13g2_decap_8 FILLER_30_2484 ();
 sg13g2_decap_8 FILLER_30_2491 ();
 sg13g2_decap_8 FILLER_30_2498 ();
 sg13g2_decap_8 FILLER_30_2505 ();
 sg13g2_decap_8 FILLER_30_2512 ();
 sg13g2_decap_8 FILLER_30_2519 ();
 sg13g2_decap_8 FILLER_30_2526 ();
 sg13g2_decap_8 FILLER_30_2533 ();
 sg13g2_decap_8 FILLER_30_2540 ();
 sg13g2_decap_8 FILLER_30_2547 ();
 sg13g2_decap_8 FILLER_30_2554 ();
 sg13g2_decap_8 FILLER_30_2561 ();
 sg13g2_decap_8 FILLER_30_2568 ();
 sg13g2_decap_8 FILLER_30_2575 ();
 sg13g2_decap_8 FILLER_30_2582 ();
 sg13g2_decap_8 FILLER_30_2589 ();
 sg13g2_decap_8 FILLER_30_2596 ();
 sg13g2_decap_4 FILLER_30_2603 ();
 sg13g2_fill_2 FILLER_30_2618 ();
 sg13g2_fill_1 FILLER_30_2620 ();
 sg13g2_decap_8 FILLER_30_2626 ();
 sg13g2_decap_8 FILLER_30_2633 ();
 sg13g2_decap_8 FILLER_30_2640 ();
 sg13g2_decap_8 FILLER_30_2647 ();
 sg13g2_decap_8 FILLER_30_2654 ();
 sg13g2_decap_8 FILLER_30_2661 ();
 sg13g2_decap_8 FILLER_30_2668 ();
 sg13g2_decap_8 FILLER_30_2675 ();
 sg13g2_decap_8 FILLER_30_2692 ();
 sg13g2_decap_4 FILLER_30_2699 ();
 sg13g2_decap_8 FILLER_30_2708 ();
 sg13g2_decap_8 FILLER_30_2715 ();
 sg13g2_decap_4 FILLER_30_2722 ();
 sg13g2_decap_8 FILLER_30_2758 ();
 sg13g2_fill_1 FILLER_30_2765 ();
 sg13g2_decap_8 FILLER_30_2776 ();
 sg13g2_fill_2 FILLER_30_2783 ();
 sg13g2_fill_1 FILLER_30_2785 ();
 sg13g2_decap_8 FILLER_30_2796 ();
 sg13g2_decap_8 FILLER_30_2803 ();
 sg13g2_decap_8 FILLER_30_2810 ();
 sg13g2_decap_4 FILLER_30_2817 ();
 sg13g2_fill_1 FILLER_30_2821 ();
 sg13g2_decap_4 FILLER_30_2848 ();
 sg13g2_fill_2 FILLER_30_2852 ();
 sg13g2_decap_8 FILLER_30_2860 ();
 sg13g2_decap_8 FILLER_30_2867 ();
 sg13g2_decap_8 FILLER_30_2874 ();
 sg13g2_fill_2 FILLER_30_2881 ();
 sg13g2_fill_1 FILLER_30_2883 ();
 sg13g2_decap_4 FILLER_30_2936 ();
 sg13g2_fill_2 FILLER_30_2940 ();
 sg13g2_decap_8 FILLER_30_2947 ();
 sg13g2_decap_8 FILLER_30_2954 ();
 sg13g2_decap_8 FILLER_30_2961 ();
 sg13g2_decap_8 FILLER_30_2968 ();
 sg13g2_decap_8 FILLER_30_2975 ();
 sg13g2_decap_8 FILLER_30_2982 ();
 sg13g2_decap_4 FILLER_30_2989 ();
 sg13g2_fill_2 FILLER_30_3003 ();
 sg13g2_decap_8 FILLER_30_3031 ();
 sg13g2_fill_2 FILLER_30_3038 ();
 sg13g2_decap_8 FILLER_30_3066 ();
 sg13g2_decap_8 FILLER_30_3073 ();
 sg13g2_decap_8 FILLER_30_3080 ();
 sg13g2_decap_8 FILLER_30_3087 ();
 sg13g2_decap_8 FILLER_30_3094 ();
 sg13g2_decap_8 FILLER_30_3101 ();
 sg13g2_decap_4 FILLER_30_3108 ();
 sg13g2_decap_8 FILLER_30_3138 ();
 sg13g2_decap_8 FILLER_30_3145 ();
 sg13g2_decap_4 FILLER_30_3152 ();
 sg13g2_fill_2 FILLER_30_3156 ();
 sg13g2_decap_8 FILLER_30_3168 ();
 sg13g2_decap_8 FILLER_30_3175 ();
 sg13g2_decap_8 FILLER_30_3182 ();
 sg13g2_decap_8 FILLER_30_3189 ();
 sg13g2_decap_8 FILLER_30_3201 ();
 sg13g2_fill_2 FILLER_30_3208 ();
 sg13g2_decap_8 FILLER_30_3236 ();
 sg13g2_decap_8 FILLER_30_3243 ();
 sg13g2_decap_8 FILLER_30_3250 ();
 sg13g2_decap_8 FILLER_30_3257 ();
 sg13g2_decap_4 FILLER_30_3264 ();
 sg13g2_decap_8 FILLER_30_3278 ();
 sg13g2_decap_8 FILLER_30_3285 ();
 sg13g2_decap_8 FILLER_30_3292 ();
 sg13g2_decap_8 FILLER_30_3299 ();
 sg13g2_decap_8 FILLER_30_3306 ();
 sg13g2_decap_8 FILLER_30_3313 ();
 sg13g2_decap_8 FILLER_30_3320 ();
 sg13g2_decap_8 FILLER_30_3327 ();
 sg13g2_decap_8 FILLER_30_3334 ();
 sg13g2_fill_1 FILLER_30_3341 ();
 sg13g2_decap_8 FILLER_30_3348 ();
 sg13g2_decap_8 FILLER_30_3355 ();
 sg13g2_decap_8 FILLER_30_3362 ();
 sg13g2_decap_8 FILLER_30_3369 ();
 sg13g2_decap_8 FILLER_30_3376 ();
 sg13g2_decap_8 FILLER_30_3383 ();
 sg13g2_decap_8 FILLER_30_3390 ();
 sg13g2_decap_8 FILLER_30_3397 ();
 sg13g2_decap_8 FILLER_30_3404 ();
 sg13g2_decap_8 FILLER_30_3411 ();
 sg13g2_decap_8 FILLER_30_3418 ();
 sg13g2_decap_8 FILLER_30_3425 ();
 sg13g2_decap_8 FILLER_30_3432 ();
 sg13g2_fill_2 FILLER_30_3439 ();
 sg13g2_decap_8 FILLER_30_3446 ();
 sg13g2_decap_8 FILLER_30_3453 ();
 sg13g2_decap_8 FILLER_30_3460 ();
 sg13g2_decap_8 FILLER_30_3467 ();
 sg13g2_decap_8 FILLER_30_3474 ();
 sg13g2_decap_8 FILLER_30_3481 ();
 sg13g2_decap_8 FILLER_30_3488 ();
 sg13g2_decap_8 FILLER_30_3495 ();
 sg13g2_decap_8 FILLER_30_3502 ();
 sg13g2_decap_8 FILLER_30_3509 ();
 sg13g2_decap_8 FILLER_30_3516 ();
 sg13g2_fill_2 FILLER_30_3528 ();
 sg13g2_fill_1 FILLER_30_3530 ();
 sg13g2_decap_4 FILLER_30_3536 ();
 sg13g2_decap_8 FILLER_30_3550 ();
 sg13g2_decap_8 FILLER_30_3557 ();
 sg13g2_decap_8 FILLER_30_3564 ();
 sg13g2_decap_8 FILLER_30_3571 ();
 sg13g2_fill_2 FILLER_30_3578 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_4 FILLER_31_21 ();
 sg13g2_fill_2 FILLER_31_25 ();
 sg13g2_fill_2 FILLER_31_31 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_4 FILLER_31_77 ();
 sg13g2_fill_1 FILLER_31_81 ();
 sg13g2_decap_4 FILLER_31_103 ();
 sg13g2_decap_8 FILLER_31_119 ();
 sg13g2_decap_8 FILLER_31_126 ();
 sg13g2_decap_8 FILLER_31_133 ();
 sg13g2_decap_8 FILLER_31_140 ();
 sg13g2_fill_1 FILLER_31_147 ();
 sg13g2_fill_1 FILLER_31_156 ();
 sg13g2_decap_8 FILLER_31_170 ();
 sg13g2_decap_8 FILLER_31_177 ();
 sg13g2_decap_8 FILLER_31_184 ();
 sg13g2_decap_8 FILLER_31_199 ();
 sg13g2_decap_8 FILLER_31_206 ();
 sg13g2_decap_8 FILLER_31_213 ();
 sg13g2_fill_2 FILLER_31_220 ();
 sg13g2_fill_1 FILLER_31_227 ();
 sg13g2_decap_8 FILLER_31_246 ();
 sg13g2_decap_8 FILLER_31_253 ();
 sg13g2_decap_4 FILLER_31_260 ();
 sg13g2_fill_2 FILLER_31_264 ();
 sg13g2_decap_8 FILLER_31_282 ();
 sg13g2_decap_8 FILLER_31_289 ();
 sg13g2_decap_8 FILLER_31_296 ();
 sg13g2_fill_1 FILLER_31_303 ();
 sg13g2_fill_1 FILLER_31_310 ();
 sg13g2_decap_4 FILLER_31_316 ();
 sg13g2_decap_8 FILLER_31_328 ();
 sg13g2_decap_8 FILLER_31_335 ();
 sg13g2_decap_8 FILLER_31_342 ();
 sg13g2_decap_8 FILLER_31_349 ();
 sg13g2_decap_8 FILLER_31_356 ();
 sg13g2_decap_4 FILLER_31_363 ();
 sg13g2_fill_2 FILLER_31_367 ();
 sg13g2_decap_8 FILLER_31_380 ();
 sg13g2_decap_8 FILLER_31_391 ();
 sg13g2_decap_8 FILLER_31_398 ();
 sg13g2_decap_8 FILLER_31_405 ();
 sg13g2_decap_8 FILLER_31_412 ();
 sg13g2_decap_8 FILLER_31_419 ();
 sg13g2_fill_1 FILLER_31_432 ();
 sg13g2_fill_1 FILLER_31_455 ();
 sg13g2_decap_4 FILLER_31_464 ();
 sg13g2_fill_1 FILLER_31_468 ();
 sg13g2_fill_1 FILLER_31_478 ();
 sg13g2_fill_2 FILLER_31_488 ();
 sg13g2_fill_1 FILLER_31_502 ();
 sg13g2_decap_4 FILLER_31_519 ();
 sg13g2_fill_2 FILLER_31_523 ();
 sg13g2_fill_2 FILLER_31_538 ();
 sg13g2_decap_8 FILLER_31_548 ();
 sg13g2_decap_8 FILLER_31_555 ();
 sg13g2_decap_8 FILLER_31_562 ();
 sg13g2_decap_8 FILLER_31_569 ();
 sg13g2_decap_8 FILLER_31_576 ();
 sg13g2_decap_8 FILLER_31_583 ();
 sg13g2_decap_4 FILLER_31_590 ();
 sg13g2_fill_2 FILLER_31_594 ();
 sg13g2_decap_4 FILLER_31_608 ();
 sg13g2_fill_1 FILLER_31_612 ();
 sg13g2_decap_8 FILLER_31_625 ();
 sg13g2_decap_8 FILLER_31_632 ();
 sg13g2_decap_4 FILLER_31_639 ();
 sg13g2_fill_2 FILLER_31_643 ();
 sg13g2_decap_4 FILLER_31_655 ();
 sg13g2_fill_2 FILLER_31_659 ();
 sg13g2_decap_8 FILLER_31_686 ();
 sg13g2_decap_8 FILLER_31_693 ();
 sg13g2_decap_8 FILLER_31_700 ();
 sg13g2_decap_8 FILLER_31_707 ();
 sg13g2_decap_4 FILLER_31_714 ();
 sg13g2_fill_1 FILLER_31_723 ();
 sg13g2_decap_8 FILLER_31_747 ();
 sg13g2_decap_4 FILLER_31_754 ();
 sg13g2_fill_1 FILLER_31_758 ();
 sg13g2_decap_8 FILLER_31_795 ();
 sg13g2_decap_8 FILLER_31_847 ();
 sg13g2_decap_8 FILLER_31_854 ();
 sg13g2_decap_8 FILLER_31_861 ();
 sg13g2_fill_2 FILLER_31_868 ();
 sg13g2_decap_4 FILLER_31_906 ();
 sg13g2_fill_1 FILLER_31_910 ();
 sg13g2_decap_8 FILLER_31_917 ();
 sg13g2_decap_8 FILLER_31_924 ();
 sg13g2_decap_8 FILLER_31_931 ();
 sg13g2_decap_8 FILLER_31_938 ();
 sg13g2_decap_8 FILLER_31_945 ();
 sg13g2_decap_8 FILLER_31_952 ();
 sg13g2_decap_8 FILLER_31_959 ();
 sg13g2_fill_2 FILLER_31_966 ();
 sg13g2_decap_4 FILLER_31_978 ();
 sg13g2_decap_8 FILLER_31_992 ();
 sg13g2_decap_8 FILLER_31_999 ();
 sg13g2_decap_8 FILLER_31_1006 ();
 sg13g2_decap_8 FILLER_31_1013 ();
 sg13g2_decap_8 FILLER_31_1020 ();
 sg13g2_decap_8 FILLER_31_1053 ();
 sg13g2_decap_4 FILLER_31_1060 ();
 sg13g2_fill_1 FILLER_31_1064 ();
 sg13g2_decap_8 FILLER_31_1075 ();
 sg13g2_decap_8 FILLER_31_1082 ();
 sg13g2_decap_8 FILLER_31_1089 ();
 sg13g2_decap_8 FILLER_31_1096 ();
 sg13g2_decap_8 FILLER_31_1103 ();
 sg13g2_decap_4 FILLER_31_1110 ();
 sg13g2_decap_8 FILLER_31_1124 ();
 sg13g2_decap_8 FILLER_31_1131 ();
 sg13g2_decap_8 FILLER_31_1138 ();
 sg13g2_decap_8 FILLER_31_1145 ();
 sg13g2_decap_8 FILLER_31_1152 ();
 sg13g2_decap_8 FILLER_31_1159 ();
 sg13g2_decap_4 FILLER_31_1166 ();
 sg13g2_fill_2 FILLER_31_1170 ();
 sg13g2_decap_8 FILLER_31_1198 ();
 sg13g2_decap_8 FILLER_31_1205 ();
 sg13g2_decap_8 FILLER_31_1212 ();
 sg13g2_fill_2 FILLER_31_1219 ();
 sg13g2_fill_1 FILLER_31_1221 ();
 sg13g2_decap_8 FILLER_31_1240 ();
 sg13g2_decap_8 FILLER_31_1247 ();
 sg13g2_decap_8 FILLER_31_1254 ();
 sg13g2_decap_8 FILLER_31_1261 ();
 sg13g2_decap_8 FILLER_31_1268 ();
 sg13g2_decap_8 FILLER_31_1275 ();
 sg13g2_decap_8 FILLER_31_1282 ();
 sg13g2_decap_4 FILLER_31_1289 ();
 sg13g2_fill_2 FILLER_31_1293 ();
 sg13g2_decap_4 FILLER_31_1321 ();
 sg13g2_fill_1 FILLER_31_1325 ();
 sg13g2_decap_8 FILLER_31_1336 ();
 sg13g2_decap_8 FILLER_31_1343 ();
 sg13g2_decap_4 FILLER_31_1350 ();
 sg13g2_decap_8 FILLER_31_1385 ();
 sg13g2_fill_2 FILLER_31_1392 ();
 sg13g2_decap_8 FILLER_31_1430 ();
 sg13g2_decap_8 FILLER_31_1447 ();
 sg13g2_decap_8 FILLER_31_1454 ();
 sg13g2_decap_8 FILLER_31_1461 ();
 sg13g2_decap_8 FILLER_31_1468 ();
 sg13g2_decap_4 FILLER_31_1475 ();
 sg13g2_decap_8 FILLER_31_1491 ();
 sg13g2_decap_8 FILLER_31_1498 ();
 sg13g2_decap_8 FILLER_31_1505 ();
 sg13g2_decap_4 FILLER_31_1512 ();
 sg13g2_fill_1 FILLER_31_1516 ();
 sg13g2_decap_8 FILLER_31_1533 ();
 sg13g2_decap_8 FILLER_31_1540 ();
 sg13g2_decap_8 FILLER_31_1547 ();
 sg13g2_decap_8 FILLER_31_1554 ();
 sg13g2_decap_8 FILLER_31_1561 ();
 sg13g2_decap_8 FILLER_31_1568 ();
 sg13g2_fill_1 FILLER_31_1575 ();
 sg13g2_fill_2 FILLER_31_1585 ();
 sg13g2_fill_1 FILLER_31_1608 ();
 sg13g2_decap_8 FILLER_31_1626 ();
 sg13g2_decap_8 FILLER_31_1633 ();
 sg13g2_fill_2 FILLER_31_1640 ();
 sg13g2_fill_1 FILLER_31_1642 ();
 sg13g2_decap_8 FILLER_31_1653 ();
 sg13g2_decap_8 FILLER_31_1660 ();
 sg13g2_fill_1 FILLER_31_1667 ();
 sg13g2_decap_8 FILLER_31_1691 ();
 sg13g2_decap_8 FILLER_31_1698 ();
 sg13g2_decap_8 FILLER_31_1705 ();
 sg13g2_fill_1 FILLER_31_1712 ();
 sg13g2_decap_8 FILLER_31_1723 ();
 sg13g2_decap_8 FILLER_31_1730 ();
 sg13g2_decap_8 FILLER_31_1737 ();
 sg13g2_fill_2 FILLER_31_1744 ();
 sg13g2_fill_1 FILLER_31_1746 ();
 sg13g2_decap_8 FILLER_31_1785 ();
 sg13g2_fill_1 FILLER_31_1792 ();
 sg13g2_decap_8 FILLER_31_1813 ();
 sg13g2_decap_4 FILLER_31_1820 ();
 sg13g2_fill_2 FILLER_31_1824 ();
 sg13g2_decap_8 FILLER_31_1862 ();
 sg13g2_decap_8 FILLER_31_1869 ();
 sg13g2_decap_8 FILLER_31_1876 ();
 sg13g2_decap_8 FILLER_31_1915 ();
 sg13g2_decap_8 FILLER_31_1922 ();
 sg13g2_decap_8 FILLER_31_1929 ();
 sg13g2_decap_8 FILLER_31_1936 ();
 sg13g2_decap_8 FILLER_31_1943 ();
 sg13g2_decap_8 FILLER_31_1950 ();
 sg13g2_decap_8 FILLER_31_1957 ();
 sg13g2_decap_8 FILLER_31_1964 ();
 sg13g2_decap_8 FILLER_31_1971 ();
 sg13g2_decap_4 FILLER_31_1978 ();
 sg13g2_decap_8 FILLER_31_1996 ();
 sg13g2_decap_8 FILLER_31_2011 ();
 sg13g2_decap_8 FILLER_31_2018 ();
 sg13g2_decap_8 FILLER_31_2025 ();
 sg13g2_decap_8 FILLER_31_2032 ();
 sg13g2_fill_1 FILLER_31_2039 ();
 sg13g2_decap_8 FILLER_31_2060 ();
 sg13g2_decap_8 FILLER_31_2067 ();
 sg13g2_decap_8 FILLER_31_2074 ();
 sg13g2_decap_8 FILLER_31_2081 ();
 sg13g2_decap_8 FILLER_31_2088 ();
 sg13g2_decap_8 FILLER_31_2131 ();
 sg13g2_decap_4 FILLER_31_2138 ();
 sg13g2_fill_1 FILLER_31_2142 ();
 sg13g2_fill_1 FILLER_31_2158 ();
 sg13g2_decap_8 FILLER_31_2171 ();
 sg13g2_decap_8 FILLER_31_2178 ();
 sg13g2_decap_4 FILLER_31_2185 ();
 sg13g2_fill_2 FILLER_31_2200 ();
 sg13g2_decap_8 FILLER_31_2213 ();
 sg13g2_decap_8 FILLER_31_2220 ();
 sg13g2_decap_8 FILLER_31_2227 ();
 sg13g2_decap_8 FILLER_31_2234 ();
 sg13g2_decap_8 FILLER_31_2262 ();
 sg13g2_fill_1 FILLER_31_2269 ();
 sg13g2_decap_4 FILLER_31_2276 ();
 sg13g2_fill_1 FILLER_31_2280 ();
 sg13g2_decap_8 FILLER_31_2289 ();
 sg13g2_decap_8 FILLER_31_2296 ();
 sg13g2_decap_8 FILLER_31_2303 ();
 sg13g2_decap_8 FILLER_31_2310 ();
 sg13g2_decap_8 FILLER_31_2317 ();
 sg13g2_decap_8 FILLER_31_2324 ();
 sg13g2_decap_4 FILLER_31_2331 ();
 sg13g2_fill_1 FILLER_31_2335 ();
 sg13g2_decap_4 FILLER_31_2347 ();
 sg13g2_fill_1 FILLER_31_2362 ();
 sg13g2_fill_1 FILLER_31_2404 ();
 sg13g2_decap_8 FILLER_31_2422 ();
 sg13g2_fill_2 FILLER_31_2429 ();
 sg13g2_fill_1 FILLER_31_2431 ();
 sg13g2_decap_8 FILLER_31_2438 ();
 sg13g2_decap_8 FILLER_31_2445 ();
 sg13g2_decap_8 FILLER_31_2452 ();
 sg13g2_decap_8 FILLER_31_2459 ();
 sg13g2_decap_4 FILLER_31_2466 ();
 sg13g2_fill_1 FILLER_31_2470 ();
 sg13g2_decap_8 FILLER_31_2476 ();
 sg13g2_decap_4 FILLER_31_2483 ();
 sg13g2_fill_1 FILLER_31_2487 ();
 sg13g2_decap_8 FILLER_31_2494 ();
 sg13g2_decap_4 FILLER_31_2501 ();
 sg13g2_decap_8 FILLER_31_2510 ();
 sg13g2_decap_8 FILLER_31_2517 ();
 sg13g2_decap_8 FILLER_31_2524 ();
 sg13g2_decap_8 FILLER_31_2531 ();
 sg13g2_decap_4 FILLER_31_2538 ();
 sg13g2_fill_1 FILLER_31_2542 ();
 sg13g2_decap_8 FILLER_31_2548 ();
 sg13g2_decap_8 FILLER_31_2555 ();
 sg13g2_decap_8 FILLER_31_2562 ();
 sg13g2_decap_8 FILLER_31_2569 ();
 sg13g2_decap_8 FILLER_31_2576 ();
 sg13g2_decap_8 FILLER_31_2583 ();
 sg13g2_decap_8 FILLER_31_2590 ();
 sg13g2_decap_8 FILLER_31_2597 ();
 sg13g2_decap_8 FILLER_31_2604 ();
 sg13g2_decap_8 FILLER_31_2611 ();
 sg13g2_decap_4 FILLER_31_2624 ();
 sg13g2_fill_2 FILLER_31_2641 ();
 sg13g2_decap_8 FILLER_31_2654 ();
 sg13g2_decap_8 FILLER_31_2661 ();
 sg13g2_decap_8 FILLER_31_2668 ();
 sg13g2_fill_1 FILLER_31_2675 ();
 sg13g2_decap_8 FILLER_31_2702 ();
 sg13g2_decap_8 FILLER_31_2709 ();
 sg13g2_fill_2 FILLER_31_2716 ();
 sg13g2_fill_1 FILLER_31_2737 ();
 sg13g2_fill_1 FILLER_31_2744 ();
 sg13g2_decap_8 FILLER_31_2755 ();
 sg13g2_decap_8 FILLER_31_2762 ();
 sg13g2_decap_8 FILLER_31_2769 ();
 sg13g2_decap_4 FILLER_31_2776 ();
 sg13g2_decap_8 FILLER_31_2806 ();
 sg13g2_decap_4 FILLER_31_2813 ();
 sg13g2_fill_2 FILLER_31_2817 ();
 sg13g2_fill_1 FILLER_31_2847 ();
 sg13g2_fill_1 FILLER_31_2860 ();
 sg13g2_decap_8 FILLER_31_2872 ();
 sg13g2_decap_8 FILLER_31_2879 ();
 sg13g2_fill_2 FILLER_31_2886 ();
 sg13g2_decap_8 FILLER_31_2902 ();
 sg13g2_decap_8 FILLER_31_2909 ();
 sg13g2_decap_8 FILLER_31_2916 ();
 sg13g2_fill_2 FILLER_31_2923 ();
 sg13g2_fill_1 FILLER_31_2925 ();
 sg13g2_decap_8 FILLER_31_2962 ();
 sg13g2_decap_8 FILLER_31_2969 ();
 sg13g2_decap_4 FILLER_31_2976 ();
 sg13g2_fill_1 FILLER_31_2980 ();
 sg13g2_decap_8 FILLER_31_3017 ();
 sg13g2_decap_8 FILLER_31_3024 ();
 sg13g2_decap_8 FILLER_31_3031 ();
 sg13g2_decap_8 FILLER_31_3038 ();
 sg13g2_decap_8 FILLER_31_3045 ();
 sg13g2_decap_8 FILLER_31_3052 ();
 sg13g2_fill_1 FILLER_31_3059 ();
 sg13g2_fill_2 FILLER_31_3073 ();
 sg13g2_fill_1 FILLER_31_3075 ();
 sg13g2_decap_8 FILLER_31_3086 ();
 sg13g2_decap_4 FILLER_31_3093 ();
 sg13g2_decap_8 FILLER_31_3107 ();
 sg13g2_decap_8 FILLER_31_3114 ();
 sg13g2_decap_8 FILLER_31_3121 ();
 sg13g2_decap_8 FILLER_31_3128 ();
 sg13g2_fill_2 FILLER_31_3135 ();
 sg13g2_fill_1 FILLER_31_3137 ();
 sg13g2_decap_8 FILLER_31_3179 ();
 sg13g2_decap_8 FILLER_31_3186 ();
 sg13g2_decap_8 FILLER_31_3193 ();
 sg13g2_decap_8 FILLER_31_3200 ();
 sg13g2_decap_8 FILLER_31_3212 ();
 sg13g2_fill_2 FILLER_31_3219 ();
 sg13g2_fill_1 FILLER_31_3221 ();
 sg13g2_decap_8 FILLER_31_3232 ();
 sg13g2_decap_4 FILLER_31_3239 ();
 sg13g2_fill_2 FILLER_31_3243 ();
 sg13g2_decap_8 FILLER_31_3253 ();
 sg13g2_decap_4 FILLER_31_3260 ();
 sg13g2_decap_8 FILLER_31_3300 ();
 sg13g2_decap_8 FILLER_31_3307 ();
 sg13g2_decap_8 FILLER_31_3314 ();
 sg13g2_decap_8 FILLER_31_3321 ();
 sg13g2_decap_8 FILLER_31_3328 ();
 sg13g2_decap_4 FILLER_31_3335 ();
 sg13g2_fill_1 FILLER_31_3339 ();
 sg13g2_decap_8 FILLER_31_3366 ();
 sg13g2_decap_8 FILLER_31_3373 ();
 sg13g2_decap_4 FILLER_31_3380 ();
 sg13g2_fill_1 FILLER_31_3384 ();
 sg13g2_decap_8 FILLER_31_3411 ();
 sg13g2_decap_8 FILLER_31_3418 ();
 sg13g2_decap_4 FILLER_31_3425 ();
 sg13g2_fill_2 FILLER_31_3429 ();
 sg13g2_decap_8 FILLER_31_3457 ();
 sg13g2_decap_8 FILLER_31_3464 ();
 sg13g2_decap_8 FILLER_31_3471 ();
 sg13g2_decap_4 FILLER_31_3478 ();
 sg13g2_fill_1 FILLER_31_3482 ();
 sg13g2_fill_2 FILLER_31_3493 ();
 sg13g2_fill_1 FILLER_31_3495 ();
 sg13g2_decap_8 FILLER_31_3500 ();
 sg13g2_decap_8 FILLER_31_3512 ();
 sg13g2_decap_8 FILLER_31_3519 ();
 sg13g2_decap_8 FILLER_31_3526 ();
 sg13g2_decap_8 FILLER_31_3533 ();
 sg13g2_decap_8 FILLER_31_3540 ();
 sg13g2_decap_4 FILLER_31_3547 ();
 sg13g2_fill_2 FILLER_31_3551 ();
 sg13g2_decap_8 FILLER_31_3561 ();
 sg13g2_decap_8 FILLER_31_3568 ();
 sg13g2_decap_4 FILLER_31_3575 ();
 sg13g2_fill_1 FILLER_31_3579 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_fill_2 FILLER_32_21 ();
 sg13g2_fill_1 FILLER_32_23 ();
 sg13g2_fill_2 FILLER_32_42 ();
 sg13g2_fill_1 FILLER_32_44 ();
 sg13g2_decap_8 FILLER_32_50 ();
 sg13g2_decap_8 FILLER_32_57 ();
 sg13g2_decap_8 FILLER_32_64 ();
 sg13g2_decap_8 FILLER_32_71 ();
 sg13g2_decap_4 FILLER_32_78 ();
 sg13g2_fill_2 FILLER_32_82 ();
 sg13g2_decap_8 FILLER_32_92 ();
 sg13g2_decap_8 FILLER_32_99 ();
 sg13g2_decap_8 FILLER_32_106 ();
 sg13g2_decap_8 FILLER_32_113 ();
 sg13g2_decap_8 FILLER_32_120 ();
 sg13g2_decap_8 FILLER_32_127 ();
 sg13g2_decap_4 FILLER_32_134 ();
 sg13g2_decap_8 FILLER_32_179 ();
 sg13g2_fill_1 FILLER_32_186 ();
 sg13g2_decap_4 FILLER_32_203 ();
 sg13g2_fill_1 FILLER_32_213 ();
 sg13g2_fill_2 FILLER_32_233 ();
 sg13g2_fill_1 FILLER_32_243 ();
 sg13g2_decap_8 FILLER_32_249 ();
 sg13g2_decap_4 FILLER_32_256 ();
 sg13g2_fill_1 FILLER_32_260 ();
 sg13g2_decap_8 FILLER_32_279 ();
 sg13g2_decap_8 FILLER_32_286 ();
 sg13g2_decap_4 FILLER_32_293 ();
 sg13g2_fill_2 FILLER_32_297 ();
 sg13g2_decap_4 FILLER_32_302 ();
 sg13g2_decap_8 FILLER_32_332 ();
 sg13g2_decap_8 FILLER_32_339 ();
 sg13g2_decap_4 FILLER_32_346 ();
 sg13g2_fill_1 FILLER_32_390 ();
 sg13g2_decap_8 FILLER_32_400 ();
 sg13g2_decap_8 FILLER_32_407 ();
 sg13g2_decap_8 FILLER_32_418 ();
 sg13g2_decap_8 FILLER_32_425 ();
 sg13g2_decap_4 FILLER_32_432 ();
 sg13g2_decap_8 FILLER_32_446 ();
 sg13g2_decap_8 FILLER_32_453 ();
 sg13g2_decap_4 FILLER_32_460 ();
 sg13g2_fill_2 FILLER_32_464 ();
 sg13g2_fill_2 FILLER_32_479 ();
 sg13g2_fill_2 FILLER_32_485 ();
 sg13g2_decap_8 FILLER_32_495 ();
 sg13g2_decap_8 FILLER_32_502 ();
 sg13g2_decap_4 FILLER_32_509 ();
 sg13g2_fill_2 FILLER_32_513 ();
 sg13g2_decap_4 FILLER_32_530 ();
 sg13g2_decap_8 FILLER_32_551 ();
 sg13g2_decap_8 FILLER_32_558 ();
 sg13g2_decap_8 FILLER_32_565 ();
 sg13g2_decap_4 FILLER_32_572 ();
 sg13g2_fill_1 FILLER_32_576 ();
 sg13g2_decap_8 FILLER_32_590 ();
 sg13g2_decap_8 FILLER_32_597 ();
 sg13g2_decap_4 FILLER_32_604 ();
 sg13g2_fill_2 FILLER_32_608 ();
 sg13g2_decap_8 FILLER_32_623 ();
 sg13g2_decap_8 FILLER_32_630 ();
 sg13g2_decap_8 FILLER_32_637 ();
 sg13g2_decap_8 FILLER_32_644 ();
 sg13g2_decap_8 FILLER_32_651 ();
 sg13g2_fill_2 FILLER_32_658 ();
 sg13g2_fill_1 FILLER_32_660 ();
 sg13g2_decap_8 FILLER_32_683 ();
 sg13g2_decap_8 FILLER_32_690 ();
 sg13g2_decap_8 FILLER_32_697 ();
 sg13g2_decap_8 FILLER_32_704 ();
 sg13g2_decap_8 FILLER_32_711 ();
 sg13g2_decap_8 FILLER_32_718 ();
 sg13g2_decap_4 FILLER_32_725 ();
 sg13g2_fill_2 FILLER_32_729 ();
 sg13g2_decap_8 FILLER_32_743 ();
 sg13g2_decap_8 FILLER_32_750 ();
 sg13g2_decap_8 FILLER_32_757 ();
 sg13g2_fill_1 FILLER_32_764 ();
 sg13g2_decap_8 FILLER_32_801 ();
 sg13g2_decap_8 FILLER_32_808 ();
 sg13g2_decap_8 FILLER_32_815 ();
 sg13g2_decap_8 FILLER_32_822 ();
 sg13g2_decap_8 FILLER_32_855 ();
 sg13g2_decap_8 FILLER_32_862 ();
 sg13g2_fill_1 FILLER_32_869 ();
 sg13g2_fill_2 FILLER_32_880 ();
 sg13g2_fill_1 FILLER_32_882 ();
 sg13g2_fill_2 FILLER_32_909 ();
 sg13g2_decap_8 FILLER_32_924 ();
 sg13g2_fill_1 FILLER_32_931 ();
 sg13g2_decap_8 FILLER_32_942 ();
 sg13g2_decap_8 FILLER_32_949 ();
 sg13g2_decap_8 FILLER_32_956 ();
 sg13g2_decap_8 FILLER_32_963 ();
 sg13g2_decap_8 FILLER_32_970 ();
 sg13g2_fill_2 FILLER_32_977 ();
 sg13g2_fill_1 FILLER_32_979 ();
 sg13g2_decap_8 FILLER_32_1006 ();
 sg13g2_decap_8 FILLER_32_1013 ();
 sg13g2_decap_8 FILLER_32_1020 ();
 sg13g2_decap_8 FILLER_32_1027 ();
 sg13g2_decap_8 FILLER_32_1034 ();
 sg13g2_fill_1 FILLER_32_1041 ();
 sg13g2_decap_8 FILLER_32_1052 ();
 sg13g2_decap_8 FILLER_32_1059 ();
 sg13g2_decap_8 FILLER_32_1066 ();
 sg13g2_decap_8 FILLER_32_1073 ();
 sg13g2_decap_8 FILLER_32_1080 ();
 sg13g2_decap_8 FILLER_32_1087 ();
 sg13g2_decap_8 FILLER_32_1094 ();
 sg13g2_decap_8 FILLER_32_1101 ();
 sg13g2_decap_8 FILLER_32_1108 ();
 sg13g2_fill_2 FILLER_32_1121 ();
 sg13g2_fill_1 FILLER_32_1123 ();
 sg13g2_decap_8 FILLER_32_1150 ();
 sg13g2_decap_8 FILLER_32_1157 ();
 sg13g2_decap_4 FILLER_32_1164 ();
 sg13g2_fill_2 FILLER_32_1168 ();
 sg13g2_decap_8 FILLER_32_1180 ();
 sg13g2_decap_8 FILLER_32_1187 ();
 sg13g2_decap_8 FILLER_32_1194 ();
 sg13g2_decap_8 FILLER_32_1201 ();
 sg13g2_decap_8 FILLER_32_1208 ();
 sg13g2_decap_8 FILLER_32_1215 ();
 sg13g2_decap_8 FILLER_32_1222 ();
 sg13g2_fill_2 FILLER_32_1229 ();
 sg13g2_decap_8 FILLER_32_1241 ();
 sg13g2_decap_4 FILLER_32_1248 ();
 sg13g2_fill_1 FILLER_32_1252 ();
 sg13g2_decap_8 FILLER_32_1259 ();
 sg13g2_decap_8 FILLER_32_1266 ();
 sg13g2_decap_8 FILLER_32_1273 ();
 sg13g2_decap_8 FILLER_32_1280 ();
 sg13g2_decap_4 FILLER_32_1287 ();
 sg13g2_decap_4 FILLER_32_1317 ();
 sg13g2_fill_1 FILLER_32_1321 ();
 sg13g2_decap_8 FILLER_32_1348 ();
 sg13g2_decap_4 FILLER_32_1355 ();
 sg13g2_fill_1 FILLER_32_1359 ();
 sg13g2_fill_2 FILLER_32_1366 ();
 sg13g2_fill_1 FILLER_32_1368 ();
 sg13g2_decap_8 FILLER_32_1375 ();
 sg13g2_decap_8 FILLER_32_1382 ();
 sg13g2_decap_8 FILLER_32_1389 ();
 sg13g2_decap_8 FILLER_32_1396 ();
 sg13g2_decap_8 FILLER_32_1433 ();
 sg13g2_decap_8 FILLER_32_1440 ();
 sg13g2_decap_8 FILLER_32_1447 ();
 sg13g2_fill_2 FILLER_32_1454 ();
 sg13g2_decap_8 FILLER_32_1482 ();
 sg13g2_decap_8 FILLER_32_1489 ();
 sg13g2_decap_8 FILLER_32_1496 ();
 sg13g2_decap_8 FILLER_32_1503 ();
 sg13g2_decap_4 FILLER_32_1510 ();
 sg13g2_fill_1 FILLER_32_1514 ();
 sg13g2_decap_8 FILLER_32_1552 ();
 sg13g2_decap_8 FILLER_32_1559 ();
 sg13g2_fill_2 FILLER_32_1566 ();
 sg13g2_decap_8 FILLER_32_1593 ();
 sg13g2_fill_2 FILLER_32_1600 ();
 sg13g2_fill_1 FILLER_32_1602 ();
 sg13g2_decap_8 FILLER_32_1609 ();
 sg13g2_decap_8 FILLER_32_1616 ();
 sg13g2_fill_2 FILLER_32_1623 ();
 sg13g2_decap_8 FILLER_32_1631 ();
 sg13g2_decap_4 FILLER_32_1638 ();
 sg13g2_decap_4 FILLER_32_1668 ();
 sg13g2_fill_1 FILLER_32_1672 ();
 sg13g2_decap_8 FILLER_32_1709 ();
 sg13g2_fill_2 FILLER_32_1716 ();
 sg13g2_fill_1 FILLER_32_1718 ();
 sg13g2_decap_8 FILLER_32_1725 ();
 sg13g2_decap_8 FILLER_32_1732 ();
 sg13g2_decap_8 FILLER_32_1739 ();
 sg13g2_decap_8 FILLER_32_1746 ();
 sg13g2_decap_8 FILLER_32_1753 ();
 sg13g2_decap_8 FILLER_32_1760 ();
 sg13g2_fill_2 FILLER_32_1767 ();
 sg13g2_decap_8 FILLER_32_1774 ();
 sg13g2_decap_8 FILLER_32_1781 ();
 sg13g2_decap_8 FILLER_32_1788 ();
 sg13g2_decap_8 FILLER_32_1795 ();
 sg13g2_decap_4 FILLER_32_1802 ();
 sg13g2_decap_4 FILLER_32_1810 ();
 sg13g2_fill_2 FILLER_32_1814 ();
 sg13g2_decap_8 FILLER_32_1820 ();
 sg13g2_decap_4 FILLER_32_1827 ();
 sg13g2_decap_8 FILLER_32_1841 ();
 sg13g2_fill_1 FILLER_32_1848 ();
 sg13g2_decap_8 FILLER_32_1855 ();
 sg13g2_decap_8 FILLER_32_1862 ();
 sg13g2_fill_2 FILLER_32_1869 ();
 sg13g2_fill_1 FILLER_32_1871 ();
 sg13g2_decap_8 FILLER_32_1878 ();
 sg13g2_decap_8 FILLER_32_1885 ();
 sg13g2_decap_8 FILLER_32_1895 ();
 sg13g2_decap_8 FILLER_32_1902 ();
 sg13g2_decap_4 FILLER_32_1909 ();
 sg13g2_fill_2 FILLER_32_1913 ();
 sg13g2_decap_8 FILLER_32_1929 ();
 sg13g2_decap_8 FILLER_32_1936 ();
 sg13g2_decap_8 FILLER_32_1943 ();
 sg13g2_fill_1 FILLER_32_1950 ();
 sg13g2_fill_1 FILLER_32_1977 ();
 sg13g2_decap_4 FILLER_32_1990 ();
 sg13g2_fill_2 FILLER_32_1994 ();
 sg13g2_decap_8 FILLER_32_2010 ();
 sg13g2_decap_8 FILLER_32_2017 ();
 sg13g2_decap_8 FILLER_32_2024 ();
 sg13g2_decap_8 FILLER_32_2031 ();
 sg13g2_decap_8 FILLER_32_2038 ();
 sg13g2_fill_2 FILLER_32_2045 ();
 sg13g2_fill_1 FILLER_32_2047 ();
 sg13g2_decap_4 FILLER_32_2063 ();
 sg13g2_decap_8 FILLER_32_2121 ();
 sg13g2_decap_8 FILLER_32_2128 ();
 sg13g2_decap_8 FILLER_32_2135 ();
 sg13g2_decap_8 FILLER_32_2142 ();
 sg13g2_decap_8 FILLER_32_2149 ();
 sg13g2_decap_8 FILLER_32_2156 ();
 sg13g2_decap_8 FILLER_32_2169 ();
 sg13g2_decap_8 FILLER_32_2176 ();
 sg13g2_decap_4 FILLER_32_2183 ();
 sg13g2_fill_2 FILLER_32_2187 ();
 sg13g2_decap_8 FILLER_32_2207 ();
 sg13g2_decap_8 FILLER_32_2219 ();
 sg13g2_decap_8 FILLER_32_2226 ();
 sg13g2_decap_4 FILLER_32_2233 ();
 sg13g2_decap_8 FILLER_32_2268 ();
 sg13g2_decap_8 FILLER_32_2275 ();
 sg13g2_decap_8 FILLER_32_2282 ();
 sg13g2_decap_8 FILLER_32_2289 ();
 sg13g2_decap_8 FILLER_32_2296 ();
 sg13g2_decap_8 FILLER_32_2303 ();
 sg13g2_decap_8 FILLER_32_2310 ();
 sg13g2_fill_2 FILLER_32_2317 ();
 sg13g2_decap_8 FILLER_32_2324 ();
 sg13g2_fill_2 FILLER_32_2331 ();
 sg13g2_fill_1 FILLER_32_2333 ();
 sg13g2_decap_8 FILLER_32_2354 ();
 sg13g2_decap_8 FILLER_32_2361 ();
 sg13g2_fill_2 FILLER_32_2368 ();
 sg13g2_decap_4 FILLER_32_2394 ();
 sg13g2_fill_1 FILLER_32_2398 ();
 sg13g2_decap_8 FILLER_32_2405 ();
 sg13g2_decap_8 FILLER_32_2412 ();
 sg13g2_decap_8 FILLER_32_2419 ();
 sg13g2_decap_8 FILLER_32_2426 ();
 sg13g2_decap_8 FILLER_32_2433 ();
 sg13g2_fill_2 FILLER_32_2440 ();
 sg13g2_decap_8 FILLER_32_2450 ();
 sg13g2_decap_8 FILLER_32_2457 ();
 sg13g2_fill_2 FILLER_32_2470 ();
 sg13g2_fill_1 FILLER_32_2472 ();
 sg13g2_fill_2 FILLER_32_2478 ();
 sg13g2_fill_1 FILLER_32_2480 ();
 sg13g2_fill_1 FILLER_32_2494 ();
 sg13g2_decap_4 FILLER_32_2504 ();
 sg13g2_fill_2 FILLER_32_2521 ();
 sg13g2_decap_4 FILLER_32_2529 ();
 sg13g2_fill_2 FILLER_32_2533 ();
 sg13g2_decap_4 FILLER_32_2558 ();
 sg13g2_fill_1 FILLER_32_2568 ();
 sg13g2_fill_2 FILLER_32_2587 ();
 sg13g2_fill_1 FILLER_32_2589 ();
 sg13g2_decap_8 FILLER_32_2595 ();
 sg13g2_decap_8 FILLER_32_2602 ();
 sg13g2_decap_4 FILLER_32_2609 ();
 sg13g2_decap_8 FILLER_32_2631 ();
 sg13g2_decap_8 FILLER_32_2664 ();
 sg13g2_decap_8 FILLER_32_2671 ();
 sg13g2_decap_8 FILLER_32_2678 ();
 sg13g2_decap_8 FILLER_32_2685 ();
 sg13g2_decap_8 FILLER_32_2692 ();
 sg13g2_decap_8 FILLER_32_2699 ();
 sg13g2_decap_8 FILLER_32_2706 ();
 sg13g2_decap_8 FILLER_32_2713 ();
 sg13g2_decap_8 FILLER_32_2720 ();
 sg13g2_decap_4 FILLER_32_2727 ();
 sg13g2_decap_8 FILLER_32_2736 ();
 sg13g2_decap_8 FILLER_32_2743 ();
 sg13g2_decap_8 FILLER_32_2750 ();
 sg13g2_decap_8 FILLER_32_2757 ();
 sg13g2_decap_8 FILLER_32_2764 ();
 sg13g2_decap_8 FILLER_32_2771 ();
 sg13g2_decap_8 FILLER_32_2778 ();
 sg13g2_decap_8 FILLER_32_2785 ();
 sg13g2_decap_8 FILLER_32_2792 ();
 sg13g2_decap_8 FILLER_32_2799 ();
 sg13g2_decap_8 FILLER_32_2806 ();
 sg13g2_decap_4 FILLER_32_2813 ();
 sg13g2_decap_8 FILLER_32_2822 ();
 sg13g2_decap_8 FILLER_32_2829 ();
 sg13g2_fill_1 FILLER_32_2836 ();
 sg13g2_fill_2 FILLER_32_2846 ();
 sg13g2_fill_1 FILLER_32_2853 ();
 sg13g2_decap_8 FILLER_32_2860 ();
 sg13g2_decap_8 FILLER_32_2867 ();
 sg13g2_decap_8 FILLER_32_2874 ();
 sg13g2_decap_8 FILLER_32_2881 ();
 sg13g2_decap_8 FILLER_32_2888 ();
 sg13g2_decap_8 FILLER_32_2895 ();
 sg13g2_decap_8 FILLER_32_2902 ();
 sg13g2_decap_8 FILLER_32_2909 ();
 sg13g2_decap_8 FILLER_32_2916 ();
 sg13g2_decap_8 FILLER_32_2923 ();
 sg13g2_decap_8 FILLER_32_2930 ();
 sg13g2_decap_4 FILLER_32_2937 ();
 sg13g2_fill_1 FILLER_32_2946 ();
 sg13g2_decap_8 FILLER_32_2962 ();
 sg13g2_decap_8 FILLER_32_2969 ();
 sg13g2_decap_8 FILLER_32_2976 ();
 sg13g2_decap_8 FILLER_32_2983 ();
 sg13g2_decap_8 FILLER_32_2990 ();
 sg13g2_decap_8 FILLER_32_2997 ();
 sg13g2_decap_8 FILLER_32_3004 ();
 sg13g2_decap_8 FILLER_32_3011 ();
 sg13g2_decap_8 FILLER_32_3018 ();
 sg13g2_decap_8 FILLER_32_3025 ();
 sg13g2_decap_8 FILLER_32_3032 ();
 sg13g2_decap_4 FILLER_32_3039 ();
 sg13g2_fill_2 FILLER_32_3043 ();
 sg13g2_decap_8 FILLER_32_3070 ();
 sg13g2_decap_4 FILLER_32_3077 ();
 sg13g2_decap_8 FILLER_32_3107 ();
 sg13g2_decap_8 FILLER_32_3114 ();
 sg13g2_decap_8 FILLER_32_3121 ();
 sg13g2_decap_8 FILLER_32_3128 ();
 sg13g2_decap_8 FILLER_32_3135 ();
 sg13g2_decap_8 FILLER_32_3142 ();
 sg13g2_decap_8 FILLER_32_3149 ();
 sg13g2_fill_1 FILLER_32_3156 ();
 sg13g2_fill_2 FILLER_32_3165 ();
 sg13g2_decap_8 FILLER_32_3193 ();
 sg13g2_decap_8 FILLER_32_3200 ();
 sg13g2_decap_8 FILLER_32_3207 ();
 sg13g2_decap_8 FILLER_32_3214 ();
 sg13g2_decap_8 FILLER_32_3231 ();
 sg13g2_decap_8 FILLER_32_3238 ();
 sg13g2_decap_8 FILLER_32_3245 ();
 sg13g2_decap_8 FILLER_32_3252 ();
 sg13g2_decap_4 FILLER_32_3259 ();
 sg13g2_fill_2 FILLER_32_3263 ();
 sg13g2_decap_8 FILLER_32_3291 ();
 sg13g2_decap_8 FILLER_32_3298 ();
 sg13g2_decap_8 FILLER_32_3305 ();
 sg13g2_decap_8 FILLER_32_3312 ();
 sg13g2_decap_8 FILLER_32_3319 ();
 sg13g2_fill_1 FILLER_32_3326 ();
 sg13g2_decap_8 FILLER_32_3363 ();
 sg13g2_decap_4 FILLER_32_3370 ();
 sg13g2_fill_2 FILLER_32_3374 ();
 sg13g2_decap_8 FILLER_32_3412 ();
 sg13g2_decap_8 FILLER_32_3419 ();
 sg13g2_fill_2 FILLER_32_3426 ();
 sg13g2_fill_1 FILLER_32_3428 ();
 sg13g2_decap_8 FILLER_32_3465 ();
 sg13g2_decap_8 FILLER_32_3472 ();
 sg13g2_decap_8 FILLER_32_3499 ();
 sg13g2_decap_8 FILLER_32_3506 ();
 sg13g2_decap_4 FILLER_32_3513 ();
 sg13g2_decap_8 FILLER_32_3562 ();
 sg13g2_decap_8 FILLER_32_3569 ();
 sg13g2_decap_4 FILLER_32_3576 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_fill_2 FILLER_33_33 ();
 sg13g2_fill_1 FILLER_33_45 ();
 sg13g2_decap_4 FILLER_33_50 ();
 sg13g2_decap_8 FILLER_33_59 ();
 sg13g2_decap_8 FILLER_33_66 ();
 sg13g2_decap_8 FILLER_33_73 ();
 sg13g2_decap_8 FILLER_33_83 ();
 sg13g2_fill_2 FILLER_33_90 ();
 sg13g2_decap_8 FILLER_33_105 ();
 sg13g2_decap_8 FILLER_33_117 ();
 sg13g2_decap_8 FILLER_33_124 ();
 sg13g2_decap_8 FILLER_33_131 ();
 sg13g2_decap_8 FILLER_33_138 ();
 sg13g2_decap_4 FILLER_33_145 ();
 sg13g2_fill_1 FILLER_33_149 ();
 sg13g2_fill_1 FILLER_33_165 ();
 sg13g2_decap_8 FILLER_33_175 ();
 sg13g2_decap_8 FILLER_33_182 ();
 sg13g2_decap_8 FILLER_33_189 ();
 sg13g2_fill_2 FILLER_33_207 ();
 sg13g2_fill_2 FILLER_33_255 ();
 sg13g2_fill_2 FILLER_33_263 ();
 sg13g2_fill_1 FILLER_33_265 ();
 sg13g2_decap_8 FILLER_33_271 ();
 sg13g2_fill_2 FILLER_33_278 ();
 sg13g2_fill_1 FILLER_33_280 ();
 sg13g2_fill_2 FILLER_33_287 ();
 sg13g2_fill_1 FILLER_33_306 ();
 sg13g2_decap_4 FILLER_33_311 ();
 sg13g2_fill_1 FILLER_33_318 ();
 sg13g2_decap_8 FILLER_33_339 ();
 sg13g2_decap_8 FILLER_33_346 ();
 sg13g2_decap_8 FILLER_33_353 ();
 sg13g2_decap_8 FILLER_33_360 ();
 sg13g2_decap_8 FILLER_33_367 ();
 sg13g2_decap_8 FILLER_33_374 ();
 sg13g2_fill_2 FILLER_33_381 ();
 sg13g2_decap_8 FILLER_33_388 ();
 sg13g2_decap_8 FILLER_33_395 ();
 sg13g2_decap_8 FILLER_33_402 ();
 sg13g2_decap_8 FILLER_33_409 ();
 sg13g2_fill_2 FILLER_33_416 ();
 sg13g2_fill_1 FILLER_33_418 ();
 sg13g2_decap_4 FILLER_33_424 ();
 sg13g2_fill_2 FILLER_33_428 ();
 sg13g2_fill_2 FILLER_33_443 ();
 sg13g2_fill_1 FILLER_33_445 ();
 sg13g2_fill_1 FILLER_33_456 ();
 sg13g2_decap_8 FILLER_33_465 ();
 sg13g2_decap_8 FILLER_33_472 ();
 sg13g2_decap_8 FILLER_33_479 ();
 sg13g2_decap_8 FILLER_33_486 ();
 sg13g2_decap_8 FILLER_33_493 ();
 sg13g2_decap_8 FILLER_33_500 ();
 sg13g2_decap_8 FILLER_33_507 ();
 sg13g2_decap_8 FILLER_33_514 ();
 sg13g2_decap_8 FILLER_33_521 ();
 sg13g2_decap_8 FILLER_33_528 ();
 sg13g2_decap_8 FILLER_33_535 ();
 sg13g2_decap_8 FILLER_33_542 ();
 sg13g2_decap_8 FILLER_33_549 ();
 sg13g2_decap_8 FILLER_33_556 ();
 sg13g2_decap_8 FILLER_33_563 ();
 sg13g2_decap_8 FILLER_33_570 ();
 sg13g2_decap_8 FILLER_33_577 ();
 sg13g2_decap_8 FILLER_33_584 ();
 sg13g2_decap_8 FILLER_33_591 ();
 sg13g2_decap_4 FILLER_33_598 ();
 sg13g2_fill_2 FILLER_33_632 ();
 sg13g2_decap_8 FILLER_33_639 ();
 sg13g2_decap_8 FILLER_33_646 ();
 sg13g2_decap_8 FILLER_33_653 ();
 sg13g2_decap_8 FILLER_33_660 ();
 sg13g2_decap_8 FILLER_33_667 ();
 sg13g2_decap_8 FILLER_33_674 ();
 sg13g2_decap_8 FILLER_33_681 ();
 sg13g2_decap_8 FILLER_33_688 ();
 sg13g2_decap_8 FILLER_33_695 ();
 sg13g2_decap_8 FILLER_33_702 ();
 sg13g2_decap_8 FILLER_33_709 ();
 sg13g2_decap_8 FILLER_33_716 ();
 sg13g2_decap_8 FILLER_33_723 ();
 sg13g2_decap_8 FILLER_33_730 ();
 sg13g2_decap_8 FILLER_33_737 ();
 sg13g2_decap_8 FILLER_33_744 ();
 sg13g2_decap_8 FILLER_33_751 ();
 sg13g2_decap_8 FILLER_33_758 ();
 sg13g2_decap_8 FILLER_33_765 ();
 sg13g2_decap_8 FILLER_33_772 ();
 sg13g2_decap_8 FILLER_33_779 ();
 sg13g2_decap_8 FILLER_33_786 ();
 sg13g2_decap_8 FILLER_33_793 ();
 sg13g2_decap_8 FILLER_33_800 ();
 sg13g2_decap_8 FILLER_33_807 ();
 sg13g2_decap_8 FILLER_33_814 ();
 sg13g2_decap_8 FILLER_33_821 ();
 sg13g2_decap_8 FILLER_33_838 ();
 sg13g2_decap_8 FILLER_33_845 ();
 sg13g2_decap_8 FILLER_33_852 ();
 sg13g2_fill_2 FILLER_33_859 ();
 sg13g2_fill_1 FILLER_33_861 ();
 sg13g2_decap_8 FILLER_33_872 ();
 sg13g2_decap_8 FILLER_33_879 ();
 sg13g2_decap_8 FILLER_33_886 ();
 sg13g2_decap_8 FILLER_33_893 ();
 sg13g2_decap_8 FILLER_33_900 ();
 sg13g2_decap_8 FILLER_33_907 ();
 sg13g2_decap_8 FILLER_33_917 ();
 sg13g2_decap_8 FILLER_33_924 ();
 sg13g2_decap_8 FILLER_33_931 ();
 sg13g2_fill_2 FILLER_33_938 ();
 sg13g2_fill_1 FILLER_33_940 ();
 sg13g2_decap_8 FILLER_33_967 ();
 sg13g2_decap_8 FILLER_33_974 ();
 sg13g2_fill_1 FILLER_33_981 ();
 sg13g2_decap_8 FILLER_33_1018 ();
 sg13g2_decap_8 FILLER_33_1025 ();
 sg13g2_decap_8 FILLER_33_1032 ();
 sg13g2_decap_8 FILLER_33_1039 ();
 sg13g2_decap_8 FILLER_33_1046 ();
 sg13g2_decap_4 FILLER_33_1053 ();
 sg13g2_decap_8 FILLER_33_1061 ();
 sg13g2_decap_8 FILLER_33_1068 ();
 sg13g2_decap_4 FILLER_33_1075 ();
 sg13g2_fill_1 FILLER_33_1079 ();
 sg13g2_decap_8 FILLER_33_1090 ();
 sg13g2_decap_8 FILLER_33_1097 ();
 sg13g2_decap_8 FILLER_33_1104 ();
 sg13g2_fill_1 FILLER_33_1111 ();
 sg13g2_decap_8 FILLER_33_1151 ();
 sg13g2_decap_8 FILLER_33_1158 ();
 sg13g2_decap_8 FILLER_33_1165 ();
 sg13g2_decap_8 FILLER_33_1172 ();
 sg13g2_decap_8 FILLER_33_1179 ();
 sg13g2_decap_8 FILLER_33_1186 ();
 sg13g2_decap_8 FILLER_33_1193 ();
 sg13g2_decap_8 FILLER_33_1200 ();
 sg13g2_decap_8 FILLER_33_1207 ();
 sg13g2_decap_8 FILLER_33_1214 ();
 sg13g2_decap_4 FILLER_33_1221 ();
 sg13g2_fill_2 FILLER_33_1225 ();
 sg13g2_decap_8 FILLER_33_1269 ();
 sg13g2_decap_8 FILLER_33_1276 ();
 sg13g2_decap_8 FILLER_33_1283 ();
 sg13g2_fill_2 FILLER_33_1290 ();
 sg13g2_decap_8 FILLER_33_1302 ();
 sg13g2_decap_8 FILLER_33_1309 ();
 sg13g2_decap_8 FILLER_33_1316 ();
 sg13g2_decap_4 FILLER_33_1323 ();
 sg13g2_fill_2 FILLER_33_1327 ();
 sg13g2_decap_8 FILLER_33_1339 ();
 sg13g2_decap_8 FILLER_33_1346 ();
 sg13g2_fill_1 FILLER_33_1353 ();
 sg13g2_decap_8 FILLER_33_1360 ();
 sg13g2_decap_8 FILLER_33_1367 ();
 sg13g2_decap_8 FILLER_33_1374 ();
 sg13g2_decap_8 FILLER_33_1381 ();
 sg13g2_decap_8 FILLER_33_1388 ();
 sg13g2_decap_8 FILLER_33_1395 ();
 sg13g2_decap_4 FILLER_33_1402 ();
 sg13g2_fill_2 FILLER_33_1406 ();
 sg13g2_decap_8 FILLER_33_1411 ();
 sg13g2_decap_4 FILLER_33_1418 ();
 sg13g2_decap_4 FILLER_33_1428 ();
 sg13g2_fill_1 FILLER_33_1432 ();
 sg13g2_decap_8 FILLER_33_1441 ();
 sg13g2_decap_8 FILLER_33_1458 ();
 sg13g2_fill_1 FILLER_33_1465 ();
 sg13g2_decap_8 FILLER_33_1498 ();
 sg13g2_decap_8 FILLER_33_1505 ();
 sg13g2_decap_8 FILLER_33_1512 ();
 sg13g2_decap_4 FILLER_33_1519 ();
 sg13g2_fill_1 FILLER_33_1523 ();
 sg13g2_decap_8 FILLER_33_1550 ();
 sg13g2_decap_8 FILLER_33_1557 ();
 sg13g2_decap_4 FILLER_33_1564 ();
 sg13g2_decap_8 FILLER_33_1600 ();
 sg13g2_decap_8 FILLER_33_1607 ();
 sg13g2_decap_8 FILLER_33_1614 ();
 sg13g2_decap_8 FILLER_33_1621 ();
 sg13g2_decap_8 FILLER_33_1628 ();
 sg13g2_decap_8 FILLER_33_1635 ();
 sg13g2_decap_8 FILLER_33_1642 ();
 sg13g2_decap_8 FILLER_33_1649 ();
 sg13g2_decap_8 FILLER_33_1656 ();
 sg13g2_decap_8 FILLER_33_1663 ();
 sg13g2_decap_8 FILLER_33_1670 ();
 sg13g2_fill_2 FILLER_33_1677 ();
 sg13g2_decap_8 FILLER_33_1705 ();
 sg13g2_decap_4 FILLER_33_1712 ();
 sg13g2_fill_1 FILLER_33_1716 ();
 sg13g2_decap_8 FILLER_33_1727 ();
 sg13g2_decap_8 FILLER_33_1734 ();
 sg13g2_decap_8 FILLER_33_1741 ();
 sg13g2_decap_4 FILLER_33_1748 ();
 sg13g2_fill_2 FILLER_33_1752 ();
 sg13g2_decap_8 FILLER_33_1760 ();
 sg13g2_decap_8 FILLER_33_1767 ();
 sg13g2_decap_8 FILLER_33_1774 ();
 sg13g2_decap_8 FILLER_33_1781 ();
 sg13g2_decap_4 FILLER_33_1788 ();
 sg13g2_fill_1 FILLER_33_1792 ();
 sg13g2_decap_8 FILLER_33_1799 ();
 sg13g2_decap_4 FILLER_33_1806 ();
 sg13g2_decap_8 FILLER_33_1816 ();
 sg13g2_decap_8 FILLER_33_1823 ();
 sg13g2_decap_8 FILLER_33_1830 ();
 sg13g2_decap_8 FILLER_33_1837 ();
 sg13g2_decap_8 FILLER_33_1844 ();
 sg13g2_decap_8 FILLER_33_1851 ();
 sg13g2_decap_8 FILLER_33_1858 ();
 sg13g2_decap_8 FILLER_33_1865 ();
 sg13g2_decap_4 FILLER_33_1872 ();
 sg13g2_fill_1 FILLER_33_1876 ();
 sg13g2_fill_1 FILLER_33_1899 ();
 sg13g2_decap_8 FILLER_33_1910 ();
 sg13g2_decap_8 FILLER_33_1917 ();
 sg13g2_decap_8 FILLER_33_1924 ();
 sg13g2_decap_8 FILLER_33_1931 ();
 sg13g2_fill_2 FILLER_33_1938 ();
 sg13g2_decap_8 FILLER_33_1958 ();
 sg13g2_decap_8 FILLER_33_1965 ();
 sg13g2_decap_8 FILLER_33_1972 ();
 sg13g2_decap_8 FILLER_33_1979 ();
 sg13g2_decap_8 FILLER_33_1986 ();
 sg13g2_decap_8 FILLER_33_2021 ();
 sg13g2_decap_8 FILLER_33_2028 ();
 sg13g2_decap_8 FILLER_33_2035 ();
 sg13g2_decap_8 FILLER_33_2042 ();
 sg13g2_decap_8 FILLER_33_2049 ();
 sg13g2_decap_8 FILLER_33_2056 ();
 sg13g2_decap_8 FILLER_33_2063 ();
 sg13g2_fill_2 FILLER_33_2070 ();
 sg13g2_fill_1 FILLER_33_2072 ();
 sg13g2_decap_8 FILLER_33_2079 ();
 sg13g2_decap_8 FILLER_33_2086 ();
 sg13g2_decap_8 FILLER_33_2093 ();
 sg13g2_fill_1 FILLER_33_2100 ();
 sg13g2_decap_8 FILLER_33_2107 ();
 sg13g2_decap_8 FILLER_33_2114 ();
 sg13g2_decap_8 FILLER_33_2121 ();
 sg13g2_decap_8 FILLER_33_2128 ();
 sg13g2_decap_4 FILLER_33_2135 ();
 sg13g2_fill_2 FILLER_33_2145 ();
 sg13g2_fill_1 FILLER_33_2147 ();
 sg13g2_decap_8 FILLER_33_2178 ();
 sg13g2_decap_8 FILLER_33_2185 ();
 sg13g2_fill_2 FILLER_33_2192 ();
 sg13g2_decap_4 FILLER_33_2202 ();
 sg13g2_decap_8 FILLER_33_2212 ();
 sg13g2_decap_8 FILLER_33_2219 ();
 sg13g2_decap_8 FILLER_33_2226 ();
 sg13g2_decap_8 FILLER_33_2233 ();
 sg13g2_decap_8 FILLER_33_2240 ();
 sg13g2_fill_1 FILLER_33_2247 ();
 sg13g2_decap_8 FILLER_33_2262 ();
 sg13g2_fill_2 FILLER_33_2269 ();
 sg13g2_fill_1 FILLER_33_2271 ();
 sg13g2_decap_4 FILLER_33_2278 ();
 sg13g2_fill_1 FILLER_33_2282 ();
 sg13g2_decap_8 FILLER_33_2294 ();
 sg13g2_decap_4 FILLER_33_2301 ();
 sg13g2_decap_8 FILLER_33_2311 ();
 sg13g2_decap_8 FILLER_33_2318 ();
 sg13g2_decap_8 FILLER_33_2325 ();
 sg13g2_decap_8 FILLER_33_2332 ();
 sg13g2_fill_2 FILLER_33_2339 ();
 sg13g2_fill_1 FILLER_33_2341 ();
 sg13g2_decap_8 FILLER_33_2347 ();
 sg13g2_decap_8 FILLER_33_2354 ();
 sg13g2_decap_8 FILLER_33_2361 ();
 sg13g2_decap_8 FILLER_33_2368 ();
 sg13g2_decap_8 FILLER_33_2375 ();
 sg13g2_decap_8 FILLER_33_2382 ();
 sg13g2_decap_8 FILLER_33_2389 ();
 sg13g2_decap_4 FILLER_33_2396 ();
 sg13g2_fill_1 FILLER_33_2400 ();
 sg13g2_decap_8 FILLER_33_2407 ();
 sg13g2_decap_8 FILLER_33_2414 ();
 sg13g2_decap_8 FILLER_33_2421 ();
 sg13g2_decap_4 FILLER_33_2442 ();
 sg13g2_fill_1 FILLER_33_2452 ();
 sg13g2_decap_4 FILLER_33_2463 ();
 sg13g2_fill_2 FILLER_33_2467 ();
 sg13g2_decap_4 FILLER_33_2474 ();
 sg13g2_fill_1 FILLER_33_2478 ();
 sg13g2_fill_1 FILLER_33_2486 ();
 sg13g2_decap_8 FILLER_33_2498 ();
 sg13g2_decap_8 FILLER_33_2505 ();
 sg13g2_fill_1 FILLER_33_2512 ();
 sg13g2_fill_1 FILLER_33_2520 ();
 sg13g2_decap_8 FILLER_33_2543 ();
 sg13g2_decap_8 FILLER_33_2550 ();
 sg13g2_fill_1 FILLER_33_2557 ();
 sg13g2_fill_2 FILLER_33_2585 ();
 sg13g2_fill_1 FILLER_33_2587 ();
 sg13g2_decap_4 FILLER_33_2600 ();
 sg13g2_fill_1 FILLER_33_2604 ();
 sg13g2_decap_4 FILLER_33_2614 ();
 sg13g2_decap_8 FILLER_33_2628 ();
 sg13g2_decap_8 FILLER_33_2635 ();
 sg13g2_decap_8 FILLER_33_2642 ();
 sg13g2_decap_8 FILLER_33_2649 ();
 sg13g2_decap_8 FILLER_33_2656 ();
 sg13g2_fill_2 FILLER_33_2663 ();
 sg13g2_fill_1 FILLER_33_2665 ();
 sg13g2_decap_4 FILLER_33_2674 ();
 sg13g2_decap_8 FILLER_33_2696 ();
 sg13g2_decap_8 FILLER_33_2703 ();
 sg13g2_fill_1 FILLER_33_2710 ();
 sg13g2_decap_8 FILLER_33_2721 ();
 sg13g2_decap_8 FILLER_33_2728 ();
 sg13g2_decap_8 FILLER_33_2735 ();
 sg13g2_decap_8 FILLER_33_2742 ();
 sg13g2_decap_8 FILLER_33_2749 ();
 sg13g2_decap_4 FILLER_33_2756 ();
 sg13g2_fill_2 FILLER_33_2760 ();
 sg13g2_decap_8 FILLER_33_2766 ();
 sg13g2_decap_8 FILLER_33_2773 ();
 sg13g2_decap_8 FILLER_33_2780 ();
 sg13g2_decap_8 FILLER_33_2787 ();
 sg13g2_decap_4 FILLER_33_2794 ();
 sg13g2_fill_1 FILLER_33_2798 ();
 sg13g2_fill_1 FILLER_33_2809 ();
 sg13g2_decap_8 FILLER_33_2815 ();
 sg13g2_decap_8 FILLER_33_2822 ();
 sg13g2_fill_2 FILLER_33_2829 ();
 sg13g2_decap_8 FILLER_33_2842 ();
 sg13g2_decap_8 FILLER_33_2849 ();
 sg13g2_decap_8 FILLER_33_2864 ();
 sg13g2_decap_8 FILLER_33_2871 ();
 sg13g2_decap_8 FILLER_33_2878 ();
 sg13g2_decap_8 FILLER_33_2885 ();
 sg13g2_decap_8 FILLER_33_2892 ();
 sg13g2_decap_8 FILLER_33_2899 ();
 sg13g2_decap_8 FILLER_33_2906 ();
 sg13g2_decap_8 FILLER_33_2913 ();
 sg13g2_decap_4 FILLER_33_2920 ();
 sg13g2_fill_1 FILLER_33_2924 ();
 sg13g2_decap_8 FILLER_33_2930 ();
 sg13g2_decap_8 FILLER_33_2937 ();
 sg13g2_decap_4 FILLER_33_2944 ();
 sg13g2_fill_1 FILLER_33_2948 ();
 sg13g2_fill_1 FILLER_33_2975 ();
 sg13g2_decap_8 FILLER_33_2986 ();
 sg13g2_decap_8 FILLER_33_2993 ();
 sg13g2_decap_8 FILLER_33_3000 ();
 sg13g2_decap_8 FILLER_33_3007 ();
 sg13g2_decap_8 FILLER_33_3014 ();
 sg13g2_fill_2 FILLER_33_3021 ();
 sg13g2_decap_8 FILLER_33_3033 ();
 sg13g2_decap_8 FILLER_33_3040 ();
 sg13g2_decap_8 FILLER_33_3047 ();
 sg13g2_decap_8 FILLER_33_3054 ();
 sg13g2_decap_8 FILLER_33_3061 ();
 sg13g2_decap_8 FILLER_33_3068 ();
 sg13g2_decap_8 FILLER_33_3075 ();
 sg13g2_decap_8 FILLER_33_3082 ();
 sg13g2_decap_8 FILLER_33_3089 ();
 sg13g2_decap_4 FILLER_33_3096 ();
 sg13g2_fill_2 FILLER_33_3100 ();
 sg13g2_decap_8 FILLER_33_3128 ();
 sg13g2_decap_8 FILLER_33_3135 ();
 sg13g2_decap_8 FILLER_33_3142 ();
 sg13g2_decap_8 FILLER_33_3149 ();
 sg13g2_decap_8 FILLER_33_3156 ();
 sg13g2_decap_4 FILLER_33_3163 ();
 sg13g2_decap_8 FILLER_33_3177 ();
 sg13g2_decap_8 FILLER_33_3184 ();
 sg13g2_decap_8 FILLER_33_3191 ();
 sg13g2_decap_8 FILLER_33_3198 ();
 sg13g2_decap_8 FILLER_33_3205 ();
 sg13g2_fill_1 FILLER_33_3212 ();
 sg13g2_decap_8 FILLER_33_3239 ();
 sg13g2_decap_8 FILLER_33_3246 ();
 sg13g2_decap_8 FILLER_33_3253 ();
 sg13g2_decap_8 FILLER_33_3260 ();
 sg13g2_fill_2 FILLER_33_3267 ();
 sg13g2_decap_8 FILLER_33_3273 ();
 sg13g2_decap_8 FILLER_33_3280 ();
 sg13g2_decap_8 FILLER_33_3287 ();
 sg13g2_decap_4 FILLER_33_3294 ();
 sg13g2_fill_1 FILLER_33_3298 ();
 sg13g2_fill_2 FILLER_33_3335 ();
 sg13g2_fill_1 FILLER_33_3347 ();
 sg13g2_decap_8 FILLER_33_3351 ();
 sg13g2_decap_8 FILLER_33_3358 ();
 sg13g2_decap_8 FILLER_33_3365 ();
 sg13g2_decap_8 FILLER_33_3372 ();
 sg13g2_decap_4 FILLER_33_3379 ();
 sg13g2_fill_2 FILLER_33_3383 ();
 sg13g2_decap_8 FILLER_33_3395 ();
 sg13g2_decap_8 FILLER_33_3402 ();
 sg13g2_decap_8 FILLER_33_3409 ();
 sg13g2_decap_8 FILLER_33_3416 ();
 sg13g2_decap_8 FILLER_33_3423 ();
 sg13g2_decap_4 FILLER_33_3430 ();
 sg13g2_fill_1 FILLER_33_3434 ();
 sg13g2_decap_8 FILLER_33_3460 ();
 sg13g2_decap_8 FILLER_33_3467 ();
 sg13g2_decap_8 FILLER_33_3474 ();
 sg13g2_fill_1 FILLER_33_3486 ();
 sg13g2_decap_8 FILLER_33_3501 ();
 sg13g2_decap_8 FILLER_33_3508 ();
 sg13g2_fill_1 FILLER_33_3515 ();
 sg13g2_fill_2 FILLER_33_3521 ();
 sg13g2_fill_2 FILLER_33_3528 ();
 sg13g2_decap_8 FILLER_33_3563 ();
 sg13g2_decap_8 FILLER_33_3570 ();
 sg13g2_fill_2 FILLER_33_3577 ();
 sg13g2_fill_1 FILLER_33_3579 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_4 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_27 ();
 sg13g2_fill_2 FILLER_34_34 ();
 sg13g2_decap_8 FILLER_34_59 ();
 sg13g2_decap_8 FILLER_34_66 ();
 sg13g2_decap_8 FILLER_34_73 ();
 sg13g2_decap_8 FILLER_34_80 ();
 sg13g2_decap_8 FILLER_34_87 ();
 sg13g2_decap_8 FILLER_34_94 ();
 sg13g2_fill_2 FILLER_34_101 ();
 sg13g2_fill_1 FILLER_34_103 ();
 sg13g2_decap_4 FILLER_34_114 ();
 sg13g2_fill_1 FILLER_34_118 ();
 sg13g2_decap_8 FILLER_34_127 ();
 sg13g2_decap_8 FILLER_34_134 ();
 sg13g2_decap_8 FILLER_34_141 ();
 sg13g2_decap_8 FILLER_34_148 ();
 sg13g2_fill_1 FILLER_34_160 ();
 sg13g2_decap_8 FILLER_34_178 ();
 sg13g2_decap_8 FILLER_34_185 ();
 sg13g2_decap_8 FILLER_34_192 ();
 sg13g2_decap_4 FILLER_34_199 ();
 sg13g2_decap_4 FILLER_34_208 ();
 sg13g2_fill_1 FILLER_34_212 ();
 sg13g2_fill_1 FILLER_34_218 ();
 sg13g2_decap_4 FILLER_34_228 ();
 sg13g2_fill_1 FILLER_34_232 ();
 sg13g2_decap_8 FILLER_34_243 ();
 sg13g2_decap_8 FILLER_34_250 ();
 sg13g2_decap_8 FILLER_34_257 ();
 sg13g2_decap_8 FILLER_34_264 ();
 sg13g2_decap_8 FILLER_34_271 ();
 sg13g2_decap_8 FILLER_34_278 ();
 sg13g2_decap_4 FILLER_34_285 ();
 sg13g2_fill_1 FILLER_34_315 ();
 sg13g2_decap_8 FILLER_34_325 ();
 sg13g2_decap_8 FILLER_34_332 ();
 sg13g2_fill_2 FILLER_34_339 ();
 sg13g2_decap_8 FILLER_34_354 ();
 sg13g2_decap_8 FILLER_34_361 ();
 sg13g2_decap_8 FILLER_34_368 ();
 sg13g2_fill_2 FILLER_34_375 ();
 sg13g2_fill_1 FILLER_34_377 ();
 sg13g2_fill_2 FILLER_34_404 ();
 sg13g2_fill_1 FILLER_34_406 ();
 sg13g2_decap_8 FILLER_34_415 ();
 sg13g2_fill_2 FILLER_34_422 ();
 sg13g2_fill_2 FILLER_34_439 ();
 sg13g2_fill_1 FILLER_34_441 ();
 sg13g2_decap_8 FILLER_34_461 ();
 sg13g2_decap_8 FILLER_34_468 ();
 sg13g2_decap_8 FILLER_34_475 ();
 sg13g2_decap_8 FILLER_34_482 ();
 sg13g2_decap_8 FILLER_34_489 ();
 sg13g2_decap_8 FILLER_34_496 ();
 sg13g2_decap_8 FILLER_34_503 ();
 sg13g2_decap_8 FILLER_34_510 ();
 sg13g2_decap_8 FILLER_34_517 ();
 sg13g2_decap_8 FILLER_34_524 ();
 sg13g2_decap_8 FILLER_34_531 ();
 sg13g2_decap_8 FILLER_34_538 ();
 sg13g2_decap_8 FILLER_34_545 ();
 sg13g2_decap_8 FILLER_34_552 ();
 sg13g2_decap_8 FILLER_34_559 ();
 sg13g2_decap_8 FILLER_34_566 ();
 sg13g2_decap_8 FILLER_34_573 ();
 sg13g2_decap_8 FILLER_34_580 ();
 sg13g2_decap_8 FILLER_34_587 ();
 sg13g2_decap_4 FILLER_34_594 ();
 sg13g2_fill_2 FILLER_34_598 ();
 sg13g2_fill_1 FILLER_34_637 ();
 sg13g2_decap_8 FILLER_34_651 ();
 sg13g2_decap_8 FILLER_34_658 ();
 sg13g2_decap_8 FILLER_34_665 ();
 sg13g2_fill_2 FILLER_34_672 ();
 sg13g2_fill_1 FILLER_34_674 ();
 sg13g2_decap_4 FILLER_34_696 ();
 sg13g2_fill_1 FILLER_34_705 ();
 sg13g2_decap_8 FILLER_34_709 ();
 sg13g2_fill_1 FILLER_34_716 ();
 sg13g2_decap_8 FILLER_34_727 ();
 sg13g2_decap_8 FILLER_34_734 ();
 sg13g2_fill_2 FILLER_34_741 ();
 sg13g2_fill_1 FILLER_34_743 ();
 sg13g2_decap_8 FILLER_34_749 ();
 sg13g2_decap_8 FILLER_34_756 ();
 sg13g2_decap_8 FILLER_34_763 ();
 sg13g2_decap_8 FILLER_34_770 ();
 sg13g2_decap_8 FILLER_34_777 ();
 sg13g2_decap_8 FILLER_34_784 ();
 sg13g2_decap_8 FILLER_34_791 ();
 sg13g2_decap_8 FILLER_34_798 ();
 sg13g2_decap_8 FILLER_34_805 ();
 sg13g2_decap_8 FILLER_34_812 ();
 sg13g2_decap_8 FILLER_34_819 ();
 sg13g2_decap_8 FILLER_34_826 ();
 sg13g2_fill_1 FILLER_34_833 ();
 sg13g2_decap_8 FILLER_34_842 ();
 sg13g2_fill_1 FILLER_34_849 ();
 sg13g2_decap_8 FILLER_34_853 ();
 sg13g2_decap_8 FILLER_34_860 ();
 sg13g2_decap_4 FILLER_34_867 ();
 sg13g2_decap_8 FILLER_34_897 ();
 sg13g2_decap_8 FILLER_34_904 ();
 sg13g2_decap_4 FILLER_34_911 ();
 sg13g2_decap_8 FILLER_34_941 ();
 sg13g2_decap_8 FILLER_34_948 ();
 sg13g2_decap_8 FILLER_34_955 ();
 sg13g2_decap_8 FILLER_34_962 ();
 sg13g2_decap_8 FILLER_34_969 ();
 sg13g2_decap_8 FILLER_34_976 ();
 sg13g2_decap_8 FILLER_34_983 ();
 sg13g2_decap_8 FILLER_34_990 ();
 sg13g2_decap_8 FILLER_34_997 ();
 sg13g2_decap_8 FILLER_34_1004 ();
 sg13g2_decap_8 FILLER_34_1011 ();
 sg13g2_decap_8 FILLER_34_1018 ();
 sg13g2_decap_8 FILLER_34_1025 ();
 sg13g2_decap_4 FILLER_34_1032 ();
 sg13g2_fill_2 FILLER_34_1036 ();
 sg13g2_fill_2 FILLER_34_1057 ();
 sg13g2_fill_1 FILLER_34_1059 ();
 sg13g2_decap_8 FILLER_34_1096 ();
 sg13g2_decap_8 FILLER_34_1103 ();
 sg13g2_decap_8 FILLER_34_1110 ();
 sg13g2_decap_8 FILLER_34_1117 ();
 sg13g2_decap_8 FILLER_34_1124 ();
 sg13g2_decap_8 FILLER_34_1131 ();
 sg13g2_decap_8 FILLER_34_1138 ();
 sg13g2_decap_8 FILLER_34_1145 ();
 sg13g2_decap_8 FILLER_34_1152 ();
 sg13g2_fill_1 FILLER_34_1159 ();
 sg13g2_decap_8 FILLER_34_1196 ();
 sg13g2_decap_8 FILLER_34_1203 ();
 sg13g2_decap_8 FILLER_34_1210 ();
 sg13g2_decap_8 FILLER_34_1217 ();
 sg13g2_decap_8 FILLER_34_1224 ();
 sg13g2_decap_8 FILLER_34_1231 ();
 sg13g2_fill_2 FILLER_34_1238 ();
 sg13g2_fill_1 FILLER_34_1240 ();
 sg13g2_fill_1 FILLER_34_1244 ();
 sg13g2_fill_2 FILLER_34_1254 ();
 sg13g2_decap_8 FILLER_34_1295 ();
 sg13g2_decap_8 FILLER_34_1302 ();
 sg13g2_decap_8 FILLER_34_1309 ();
 sg13g2_decap_8 FILLER_34_1316 ();
 sg13g2_decap_4 FILLER_34_1323 ();
 sg13g2_fill_1 FILLER_34_1327 ();
 sg13g2_decap_8 FILLER_34_1333 ();
 sg13g2_decap_8 FILLER_34_1340 ();
 sg13g2_decap_4 FILLER_34_1347 ();
 sg13g2_fill_2 FILLER_34_1351 ();
 sg13g2_decap_4 FILLER_34_1359 ();
 sg13g2_decap_8 FILLER_34_1407 ();
 sg13g2_decap_8 FILLER_34_1414 ();
 sg13g2_decap_8 FILLER_34_1421 ();
 sg13g2_decap_8 FILLER_34_1428 ();
 sg13g2_decap_8 FILLER_34_1435 ();
 sg13g2_decap_8 FILLER_34_1442 ();
 sg13g2_decap_8 FILLER_34_1449 ();
 sg13g2_decap_8 FILLER_34_1456 ();
 sg13g2_decap_8 FILLER_34_1463 ();
 sg13g2_fill_1 FILLER_34_1470 ();
 sg13g2_decap_8 FILLER_34_1481 ();
 sg13g2_decap_4 FILLER_34_1488 ();
 sg13g2_decap_8 FILLER_34_1503 ();
 sg13g2_decap_8 FILLER_34_1510 ();
 sg13g2_decap_4 FILLER_34_1517 ();
 sg13g2_fill_2 FILLER_34_1521 ();
 sg13g2_decap_8 FILLER_34_1543 ();
 sg13g2_decap_8 FILLER_34_1550 ();
 sg13g2_decap_8 FILLER_34_1557 ();
 sg13g2_decap_8 FILLER_34_1564 ();
 sg13g2_decap_8 FILLER_34_1571 ();
 sg13g2_decap_4 FILLER_34_1578 ();
 sg13g2_decap_4 FILLER_34_1590 ();
 sg13g2_fill_2 FILLER_34_1594 ();
 sg13g2_decap_8 FILLER_34_1602 ();
 sg13g2_decap_4 FILLER_34_1609 ();
 sg13g2_fill_2 FILLER_34_1613 ();
 sg13g2_decap_8 FILLER_34_1628 ();
 sg13g2_decap_4 FILLER_34_1635 ();
 sg13g2_fill_2 FILLER_34_1639 ();
 sg13g2_decap_8 FILLER_34_1662 ();
 sg13g2_fill_2 FILLER_34_1669 ();
 sg13g2_fill_1 FILLER_34_1671 ();
 sg13g2_decap_8 FILLER_34_1682 ();
 sg13g2_decap_8 FILLER_34_1689 ();
 sg13g2_decap_8 FILLER_34_1696 ();
 sg13g2_decap_4 FILLER_34_1703 ();
 sg13g2_fill_1 FILLER_34_1707 ();
 sg13g2_decap_8 FILLER_34_1740 ();
 sg13g2_decap_8 FILLER_34_1757 ();
 sg13g2_decap_8 FILLER_34_1764 ();
 sg13g2_decap_8 FILLER_34_1771 ();
 sg13g2_fill_1 FILLER_34_1778 ();
 sg13g2_fill_2 FILLER_34_1815 ();
 sg13g2_fill_1 FILLER_34_1817 ();
 sg13g2_decap_8 FILLER_34_1828 ();
 sg13g2_decap_8 FILLER_34_1861 ();
 sg13g2_decap_8 FILLER_34_1868 ();
 sg13g2_decap_8 FILLER_34_1875 ();
 sg13g2_decap_4 FILLER_34_1882 ();
 sg13g2_decap_4 FILLER_34_1924 ();
 sg13g2_fill_2 FILLER_34_1928 ();
 sg13g2_decap_8 FILLER_34_1969 ();
 sg13g2_decap_8 FILLER_34_1976 ();
 sg13g2_decap_8 FILLER_34_1983 ();
 sg13g2_decap_8 FILLER_34_1990 ();
 sg13g2_decap_8 FILLER_34_1997 ();
 sg13g2_decap_8 FILLER_34_2004 ();
 sg13g2_decap_4 FILLER_34_2011 ();
 sg13g2_decap_4 FILLER_34_2020 ();
 sg13g2_fill_1 FILLER_34_2024 ();
 sg13g2_fill_2 FILLER_34_2033 ();
 sg13g2_fill_2 FILLER_34_2045 ();
 sg13g2_fill_2 FILLER_34_2073 ();
 sg13g2_fill_1 FILLER_34_2075 ();
 sg13g2_decap_8 FILLER_34_2091 ();
 sg13g2_decap_8 FILLER_34_2098 ();
 sg13g2_decap_4 FILLER_34_2105 ();
 sg13g2_fill_2 FILLER_34_2109 ();
 sg13g2_decap_8 FILLER_34_2115 ();
 sg13g2_fill_2 FILLER_34_2122 ();
 sg13g2_fill_1 FILLER_34_2124 ();
 sg13g2_decap_8 FILLER_34_2131 ();
 sg13g2_decap_8 FILLER_34_2138 ();
 sg13g2_decap_8 FILLER_34_2145 ();
 sg13g2_decap_8 FILLER_34_2152 ();
 sg13g2_decap_8 FILLER_34_2159 ();
 sg13g2_decap_8 FILLER_34_2166 ();
 sg13g2_decap_4 FILLER_34_2173 ();
 sg13g2_fill_2 FILLER_34_2207 ();
 sg13g2_fill_1 FILLER_34_2218 ();
 sg13g2_decap_8 FILLER_34_2236 ();
 sg13g2_fill_2 FILLER_34_2243 ();
 sg13g2_fill_1 FILLER_34_2250 ();
 sg13g2_decap_8 FILLER_34_2257 ();
 sg13g2_fill_2 FILLER_34_2264 ();
 sg13g2_fill_1 FILLER_34_2266 ();
 sg13g2_fill_1 FILLER_34_2275 ();
 sg13g2_fill_2 FILLER_34_2282 ();
 sg13g2_fill_1 FILLER_34_2284 ();
 sg13g2_fill_2 FILLER_34_2297 ();
 sg13g2_fill_1 FILLER_34_2299 ();
 sg13g2_fill_1 FILLER_34_2320 ();
 sg13g2_decap_4 FILLER_34_2347 ();
 sg13g2_decap_4 FILLER_34_2357 ();
 sg13g2_decap_4 FILLER_34_2375 ();
 sg13g2_fill_1 FILLER_34_2379 ();
 sg13g2_decap_8 FILLER_34_2388 ();
 sg13g2_fill_2 FILLER_34_2401 ();
 sg13g2_fill_1 FILLER_34_2403 ();
 sg13g2_decap_8 FILLER_34_2418 ();
 sg13g2_decap_8 FILLER_34_2425 ();
 sg13g2_fill_1 FILLER_34_2432 ();
 sg13g2_decap_8 FILLER_34_2439 ();
 sg13g2_decap_4 FILLER_34_2446 ();
 sg13g2_decap_8 FILLER_34_2478 ();
 sg13g2_decap_8 FILLER_34_2485 ();
 sg13g2_fill_2 FILLER_34_2492 ();
 sg13g2_fill_1 FILLER_34_2494 ();
 sg13g2_decap_8 FILLER_34_2501 ();
 sg13g2_decap_8 FILLER_34_2508 ();
 sg13g2_fill_1 FILLER_34_2515 ();
 sg13g2_decap_8 FILLER_34_2527 ();
 sg13g2_decap_8 FILLER_34_2534 ();
 sg13g2_fill_2 FILLER_34_2541 ();
 sg13g2_decap_8 FILLER_34_2549 ();
 sg13g2_decap_4 FILLER_34_2556 ();
 sg13g2_fill_1 FILLER_34_2560 ();
 sg13g2_fill_2 FILLER_34_2567 ();
 sg13g2_fill_1 FILLER_34_2569 ();
 sg13g2_decap_8 FILLER_34_2575 ();
 sg13g2_fill_2 FILLER_34_2582 ();
 sg13g2_fill_1 FILLER_34_2613 ();
 sg13g2_decap_8 FILLER_34_2619 ();
 sg13g2_decap_8 FILLER_34_2626 ();
 sg13g2_decap_8 FILLER_34_2633 ();
 sg13g2_decap_8 FILLER_34_2643 ();
 sg13g2_decap_8 FILLER_34_2650 ();
 sg13g2_decap_8 FILLER_34_2657 ();
 sg13g2_fill_2 FILLER_34_2664 ();
 sg13g2_decap_8 FILLER_34_2695 ();
 sg13g2_decap_4 FILLER_34_2702 ();
 sg13g2_fill_2 FILLER_34_2706 ();
 sg13g2_decap_8 FILLER_34_2768 ();
 sg13g2_fill_1 FILLER_34_2775 ();
 sg13g2_decap_4 FILLER_34_2788 ();
 sg13g2_fill_2 FILLER_34_2792 ();
 sg13g2_decap_8 FILLER_34_2820 ();
 sg13g2_decap_8 FILLER_34_2827 ();
 sg13g2_decap_8 FILLER_34_2834 ();
 sg13g2_decap_8 FILLER_34_2841 ();
 sg13g2_decap_8 FILLER_34_2848 ();
 sg13g2_fill_2 FILLER_34_2855 ();
 sg13g2_fill_1 FILLER_34_2867 ();
 sg13g2_decap_8 FILLER_34_2894 ();
 sg13g2_decap_8 FILLER_34_2901 ();
 sg13g2_fill_1 FILLER_34_2908 ();
 sg13g2_fill_1 FILLER_34_2914 ();
 sg13g2_decap_8 FILLER_34_2936 ();
 sg13g2_decap_8 FILLER_34_2943 ();
 sg13g2_decap_8 FILLER_34_2950 ();
 sg13g2_decap_4 FILLER_34_2957 ();
 sg13g2_decap_8 FILLER_34_2966 ();
 sg13g2_decap_8 FILLER_34_2973 ();
 sg13g2_fill_2 FILLER_34_2980 ();
 sg13g2_decap_8 FILLER_34_3008 ();
 sg13g2_decap_8 FILLER_34_3015 ();
 sg13g2_decap_4 FILLER_34_3022 ();
 sg13g2_fill_1 FILLER_34_3026 ();
 sg13g2_decap_8 FILLER_34_3061 ();
 sg13g2_decap_8 FILLER_34_3068 ();
 sg13g2_decap_8 FILLER_34_3075 ();
 sg13g2_decap_8 FILLER_34_3082 ();
 sg13g2_decap_8 FILLER_34_3089 ();
 sg13g2_decap_8 FILLER_34_3096 ();
 sg13g2_decap_8 FILLER_34_3103 ();
 sg13g2_decap_8 FILLER_34_3110 ();
 sg13g2_decap_8 FILLER_34_3117 ();
 sg13g2_decap_8 FILLER_34_3124 ();
 sg13g2_decap_8 FILLER_34_3131 ();
 sg13g2_decap_8 FILLER_34_3138 ();
 sg13g2_decap_8 FILLER_34_3145 ();
 sg13g2_decap_8 FILLER_34_3152 ();
 sg13g2_decap_4 FILLER_34_3159 ();
 sg13g2_fill_2 FILLER_34_3163 ();
 sg13g2_decap_8 FILLER_34_3170 ();
 sg13g2_decap_8 FILLER_34_3177 ();
 sg13g2_decap_8 FILLER_34_3184 ();
 sg13g2_decap_8 FILLER_34_3191 ();
 sg13g2_decap_8 FILLER_34_3198 ();
 sg13g2_decap_8 FILLER_34_3205 ();
 sg13g2_decap_8 FILLER_34_3212 ();
 sg13g2_decap_4 FILLER_34_3219 ();
 sg13g2_decap_8 FILLER_34_3229 ();
 sg13g2_decap_8 FILLER_34_3236 ();
 sg13g2_decap_8 FILLER_34_3243 ();
 sg13g2_fill_2 FILLER_34_3250 ();
 sg13g2_decap_8 FILLER_34_3288 ();
 sg13g2_decap_8 FILLER_34_3295 ();
 sg13g2_decap_8 FILLER_34_3302 ();
 sg13g2_decap_8 FILLER_34_3309 ();
 sg13g2_decap_8 FILLER_34_3316 ();
 sg13g2_decap_8 FILLER_34_3323 ();
 sg13g2_decap_8 FILLER_34_3330 ();
 sg13g2_decap_8 FILLER_34_3337 ();
 sg13g2_decap_8 FILLER_34_3344 ();
 sg13g2_decap_8 FILLER_34_3351 ();
 sg13g2_fill_1 FILLER_34_3358 ();
 sg13g2_decap_8 FILLER_34_3367 ();
 sg13g2_decap_8 FILLER_34_3374 ();
 sg13g2_decap_8 FILLER_34_3381 ();
 sg13g2_decap_8 FILLER_34_3388 ();
 sg13g2_fill_2 FILLER_34_3395 ();
 sg13g2_decap_8 FILLER_34_3402 ();
 sg13g2_decap_8 FILLER_34_3409 ();
 sg13g2_decap_8 FILLER_34_3416 ();
 sg13g2_decap_8 FILLER_34_3423 ();
 sg13g2_decap_8 FILLER_34_3430 ();
 sg13g2_decap_4 FILLER_34_3437 ();
 sg13g2_fill_1 FILLER_34_3446 ();
 sg13g2_fill_1 FILLER_34_3452 ();
 sg13g2_decap_8 FILLER_34_3458 ();
 sg13g2_decap_8 FILLER_34_3465 ();
 sg13g2_decap_8 FILLER_34_3472 ();
 sg13g2_fill_1 FILLER_34_3479 ();
 sg13g2_fill_1 FILLER_34_3485 ();
 sg13g2_decap_4 FILLER_34_3491 ();
 sg13g2_decap_8 FILLER_34_3500 ();
 sg13g2_decap_8 FILLER_34_3507 ();
 sg13g2_decap_8 FILLER_34_3514 ();
 sg13g2_decap_8 FILLER_34_3521 ();
 sg13g2_fill_2 FILLER_34_3540 ();
 sg13g2_fill_1 FILLER_34_3542 ();
 sg13g2_decap_8 FILLER_34_3553 ();
 sg13g2_decap_8 FILLER_34_3560 ();
 sg13g2_decap_8 FILLER_34_3567 ();
 sg13g2_decap_4 FILLER_34_3574 ();
 sg13g2_fill_2 FILLER_34_3578 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_fill_1 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_50 ();
 sg13g2_decap_8 FILLER_35_57 ();
 sg13g2_decap_4 FILLER_35_64 ();
 sg13g2_fill_2 FILLER_35_68 ();
 sg13g2_fill_2 FILLER_35_83 ();
 sg13g2_fill_1 FILLER_35_85 ();
 sg13g2_decap_4 FILLER_35_99 ();
 sg13g2_decap_8 FILLER_35_113 ();
 sg13g2_decap_8 FILLER_35_120 ();
 sg13g2_decap_4 FILLER_35_127 ();
 sg13g2_fill_2 FILLER_35_131 ();
 sg13g2_decap_8 FILLER_35_138 ();
 sg13g2_decap_8 FILLER_35_145 ();
 sg13g2_decap_8 FILLER_35_152 ();
 sg13g2_decap_8 FILLER_35_164 ();
 sg13g2_decap_8 FILLER_35_171 ();
 sg13g2_decap_8 FILLER_35_178 ();
 sg13g2_decap_8 FILLER_35_185 ();
 sg13g2_decap_8 FILLER_35_192 ();
 sg13g2_decap_8 FILLER_35_199 ();
 sg13g2_decap_8 FILLER_35_206 ();
 sg13g2_fill_2 FILLER_35_213 ();
 sg13g2_fill_1 FILLER_35_215 ();
 sg13g2_decap_8 FILLER_35_221 ();
 sg13g2_fill_2 FILLER_35_228 ();
 sg13g2_decap_4 FILLER_35_234 ();
 sg13g2_decap_8 FILLER_35_247 ();
 sg13g2_decap_8 FILLER_35_254 ();
 sg13g2_fill_1 FILLER_35_261 ();
 sg13g2_decap_8 FILLER_35_267 ();
 sg13g2_decap_8 FILLER_35_274 ();
 sg13g2_decap_8 FILLER_35_281 ();
 sg13g2_decap_8 FILLER_35_288 ();
 sg13g2_fill_1 FILLER_35_295 ();
 sg13g2_decap_4 FILLER_35_301 ();
 sg13g2_decap_8 FILLER_35_313 ();
 sg13g2_decap_8 FILLER_35_320 ();
 sg13g2_decap_4 FILLER_35_327 ();
 sg13g2_fill_1 FILLER_35_331 ();
 sg13g2_decap_8 FILLER_35_366 ();
 sg13g2_fill_2 FILLER_35_373 ();
 sg13g2_decap_8 FILLER_35_381 ();
 sg13g2_decap_4 FILLER_35_388 ();
 sg13g2_decap_8 FILLER_35_401 ();
 sg13g2_decap_8 FILLER_35_408 ();
 sg13g2_fill_2 FILLER_35_415 ();
 sg13g2_decap_8 FILLER_35_428 ();
 sg13g2_decap_8 FILLER_35_435 ();
 sg13g2_fill_1 FILLER_35_442 ();
 sg13g2_decap_8 FILLER_35_453 ();
 sg13g2_decap_8 FILLER_35_460 ();
 sg13g2_decap_8 FILLER_35_467 ();
 sg13g2_decap_8 FILLER_35_474 ();
 sg13g2_fill_2 FILLER_35_481 ();
 sg13g2_fill_1 FILLER_35_483 ();
 sg13g2_decap_8 FILLER_35_487 ();
 sg13g2_decap_8 FILLER_35_494 ();
 sg13g2_decap_8 FILLER_35_501 ();
 sg13g2_decap_8 FILLER_35_508 ();
 sg13g2_decap_8 FILLER_35_515 ();
 sg13g2_decap_8 FILLER_35_522 ();
 sg13g2_decap_4 FILLER_35_529 ();
 sg13g2_fill_1 FILLER_35_533 ();
 sg13g2_fill_2 FILLER_35_560 ();
 sg13g2_decap_8 FILLER_35_583 ();
 sg13g2_decap_8 FILLER_35_590 ();
 sg13g2_decap_8 FILLER_35_597 ();
 sg13g2_decap_4 FILLER_35_604 ();
 sg13g2_fill_1 FILLER_35_608 ();
 sg13g2_fill_2 FILLER_35_630 ();
 sg13g2_fill_1 FILLER_35_632 ();
 sg13g2_decap_8 FILLER_35_641 ();
 sg13g2_decap_8 FILLER_35_648 ();
 sg13g2_fill_2 FILLER_35_655 ();
 sg13g2_fill_2 FILLER_35_695 ();
 sg13g2_fill_1 FILLER_35_723 ();
 sg13g2_decap_4 FILLER_35_731 ();
 sg13g2_fill_2 FILLER_35_735 ();
 sg13g2_fill_1 FILLER_35_749 ();
 sg13g2_decap_4 FILLER_35_755 ();
 sg13g2_fill_1 FILLER_35_759 ();
 sg13g2_decap_8 FILLER_35_780 ();
 sg13g2_fill_2 FILLER_35_787 ();
 sg13g2_decap_8 FILLER_35_796 ();
 sg13g2_decap_8 FILLER_35_803 ();
 sg13g2_decap_8 FILLER_35_810 ();
 sg13g2_fill_1 FILLER_35_817 ();
 sg13g2_decap_8 FILLER_35_848 ();
 sg13g2_decap_8 FILLER_35_855 ();
 sg13g2_decap_8 FILLER_35_862 ();
 sg13g2_decap_8 FILLER_35_869 ();
 sg13g2_decap_8 FILLER_35_876 ();
 sg13g2_decap_8 FILLER_35_883 ();
 sg13g2_decap_8 FILLER_35_890 ();
 sg13g2_decap_8 FILLER_35_897 ();
 sg13g2_decap_8 FILLER_35_904 ();
 sg13g2_decap_8 FILLER_35_911 ();
 sg13g2_decap_8 FILLER_35_918 ();
 sg13g2_decap_8 FILLER_35_925 ();
 sg13g2_fill_2 FILLER_35_932 ();
 sg13g2_fill_1 FILLER_35_934 ();
 sg13g2_fill_2 FILLER_35_940 ();
 sg13g2_decap_8 FILLER_35_950 ();
 sg13g2_decap_8 FILLER_35_957 ();
 sg13g2_fill_2 FILLER_35_964 ();
 sg13g2_fill_1 FILLER_35_966 ();
 sg13g2_decap_8 FILLER_35_995 ();
 sg13g2_decap_8 FILLER_35_1002 ();
 sg13g2_decap_8 FILLER_35_1009 ();
 sg13g2_decap_8 FILLER_35_1016 ();
 sg13g2_decap_4 FILLER_35_1023 ();
 sg13g2_decap_4 FILLER_35_1051 ();
 sg13g2_fill_1 FILLER_35_1055 ();
 sg13g2_decap_8 FILLER_35_1060 ();
 sg13g2_decap_8 FILLER_35_1067 ();
 sg13g2_decap_8 FILLER_35_1074 ();
 sg13g2_decap_8 FILLER_35_1081 ();
 sg13g2_decap_8 FILLER_35_1088 ();
 sg13g2_decap_8 FILLER_35_1095 ();
 sg13g2_decap_8 FILLER_35_1102 ();
 sg13g2_decap_8 FILLER_35_1109 ();
 sg13g2_decap_8 FILLER_35_1121 ();
 sg13g2_decap_8 FILLER_35_1128 ();
 sg13g2_decap_8 FILLER_35_1135 ();
 sg13g2_decap_8 FILLER_35_1142 ();
 sg13g2_decap_4 FILLER_35_1149 ();
 sg13g2_decap_8 FILLER_35_1173 ();
 sg13g2_decap_8 FILLER_35_1180 ();
 sg13g2_decap_8 FILLER_35_1187 ();
 sg13g2_decap_8 FILLER_35_1194 ();
 sg13g2_decap_4 FILLER_35_1201 ();
 sg13g2_fill_2 FILLER_35_1258 ();
 sg13g2_decap_8 FILLER_35_1281 ();
 sg13g2_decap_8 FILLER_35_1288 ();
 sg13g2_decap_8 FILLER_35_1295 ();
 sg13g2_decap_8 FILLER_35_1302 ();
 sg13g2_fill_2 FILLER_35_1309 ();
 sg13g2_fill_2 FILLER_35_1325 ();
 sg13g2_decap_8 FILLER_35_1340 ();
 sg13g2_decap_8 FILLER_35_1347 ();
 sg13g2_decap_8 FILLER_35_1354 ();
 sg13g2_decap_8 FILLER_35_1361 ();
 sg13g2_decap_8 FILLER_35_1368 ();
 sg13g2_decap_8 FILLER_35_1375 ();
 sg13g2_decap_8 FILLER_35_1382 ();
 sg13g2_decap_8 FILLER_35_1389 ();
 sg13g2_decap_8 FILLER_35_1396 ();
 sg13g2_decap_8 FILLER_35_1403 ();
 sg13g2_fill_2 FILLER_35_1410 ();
 sg13g2_decap_8 FILLER_35_1422 ();
 sg13g2_decap_8 FILLER_35_1429 ();
 sg13g2_fill_2 FILLER_35_1436 ();
 sg13g2_decap_8 FILLER_35_1450 ();
 sg13g2_decap_8 FILLER_35_1457 ();
 sg13g2_decap_8 FILLER_35_1464 ();
 sg13g2_decap_8 FILLER_35_1476 ();
 sg13g2_decap_4 FILLER_35_1483 ();
 sg13g2_fill_1 FILLER_35_1487 ();
 sg13g2_decap_8 FILLER_35_1491 ();
 sg13g2_decap_8 FILLER_35_1498 ();
 sg13g2_decap_8 FILLER_35_1505 ();
 sg13g2_decap_8 FILLER_35_1522 ();
 sg13g2_decap_8 FILLER_35_1529 ();
 sg13g2_decap_8 FILLER_35_1536 ();
 sg13g2_decap_8 FILLER_35_1543 ();
 sg13g2_decap_8 FILLER_35_1550 ();
 sg13g2_decap_8 FILLER_35_1557 ();
 sg13g2_decap_8 FILLER_35_1564 ();
 sg13g2_decap_8 FILLER_35_1571 ();
 sg13g2_decap_8 FILLER_35_1578 ();
 sg13g2_decap_4 FILLER_35_1585 ();
 sg13g2_fill_1 FILLER_35_1589 ();
 sg13g2_decap_8 FILLER_35_1596 ();
 sg13g2_fill_1 FILLER_35_1603 ();
 sg13g2_decap_8 FILLER_35_1610 ();
 sg13g2_decap_8 FILLER_35_1617 ();
 sg13g2_decap_8 FILLER_35_1624 ();
 sg13g2_decap_4 FILLER_35_1631 ();
 sg13g2_fill_2 FILLER_35_1635 ();
 sg13g2_decap_8 FILLER_35_1662 ();
 sg13g2_decap_8 FILLER_35_1669 ();
 sg13g2_decap_8 FILLER_35_1676 ();
 sg13g2_decap_8 FILLER_35_1683 ();
 sg13g2_decap_8 FILLER_35_1690 ();
 sg13g2_decap_8 FILLER_35_1697 ();
 sg13g2_decap_8 FILLER_35_1704 ();
 sg13g2_decap_4 FILLER_35_1711 ();
 sg13g2_decap_8 FILLER_35_1721 ();
 sg13g2_decap_8 FILLER_35_1728 ();
 sg13g2_decap_8 FILLER_35_1735 ();
 sg13g2_decap_8 FILLER_35_1742 ();
 sg13g2_decap_4 FILLER_35_1781 ();
 sg13g2_fill_2 FILLER_35_1785 ();
 sg13g2_decap_8 FILLER_35_1793 ();
 sg13g2_decap_8 FILLER_35_1800 ();
 sg13g2_decap_8 FILLER_35_1807 ();
 sg13g2_fill_2 FILLER_35_1814 ();
 sg13g2_fill_1 FILLER_35_1816 ();
 sg13g2_decap_4 FILLER_35_1827 ();
 sg13g2_fill_1 FILLER_35_1831 ();
 sg13g2_decap_8 FILLER_35_1858 ();
 sg13g2_decap_8 FILLER_35_1865 ();
 sg13g2_decap_8 FILLER_35_1872 ();
 sg13g2_decap_8 FILLER_35_1879 ();
 sg13g2_decap_4 FILLER_35_1886 ();
 sg13g2_fill_2 FILLER_35_1890 ();
 sg13g2_decap_8 FILLER_35_1903 ();
 sg13g2_decap_8 FILLER_35_1910 ();
 sg13g2_decap_8 FILLER_35_1938 ();
 sg13g2_decap_8 FILLER_35_1951 ();
 sg13g2_fill_2 FILLER_35_1958 ();
 sg13g2_fill_1 FILLER_35_1960 ();
 sg13g2_decap_4 FILLER_35_1967 ();
 sg13g2_fill_2 FILLER_35_1971 ();
 sg13g2_decap_4 FILLER_35_1985 ();
 sg13g2_decap_8 FILLER_35_1995 ();
 sg13g2_decap_8 FILLER_35_2002 ();
 sg13g2_fill_2 FILLER_35_2009 ();
 sg13g2_fill_2 FILLER_35_2025 ();
 sg13g2_fill_1 FILLER_35_2027 ();
 sg13g2_decap_8 FILLER_35_2058 ();
 sg13g2_decap_8 FILLER_35_2065 ();
 sg13g2_decap_8 FILLER_35_2072 ();
 sg13g2_decap_8 FILLER_35_2079 ();
 sg13g2_decap_8 FILLER_35_2086 ();
 sg13g2_fill_1 FILLER_35_2093 ();
 sg13g2_fill_1 FILLER_35_2097 ();
 sg13g2_decap_8 FILLER_35_2104 ();
 sg13g2_decap_4 FILLER_35_2111 ();
 sg13g2_decap_8 FILLER_35_2127 ();
 sg13g2_decap_4 FILLER_35_2134 ();
 sg13g2_fill_1 FILLER_35_2138 ();
 sg13g2_fill_2 FILLER_35_2151 ();
 sg13g2_decap_4 FILLER_35_2165 ();
 sg13g2_fill_2 FILLER_35_2169 ();
 sg13g2_fill_2 FILLER_35_2177 ();
 sg13g2_fill_1 FILLER_35_2179 ();
 sg13g2_decap_8 FILLER_35_2186 ();
 sg13g2_decap_8 FILLER_35_2193 ();
 sg13g2_decap_8 FILLER_35_2200 ();
 sg13g2_decap_8 FILLER_35_2207 ();
 sg13g2_fill_1 FILLER_35_2214 ();
 sg13g2_decap_8 FILLER_35_2221 ();
 sg13g2_decap_4 FILLER_35_2228 ();
 sg13g2_fill_1 FILLER_35_2232 ();
 sg13g2_decap_8 FILLER_35_2251 ();
 sg13g2_fill_1 FILLER_35_2258 ();
 sg13g2_decap_8 FILLER_35_2265 ();
 sg13g2_decap_8 FILLER_35_2272 ();
 sg13g2_fill_1 FILLER_35_2285 ();
 sg13g2_fill_1 FILLER_35_2292 ();
 sg13g2_decap_8 FILLER_35_2299 ();
 sg13g2_decap_8 FILLER_35_2306 ();
 sg13g2_decap_8 FILLER_35_2313 ();
 sg13g2_decap_4 FILLER_35_2320 ();
 sg13g2_fill_1 FILLER_35_2324 ();
 sg13g2_decap_8 FILLER_35_2331 ();
 sg13g2_decap_8 FILLER_35_2338 ();
 sg13g2_fill_2 FILLER_35_2345 ();
 sg13g2_decap_8 FILLER_35_2359 ();
 sg13g2_decap_4 FILLER_35_2366 ();
 sg13g2_decap_8 FILLER_35_2376 ();
 sg13g2_decap_4 FILLER_35_2383 ();
 sg13g2_fill_1 FILLER_35_2387 ();
 sg13g2_fill_2 FILLER_35_2394 ();
 sg13g2_fill_1 FILLER_35_2396 ();
 sg13g2_decap_8 FILLER_35_2415 ();
 sg13g2_decap_8 FILLER_35_2422 ();
 sg13g2_decap_4 FILLER_35_2429 ();
 sg13g2_fill_1 FILLER_35_2433 ();
 sg13g2_decap_4 FILLER_35_2446 ();
 sg13g2_fill_2 FILLER_35_2450 ();
 sg13g2_fill_2 FILLER_35_2463 ();
 sg13g2_fill_1 FILLER_35_2465 ();
 sg13g2_decap_8 FILLER_35_2473 ();
 sg13g2_decap_8 FILLER_35_2480 ();
 sg13g2_decap_8 FILLER_35_2487 ();
 sg13g2_decap_8 FILLER_35_2494 ();
 sg13g2_decap_8 FILLER_35_2501 ();
 sg13g2_decap_8 FILLER_35_2508 ();
 sg13g2_decap_8 FILLER_35_2515 ();
 sg13g2_decap_8 FILLER_35_2527 ();
 sg13g2_decap_8 FILLER_35_2534 ();
 sg13g2_decap_8 FILLER_35_2541 ();
 sg13g2_decap_4 FILLER_35_2556 ();
 sg13g2_fill_2 FILLER_35_2566 ();
 sg13g2_fill_1 FILLER_35_2568 ();
 sg13g2_decap_8 FILLER_35_2574 ();
 sg13g2_decap_8 FILLER_35_2581 ();
 sg13g2_decap_4 FILLER_35_2588 ();
 sg13g2_fill_1 FILLER_35_2592 ();
 sg13g2_decap_8 FILLER_35_2599 ();
 sg13g2_fill_1 FILLER_35_2606 ();
 sg13g2_fill_1 FILLER_35_2610 ();
 sg13g2_fill_1 FILLER_35_2617 ();
 sg13g2_fill_2 FILLER_35_2624 ();
 sg13g2_fill_2 FILLER_35_2669 ();
 sg13g2_decap_8 FILLER_35_2676 ();
 sg13g2_decap_8 FILLER_35_2683 ();
 sg13g2_decap_8 FILLER_35_2690 ();
 sg13g2_decap_8 FILLER_35_2697 ();
 sg13g2_decap_4 FILLER_35_2704 ();
 sg13g2_fill_2 FILLER_35_2708 ();
 sg13g2_decap_8 FILLER_35_2716 ();
 sg13g2_decap_8 FILLER_35_2723 ();
 sg13g2_decap_8 FILLER_35_2730 ();
 sg13g2_decap_8 FILLER_35_2737 ();
 sg13g2_decap_8 FILLER_35_2744 ();
 sg13g2_decap_8 FILLER_35_2751 ();
 sg13g2_fill_2 FILLER_35_2779 ();
 sg13g2_fill_1 FILLER_35_2801 ();
 sg13g2_decap_8 FILLER_35_2812 ();
 sg13g2_decap_8 FILLER_35_2829 ();
 sg13g2_fill_2 FILLER_35_2836 ();
 sg13g2_fill_1 FILLER_35_2838 ();
 sg13g2_decap_8 FILLER_35_2844 ();
 sg13g2_decap_4 FILLER_35_2851 ();
 sg13g2_fill_2 FILLER_35_2855 ();
 sg13g2_decap_8 FILLER_35_2934 ();
 sg13g2_decap_8 FILLER_35_2941 ();
 sg13g2_decap_8 FILLER_35_2948 ();
 sg13g2_decap_4 FILLER_35_2955 ();
 sg13g2_fill_1 FILLER_35_2959 ();
 sg13g2_decap_8 FILLER_35_2965 ();
 sg13g2_decap_8 FILLER_35_2972 ();
 sg13g2_decap_8 FILLER_35_2979 ();
 sg13g2_decap_8 FILLER_35_2986 ();
 sg13g2_decap_4 FILLER_35_2993 ();
 sg13g2_fill_1 FILLER_35_2997 ();
 sg13g2_decap_8 FILLER_35_3008 ();
 sg13g2_decap_8 FILLER_35_3015 ();
 sg13g2_decap_8 FILLER_35_3022 ();
 sg13g2_fill_2 FILLER_35_3029 ();
 sg13g2_decap_8 FILLER_35_3057 ();
 sg13g2_decap_8 FILLER_35_3064 ();
 sg13g2_decap_8 FILLER_35_3071 ();
 sg13g2_decap_4 FILLER_35_3104 ();
 sg13g2_fill_1 FILLER_35_3108 ();
 sg13g2_decap_8 FILLER_35_3145 ();
 sg13g2_decap_8 FILLER_35_3152 ();
 sg13g2_decap_8 FILLER_35_3159 ();
 sg13g2_fill_2 FILLER_35_3166 ();
 sg13g2_decap_8 FILLER_35_3194 ();
 sg13g2_decap_8 FILLER_35_3201 ();
 sg13g2_decap_8 FILLER_35_3208 ();
 sg13g2_decap_8 FILLER_35_3215 ();
 sg13g2_fill_2 FILLER_35_3222 ();
 sg13g2_decap_4 FILLER_35_3234 ();
 sg13g2_fill_2 FILLER_35_3238 ();
 sg13g2_decap_8 FILLER_35_3248 ();
 sg13g2_decap_8 FILLER_35_3255 ();
 sg13g2_decap_8 FILLER_35_3262 ();
 sg13g2_decap_8 FILLER_35_3269 ();
 sg13g2_decap_8 FILLER_35_3276 ();
 sg13g2_decap_8 FILLER_35_3283 ();
 sg13g2_decap_4 FILLER_35_3290 ();
 sg13g2_fill_1 FILLER_35_3294 ();
 sg13g2_decap_8 FILLER_35_3331 ();
 sg13g2_decap_8 FILLER_35_3338 ();
 sg13g2_decap_8 FILLER_35_3345 ();
 sg13g2_decap_8 FILLER_35_3352 ();
 sg13g2_decap_8 FILLER_35_3359 ();
 sg13g2_decap_8 FILLER_35_3366 ();
 sg13g2_decap_8 FILLER_35_3373 ();
 sg13g2_decap_4 FILLER_35_3380 ();
 sg13g2_fill_2 FILLER_35_3384 ();
 sg13g2_fill_2 FILLER_35_3400 ();
 sg13g2_decap_8 FILLER_35_3428 ();
 sg13g2_decap_8 FILLER_35_3435 ();
 sg13g2_decap_8 FILLER_35_3442 ();
 sg13g2_fill_2 FILLER_35_3449 ();
 sg13g2_decap_4 FILLER_35_3456 ();
 sg13g2_fill_1 FILLER_35_3460 ();
 sg13g2_decap_8 FILLER_35_3466 ();
 sg13g2_decap_8 FILLER_35_3477 ();
 sg13g2_decap_8 FILLER_35_3484 ();
 sg13g2_decap_8 FILLER_35_3491 ();
 sg13g2_decap_8 FILLER_35_3498 ();
 sg13g2_decap_8 FILLER_35_3505 ();
 sg13g2_fill_2 FILLER_35_3512 ();
 sg13g2_fill_1 FILLER_35_3514 ();
 sg13g2_decap_8 FILLER_35_3518 ();
 sg13g2_decap_4 FILLER_35_3525 ();
 sg13g2_fill_1 FILLER_35_3529 ();
 sg13g2_decap_8 FILLER_35_3535 ();
 sg13g2_decap_8 FILLER_35_3542 ();
 sg13g2_fill_1 FILLER_35_3549 ();
 sg13g2_decap_8 FILLER_35_3555 ();
 sg13g2_decap_8 FILLER_35_3562 ();
 sg13g2_decap_8 FILLER_35_3569 ();
 sg13g2_decap_4 FILLER_35_3576 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_fill_1 FILLER_36_78 ();
 sg13g2_fill_1 FILLER_36_90 ();
 sg13g2_decap_4 FILLER_36_101 ();
 sg13g2_fill_1 FILLER_36_105 ();
 sg13g2_decap_8 FILLER_36_114 ();
 sg13g2_decap_4 FILLER_36_121 ();
 sg13g2_fill_2 FILLER_36_125 ();
 sg13g2_fill_1 FILLER_36_143 ();
 sg13g2_decap_8 FILLER_36_171 ();
 sg13g2_decap_8 FILLER_36_178 ();
 sg13g2_decap_8 FILLER_36_185 ();
 sg13g2_decap_8 FILLER_36_192 ();
 sg13g2_decap_8 FILLER_36_199 ();
 sg13g2_decap_8 FILLER_36_206 ();
 sg13g2_decap_4 FILLER_36_213 ();
 sg13g2_fill_2 FILLER_36_217 ();
 sg13g2_fill_2 FILLER_36_266 ();
 sg13g2_fill_1 FILLER_36_268 ();
 sg13g2_decap_8 FILLER_36_282 ();
 sg13g2_decap_8 FILLER_36_289 ();
 sg13g2_decap_8 FILLER_36_296 ();
 sg13g2_decap_8 FILLER_36_303 ();
 sg13g2_decap_8 FILLER_36_310 ();
 sg13g2_decap_8 FILLER_36_317 ();
 sg13g2_decap_8 FILLER_36_324 ();
 sg13g2_decap_8 FILLER_36_331 ();
 sg13g2_decap_8 FILLER_36_338 ();
 sg13g2_decap_8 FILLER_36_345 ();
 sg13g2_decap_8 FILLER_36_352 ();
 sg13g2_decap_8 FILLER_36_359 ();
 sg13g2_fill_2 FILLER_36_366 ();
 sg13g2_fill_1 FILLER_36_368 ();
 sg13g2_decap_8 FILLER_36_393 ();
 sg13g2_fill_2 FILLER_36_400 ();
 sg13g2_fill_1 FILLER_36_402 ();
 sg13g2_decap_8 FILLER_36_443 ();
 sg13g2_decap_8 FILLER_36_450 ();
 sg13g2_decap_8 FILLER_36_457 ();
 sg13g2_decap_8 FILLER_36_464 ();
 sg13g2_decap_8 FILLER_36_471 ();
 sg13g2_decap_8 FILLER_36_521 ();
 sg13g2_decap_8 FILLER_36_528 ();
 sg13g2_decap_8 FILLER_36_535 ();
 sg13g2_decap_4 FILLER_36_542 ();
 sg13g2_fill_2 FILLER_36_546 ();
 sg13g2_decap_4 FILLER_36_554 ();
 sg13g2_fill_2 FILLER_36_558 ();
 sg13g2_decap_8 FILLER_36_584 ();
 sg13g2_decap_8 FILLER_36_596 ();
 sg13g2_decap_8 FILLER_36_603 ();
 sg13g2_decap_8 FILLER_36_610 ();
 sg13g2_decap_8 FILLER_36_620 ();
 sg13g2_decap_8 FILLER_36_627 ();
 sg13g2_fill_1 FILLER_36_634 ();
 sg13g2_decap_8 FILLER_36_645 ();
 sg13g2_decap_8 FILLER_36_652 ();
 sg13g2_decap_4 FILLER_36_659 ();
 sg13g2_fill_1 FILLER_36_663 ();
 sg13g2_fill_1 FILLER_36_696 ();
 sg13g2_decap_8 FILLER_36_702 ();
 sg13g2_decap_8 FILLER_36_709 ();
 sg13g2_decap_4 FILLER_36_724 ();
 sg13g2_decap_8 FILLER_36_736 ();
 sg13g2_fill_1 FILLER_36_743 ();
 sg13g2_fill_2 FILLER_36_773 ();
 sg13g2_fill_1 FILLER_36_775 ();
 sg13g2_decap_8 FILLER_36_804 ();
 sg13g2_decap_4 FILLER_36_811 ();
 sg13g2_fill_2 FILLER_36_831 ();
 sg13g2_fill_1 FILLER_36_833 ();
 sg13g2_decap_8 FILLER_36_860 ();
 sg13g2_decap_8 FILLER_36_867 ();
 sg13g2_decap_8 FILLER_36_874 ();
 sg13g2_decap_8 FILLER_36_881 ();
 sg13g2_decap_8 FILLER_36_914 ();
 sg13g2_decap_8 FILLER_36_921 ();
 sg13g2_decap_8 FILLER_36_928 ();
 sg13g2_decap_8 FILLER_36_971 ();
 sg13g2_decap_8 FILLER_36_978 ();
 sg13g2_fill_1 FILLER_36_985 ();
 sg13g2_decap_4 FILLER_36_1012 ();
 sg13g2_fill_1 FILLER_36_1016 ();
 sg13g2_decap_8 FILLER_36_1042 ();
 sg13g2_decap_8 FILLER_36_1049 ();
 sg13g2_decap_8 FILLER_36_1056 ();
 sg13g2_decap_8 FILLER_36_1063 ();
 sg13g2_decap_8 FILLER_36_1070 ();
 sg13g2_fill_2 FILLER_36_1077 ();
 sg13g2_fill_1 FILLER_36_1079 ();
 sg13g2_decap_8 FILLER_36_1128 ();
 sg13g2_decap_8 FILLER_36_1135 ();
 sg13g2_decap_8 FILLER_36_1142 ();
 sg13g2_decap_8 FILLER_36_1149 ();
 sg13g2_decap_8 FILLER_36_1156 ();
 sg13g2_decap_8 FILLER_36_1189 ();
 sg13g2_decap_8 FILLER_36_1196 ();
 sg13g2_fill_1 FILLER_36_1203 ();
 sg13g2_decap_8 FILLER_36_1225 ();
 sg13g2_decap_8 FILLER_36_1232 ();
 sg13g2_fill_2 FILLER_36_1274 ();
 sg13g2_fill_2 FILLER_36_1285 ();
 sg13g2_decap_4 FILLER_36_1295 ();
 sg13g2_fill_2 FILLER_36_1299 ();
 sg13g2_decap_4 FILLER_36_1310 ();
 sg13g2_fill_1 FILLER_36_1314 ();
 sg13g2_fill_2 FILLER_36_1323 ();
 sg13g2_fill_1 FILLER_36_1325 ();
 sg13g2_decap_8 FILLER_36_1355 ();
 sg13g2_decap_8 FILLER_36_1362 ();
 sg13g2_decap_8 FILLER_36_1369 ();
 sg13g2_fill_2 FILLER_36_1376 ();
 sg13g2_fill_1 FILLER_36_1378 ();
 sg13g2_decap_8 FILLER_36_1390 ();
 sg13g2_decap_8 FILLER_36_1397 ();
 sg13g2_fill_2 FILLER_36_1404 ();
 sg13g2_fill_1 FILLER_36_1406 ();
 sg13g2_decap_8 FILLER_36_1433 ();
 sg13g2_decap_8 FILLER_36_1446 ();
 sg13g2_decap_8 FILLER_36_1453 ();
 sg13g2_decap_8 FILLER_36_1460 ();
 sg13g2_decap_8 FILLER_36_1467 ();
 sg13g2_fill_1 FILLER_36_1474 ();
 sg13g2_decap_8 FILLER_36_1478 ();
 sg13g2_decap_4 FILLER_36_1485 ();
 sg13g2_fill_1 FILLER_36_1489 ();
 sg13g2_decap_8 FILLER_36_1502 ();
 sg13g2_decap_8 FILLER_36_1509 ();
 sg13g2_fill_1 FILLER_36_1516 ();
 sg13g2_decap_4 FILLER_36_1520 ();
 sg13g2_decap_8 FILLER_36_1550 ();
 sg13g2_decap_8 FILLER_36_1557 ();
 sg13g2_decap_8 FILLER_36_1564 ();
 sg13g2_decap_8 FILLER_36_1571 ();
 sg13g2_decap_8 FILLER_36_1578 ();
 sg13g2_decap_8 FILLER_36_1585 ();
 sg13g2_decap_8 FILLER_36_1592 ();
 sg13g2_decap_8 FILLER_36_1599 ();
 sg13g2_decap_8 FILLER_36_1606 ();
 sg13g2_decap_8 FILLER_36_1613 ();
 sg13g2_decap_8 FILLER_36_1620 ();
 sg13g2_fill_2 FILLER_36_1627 ();
 sg13g2_fill_1 FILLER_36_1629 ();
 sg13g2_decap_8 FILLER_36_1656 ();
 sg13g2_decap_8 FILLER_36_1663 ();
 sg13g2_decap_8 FILLER_36_1670 ();
 sg13g2_decap_8 FILLER_36_1677 ();
 sg13g2_decap_8 FILLER_36_1684 ();
 sg13g2_decap_8 FILLER_36_1691 ();
 sg13g2_decap_8 FILLER_36_1698 ();
 sg13g2_decap_8 FILLER_36_1705 ();
 sg13g2_decap_8 FILLER_36_1712 ();
 sg13g2_decap_8 FILLER_36_1739 ();
 sg13g2_fill_2 FILLER_36_1746 ();
 sg13g2_decap_8 FILLER_36_1754 ();
 sg13g2_decap_8 FILLER_36_1761 ();
 sg13g2_decap_8 FILLER_36_1768 ();
 sg13g2_decap_8 FILLER_36_1775 ();
 sg13g2_decap_8 FILLER_36_1782 ();
 sg13g2_decap_8 FILLER_36_1795 ();
 sg13g2_decap_8 FILLER_36_1802 ();
 sg13g2_decap_8 FILLER_36_1809 ();
 sg13g2_decap_8 FILLER_36_1816 ();
 sg13g2_decap_8 FILLER_36_1823 ();
 sg13g2_decap_8 FILLER_36_1830 ();
 sg13g2_decap_8 FILLER_36_1837 ();
 sg13g2_decap_4 FILLER_36_1844 ();
 sg13g2_decap_8 FILLER_36_1859 ();
 sg13g2_decap_4 FILLER_36_1866 ();
 sg13g2_fill_2 FILLER_36_1870 ();
 sg13g2_fill_1 FILLER_36_1880 ();
 sg13g2_decap_8 FILLER_36_1890 ();
 sg13g2_decap_8 FILLER_36_1897 ();
 sg13g2_decap_8 FILLER_36_1904 ();
 sg13g2_decap_4 FILLER_36_1911 ();
 sg13g2_fill_1 FILLER_36_1915 ();
 sg13g2_decap_8 FILLER_36_1938 ();
 sg13g2_decap_8 FILLER_36_1945 ();
 sg13g2_decap_8 FILLER_36_1952 ();
 sg13g2_decap_8 FILLER_36_1959 ();
 sg13g2_decap_4 FILLER_36_1966 ();
 sg13g2_fill_1 FILLER_36_1970 ();
 sg13g2_decap_8 FILLER_36_2029 ();
 sg13g2_decap_8 FILLER_36_2036 ();
 sg13g2_decap_4 FILLER_36_2043 ();
 sg13g2_fill_1 FILLER_36_2047 ();
 sg13g2_decap_8 FILLER_36_2074 ();
 sg13g2_decap_4 FILLER_36_2081 ();
 sg13g2_fill_1 FILLER_36_2097 ();
 sg13g2_decap_8 FILLER_36_2104 ();
 sg13g2_fill_2 FILLER_36_2111 ();
 sg13g2_fill_1 FILLER_36_2113 ();
 sg13g2_decap_4 FILLER_36_2120 ();
 sg13g2_fill_1 FILLER_36_2124 ();
 sg13g2_decap_8 FILLER_36_2158 ();
 sg13g2_decap_8 FILLER_36_2165 ();
 sg13g2_decap_8 FILLER_36_2172 ();
 sg13g2_decap_4 FILLER_36_2179 ();
 sg13g2_fill_2 FILLER_36_2183 ();
 sg13g2_decap_8 FILLER_36_2191 ();
 sg13g2_decap_8 FILLER_36_2198 ();
 sg13g2_decap_8 FILLER_36_2205 ();
 sg13g2_fill_2 FILLER_36_2212 ();
 sg13g2_fill_1 FILLER_36_2214 ();
 sg13g2_fill_1 FILLER_36_2218 ();
 sg13g2_fill_2 FILLER_36_2239 ();
 sg13g2_fill_1 FILLER_36_2241 ();
 sg13g2_decap_8 FILLER_36_2248 ();
 sg13g2_fill_2 FILLER_36_2255 ();
 sg13g2_decap_8 FILLER_36_2263 ();
 sg13g2_decap_8 FILLER_36_2270 ();
 sg13g2_decap_8 FILLER_36_2277 ();
 sg13g2_decap_8 FILLER_36_2284 ();
 sg13g2_decap_8 FILLER_36_2291 ();
 sg13g2_fill_2 FILLER_36_2298 ();
 sg13g2_decap_8 FILLER_36_2306 ();
 sg13g2_decap_8 FILLER_36_2313 ();
 sg13g2_decap_8 FILLER_36_2320 ();
 sg13g2_decap_8 FILLER_36_2333 ();
 sg13g2_fill_1 FILLER_36_2340 ();
 sg13g2_decap_4 FILLER_36_2347 ();
 sg13g2_fill_1 FILLER_36_2351 ();
 sg13g2_decap_8 FILLER_36_2366 ();
 sg13g2_decap_4 FILLER_36_2373 ();
 sg13g2_decap_4 FILLER_36_2383 ();
 sg13g2_fill_2 FILLER_36_2387 ();
 sg13g2_fill_2 FILLER_36_2407 ();
 sg13g2_decap_8 FILLER_36_2417 ();
 sg13g2_decap_8 FILLER_36_2424 ();
 sg13g2_decap_8 FILLER_36_2431 ();
 sg13g2_decap_8 FILLER_36_2438 ();
 sg13g2_fill_1 FILLER_36_2449 ();
 sg13g2_decap_8 FILLER_36_2456 ();
 sg13g2_fill_2 FILLER_36_2467 ();
 sg13g2_decap_8 FILLER_36_2477 ();
 sg13g2_decap_4 FILLER_36_2484 ();
 sg13g2_fill_2 FILLER_36_2488 ();
 sg13g2_decap_8 FILLER_36_2498 ();
 sg13g2_decap_8 FILLER_36_2505 ();
 sg13g2_decap_8 FILLER_36_2512 ();
 sg13g2_fill_1 FILLER_36_2519 ();
 sg13g2_decap_8 FILLER_36_2533 ();
 sg13g2_decap_8 FILLER_36_2540 ();
 sg13g2_decap_8 FILLER_36_2547 ();
 sg13g2_fill_2 FILLER_36_2554 ();
 sg13g2_decap_4 FILLER_36_2562 ();
 sg13g2_decap_8 FILLER_36_2572 ();
 sg13g2_decap_8 FILLER_36_2579 ();
 sg13g2_decap_8 FILLER_36_2586 ();
 sg13g2_decap_8 FILLER_36_2593 ();
 sg13g2_decap_8 FILLER_36_2600 ();
 sg13g2_decap_4 FILLER_36_2607 ();
 sg13g2_fill_1 FILLER_36_2621 ();
 sg13g2_decap_8 FILLER_36_2633 ();
 sg13g2_decap_8 FILLER_36_2640 ();
 sg13g2_decap_8 FILLER_36_2647 ();
 sg13g2_decap_8 FILLER_36_2654 ();
 sg13g2_decap_8 FILLER_36_2661 ();
 sg13g2_decap_8 FILLER_36_2668 ();
 sg13g2_decap_8 FILLER_36_2675 ();
 sg13g2_decap_8 FILLER_36_2682 ();
 sg13g2_decap_8 FILLER_36_2689 ();
 sg13g2_decap_8 FILLER_36_2696 ();
 sg13g2_fill_1 FILLER_36_2703 ();
 sg13g2_decap_8 FILLER_36_2709 ();
 sg13g2_decap_8 FILLER_36_2716 ();
 sg13g2_decap_8 FILLER_36_2723 ();
 sg13g2_decap_8 FILLER_36_2745 ();
 sg13g2_decap_8 FILLER_36_2752 ();
 sg13g2_decap_8 FILLER_36_2759 ();
 sg13g2_decap_8 FILLER_36_2766 ();
 sg13g2_fill_2 FILLER_36_2773 ();
 sg13g2_fill_2 FILLER_36_2780 ();
 sg13g2_decap_8 FILLER_36_2786 ();
 sg13g2_decap_4 FILLER_36_2793 ();
 sg13g2_decap_8 FILLER_36_2849 ();
 sg13g2_decap_8 FILLER_36_2856 ();
 sg13g2_decap_4 FILLER_36_2863 ();
 sg13g2_decap_8 FILLER_36_2887 ();
 sg13g2_decap_8 FILLER_36_2894 ();
 sg13g2_decap_8 FILLER_36_2901 ();
 sg13g2_decap_4 FILLER_36_2908 ();
 sg13g2_fill_2 FILLER_36_2912 ();
 sg13g2_fill_2 FILLER_36_2929 ();
 sg13g2_decap_4 FILLER_36_2935 ();
 sg13g2_fill_1 FILLER_36_2939 ();
 sg13g2_decap_4 FILLER_36_2950 ();
 sg13g2_decap_8 FILLER_36_2964 ();
 sg13g2_decap_8 FILLER_36_2971 ();
 sg13g2_decap_8 FILLER_36_2978 ();
 sg13g2_fill_2 FILLER_36_2985 ();
 sg13g2_fill_1 FILLER_36_2987 ();
 sg13g2_decap_8 FILLER_36_2996 ();
 sg13g2_fill_1 FILLER_36_3003 ();
 sg13g2_decap_8 FILLER_36_3012 ();
 sg13g2_decap_8 FILLER_36_3019 ();
 sg13g2_decap_8 FILLER_36_3026 ();
 sg13g2_decap_4 FILLER_36_3033 ();
 sg13g2_fill_2 FILLER_36_3037 ();
 sg13g2_decap_8 FILLER_36_3049 ();
 sg13g2_decap_8 FILLER_36_3056 ();
 sg13g2_fill_1 FILLER_36_3063 ();
 sg13g2_decap_4 FILLER_36_3100 ();
 sg13g2_fill_1 FILLER_36_3104 ();
 sg13g2_decap_8 FILLER_36_3141 ();
 sg13g2_decap_8 FILLER_36_3148 ();
 sg13g2_decap_8 FILLER_36_3155 ();
 sg13g2_decap_4 FILLER_36_3162 ();
 sg13g2_decap_8 FILLER_36_3202 ();
 sg13g2_decap_8 FILLER_36_3209 ();
 sg13g2_fill_1 FILLER_36_3216 ();
 sg13g2_decap_8 FILLER_36_3243 ();
 sg13g2_decap_8 FILLER_36_3250 ();
 sg13g2_decap_8 FILLER_36_3267 ();
 sg13g2_decap_8 FILLER_36_3274 ();
 sg13g2_fill_2 FILLER_36_3281 ();
 sg13g2_fill_1 FILLER_36_3283 ();
 sg13g2_decap_8 FILLER_36_3294 ();
 sg13g2_fill_2 FILLER_36_3301 ();
 sg13g2_decap_8 FILLER_36_3311 ();
 sg13g2_decap_8 FILLER_36_3318 ();
 sg13g2_decap_8 FILLER_36_3325 ();
 sg13g2_decap_4 FILLER_36_3332 ();
 sg13g2_decap_8 FILLER_36_3356 ();
 sg13g2_decap_8 FILLER_36_3363 ();
 sg13g2_decap_8 FILLER_36_3370 ();
 sg13g2_decap_4 FILLER_36_3377 ();
 sg13g2_fill_1 FILLER_36_3381 ();
 sg13g2_decap_4 FILLER_36_3392 ();
 sg13g2_fill_1 FILLER_36_3396 ();
 sg13g2_decap_8 FILLER_36_3423 ();
 sg13g2_decap_8 FILLER_36_3430 ();
 sg13g2_decap_8 FILLER_36_3437 ();
 sg13g2_fill_2 FILLER_36_3444 ();
 sg13g2_decap_8 FILLER_36_3451 ();
 sg13g2_decap_8 FILLER_36_3458 ();
 sg13g2_decap_8 FILLER_36_3500 ();
 sg13g2_decap_8 FILLER_36_3507 ();
 sg13g2_decap_8 FILLER_36_3514 ();
 sg13g2_decap_4 FILLER_36_3521 ();
 sg13g2_fill_2 FILLER_36_3525 ();
 sg13g2_decap_8 FILLER_36_3545 ();
 sg13g2_decap_8 FILLER_36_3552 ();
 sg13g2_decap_8 FILLER_36_3559 ();
 sg13g2_decap_8 FILLER_36_3566 ();
 sg13g2_decap_8 FILLER_36_3573 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_4 FILLER_37_14 ();
 sg13g2_fill_1 FILLER_37_18 ();
 sg13g2_decap_8 FILLER_37_27 ();
 sg13g2_decap_8 FILLER_37_34 ();
 sg13g2_decap_8 FILLER_37_41 ();
 sg13g2_decap_8 FILLER_37_48 ();
 sg13g2_decap_8 FILLER_37_55 ();
 sg13g2_decap_4 FILLER_37_62 ();
 sg13g2_decap_8 FILLER_37_102 ();
 sg13g2_decap_8 FILLER_37_109 ();
 sg13g2_decap_8 FILLER_37_116 ();
 sg13g2_decap_8 FILLER_37_123 ();
 sg13g2_decap_8 FILLER_37_130 ();
 sg13g2_fill_2 FILLER_37_137 ();
 sg13g2_fill_2 FILLER_37_147 ();
 sg13g2_decap_8 FILLER_37_179 ();
 sg13g2_decap_8 FILLER_37_186 ();
 sg13g2_decap_8 FILLER_37_193 ();
 sg13g2_decap_8 FILLER_37_200 ();
 sg13g2_decap_4 FILLER_37_207 ();
 sg13g2_fill_2 FILLER_37_211 ();
 sg13g2_decap_8 FILLER_37_221 ();
 sg13g2_decap_8 FILLER_37_228 ();
 sg13g2_decap_8 FILLER_37_235 ();
 sg13g2_decap_8 FILLER_37_242 ();
 sg13g2_decap_8 FILLER_37_249 ();
 sg13g2_fill_2 FILLER_37_256 ();
 sg13g2_fill_1 FILLER_37_266 ();
 sg13g2_decap_8 FILLER_37_275 ();
 sg13g2_decap_8 FILLER_37_282 ();
 sg13g2_decap_8 FILLER_37_289 ();
 sg13g2_decap_8 FILLER_37_296 ();
 sg13g2_decap_8 FILLER_37_303 ();
 sg13g2_decap_8 FILLER_37_310 ();
 sg13g2_decap_8 FILLER_37_317 ();
 sg13g2_decap_8 FILLER_37_324 ();
 sg13g2_decap_8 FILLER_37_331 ();
 sg13g2_fill_1 FILLER_37_338 ();
 sg13g2_decap_8 FILLER_37_365 ();
 sg13g2_decap_8 FILLER_37_372 ();
 sg13g2_decap_8 FILLER_37_384 ();
 sg13g2_decap_8 FILLER_37_391 ();
 sg13g2_decap_8 FILLER_37_398 ();
 sg13g2_decap_8 FILLER_37_405 ();
 sg13g2_decap_8 FILLER_37_412 ();
 sg13g2_decap_8 FILLER_37_427 ();
 sg13g2_decap_8 FILLER_37_434 ();
 sg13g2_decap_8 FILLER_37_441 ();
 sg13g2_decap_8 FILLER_37_448 ();
 sg13g2_decap_8 FILLER_37_455 ();
 sg13g2_fill_1 FILLER_37_462 ();
 sg13g2_decap_4 FILLER_37_471 ();
 sg13g2_fill_1 FILLER_37_475 ();
 sg13g2_decap_8 FILLER_37_517 ();
 sg13g2_decap_8 FILLER_37_524 ();
 sg13g2_decap_8 FILLER_37_531 ();
 sg13g2_decap_8 FILLER_37_538 ();
 sg13g2_fill_2 FILLER_37_545 ();
 sg13g2_fill_1 FILLER_37_547 ();
 sg13g2_fill_2 FILLER_37_573 ();
 sg13g2_fill_1 FILLER_37_575 ();
 sg13g2_decap_8 FILLER_37_588 ();
 sg13g2_decap_8 FILLER_37_595 ();
 sg13g2_fill_1 FILLER_37_602 ();
 sg13g2_decap_4 FILLER_37_611 ();
 sg13g2_fill_2 FILLER_37_615 ();
 sg13g2_decap_8 FILLER_37_622 ();
 sg13g2_decap_8 FILLER_37_629 ();
 sg13g2_decap_8 FILLER_37_636 ();
 sg13g2_decap_8 FILLER_37_643 ();
 sg13g2_decap_8 FILLER_37_650 ();
 sg13g2_decap_8 FILLER_37_657 ();
 sg13g2_decap_8 FILLER_37_664 ();
 sg13g2_fill_1 FILLER_37_671 ();
 sg13g2_decap_8 FILLER_37_693 ();
 sg13g2_decap_8 FILLER_37_700 ();
 sg13g2_decap_8 FILLER_37_707 ();
 sg13g2_decap_8 FILLER_37_714 ();
 sg13g2_decap_8 FILLER_37_726 ();
 sg13g2_decap_8 FILLER_37_733 ();
 sg13g2_decap_8 FILLER_37_740 ();
 sg13g2_decap_8 FILLER_37_747 ();
 sg13g2_decap_8 FILLER_37_754 ();
 sg13g2_decap_8 FILLER_37_761 ();
 sg13g2_fill_1 FILLER_37_768 ();
 sg13g2_decap_4 FILLER_37_773 ();
 sg13g2_fill_2 FILLER_37_777 ();
 sg13g2_fill_2 FILLER_37_784 ();
 sg13g2_fill_1 FILLER_37_786 ();
 sg13g2_decap_8 FILLER_37_791 ();
 sg13g2_fill_2 FILLER_37_798 ();
 sg13g2_decap_8 FILLER_37_864 ();
 sg13g2_decap_8 FILLER_37_871 ();
 sg13g2_decap_8 FILLER_37_878 ();
 sg13g2_decap_8 FILLER_37_885 ();
 sg13g2_fill_2 FILLER_37_892 ();
 sg13g2_fill_1 FILLER_37_894 ();
 sg13g2_decap_8 FILLER_37_905 ();
 sg13g2_fill_2 FILLER_37_912 ();
 sg13g2_decap_8 FILLER_37_920 ();
 sg13g2_decap_8 FILLER_37_930 ();
 sg13g2_decap_8 FILLER_37_937 ();
 sg13g2_decap_8 FILLER_37_944 ();
 sg13g2_decap_8 FILLER_37_951 ();
 sg13g2_decap_8 FILLER_37_958 ();
 sg13g2_decap_8 FILLER_37_965 ();
 sg13g2_decap_8 FILLER_37_972 ();
 sg13g2_decap_8 FILLER_37_979 ();
 sg13g2_decap_8 FILLER_37_994 ();
 sg13g2_decap_8 FILLER_37_1001 ();
 sg13g2_decap_8 FILLER_37_1008 ();
 sg13g2_decap_8 FILLER_37_1015 ();
 sg13g2_decap_8 FILLER_37_1022 ();
 sg13g2_decap_8 FILLER_37_1029 ();
 sg13g2_decap_8 FILLER_37_1036 ();
 sg13g2_decap_8 FILLER_37_1043 ();
 sg13g2_decap_8 FILLER_37_1050 ();
 sg13g2_decap_4 FILLER_37_1057 ();
 sg13g2_fill_2 FILLER_37_1061 ();
 sg13g2_decap_8 FILLER_37_1076 ();
 sg13g2_decap_4 FILLER_37_1083 ();
 sg13g2_decap_8 FILLER_37_1113 ();
 sg13g2_decap_8 FILLER_37_1120 ();
 sg13g2_decap_8 FILLER_37_1127 ();
 sg13g2_decap_8 FILLER_37_1134 ();
 sg13g2_decap_8 FILLER_37_1141 ();
 sg13g2_fill_2 FILLER_37_1148 ();
 sg13g2_decap_8 FILLER_37_1160 ();
 sg13g2_decap_8 FILLER_37_1167 ();
 sg13g2_decap_8 FILLER_37_1174 ();
 sg13g2_decap_8 FILLER_37_1181 ();
 sg13g2_decap_8 FILLER_37_1198 ();
 sg13g2_decap_8 FILLER_37_1213 ();
 sg13g2_decap_8 FILLER_37_1220 ();
 sg13g2_decap_8 FILLER_37_1227 ();
 sg13g2_decap_8 FILLER_37_1234 ();
 sg13g2_decap_8 FILLER_37_1241 ();
 sg13g2_fill_2 FILLER_37_1248 ();
 sg13g2_decap_8 FILLER_37_1274 ();
 sg13g2_decap_8 FILLER_37_1281 ();
 sg13g2_decap_8 FILLER_37_1288 ();
 sg13g2_decap_8 FILLER_37_1295 ();
 sg13g2_decap_8 FILLER_37_1302 ();
 sg13g2_fill_1 FILLER_37_1309 ();
 sg13g2_decap_4 FILLER_37_1322 ();
 sg13g2_decap_8 FILLER_37_1352 ();
 sg13g2_decap_8 FILLER_37_1359 ();
 sg13g2_fill_2 FILLER_37_1366 ();
 sg13g2_decap_8 FILLER_37_1395 ();
 sg13g2_decap_8 FILLER_37_1402 ();
 sg13g2_decap_8 FILLER_37_1409 ();
 sg13g2_decap_8 FILLER_37_1416 ();
 sg13g2_decap_8 FILLER_37_1423 ();
 sg13g2_fill_2 FILLER_37_1430 ();
 sg13g2_fill_2 FILLER_37_1453 ();
 sg13g2_fill_1 FILLER_37_1455 ();
 sg13g2_decap_8 FILLER_37_1462 ();
 sg13g2_decap_4 FILLER_37_1486 ();
 sg13g2_fill_1 FILLER_37_1496 ();
 sg13g2_decap_8 FILLER_37_1502 ();
 sg13g2_decap_8 FILLER_37_1509 ();
 sg13g2_fill_1 FILLER_37_1516 ();
 sg13g2_fill_2 FILLER_37_1523 ();
 sg13g2_fill_2 FILLER_37_1571 ();
 sg13g2_fill_1 FILLER_37_1573 ();
 sg13g2_decap_8 FILLER_37_1600 ();
 sg13g2_decap_8 FILLER_37_1607 ();
 sg13g2_decap_8 FILLER_37_1614 ();
 sg13g2_decap_8 FILLER_37_1621 ();
 sg13g2_decap_8 FILLER_37_1650 ();
 sg13g2_decap_8 FILLER_37_1657 ();
 sg13g2_decap_8 FILLER_37_1664 ();
 sg13g2_decap_8 FILLER_37_1671 ();
 sg13g2_fill_1 FILLER_37_1678 ();
 sg13g2_decap_8 FILLER_37_1693 ();
 sg13g2_decap_8 FILLER_37_1700 ();
 sg13g2_fill_2 FILLER_37_1707 ();
 sg13g2_decap_8 FILLER_37_1736 ();
 sg13g2_decap_4 FILLER_37_1743 ();
 sg13g2_fill_1 FILLER_37_1747 ();
 sg13g2_decap_8 FILLER_37_1759 ();
 sg13g2_decap_8 FILLER_37_1766 ();
 sg13g2_fill_2 FILLER_37_1773 ();
 sg13g2_fill_1 FILLER_37_1775 ();
 sg13g2_decap_8 FILLER_37_1782 ();
 sg13g2_decap_8 FILLER_37_1789 ();
 sg13g2_decap_8 FILLER_37_1796 ();
 sg13g2_fill_2 FILLER_37_1803 ();
 sg13g2_fill_2 FILLER_37_1811 ();
 sg13g2_decap_8 FILLER_37_1819 ();
 sg13g2_decap_8 FILLER_37_1826 ();
 sg13g2_decap_8 FILLER_37_1833 ();
 sg13g2_decap_8 FILLER_37_1840 ();
 sg13g2_decap_8 FILLER_37_1847 ();
 sg13g2_decap_8 FILLER_37_1854 ();
 sg13g2_fill_2 FILLER_37_1861 ();
 sg13g2_fill_1 FILLER_37_1863 ();
 sg13g2_fill_1 FILLER_37_1872 ();
 sg13g2_fill_2 FILLER_37_1881 ();
 sg13g2_decap_8 FILLER_37_1902 ();
 sg13g2_decap_8 FILLER_37_1936 ();
 sg13g2_decap_8 FILLER_37_1943 ();
 sg13g2_decap_8 FILLER_37_1950 ();
 sg13g2_decap_8 FILLER_37_1957 ();
 sg13g2_decap_8 FILLER_37_1964 ();
 sg13g2_decap_8 FILLER_37_1971 ();
 sg13g2_decap_4 FILLER_37_1978 ();
 sg13g2_fill_1 FILLER_37_1982 ();
 sg13g2_decap_8 FILLER_37_2007 ();
 sg13g2_decap_8 FILLER_37_2014 ();
 sg13g2_decap_8 FILLER_37_2021 ();
 sg13g2_decap_4 FILLER_37_2028 ();
 sg13g2_fill_2 FILLER_37_2032 ();
 sg13g2_decap_8 FILLER_37_2044 ();
 sg13g2_decap_8 FILLER_37_2051 ();
 sg13g2_decap_8 FILLER_37_2058 ();
 sg13g2_decap_8 FILLER_37_2065 ();
 sg13g2_decap_8 FILLER_37_2072 ();
 sg13g2_decap_8 FILLER_37_2079 ();
 sg13g2_decap_8 FILLER_37_2086 ();
 sg13g2_decap_8 FILLER_37_2093 ();
 sg13g2_fill_1 FILLER_37_2112 ();
 sg13g2_decap_8 FILLER_37_2119 ();
 sg13g2_decap_8 FILLER_37_2126 ();
 sg13g2_decap_8 FILLER_37_2133 ();
 sg13g2_fill_2 FILLER_37_2140 ();
 sg13g2_decap_8 FILLER_37_2148 ();
 sg13g2_decap_8 FILLER_37_2155 ();
 sg13g2_decap_8 FILLER_37_2162 ();
 sg13g2_decap_8 FILLER_37_2169 ();
 sg13g2_decap_8 FILLER_37_2197 ();
 sg13g2_decap_8 FILLER_37_2204 ();
 sg13g2_fill_1 FILLER_37_2232 ();
 sg13g2_fill_1 FILLER_37_2239 ();
 sg13g2_fill_1 FILLER_37_2243 ();
 sg13g2_decap_8 FILLER_37_2250 ();
 sg13g2_decap_8 FILLER_37_2257 ();
 sg13g2_decap_4 FILLER_37_2264 ();
 sg13g2_fill_2 FILLER_37_2268 ();
 sg13g2_decap_8 FILLER_37_2278 ();
 sg13g2_fill_2 FILLER_37_2285 ();
 sg13g2_fill_1 FILLER_37_2287 ();
 sg13g2_fill_1 FILLER_37_2294 ();
 sg13g2_decap_8 FILLER_37_2298 ();
 sg13g2_decap_4 FILLER_37_2305 ();
 sg13g2_fill_2 FILLER_37_2309 ();
 sg13g2_decap_8 FILLER_37_2317 ();
 sg13g2_decap_8 FILLER_37_2343 ();
 sg13g2_decap_8 FILLER_37_2350 ();
 sg13g2_decap_8 FILLER_37_2357 ();
 sg13g2_decap_8 FILLER_37_2364 ();
 sg13g2_fill_1 FILLER_37_2371 ();
 sg13g2_decap_8 FILLER_37_2378 ();
 sg13g2_decap_8 FILLER_37_2385 ();
 sg13g2_decap_8 FILLER_37_2392 ();
 sg13g2_fill_2 FILLER_37_2399 ();
 sg13g2_decap_8 FILLER_37_2413 ();
 sg13g2_decap_4 FILLER_37_2420 ();
 sg13g2_fill_1 FILLER_37_2424 ();
 sg13g2_decap_8 FILLER_37_2433 ();
 sg13g2_decap_8 FILLER_37_2440 ();
 sg13g2_decap_8 FILLER_37_2447 ();
 sg13g2_decap_4 FILLER_37_2454 ();
 sg13g2_fill_1 FILLER_37_2458 ();
 sg13g2_fill_2 FILLER_37_2465 ();
 sg13g2_fill_1 FILLER_37_2467 ();
 sg13g2_decap_8 FILLER_37_2474 ();
 sg13g2_decap_4 FILLER_37_2487 ();
 sg13g2_decap_8 FILLER_37_2506 ();
 sg13g2_decap_8 FILLER_37_2513 ();
 sg13g2_fill_2 FILLER_37_2520 ();
 sg13g2_decap_8 FILLER_37_2527 ();
 sg13g2_decap_8 FILLER_37_2534 ();
 sg13g2_decap_8 FILLER_37_2541 ();
 sg13g2_decap_8 FILLER_37_2548 ();
 sg13g2_decap_4 FILLER_37_2555 ();
 sg13g2_decap_8 FILLER_37_2565 ();
 sg13g2_decap_8 FILLER_37_2572 ();
 sg13g2_fill_2 FILLER_37_2579 ();
 sg13g2_decap_8 FILLER_37_2587 ();
 sg13g2_decap_8 FILLER_37_2594 ();
 sg13g2_decap_4 FILLER_37_2601 ();
 sg13g2_fill_1 FILLER_37_2605 ();
 sg13g2_decap_8 FILLER_37_2632 ();
 sg13g2_decap_8 FILLER_37_2639 ();
 sg13g2_fill_2 FILLER_37_2646 ();
 sg13g2_fill_1 FILLER_37_2648 ();
 sg13g2_decap_4 FILLER_37_2655 ();
 sg13g2_fill_1 FILLER_37_2659 ();
 sg13g2_decap_8 FILLER_37_2665 ();
 sg13g2_decap_8 FILLER_37_2672 ();
 sg13g2_decap_8 FILLER_37_2679 ();
 sg13g2_fill_1 FILLER_37_2686 ();
 sg13g2_decap_8 FILLER_37_2697 ();
 sg13g2_decap_8 FILLER_37_2704 ();
 sg13g2_decap_8 FILLER_37_2711 ();
 sg13g2_decap_8 FILLER_37_2718 ();
 sg13g2_decap_8 FILLER_37_2725 ();
 sg13g2_decap_8 FILLER_37_2732 ();
 sg13g2_fill_1 FILLER_37_2739 ();
 sg13g2_decap_8 FILLER_37_2766 ();
 sg13g2_decap_8 FILLER_37_2773 ();
 sg13g2_decap_8 FILLER_37_2780 ();
 sg13g2_decap_8 FILLER_37_2787 ();
 sg13g2_decap_8 FILLER_37_2794 ();
 sg13g2_decap_4 FILLER_37_2801 ();
 sg13g2_fill_2 FILLER_37_2805 ();
 sg13g2_decap_4 FILLER_37_2811 ();
 sg13g2_fill_1 FILLER_37_2815 ();
 sg13g2_decap_8 FILLER_37_2834 ();
 sg13g2_decap_8 FILLER_37_2841 ();
 sg13g2_decap_8 FILLER_37_2848 ();
 sg13g2_decap_8 FILLER_37_2855 ();
 sg13g2_decap_8 FILLER_37_2862 ();
 sg13g2_decap_8 FILLER_37_2869 ();
 sg13g2_decap_8 FILLER_37_2876 ();
 sg13g2_decap_8 FILLER_37_2883 ();
 sg13g2_decap_8 FILLER_37_2890 ();
 sg13g2_decap_8 FILLER_37_2897 ();
 sg13g2_decap_8 FILLER_37_2904 ();
 sg13g2_decap_8 FILLER_37_2911 ();
 sg13g2_decap_8 FILLER_37_2918 ();
 sg13g2_decap_8 FILLER_37_2925 ();
 sg13g2_decap_4 FILLER_37_2932 ();
 sg13g2_fill_1 FILLER_37_2936 ();
 sg13g2_fill_2 FILLER_37_2942 ();
 sg13g2_fill_1 FILLER_37_2948 ();
 sg13g2_decap_8 FILLER_37_2959 ();
 sg13g2_fill_1 FILLER_37_2966 ();
 sg13g2_fill_2 FILLER_37_2977 ();
 sg13g2_fill_1 FILLER_37_2979 ();
 sg13g2_decap_8 FILLER_37_3006 ();
 sg13g2_decap_8 FILLER_37_3031 ();
 sg13g2_decap_8 FILLER_37_3038 ();
 sg13g2_decap_8 FILLER_37_3045 ();
 sg13g2_decap_8 FILLER_37_3052 ();
 sg13g2_decap_8 FILLER_37_3059 ();
 sg13g2_decap_4 FILLER_37_3066 ();
 sg13g2_fill_2 FILLER_37_3070 ();
 sg13g2_decap_8 FILLER_37_3082 ();
 sg13g2_decap_8 FILLER_37_3089 ();
 sg13g2_decap_8 FILLER_37_3096 ();
 sg13g2_decap_8 FILLER_37_3103 ();
 sg13g2_decap_8 FILLER_37_3110 ();
 sg13g2_decap_8 FILLER_37_3117 ();
 sg13g2_decap_8 FILLER_37_3124 ();
 sg13g2_decap_8 FILLER_37_3131 ();
 sg13g2_decap_8 FILLER_37_3138 ();
 sg13g2_decap_8 FILLER_37_3145 ();
 sg13g2_decap_8 FILLER_37_3152 ();
 sg13g2_decap_8 FILLER_37_3159 ();
 sg13g2_decap_8 FILLER_37_3166 ();
 sg13g2_fill_1 FILLER_37_3173 ();
 sg13g2_decap_4 FILLER_37_3184 ();
 sg13g2_fill_1 FILLER_37_3188 ();
 sg13g2_decap_8 FILLER_37_3192 ();
 sg13g2_decap_8 FILLER_37_3199 ();
 sg13g2_decap_8 FILLER_37_3206 ();
 sg13g2_decap_8 FILLER_37_3213 ();
 sg13g2_decap_8 FILLER_37_3220 ();
 sg13g2_decap_8 FILLER_37_3227 ();
 sg13g2_decap_8 FILLER_37_3234 ();
 sg13g2_decap_8 FILLER_37_3241 ();
 sg13g2_decap_8 FILLER_37_3248 ();
 sg13g2_decap_8 FILLER_37_3255 ();
 sg13g2_fill_2 FILLER_37_3262 ();
 sg13g2_fill_1 FILLER_37_3290 ();
 sg13g2_decap_8 FILLER_37_3317 ();
 sg13g2_fill_1 FILLER_37_3324 ();
 sg13g2_decap_8 FILLER_37_3361 ();
 sg13g2_decap_4 FILLER_37_3368 ();
 sg13g2_fill_1 FILLER_37_3372 ();
 sg13g2_decap_8 FILLER_37_3407 ();
 sg13g2_decap_8 FILLER_37_3414 ();
 sg13g2_decap_8 FILLER_37_3421 ();
 sg13g2_decap_8 FILLER_37_3428 ();
 sg13g2_decap_8 FILLER_37_3435 ();
 sg13g2_decap_8 FILLER_37_3442 ();
 sg13g2_decap_8 FILLER_37_3449 ();
 sg13g2_fill_2 FILLER_37_3456 ();
 sg13g2_decap_8 FILLER_37_3462 ();
 sg13g2_decap_8 FILLER_37_3469 ();
 sg13g2_decap_8 FILLER_37_3495 ();
 sg13g2_decap_8 FILLER_37_3502 ();
 sg13g2_decap_8 FILLER_37_3509 ();
 sg13g2_decap_8 FILLER_37_3516 ();
 sg13g2_decap_4 FILLER_37_3523 ();
 sg13g2_fill_2 FILLER_37_3527 ();
 sg13g2_decap_8 FILLER_37_3563 ();
 sg13g2_decap_8 FILLER_37_3570 ();
 sg13g2_fill_2 FILLER_37_3577 ();
 sg13g2_fill_1 FILLER_37_3579 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_40 ();
 sg13g2_decap_8 FILLER_38_47 ();
 sg13g2_decap_4 FILLER_38_54 ();
 sg13g2_fill_1 FILLER_38_58 ();
 sg13g2_decap_8 FILLER_38_63 ();
 sg13g2_decap_4 FILLER_38_70 ();
 sg13g2_fill_1 FILLER_38_74 ();
 sg13g2_fill_2 FILLER_38_87 ();
 sg13g2_fill_1 FILLER_38_89 ();
 sg13g2_decap_8 FILLER_38_95 ();
 sg13g2_fill_2 FILLER_38_102 ();
 sg13g2_decap_8 FILLER_38_114 ();
 sg13g2_decap_8 FILLER_38_121 ();
 sg13g2_decap_8 FILLER_38_128 ();
 sg13g2_decap_8 FILLER_38_135 ();
 sg13g2_fill_1 FILLER_38_142 ();
 sg13g2_decap_8 FILLER_38_152 ();
 sg13g2_fill_2 FILLER_38_159 ();
 sg13g2_fill_1 FILLER_38_161 ();
 sg13g2_decap_8 FILLER_38_170 ();
 sg13g2_decap_4 FILLER_38_177 ();
 sg13g2_decap_8 FILLER_38_193 ();
 sg13g2_fill_2 FILLER_38_200 ();
 sg13g2_fill_1 FILLER_38_202 ();
 sg13g2_decap_8 FILLER_38_208 ();
 sg13g2_decap_8 FILLER_38_215 ();
 sg13g2_fill_1 FILLER_38_222 ();
 sg13g2_decap_8 FILLER_38_231 ();
 sg13g2_decap_8 FILLER_38_238 ();
 sg13g2_decap_8 FILLER_38_245 ();
 sg13g2_decap_4 FILLER_38_252 ();
 sg13g2_fill_2 FILLER_38_256 ();
 sg13g2_fill_2 FILLER_38_271 ();
 sg13g2_decap_4 FILLER_38_281 ();
 sg13g2_fill_1 FILLER_38_285 ();
 sg13g2_decap_8 FILLER_38_302 ();
 sg13g2_decap_8 FILLER_38_309 ();
 sg13g2_decap_8 FILLER_38_316 ();
 sg13g2_decap_4 FILLER_38_323 ();
 sg13g2_decap_8 FILLER_38_337 ();
 sg13g2_fill_1 FILLER_38_344 ();
 sg13g2_decap_8 FILLER_38_371 ();
 sg13g2_decap_8 FILLER_38_378 ();
 sg13g2_decap_8 FILLER_38_385 ();
 sg13g2_decap_8 FILLER_38_392 ();
 sg13g2_decap_8 FILLER_38_399 ();
 sg13g2_decap_8 FILLER_38_406 ();
 sg13g2_decap_8 FILLER_38_413 ();
 sg13g2_decap_8 FILLER_38_420 ();
 sg13g2_decap_8 FILLER_38_427 ();
 sg13g2_decap_8 FILLER_38_434 ();
 sg13g2_fill_1 FILLER_38_441 ();
 sg13g2_decap_8 FILLER_38_445 ();
 sg13g2_decap_8 FILLER_38_452 ();
 sg13g2_decap_8 FILLER_38_464 ();
 sg13g2_decap_8 FILLER_38_471 ();
 sg13g2_decap_8 FILLER_38_478 ();
 sg13g2_decap_4 FILLER_38_485 ();
 sg13g2_fill_1 FILLER_38_515 ();
 sg13g2_decap_8 FILLER_38_542 ();
 sg13g2_decap_8 FILLER_38_549 ();
 sg13g2_fill_1 FILLER_38_556 ();
 sg13g2_decap_4 FILLER_38_563 ();
 sg13g2_fill_2 FILLER_38_576 ();
 sg13g2_decap_4 FILLER_38_591 ();
 sg13g2_decap_4 FILLER_38_602 ();
 sg13g2_fill_1 FILLER_38_606 ();
 sg13g2_decap_4 FILLER_38_612 ();
 sg13g2_decap_8 FILLER_38_620 ();
 sg13g2_decap_8 FILLER_38_627 ();
 sg13g2_decap_8 FILLER_38_634 ();
 sg13g2_decap_8 FILLER_38_641 ();
 sg13g2_decap_8 FILLER_38_648 ();
 sg13g2_decap_8 FILLER_38_655 ();
 sg13g2_decap_8 FILLER_38_662 ();
 sg13g2_decap_8 FILLER_38_669 ();
 sg13g2_decap_8 FILLER_38_676 ();
 sg13g2_decap_8 FILLER_38_683 ();
 sg13g2_decap_8 FILLER_38_690 ();
 sg13g2_decap_4 FILLER_38_697 ();
 sg13g2_fill_1 FILLER_38_701 ();
 sg13g2_decap_8 FILLER_38_705 ();
 sg13g2_decap_8 FILLER_38_712 ();
 sg13g2_decap_8 FILLER_38_719 ();
 sg13g2_decap_8 FILLER_38_726 ();
 sg13g2_decap_8 FILLER_38_733 ();
 sg13g2_decap_8 FILLER_38_740 ();
 sg13g2_decap_8 FILLER_38_747 ();
 sg13g2_decap_8 FILLER_38_754 ();
 sg13g2_decap_8 FILLER_38_761 ();
 sg13g2_decap_8 FILLER_38_768 ();
 sg13g2_decap_8 FILLER_38_775 ();
 sg13g2_decap_8 FILLER_38_782 ();
 sg13g2_decap_8 FILLER_38_789 ();
 sg13g2_decap_8 FILLER_38_796 ();
 sg13g2_fill_2 FILLER_38_816 ();
 sg13g2_fill_1 FILLER_38_818 ();
 sg13g2_decap_4 FILLER_38_831 ();
 sg13g2_decap_8 FILLER_38_841 ();
 sg13g2_decap_8 FILLER_38_848 ();
 sg13g2_decap_8 FILLER_38_855 ();
 sg13g2_decap_8 FILLER_38_862 ();
 sg13g2_decap_8 FILLER_38_869 ();
 sg13g2_decap_8 FILLER_38_876 ();
 sg13g2_decap_8 FILLER_38_883 ();
 sg13g2_fill_2 FILLER_38_890 ();
 sg13g2_fill_1 FILLER_38_892 ();
 sg13g2_fill_2 FILLER_38_912 ();
 sg13g2_decap_8 FILLER_38_962 ();
 sg13g2_decap_8 FILLER_38_969 ();
 sg13g2_decap_8 FILLER_38_976 ();
 sg13g2_fill_1 FILLER_38_983 ();
 sg13g2_decap_8 FILLER_38_1014 ();
 sg13g2_decap_8 FILLER_38_1021 ();
 sg13g2_decap_8 FILLER_38_1028 ();
 sg13g2_decap_8 FILLER_38_1035 ();
 sg13g2_decap_4 FILLER_38_1042 ();
 sg13g2_decap_8 FILLER_38_1066 ();
 sg13g2_decap_8 FILLER_38_1073 ();
 sg13g2_fill_2 FILLER_38_1080 ();
 sg13g2_fill_1 FILLER_38_1082 ();
 sg13g2_decap_8 FILLER_38_1093 ();
 sg13g2_decap_8 FILLER_38_1100 ();
 sg13g2_decap_8 FILLER_38_1107 ();
 sg13g2_decap_4 FILLER_38_1114 ();
 sg13g2_fill_2 FILLER_38_1118 ();
 sg13g2_decap_8 FILLER_38_1130 ();
 sg13g2_fill_2 FILLER_38_1137 ();
 sg13g2_fill_1 FILLER_38_1139 ();
 sg13g2_decap_8 FILLER_38_1166 ();
 sg13g2_decap_8 FILLER_38_1173 ();
 sg13g2_decap_8 FILLER_38_1180 ();
 sg13g2_decap_8 FILLER_38_1187 ();
 sg13g2_fill_1 FILLER_38_1194 ();
 sg13g2_decap_8 FILLER_38_1221 ();
 sg13g2_decap_8 FILLER_38_1228 ();
 sg13g2_decap_8 FILLER_38_1235 ();
 sg13g2_decap_8 FILLER_38_1242 ();
 sg13g2_decap_8 FILLER_38_1249 ();
 sg13g2_fill_2 FILLER_38_1256 ();
 sg13g2_decap_8 FILLER_38_1261 ();
 sg13g2_decap_8 FILLER_38_1268 ();
 sg13g2_decap_8 FILLER_38_1275 ();
 sg13g2_decap_8 FILLER_38_1282 ();
 sg13g2_decap_8 FILLER_38_1289 ();
 sg13g2_decap_8 FILLER_38_1296 ();
 sg13g2_decap_8 FILLER_38_1303 ();
 sg13g2_decap_8 FILLER_38_1310 ();
 sg13g2_decap_8 FILLER_38_1317 ();
 sg13g2_decap_8 FILLER_38_1324 ();
 sg13g2_decap_8 FILLER_38_1331 ();
 sg13g2_fill_1 FILLER_38_1338 ();
 sg13g2_decap_8 FILLER_38_1345 ();
 sg13g2_decap_8 FILLER_38_1352 ();
 sg13g2_decap_8 FILLER_38_1359 ();
 sg13g2_decap_8 FILLER_38_1366 ();
 sg13g2_decap_4 FILLER_38_1373 ();
 sg13g2_fill_2 FILLER_38_1377 ();
 sg13g2_fill_1 FILLER_38_1385 ();
 sg13g2_decap_8 FILLER_38_1400 ();
 sg13g2_decap_8 FILLER_38_1407 ();
 sg13g2_decap_8 FILLER_38_1414 ();
 sg13g2_decap_8 FILLER_38_1421 ();
 sg13g2_decap_8 FILLER_38_1428 ();
 sg13g2_fill_2 FILLER_38_1435 ();
 sg13g2_fill_1 FILLER_38_1437 ();
 sg13g2_decap_8 FILLER_38_1441 ();
 sg13g2_decap_8 FILLER_38_1448 ();
 sg13g2_decap_8 FILLER_38_1455 ();
 sg13g2_fill_2 FILLER_38_1462 ();
 sg13g2_fill_2 FILLER_38_1478 ();
 sg13g2_fill_1 FILLER_38_1486 ();
 sg13g2_decap_8 FILLER_38_1493 ();
 sg13g2_decap_8 FILLER_38_1500 ();
 sg13g2_decap_8 FILLER_38_1507 ();
 sg13g2_decap_8 FILLER_38_1514 ();
 sg13g2_decap_8 FILLER_38_1521 ();
 sg13g2_decap_8 FILLER_38_1528 ();
 sg13g2_decap_4 FILLER_38_1535 ();
 sg13g2_decap_8 FILLER_38_1549 ();
 sg13g2_decap_4 FILLER_38_1559 ();
 sg13g2_fill_1 FILLER_38_1563 ();
 sg13g2_decap_8 FILLER_38_1568 ();
 sg13g2_decap_8 FILLER_38_1575 ();
 sg13g2_decap_8 FILLER_38_1582 ();
 sg13g2_fill_2 FILLER_38_1589 ();
 sg13g2_fill_1 FILLER_38_1591 ();
 sg13g2_decap_8 FILLER_38_1596 ();
 sg13g2_decap_8 FILLER_38_1603 ();
 sg13g2_decap_8 FILLER_38_1610 ();
 sg13g2_fill_2 FILLER_38_1617 ();
 sg13g2_fill_1 FILLER_38_1619 ();
 sg13g2_decap_8 FILLER_38_1647 ();
 sg13g2_decap_8 FILLER_38_1654 ();
 sg13g2_decap_8 FILLER_38_1661 ();
 sg13g2_fill_2 FILLER_38_1668 ();
 sg13g2_decap_8 FILLER_38_1687 ();
 sg13g2_decap_8 FILLER_38_1694 ();
 sg13g2_decap_8 FILLER_38_1701 ();
 sg13g2_decap_8 FILLER_38_1708 ();
 sg13g2_fill_2 FILLER_38_1715 ();
 sg13g2_fill_1 FILLER_38_1717 ();
 sg13g2_decap_8 FILLER_38_1727 ();
 sg13g2_decap_8 FILLER_38_1734 ();
 sg13g2_decap_8 FILLER_38_1741 ();
 sg13g2_decap_8 FILLER_38_1748 ();
 sg13g2_fill_1 FILLER_38_1755 ();
 sg13g2_decap_8 FILLER_38_1761 ();
 sg13g2_decap_8 FILLER_38_1768 ();
 sg13g2_decap_8 FILLER_38_1775 ();
 sg13g2_decap_4 FILLER_38_1782 ();
 sg13g2_fill_2 FILLER_38_1786 ();
 sg13g2_decap_8 FILLER_38_1794 ();
 sg13g2_decap_8 FILLER_38_1801 ();
 sg13g2_decap_8 FILLER_38_1808 ();
 sg13g2_decap_8 FILLER_38_1815 ();
 sg13g2_decap_8 FILLER_38_1822 ();
 sg13g2_decap_8 FILLER_38_1829 ();
 sg13g2_decap_4 FILLER_38_1836 ();
 sg13g2_fill_2 FILLER_38_1840 ();
 sg13g2_decap_8 FILLER_38_1848 ();
 sg13g2_decap_4 FILLER_38_1855 ();
 sg13g2_fill_2 FILLER_38_1859 ();
 sg13g2_decap_4 FILLER_38_1877 ();
 sg13g2_fill_2 FILLER_38_1881 ();
 sg13g2_decap_8 FILLER_38_1886 ();
 sg13g2_decap_8 FILLER_38_1893 ();
 sg13g2_decap_8 FILLER_38_1900 ();
 sg13g2_decap_8 FILLER_38_1927 ();
 sg13g2_decap_8 FILLER_38_1934 ();
 sg13g2_decap_8 FILLER_38_1941 ();
 sg13g2_decap_8 FILLER_38_1948 ();
 sg13g2_decap_4 FILLER_38_1955 ();
 sg13g2_fill_1 FILLER_38_1959 ();
 sg13g2_decap_4 FILLER_38_1984 ();
 sg13g2_fill_1 FILLER_38_1988 ();
 sg13g2_decap_8 FILLER_38_1995 ();
 sg13g2_decap_8 FILLER_38_2002 ();
 sg13g2_decap_8 FILLER_38_2009 ();
 sg13g2_decap_8 FILLER_38_2016 ();
 sg13g2_decap_4 FILLER_38_2023 ();
 sg13g2_fill_2 FILLER_38_2027 ();
 sg13g2_decap_8 FILLER_38_2039 ();
 sg13g2_decap_8 FILLER_38_2046 ();
 sg13g2_decap_8 FILLER_38_2053 ();
 sg13g2_decap_8 FILLER_38_2060 ();
 sg13g2_decap_8 FILLER_38_2067 ();
 sg13g2_fill_2 FILLER_38_2074 ();
 sg13g2_fill_1 FILLER_38_2076 ();
 sg13g2_decap_8 FILLER_38_2089 ();
 sg13g2_decap_8 FILLER_38_2096 ();
 sg13g2_decap_8 FILLER_38_2103 ();
 sg13g2_decap_8 FILLER_38_2110 ();
 sg13g2_decap_4 FILLER_38_2117 ();
 sg13g2_fill_2 FILLER_38_2121 ();
 sg13g2_decap_8 FILLER_38_2132 ();
 sg13g2_decap_8 FILLER_38_2139 ();
 sg13g2_decap_8 FILLER_38_2146 ();
 sg13g2_decap_8 FILLER_38_2153 ();
 sg13g2_decap_8 FILLER_38_2160 ();
 sg13g2_decap_8 FILLER_38_2167 ();
 sg13g2_decap_4 FILLER_38_2174 ();
 sg13g2_fill_2 FILLER_38_2210 ();
 sg13g2_fill_1 FILLER_38_2212 ();
 sg13g2_fill_1 FILLER_38_2219 ();
 sg13g2_fill_1 FILLER_38_2232 ();
 sg13g2_fill_1 FILLER_38_2243 ();
 sg13g2_decap_8 FILLER_38_2255 ();
 sg13g2_decap_8 FILLER_38_2276 ();
 sg13g2_fill_1 FILLER_38_2283 ();
 sg13g2_fill_2 FILLER_38_2305 ();
 sg13g2_fill_1 FILLER_38_2307 ();
 sg13g2_decap_8 FILLER_38_2314 ();
 sg13g2_decap_8 FILLER_38_2321 ();
 sg13g2_decap_8 FILLER_38_2328 ();
 sg13g2_fill_1 FILLER_38_2335 ();
 sg13g2_decap_8 FILLER_38_2342 ();
 sg13g2_fill_2 FILLER_38_2349 ();
 sg13g2_decap_4 FILLER_38_2357 ();
 sg13g2_decap_4 FILLER_38_2367 ();
 sg13g2_decap_4 FILLER_38_2376 ();
 sg13g2_decap_8 FILLER_38_2386 ();
 sg13g2_decap_8 FILLER_38_2393 ();
 sg13g2_decap_8 FILLER_38_2405 ();
 sg13g2_decap_8 FILLER_38_2412 ();
 sg13g2_decap_8 FILLER_38_2419 ();
 sg13g2_decap_4 FILLER_38_2426 ();
 sg13g2_fill_1 FILLER_38_2430 ();
 sg13g2_decap_8 FILLER_38_2437 ();
 sg13g2_decap_4 FILLER_38_2444 ();
 sg13g2_fill_2 FILLER_38_2448 ();
 sg13g2_decap_8 FILLER_38_2458 ();
 sg13g2_decap_8 FILLER_38_2465 ();
 sg13g2_decap_8 FILLER_38_2472 ();
 sg13g2_decap_8 FILLER_38_2479 ();
 sg13g2_decap_8 FILLER_38_2486 ();
 sg13g2_decap_8 FILLER_38_2499 ();
 sg13g2_decap_8 FILLER_38_2506 ();
 sg13g2_decap_4 FILLER_38_2513 ();
 sg13g2_decap_8 FILLER_38_2541 ();
 sg13g2_decap_8 FILLER_38_2548 ();
 sg13g2_fill_2 FILLER_38_2555 ();
 sg13g2_decap_8 FILLER_38_2589 ();
 sg13g2_decap_8 FILLER_38_2596 ();
 sg13g2_decap_8 FILLER_38_2603 ();
 sg13g2_decap_8 FILLER_38_2620 ();
 sg13g2_decap_8 FILLER_38_2627 ();
 sg13g2_fill_2 FILLER_38_2634 ();
 sg13g2_decap_8 FILLER_38_2644 ();
 sg13g2_decap_4 FILLER_38_2651 ();
 sg13g2_fill_2 FILLER_38_2655 ();
 sg13g2_decap_8 FILLER_38_2668 ();
 sg13g2_decap_8 FILLER_38_2675 ();
 sg13g2_fill_2 FILLER_38_2682 ();
 sg13g2_decap_8 FILLER_38_2727 ();
 sg13g2_decap_8 FILLER_38_2734 ();
 sg13g2_decap_8 FILLER_38_2741 ();
 sg13g2_decap_8 FILLER_38_2748 ();
 sg13g2_decap_4 FILLER_38_2755 ();
 sg13g2_fill_1 FILLER_38_2759 ();
 sg13g2_decap_8 FILLER_38_2765 ();
 sg13g2_decap_8 FILLER_38_2772 ();
 sg13g2_decap_8 FILLER_38_2779 ();
 sg13g2_decap_8 FILLER_38_2786 ();
 sg13g2_decap_8 FILLER_38_2793 ();
 sg13g2_decap_8 FILLER_38_2800 ();
 sg13g2_decap_8 FILLER_38_2807 ();
 sg13g2_decap_8 FILLER_38_2814 ();
 sg13g2_fill_2 FILLER_38_2821 ();
 sg13g2_decap_8 FILLER_38_2833 ();
 sg13g2_decap_8 FILLER_38_2840 ();
 sg13g2_decap_8 FILLER_38_2847 ();
 sg13g2_decap_8 FILLER_38_2854 ();
 sg13g2_decap_8 FILLER_38_2861 ();
 sg13g2_decap_8 FILLER_38_2868 ();
 sg13g2_decap_8 FILLER_38_2875 ();
 sg13g2_decap_8 FILLER_38_2882 ();
 sg13g2_decap_8 FILLER_38_2889 ();
 sg13g2_decap_8 FILLER_38_2896 ();
 sg13g2_decap_8 FILLER_38_2903 ();
 sg13g2_decap_8 FILLER_38_2910 ();
 sg13g2_decap_8 FILLER_38_2917 ();
 sg13g2_decap_8 FILLER_38_2924 ();
 sg13g2_decap_8 FILLER_38_2931 ();
 sg13g2_decap_8 FILLER_38_2938 ();
 sg13g2_decap_8 FILLER_38_2945 ();
 sg13g2_decap_8 FILLER_38_2952 ();
 sg13g2_decap_8 FILLER_38_2959 ();
 sg13g2_decap_8 FILLER_38_2966 ();
 sg13g2_decap_8 FILLER_38_2973 ();
 sg13g2_decap_8 FILLER_38_2980 ();
 sg13g2_decap_4 FILLER_38_2987 ();
 sg13g2_decap_4 FILLER_38_3001 ();
 sg13g2_fill_1 FILLER_38_3005 ();
 sg13g2_decap_8 FILLER_38_3032 ();
 sg13g2_decap_8 FILLER_38_3039 ();
 sg13g2_decap_8 FILLER_38_3046 ();
 sg13g2_decap_8 FILLER_38_3053 ();
 sg13g2_decap_4 FILLER_38_3060 ();
 sg13g2_fill_1 FILLER_38_3064 ();
 sg13g2_decap_8 FILLER_38_3085 ();
 sg13g2_decap_8 FILLER_38_3092 ();
 sg13g2_decap_8 FILLER_38_3099 ();
 sg13g2_decap_8 FILLER_38_3106 ();
 sg13g2_decap_8 FILLER_38_3113 ();
 sg13g2_decap_8 FILLER_38_3120 ();
 sg13g2_decap_8 FILLER_38_3127 ();
 sg13g2_decap_8 FILLER_38_3134 ();
 sg13g2_decap_8 FILLER_38_3141 ();
 sg13g2_fill_2 FILLER_38_3148 ();
 sg13g2_decap_8 FILLER_38_3176 ();
 sg13g2_decap_4 FILLER_38_3183 ();
 sg13g2_fill_2 FILLER_38_3187 ();
 sg13g2_decap_4 FILLER_38_3199 ();
 sg13g2_decap_8 FILLER_38_3229 ();
 sg13g2_decap_8 FILLER_38_3236 ();
 sg13g2_decap_8 FILLER_38_3243 ();
 sg13g2_decap_4 FILLER_38_3250 ();
 sg13g2_decap_4 FILLER_38_3260 ();
 sg13g2_decap_8 FILLER_38_3272 ();
 sg13g2_decap_8 FILLER_38_3279 ();
 sg13g2_decap_8 FILLER_38_3286 ();
 sg13g2_decap_4 FILLER_38_3293 ();
 sg13g2_fill_1 FILLER_38_3297 ();
 sg13g2_decap_8 FILLER_38_3303 ();
 sg13g2_decap_8 FILLER_38_3310 ();
 sg13g2_decap_8 FILLER_38_3317 ();
 sg13g2_decap_8 FILLER_38_3324 ();
 sg13g2_decap_8 FILLER_38_3331 ();
 sg13g2_fill_2 FILLER_38_3338 ();
 sg13g2_fill_1 FILLER_38_3340 ();
 sg13g2_decap_8 FILLER_38_3349 ();
 sg13g2_decap_4 FILLER_38_3356 ();
 sg13g2_fill_2 FILLER_38_3360 ();
 sg13g2_decap_8 FILLER_38_3367 ();
 sg13g2_decap_8 FILLER_38_3374 ();
 sg13g2_decap_8 FILLER_38_3381 ();
 sg13g2_decap_8 FILLER_38_3388 ();
 sg13g2_decap_8 FILLER_38_3395 ();
 sg13g2_decap_8 FILLER_38_3402 ();
 sg13g2_decap_8 FILLER_38_3409 ();
 sg13g2_decap_8 FILLER_38_3416 ();
 sg13g2_decap_8 FILLER_38_3423 ();
 sg13g2_decap_8 FILLER_38_3430 ();
 sg13g2_fill_2 FILLER_38_3437 ();
 sg13g2_decap_8 FILLER_38_3473 ();
 sg13g2_fill_1 FILLER_38_3480 ();
 sg13g2_decap_8 FILLER_38_3507 ();
 sg13g2_decap_8 FILLER_38_3523 ();
 sg13g2_decap_4 FILLER_38_3530 ();
 sg13g2_fill_1 FILLER_38_3534 ();
 sg13g2_decap_8 FILLER_38_3569 ();
 sg13g2_decap_4 FILLER_38_3576 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_50 ();
 sg13g2_decap_8 FILLER_39_57 ();
 sg13g2_decap_8 FILLER_39_64 ();
 sg13g2_decap_8 FILLER_39_71 ();
 sg13g2_fill_2 FILLER_39_78 ();
 sg13g2_decap_4 FILLER_39_84 ();
 sg13g2_fill_1 FILLER_39_88 ();
 sg13g2_decap_8 FILLER_39_112 ();
 sg13g2_decap_8 FILLER_39_119 ();
 sg13g2_decap_8 FILLER_39_126 ();
 sg13g2_decap_8 FILLER_39_133 ();
 sg13g2_decap_8 FILLER_39_140 ();
 sg13g2_decap_8 FILLER_39_147 ();
 sg13g2_decap_4 FILLER_39_154 ();
 sg13g2_fill_1 FILLER_39_158 ();
 sg13g2_fill_2 FILLER_39_164 ();
 sg13g2_decap_8 FILLER_39_170 ();
 sg13g2_decap_8 FILLER_39_177 ();
 sg13g2_decap_4 FILLER_39_184 ();
 sg13g2_fill_2 FILLER_39_188 ();
 sg13g2_decap_8 FILLER_39_198 ();
 sg13g2_decap_8 FILLER_39_205 ();
 sg13g2_fill_2 FILLER_39_212 ();
 sg13g2_decap_8 FILLER_39_224 ();
 sg13g2_decap_8 FILLER_39_231 ();
 sg13g2_decap_8 FILLER_39_238 ();
 sg13g2_decap_8 FILLER_39_245 ();
 sg13g2_decap_8 FILLER_39_252 ();
 sg13g2_decap_8 FILLER_39_259 ();
 sg13g2_fill_2 FILLER_39_266 ();
 sg13g2_fill_1 FILLER_39_268 ();
 sg13g2_decap_4 FILLER_39_282 ();
 sg13g2_decap_4 FILLER_39_299 ();
 sg13g2_decap_8 FILLER_39_329 ();
 sg13g2_decap_8 FILLER_39_362 ();
 sg13g2_decap_4 FILLER_39_369 ();
 sg13g2_decap_8 FILLER_39_381 ();
 sg13g2_decap_8 FILLER_39_388 ();
 sg13g2_decap_8 FILLER_39_395 ();
 sg13g2_fill_2 FILLER_39_402 ();
 sg13g2_fill_1 FILLER_39_404 ();
 sg13g2_decap_4 FILLER_39_437 ();
 sg13g2_fill_2 FILLER_39_441 ();
 sg13g2_decap_8 FILLER_39_448 ();
 sg13g2_decap_8 FILLER_39_455 ();
 sg13g2_fill_2 FILLER_39_462 ();
 sg13g2_decap_4 FILLER_39_472 ();
 sg13g2_fill_2 FILLER_39_476 ();
 sg13g2_decap_8 FILLER_39_486 ();
 sg13g2_decap_4 FILLER_39_493 ();
 sg13g2_fill_2 FILLER_39_497 ();
 sg13g2_decap_8 FILLER_39_521 ();
 sg13g2_fill_1 FILLER_39_528 ();
 sg13g2_decap_8 FILLER_39_538 ();
 sg13g2_decap_8 FILLER_39_545 ();
 sg13g2_fill_2 FILLER_39_552 ();
 sg13g2_fill_1 FILLER_39_554 ();
 sg13g2_fill_1 FILLER_39_561 ();
 sg13g2_fill_1 FILLER_39_582 ();
 sg13g2_decap_8 FILLER_39_590 ();
 sg13g2_decap_8 FILLER_39_597 ();
 sg13g2_decap_4 FILLER_39_604 ();
 sg13g2_fill_1 FILLER_39_634 ();
 sg13g2_decap_8 FILLER_39_643 ();
 sg13g2_decap_8 FILLER_39_650 ();
 sg13g2_decap_8 FILLER_39_657 ();
 sg13g2_decap_8 FILLER_39_664 ();
 sg13g2_decap_8 FILLER_39_671 ();
 sg13g2_decap_8 FILLER_39_678 ();
 sg13g2_decap_8 FILLER_39_685 ();
 sg13g2_decap_8 FILLER_39_692 ();
 sg13g2_decap_8 FILLER_39_708 ();
 sg13g2_decap_8 FILLER_39_715 ();
 sg13g2_decap_8 FILLER_39_722 ();
 sg13g2_decap_8 FILLER_39_729 ();
 sg13g2_decap_8 FILLER_39_736 ();
 sg13g2_decap_8 FILLER_39_743 ();
 sg13g2_fill_2 FILLER_39_750 ();
 sg13g2_fill_1 FILLER_39_752 ();
 sg13g2_fill_1 FILLER_39_760 ();
 sg13g2_decap_8 FILLER_39_768 ();
 sg13g2_decap_8 FILLER_39_779 ();
 sg13g2_decap_8 FILLER_39_786 ();
 sg13g2_decap_8 FILLER_39_793 ();
 sg13g2_decap_8 FILLER_39_800 ();
 sg13g2_decap_8 FILLER_39_807 ();
 sg13g2_decap_8 FILLER_39_814 ();
 sg13g2_decap_8 FILLER_39_821 ();
 sg13g2_decap_8 FILLER_39_828 ();
 sg13g2_decap_8 FILLER_39_835 ();
 sg13g2_decap_8 FILLER_39_842 ();
 sg13g2_decap_8 FILLER_39_849 ();
 sg13g2_decap_4 FILLER_39_856 ();
 sg13g2_fill_2 FILLER_39_864 ();
 sg13g2_fill_2 FILLER_39_875 ();
 sg13g2_decap_4 FILLER_39_890 ();
 sg13g2_fill_1 FILLER_39_894 ();
 sg13g2_decap_8 FILLER_39_908 ();
 sg13g2_decap_8 FILLER_39_915 ();
 sg13g2_decap_8 FILLER_39_922 ();
 sg13g2_decap_4 FILLER_39_929 ();
 sg13g2_decap_4 FILLER_39_941 ();
 sg13g2_decap_8 FILLER_39_950 ();
 sg13g2_decap_8 FILLER_39_957 ();
 sg13g2_decap_8 FILLER_39_964 ();
 sg13g2_decap_4 FILLER_39_971 ();
 sg13g2_fill_1 FILLER_39_975 ();
 sg13g2_decap_8 FILLER_39_986 ();
 sg13g2_decap_4 FILLER_39_993 ();
 sg13g2_fill_2 FILLER_39_997 ();
 sg13g2_decap_8 FILLER_39_1027 ();
 sg13g2_decap_8 FILLER_39_1034 ();
 sg13g2_fill_2 FILLER_39_1041 ();
 sg13g2_decap_8 FILLER_39_1069 ();
 sg13g2_decap_8 FILLER_39_1076 ();
 sg13g2_decap_8 FILLER_39_1083 ();
 sg13g2_decap_8 FILLER_39_1090 ();
 sg13g2_fill_2 FILLER_39_1097 ();
 sg13g2_fill_2 FILLER_39_1107 ();
 sg13g2_fill_1 FILLER_39_1109 ();
 sg13g2_fill_1 FILLER_39_1118 ();
 sg13g2_decap_8 FILLER_39_1132 ();
 sg13g2_fill_1 FILLER_39_1139 ();
 sg13g2_decap_8 FILLER_39_1166 ();
 sg13g2_decap_8 FILLER_39_1173 ();
 sg13g2_decap_8 FILLER_39_1180 ();
 sg13g2_decap_8 FILLER_39_1187 ();
 sg13g2_decap_8 FILLER_39_1194 ();
 sg13g2_decap_8 FILLER_39_1201 ();
 sg13g2_decap_8 FILLER_39_1208 ();
 sg13g2_fill_2 FILLER_39_1215 ();
 sg13g2_fill_1 FILLER_39_1217 ();
 sg13g2_decap_8 FILLER_39_1228 ();
 sg13g2_decap_8 FILLER_39_1235 ();
 sg13g2_decap_8 FILLER_39_1242 ();
 sg13g2_decap_8 FILLER_39_1249 ();
 sg13g2_decap_8 FILLER_39_1256 ();
 sg13g2_decap_8 FILLER_39_1263 ();
 sg13g2_fill_1 FILLER_39_1270 ();
 sg13g2_fill_2 FILLER_39_1281 ();
 sg13g2_fill_1 FILLER_39_1283 ();
 sg13g2_decap_8 FILLER_39_1315 ();
 sg13g2_decap_8 FILLER_39_1322 ();
 sg13g2_decap_8 FILLER_39_1329 ();
 sg13g2_decap_8 FILLER_39_1336 ();
 sg13g2_decap_8 FILLER_39_1343 ();
 sg13g2_decap_8 FILLER_39_1350 ();
 sg13g2_decap_8 FILLER_39_1369 ();
 sg13g2_decap_8 FILLER_39_1376 ();
 sg13g2_decap_8 FILLER_39_1383 ();
 sg13g2_decap_8 FILLER_39_1390 ();
 sg13g2_decap_8 FILLER_39_1397 ();
 sg13g2_decap_8 FILLER_39_1430 ();
 sg13g2_fill_1 FILLER_39_1437 ();
 sg13g2_fill_1 FILLER_39_1457 ();
 sg13g2_decap_8 FILLER_39_1466 ();
 sg13g2_decap_4 FILLER_39_1473 ();
 sg13g2_fill_1 FILLER_39_1477 ();
 sg13g2_decap_8 FILLER_39_1482 ();
 sg13g2_decap_8 FILLER_39_1489 ();
 sg13g2_fill_2 FILLER_39_1496 ();
 sg13g2_decap_8 FILLER_39_1504 ();
 sg13g2_decap_8 FILLER_39_1511 ();
 sg13g2_decap_8 FILLER_39_1518 ();
 sg13g2_decap_8 FILLER_39_1525 ();
 sg13g2_decap_8 FILLER_39_1532 ();
 sg13g2_decap_8 FILLER_39_1539 ();
 sg13g2_decap_8 FILLER_39_1546 ();
 sg13g2_decap_8 FILLER_39_1553 ();
 sg13g2_decap_8 FILLER_39_1560 ();
 sg13g2_decap_8 FILLER_39_1567 ();
 sg13g2_decap_8 FILLER_39_1574 ();
 sg13g2_decap_8 FILLER_39_1581 ();
 sg13g2_decap_8 FILLER_39_1588 ();
 sg13g2_decap_8 FILLER_39_1595 ();
 sg13g2_decap_8 FILLER_39_1602 ();
 sg13g2_decap_8 FILLER_39_1609 ();
 sg13g2_fill_1 FILLER_39_1616 ();
 sg13g2_decap_8 FILLER_39_1651 ();
 sg13g2_decap_8 FILLER_39_1658 ();
 sg13g2_decap_4 FILLER_39_1665 ();
 sg13g2_fill_1 FILLER_39_1669 ();
 sg13g2_decap_8 FILLER_39_1681 ();
 sg13g2_fill_1 FILLER_39_1688 ();
 sg13g2_decap_4 FILLER_39_1711 ();
 sg13g2_fill_2 FILLER_39_1715 ();
 sg13g2_decap_8 FILLER_39_1723 ();
 sg13g2_decap_8 FILLER_39_1730 ();
 sg13g2_decap_8 FILLER_39_1737 ();
 sg13g2_fill_2 FILLER_39_1744 ();
 sg13g2_fill_1 FILLER_39_1746 ();
 sg13g2_decap_8 FILLER_39_1782 ();
 sg13g2_decap_8 FILLER_39_1789 ();
 sg13g2_decap_8 FILLER_39_1796 ();
 sg13g2_decap_8 FILLER_39_1835 ();
 sg13g2_decap_8 FILLER_39_1842 ();
 sg13g2_decap_8 FILLER_39_1849 ();
 sg13g2_fill_2 FILLER_39_1856 ();
 sg13g2_fill_1 FILLER_39_1858 ();
 sg13g2_fill_2 FILLER_39_1879 ();
 sg13g2_fill_1 FILLER_39_1881 ();
 sg13g2_fill_1 FILLER_39_1895 ();
 sg13g2_decap_8 FILLER_39_1902 ();
 sg13g2_decap_4 FILLER_39_1909 ();
 sg13g2_fill_1 FILLER_39_1919 ();
 sg13g2_decap_8 FILLER_39_1926 ();
 sg13g2_decap_4 FILLER_39_1933 ();
 sg13g2_fill_1 FILLER_39_1937 ();
 sg13g2_decap_8 FILLER_39_1941 ();
 sg13g2_fill_2 FILLER_39_1948 ();
 sg13g2_decap_4 FILLER_39_1959 ();
 sg13g2_fill_1 FILLER_39_1963 ();
 sg13g2_decap_8 FILLER_39_1967 ();
 sg13g2_fill_1 FILLER_39_1974 ();
 sg13g2_decap_8 FILLER_39_1981 ();
 sg13g2_fill_2 FILLER_39_1988 ();
 sg13g2_fill_1 FILLER_39_1990 ();
 sg13g2_decap_8 FILLER_39_1997 ();
 sg13g2_decap_8 FILLER_39_2004 ();
 sg13g2_decap_8 FILLER_39_2011 ();
 sg13g2_fill_2 FILLER_39_2018 ();
 sg13g2_fill_1 FILLER_39_2020 ();
 sg13g2_decap_8 FILLER_39_2024 ();
 sg13g2_fill_1 FILLER_39_2031 ();
 sg13g2_fill_1 FILLER_39_2066 ();
 sg13g2_decap_4 FILLER_39_2073 ();
 sg13g2_decap_4 FILLER_39_2082 ();
 sg13g2_fill_1 FILLER_39_2086 ();
 sg13g2_decap_8 FILLER_39_2093 ();
 sg13g2_decap_8 FILLER_39_2100 ();
 sg13g2_decap_8 FILLER_39_2107 ();
 sg13g2_fill_2 FILLER_39_2114 ();
 sg13g2_fill_1 FILLER_39_2116 ();
 sg13g2_fill_1 FILLER_39_2135 ();
 sg13g2_fill_2 FILLER_39_2154 ();
 sg13g2_fill_1 FILLER_39_2156 ();
 sg13g2_decap_8 FILLER_39_2163 ();
 sg13g2_fill_2 FILLER_39_2170 ();
 sg13g2_fill_2 FILLER_39_2195 ();
 sg13g2_fill_1 FILLER_39_2197 ();
 sg13g2_decap_8 FILLER_39_2204 ();
 sg13g2_decap_8 FILLER_39_2211 ();
 sg13g2_fill_2 FILLER_39_2218 ();
 sg13g2_fill_1 FILLER_39_2220 ();
 sg13g2_decap_8 FILLER_39_2254 ();
 sg13g2_decap_8 FILLER_39_2261 ();
 sg13g2_fill_2 FILLER_39_2280 ();
 sg13g2_fill_1 FILLER_39_2294 ();
 sg13g2_decap_8 FILLER_39_2301 ();
 sg13g2_decap_8 FILLER_39_2308 ();
 sg13g2_decap_8 FILLER_39_2315 ();
 sg13g2_decap_8 FILLER_39_2322 ();
 sg13g2_decap_8 FILLER_39_2329 ();
 sg13g2_fill_2 FILLER_39_2336 ();
 sg13g2_fill_1 FILLER_39_2338 ();
 sg13g2_decap_4 FILLER_39_2347 ();
 sg13g2_decap_8 FILLER_39_2363 ();
 sg13g2_decap_8 FILLER_39_2370 ();
 sg13g2_decap_8 FILLER_39_2377 ();
 sg13g2_fill_1 FILLER_39_2384 ();
 sg13g2_fill_2 FILLER_39_2403 ();
 sg13g2_decap_8 FILLER_39_2431 ();
 sg13g2_fill_2 FILLER_39_2438 ();
 sg13g2_fill_1 FILLER_39_2440 ();
 sg13g2_decap_8 FILLER_39_2447 ();
 sg13g2_decap_8 FILLER_39_2454 ();
 sg13g2_decap_4 FILLER_39_2461 ();
 sg13g2_fill_1 FILLER_39_2465 ();
 sg13g2_decap_8 FILLER_39_2482 ();
 sg13g2_decap_8 FILLER_39_2489 ();
 sg13g2_decap_8 FILLER_39_2496 ();
 sg13g2_decap_8 FILLER_39_2503 ();
 sg13g2_decap_8 FILLER_39_2529 ();
 sg13g2_decap_4 FILLER_39_2536 ();
 sg13g2_fill_1 FILLER_39_2540 ();
 sg13g2_decap_8 FILLER_39_2547 ();
 sg13g2_decap_8 FILLER_39_2554 ();
 sg13g2_decap_4 FILLER_39_2561 ();
 sg13g2_fill_2 FILLER_39_2565 ();
 sg13g2_decap_8 FILLER_39_2577 ();
 sg13g2_decap_8 FILLER_39_2584 ();
 sg13g2_decap_8 FILLER_39_2591 ();
 sg13g2_decap_4 FILLER_39_2604 ();
 sg13g2_decap_8 FILLER_39_2634 ();
 sg13g2_decap_8 FILLER_39_2641 ();
 sg13g2_decap_8 FILLER_39_2648 ();
 sg13g2_fill_1 FILLER_39_2655 ();
 sg13g2_fill_2 FILLER_39_2682 ();
 sg13g2_decap_4 FILLER_39_2735 ();
 sg13g2_decap_8 FILLER_39_2742 ();
 sg13g2_decap_8 FILLER_39_2749 ();
 sg13g2_decap_4 FILLER_39_2756 ();
 sg13g2_decap_8 FILLER_39_2781 ();
 sg13g2_decap_8 FILLER_39_2788 ();
 sg13g2_decap_8 FILLER_39_2795 ();
 sg13g2_decap_8 FILLER_39_2802 ();
 sg13g2_decap_8 FILLER_39_2809 ();
 sg13g2_decap_8 FILLER_39_2816 ();
 sg13g2_decap_8 FILLER_39_2823 ();
 sg13g2_decap_8 FILLER_39_2830 ();
 sg13g2_decap_8 FILLER_39_2837 ();
 sg13g2_decap_8 FILLER_39_2844 ();
 sg13g2_fill_2 FILLER_39_2851 ();
 sg13g2_fill_1 FILLER_39_2853 ();
 sg13g2_fill_1 FILLER_39_2859 ();
 sg13g2_decap_8 FILLER_39_2875 ();
 sg13g2_decap_8 FILLER_39_2882 ();
 sg13g2_decap_8 FILLER_39_2889 ();
 sg13g2_fill_2 FILLER_39_2896 ();
 sg13g2_fill_1 FILLER_39_2898 ();
 sg13g2_decap_8 FILLER_39_2935 ();
 sg13g2_fill_1 FILLER_39_2942 ();
 sg13g2_fill_1 FILLER_39_2968 ();
 sg13g2_decap_8 FILLER_39_2977 ();
 sg13g2_decap_8 FILLER_39_2984 ();
 sg13g2_decap_4 FILLER_39_2991 ();
 sg13g2_fill_1 FILLER_39_2995 ();
 sg13g2_fill_2 FILLER_39_3006 ();
 sg13g2_decap_8 FILLER_39_3034 ();
 sg13g2_decap_8 FILLER_39_3041 ();
 sg13g2_decap_8 FILLER_39_3048 ();
 sg13g2_fill_1 FILLER_39_3055 ();
 sg13g2_fill_2 FILLER_39_3089 ();
 sg13g2_fill_1 FILLER_39_3091 ();
 sg13g2_decap_8 FILLER_39_3109 ();
 sg13g2_decap_8 FILLER_39_3133 ();
 sg13g2_decap_8 FILLER_39_3140 ();
 sg13g2_fill_1 FILLER_39_3147 ();
 sg13g2_fill_1 FILLER_39_3174 ();
 sg13g2_decap_8 FILLER_39_3211 ();
 sg13g2_decap_4 FILLER_39_3218 ();
 sg13g2_fill_2 FILLER_39_3222 ();
 sg13g2_decap_8 FILLER_39_3229 ();
 sg13g2_decap_8 FILLER_39_3236 ();
 sg13g2_decap_8 FILLER_39_3243 ();
 sg13g2_decap_8 FILLER_39_3250 ();
 sg13g2_decap_8 FILLER_39_3257 ();
 sg13g2_decap_8 FILLER_39_3264 ();
 sg13g2_decap_8 FILLER_39_3271 ();
 sg13g2_decap_8 FILLER_39_3278 ();
 sg13g2_decap_8 FILLER_39_3285 ();
 sg13g2_decap_4 FILLER_39_3292 ();
 sg13g2_decap_8 FILLER_39_3301 ();
 sg13g2_decap_8 FILLER_39_3308 ();
 sg13g2_decap_8 FILLER_39_3315 ();
 sg13g2_decap_8 FILLER_39_3322 ();
 sg13g2_decap_8 FILLER_39_3329 ();
 sg13g2_fill_1 FILLER_39_3336 ();
 sg13g2_decap_8 FILLER_39_3363 ();
 sg13g2_decap_8 FILLER_39_3370 ();
 sg13g2_decap_8 FILLER_39_3377 ();
 sg13g2_decap_8 FILLER_39_3384 ();
 sg13g2_decap_8 FILLER_39_3391 ();
 sg13g2_decap_8 FILLER_39_3398 ();
 sg13g2_decap_8 FILLER_39_3405 ();
 sg13g2_decap_8 FILLER_39_3412 ();
 sg13g2_decap_8 FILLER_39_3419 ();
 sg13g2_decap_8 FILLER_39_3426 ();
 sg13g2_fill_2 FILLER_39_3433 ();
 sg13g2_fill_1 FILLER_39_3435 ();
 sg13g2_decap_8 FILLER_39_3439 ();
 sg13g2_decap_8 FILLER_39_3446 ();
 sg13g2_decap_8 FILLER_39_3453 ();
 sg13g2_fill_2 FILLER_39_3479 ();
 sg13g2_decap_4 FILLER_39_3490 ();
 sg13g2_fill_1 FILLER_39_3494 ();
 sg13g2_decap_4 FILLER_39_3500 ();
 sg13g2_fill_2 FILLER_39_3504 ();
 sg13g2_decap_8 FILLER_39_3509 ();
 sg13g2_decap_8 FILLER_39_3516 ();
 sg13g2_decap_8 FILLER_39_3523 ();
 sg13g2_fill_2 FILLER_39_3530 ();
 sg13g2_fill_1 FILLER_39_3532 ();
 sg13g2_decap_4 FILLER_39_3543 ();
 sg13g2_decap_8 FILLER_39_3573 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_fill_1 FILLER_40_14 ();
 sg13g2_fill_2 FILLER_40_29 ();
 sg13g2_fill_1 FILLER_40_31 ();
 sg13g2_decap_8 FILLER_40_53 ();
 sg13g2_decap_8 FILLER_40_60 ();
 sg13g2_decap_8 FILLER_40_67 ();
 sg13g2_decap_8 FILLER_40_74 ();
 sg13g2_decap_8 FILLER_40_81 ();
 sg13g2_decap_8 FILLER_40_88 ();
 sg13g2_decap_8 FILLER_40_95 ();
 sg13g2_decap_4 FILLER_40_102 ();
 sg13g2_fill_2 FILLER_40_106 ();
 sg13g2_decap_8 FILLER_40_121 ();
 sg13g2_decap_8 FILLER_40_128 ();
 sg13g2_decap_8 FILLER_40_135 ();
 sg13g2_fill_2 FILLER_40_142 ();
 sg13g2_fill_1 FILLER_40_149 ();
 sg13g2_decap_8 FILLER_40_158 ();
 sg13g2_fill_2 FILLER_40_165 ();
 sg13g2_decap_8 FILLER_40_171 ();
 sg13g2_fill_2 FILLER_40_178 ();
 sg13g2_fill_1 FILLER_40_180 ();
 sg13g2_decap_4 FILLER_40_186 ();
 sg13g2_decap_8 FILLER_40_195 ();
 sg13g2_fill_1 FILLER_40_202 ();
 sg13g2_fill_2 FILLER_40_229 ();
 sg13g2_fill_1 FILLER_40_231 ();
 sg13g2_decap_8 FILLER_40_237 ();
 sg13g2_decap_8 FILLER_40_244 ();
 sg13g2_decap_8 FILLER_40_251 ();
 sg13g2_decap_8 FILLER_40_258 ();
 sg13g2_decap_8 FILLER_40_265 ();
 sg13g2_decap_8 FILLER_40_272 ();
 sg13g2_decap_8 FILLER_40_279 ();
 sg13g2_decap_8 FILLER_40_286 ();
 sg13g2_decap_8 FILLER_40_293 ();
 sg13g2_decap_8 FILLER_40_300 ();
 sg13g2_decap_8 FILLER_40_307 ();
 sg13g2_decap_8 FILLER_40_314 ();
 sg13g2_decap_8 FILLER_40_321 ();
 sg13g2_fill_2 FILLER_40_328 ();
 sg13g2_decap_8 FILLER_40_339 ();
 sg13g2_fill_1 FILLER_40_346 ();
 sg13g2_decap_8 FILLER_40_350 ();
 sg13g2_decap_8 FILLER_40_357 ();
 sg13g2_decap_8 FILLER_40_364 ();
 sg13g2_decap_8 FILLER_40_371 ();
 sg13g2_fill_2 FILLER_40_378 ();
 sg13g2_decap_8 FILLER_40_406 ();
 sg13g2_decap_8 FILLER_40_413 ();
 sg13g2_decap_8 FILLER_40_420 ();
 sg13g2_fill_2 FILLER_40_427 ();
 sg13g2_decap_8 FILLER_40_449 ();
 sg13g2_decap_8 FILLER_40_456 ();
 sg13g2_decap_8 FILLER_40_463 ();
 sg13g2_decap_8 FILLER_40_470 ();
 sg13g2_decap_8 FILLER_40_477 ();
 sg13g2_decap_8 FILLER_40_484 ();
 sg13g2_decap_8 FILLER_40_491 ();
 sg13g2_decap_8 FILLER_40_498 ();
 sg13g2_decap_8 FILLER_40_505 ();
 sg13g2_decap_8 FILLER_40_512 ();
 sg13g2_decap_4 FILLER_40_519 ();
 sg13g2_fill_1 FILLER_40_523 ();
 sg13g2_fill_1 FILLER_40_536 ();
 sg13g2_fill_2 FILLER_40_542 ();
 sg13g2_fill_1 FILLER_40_544 ();
 sg13g2_decap_4 FILLER_40_558 ();
 sg13g2_decap_8 FILLER_40_572 ();
 sg13g2_decap_4 FILLER_40_579 ();
 sg13g2_decap_4 FILLER_40_588 ();
 sg13g2_fill_2 FILLER_40_592 ();
 sg13g2_decap_8 FILLER_40_603 ();
 sg13g2_decap_4 FILLER_40_610 ();
 sg13g2_fill_2 FILLER_40_614 ();
 sg13g2_decap_4 FILLER_40_640 ();
 sg13g2_fill_1 FILLER_40_644 ();
 sg13g2_fill_1 FILLER_40_671 ();
 sg13g2_decap_8 FILLER_40_698 ();
 sg13g2_fill_1 FILLER_40_705 ();
 sg13g2_decap_8 FILLER_40_712 ();
 sg13g2_decap_8 FILLER_40_731 ();
 sg13g2_decap_4 FILLER_40_738 ();
 sg13g2_fill_1 FILLER_40_742 ();
 sg13g2_fill_2 FILLER_40_764 ();
 sg13g2_fill_1 FILLER_40_766 ();
 sg13g2_decap_8 FILLER_40_785 ();
 sg13g2_decap_8 FILLER_40_792 ();
 sg13g2_decap_8 FILLER_40_799 ();
 sg13g2_decap_8 FILLER_40_806 ();
 sg13g2_decap_8 FILLER_40_813 ();
 sg13g2_decap_4 FILLER_40_820 ();
 sg13g2_decap_8 FILLER_40_827 ();
 sg13g2_decap_8 FILLER_40_834 ();
 sg13g2_fill_1 FILLER_40_841 ();
 sg13g2_fill_1 FILLER_40_855 ();
 sg13g2_decap_8 FILLER_40_880 ();
 sg13g2_decap_8 FILLER_40_887 ();
 sg13g2_decap_8 FILLER_40_894 ();
 sg13g2_fill_2 FILLER_40_901 ();
 sg13g2_fill_1 FILLER_40_903 ();
 sg13g2_decap_8 FILLER_40_907 ();
 sg13g2_decap_8 FILLER_40_914 ();
 sg13g2_decap_8 FILLER_40_921 ();
 sg13g2_decap_4 FILLER_40_928 ();
 sg13g2_decap_8 FILLER_40_941 ();
 sg13g2_decap_8 FILLER_40_948 ();
 sg13g2_decap_8 FILLER_40_955 ();
 sg13g2_decap_8 FILLER_40_975 ();
 sg13g2_decap_8 FILLER_40_982 ();
 sg13g2_decap_8 FILLER_40_989 ();
 sg13g2_decap_8 FILLER_40_996 ();
 sg13g2_fill_2 FILLER_40_1003 ();
 sg13g2_fill_1 FILLER_40_1005 ();
 sg13g2_decap_8 FILLER_40_1019 ();
 sg13g2_decap_8 FILLER_40_1026 ();
 sg13g2_decap_8 FILLER_40_1033 ();
 sg13g2_decap_8 FILLER_40_1040 ();
 sg13g2_decap_8 FILLER_40_1047 ();
 sg13g2_fill_2 FILLER_40_1054 ();
 sg13g2_decap_8 FILLER_40_1069 ();
 sg13g2_decap_8 FILLER_40_1076 ();
 sg13g2_decap_8 FILLER_40_1083 ();
 sg13g2_decap_8 FILLER_40_1090 ();
 sg13g2_decap_4 FILLER_40_1097 ();
 sg13g2_decap_8 FILLER_40_1111 ();
 sg13g2_fill_1 FILLER_40_1118 ();
 sg13g2_decap_8 FILLER_40_1125 ();
 sg13g2_decap_8 FILLER_40_1132 ();
 sg13g2_decap_8 FILLER_40_1139 ();
 sg13g2_decap_8 FILLER_40_1146 ();
 sg13g2_decap_8 FILLER_40_1153 ();
 sg13g2_decap_8 FILLER_40_1160 ();
 sg13g2_decap_8 FILLER_40_1167 ();
 sg13g2_decap_8 FILLER_40_1174 ();
 sg13g2_decap_8 FILLER_40_1181 ();
 sg13g2_decap_8 FILLER_40_1188 ();
 sg13g2_decap_4 FILLER_40_1195 ();
 sg13g2_fill_2 FILLER_40_1199 ();
 sg13g2_decap_8 FILLER_40_1204 ();
 sg13g2_decap_8 FILLER_40_1211 ();
 sg13g2_fill_2 FILLER_40_1218 ();
 sg13g2_decap_8 FILLER_40_1246 ();
 sg13g2_decap_8 FILLER_40_1253 ();
 sg13g2_decap_8 FILLER_40_1260 ();
 sg13g2_decap_4 FILLER_40_1293 ();
 sg13g2_fill_1 FILLER_40_1297 ();
 sg13g2_decap_8 FILLER_40_1324 ();
 sg13g2_decap_8 FILLER_40_1331 ();
 sg13g2_decap_8 FILLER_40_1338 ();
 sg13g2_decap_8 FILLER_40_1355 ();
 sg13g2_fill_2 FILLER_40_1362 ();
 sg13g2_decap_8 FILLER_40_1380 ();
 sg13g2_decap_8 FILLER_40_1387 ();
 sg13g2_decap_4 FILLER_40_1394 ();
 sg13g2_decap_8 FILLER_40_1408 ();
 sg13g2_decap_8 FILLER_40_1415 ();
 sg13g2_decap_8 FILLER_40_1422 ();
 sg13g2_decap_8 FILLER_40_1429 ();
 sg13g2_decap_8 FILLER_40_1436 ();
 sg13g2_decap_8 FILLER_40_1443 ();
 sg13g2_decap_8 FILLER_40_1450 ();
 sg13g2_decap_8 FILLER_40_1457 ();
 sg13g2_decap_8 FILLER_40_1464 ();
 sg13g2_decap_8 FILLER_40_1471 ();
 sg13g2_decap_8 FILLER_40_1478 ();
 sg13g2_fill_1 FILLER_40_1495 ();
 sg13g2_fill_1 FILLER_40_1501 ();
 sg13g2_decap_8 FILLER_40_1510 ();
 sg13g2_decap_4 FILLER_40_1517 ();
 sg13g2_fill_1 FILLER_40_1521 ();
 sg13g2_decap_4 FILLER_40_1526 ();
 sg13g2_decap_8 FILLER_40_1542 ();
 sg13g2_decap_8 FILLER_40_1549 ();
 sg13g2_fill_2 FILLER_40_1562 ();
 sg13g2_decap_8 FILLER_40_1570 ();
 sg13g2_fill_2 FILLER_40_1577 ();
 sg13g2_decap_8 FILLER_40_1591 ();
 sg13g2_decap_8 FILLER_40_1598 ();
 sg13g2_decap_4 FILLER_40_1605 ();
 sg13g2_fill_2 FILLER_40_1609 ();
 sg13g2_fill_1 FILLER_40_1625 ();
 sg13g2_decap_8 FILLER_40_1646 ();
 sg13g2_decap_8 FILLER_40_1653 ();
 sg13g2_decap_8 FILLER_40_1660 ();
 sg13g2_decap_4 FILLER_40_1667 ();
 sg13g2_fill_2 FILLER_40_1671 ();
 sg13g2_fill_1 FILLER_40_1705 ();
 sg13g2_decap_8 FILLER_40_1715 ();
 sg13g2_decap_8 FILLER_40_1722 ();
 sg13g2_decap_8 FILLER_40_1729 ();
 sg13g2_decap_8 FILLER_40_1736 ();
 sg13g2_decap_8 FILLER_40_1743 ();
 sg13g2_fill_2 FILLER_40_1750 ();
 sg13g2_fill_1 FILLER_40_1752 ();
 sg13g2_decap_8 FILLER_40_1787 ();
 sg13g2_fill_2 FILLER_40_1794 ();
 sg13g2_fill_1 FILLER_40_1796 ();
 sg13g2_decap_8 FILLER_40_1833 ();
 sg13g2_fill_1 FILLER_40_1840 ();
 sg13g2_decap_8 FILLER_40_1847 ();
 sg13g2_decap_8 FILLER_40_1854 ();
 sg13g2_decap_8 FILLER_40_1861 ();
 sg13g2_fill_1 FILLER_40_1868 ();
 sg13g2_decap_8 FILLER_40_1885 ();
 sg13g2_decap_8 FILLER_40_1892 ();
 sg13g2_decap_8 FILLER_40_1899 ();
 sg13g2_decap_8 FILLER_40_1906 ();
 sg13g2_decap_4 FILLER_40_1913 ();
 sg13g2_fill_2 FILLER_40_1917 ();
 sg13g2_fill_2 FILLER_40_1936 ();
 sg13g2_decap_8 FILLER_40_1987 ();
 sg13g2_fill_2 FILLER_40_1994 ();
 sg13g2_fill_2 FILLER_40_2002 ();
 sg13g2_decap_8 FILLER_40_2036 ();
 sg13g2_decap_8 FILLER_40_2043 ();
 sg13g2_decap_8 FILLER_40_2050 ();
 sg13g2_decap_8 FILLER_40_2057 ();
 sg13g2_decap_8 FILLER_40_2064 ();
 sg13g2_decap_8 FILLER_40_2071 ();
 sg13g2_decap_8 FILLER_40_2078 ();
 sg13g2_decap_8 FILLER_40_2085 ();
 sg13g2_decap_8 FILLER_40_2092 ();
 sg13g2_decap_8 FILLER_40_2099 ();
 sg13g2_decap_8 FILLER_40_2106 ();
 sg13g2_decap_4 FILLER_40_2113 ();
 sg13g2_fill_1 FILLER_40_2117 ();
 sg13g2_fill_2 FILLER_40_2124 ();
 sg13g2_fill_1 FILLER_40_2126 ();
 sg13g2_decap_8 FILLER_40_2154 ();
 sg13g2_decap_4 FILLER_40_2161 ();
 sg13g2_fill_2 FILLER_40_2180 ();
 sg13g2_decap_8 FILLER_40_2206 ();
 sg13g2_decap_8 FILLER_40_2213 ();
 sg13g2_decap_8 FILLER_40_2220 ();
 sg13g2_fill_2 FILLER_40_2227 ();
 sg13g2_fill_1 FILLER_40_2229 ();
 sg13g2_fill_1 FILLER_40_2248 ();
 sg13g2_decap_8 FILLER_40_2258 ();
 sg13g2_fill_2 FILLER_40_2265 ();
 sg13g2_fill_1 FILLER_40_2267 ();
 sg13g2_decap_8 FILLER_40_2301 ();
 sg13g2_decap_8 FILLER_40_2308 ();
 sg13g2_fill_1 FILLER_40_2315 ();
 sg13g2_decap_8 FILLER_40_2322 ();
 sg13g2_decap_4 FILLER_40_2329 ();
 sg13g2_fill_1 FILLER_40_2333 ();
 sg13g2_decap_8 FILLER_40_2367 ();
 sg13g2_decap_8 FILLER_40_2374 ();
 sg13g2_fill_2 FILLER_40_2381 ();
 sg13g2_decap_8 FILLER_40_2386 ();
 sg13g2_fill_1 FILLER_40_2393 ();
 sg13g2_fill_2 FILLER_40_2397 ();
 sg13g2_decap_4 FILLER_40_2414 ();
 sg13g2_fill_1 FILLER_40_2418 ();
 sg13g2_decap_8 FILLER_40_2431 ();
 sg13g2_decap_8 FILLER_40_2438 ();
 sg13g2_fill_2 FILLER_40_2445 ();
 sg13g2_fill_1 FILLER_40_2447 ();
 sg13g2_decap_4 FILLER_40_2454 ();
 sg13g2_decap_8 FILLER_40_2476 ();
 sg13g2_decap_4 FILLER_40_2483 ();
 sg13g2_fill_1 FILLER_40_2487 ();
 sg13g2_fill_2 FILLER_40_2494 ();
 sg13g2_fill_1 FILLER_40_2496 ();
 sg13g2_decap_4 FILLER_40_2514 ();
 sg13g2_fill_2 FILLER_40_2518 ();
 sg13g2_decap_8 FILLER_40_2538 ();
 sg13g2_decap_8 FILLER_40_2545 ();
 sg13g2_fill_2 FILLER_40_2552 ();
 sg13g2_decap_4 FILLER_40_2566 ();
 sg13g2_fill_1 FILLER_40_2570 ();
 sg13g2_decap_8 FILLER_40_2592 ();
 sg13g2_decap_8 FILLER_40_2599 ();
 sg13g2_fill_2 FILLER_40_2606 ();
 sg13g2_decap_4 FILLER_40_2618 ();
 sg13g2_fill_1 FILLER_40_2622 ();
 sg13g2_decap_8 FILLER_40_2629 ();
 sg13g2_decap_8 FILLER_40_2636 ();
 sg13g2_decap_8 FILLER_40_2643 ();
 sg13g2_fill_2 FILLER_40_2650 ();
 sg13g2_decap_8 FILLER_40_2662 ();
 sg13g2_decap_4 FILLER_40_2669 ();
 sg13g2_decap_8 FILLER_40_2676 ();
 sg13g2_decap_8 FILLER_40_2683 ();
 sg13g2_decap_4 FILLER_40_2690 ();
 sg13g2_fill_1 FILLER_40_2694 ();
 sg13g2_fill_2 FILLER_40_2701 ();
 sg13g2_fill_1 FILLER_40_2703 ();
 sg13g2_fill_2 FILLER_40_2731 ();
 sg13g2_fill_1 FILLER_40_2733 ();
 sg13g2_decap_8 FILLER_40_2745 ();
 sg13g2_decap_8 FILLER_40_2752 ();
 sg13g2_fill_2 FILLER_40_2759 ();
 sg13g2_fill_1 FILLER_40_2782 ();
 sg13g2_decap_4 FILLER_40_2808 ();
 sg13g2_fill_2 FILLER_40_2812 ();
 sg13g2_decap_8 FILLER_40_2819 ();
 sg13g2_decap_8 FILLER_40_2826 ();
 sg13g2_fill_2 FILLER_40_2833 ();
 sg13g2_fill_1 FILLER_40_2856 ();
 sg13g2_decap_8 FILLER_40_2883 ();
 sg13g2_decap_8 FILLER_40_2890 ();
 sg13g2_fill_2 FILLER_40_2897 ();
 sg13g2_fill_1 FILLER_40_2899 ();
 sg13g2_decap_8 FILLER_40_2908 ();
 sg13g2_decap_8 FILLER_40_2915 ();
 sg13g2_decap_8 FILLER_40_2922 ();
 sg13g2_fill_1 FILLER_40_2929 ();
 sg13g2_decap_8 FILLER_40_2982 ();
 sg13g2_decap_8 FILLER_40_2989 ();
 sg13g2_decap_8 FILLER_40_2996 ();
 sg13g2_decap_8 FILLER_40_3003 ();
 sg13g2_decap_8 FILLER_40_3010 ();
 sg13g2_decap_8 FILLER_40_3017 ();
 sg13g2_decap_8 FILLER_40_3024 ();
 sg13g2_decap_8 FILLER_40_3048 ();
 sg13g2_decap_8 FILLER_40_3055 ();
 sg13g2_decap_4 FILLER_40_3062 ();
 sg13g2_fill_1 FILLER_40_3066 ();
 sg13g2_decap_8 FILLER_40_3081 ();
 sg13g2_decap_8 FILLER_40_3088 ();
 sg13g2_decap_8 FILLER_40_3095 ();
 sg13g2_fill_2 FILLER_40_3102 ();
 sg13g2_decap_8 FILLER_40_3110 ();
 sg13g2_fill_2 FILLER_40_3117 ();
 sg13g2_decap_8 FILLER_40_3125 ();
 sg13g2_decap_8 FILLER_40_3132 ();
 sg13g2_decap_8 FILLER_40_3139 ();
 sg13g2_decap_8 FILLER_40_3146 ();
 sg13g2_decap_8 FILLER_40_3153 ();
 sg13g2_fill_1 FILLER_40_3160 ();
 sg13g2_decap_8 FILLER_40_3181 ();
 sg13g2_decap_8 FILLER_40_3188 ();
 sg13g2_decap_8 FILLER_40_3195 ();
 sg13g2_decap_8 FILLER_40_3202 ();
 sg13g2_decap_8 FILLER_40_3209 ();
 sg13g2_decap_8 FILLER_40_3216 ();
 sg13g2_decap_8 FILLER_40_3223 ();
 sg13g2_decap_4 FILLER_40_3230 ();
 sg13g2_fill_2 FILLER_40_3234 ();
 sg13g2_decap_8 FILLER_40_3275 ();
 sg13g2_decap_8 FILLER_40_3282 ();
 sg13g2_fill_2 FILLER_40_3289 ();
 sg13g2_decap_8 FILLER_40_3317 ();
 sg13g2_decap_8 FILLER_40_3324 ();
 sg13g2_decap_4 FILLER_40_3331 ();
 sg13g2_fill_2 FILLER_40_3335 ();
 sg13g2_decap_8 FILLER_40_3342 ();
 sg13g2_decap_8 FILLER_40_3349 ();
 sg13g2_decap_8 FILLER_40_3356 ();
 sg13g2_fill_2 FILLER_40_3363 ();
 sg13g2_decap_8 FILLER_40_3399 ();
 sg13g2_decap_8 FILLER_40_3406 ();
 sg13g2_decap_8 FILLER_40_3413 ();
 sg13g2_decap_8 FILLER_40_3420 ();
 sg13g2_decap_8 FILLER_40_3427 ();
 sg13g2_fill_2 FILLER_40_3434 ();
 sg13g2_decap_8 FILLER_40_3444 ();
 sg13g2_decap_8 FILLER_40_3451 ();
 sg13g2_decap_8 FILLER_40_3458 ();
 sg13g2_fill_2 FILLER_40_3465 ();
 sg13g2_fill_2 FILLER_40_3493 ();
 sg13g2_decap_8 FILLER_40_3530 ();
 sg13g2_decap_8 FILLER_40_3551 ();
 sg13g2_fill_1 FILLER_40_3558 ();
 sg13g2_decap_4 FILLER_40_3562 ();
 sg13g2_fill_1 FILLER_40_3566 ();
 sg13g2_decap_4 FILLER_40_3576 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_fill_2 FILLER_41_14 ();
 sg13g2_decap_8 FILLER_41_43 ();
 sg13g2_decap_8 FILLER_41_50 ();
 sg13g2_decap_8 FILLER_41_57 ();
 sg13g2_decap_8 FILLER_41_64 ();
 sg13g2_decap_4 FILLER_41_71 ();
 sg13g2_fill_1 FILLER_41_75 ();
 sg13g2_decap_8 FILLER_41_81 ();
 sg13g2_decap_4 FILLER_41_88 ();
 sg13g2_decap_4 FILLER_41_100 ();
 sg13g2_fill_2 FILLER_41_104 ();
 sg13g2_decap_8 FILLER_41_115 ();
 sg13g2_decap_8 FILLER_41_122 ();
 sg13g2_decap_8 FILLER_41_129 ();
 sg13g2_decap_8 FILLER_41_136 ();
 sg13g2_decap_8 FILLER_41_143 ();
 sg13g2_decap_4 FILLER_41_150 ();
 sg13g2_fill_2 FILLER_41_154 ();
 sg13g2_decap_8 FILLER_41_169 ();
 sg13g2_decap_8 FILLER_41_176 ();
 sg13g2_decap_8 FILLER_41_183 ();
 sg13g2_decap_8 FILLER_41_190 ();
 sg13g2_fill_1 FILLER_41_197 ();
 sg13g2_decap_4 FILLER_41_212 ();
 sg13g2_decap_8 FILLER_41_227 ();
 sg13g2_decap_8 FILLER_41_234 ();
 sg13g2_decap_8 FILLER_41_264 ();
 sg13g2_decap_8 FILLER_41_271 ();
 sg13g2_fill_2 FILLER_41_278 ();
 sg13g2_fill_1 FILLER_41_280 ();
 sg13g2_decap_8 FILLER_41_297 ();
 sg13g2_decap_8 FILLER_41_304 ();
 sg13g2_decap_8 FILLER_41_311 ();
 sg13g2_decap_4 FILLER_41_318 ();
 sg13g2_fill_2 FILLER_41_322 ();
 sg13g2_decap_8 FILLER_41_366 ();
 sg13g2_decap_8 FILLER_41_373 ();
 sg13g2_decap_8 FILLER_41_380 ();
 sg13g2_fill_2 FILLER_41_387 ();
 sg13g2_fill_1 FILLER_41_389 ();
 sg13g2_fill_2 FILLER_41_394 ();
 sg13g2_decap_8 FILLER_41_418 ();
 sg13g2_decap_8 FILLER_41_425 ();
 sg13g2_decap_8 FILLER_41_440 ();
 sg13g2_decap_4 FILLER_41_447 ();
 sg13g2_fill_2 FILLER_41_451 ();
 sg13g2_fill_1 FILLER_41_461 ();
 sg13g2_decap_4 FILLER_41_470 ();
 sg13g2_fill_1 FILLER_41_474 ();
 sg13g2_decap_8 FILLER_41_519 ();
 sg13g2_decap_4 FILLER_41_526 ();
 sg13g2_fill_1 FILLER_41_538 ();
 sg13g2_fill_2 FILLER_41_549 ();
 sg13g2_fill_2 FILLER_41_556 ();
 sg13g2_decap_8 FILLER_41_566 ();
 sg13g2_decap_8 FILLER_41_573 ();
 sg13g2_decap_8 FILLER_41_599 ();
 sg13g2_decap_4 FILLER_41_606 ();
 sg13g2_fill_1 FILLER_41_610 ();
 sg13g2_decap_8 FILLER_41_630 ();
 sg13g2_decap_8 FILLER_41_637 ();
 sg13g2_decap_8 FILLER_41_644 ();
 sg13g2_decap_8 FILLER_41_651 ();
 sg13g2_decap_8 FILLER_41_658 ();
 sg13g2_decap_8 FILLER_41_665 ();
 sg13g2_decap_8 FILLER_41_672 ();
 sg13g2_decap_8 FILLER_41_679 ();
 sg13g2_decap_8 FILLER_41_686 ();
 sg13g2_decap_8 FILLER_41_693 ();
 sg13g2_decap_8 FILLER_41_700 ();
 sg13g2_decap_8 FILLER_41_707 ();
 sg13g2_decap_4 FILLER_41_714 ();
 sg13g2_fill_2 FILLER_41_718 ();
 sg13g2_decap_4 FILLER_41_724 ();
 sg13g2_decap_8 FILLER_41_770 ();
 sg13g2_decap_8 FILLER_41_790 ();
 sg13g2_decap_8 FILLER_41_797 ();
 sg13g2_fill_2 FILLER_41_804 ();
 sg13g2_fill_2 FILLER_41_833 ();
 sg13g2_fill_2 FILLER_41_846 ();
 sg13g2_decap_4 FILLER_41_870 ();
 sg13g2_fill_2 FILLER_41_874 ();
 sg13g2_decap_8 FILLER_41_961 ();
 sg13g2_decap_8 FILLER_41_968 ();
 sg13g2_decap_8 FILLER_41_975 ();
 sg13g2_decap_8 FILLER_41_982 ();
 sg13g2_decap_4 FILLER_41_989 ();
 sg13g2_fill_2 FILLER_41_993 ();
 sg13g2_decap_4 FILLER_41_999 ();
 sg13g2_decap_8 FILLER_41_1006 ();
 sg13g2_decap_8 FILLER_41_1026 ();
 sg13g2_decap_4 FILLER_41_1033 ();
 sg13g2_fill_2 FILLER_41_1037 ();
 sg13g2_decap_8 FILLER_41_1056 ();
 sg13g2_decap_8 FILLER_41_1063 ();
 sg13g2_decap_8 FILLER_41_1070 ();
 sg13g2_decap_8 FILLER_41_1077 ();
 sg13g2_decap_8 FILLER_41_1084 ();
 sg13g2_fill_2 FILLER_41_1091 ();
 sg13g2_fill_2 FILLER_41_1101 ();
 sg13g2_decap_8 FILLER_41_1116 ();
 sg13g2_decap_8 FILLER_41_1123 ();
 sg13g2_decap_8 FILLER_41_1130 ();
 sg13g2_decap_4 FILLER_41_1137 ();
 sg13g2_decap_8 FILLER_41_1182 ();
 sg13g2_decap_8 FILLER_41_1189 ();
 sg13g2_decap_4 FILLER_41_1196 ();
 sg13g2_decap_8 FILLER_41_1210 ();
 sg13g2_decap_8 FILLER_41_1217 ();
 sg13g2_decap_8 FILLER_41_1224 ();
 sg13g2_decap_8 FILLER_41_1267 ();
 sg13g2_decap_8 FILLER_41_1274 ();
 sg13g2_decap_8 FILLER_41_1281 ();
 sg13g2_decap_4 FILLER_41_1288 ();
 sg13g2_fill_1 FILLER_41_1292 ();
 sg13g2_decap_4 FILLER_41_1301 ();
 sg13g2_fill_1 FILLER_41_1305 ();
 sg13g2_decap_8 FILLER_41_1316 ();
 sg13g2_decap_8 FILLER_41_1323 ();
 sg13g2_decap_8 FILLER_41_1330 ();
 sg13g2_decap_8 FILLER_41_1337 ();
 sg13g2_decap_8 FILLER_41_1344 ();
 sg13g2_decap_8 FILLER_41_1351 ();
 sg13g2_decap_8 FILLER_41_1358 ();
 sg13g2_decap_8 FILLER_41_1365 ();
 sg13g2_decap_8 FILLER_41_1372 ();
 sg13g2_decap_8 FILLER_41_1379 ();
 sg13g2_fill_1 FILLER_41_1386 ();
 sg13g2_decap_8 FILLER_41_1397 ();
 sg13g2_decap_4 FILLER_41_1404 ();
 sg13g2_fill_1 FILLER_41_1408 ();
 sg13g2_fill_1 FILLER_41_1415 ();
 sg13g2_decap_8 FILLER_41_1422 ();
 sg13g2_decap_8 FILLER_41_1429 ();
 sg13g2_decap_4 FILLER_41_1436 ();
 sg13g2_fill_2 FILLER_41_1440 ();
 sg13g2_decap_8 FILLER_41_1447 ();
 sg13g2_decap_8 FILLER_41_1454 ();
 sg13g2_decap_8 FILLER_41_1461 ();
 sg13g2_decap_8 FILLER_41_1468 ();
 sg13g2_decap_4 FILLER_41_1475 ();
 sg13g2_fill_1 FILLER_41_1520 ();
 sg13g2_fill_2 FILLER_41_1529 ();
 sg13g2_fill_1 FILLER_41_1531 ();
 sg13g2_fill_2 FILLER_41_1540 ();
 sg13g2_decap_8 FILLER_41_1552 ();
 sg13g2_decap_8 FILLER_41_1559 ();
 sg13g2_decap_8 FILLER_41_1566 ();
 sg13g2_decap_8 FILLER_41_1573 ();
 sg13g2_decap_8 FILLER_41_1580 ();
 sg13g2_decap_8 FILLER_41_1587 ();
 sg13g2_decap_8 FILLER_41_1594 ();
 sg13g2_decap_8 FILLER_41_1601 ();
 sg13g2_decap_8 FILLER_41_1608 ();
 sg13g2_fill_2 FILLER_41_1615 ();
 sg13g2_decap_8 FILLER_41_1622 ();
 sg13g2_fill_1 FILLER_41_1629 ();
 sg13g2_decap_8 FILLER_41_1635 ();
 sg13g2_decap_8 FILLER_41_1642 ();
 sg13g2_decap_8 FILLER_41_1649 ();
 sg13g2_decap_8 FILLER_41_1656 ();
 sg13g2_decap_4 FILLER_41_1663 ();
 sg13g2_fill_2 FILLER_41_1667 ();
 sg13g2_fill_1 FILLER_41_1675 ();
 sg13g2_decap_4 FILLER_41_1684 ();
 sg13g2_fill_1 FILLER_41_1701 ();
 sg13g2_fill_2 FILLER_41_1722 ();
 sg13g2_fill_1 FILLER_41_1724 ();
 sg13g2_decap_8 FILLER_41_1733 ();
 sg13g2_fill_1 FILLER_41_1740 ();
 sg13g2_decap_8 FILLER_41_1752 ();
 sg13g2_fill_1 FILLER_41_1759 ();
 sg13g2_decap_8 FILLER_41_1772 ();
 sg13g2_decap_8 FILLER_41_1779 ();
 sg13g2_decap_8 FILLER_41_1786 ();
 sg13g2_decap_8 FILLER_41_1793 ();
 sg13g2_fill_1 FILLER_41_1800 ();
 sg13g2_decap_8 FILLER_41_1811 ();
 sg13g2_decap_8 FILLER_41_1818 ();
 sg13g2_decap_8 FILLER_41_1825 ();
 sg13g2_decap_8 FILLER_41_1832 ();
 sg13g2_decap_8 FILLER_41_1839 ();
 sg13g2_decap_8 FILLER_41_1846 ();
 sg13g2_decap_8 FILLER_41_1863 ();
 sg13g2_decap_8 FILLER_41_1870 ();
 sg13g2_decap_8 FILLER_41_1877 ();
 sg13g2_decap_8 FILLER_41_1884 ();
 sg13g2_decap_8 FILLER_41_1891 ();
 sg13g2_decap_8 FILLER_41_1898 ();
 sg13g2_decap_4 FILLER_41_1905 ();
 sg13g2_fill_2 FILLER_41_1909 ();
 sg13g2_decap_4 FILLER_41_1921 ();
 sg13g2_decap_8 FILLER_41_1931 ();
 sg13g2_decap_8 FILLER_41_1938 ();
 sg13g2_decap_8 FILLER_41_1945 ();
 sg13g2_decap_8 FILLER_41_1952 ();
 sg13g2_decap_4 FILLER_41_1959 ();
 sg13g2_fill_2 FILLER_41_1963 ();
 sg13g2_decap_8 FILLER_41_1971 ();
 sg13g2_decap_8 FILLER_41_1978 ();
 sg13g2_decap_8 FILLER_41_1985 ();
 sg13g2_decap_8 FILLER_41_1992 ();
 sg13g2_decap_8 FILLER_41_1999 ();
 sg13g2_decap_8 FILLER_41_2041 ();
 sg13g2_decap_8 FILLER_41_2048 ();
 sg13g2_decap_8 FILLER_41_2055 ();
 sg13g2_decap_4 FILLER_41_2062 ();
 sg13g2_fill_1 FILLER_41_2066 ();
 sg13g2_decap_4 FILLER_41_2079 ();
 sg13g2_fill_1 FILLER_41_2083 ();
 sg13g2_decap_8 FILLER_41_2097 ();
 sg13g2_fill_2 FILLER_41_2104 ();
 sg13g2_fill_1 FILLER_41_2106 ();
 sg13g2_decap_4 FILLER_41_2122 ();
 sg13g2_fill_2 FILLER_41_2136 ();
 sg13g2_fill_1 FILLER_41_2138 ();
 sg13g2_decap_4 FILLER_41_2142 ();
 sg13g2_fill_1 FILLER_41_2146 ();
 sg13g2_fill_2 FILLER_41_2197 ();
 sg13g2_decap_8 FILLER_41_2216 ();
 sg13g2_fill_2 FILLER_41_2223 ();
 sg13g2_fill_2 FILLER_41_2240 ();
 sg13g2_decap_8 FILLER_41_2254 ();
 sg13g2_decap_8 FILLER_41_2261 ();
 sg13g2_decap_8 FILLER_41_2268 ();
 sg13g2_decap_4 FILLER_41_2275 ();
 sg13g2_decap_8 FILLER_41_2297 ();
 sg13g2_decap_8 FILLER_41_2304 ();
 sg13g2_decap_8 FILLER_41_2311 ();
 sg13g2_decap_8 FILLER_41_2318 ();
 sg13g2_decap_8 FILLER_41_2325 ();
 sg13g2_fill_1 FILLER_41_2332 ();
 sg13g2_fill_1 FILLER_41_2338 ();
 sg13g2_decap_8 FILLER_41_2361 ();
 sg13g2_fill_1 FILLER_41_2382 ();
 sg13g2_fill_2 FILLER_41_2392 ();
 sg13g2_decap_8 FILLER_41_2418 ();
 sg13g2_decap_4 FILLER_41_2425 ();
 sg13g2_decap_8 FILLER_41_2447 ();
 sg13g2_decap_8 FILLER_41_2454 ();
 sg13g2_fill_2 FILLER_41_2461 ();
 sg13g2_fill_1 FILLER_41_2463 ();
 sg13g2_decap_8 FILLER_41_2470 ();
 sg13g2_decap_4 FILLER_41_2477 ();
 sg13g2_fill_1 FILLER_41_2481 ();
 sg13g2_decap_8 FILLER_41_2496 ();
 sg13g2_decap_8 FILLER_41_2503 ();
 sg13g2_decap_8 FILLER_41_2510 ();
 sg13g2_decap_4 FILLER_41_2517 ();
 sg13g2_decap_8 FILLER_41_2540 ();
 sg13g2_decap_8 FILLER_41_2547 ();
 sg13g2_decap_8 FILLER_41_2554 ();
 sg13g2_decap_8 FILLER_41_2561 ();
 sg13g2_fill_1 FILLER_41_2574 ();
 sg13g2_decap_8 FILLER_41_2585 ();
 sg13g2_decap_8 FILLER_41_2597 ();
 sg13g2_decap_4 FILLER_41_2604 ();
 sg13g2_fill_1 FILLER_41_2608 ();
 sg13g2_decap_8 FILLER_41_2635 ();
 sg13g2_decap_4 FILLER_41_2642 ();
 sg13g2_fill_1 FILLER_41_2646 ();
 sg13g2_decap_8 FILLER_41_2658 ();
 sg13g2_decap_8 FILLER_41_2665 ();
 sg13g2_fill_1 FILLER_41_2672 ();
 sg13g2_decap_8 FILLER_41_2679 ();
 sg13g2_decap_8 FILLER_41_2686 ();
 sg13g2_decap_8 FILLER_41_2693 ();
 sg13g2_decap_8 FILLER_41_2700 ();
 sg13g2_decap_8 FILLER_41_2707 ();
 sg13g2_fill_2 FILLER_41_2714 ();
 sg13g2_fill_1 FILLER_41_2716 ();
 sg13g2_decap_8 FILLER_41_2723 ();
 sg13g2_decap_8 FILLER_41_2730 ();
 sg13g2_decap_8 FILLER_41_2737 ();
 sg13g2_decap_4 FILLER_41_2744 ();
 sg13g2_decap_8 FILLER_41_2754 ();
 sg13g2_decap_8 FILLER_41_2761 ();
 sg13g2_decap_8 FILLER_41_2768 ();
 sg13g2_fill_2 FILLER_41_2809 ();
 sg13g2_fill_1 FILLER_41_2811 ();
 sg13g2_decap_8 FILLER_41_2832 ();
 sg13g2_decap_8 FILLER_41_2839 ();
 sg13g2_fill_1 FILLER_41_2846 ();
 sg13g2_fill_2 FILLER_41_2867 ();
 sg13g2_decap_8 FILLER_41_2892 ();
 sg13g2_decap_8 FILLER_41_2899 ();
 sg13g2_fill_2 FILLER_41_2906 ();
 sg13g2_decap_8 FILLER_41_2914 ();
 sg13g2_decap_8 FILLER_41_2921 ();
 sg13g2_fill_2 FILLER_41_2928 ();
 sg13g2_decap_8 FILLER_41_2938 ();
 sg13g2_decap_8 FILLER_41_2945 ();
 sg13g2_decap_8 FILLER_41_2961 ();
 sg13g2_decap_4 FILLER_41_2968 ();
 sg13g2_fill_1 FILLER_41_2972 ();
 sg13g2_decap_8 FILLER_41_2979 ();
 sg13g2_decap_8 FILLER_41_2986 ();
 sg13g2_decap_8 FILLER_41_2993 ();
 sg13g2_decap_8 FILLER_41_3000 ();
 sg13g2_decap_8 FILLER_41_3007 ();
 sg13g2_decap_8 FILLER_41_3014 ();
 sg13g2_decap_8 FILLER_41_3021 ();
 sg13g2_decap_8 FILLER_41_3028 ();
 sg13g2_decap_4 FILLER_41_3035 ();
 sg13g2_fill_2 FILLER_41_3045 ();
 sg13g2_fill_1 FILLER_41_3047 ();
 sg13g2_decap_8 FILLER_41_3051 ();
 sg13g2_decap_8 FILLER_41_3058 ();
 sg13g2_decap_4 FILLER_41_3065 ();
 sg13g2_fill_1 FILLER_41_3069 ();
 sg13g2_decap_8 FILLER_41_3079 ();
 sg13g2_decap_8 FILLER_41_3086 ();
 sg13g2_decap_8 FILLER_41_3093 ();
 sg13g2_decap_8 FILLER_41_3100 ();
 sg13g2_decap_8 FILLER_41_3107 ();
 sg13g2_decap_8 FILLER_41_3114 ();
 sg13g2_decap_8 FILLER_41_3121 ();
 sg13g2_decap_8 FILLER_41_3128 ();
 sg13g2_decap_8 FILLER_41_3135 ();
 sg13g2_decap_8 FILLER_41_3142 ();
 sg13g2_decap_8 FILLER_41_3149 ();
 sg13g2_decap_8 FILLER_41_3156 ();
 sg13g2_decap_8 FILLER_41_3163 ();
 sg13g2_decap_8 FILLER_41_3170 ();
 sg13g2_decap_8 FILLER_41_3177 ();
 sg13g2_decap_8 FILLER_41_3184 ();
 sg13g2_decap_8 FILLER_41_3191 ();
 sg13g2_fill_2 FILLER_41_3198 ();
 sg13g2_decap_8 FILLER_41_3205 ();
 sg13g2_decap_8 FILLER_41_3215 ();
 sg13g2_decap_4 FILLER_41_3222 ();
 sg13g2_decap_8 FILLER_41_3231 ();
 sg13g2_decap_8 FILLER_41_3238 ();
 sg13g2_decap_4 FILLER_41_3245 ();
 sg13g2_decap_8 FILLER_41_3259 ();
 sg13g2_fill_2 FILLER_41_3266 ();
 sg13g2_fill_1 FILLER_41_3268 ();
 sg13g2_decap_8 FILLER_41_3305 ();
 sg13g2_decap_8 FILLER_41_3312 ();
 sg13g2_decap_8 FILLER_41_3319 ();
 sg13g2_decap_8 FILLER_41_3326 ();
 sg13g2_decap_8 FILLER_41_3333 ();
 sg13g2_decap_8 FILLER_41_3340 ();
 sg13g2_decap_8 FILLER_41_3347 ();
 sg13g2_decap_8 FILLER_41_3354 ();
 sg13g2_fill_2 FILLER_41_3361 ();
 sg13g2_decap_8 FILLER_41_3373 ();
 sg13g2_decap_8 FILLER_41_3380 ();
 sg13g2_decap_8 FILLER_41_3387 ();
 sg13g2_decap_8 FILLER_41_3394 ();
 sg13g2_fill_1 FILLER_41_3401 ();
 sg13g2_decap_8 FILLER_41_3428 ();
 sg13g2_decap_8 FILLER_41_3435 ();
 sg13g2_decap_8 FILLER_41_3442 ();
 sg13g2_decap_8 FILLER_41_3449 ();
 sg13g2_decap_8 FILLER_41_3456 ();
 sg13g2_decap_4 FILLER_41_3463 ();
 sg13g2_fill_2 FILLER_41_3467 ();
 sg13g2_decap_8 FILLER_41_3477 ();
 sg13g2_decap_8 FILLER_41_3484 ();
 sg13g2_decap_8 FILLER_41_3491 ();
 sg13g2_fill_2 FILLER_41_3498 ();
 sg13g2_decap_8 FILLER_41_3536 ();
 sg13g2_fill_2 FILLER_41_3543 ();
 sg13g2_decap_8 FILLER_41_3563 ();
 sg13g2_decap_8 FILLER_41_3570 ();
 sg13g2_fill_2 FILLER_41_3577 ();
 sg13g2_fill_1 FILLER_41_3579 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_decap_8 FILLER_42_14 ();
 sg13g2_decap_4 FILLER_42_21 ();
 sg13g2_decap_8 FILLER_42_39 ();
 sg13g2_decap_8 FILLER_42_46 ();
 sg13g2_decap_8 FILLER_42_53 ();
 sg13g2_decap_8 FILLER_42_60 ();
 sg13g2_decap_8 FILLER_42_67 ();
 sg13g2_decap_8 FILLER_42_74 ();
 sg13g2_decap_4 FILLER_42_81 ();
 sg13g2_fill_2 FILLER_42_85 ();
 sg13g2_fill_1 FILLER_42_94 ();
 sg13g2_decap_8 FILLER_42_123 ();
 sg13g2_decap_8 FILLER_42_130 ();
 sg13g2_decap_8 FILLER_42_137 ();
 sg13g2_fill_2 FILLER_42_144 ();
 sg13g2_fill_1 FILLER_42_146 ();
 sg13g2_decap_8 FILLER_42_169 ();
 sg13g2_fill_2 FILLER_42_176 ();
 sg13g2_decap_4 FILLER_42_185 ();
 sg13g2_fill_2 FILLER_42_189 ();
 sg13g2_decap_8 FILLER_42_230 ();
 sg13g2_decap_4 FILLER_42_237 ();
 sg13g2_fill_1 FILLER_42_241 ();
 sg13g2_decap_8 FILLER_42_294 ();
 sg13g2_decap_8 FILLER_42_301 ();
 sg13g2_fill_2 FILLER_42_308 ();
 sg13g2_fill_1 FILLER_42_310 ();
 sg13g2_fill_1 FILLER_42_337 ();
 sg13g2_decap_8 FILLER_42_366 ();
 sg13g2_decap_8 FILLER_42_373 ();
 sg13g2_decap_8 FILLER_42_380 ();
 sg13g2_decap_8 FILLER_42_391 ();
 sg13g2_decap_8 FILLER_42_398 ();
 sg13g2_decap_8 FILLER_42_405 ();
 sg13g2_decap_8 FILLER_42_412 ();
 sg13g2_decap_8 FILLER_42_419 ();
 sg13g2_decap_4 FILLER_42_426 ();
 sg13g2_fill_1 FILLER_42_430 ();
 sg13g2_decap_4 FILLER_42_435 ();
 sg13g2_fill_1 FILLER_42_439 ();
 sg13g2_decap_8 FILLER_42_446 ();
 sg13g2_decap_8 FILLER_42_453 ();
 sg13g2_decap_8 FILLER_42_468 ();
 sg13g2_decap_8 FILLER_42_475 ();
 sg13g2_decap_8 FILLER_42_482 ();
 sg13g2_decap_8 FILLER_42_489 ();
 sg13g2_decap_4 FILLER_42_496 ();
 sg13g2_fill_2 FILLER_42_500 ();
 sg13g2_decap_8 FILLER_42_516 ();
 sg13g2_decap_8 FILLER_42_523 ();
 sg13g2_decap_8 FILLER_42_530 ();
 sg13g2_decap_8 FILLER_42_537 ();
 sg13g2_decap_8 FILLER_42_544 ();
 sg13g2_decap_8 FILLER_42_551 ();
 sg13g2_fill_2 FILLER_42_558 ();
 sg13g2_decap_8 FILLER_42_563 ();
 sg13g2_decap_4 FILLER_42_570 ();
 sg13g2_decap_8 FILLER_42_600 ();
 sg13g2_decap_8 FILLER_42_607 ();
 sg13g2_fill_1 FILLER_42_614 ();
 sg13g2_decap_8 FILLER_42_624 ();
 sg13g2_decap_8 FILLER_42_631 ();
 sg13g2_decap_8 FILLER_42_638 ();
 sg13g2_decap_8 FILLER_42_645 ();
 sg13g2_decap_8 FILLER_42_652 ();
 sg13g2_decap_8 FILLER_42_659 ();
 sg13g2_decap_8 FILLER_42_666 ();
 sg13g2_decap_8 FILLER_42_673 ();
 sg13g2_decap_4 FILLER_42_680 ();
 sg13g2_fill_2 FILLER_42_684 ();
 sg13g2_decap_8 FILLER_42_691 ();
 sg13g2_decap_8 FILLER_42_698 ();
 sg13g2_decap_8 FILLER_42_705 ();
 sg13g2_fill_1 FILLER_42_712 ();
 sg13g2_fill_2 FILLER_42_721 ();
 sg13g2_decap_8 FILLER_42_730 ();
 sg13g2_decap_8 FILLER_42_737 ();
 sg13g2_fill_2 FILLER_42_744 ();
 sg13g2_fill_1 FILLER_42_746 ();
 sg13g2_fill_2 FILLER_42_757 ();
 sg13g2_decap_8 FILLER_42_763 ();
 sg13g2_decap_8 FILLER_42_770 ();
 sg13g2_decap_8 FILLER_42_777 ();
 sg13g2_decap_8 FILLER_42_784 ();
 sg13g2_decap_8 FILLER_42_791 ();
 sg13g2_decap_4 FILLER_42_798 ();
 sg13g2_fill_2 FILLER_42_805 ();
 sg13g2_fill_1 FILLER_42_807 ();
 sg13g2_fill_2 FILLER_42_841 ();
 sg13g2_fill_1 FILLER_42_857 ();
 sg13g2_decap_8 FILLER_42_883 ();
 sg13g2_decap_8 FILLER_42_890 ();
 sg13g2_decap_4 FILLER_42_897 ();
 sg13g2_fill_1 FILLER_42_901 ();
 sg13g2_decap_8 FILLER_42_928 ();
 sg13g2_decap_8 FILLER_42_935 ();
 sg13g2_decap_8 FILLER_42_942 ();
 sg13g2_decap_4 FILLER_42_949 ();
 sg13g2_decap_8 FILLER_42_957 ();
 sg13g2_decap_8 FILLER_42_964 ();
 sg13g2_decap_8 FILLER_42_971 ();
 sg13g2_decap_8 FILLER_42_978 ();
 sg13g2_fill_2 FILLER_42_985 ();
 sg13g2_fill_1 FILLER_42_987 ();
 sg13g2_decap_4 FILLER_42_1005 ();
 sg13g2_fill_1 FILLER_42_1009 ();
 sg13g2_decap_8 FILLER_42_1019 ();
 sg13g2_decap_8 FILLER_42_1026 ();
 sg13g2_decap_8 FILLER_42_1033 ();
 sg13g2_decap_8 FILLER_42_1040 ();
 sg13g2_decap_8 FILLER_42_1047 ();
 sg13g2_decap_8 FILLER_42_1054 ();
 sg13g2_decap_8 FILLER_42_1061 ();
 sg13g2_fill_2 FILLER_42_1068 ();
 sg13g2_decap_8 FILLER_42_1078 ();
 sg13g2_fill_2 FILLER_42_1085 ();
 sg13g2_fill_1 FILLER_42_1087 ();
 sg13g2_decap_8 FILLER_42_1110 ();
 sg13g2_fill_2 FILLER_42_1117 ();
 sg13g2_decap_8 FILLER_42_1129 ();
 sg13g2_decap_8 FILLER_42_1136 ();
 sg13g2_decap_8 FILLER_42_1143 ();
 sg13g2_decap_8 FILLER_42_1150 ();
 sg13g2_decap_8 FILLER_42_1157 ();
 sg13g2_decap_4 FILLER_42_1164 ();
 sg13g2_decap_8 FILLER_42_1224 ();
 sg13g2_decap_8 FILLER_42_1231 ();
 sg13g2_decap_8 FILLER_42_1238 ();
 sg13g2_decap_8 FILLER_42_1245 ();
 sg13g2_decap_8 FILLER_42_1252 ();
 sg13g2_fill_2 FILLER_42_1259 ();
 sg13g2_decap_8 FILLER_42_1266 ();
 sg13g2_decap_8 FILLER_42_1273 ();
 sg13g2_decap_8 FILLER_42_1280 ();
 sg13g2_decap_8 FILLER_42_1287 ();
 sg13g2_decap_8 FILLER_42_1294 ();
 sg13g2_decap_8 FILLER_42_1301 ();
 sg13g2_decap_8 FILLER_42_1308 ();
 sg13g2_decap_8 FILLER_42_1315 ();
 sg13g2_decap_8 FILLER_42_1322 ();
 sg13g2_decap_8 FILLER_42_1329 ();
 sg13g2_decap_4 FILLER_42_1336 ();
 sg13g2_fill_1 FILLER_42_1340 ();
 sg13g2_decap_8 FILLER_42_1377 ();
 sg13g2_fill_2 FILLER_42_1384 ();
 sg13g2_fill_1 FILLER_42_1386 ();
 sg13g2_decap_8 FILLER_42_1413 ();
 sg13g2_fill_1 FILLER_42_1420 ();
 sg13g2_decap_4 FILLER_42_1431 ();
 sg13g2_decap_8 FILLER_42_1441 ();
 sg13g2_decap_8 FILLER_42_1448 ();
 sg13g2_decap_8 FILLER_42_1455 ();
 sg13g2_decap_4 FILLER_42_1462 ();
 sg13g2_fill_1 FILLER_42_1500 ();
 sg13g2_decap_8 FILLER_42_1506 ();
 sg13g2_decap_8 FILLER_42_1513 ();
 sg13g2_decap_8 FILLER_42_1520 ();
 sg13g2_decap_8 FILLER_42_1527 ();
 sg13g2_decap_8 FILLER_42_1534 ();
 sg13g2_fill_1 FILLER_42_1541 ();
 sg13g2_decap_8 FILLER_42_1574 ();
 sg13g2_decap_8 FILLER_42_1581 ();
 sg13g2_decap_8 FILLER_42_1588 ();
 sg13g2_decap_8 FILLER_42_1595 ();
 sg13g2_decap_8 FILLER_42_1602 ();
 sg13g2_decap_8 FILLER_42_1609 ();
 sg13g2_decap_8 FILLER_42_1616 ();
 sg13g2_decap_8 FILLER_42_1623 ();
 sg13g2_decap_8 FILLER_42_1630 ();
 sg13g2_decap_8 FILLER_42_1637 ();
 sg13g2_decap_8 FILLER_42_1644 ();
 sg13g2_decap_8 FILLER_42_1651 ();
 sg13g2_decap_8 FILLER_42_1658 ();
 sg13g2_decap_8 FILLER_42_1665 ();
 sg13g2_decap_8 FILLER_42_1672 ();
 sg13g2_decap_8 FILLER_42_1679 ();
 sg13g2_decap_8 FILLER_42_1686 ();
 sg13g2_decap_8 FILLER_42_1693 ();
 sg13g2_decap_8 FILLER_42_1700 ();
 sg13g2_decap_8 FILLER_42_1707 ();
 sg13g2_fill_2 FILLER_42_1714 ();
 sg13g2_fill_1 FILLER_42_1716 ();
 sg13g2_decap_4 FILLER_42_1727 ();
 sg13g2_fill_1 FILLER_42_1731 ();
 sg13g2_decap_8 FILLER_42_1738 ();
 sg13g2_fill_1 FILLER_42_1745 ();
 sg13g2_decap_8 FILLER_42_1754 ();
 sg13g2_decap_8 FILLER_42_1761 ();
 sg13g2_decap_8 FILLER_42_1768 ();
 sg13g2_decap_8 FILLER_42_1775 ();
 sg13g2_decap_8 FILLER_42_1782 ();
 sg13g2_decap_8 FILLER_42_1789 ();
 sg13g2_decap_8 FILLER_42_1796 ();
 sg13g2_decap_8 FILLER_42_1803 ();
 sg13g2_decap_8 FILLER_42_1820 ();
 sg13g2_decap_8 FILLER_42_1827 ();
 sg13g2_decap_8 FILLER_42_1834 ();
 sg13g2_decap_8 FILLER_42_1841 ();
 sg13g2_decap_8 FILLER_42_1848 ();
 sg13g2_decap_8 FILLER_42_1855 ();
 sg13g2_decap_8 FILLER_42_1888 ();
 sg13g2_decap_8 FILLER_42_1895 ();
 sg13g2_decap_4 FILLER_42_1902 ();
 sg13g2_fill_1 FILLER_42_1906 ();
 sg13g2_decap_8 FILLER_42_1933 ();
 sg13g2_decap_8 FILLER_42_1940 ();
 sg13g2_decap_8 FILLER_42_1947 ();
 sg13g2_decap_8 FILLER_42_1954 ();
 sg13g2_decap_8 FILLER_42_1961 ();
 sg13g2_decap_8 FILLER_42_1968 ();
 sg13g2_decap_8 FILLER_42_1975 ();
 sg13g2_decap_8 FILLER_42_1982 ();
 sg13g2_decap_8 FILLER_42_1989 ();
 sg13g2_decap_4 FILLER_42_2022 ();
 sg13g2_fill_2 FILLER_42_2029 ();
 sg13g2_decap_8 FILLER_42_2043 ();
 sg13g2_decap_8 FILLER_42_2050 ();
 sg13g2_decap_8 FILLER_42_2057 ();
 sg13g2_decap_8 FILLER_42_2064 ();
 sg13g2_fill_1 FILLER_42_2071 ();
 sg13g2_fill_2 FILLER_42_2087 ();
 sg13g2_decap_8 FILLER_42_2101 ();
 sg13g2_fill_2 FILLER_42_2108 ();
 sg13g2_decap_8 FILLER_42_2113 ();
 sg13g2_decap_8 FILLER_42_2120 ();
 sg13g2_decap_8 FILLER_42_2127 ();
 sg13g2_decap_8 FILLER_42_2134 ();
 sg13g2_decap_8 FILLER_42_2141 ();
 sg13g2_decap_8 FILLER_42_2148 ();
 sg13g2_decap_4 FILLER_42_2155 ();
 sg13g2_fill_1 FILLER_42_2159 ();
 sg13g2_fill_1 FILLER_42_2193 ();
 sg13g2_fill_2 FILLER_42_2209 ();
 sg13g2_fill_1 FILLER_42_2211 ();
 sg13g2_decap_8 FILLER_42_2220 ();
 sg13g2_decap_8 FILLER_42_2227 ();
 sg13g2_decap_4 FILLER_42_2234 ();
 sg13g2_fill_1 FILLER_42_2238 ();
 sg13g2_decap_8 FILLER_42_2253 ();
 sg13g2_decap_8 FILLER_42_2260 ();
 sg13g2_fill_2 FILLER_42_2267 ();
 sg13g2_decap_4 FILLER_42_2273 ();
 sg13g2_fill_1 FILLER_42_2292 ();
 sg13g2_decap_8 FILLER_42_2299 ();
 sg13g2_fill_2 FILLER_42_2306 ();
 sg13g2_fill_2 FILLER_42_2316 ();
 sg13g2_fill_1 FILLER_42_2318 ();
 sg13g2_decap_8 FILLER_42_2327 ();
 sg13g2_decap_8 FILLER_42_2334 ();
 sg13g2_fill_1 FILLER_42_2341 ();
 sg13g2_decap_4 FILLER_42_2347 ();
 sg13g2_fill_1 FILLER_42_2351 ();
 sg13g2_fill_2 FILLER_42_2360 ();
 sg13g2_decap_8 FILLER_42_2365 ();
 sg13g2_decap_8 FILLER_42_2380 ();
 sg13g2_decap_8 FILLER_42_2387 ();
 sg13g2_decap_8 FILLER_42_2397 ();
 sg13g2_decap_8 FILLER_42_2404 ();
 sg13g2_decap_8 FILLER_42_2411 ();
 sg13g2_decap_8 FILLER_42_2418 ();
 sg13g2_fill_2 FILLER_42_2425 ();
 sg13g2_decap_8 FILLER_42_2452 ();
 sg13g2_decap_4 FILLER_42_2459 ();
 sg13g2_decap_8 FILLER_42_2478 ();
 sg13g2_decap_8 FILLER_42_2485 ();
 sg13g2_decap_8 FILLER_42_2492 ();
 sg13g2_decap_8 FILLER_42_2499 ();
 sg13g2_decap_8 FILLER_42_2506 ();
 sg13g2_decap_8 FILLER_42_2513 ();
 sg13g2_decap_4 FILLER_42_2520 ();
 sg13g2_fill_2 FILLER_42_2524 ();
 sg13g2_decap_8 FILLER_42_2537 ();
 sg13g2_fill_1 FILLER_42_2544 ();
 sg13g2_decap_8 FILLER_42_2555 ();
 sg13g2_decap_8 FILLER_42_2562 ();
 sg13g2_fill_2 FILLER_42_2569 ();
 sg13g2_decap_8 FILLER_42_2579 ();
 sg13g2_decap_8 FILLER_42_2586 ();
 sg13g2_decap_8 FILLER_42_2593 ();
 sg13g2_decap_8 FILLER_42_2600 ();
 sg13g2_decap_8 FILLER_42_2607 ();
 sg13g2_decap_8 FILLER_42_2614 ();
 sg13g2_decap_8 FILLER_42_2621 ();
 sg13g2_decap_8 FILLER_42_2628 ();
 sg13g2_decap_8 FILLER_42_2635 ();
 sg13g2_decap_8 FILLER_42_2642 ();
 sg13g2_decap_4 FILLER_42_2649 ();
 sg13g2_fill_1 FILLER_42_2653 ();
 sg13g2_decap_4 FILLER_42_2662 ();
 sg13g2_fill_1 FILLER_42_2666 ();
 sg13g2_decap_8 FILLER_42_2670 ();
 sg13g2_decap_8 FILLER_42_2677 ();
 sg13g2_decap_8 FILLER_42_2684 ();
 sg13g2_decap_8 FILLER_42_2691 ();
 sg13g2_decap_8 FILLER_42_2698 ();
 sg13g2_decap_8 FILLER_42_2759 ();
 sg13g2_decap_8 FILLER_42_2766 ();
 sg13g2_fill_2 FILLER_42_2773 ();
 sg13g2_decap_8 FILLER_42_2798 ();
 sg13g2_decap_4 FILLER_42_2805 ();
 sg13g2_fill_2 FILLER_42_2814 ();
 sg13g2_fill_1 FILLER_42_2816 ();
 sg13g2_decap_8 FILLER_42_2822 ();
 sg13g2_decap_8 FILLER_42_2829 ();
 sg13g2_decap_8 FILLER_42_2836 ();
 sg13g2_decap_8 FILLER_42_2843 ();
 sg13g2_fill_2 FILLER_42_2850 ();
 sg13g2_fill_1 FILLER_42_2852 ();
 sg13g2_decap_8 FILLER_42_2888 ();
 sg13g2_fill_1 FILLER_42_2895 ();
 sg13g2_decap_8 FILLER_42_2906 ();
 sg13g2_decap_8 FILLER_42_2913 ();
 sg13g2_decap_8 FILLER_42_2920 ();
 sg13g2_decap_8 FILLER_42_2927 ();
 sg13g2_decap_8 FILLER_42_2934 ();
 sg13g2_decap_8 FILLER_42_2941 ();
 sg13g2_decap_8 FILLER_42_2948 ();
 sg13g2_decap_8 FILLER_42_2955 ();
 sg13g2_decap_8 FILLER_42_2962 ();
 sg13g2_decap_8 FILLER_42_2969 ();
 sg13g2_decap_8 FILLER_42_2976 ();
 sg13g2_decap_4 FILLER_42_2983 ();
 sg13g2_fill_1 FILLER_42_2987 ();
 sg13g2_decap_4 FILLER_42_2994 ();
 sg13g2_fill_1 FILLER_42_2998 ();
 sg13g2_decap_8 FILLER_42_3003 ();
 sg13g2_decap_8 FILLER_42_3010 ();
 sg13g2_decap_8 FILLER_42_3017 ();
 sg13g2_decap_8 FILLER_42_3024 ();
 sg13g2_fill_2 FILLER_42_3031 ();
 sg13g2_decap_8 FILLER_42_3065 ();
 sg13g2_decap_8 FILLER_42_3072 ();
 sg13g2_decap_4 FILLER_42_3079 ();
 sg13g2_fill_2 FILLER_42_3083 ();
 sg13g2_fill_2 FILLER_42_3090 ();
 sg13g2_decap_8 FILLER_42_3103 ();
 sg13g2_fill_1 FILLER_42_3110 ();
 sg13g2_decap_8 FILLER_42_3116 ();
 sg13g2_decap_8 FILLER_42_3123 ();
 sg13g2_decap_4 FILLER_42_3130 ();
 sg13g2_decap_8 FILLER_42_3145 ();
 sg13g2_fill_2 FILLER_42_3152 ();
 sg13g2_fill_1 FILLER_42_3154 ();
 sg13g2_decap_4 FILLER_42_3158 ();
 sg13g2_fill_2 FILLER_42_3162 ();
 sg13g2_decap_8 FILLER_42_3167 ();
 sg13g2_decap_8 FILLER_42_3174 ();
 sg13g2_fill_2 FILLER_42_3181 ();
 sg13g2_decap_4 FILLER_42_3186 ();
 sg13g2_fill_2 FILLER_42_3190 ();
 sg13g2_fill_2 FILLER_42_3197 ();
 sg13g2_decap_8 FILLER_42_3221 ();
 sg13g2_decap_8 FILLER_42_3228 ();
 sg13g2_fill_1 FILLER_42_3235 ();
 sg13g2_decap_8 FILLER_42_3262 ();
 sg13g2_decap_8 FILLER_42_3269 ();
 sg13g2_decap_8 FILLER_42_3276 ();
 sg13g2_decap_8 FILLER_42_3283 ();
 sg13g2_decap_8 FILLER_42_3290 ();
 sg13g2_decap_8 FILLER_42_3307 ();
 sg13g2_decap_8 FILLER_42_3314 ();
 sg13g2_decap_8 FILLER_42_3321 ();
 sg13g2_fill_2 FILLER_42_3328 ();
 sg13g2_fill_1 FILLER_42_3330 ();
 sg13g2_fill_2 FILLER_42_3361 ();
 sg13g2_fill_1 FILLER_42_3363 ();
 sg13g2_decap_8 FILLER_42_3369 ();
 sg13g2_decap_8 FILLER_42_3376 ();
 sg13g2_decap_8 FILLER_42_3383 ();
 sg13g2_decap_8 FILLER_42_3390 ();
 sg13g2_decap_8 FILLER_42_3407 ();
 sg13g2_fill_2 FILLER_42_3414 ();
 sg13g2_decap_8 FILLER_42_3442 ();
 sg13g2_decap_8 FILLER_42_3449 ();
 sg13g2_decap_8 FILLER_42_3456 ();
 sg13g2_decap_8 FILLER_42_3463 ();
 sg13g2_decap_8 FILLER_42_3470 ();
 sg13g2_decap_8 FILLER_42_3477 ();
 sg13g2_decap_8 FILLER_42_3484 ();
 sg13g2_decap_8 FILLER_42_3491 ();
 sg13g2_decap_8 FILLER_42_3498 ();
 sg13g2_fill_2 FILLER_42_3505 ();
 sg13g2_fill_1 FILLER_42_3507 ();
 sg13g2_decap_8 FILLER_42_3517 ();
 sg13g2_decap_8 FILLER_42_3524 ();
 sg13g2_decap_8 FILLER_42_3531 ();
 sg13g2_fill_1 FILLER_42_3538 ();
 sg13g2_decap_8 FILLER_42_3573 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_4 FILLER_43_7 ();
 sg13g2_fill_1 FILLER_43_11 ();
 sg13g2_decap_8 FILLER_43_47 ();
 sg13g2_decap_8 FILLER_43_54 ();
 sg13g2_decap_8 FILLER_43_61 ();
 sg13g2_decap_4 FILLER_43_68 ();
 sg13g2_decap_8 FILLER_43_108 ();
 sg13g2_decap_4 FILLER_43_115 ();
 sg13g2_fill_2 FILLER_43_119 ();
 sg13g2_decap_8 FILLER_43_124 ();
 sg13g2_decap_8 FILLER_43_131 ();
 sg13g2_decap_4 FILLER_43_138 ();
 sg13g2_decap_8 FILLER_43_176 ();
 sg13g2_decap_8 FILLER_43_183 ();
 sg13g2_decap_8 FILLER_43_190 ();
 sg13g2_decap_8 FILLER_43_197 ();
 sg13g2_decap_4 FILLER_43_204 ();
 sg13g2_decap_8 FILLER_43_234 ();
 sg13g2_decap_4 FILLER_43_241 ();
 sg13g2_decap_4 FILLER_43_248 ();
 sg13g2_decap_8 FILLER_43_265 ();
 sg13g2_decap_8 FILLER_43_272 ();
 sg13g2_decap_8 FILLER_43_279 ();
 sg13g2_decap_8 FILLER_43_286 ();
 sg13g2_decap_8 FILLER_43_293 ();
 sg13g2_decap_8 FILLER_43_300 ();
 sg13g2_decap_8 FILLER_43_307 ();
 sg13g2_fill_1 FILLER_43_346 ();
 sg13g2_decap_8 FILLER_43_367 ();
 sg13g2_decap_8 FILLER_43_374 ();
 sg13g2_decap_8 FILLER_43_381 ();
 sg13g2_decap_8 FILLER_43_388 ();
 sg13g2_fill_2 FILLER_43_395 ();
 sg13g2_fill_1 FILLER_43_397 ();
 sg13g2_fill_1 FILLER_43_412 ();
 sg13g2_decap_8 FILLER_43_419 ();
 sg13g2_decap_8 FILLER_43_426 ();
 sg13g2_decap_8 FILLER_43_439 ();
 sg13g2_fill_2 FILLER_43_446 ();
 sg13g2_decap_8 FILLER_43_459 ();
 sg13g2_decap_8 FILLER_43_466 ();
 sg13g2_decap_8 FILLER_43_473 ();
 sg13g2_decap_8 FILLER_43_480 ();
 sg13g2_decap_8 FILLER_43_487 ();
 sg13g2_decap_8 FILLER_43_494 ();
 sg13g2_fill_1 FILLER_43_501 ();
 sg13g2_fill_2 FILLER_43_507 ();
 sg13g2_decap_8 FILLER_43_528 ();
 sg13g2_decap_8 FILLER_43_535 ();
 sg13g2_fill_1 FILLER_43_542 ();
 sg13g2_decap_4 FILLER_43_552 ();
 sg13g2_fill_1 FILLER_43_556 ();
 sg13g2_decap_8 FILLER_43_588 ();
 sg13g2_decap_8 FILLER_43_595 ();
 sg13g2_decap_8 FILLER_43_602 ();
 sg13g2_decap_8 FILLER_43_609 ();
 sg13g2_decap_8 FILLER_43_616 ();
 sg13g2_decap_8 FILLER_43_623 ();
 sg13g2_decap_8 FILLER_43_630 ();
 sg13g2_decap_8 FILLER_43_637 ();
 sg13g2_decap_8 FILLER_43_644 ();
 sg13g2_decap_8 FILLER_43_651 ();
 sg13g2_decap_8 FILLER_43_658 ();
 sg13g2_decap_4 FILLER_43_665 ();
 sg13g2_fill_1 FILLER_43_669 ();
 sg13g2_fill_2 FILLER_43_696 ();
 sg13g2_decap_4 FILLER_43_702 ();
 sg13g2_fill_2 FILLER_43_710 ();
 sg13g2_decap_8 FILLER_43_720 ();
 sg13g2_fill_2 FILLER_43_727 ();
 sg13g2_fill_1 FILLER_43_729 ();
 sg13g2_decap_8 FILLER_43_736 ();
 sg13g2_decap_8 FILLER_43_743 ();
 sg13g2_fill_2 FILLER_43_750 ();
 sg13g2_fill_1 FILLER_43_752 ();
 sg13g2_decap_8 FILLER_43_758 ();
 sg13g2_decap_8 FILLER_43_765 ();
 sg13g2_decap_8 FILLER_43_772 ();
 sg13g2_decap_4 FILLER_43_779 ();
 sg13g2_fill_2 FILLER_43_783 ();
 sg13g2_decap_4 FILLER_43_790 ();
 sg13g2_fill_1 FILLER_43_794 ();
 sg13g2_fill_2 FILLER_43_807 ();
 sg13g2_fill_1 FILLER_43_846 ();
 sg13g2_fill_1 FILLER_43_873 ();
 sg13g2_decap_8 FILLER_43_900 ();
 sg13g2_decap_8 FILLER_43_907 ();
 sg13g2_decap_8 FILLER_43_914 ();
 sg13g2_decap_8 FILLER_43_921 ();
 sg13g2_decap_8 FILLER_43_928 ();
 sg13g2_decap_8 FILLER_43_935 ();
 sg13g2_fill_2 FILLER_43_942 ();
 sg13g2_decap_8 FILLER_43_963 ();
 sg13g2_decap_8 FILLER_43_970 ();
 sg13g2_decap_8 FILLER_43_977 ();
 sg13g2_decap_8 FILLER_43_984 ();
 sg13g2_fill_2 FILLER_43_991 ();
 sg13g2_fill_1 FILLER_43_993 ();
 sg13g2_decap_4 FILLER_43_1007 ();
 sg13g2_fill_2 FILLER_43_1011 ();
 sg13g2_decap_8 FILLER_43_1021 ();
 sg13g2_fill_1 FILLER_43_1028 ();
 sg13g2_decap_8 FILLER_43_1049 ();
 sg13g2_decap_8 FILLER_43_1056 ();
 sg13g2_decap_8 FILLER_43_1063 ();
 sg13g2_fill_2 FILLER_43_1070 ();
 sg13g2_decap_4 FILLER_43_1086 ();
 sg13g2_decap_8 FILLER_43_1104 ();
 sg13g2_decap_4 FILLER_43_1111 ();
 sg13g2_fill_1 FILLER_43_1115 ();
 sg13g2_decap_8 FILLER_43_1122 ();
 sg13g2_decap_8 FILLER_43_1129 ();
 sg13g2_decap_8 FILLER_43_1136 ();
 sg13g2_decap_8 FILLER_43_1143 ();
 sg13g2_decap_8 FILLER_43_1150 ();
 sg13g2_decap_8 FILLER_43_1157 ();
 sg13g2_decap_8 FILLER_43_1164 ();
 sg13g2_decap_8 FILLER_43_1171 ();
 sg13g2_decap_8 FILLER_43_1183 ();
 sg13g2_decap_8 FILLER_43_1190 ();
 sg13g2_decap_8 FILLER_43_1197 ();
 sg13g2_decap_8 FILLER_43_1204 ();
 sg13g2_decap_8 FILLER_43_1211 ();
 sg13g2_decap_8 FILLER_43_1218 ();
 sg13g2_decap_8 FILLER_43_1225 ();
 sg13g2_decap_8 FILLER_43_1232 ();
 sg13g2_fill_1 FILLER_43_1239 ();
 sg13g2_decap_8 FILLER_43_1253 ();
 sg13g2_decap_8 FILLER_43_1260 ();
 sg13g2_decap_8 FILLER_43_1267 ();
 sg13g2_decap_8 FILLER_43_1274 ();
 sg13g2_decap_8 FILLER_43_1281 ();
 sg13g2_decap_8 FILLER_43_1288 ();
 sg13g2_decap_4 FILLER_43_1295 ();
 sg13g2_fill_1 FILLER_43_1299 ();
 sg13g2_decap_4 FILLER_43_1308 ();
 sg13g2_fill_1 FILLER_43_1312 ();
 sg13g2_decap_8 FILLER_43_1319 ();
 sg13g2_decap_8 FILLER_43_1326 ();
 sg13g2_decap_4 FILLER_43_1333 ();
 sg13g2_decap_8 FILLER_43_1373 ();
 sg13g2_decap_8 FILLER_43_1380 ();
 sg13g2_decap_8 FILLER_43_1387 ();
 sg13g2_decap_8 FILLER_43_1394 ();
 sg13g2_decap_8 FILLER_43_1401 ();
 sg13g2_decap_8 FILLER_43_1408 ();
 sg13g2_decap_4 FILLER_43_1415 ();
 sg13g2_fill_2 FILLER_43_1419 ();
 sg13g2_decap_8 FILLER_43_1452 ();
 sg13g2_decap_8 FILLER_43_1459 ();
 sg13g2_decap_8 FILLER_43_1466 ();
 sg13g2_fill_1 FILLER_43_1473 ();
 sg13g2_decap_8 FILLER_43_1497 ();
 sg13g2_decap_8 FILLER_43_1504 ();
 sg13g2_decap_8 FILLER_43_1511 ();
 sg13g2_decap_8 FILLER_43_1518 ();
 sg13g2_decap_8 FILLER_43_1525 ();
 sg13g2_decap_4 FILLER_43_1532 ();
 sg13g2_decap_8 FILLER_43_1562 ();
 sg13g2_decap_8 FILLER_43_1569 ();
 sg13g2_fill_2 FILLER_43_1576 ();
 sg13g2_fill_1 FILLER_43_1578 ();
 sg13g2_decap_4 FILLER_43_1585 ();
 sg13g2_decap_8 FILLER_43_1615 ();
 sg13g2_decap_8 FILLER_43_1622 ();
 sg13g2_decap_8 FILLER_43_1629 ();
 sg13g2_decap_8 FILLER_43_1636 ();
 sg13g2_decap_8 FILLER_43_1643 ();
 sg13g2_decap_8 FILLER_43_1650 ();
 sg13g2_fill_2 FILLER_43_1657 ();
 sg13g2_fill_1 FILLER_43_1659 ();
 sg13g2_decap_8 FILLER_43_1668 ();
 sg13g2_decap_8 FILLER_43_1675 ();
 sg13g2_decap_8 FILLER_43_1682 ();
 sg13g2_decap_8 FILLER_43_1689 ();
 sg13g2_decap_8 FILLER_43_1696 ();
 sg13g2_decap_8 FILLER_43_1703 ();
 sg13g2_decap_8 FILLER_43_1710 ();
 sg13g2_fill_1 FILLER_43_1717 ();
 sg13g2_decap_8 FILLER_43_1744 ();
 sg13g2_fill_1 FILLER_43_1751 ();
 sg13g2_decap_4 FILLER_43_1762 ();
 sg13g2_decap_8 FILLER_43_1772 ();
 sg13g2_decap_8 FILLER_43_1779 ();
 sg13g2_decap_8 FILLER_43_1786 ();
 sg13g2_decap_8 FILLER_43_1793 ();
 sg13g2_decap_4 FILLER_43_1800 ();
 sg13g2_decap_8 FILLER_43_1814 ();
 sg13g2_decap_8 FILLER_43_1821 ();
 sg13g2_decap_8 FILLER_43_1828 ();
 sg13g2_decap_8 FILLER_43_1835 ();
 sg13g2_decap_8 FILLER_43_1842 ();
 sg13g2_decap_8 FILLER_43_1849 ();
 sg13g2_decap_4 FILLER_43_1856 ();
 sg13g2_fill_2 FILLER_43_1860 ();
 sg13g2_decap_8 FILLER_43_1888 ();
 sg13g2_decap_8 FILLER_43_1895 ();
 sg13g2_decap_8 FILLER_43_1902 ();
 sg13g2_fill_2 FILLER_43_1909 ();
 sg13g2_decap_8 FILLER_43_1919 ();
 sg13g2_decap_8 FILLER_43_1926 ();
 sg13g2_decap_8 FILLER_43_1933 ();
 sg13g2_decap_8 FILLER_43_1940 ();
 sg13g2_decap_8 FILLER_43_1947 ();
 sg13g2_decap_8 FILLER_43_1954 ();
 sg13g2_fill_2 FILLER_43_1961 ();
 sg13g2_fill_1 FILLER_43_1963 ();
 sg13g2_decap_4 FILLER_43_1970 ();
 sg13g2_fill_1 FILLER_43_1974 ();
 sg13g2_fill_2 FILLER_43_1978 ();
 sg13g2_decap_4 FILLER_43_1999 ();
 sg13g2_fill_1 FILLER_43_2003 ();
 sg13g2_decap_8 FILLER_43_2010 ();
 sg13g2_decap_8 FILLER_43_2017 ();
 sg13g2_decap_8 FILLER_43_2024 ();
 sg13g2_decap_8 FILLER_43_2031 ();
 sg13g2_decap_8 FILLER_43_2046 ();
 sg13g2_decap_4 FILLER_43_2053 ();
 sg13g2_fill_1 FILLER_43_2057 ();
 sg13g2_decap_4 FILLER_43_2064 ();
 sg13g2_fill_1 FILLER_43_2068 ();
 sg13g2_decap_8 FILLER_43_2081 ();
 sg13g2_decap_4 FILLER_43_2088 ();
 sg13g2_decap_4 FILLER_43_2097 ();
 sg13g2_fill_2 FILLER_43_2119 ();
 sg13g2_decap_4 FILLER_43_2127 ();
 sg13g2_fill_1 FILLER_43_2131 ();
 sg13g2_fill_2 FILLER_43_2138 ();
 sg13g2_fill_1 FILLER_43_2140 ();
 sg13g2_fill_2 FILLER_43_2153 ();
 sg13g2_decap_4 FILLER_43_2178 ();
 sg13g2_decap_8 FILLER_43_2194 ();
 sg13g2_decap_8 FILLER_43_2201 ();
 sg13g2_decap_8 FILLER_43_2208 ();
 sg13g2_decap_8 FILLER_43_2215 ();
 sg13g2_decap_8 FILLER_43_2222 ();
 sg13g2_fill_2 FILLER_43_2238 ();
 sg13g2_fill_1 FILLER_43_2240 ();
 sg13g2_fill_1 FILLER_43_2246 ();
 sg13g2_decap_8 FILLER_43_2251 ();
 sg13g2_decap_4 FILLER_43_2258 ();
 sg13g2_decap_8 FILLER_43_2280 ();
 sg13g2_decap_8 FILLER_43_2287 ();
 sg13g2_decap_8 FILLER_43_2294 ();
 sg13g2_decap_8 FILLER_43_2301 ();
 sg13g2_decap_8 FILLER_43_2308 ();
 sg13g2_decap_8 FILLER_43_2315 ();
 sg13g2_decap_4 FILLER_43_2322 ();
 sg13g2_fill_1 FILLER_43_2326 ();
 sg13g2_decap_8 FILLER_43_2333 ();
 sg13g2_decap_8 FILLER_43_2340 ();
 sg13g2_decap_8 FILLER_43_2347 ();
 sg13g2_decap_8 FILLER_43_2354 ();
 sg13g2_decap_8 FILLER_43_2361 ();
 sg13g2_decap_8 FILLER_43_2368 ();
 sg13g2_decap_8 FILLER_43_2375 ();
 sg13g2_fill_1 FILLER_43_2382 ();
 sg13g2_decap_8 FILLER_43_2406 ();
 sg13g2_fill_1 FILLER_43_2413 ();
 sg13g2_decap_8 FILLER_43_2431 ();
 sg13g2_decap_4 FILLER_43_2438 ();
 sg13g2_fill_2 FILLER_43_2442 ();
 sg13g2_decap_8 FILLER_43_2450 ();
 sg13g2_fill_2 FILLER_43_2457 ();
 sg13g2_decap_8 FILLER_43_2467 ();
 sg13g2_fill_1 FILLER_43_2474 ();
 sg13g2_decap_8 FILLER_43_2493 ();
 sg13g2_decap_8 FILLER_43_2500 ();
 sg13g2_decap_4 FILLER_43_2507 ();
 sg13g2_fill_2 FILLER_43_2511 ();
 sg13g2_fill_2 FILLER_43_2524 ();
 sg13g2_decap_8 FILLER_43_2569 ();
 sg13g2_decap_8 FILLER_43_2576 ();
 sg13g2_decap_8 FILLER_43_2583 ();
 sg13g2_decap_4 FILLER_43_2590 ();
 sg13g2_fill_1 FILLER_43_2594 ();
 sg13g2_fill_2 FILLER_43_2603 ();
 sg13g2_decap_4 FILLER_43_2611 ();
 sg13g2_decap_8 FILLER_43_2625 ();
 sg13g2_decap_8 FILLER_43_2632 ();
 sg13g2_decap_8 FILLER_43_2639 ();
 sg13g2_decap_8 FILLER_43_2646 ();
 sg13g2_decap_8 FILLER_43_2653 ();
 sg13g2_fill_1 FILLER_43_2660 ();
 sg13g2_decap_8 FILLER_43_2687 ();
 sg13g2_fill_2 FILLER_43_2720 ();
 sg13g2_fill_1 FILLER_43_2722 ();
 sg13g2_decap_8 FILLER_43_2728 ();
 sg13g2_decap_8 FILLER_43_2735 ();
 sg13g2_decap_8 FILLER_43_2742 ();
 sg13g2_decap_8 FILLER_43_2749 ();
 sg13g2_decap_4 FILLER_43_2756 ();
 sg13g2_fill_1 FILLER_43_2760 ();
 sg13g2_decap_8 FILLER_43_2764 ();
 sg13g2_decap_4 FILLER_43_2771 ();
 sg13g2_fill_1 FILLER_43_2775 ();
 sg13g2_decap_8 FILLER_43_2781 ();
 sg13g2_decap_8 FILLER_43_2788 ();
 sg13g2_decap_8 FILLER_43_2795 ();
 sg13g2_decap_8 FILLER_43_2802 ();
 sg13g2_decap_8 FILLER_43_2809 ();
 sg13g2_decap_4 FILLER_43_2816 ();
 sg13g2_decap_8 FILLER_43_2825 ();
 sg13g2_decap_8 FILLER_43_2832 ();
 sg13g2_decap_8 FILLER_43_2839 ();
 sg13g2_decap_8 FILLER_43_2846 ();
 sg13g2_decap_8 FILLER_43_2853 ();
 sg13g2_decap_8 FILLER_43_2860 ();
 sg13g2_decap_8 FILLER_43_2867 ();
 sg13g2_decap_8 FILLER_43_2874 ();
 sg13g2_decap_8 FILLER_43_2881 ();
 sg13g2_decap_8 FILLER_43_2888 ();
 sg13g2_fill_2 FILLER_43_2895 ();
 sg13g2_decap_8 FILLER_43_2923 ();
 sg13g2_decap_8 FILLER_43_2930 ();
 sg13g2_decap_8 FILLER_43_2937 ();
 sg13g2_decap_8 FILLER_43_2944 ();
 sg13g2_fill_1 FILLER_43_2977 ();
 sg13g2_fill_2 FILLER_43_2986 ();
 sg13g2_fill_1 FILLER_43_2988 ();
 sg13g2_decap_8 FILLER_43_3015 ();
 sg13g2_decap_8 FILLER_43_3022 ();
 sg13g2_decap_8 FILLER_43_3055 ();
 sg13g2_decap_8 FILLER_43_3062 ();
 sg13g2_decap_8 FILLER_43_3069 ();
 sg13g2_decap_4 FILLER_43_3076 ();
 sg13g2_fill_1 FILLER_43_3080 ();
 sg13g2_decap_8 FILLER_43_3096 ();
 sg13g2_decap_4 FILLER_43_3103 ();
 sg13g2_fill_1 FILLER_43_3112 ();
 sg13g2_decap_8 FILLER_43_3128 ();
 sg13g2_decap_8 FILLER_43_3135 ();
 sg13g2_decap_8 FILLER_43_3142 ();
 sg13g2_decap_4 FILLER_43_3149 ();
 sg13g2_fill_2 FILLER_43_3153 ();
 sg13g2_decap_4 FILLER_43_3160 ();
 sg13g2_decap_8 FILLER_43_3169 ();
 sg13g2_decap_8 FILLER_43_3176 ();
 sg13g2_fill_1 FILLER_43_3198 ();
 sg13g2_decap_4 FILLER_43_3214 ();
 sg13g2_decap_8 FILLER_43_3226 ();
 sg13g2_decap_4 FILLER_43_3233 ();
 sg13g2_decap_8 FILLER_43_3258 ();
 sg13g2_decap_8 FILLER_43_3265 ();
 sg13g2_decap_8 FILLER_43_3272 ();
 sg13g2_decap_8 FILLER_43_3279 ();
 sg13g2_decap_8 FILLER_43_3286 ();
 sg13g2_decap_4 FILLER_43_3293 ();
 sg13g2_fill_1 FILLER_43_3297 ();
 sg13g2_fill_2 FILLER_43_3304 ();
 sg13g2_fill_1 FILLER_43_3316 ();
 sg13g2_decap_8 FILLER_43_3327 ();
 sg13g2_decap_8 FILLER_43_3334 ();
 sg13g2_decap_8 FILLER_43_3341 ();
 sg13g2_decap_8 FILLER_43_3348 ();
 sg13g2_decap_4 FILLER_43_3355 ();
 sg13g2_fill_1 FILLER_43_3359 ();
 sg13g2_decap_4 FILLER_43_3370 ();
 sg13g2_decap_8 FILLER_43_3400 ();
 sg13g2_decap_8 FILLER_43_3443 ();
 sg13g2_decap_8 FILLER_43_3450 ();
 sg13g2_decap_8 FILLER_43_3457 ();
 sg13g2_decap_8 FILLER_43_3464 ();
 sg13g2_decap_8 FILLER_43_3471 ();
 sg13g2_decap_4 FILLER_43_3478 ();
 sg13g2_fill_1 FILLER_43_3482 ();
 sg13g2_decap_8 FILLER_43_3509 ();
 sg13g2_decap_8 FILLER_43_3516 ();
 sg13g2_decap_8 FILLER_43_3523 ();
 sg13g2_decap_8 FILLER_43_3530 ();
 sg13g2_decap_8 FILLER_43_3537 ();
 sg13g2_decap_8 FILLER_43_3544 ();
 sg13g2_decap_8 FILLER_43_3551 ();
 sg13g2_decap_8 FILLER_43_3558 ();
 sg13g2_decap_8 FILLER_43_3565 ();
 sg13g2_decap_8 FILLER_43_3572 ();
 sg13g2_fill_1 FILLER_43_3579 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_fill_2 FILLER_44_14 ();
 sg13g2_fill_1 FILLER_44_30 ();
 sg13g2_decap_8 FILLER_44_49 ();
 sg13g2_decap_8 FILLER_44_56 ();
 sg13g2_decap_4 FILLER_44_63 ();
 sg13g2_decap_4 FILLER_44_93 ();
 sg13g2_decap_8 FILLER_44_106 ();
 sg13g2_decap_4 FILLER_44_149 ();
 sg13g2_decap_8 FILLER_44_166 ();
 sg13g2_fill_1 FILLER_44_173 ();
 sg13g2_decap_8 FILLER_44_183 ();
 sg13g2_decap_8 FILLER_44_190 ();
 sg13g2_decap_8 FILLER_44_197 ();
 sg13g2_decap_8 FILLER_44_204 ();
 sg13g2_decap_4 FILLER_44_211 ();
 sg13g2_fill_2 FILLER_44_215 ();
 sg13g2_decap_8 FILLER_44_227 ();
 sg13g2_decap_4 FILLER_44_234 ();
 sg13g2_fill_2 FILLER_44_238 ();
 sg13g2_decap_8 FILLER_44_249 ();
 sg13g2_decap_8 FILLER_44_256 ();
 sg13g2_decap_8 FILLER_44_263 ();
 sg13g2_decap_8 FILLER_44_270 ();
 sg13g2_decap_8 FILLER_44_277 ();
 sg13g2_decap_8 FILLER_44_284 ();
 sg13g2_decap_8 FILLER_44_291 ();
 sg13g2_decap_8 FILLER_44_298 ();
 sg13g2_decap_4 FILLER_44_305 ();
 sg13g2_fill_2 FILLER_44_347 ();
 sg13g2_fill_1 FILLER_44_349 ();
 sg13g2_decap_8 FILLER_44_357 ();
 sg13g2_decap_4 FILLER_44_364 ();
 sg13g2_decap_8 FILLER_44_394 ();
 sg13g2_decap_8 FILLER_44_401 ();
 sg13g2_decap_8 FILLER_44_408 ();
 sg13g2_decap_4 FILLER_44_415 ();
 sg13g2_decap_8 FILLER_44_425 ();
 sg13g2_decap_8 FILLER_44_432 ();
 sg13g2_decap_8 FILLER_44_445 ();
 sg13g2_fill_2 FILLER_44_452 ();
 sg13g2_fill_1 FILLER_44_454 ();
 sg13g2_decap_4 FILLER_44_463 ();
 sg13g2_fill_1 FILLER_44_467 ();
 sg13g2_decap_4 FILLER_44_477 ();
 sg13g2_decap_8 FILLER_44_485 ();
 sg13g2_decap_8 FILLER_44_492 ();
 sg13g2_decap_4 FILLER_44_499 ();
 sg13g2_fill_1 FILLER_44_503 ();
 sg13g2_fill_1 FILLER_44_532 ();
 sg13g2_fill_1 FILLER_44_558 ();
 sg13g2_decap_8 FILLER_44_585 ();
 sg13g2_decap_8 FILLER_44_592 ();
 sg13g2_decap_8 FILLER_44_599 ();
 sg13g2_decap_8 FILLER_44_606 ();
 sg13g2_decap_8 FILLER_44_613 ();
 sg13g2_decap_8 FILLER_44_620 ();
 sg13g2_fill_1 FILLER_44_627 ();
 sg13g2_decap_4 FILLER_44_634 ();
 sg13g2_fill_1 FILLER_44_638 ();
 sg13g2_decap_4 FILLER_44_644 ();
 sg13g2_fill_1 FILLER_44_648 ();
 sg13g2_fill_2 FILLER_44_657 ();
 sg13g2_fill_2 FILLER_44_665 ();
 sg13g2_fill_1 FILLER_44_667 ();
 sg13g2_decap_8 FILLER_44_691 ();
 sg13g2_decap_8 FILLER_44_698 ();
 sg13g2_decap_8 FILLER_44_705 ();
 sg13g2_decap_8 FILLER_44_727 ();
 sg13g2_decap_4 FILLER_44_734 ();
 sg13g2_fill_2 FILLER_44_738 ();
 sg13g2_decap_4 FILLER_44_745 ();
 sg13g2_fill_2 FILLER_44_749 ();
 sg13g2_fill_2 FILLER_44_756 ();
 sg13g2_fill_1 FILLER_44_758 ();
 sg13g2_decap_8 FILLER_44_762 ();
 sg13g2_decap_4 FILLER_44_769 ();
 sg13g2_fill_2 FILLER_44_783 ();
 sg13g2_fill_1 FILLER_44_785 ();
 sg13g2_decap_8 FILLER_44_803 ();
 sg13g2_decap_4 FILLER_44_810 ();
 sg13g2_decap_8 FILLER_44_818 ();
 sg13g2_decap_4 FILLER_44_825 ();
 sg13g2_fill_1 FILLER_44_829 ();
 sg13g2_fill_2 FILLER_44_843 ();
 sg13g2_decap_8 FILLER_44_853 ();
 sg13g2_decap_8 FILLER_44_860 ();
 sg13g2_decap_8 FILLER_44_867 ();
 sg13g2_decap_8 FILLER_44_874 ();
 sg13g2_fill_1 FILLER_44_881 ();
 sg13g2_decap_8 FILLER_44_895 ();
 sg13g2_decap_8 FILLER_44_902 ();
 sg13g2_decap_8 FILLER_44_909 ();
 sg13g2_decap_8 FILLER_44_916 ();
 sg13g2_decap_8 FILLER_44_923 ();
 sg13g2_decap_8 FILLER_44_930 ();
 sg13g2_fill_2 FILLER_44_937 ();
 sg13g2_fill_1 FILLER_44_955 ();
 sg13g2_fill_2 FILLER_44_969 ();
 sg13g2_decap_8 FILLER_44_976 ();
 sg13g2_fill_2 FILLER_44_983 ();
 sg13g2_fill_1 FILLER_44_985 ();
 sg13g2_decap_8 FILLER_44_993 ();
 sg13g2_decap_8 FILLER_44_1000 ();
 sg13g2_decap_8 FILLER_44_1007 ();
 sg13g2_decap_8 FILLER_44_1014 ();
 sg13g2_decap_8 FILLER_44_1021 ();
 sg13g2_decap_8 FILLER_44_1028 ();
 sg13g2_decap_8 FILLER_44_1035 ();
 sg13g2_decap_8 FILLER_44_1042 ();
 sg13g2_decap_8 FILLER_44_1049 ();
 sg13g2_fill_2 FILLER_44_1056 ();
 sg13g2_decap_8 FILLER_44_1089 ();
 sg13g2_decap_8 FILLER_44_1096 ();
 sg13g2_decap_8 FILLER_44_1103 ();
 sg13g2_fill_2 FILLER_44_1110 ();
 sg13g2_fill_1 FILLER_44_1112 ();
 sg13g2_decap_8 FILLER_44_1152 ();
 sg13g2_decap_8 FILLER_44_1159 ();
 sg13g2_decap_8 FILLER_44_1166 ();
 sg13g2_decap_8 FILLER_44_1173 ();
 sg13g2_decap_4 FILLER_44_1180 ();
 sg13g2_fill_1 FILLER_44_1184 ();
 sg13g2_decap_8 FILLER_44_1188 ();
 sg13g2_decap_8 FILLER_44_1195 ();
 sg13g2_decap_8 FILLER_44_1202 ();
 sg13g2_decap_8 FILLER_44_1209 ();
 sg13g2_decap_8 FILLER_44_1216 ();
 sg13g2_fill_2 FILLER_44_1223 ();
 sg13g2_fill_1 FILLER_44_1225 ();
 sg13g2_decap_8 FILLER_44_1262 ();
 sg13g2_decap_8 FILLER_44_1269 ();
 sg13g2_decap_8 FILLER_44_1276 ();
 sg13g2_fill_2 FILLER_44_1283 ();
 sg13g2_decap_8 FILLER_44_1311 ();
 sg13g2_decap_8 FILLER_44_1318 ();
 sg13g2_decap_8 FILLER_44_1325 ();
 sg13g2_decap_8 FILLER_44_1332 ();
 sg13g2_decap_8 FILLER_44_1339 ();
 sg13g2_fill_1 FILLER_44_1346 ();
 sg13g2_decap_4 FILLER_44_1358 ();
 sg13g2_decap_8 FILLER_44_1368 ();
 sg13g2_decap_8 FILLER_44_1375 ();
 sg13g2_decap_8 FILLER_44_1382 ();
 sg13g2_fill_2 FILLER_44_1389 ();
 sg13g2_fill_1 FILLER_44_1391 ();
 sg13g2_decap_8 FILLER_44_1400 ();
 sg13g2_decap_8 FILLER_44_1407 ();
 sg13g2_decap_8 FILLER_44_1414 ();
 sg13g2_decap_8 FILLER_44_1421 ();
 sg13g2_decap_8 FILLER_44_1428 ();
 sg13g2_decap_8 FILLER_44_1435 ();
 sg13g2_decap_8 FILLER_44_1456 ();
 sg13g2_decap_8 FILLER_44_1463 ();
 sg13g2_decap_8 FILLER_44_1470 ();
 sg13g2_decap_8 FILLER_44_1477 ();
 sg13g2_decap_8 FILLER_44_1484 ();
 sg13g2_decap_8 FILLER_44_1491 ();
 sg13g2_decap_8 FILLER_44_1498 ();
 sg13g2_decap_8 FILLER_44_1505 ();
 sg13g2_decap_8 FILLER_44_1512 ();
 sg13g2_decap_8 FILLER_44_1519 ();
 sg13g2_decap_8 FILLER_44_1526 ();
 sg13g2_decap_4 FILLER_44_1533 ();
 sg13g2_fill_1 FILLER_44_1537 ();
 sg13g2_decap_8 FILLER_44_1548 ();
 sg13g2_decap_8 FILLER_44_1555 ();
 sg13g2_decap_8 FILLER_44_1562 ();
 sg13g2_fill_2 FILLER_44_1569 ();
 sg13g2_fill_1 FILLER_44_1571 ();
 sg13g2_decap_8 FILLER_44_1619 ();
 sg13g2_fill_2 FILLER_44_1626 ();
 sg13g2_fill_1 FILLER_44_1628 ();
 sg13g2_decap_4 FILLER_44_1665 ();
 sg13g2_fill_1 FILLER_44_1669 ();
 sg13g2_decap_8 FILLER_44_1691 ();
 sg13g2_fill_1 FILLER_44_1698 ();
 sg13g2_decap_8 FILLER_44_1715 ();
 sg13g2_decap_8 FILLER_44_1722 ();
 sg13g2_decap_8 FILLER_44_1729 ();
 sg13g2_decap_8 FILLER_44_1736 ();
 sg13g2_decap_8 FILLER_44_1743 ();
 sg13g2_fill_1 FILLER_44_1750 ();
 sg13g2_decap_8 FILLER_44_1777 ();
 sg13g2_decap_8 FILLER_44_1784 ();
 sg13g2_decap_8 FILLER_44_1791 ();
 sg13g2_fill_2 FILLER_44_1798 ();
 sg13g2_fill_1 FILLER_44_1800 ();
 sg13g2_decap_8 FILLER_44_1838 ();
 sg13g2_decap_8 FILLER_44_1845 ();
 sg13g2_decap_8 FILLER_44_1852 ();
 sg13g2_decap_8 FILLER_44_1859 ();
 sg13g2_decap_8 FILLER_44_1866 ();
 sg13g2_decap_8 FILLER_44_1873 ();
 sg13g2_decap_8 FILLER_44_1880 ();
 sg13g2_decap_8 FILLER_44_1887 ();
 sg13g2_decap_8 FILLER_44_1894 ();
 sg13g2_decap_8 FILLER_44_1901 ();
 sg13g2_fill_2 FILLER_44_1919 ();
 sg13g2_fill_1 FILLER_44_1921 ();
 sg13g2_decap_8 FILLER_44_1928 ();
 sg13g2_decap_8 FILLER_44_1935 ();
 sg13g2_fill_2 FILLER_44_1942 ();
 sg13g2_decap_8 FILLER_44_1954 ();
 sg13g2_fill_1 FILLER_44_1961 ();
 sg13g2_decap_8 FILLER_44_2002 ();
 sg13g2_decap_8 FILLER_44_2009 ();
 sg13g2_decap_8 FILLER_44_2016 ();
 sg13g2_fill_1 FILLER_44_2023 ();
 sg13g2_decap_8 FILLER_44_2039 ();
 sg13g2_fill_1 FILLER_44_2046 ();
 sg13g2_decap_8 FILLER_44_2057 ();
 sg13g2_decap_8 FILLER_44_2064 ();
 sg13g2_decap_8 FILLER_44_2071 ();
 sg13g2_decap_8 FILLER_44_2078 ();
 sg13g2_fill_2 FILLER_44_2095 ();
 sg13g2_fill_1 FILLER_44_2097 ();
 sg13g2_decap_8 FILLER_44_2104 ();
 sg13g2_decap_8 FILLER_44_2111 ();
 sg13g2_fill_2 FILLER_44_2118 ();
 sg13g2_decap_8 FILLER_44_2128 ();
 sg13g2_decap_8 FILLER_44_2156 ();
 sg13g2_fill_2 FILLER_44_2163 ();
 sg13g2_fill_1 FILLER_44_2165 ();
 sg13g2_decap_8 FILLER_44_2169 ();
 sg13g2_decap_8 FILLER_44_2176 ();
 sg13g2_decap_8 FILLER_44_2183 ();
 sg13g2_decap_8 FILLER_44_2190 ();
 sg13g2_decap_4 FILLER_44_2197 ();
 sg13g2_decap_8 FILLER_44_2221 ();
 sg13g2_fill_1 FILLER_44_2228 ();
 sg13g2_fill_2 FILLER_44_2241 ();
 sg13g2_decap_4 FILLER_44_2257 ();
 sg13g2_decap_8 FILLER_44_2264 ();
 sg13g2_fill_2 FILLER_44_2271 ();
 sg13g2_decap_8 FILLER_44_2277 ();
 sg13g2_decap_8 FILLER_44_2284 ();
 sg13g2_fill_2 FILLER_44_2291 ();
 sg13g2_decap_8 FILLER_44_2296 ();
 sg13g2_decap_8 FILLER_44_2303 ();
 sg13g2_decap_4 FILLER_44_2310 ();
 sg13g2_fill_1 FILLER_44_2314 ();
 sg13g2_decap_8 FILLER_44_2340 ();
 sg13g2_decap_8 FILLER_44_2365 ();
 sg13g2_fill_2 FILLER_44_2372 ();
 sg13g2_fill_2 FILLER_44_2380 ();
 sg13g2_fill_1 FILLER_44_2382 ();
 sg13g2_decap_8 FILLER_44_2419 ();
 sg13g2_decap_8 FILLER_44_2426 ();
 sg13g2_decap_8 FILLER_44_2433 ();
 sg13g2_decap_4 FILLER_44_2440 ();
 sg13g2_fill_2 FILLER_44_2444 ();
 sg13g2_decap_8 FILLER_44_2456 ();
 sg13g2_decap_4 FILLER_44_2463 ();
 sg13g2_fill_2 FILLER_44_2467 ();
 sg13g2_fill_1 FILLER_44_2475 ();
 sg13g2_decap_4 FILLER_44_2482 ();
 sg13g2_decap_8 FILLER_44_2492 ();
 sg13g2_decap_8 FILLER_44_2499 ();
 sg13g2_decap_4 FILLER_44_2506 ();
 sg13g2_decap_8 FILLER_44_2519 ();
 sg13g2_decap_4 FILLER_44_2529 ();
 sg13g2_fill_2 FILLER_44_2533 ();
 sg13g2_decap_8 FILLER_44_2541 ();
 sg13g2_decap_8 FILLER_44_2548 ();
 sg13g2_decap_8 FILLER_44_2555 ();
 sg13g2_decap_8 FILLER_44_2562 ();
 sg13g2_decap_8 FILLER_44_2569 ();
 sg13g2_fill_2 FILLER_44_2576 ();
 sg13g2_decap_8 FILLER_44_2583 ();
 sg13g2_decap_8 FILLER_44_2590 ();
 sg13g2_decap_8 FILLER_44_2597 ();
 sg13g2_decap_8 FILLER_44_2604 ();
 sg13g2_decap_8 FILLER_44_2641 ();
 sg13g2_fill_1 FILLER_44_2648 ();
 sg13g2_decap_8 FILLER_44_2655 ();
 sg13g2_decap_8 FILLER_44_2672 ();
 sg13g2_decap_8 FILLER_44_2679 ();
 sg13g2_decap_8 FILLER_44_2686 ();
 sg13g2_decap_8 FILLER_44_2693 ();
 sg13g2_decap_8 FILLER_44_2700 ();
 sg13g2_decap_8 FILLER_44_2707 ();
 sg13g2_decap_4 FILLER_44_2714 ();
 sg13g2_decap_8 FILLER_44_2744 ();
 sg13g2_decap_8 FILLER_44_2751 ();
 sg13g2_decap_8 FILLER_44_2758 ();
 sg13g2_decap_8 FILLER_44_2765 ();
 sg13g2_decap_4 FILLER_44_2772 ();
 sg13g2_decap_8 FILLER_44_2786 ();
 sg13g2_decap_8 FILLER_44_2793 ();
 sg13g2_decap_8 FILLER_44_2800 ();
 sg13g2_decap_8 FILLER_44_2807 ();
 sg13g2_decap_8 FILLER_44_2814 ();
 sg13g2_fill_2 FILLER_44_2821 ();
 sg13g2_decap_8 FILLER_44_2827 ();
 sg13g2_decap_8 FILLER_44_2834 ();
 sg13g2_decap_8 FILLER_44_2841 ();
 sg13g2_decap_8 FILLER_44_2848 ();
 sg13g2_decap_8 FILLER_44_2855 ();
 sg13g2_decap_8 FILLER_44_2862 ();
 sg13g2_decap_4 FILLER_44_2869 ();
 sg13g2_decap_8 FILLER_44_2919 ();
 sg13g2_decap_4 FILLER_44_2926 ();
 sg13g2_fill_1 FILLER_44_2930 ();
 sg13g2_decap_8 FILLER_44_2941 ();
 sg13g2_decap_8 FILLER_44_2948 ();
 sg13g2_decap_8 FILLER_44_2955 ();
 sg13g2_fill_2 FILLER_44_2962 ();
 sg13g2_fill_1 FILLER_44_3000 ();
 sg13g2_decap_8 FILLER_44_3013 ();
 sg13g2_decap_8 FILLER_44_3020 ();
 sg13g2_fill_2 FILLER_44_3027 ();
 sg13g2_fill_1 FILLER_44_3029 ();
 sg13g2_decap_8 FILLER_44_3050 ();
 sg13g2_decap_8 FILLER_44_3057 ();
 sg13g2_decap_8 FILLER_44_3064 ();
 sg13g2_decap_8 FILLER_44_3071 ();
 sg13g2_decap_8 FILLER_44_3140 ();
 sg13g2_fill_2 FILLER_44_3147 ();
 sg13g2_fill_1 FILLER_44_3149 ();
 sg13g2_fill_2 FILLER_44_3155 ();
 sg13g2_fill_1 FILLER_44_3178 ();
 sg13g2_decap_8 FILLER_44_3209 ();
 sg13g2_decap_8 FILLER_44_3216 ();
 sg13g2_decap_8 FILLER_44_3223 ();
 sg13g2_decap_8 FILLER_44_3230 ();
 sg13g2_decap_8 FILLER_44_3237 ();
 sg13g2_decap_8 FILLER_44_3244 ();
 sg13g2_decap_8 FILLER_44_3251 ();
 sg13g2_decap_8 FILLER_44_3258 ();
 sg13g2_decap_8 FILLER_44_3265 ();
 sg13g2_decap_8 FILLER_44_3272 ();
 sg13g2_decap_8 FILLER_44_3279 ();
 sg13g2_decap_8 FILLER_44_3286 ();
 sg13g2_decap_8 FILLER_44_3293 ();
 sg13g2_decap_4 FILLER_44_3314 ();
 sg13g2_decap_4 FILLER_44_3328 ();
 sg13g2_fill_1 FILLER_44_3358 ();
 sg13g2_decap_8 FILLER_44_3385 ();
 sg13g2_decap_8 FILLER_44_3392 ();
 sg13g2_decap_8 FILLER_44_3399 ();
 sg13g2_decap_4 FILLER_44_3406 ();
 sg13g2_fill_1 FILLER_44_3410 ();
 sg13g2_decap_8 FILLER_44_3421 ();
 sg13g2_decap_8 FILLER_44_3428 ();
 sg13g2_decap_8 FILLER_44_3435 ();
 sg13g2_decap_8 FILLER_44_3442 ();
 sg13g2_decap_8 FILLER_44_3449 ();
 sg13g2_decap_8 FILLER_44_3456 ();
 sg13g2_decap_8 FILLER_44_3463 ();
 sg13g2_decap_4 FILLER_44_3470 ();
 sg13g2_decap_8 FILLER_44_3504 ();
 sg13g2_decap_8 FILLER_44_3511 ();
 sg13g2_decap_8 FILLER_44_3518 ();
 sg13g2_decap_8 FILLER_44_3525 ();
 sg13g2_decap_8 FILLER_44_3532 ();
 sg13g2_decap_8 FILLER_44_3539 ();
 sg13g2_decap_8 FILLER_44_3572 ();
 sg13g2_fill_1 FILLER_44_3579 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_7 ();
 sg13g2_decap_4 FILLER_45_14 ();
 sg13g2_fill_2 FILLER_45_18 ();
 sg13g2_fill_1 FILLER_45_34 ();
 sg13g2_decap_8 FILLER_45_40 ();
 sg13g2_decap_8 FILLER_45_47 ();
 sg13g2_decap_8 FILLER_45_54 ();
 sg13g2_decap_8 FILLER_45_61 ();
 sg13g2_decap_8 FILLER_45_68 ();
 sg13g2_decap_8 FILLER_45_75 ();
 sg13g2_decap_8 FILLER_45_82 ();
 sg13g2_decap_8 FILLER_45_94 ();
 sg13g2_decap_4 FILLER_45_101 ();
 sg13g2_fill_1 FILLER_45_105 ();
 sg13g2_decap_8 FILLER_45_146 ();
 sg13g2_decap_8 FILLER_45_153 ();
 sg13g2_decap_8 FILLER_45_160 ();
 sg13g2_decap_8 FILLER_45_167 ();
 sg13g2_decap_8 FILLER_45_174 ();
 sg13g2_decap_8 FILLER_45_181 ();
 sg13g2_decap_8 FILLER_45_188 ();
 sg13g2_decap_8 FILLER_45_195 ();
 sg13g2_decap_8 FILLER_45_202 ();
 sg13g2_decap_8 FILLER_45_209 ();
 sg13g2_decap_8 FILLER_45_216 ();
 sg13g2_decap_8 FILLER_45_223 ();
 sg13g2_decap_8 FILLER_45_230 ();
 sg13g2_decap_8 FILLER_45_237 ();
 sg13g2_decap_8 FILLER_45_244 ();
 sg13g2_decap_8 FILLER_45_251 ();
 sg13g2_decap_8 FILLER_45_258 ();
 sg13g2_decap_4 FILLER_45_265 ();
 sg13g2_fill_2 FILLER_45_269 ();
 sg13g2_decap_8 FILLER_45_287 ();
 sg13g2_decap_8 FILLER_45_294 ();
 sg13g2_decap_8 FILLER_45_301 ();
 sg13g2_decap_8 FILLER_45_308 ();
 sg13g2_decap_8 FILLER_45_315 ();
 sg13g2_decap_8 FILLER_45_322 ();
 sg13g2_decap_8 FILLER_45_338 ();
 sg13g2_decap_8 FILLER_45_345 ();
 sg13g2_fill_2 FILLER_45_352 ();
 sg13g2_decap_8 FILLER_45_361 ();
 sg13g2_decap_8 FILLER_45_368 ();
 sg13g2_decap_8 FILLER_45_375 ();
 sg13g2_decap_4 FILLER_45_382 ();
 sg13g2_fill_1 FILLER_45_386 ();
 sg13g2_decap_8 FILLER_45_399 ();
 sg13g2_decap_8 FILLER_45_406 ();
 sg13g2_fill_1 FILLER_45_413 ();
 sg13g2_decap_4 FILLER_45_420 ();
 sg13g2_fill_1 FILLER_45_424 ();
 sg13g2_decap_4 FILLER_45_431 ();
 sg13g2_fill_1 FILLER_45_435 ();
 sg13g2_fill_2 FILLER_45_466 ();
 sg13g2_decap_8 FILLER_45_492 ();
 sg13g2_decap_8 FILLER_45_499 ();
 sg13g2_decap_4 FILLER_45_506 ();
 sg13g2_fill_1 FILLER_45_510 ();
 sg13g2_fill_1 FILLER_45_548 ();
 sg13g2_decap_8 FILLER_45_602 ();
 sg13g2_decap_8 FILLER_45_609 ();
 sg13g2_decap_4 FILLER_45_616 ();
 sg13g2_fill_1 FILLER_45_620 ();
 sg13g2_decap_4 FILLER_45_624 ();
 sg13g2_fill_2 FILLER_45_628 ();
 sg13g2_decap_8 FILLER_45_655 ();
 sg13g2_decap_8 FILLER_45_662 ();
 sg13g2_decap_4 FILLER_45_669 ();
 sg13g2_decap_8 FILLER_45_699 ();
 sg13g2_decap_4 FILLER_45_706 ();
 sg13g2_decap_8 FILLER_45_718 ();
 sg13g2_decap_8 FILLER_45_725 ();
 sg13g2_decap_8 FILLER_45_732 ();
 sg13g2_decap_8 FILLER_45_739 ();
 sg13g2_fill_1 FILLER_45_746 ();
 sg13g2_decap_4 FILLER_45_755 ();
 sg13g2_decap_8 FILLER_45_764 ();
 sg13g2_decap_8 FILLER_45_771 ();
 sg13g2_decap_8 FILLER_45_778 ();
 sg13g2_decap_8 FILLER_45_785 ();
 sg13g2_decap_8 FILLER_45_792 ();
 sg13g2_decap_8 FILLER_45_799 ();
 sg13g2_decap_8 FILLER_45_806 ();
 sg13g2_decap_8 FILLER_45_813 ();
 sg13g2_fill_1 FILLER_45_820 ();
 sg13g2_decap_8 FILLER_45_847 ();
 sg13g2_decap_8 FILLER_45_854 ();
 sg13g2_decap_8 FILLER_45_861 ();
 sg13g2_decap_8 FILLER_45_868 ();
 sg13g2_decap_8 FILLER_45_875 ();
 sg13g2_decap_8 FILLER_45_882 ();
 sg13g2_decap_8 FILLER_45_889 ();
 sg13g2_decap_8 FILLER_45_896 ();
 sg13g2_decap_4 FILLER_45_903 ();
 sg13g2_fill_1 FILLER_45_907 ();
 sg13g2_decap_8 FILLER_45_921 ();
 sg13g2_fill_2 FILLER_45_928 ();
 sg13g2_fill_1 FILLER_45_930 ();
 sg13g2_decap_8 FILLER_45_935 ();
 sg13g2_fill_2 FILLER_45_942 ();
 sg13g2_fill_1 FILLER_45_944 ();
 sg13g2_decap_8 FILLER_45_980 ();
 sg13g2_fill_2 FILLER_45_987 ();
 sg13g2_decap_8 FILLER_45_997 ();
 sg13g2_decap_8 FILLER_45_1004 ();
 sg13g2_decap_4 FILLER_45_1011 ();
 sg13g2_fill_1 FILLER_45_1015 ();
 sg13g2_decap_8 FILLER_45_1028 ();
 sg13g2_decap_8 FILLER_45_1035 ();
 sg13g2_decap_8 FILLER_45_1042 ();
 sg13g2_fill_2 FILLER_45_1049 ();
 sg13g2_fill_1 FILLER_45_1051 ();
 sg13g2_decap_4 FILLER_45_1057 ();
 sg13g2_fill_2 FILLER_45_1061 ();
 sg13g2_decap_8 FILLER_45_1098 ();
 sg13g2_decap_8 FILLER_45_1105 ();
 sg13g2_decap_4 FILLER_45_1112 ();
 sg13g2_decap_8 FILLER_45_1142 ();
 sg13g2_decap_8 FILLER_45_1168 ();
 sg13g2_decap_8 FILLER_45_1175 ();
 sg13g2_decap_8 FILLER_45_1199 ();
 sg13g2_decap_8 FILLER_45_1206 ();
 sg13g2_decap_8 FILLER_45_1213 ();
 sg13g2_decap_4 FILLER_45_1220 ();
 sg13g2_fill_1 FILLER_45_1224 ();
 sg13g2_fill_2 FILLER_45_1230 ();
 sg13g2_fill_1 FILLER_45_1232 ();
 sg13g2_decap_8 FILLER_45_1243 ();
 sg13g2_decap_8 FILLER_45_1250 ();
 sg13g2_decap_8 FILLER_45_1257 ();
 sg13g2_decap_4 FILLER_45_1264 ();
 sg13g2_fill_1 FILLER_45_1268 ();
 sg13g2_fill_2 FILLER_45_1289 ();
 sg13g2_fill_1 FILLER_45_1291 ();
 sg13g2_decap_8 FILLER_45_1318 ();
 sg13g2_decap_8 FILLER_45_1325 ();
 sg13g2_decap_8 FILLER_45_1332 ();
 sg13g2_decap_8 FILLER_45_1365 ();
 sg13g2_decap_8 FILLER_45_1372 ();
 sg13g2_decap_8 FILLER_45_1379 ();
 sg13g2_decap_8 FILLER_45_1386 ();
 sg13g2_decap_4 FILLER_45_1393 ();
 sg13g2_fill_2 FILLER_45_1397 ();
 sg13g2_decap_8 FILLER_45_1404 ();
 sg13g2_decap_8 FILLER_45_1411 ();
 sg13g2_decap_8 FILLER_45_1428 ();
 sg13g2_decap_8 FILLER_45_1435 ();
 sg13g2_decap_8 FILLER_45_1442 ();
 sg13g2_decap_8 FILLER_45_1449 ();
 sg13g2_decap_8 FILLER_45_1456 ();
 sg13g2_fill_2 FILLER_45_1463 ();
 sg13g2_decap_8 FILLER_45_1501 ();
 sg13g2_decap_8 FILLER_45_1508 ();
 sg13g2_decap_8 FILLER_45_1515 ();
 sg13g2_decap_8 FILLER_45_1522 ();
 sg13g2_decap_8 FILLER_45_1529 ();
 sg13g2_decap_8 FILLER_45_1536 ();
 sg13g2_decap_8 FILLER_45_1543 ();
 sg13g2_decap_8 FILLER_45_1550 ();
 sg13g2_decap_8 FILLER_45_1557 ();
 sg13g2_decap_8 FILLER_45_1564 ();
 sg13g2_decap_8 FILLER_45_1571 ();
 sg13g2_decap_8 FILLER_45_1578 ();
 sg13g2_decap_8 FILLER_45_1585 ();
 sg13g2_decap_4 FILLER_45_1592 ();
 sg13g2_decap_8 FILLER_45_1612 ();
 sg13g2_decap_8 FILLER_45_1619 ();
 sg13g2_decap_8 FILLER_45_1626 ();
 sg13g2_fill_1 FILLER_45_1633 ();
 sg13g2_decap_8 FILLER_45_1670 ();
 sg13g2_decap_8 FILLER_45_1677 ();
 sg13g2_decap_8 FILLER_45_1684 ();
 sg13g2_decap_8 FILLER_45_1691 ();
 sg13g2_fill_1 FILLER_45_1698 ();
 sg13g2_decap_8 FILLER_45_1725 ();
 sg13g2_decap_8 FILLER_45_1732 ();
 sg13g2_decap_8 FILLER_45_1739 ();
 sg13g2_decap_8 FILLER_45_1746 ();
 sg13g2_decap_8 FILLER_45_1753 ();
 sg13g2_fill_2 FILLER_45_1760 ();
 sg13g2_fill_1 FILLER_45_1762 ();
 sg13g2_decap_8 FILLER_45_1773 ();
 sg13g2_decap_8 FILLER_45_1780 ();
 sg13g2_decap_8 FILLER_45_1787 ();
 sg13g2_decap_4 FILLER_45_1799 ();
 sg13g2_decap_8 FILLER_45_1813 ();
 sg13g2_decap_8 FILLER_45_1820 ();
 sg13g2_fill_2 FILLER_45_1837 ();
 sg13g2_fill_1 FILLER_45_1839 ();
 sg13g2_decap_4 FILLER_45_1850 ();
 sg13g2_fill_2 FILLER_45_1854 ();
 sg13g2_decap_8 FILLER_45_1882 ();
 sg13g2_decap_8 FILLER_45_1889 ();
 sg13g2_fill_2 FILLER_45_1896 ();
 sg13g2_fill_1 FILLER_45_1898 ();
 sg13g2_fill_2 FILLER_45_1922 ();
 sg13g2_fill_1 FILLER_45_1924 ();
 sg13g2_decap_4 FILLER_45_1937 ();
 sg13g2_fill_2 FILLER_45_1941 ();
 sg13g2_fill_1 FILLER_45_1969 ();
 sg13g2_decap_8 FILLER_45_1996 ();
 sg13g2_decap_8 FILLER_45_2003 ();
 sg13g2_decap_8 FILLER_45_2010 ();
 sg13g2_decap_8 FILLER_45_2027 ();
 sg13g2_decap_8 FILLER_45_2034 ();
 sg13g2_fill_1 FILLER_45_2041 ();
 sg13g2_fill_2 FILLER_45_2068 ();
 sg13g2_fill_1 FILLER_45_2070 ();
 sg13g2_decap_8 FILLER_45_2077 ();
 sg13g2_decap_8 FILLER_45_2084 ();
 sg13g2_fill_1 FILLER_45_2091 ();
 sg13g2_decap_8 FILLER_45_2118 ();
 sg13g2_decap_8 FILLER_45_2125 ();
 sg13g2_decap_4 FILLER_45_2132 ();
 sg13g2_fill_2 FILLER_45_2136 ();
 sg13g2_decap_4 FILLER_45_2190 ();
 sg13g2_fill_1 FILLER_45_2194 ();
 sg13g2_decap_8 FILLER_45_2224 ();
 sg13g2_decap_8 FILLER_45_2231 ();
 sg13g2_decap_8 FILLER_45_2238 ();
 sg13g2_fill_1 FILLER_45_2245 ();
 sg13g2_fill_1 FILLER_45_2251 ();
 sg13g2_fill_1 FILLER_45_2277 ();
 sg13g2_fill_2 FILLER_45_2291 ();
 sg13g2_fill_1 FILLER_45_2308 ();
 sg13g2_fill_2 FILLER_45_2340 ();
 sg13g2_fill_1 FILLER_45_2342 ();
 sg13g2_decap_8 FILLER_45_2363 ();
 sg13g2_decap_8 FILLER_45_2370 ();
 sg13g2_fill_2 FILLER_45_2377 ();
 sg13g2_fill_1 FILLER_45_2379 ();
 sg13g2_fill_2 FILLER_45_2410 ();
 sg13g2_decap_8 FILLER_45_2425 ();
 sg13g2_decap_8 FILLER_45_2432 ();
 sg13g2_decap_8 FILLER_45_2439 ();
 sg13g2_fill_2 FILLER_45_2446 ();
 sg13g2_decap_8 FILLER_45_2480 ();
 sg13g2_decap_8 FILLER_45_2487 ();
 sg13g2_decap_8 FILLER_45_2494 ();
 sg13g2_decap_8 FILLER_45_2522 ();
 sg13g2_decap_8 FILLER_45_2529 ();
 sg13g2_decap_8 FILLER_45_2536 ();
 sg13g2_decap_8 FILLER_45_2543 ();
 sg13g2_decap_8 FILLER_45_2550 ();
 sg13g2_decap_8 FILLER_45_2557 ();
 sg13g2_decap_8 FILLER_45_2564 ();
 sg13g2_decap_8 FILLER_45_2571 ();
 sg13g2_decap_4 FILLER_45_2578 ();
 sg13g2_fill_1 FILLER_45_2587 ();
 sg13g2_decap_8 FILLER_45_2606 ();
 sg13g2_decap_8 FILLER_45_2613 ();
 sg13g2_decap_8 FILLER_45_2620 ();
 sg13g2_decap_8 FILLER_45_2627 ();
 sg13g2_decap_8 FILLER_45_2634 ();
 sg13g2_decap_8 FILLER_45_2641 ();
 sg13g2_decap_8 FILLER_45_2684 ();
 sg13g2_decap_8 FILLER_45_2691 ();
 sg13g2_decap_8 FILLER_45_2698 ();
 sg13g2_decap_8 FILLER_45_2705 ();
 sg13g2_decap_8 FILLER_45_2712 ();
 sg13g2_fill_2 FILLER_45_2719 ();
 sg13g2_fill_1 FILLER_45_2721 ();
 sg13g2_decap_8 FILLER_45_2726 ();
 sg13g2_decap_8 FILLER_45_2733 ();
 sg13g2_decap_8 FILLER_45_2740 ();
 sg13g2_decap_8 FILLER_45_2747 ();
 sg13g2_decap_8 FILLER_45_2754 ();
 sg13g2_decap_8 FILLER_45_2761 ();
 sg13g2_decap_8 FILLER_45_2768 ();
 sg13g2_decap_8 FILLER_45_2794 ();
 sg13g2_decap_8 FILLER_45_2801 ();
 sg13g2_decap_8 FILLER_45_2808 ();
 sg13g2_decap_8 FILLER_45_2850 ();
 sg13g2_decap_8 FILLER_45_2857 ();
 sg13g2_decap_8 FILLER_45_2864 ();
 sg13g2_decap_4 FILLER_45_2871 ();
 sg13g2_decap_8 FILLER_45_2901 ();
 sg13g2_decap_8 FILLER_45_2908 ();
 sg13g2_decap_8 FILLER_45_2915 ();
 sg13g2_decap_8 FILLER_45_2922 ();
 sg13g2_decap_4 FILLER_45_2929 ();
 sg13g2_fill_2 FILLER_45_2933 ();
 sg13g2_decap_8 FILLER_45_2943 ();
 sg13g2_decap_8 FILLER_45_2950 ();
 sg13g2_decap_8 FILLER_45_2957 ();
 sg13g2_decap_8 FILLER_45_2974 ();
 sg13g2_decap_8 FILLER_45_2981 ();
 sg13g2_decap_8 FILLER_45_2988 ();
 sg13g2_decap_4 FILLER_45_2995 ();
 sg13g2_fill_2 FILLER_45_2999 ();
 sg13g2_decap_8 FILLER_45_3006 ();
 sg13g2_fill_2 FILLER_45_3013 ();
 sg13g2_fill_1 FILLER_45_3015 ();
 sg13g2_decap_8 FILLER_45_3060 ();
 sg13g2_decap_8 FILLER_45_3067 ();
 sg13g2_decap_8 FILLER_45_3074 ();
 sg13g2_fill_2 FILLER_45_3081 ();
 sg13g2_fill_1 FILLER_45_3083 ();
 sg13g2_decap_8 FILLER_45_3099 ();
 sg13g2_decap_8 FILLER_45_3106 ();
 sg13g2_decap_8 FILLER_45_3113 ();
 sg13g2_decap_8 FILLER_45_3120 ();
 sg13g2_decap_8 FILLER_45_3127 ();
 sg13g2_decap_4 FILLER_45_3134 ();
 sg13g2_fill_1 FILLER_45_3138 ();
 sg13g2_decap_8 FILLER_45_3165 ();
 sg13g2_decap_4 FILLER_45_3172 ();
 sg13g2_fill_2 FILLER_45_3176 ();
 sg13g2_decap_8 FILLER_45_3186 ();
 sg13g2_decap_4 FILLER_45_3198 ();
 sg13g2_fill_2 FILLER_45_3202 ();
 sg13g2_decap_8 FILLER_45_3207 ();
 sg13g2_decap_8 FILLER_45_3214 ();
 sg13g2_decap_8 FILLER_45_3221 ();
 sg13g2_decap_4 FILLER_45_3228 ();
 sg13g2_fill_2 FILLER_45_3232 ();
 sg13g2_decap_8 FILLER_45_3242 ();
 sg13g2_fill_2 FILLER_45_3249 ();
 sg13g2_decap_8 FILLER_45_3287 ();
 sg13g2_decap_8 FILLER_45_3294 ();
 sg13g2_decap_8 FILLER_45_3301 ();
 sg13g2_decap_8 FILLER_45_3308 ();
 sg13g2_decap_8 FILLER_45_3315 ();
 sg13g2_decap_8 FILLER_45_3322 ();
 sg13g2_decap_8 FILLER_45_3329 ();
 sg13g2_decap_8 FILLER_45_3336 ();
 sg13g2_decap_8 FILLER_45_3343 ();
 sg13g2_decap_8 FILLER_45_3350 ();
 sg13g2_decap_8 FILLER_45_3357 ();
 sg13g2_decap_8 FILLER_45_3364 ();
 sg13g2_fill_2 FILLER_45_3371 ();
 sg13g2_decap_8 FILLER_45_3383 ();
 sg13g2_decap_8 FILLER_45_3390 ();
 sg13g2_decap_8 FILLER_45_3397 ();
 sg13g2_decap_8 FILLER_45_3404 ();
 sg13g2_decap_8 FILLER_45_3411 ();
 sg13g2_decap_8 FILLER_45_3418 ();
 sg13g2_decap_8 FILLER_45_3425 ();
 sg13g2_decap_8 FILLER_45_3432 ();
 sg13g2_fill_2 FILLER_45_3439 ();
 sg13g2_decap_8 FILLER_45_3456 ();
 sg13g2_decap_8 FILLER_45_3463 ();
 sg13g2_decap_4 FILLER_45_3470 ();
 sg13g2_fill_1 FILLER_45_3474 ();
 sg13g2_decap_8 FILLER_45_3495 ();
 sg13g2_decap_8 FILLER_45_3502 ();
 sg13g2_decap_8 FILLER_45_3509 ();
 sg13g2_fill_2 FILLER_45_3516 ();
 sg13g2_decap_4 FILLER_45_3528 ();
 sg13g2_decap_8 FILLER_45_3558 ();
 sg13g2_decap_8 FILLER_45_3565 ();
 sg13g2_decap_8 FILLER_45_3572 ();
 sg13g2_fill_1 FILLER_45_3579 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_fill_1 FILLER_46_7 ();
 sg13g2_fill_1 FILLER_46_58 ();
 sg13g2_fill_2 FILLER_46_64 ();
 sg13g2_fill_1 FILLER_46_75 ();
 sg13g2_decap_8 FILLER_46_83 ();
 sg13g2_decap_8 FILLER_46_90 ();
 sg13g2_decap_8 FILLER_46_97 ();
 sg13g2_decap_8 FILLER_46_104 ();
 sg13g2_decap_8 FILLER_46_111 ();
 sg13g2_decap_8 FILLER_46_118 ();
 sg13g2_decap_8 FILLER_46_125 ();
 sg13g2_decap_8 FILLER_46_132 ();
 sg13g2_decap_8 FILLER_46_139 ();
 sg13g2_decap_8 FILLER_46_146 ();
 sg13g2_decap_8 FILLER_46_153 ();
 sg13g2_decap_8 FILLER_46_160 ();
 sg13g2_decap_8 FILLER_46_167 ();
 sg13g2_decap_8 FILLER_46_174 ();
 sg13g2_decap_4 FILLER_46_181 ();
 sg13g2_fill_2 FILLER_46_185 ();
 sg13g2_decap_4 FILLER_46_213 ();
 sg13g2_decap_4 FILLER_46_222 ();
 sg13g2_fill_1 FILLER_46_235 ();
 sg13g2_fill_2 FILLER_46_241 ();
 sg13g2_decap_8 FILLER_46_248 ();
 sg13g2_decap_8 FILLER_46_255 ();
 sg13g2_decap_4 FILLER_46_262 ();
 sg13g2_fill_2 FILLER_46_282 ();
 sg13g2_fill_2 FILLER_46_295 ();
 sg13g2_fill_1 FILLER_46_297 ();
 sg13g2_decap_8 FILLER_46_305 ();
 sg13g2_decap_8 FILLER_46_312 ();
 sg13g2_decap_8 FILLER_46_319 ();
 sg13g2_decap_8 FILLER_46_326 ();
 sg13g2_decap_8 FILLER_46_333 ();
 sg13g2_decap_8 FILLER_46_340 ();
 sg13g2_decap_8 FILLER_46_347 ();
 sg13g2_decap_8 FILLER_46_354 ();
 sg13g2_decap_8 FILLER_46_361 ();
 sg13g2_decap_4 FILLER_46_368 ();
 sg13g2_fill_2 FILLER_46_372 ();
 sg13g2_fill_1 FILLER_46_386 ();
 sg13g2_decap_8 FILLER_46_401 ();
 sg13g2_decap_8 FILLER_46_408 ();
 sg13g2_decap_8 FILLER_46_415 ();
 sg13g2_decap_4 FILLER_46_422 ();
 sg13g2_fill_1 FILLER_46_426 ();
 sg13g2_decap_4 FILLER_46_439 ();
 sg13g2_fill_2 FILLER_46_443 ();
 sg13g2_fill_2 FILLER_46_456 ();
 sg13g2_fill_1 FILLER_46_458 ();
 sg13g2_decap_8 FILLER_46_465 ();
 sg13g2_decap_8 FILLER_46_472 ();
 sg13g2_decap_8 FILLER_46_479 ();
 sg13g2_decap_4 FILLER_46_486 ();
 sg13g2_fill_1 FILLER_46_490 ();
 sg13g2_decap_8 FILLER_46_503 ();
 sg13g2_decap_8 FILLER_46_510 ();
 sg13g2_decap_4 FILLER_46_517 ();
 sg13g2_decap_8 FILLER_46_547 ();
 sg13g2_decap_8 FILLER_46_554 ();
 sg13g2_decap_8 FILLER_46_561 ();
 sg13g2_decap_8 FILLER_46_583 ();
 sg13g2_decap_4 FILLER_46_590 ();
 sg13g2_fill_2 FILLER_46_603 ();
 sg13g2_fill_1 FILLER_46_605 ();
 sg13g2_decap_8 FILLER_46_614 ();
 sg13g2_decap_8 FILLER_46_668 ();
 sg13g2_fill_1 FILLER_46_675 ();
 sg13g2_decap_8 FILLER_46_685 ();
 sg13g2_decap_8 FILLER_46_692 ();
 sg13g2_decap_8 FILLER_46_699 ();
 sg13g2_fill_2 FILLER_46_706 ();
 sg13g2_decap_8 FILLER_46_714 ();
 sg13g2_decap_8 FILLER_46_721 ();
 sg13g2_decap_4 FILLER_46_728 ();
 sg13g2_fill_1 FILLER_46_732 ();
 sg13g2_decap_8 FILLER_46_753 ();
 sg13g2_fill_2 FILLER_46_764 ();
 sg13g2_fill_1 FILLER_46_774 ();
 sg13g2_decap_8 FILLER_46_801 ();
 sg13g2_decap_8 FILLER_46_808 ();
 sg13g2_decap_8 FILLER_46_815 ();
 sg13g2_decap_8 FILLER_46_822 ();
 sg13g2_decap_8 FILLER_46_829 ();
 sg13g2_decap_8 FILLER_46_836 ();
 sg13g2_decap_8 FILLER_46_843 ();
 sg13g2_decap_8 FILLER_46_850 ();
 sg13g2_decap_8 FILLER_46_857 ();
 sg13g2_decap_8 FILLER_46_864 ();
 sg13g2_decap_8 FILLER_46_897 ();
 sg13g2_decap_8 FILLER_46_904 ();
 sg13g2_decap_8 FILLER_46_911 ();
 sg13g2_decap_8 FILLER_46_918 ();
 sg13g2_fill_2 FILLER_46_925 ();
 sg13g2_decap_8 FILLER_46_945 ();
 sg13g2_decap_8 FILLER_46_952 ();
 sg13g2_decap_8 FILLER_46_959 ();
 sg13g2_fill_2 FILLER_46_966 ();
 sg13g2_decap_8 FILLER_46_976 ();
 sg13g2_decap_8 FILLER_46_983 ();
 sg13g2_decap_8 FILLER_46_995 ();
 sg13g2_decap_8 FILLER_46_1002 ();
 sg13g2_decap_8 FILLER_46_1014 ();
 sg13g2_decap_8 FILLER_46_1038 ();
 sg13g2_decap_8 FILLER_46_1045 ();
 sg13g2_decap_8 FILLER_46_1052 ();
 sg13g2_decap_8 FILLER_46_1059 ();
 sg13g2_decap_8 FILLER_46_1066 ();
 sg13g2_fill_2 FILLER_46_1073 ();
 sg13g2_fill_1 FILLER_46_1075 ();
 sg13g2_decap_8 FILLER_46_1098 ();
 sg13g2_decap_8 FILLER_46_1105 ();
 sg13g2_decap_4 FILLER_46_1112 ();
 sg13g2_fill_1 FILLER_46_1116 ();
 sg13g2_decap_4 FILLER_46_1126 ();
 sg13g2_fill_1 FILLER_46_1130 ();
 sg13g2_decap_8 FILLER_46_1140 ();
 sg13g2_decap_8 FILLER_46_1147 ();
 sg13g2_decap_8 FILLER_46_1154 ();
 sg13g2_fill_2 FILLER_46_1161 ();
 sg13g2_fill_2 FILLER_46_1172 ();
 sg13g2_fill_1 FILLER_46_1183 ();
 sg13g2_fill_2 FILLER_46_1194 ();
 sg13g2_decap_8 FILLER_46_1204 ();
 sg13g2_decap_4 FILLER_46_1211 ();
 sg13g2_fill_1 FILLER_46_1215 ();
 sg13g2_decap_8 FILLER_46_1246 ();
 sg13g2_decap_8 FILLER_46_1253 ();
 sg13g2_decap_8 FILLER_46_1260 ();
 sg13g2_decap_8 FILLER_46_1267 ();
 sg13g2_decap_8 FILLER_46_1274 ();
 sg13g2_decap_8 FILLER_46_1307 ();
 sg13g2_decap_8 FILLER_46_1314 ();
 sg13g2_decap_8 FILLER_46_1321 ();
 sg13g2_decap_8 FILLER_46_1328 ();
 sg13g2_decap_8 FILLER_46_1335 ();
 sg13g2_decap_4 FILLER_46_1342 ();
 sg13g2_decap_8 FILLER_46_1367 ();
 sg13g2_decap_8 FILLER_46_1374 ();
 sg13g2_decap_8 FILLER_46_1381 ();
 sg13g2_decap_8 FILLER_46_1388 ();
 sg13g2_decap_8 FILLER_46_1395 ();
 sg13g2_fill_1 FILLER_46_1402 ();
 sg13g2_decap_8 FILLER_46_1429 ();
 sg13g2_fill_1 FILLER_46_1436 ();
 sg13g2_decap_4 FILLER_46_1440 ();
 sg13g2_fill_2 FILLER_46_1444 ();
 sg13g2_decap_8 FILLER_46_1472 ();
 sg13g2_decap_8 FILLER_46_1479 ();
 sg13g2_decap_8 FILLER_46_1486 ();
 sg13g2_decap_8 FILLER_46_1493 ();
 sg13g2_decap_8 FILLER_46_1500 ();
 sg13g2_fill_2 FILLER_46_1507 ();
 sg13g2_fill_1 FILLER_46_1509 ();
 sg13g2_decap_8 FILLER_46_1520 ();
 sg13g2_fill_2 FILLER_46_1527 ();
 sg13g2_fill_1 FILLER_46_1529 ();
 sg13g2_decap_8 FILLER_46_1543 ();
 sg13g2_decap_8 FILLER_46_1550 ();
 sg13g2_decap_8 FILLER_46_1583 ();
 sg13g2_decap_8 FILLER_46_1590 ();
 sg13g2_decap_8 FILLER_46_1597 ();
 sg13g2_decap_8 FILLER_46_1604 ();
 sg13g2_decap_8 FILLER_46_1611 ();
 sg13g2_decap_8 FILLER_46_1618 ();
 sg13g2_fill_1 FILLER_46_1625 ();
 sg13g2_decap_4 FILLER_46_1632 ();
 sg13g2_fill_1 FILLER_46_1636 ();
 sg13g2_decap_8 FILLER_46_1643 ();
 sg13g2_decap_8 FILLER_46_1650 ();
 sg13g2_decap_8 FILLER_46_1657 ();
 sg13g2_decap_8 FILLER_46_1664 ();
 sg13g2_decap_8 FILLER_46_1671 ();
 sg13g2_decap_8 FILLER_46_1678 ();
 sg13g2_decap_8 FILLER_46_1721 ();
 sg13g2_decap_8 FILLER_46_1728 ();
 sg13g2_decap_8 FILLER_46_1735 ();
 sg13g2_decap_8 FILLER_46_1742 ();
 sg13g2_decap_8 FILLER_46_1749 ();
 sg13g2_fill_1 FILLER_46_1756 ();
 sg13g2_decap_8 FILLER_46_1783 ();
 sg13g2_decap_8 FILLER_46_1790 ();
 sg13g2_decap_8 FILLER_46_1797 ();
 sg13g2_fill_2 FILLER_46_1804 ();
 sg13g2_fill_1 FILLER_46_1806 ();
 sg13g2_fill_2 FILLER_46_1839 ();
 sg13g2_decap_8 FILLER_46_1867 ();
 sg13g2_decap_4 FILLER_46_1874 ();
 sg13g2_fill_2 FILLER_46_1878 ();
 sg13g2_fill_2 FILLER_46_1888 ();
 sg13g2_fill_2 FILLER_46_1905 ();
 sg13g2_fill_1 FILLER_46_1907 ();
 sg13g2_decap_8 FILLER_46_1926 ();
 sg13g2_decap_8 FILLER_46_1933 ();
 sg13g2_decap_8 FILLER_46_1940 ();
 sg13g2_decap_8 FILLER_46_1947 ();
 sg13g2_decap_8 FILLER_46_1954 ();
 sg13g2_decap_8 FILLER_46_1961 ();
 sg13g2_decap_8 FILLER_46_1968 ();
 sg13g2_decap_8 FILLER_46_1975 ();
 sg13g2_fill_1 FILLER_46_1982 ();
 sg13g2_decap_8 FILLER_46_1997 ();
 sg13g2_decap_8 FILLER_46_2044 ();
 sg13g2_decap_8 FILLER_46_2051 ();
 sg13g2_decap_8 FILLER_46_2058 ();
 sg13g2_decap_8 FILLER_46_2065 ();
 sg13g2_decap_8 FILLER_46_2072 ();
 sg13g2_decap_8 FILLER_46_2079 ();
 sg13g2_decap_4 FILLER_46_2086 ();
 sg13g2_decap_4 FILLER_46_2096 ();
 sg13g2_fill_1 FILLER_46_2100 ();
 sg13g2_decap_8 FILLER_46_2107 ();
 sg13g2_decap_8 FILLER_46_2114 ();
 sg13g2_decap_8 FILLER_46_2121 ();
 sg13g2_decap_8 FILLER_46_2128 ();
 sg13g2_decap_8 FILLER_46_2135 ();
 sg13g2_fill_1 FILLER_46_2159 ();
 sg13g2_decap_8 FILLER_46_2166 ();
 sg13g2_decap_8 FILLER_46_2173 ();
 sg13g2_decap_8 FILLER_46_2180 ();
 sg13g2_decap_8 FILLER_46_2187 ();
 sg13g2_fill_1 FILLER_46_2194 ();
 sg13g2_decap_4 FILLER_46_2198 ();
 sg13g2_fill_1 FILLER_46_2202 ();
 sg13g2_decap_8 FILLER_46_2217 ();
 sg13g2_decap_8 FILLER_46_2224 ();
 sg13g2_decap_8 FILLER_46_2231 ();
 sg13g2_decap_8 FILLER_46_2238 ();
 sg13g2_decap_8 FILLER_46_2245 ();
 sg13g2_fill_1 FILLER_46_2252 ();
 sg13g2_fill_2 FILLER_46_2258 ();
 sg13g2_fill_1 FILLER_46_2260 ();
 sg13g2_decap_8 FILLER_46_2273 ();
 sg13g2_decap_8 FILLER_46_2280 ();
 sg13g2_decap_4 FILLER_46_2287 ();
 sg13g2_fill_2 FILLER_46_2291 ();
 sg13g2_decap_8 FILLER_46_2296 ();
 sg13g2_decap_8 FILLER_46_2303 ();
 sg13g2_decap_8 FILLER_46_2310 ();
 sg13g2_decap_8 FILLER_46_2317 ();
 sg13g2_decap_4 FILLER_46_2324 ();
 sg13g2_fill_1 FILLER_46_2341 ();
 sg13g2_decap_8 FILLER_46_2357 ();
 sg13g2_decap_8 FILLER_46_2364 ();
 sg13g2_decap_8 FILLER_46_2371 ();
 sg13g2_decap_8 FILLER_46_2378 ();
 sg13g2_fill_2 FILLER_46_2385 ();
 sg13g2_fill_1 FILLER_46_2387 ();
 sg13g2_fill_2 FILLER_46_2404 ();
 sg13g2_decap_8 FILLER_46_2417 ();
 sg13g2_decap_8 FILLER_46_2424 ();
 sg13g2_decap_8 FILLER_46_2431 ();
 sg13g2_decap_8 FILLER_46_2438 ();
 sg13g2_decap_8 FILLER_46_2445 ();
 sg13g2_decap_8 FILLER_46_2452 ();
 sg13g2_decap_8 FILLER_46_2459 ();
 sg13g2_decap_8 FILLER_46_2466 ();
 sg13g2_decap_4 FILLER_46_2473 ();
 sg13g2_decap_8 FILLER_46_2497 ();
 sg13g2_fill_2 FILLER_46_2513 ();
 sg13g2_decap_8 FILLER_46_2541 ();
 sg13g2_fill_1 FILLER_46_2548 ();
 sg13g2_fill_1 FILLER_46_2559 ();
 sg13g2_decap_8 FILLER_46_2571 ();
 sg13g2_decap_8 FILLER_46_2578 ();
 sg13g2_decap_4 FILLER_46_2585 ();
 sg13g2_fill_1 FILLER_46_2589 ();
 sg13g2_decap_8 FILLER_46_2624 ();
 sg13g2_fill_1 FILLER_46_2631 ();
 sg13g2_decap_8 FILLER_46_2649 ();
 sg13g2_decap_8 FILLER_46_2656 ();
 sg13g2_fill_2 FILLER_46_2663 ();
 sg13g2_fill_1 FILLER_46_2665 ();
 sg13g2_decap_8 FILLER_46_2674 ();
 sg13g2_decap_8 FILLER_46_2681 ();
 sg13g2_decap_8 FILLER_46_2688 ();
 sg13g2_decap_8 FILLER_46_2695 ();
 sg13g2_decap_8 FILLER_46_2702 ();
 sg13g2_decap_8 FILLER_46_2719 ();
 sg13g2_decap_4 FILLER_46_2726 ();
 sg13g2_decap_8 FILLER_46_2740 ();
 sg13g2_decap_8 FILLER_46_2747 ();
 sg13g2_decap_4 FILLER_46_2754 ();
 sg13g2_fill_1 FILLER_46_2758 ();
 sg13g2_fill_2 FILLER_46_2794 ();
 sg13g2_decap_8 FILLER_46_2800 ();
 sg13g2_decap_4 FILLER_46_2807 ();
 sg13g2_fill_1 FILLER_46_2811 ();
 sg13g2_fill_2 FILLER_46_2820 ();
 sg13g2_decap_8 FILLER_46_2848 ();
 sg13g2_decap_8 FILLER_46_2855 ();
 sg13g2_decap_4 FILLER_46_2862 ();
 sg13g2_fill_2 FILLER_46_2866 ();
 sg13g2_decap_8 FILLER_46_2894 ();
 sg13g2_decap_8 FILLER_46_2901 ();
 sg13g2_decap_8 FILLER_46_2908 ();
 sg13g2_decap_8 FILLER_46_2915 ();
 sg13g2_decap_8 FILLER_46_2922 ();
 sg13g2_decap_8 FILLER_46_2929 ();
 sg13g2_decap_8 FILLER_46_2936 ();
 sg13g2_decap_8 FILLER_46_2943 ();
 sg13g2_decap_8 FILLER_46_2950 ();
 sg13g2_decap_8 FILLER_46_2957 ();
 sg13g2_decap_8 FILLER_46_2964 ();
 sg13g2_decap_4 FILLER_46_2971 ();
 sg13g2_decap_8 FILLER_46_2985 ();
 sg13g2_decap_8 FILLER_46_2992 ();
 sg13g2_decap_8 FILLER_46_2999 ();
 sg13g2_decap_8 FILLER_46_3006 ();
 sg13g2_decap_8 FILLER_46_3013 ();
 sg13g2_decap_8 FILLER_46_3020 ();
 sg13g2_decap_8 FILLER_46_3027 ();
 sg13g2_decap_8 FILLER_46_3045 ();
 sg13g2_decap_8 FILLER_46_3052 ();
 sg13g2_decap_8 FILLER_46_3059 ();
 sg13g2_decap_8 FILLER_46_3066 ();
 sg13g2_decap_8 FILLER_46_3073 ();
 sg13g2_decap_4 FILLER_46_3080 ();
 sg13g2_fill_2 FILLER_46_3084 ();
 sg13g2_decap_8 FILLER_46_3125 ();
 sg13g2_decap_8 FILLER_46_3132 ();
 sg13g2_decap_8 FILLER_46_3139 ();
 sg13g2_decap_8 FILLER_46_3150 ();
 sg13g2_decap_8 FILLER_46_3166 ();
 sg13g2_decap_8 FILLER_46_3173 ();
 sg13g2_decap_8 FILLER_46_3180 ();
 sg13g2_decap_4 FILLER_46_3187 ();
 sg13g2_fill_1 FILLER_46_3191 ();
 sg13g2_decap_8 FILLER_46_3218 ();
 sg13g2_decap_8 FILLER_46_3225 ();
 sg13g2_decap_8 FILLER_46_3232 ();
 sg13g2_decap_8 FILLER_46_3239 ();
 sg13g2_fill_2 FILLER_46_3246 ();
 sg13g2_decap_8 FILLER_46_3274 ();
 sg13g2_decap_8 FILLER_46_3281 ();
 sg13g2_decap_4 FILLER_46_3288 ();
 sg13g2_fill_2 FILLER_46_3292 ();
 sg13g2_decap_8 FILLER_46_3300 ();
 sg13g2_decap_4 FILLER_46_3307 ();
 sg13g2_fill_1 FILLER_46_3311 ();
 sg13g2_decap_8 FILLER_46_3322 ();
 sg13g2_decap_8 FILLER_46_3329 ();
 sg13g2_decap_8 FILLER_46_3336 ();
 sg13g2_decap_8 FILLER_46_3343 ();
 sg13g2_decap_8 FILLER_46_3350 ();
 sg13g2_decap_8 FILLER_46_3357 ();
 sg13g2_decap_8 FILLER_46_3364 ();
 sg13g2_decap_8 FILLER_46_3371 ();
 sg13g2_decap_8 FILLER_46_3378 ();
 sg13g2_decap_8 FILLER_46_3385 ();
 sg13g2_decap_8 FILLER_46_3392 ();
 sg13g2_fill_1 FILLER_46_3399 ();
 sg13g2_decap_4 FILLER_46_3405 ();
 sg13g2_decap_8 FILLER_46_3424 ();
 sg13g2_decap_4 FILLER_46_3431 ();
 sg13g2_decap_8 FILLER_46_3455 ();
 sg13g2_decap_8 FILLER_46_3462 ();
 sg13g2_decap_8 FILLER_46_3469 ();
 sg13g2_decap_4 FILLER_46_3476 ();
 sg13g2_fill_1 FILLER_46_3480 ();
 sg13g2_fill_1 FILLER_46_3501 ();
 sg13g2_decap_8 FILLER_46_3507 ();
 sg13g2_decap_8 FILLER_46_3514 ();
 sg13g2_decap_4 FILLER_46_3521 ();
 sg13g2_fill_2 FILLER_46_3530 ();
 sg13g2_decap_8 FILLER_46_3552 ();
 sg13g2_decap_8 FILLER_46_3559 ();
 sg13g2_decap_8 FILLER_46_3566 ();
 sg13g2_decap_8 FILLER_46_3573 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_7 ();
 sg13g2_fill_2 FILLER_47_14 ();
 sg13g2_fill_1 FILLER_47_16 ();
 sg13g2_decap_4 FILLER_47_26 ();
 sg13g2_fill_2 FILLER_47_30 ();
 sg13g2_decap_8 FILLER_47_37 ();
 sg13g2_decap_8 FILLER_47_44 ();
 sg13g2_fill_2 FILLER_47_51 ();
 sg13g2_decap_8 FILLER_47_100 ();
 sg13g2_decap_8 FILLER_47_107 ();
 sg13g2_decap_8 FILLER_47_114 ();
 sg13g2_decap_8 FILLER_47_121 ();
 sg13g2_decap_8 FILLER_47_128 ();
 sg13g2_fill_2 FILLER_47_135 ();
 sg13g2_decap_4 FILLER_47_155 ();
 sg13g2_fill_2 FILLER_47_159 ();
 sg13g2_decap_8 FILLER_47_164 ();
 sg13g2_decap_4 FILLER_47_171 ();
 sg13g2_decap_8 FILLER_47_180 ();
 sg13g2_fill_2 FILLER_47_187 ();
 sg13g2_fill_2 FILLER_47_200 ();
 sg13g2_fill_1 FILLER_47_252 ();
 sg13g2_fill_2 FILLER_47_261 ();
 sg13g2_fill_1 FILLER_47_292 ();
 sg13g2_decap_8 FILLER_47_314 ();
 sg13g2_fill_1 FILLER_47_326 ();
 sg13g2_decap_4 FILLER_47_335 ();
 sg13g2_decap_8 FILLER_47_350 ();
 sg13g2_decap_8 FILLER_47_357 ();
 sg13g2_decap_8 FILLER_47_364 ();
 sg13g2_decap_8 FILLER_47_371 ();
 sg13g2_decap_8 FILLER_47_378 ();
 sg13g2_decap_8 FILLER_47_385 ();
 sg13g2_decap_4 FILLER_47_392 ();
 sg13g2_fill_1 FILLER_47_396 ();
 sg13g2_decap_8 FILLER_47_403 ();
 sg13g2_decap_8 FILLER_47_410 ();
 sg13g2_fill_2 FILLER_47_417 ();
 sg13g2_fill_1 FILLER_47_419 ();
 sg13g2_fill_2 FILLER_47_426 ();
 sg13g2_decap_4 FILLER_47_434 ();
 sg13g2_fill_1 FILLER_47_438 ();
 sg13g2_decap_8 FILLER_47_450 ();
 sg13g2_decap_8 FILLER_47_457 ();
 sg13g2_decap_8 FILLER_47_470 ();
 sg13g2_fill_2 FILLER_47_477 ();
 sg13g2_decap_8 FILLER_47_486 ();
 sg13g2_fill_2 FILLER_47_493 ();
 sg13g2_decap_4 FILLER_47_515 ();
 sg13g2_fill_2 FILLER_47_519 ();
 sg13g2_decap_8 FILLER_47_526 ();
 sg13g2_decap_8 FILLER_47_533 ();
 sg13g2_decap_8 FILLER_47_540 ();
 sg13g2_decap_8 FILLER_47_547 ();
 sg13g2_decap_8 FILLER_47_554 ();
 sg13g2_decap_8 FILLER_47_561 ();
 sg13g2_decap_8 FILLER_47_568 ();
 sg13g2_decap_8 FILLER_47_575 ();
 sg13g2_fill_2 FILLER_47_582 ();
 sg13g2_decap_8 FILLER_47_589 ();
 sg13g2_decap_8 FILLER_47_596 ();
 sg13g2_decap_8 FILLER_47_603 ();
 sg13g2_fill_2 FILLER_47_610 ();
 sg13g2_fill_1 FILLER_47_612 ();
 sg13g2_decap_8 FILLER_47_620 ();
 sg13g2_decap_8 FILLER_47_627 ();
 sg13g2_decap_4 FILLER_47_634 ();
 sg13g2_decap_8 FILLER_47_657 ();
 sg13g2_fill_2 FILLER_47_670 ();
 sg13g2_fill_1 FILLER_47_672 ();
 sg13g2_decap_8 FILLER_47_682 ();
 sg13g2_decap_8 FILLER_47_689 ();
 sg13g2_decap_8 FILLER_47_696 ();
 sg13g2_decap_8 FILLER_47_703 ();
 sg13g2_decap_4 FILLER_47_710 ();
 sg13g2_fill_1 FILLER_47_714 ();
 sg13g2_fill_1 FILLER_47_725 ();
 sg13g2_decap_8 FILLER_47_739 ();
 sg13g2_fill_2 FILLER_47_751 ();
 sg13g2_fill_1 FILLER_47_753 ();
 sg13g2_decap_8 FILLER_47_767 ();
 sg13g2_decap_8 FILLER_47_774 ();
 sg13g2_decap_8 FILLER_47_781 ();
 sg13g2_decap_8 FILLER_47_788 ();
 sg13g2_decap_8 FILLER_47_795 ();
 sg13g2_decap_8 FILLER_47_802 ();
 sg13g2_decap_8 FILLER_47_809 ();
 sg13g2_decap_8 FILLER_47_816 ();
 sg13g2_decap_8 FILLER_47_823 ();
 sg13g2_decap_8 FILLER_47_830 ();
 sg13g2_decap_4 FILLER_47_837 ();
 sg13g2_fill_2 FILLER_47_841 ();
 sg13g2_decap_8 FILLER_47_877 ();
 sg13g2_decap_8 FILLER_47_884 ();
 sg13g2_fill_2 FILLER_47_891 ();
 sg13g2_decap_8 FILLER_47_898 ();
 sg13g2_decap_8 FILLER_47_905 ();
 sg13g2_decap_4 FILLER_47_912 ();
 sg13g2_fill_2 FILLER_47_916 ();
 sg13g2_decap_8 FILLER_47_941 ();
 sg13g2_decap_8 FILLER_47_948 ();
 sg13g2_decap_8 FILLER_47_955 ();
 sg13g2_decap_8 FILLER_47_962 ();
 sg13g2_decap_8 FILLER_47_969 ();
 sg13g2_decap_8 FILLER_47_976 ();
 sg13g2_fill_1 FILLER_47_983 ();
 sg13g2_fill_2 FILLER_47_1005 ();
 sg13g2_decap_8 FILLER_47_1015 ();
 sg13g2_decap_8 FILLER_47_1022 ();
 sg13g2_decap_8 FILLER_47_1029 ();
 sg13g2_decap_8 FILLER_47_1036 ();
 sg13g2_decap_8 FILLER_47_1043 ();
 sg13g2_decap_8 FILLER_47_1050 ();
 sg13g2_decap_4 FILLER_47_1057 ();
 sg13g2_decap_8 FILLER_47_1074 ();
 sg13g2_decap_8 FILLER_47_1081 ();
 sg13g2_decap_4 FILLER_47_1088 ();
 sg13g2_fill_1 FILLER_47_1092 ();
 sg13g2_decap_8 FILLER_47_1098 ();
 sg13g2_decap_8 FILLER_47_1105 ();
 sg13g2_decap_8 FILLER_47_1112 ();
 sg13g2_decap_8 FILLER_47_1119 ();
 sg13g2_decap_8 FILLER_47_1126 ();
 sg13g2_decap_4 FILLER_47_1133 ();
 sg13g2_fill_2 FILLER_47_1137 ();
 sg13g2_decap_8 FILLER_47_1203 ();
 sg13g2_decap_8 FILLER_47_1210 ();
 sg13g2_decap_4 FILLER_47_1217 ();
 sg13g2_decap_8 FILLER_47_1226 ();
 sg13g2_decap_8 FILLER_47_1242 ();
 sg13g2_decap_8 FILLER_47_1249 ();
 sg13g2_decap_8 FILLER_47_1256 ();
 sg13g2_decap_8 FILLER_47_1263 ();
 sg13g2_decap_8 FILLER_47_1270 ();
 sg13g2_decap_8 FILLER_47_1277 ();
 sg13g2_fill_2 FILLER_47_1284 ();
 sg13g2_decap_8 FILLER_47_1296 ();
 sg13g2_decap_8 FILLER_47_1303 ();
 sg13g2_decap_8 FILLER_47_1310 ();
 sg13g2_decap_8 FILLER_47_1317 ();
 sg13g2_decap_8 FILLER_47_1324 ();
 sg13g2_decap_8 FILLER_47_1331 ();
 sg13g2_decap_8 FILLER_47_1338 ();
 sg13g2_decap_8 FILLER_47_1345 ();
 sg13g2_decap_4 FILLER_47_1352 ();
 sg13g2_decap_8 FILLER_47_1366 ();
 sg13g2_decap_8 FILLER_47_1373 ();
 sg13g2_decap_8 FILLER_47_1380 ();
 sg13g2_decap_8 FILLER_47_1387 ();
 sg13g2_fill_1 FILLER_47_1394 ();
 sg13g2_decap_8 FILLER_47_1431 ();
 sg13g2_decap_8 FILLER_47_1438 ();
 sg13g2_decap_8 FILLER_47_1445 ();
 sg13g2_decap_8 FILLER_47_1452 ();
 sg13g2_decap_8 FILLER_47_1459 ();
 sg13g2_decap_8 FILLER_47_1466 ();
 sg13g2_decap_8 FILLER_47_1473 ();
 sg13g2_decap_8 FILLER_47_1480 ();
 sg13g2_decap_4 FILLER_47_1513 ();
 sg13g2_fill_1 FILLER_47_1517 ();
 sg13g2_decap_8 FILLER_47_1544 ();
 sg13g2_decap_8 FILLER_47_1551 ();
 sg13g2_decap_4 FILLER_47_1558 ();
 sg13g2_fill_2 FILLER_47_1562 ();
 sg13g2_decap_8 FILLER_47_1574 ();
 sg13g2_fill_2 FILLER_47_1581 ();
 sg13g2_decap_8 FILLER_47_1588 ();
 sg13g2_decap_8 FILLER_47_1595 ();
 sg13g2_decap_8 FILLER_47_1602 ();
 sg13g2_decap_8 FILLER_47_1609 ();
 sg13g2_decap_8 FILLER_47_1616 ();
 sg13g2_decap_8 FILLER_47_1649 ();
 sg13g2_decap_8 FILLER_47_1656 ();
 sg13g2_decap_8 FILLER_47_1663 ();
 sg13g2_decap_8 FILLER_47_1670 ();
 sg13g2_decap_8 FILLER_47_1677 ();
 sg13g2_decap_8 FILLER_47_1684 ();
 sg13g2_decap_8 FILLER_47_1691 ();
 sg13g2_decap_8 FILLER_47_1698 ();
 sg13g2_decap_8 FILLER_47_1721 ();
 sg13g2_decap_8 FILLER_47_1728 ();
 sg13g2_decap_8 FILLER_47_1735 ();
 sg13g2_decap_8 FILLER_47_1742 ();
 sg13g2_decap_8 FILLER_47_1749 ();
 sg13g2_decap_8 FILLER_47_1756 ();
 sg13g2_decap_8 FILLER_47_1763 ();
 sg13g2_decap_8 FILLER_47_1770 ();
 sg13g2_fill_2 FILLER_47_1777 ();
 sg13g2_decap_8 FILLER_47_1787 ();
 sg13g2_decap_8 FILLER_47_1794 ();
 sg13g2_decap_8 FILLER_47_1801 ();
 sg13g2_decap_8 FILLER_47_1808 ();
 sg13g2_decap_8 FILLER_47_1815 ();
 sg13g2_decap_8 FILLER_47_1822 ();
 sg13g2_decap_8 FILLER_47_1829 ();
 sg13g2_decap_8 FILLER_47_1836 ();
 sg13g2_decap_8 FILLER_47_1843 ();
 sg13g2_decap_8 FILLER_47_1850 ();
 sg13g2_decap_8 FILLER_47_1857 ();
 sg13g2_decap_8 FILLER_47_1864 ();
 sg13g2_decap_8 FILLER_47_1871 ();
 sg13g2_fill_1 FILLER_47_1878 ();
 sg13g2_fill_1 FILLER_47_1892 ();
 sg13g2_decap_8 FILLER_47_1906 ();
 sg13g2_decap_8 FILLER_47_1913 ();
 sg13g2_fill_1 FILLER_47_1920 ();
 sg13g2_decap_8 FILLER_47_1934 ();
 sg13g2_decap_8 FILLER_47_1941 ();
 sg13g2_decap_8 FILLER_47_1948 ();
 sg13g2_decap_8 FILLER_47_1955 ();
 sg13g2_decap_8 FILLER_47_1962 ();
 sg13g2_decap_4 FILLER_47_1969 ();
 sg13g2_fill_1 FILLER_47_1983 ();
 sg13g2_decap_8 FILLER_47_2029 ();
 sg13g2_decap_8 FILLER_47_2036 ();
 sg13g2_decap_8 FILLER_47_2043 ();
 sg13g2_decap_8 FILLER_47_2050 ();
 sg13g2_decap_8 FILLER_47_2057 ();
 sg13g2_decap_8 FILLER_47_2064 ();
 sg13g2_decap_4 FILLER_47_2071 ();
 sg13g2_fill_2 FILLER_47_2075 ();
 sg13g2_decap_8 FILLER_47_2113 ();
 sg13g2_decap_8 FILLER_47_2120 ();
 sg13g2_decap_8 FILLER_47_2127 ();
 sg13g2_decap_8 FILLER_47_2134 ();
 sg13g2_decap_8 FILLER_47_2147 ();
 sg13g2_decap_8 FILLER_47_2154 ();
 sg13g2_decap_8 FILLER_47_2161 ();
 sg13g2_decap_8 FILLER_47_2168 ();
 sg13g2_decap_8 FILLER_47_2175 ();
 sg13g2_decap_8 FILLER_47_2182 ();
 sg13g2_decap_8 FILLER_47_2213 ();
 sg13g2_decap_8 FILLER_47_2220 ();
 sg13g2_decap_8 FILLER_47_2227 ();
 sg13g2_fill_2 FILLER_47_2234 ();
 sg13g2_decap_4 FILLER_47_2251 ();
 sg13g2_decap_8 FILLER_47_2261 ();
 sg13g2_decap_8 FILLER_47_2268 ();
 sg13g2_decap_8 FILLER_47_2275 ();
 sg13g2_decap_8 FILLER_47_2282 ();
 sg13g2_decap_8 FILLER_47_2289 ();
 sg13g2_decap_8 FILLER_47_2296 ();
 sg13g2_decap_8 FILLER_47_2303 ();
 sg13g2_decap_8 FILLER_47_2310 ();
 sg13g2_fill_1 FILLER_47_2317 ();
 sg13g2_decap_8 FILLER_47_2323 ();
 sg13g2_decap_8 FILLER_47_2330 ();
 sg13g2_decap_8 FILLER_47_2337 ();
 sg13g2_decap_8 FILLER_47_2344 ();
 sg13g2_decap_8 FILLER_47_2351 ();
 sg13g2_decap_8 FILLER_47_2358 ();
 sg13g2_decap_8 FILLER_47_2365 ();
 sg13g2_decap_8 FILLER_47_2372 ();
 sg13g2_decap_8 FILLER_47_2379 ();
 sg13g2_decap_8 FILLER_47_2386 ();
 sg13g2_fill_1 FILLER_47_2403 ();
 sg13g2_fill_2 FILLER_47_2410 ();
 sg13g2_decap_8 FILLER_47_2418 ();
 sg13g2_decap_8 FILLER_47_2425 ();
 sg13g2_decap_8 FILLER_47_2432 ();
 sg13g2_decap_8 FILLER_47_2439 ();
 sg13g2_fill_2 FILLER_47_2446 ();
 sg13g2_fill_1 FILLER_47_2448 ();
 sg13g2_decap_8 FILLER_47_2475 ();
 sg13g2_fill_1 FILLER_47_2482 ();
 sg13g2_decap_8 FILLER_47_2486 ();
 sg13g2_decap_8 FILLER_47_2493 ();
 sg13g2_decap_8 FILLER_47_2500 ();
 sg13g2_decap_4 FILLER_47_2507 ();
 sg13g2_decap_8 FILLER_47_2537 ();
 sg13g2_decap_4 FILLER_47_2544 ();
 sg13g2_fill_2 FILLER_47_2548 ();
 sg13g2_decap_8 FILLER_47_2576 ();
 sg13g2_decap_8 FILLER_47_2583 ();
 sg13g2_fill_2 FILLER_47_2590 ();
 sg13g2_decap_8 FILLER_47_2598 ();
 sg13g2_decap_8 FILLER_47_2605 ();
 sg13g2_decap_8 FILLER_47_2612 ();
 sg13g2_decap_8 FILLER_47_2619 ();
 sg13g2_decap_8 FILLER_47_2626 ();
 sg13g2_decap_8 FILLER_47_2633 ();
 sg13g2_decap_8 FILLER_47_2640 ();
 sg13g2_decap_8 FILLER_47_2647 ();
 sg13g2_decap_8 FILLER_47_2654 ();
 sg13g2_decap_8 FILLER_47_2661 ();
 sg13g2_decap_8 FILLER_47_2668 ();
 sg13g2_decap_8 FILLER_47_2675 ();
 sg13g2_decap_8 FILLER_47_2682 ();
 sg13g2_decap_8 FILLER_47_2689 ();
 sg13g2_decap_4 FILLER_47_2696 ();
 sg13g2_fill_1 FILLER_47_2700 ();
 sg13g2_decap_8 FILLER_47_2753 ();
 sg13g2_decap_8 FILLER_47_2760 ();
 sg13g2_fill_2 FILLER_47_2840 ();
 sg13g2_fill_1 FILLER_47_2842 ();
 sg13g2_decap_8 FILLER_47_2851 ();
 sg13g2_decap_8 FILLER_47_2858 ();
 sg13g2_decap_4 FILLER_47_2865 ();
 sg13g2_fill_1 FILLER_47_2869 ();
 sg13g2_decap_8 FILLER_47_2880 ();
 sg13g2_decap_8 FILLER_47_2887 ();
 sg13g2_decap_8 FILLER_47_2894 ();
 sg13g2_decap_8 FILLER_47_2901 ();
 sg13g2_decap_8 FILLER_47_2908 ();
 sg13g2_decap_8 FILLER_47_2915 ();
 sg13g2_fill_2 FILLER_47_2922 ();
 sg13g2_fill_1 FILLER_47_2924 ();
 sg13g2_fill_1 FILLER_47_2935 ();
 sg13g2_decap_8 FILLER_47_3012 ();
 sg13g2_decap_8 FILLER_47_3019 ();
 sg13g2_decap_8 FILLER_47_3026 ();
 sg13g2_decap_8 FILLER_47_3033 ();
 sg13g2_decap_8 FILLER_47_3040 ();
 sg13g2_decap_8 FILLER_47_3047 ();
 sg13g2_decap_8 FILLER_47_3054 ();
 sg13g2_decap_8 FILLER_47_3061 ();
 sg13g2_decap_8 FILLER_47_3068 ();
 sg13g2_decap_8 FILLER_47_3075 ();
 sg13g2_decap_8 FILLER_47_3082 ();
 sg13g2_decap_8 FILLER_47_3089 ();
 sg13g2_decap_8 FILLER_47_3096 ();
 sg13g2_decap_8 FILLER_47_3103 ();
 sg13g2_decap_8 FILLER_47_3110 ();
 sg13g2_fill_2 FILLER_47_3117 ();
 sg13g2_decap_8 FILLER_47_3128 ();
 sg13g2_decap_8 FILLER_47_3135 ();
 sg13g2_decap_8 FILLER_47_3142 ();
 sg13g2_decap_8 FILLER_47_3149 ();
 sg13g2_decap_8 FILLER_47_3156 ();
 sg13g2_decap_8 FILLER_47_3163 ();
 sg13g2_decap_8 FILLER_47_3170 ();
 sg13g2_decap_8 FILLER_47_3177 ();
 sg13g2_decap_8 FILLER_47_3184 ();
 sg13g2_decap_4 FILLER_47_3191 ();
 sg13g2_fill_1 FILLER_47_3195 ();
 sg13g2_decap_8 FILLER_47_3200 ();
 sg13g2_fill_1 FILLER_47_3207 ();
 sg13g2_decap_8 FILLER_47_3217 ();
 sg13g2_decap_8 FILLER_47_3224 ();
 sg13g2_decap_8 FILLER_47_3231 ();
 sg13g2_decap_8 FILLER_47_3238 ();
 sg13g2_decap_8 FILLER_47_3245 ();
 sg13g2_decap_8 FILLER_47_3252 ();
 sg13g2_fill_2 FILLER_47_3259 ();
 sg13g2_decap_8 FILLER_47_3271 ();
 sg13g2_fill_2 FILLER_47_3278 ();
 sg13g2_decap_8 FILLER_47_3306 ();
 sg13g2_decap_8 FILLER_47_3313 ();
 sg13g2_fill_2 FILLER_47_3320 ();
 sg13g2_decap_8 FILLER_47_3348 ();
 sg13g2_decap_8 FILLER_47_3355 ();
 sg13g2_decap_8 FILLER_47_3362 ();
 sg13g2_decap_8 FILLER_47_3369 ();
 sg13g2_decap_8 FILLER_47_3376 ();
 sg13g2_decap_8 FILLER_47_3383 ();
 sg13g2_decap_8 FILLER_47_3390 ();
 sg13g2_fill_2 FILLER_47_3397 ();
 sg13g2_decap_8 FILLER_47_3429 ();
 sg13g2_fill_2 FILLER_47_3436 ();
 sg13g2_fill_1 FILLER_47_3438 ();
 sg13g2_decap_8 FILLER_47_3464 ();
 sg13g2_decap_8 FILLER_47_3471 ();
 sg13g2_decap_8 FILLER_47_3478 ();
 sg13g2_decap_8 FILLER_47_3485 ();
 sg13g2_decap_8 FILLER_47_3492 ();
 sg13g2_decap_8 FILLER_47_3499 ();
 sg13g2_decap_8 FILLER_47_3506 ();
 sg13g2_decap_8 FILLER_47_3513 ();
 sg13g2_decap_8 FILLER_47_3520 ();
 sg13g2_decap_4 FILLER_47_3527 ();
 sg13g2_decap_8 FILLER_47_3551 ();
 sg13g2_decap_8 FILLER_47_3558 ();
 sg13g2_decap_8 FILLER_47_3565 ();
 sg13g2_decap_8 FILLER_47_3572 ();
 sg13g2_fill_1 FILLER_47_3579 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_decap_8 FILLER_48_14 ();
 sg13g2_decap_8 FILLER_48_21 ();
 sg13g2_decap_8 FILLER_48_28 ();
 sg13g2_decap_8 FILLER_48_35 ();
 sg13g2_decap_8 FILLER_48_42 ();
 sg13g2_decap_8 FILLER_48_49 ();
 sg13g2_decap_4 FILLER_48_56 ();
 sg13g2_fill_1 FILLER_48_60 ();
 sg13g2_fill_2 FILLER_48_66 ();
 sg13g2_fill_1 FILLER_48_68 ();
 sg13g2_decap_8 FILLER_48_79 ();
 sg13g2_decap_8 FILLER_48_86 ();
 sg13g2_decap_8 FILLER_48_93 ();
 sg13g2_decap_8 FILLER_48_100 ();
 sg13g2_decap_8 FILLER_48_107 ();
 sg13g2_decap_8 FILLER_48_114 ();
 sg13g2_decap_8 FILLER_48_121 ();
 sg13g2_decap_4 FILLER_48_128 ();
 sg13g2_fill_1 FILLER_48_132 ();
 sg13g2_fill_1 FILLER_48_138 ();
 sg13g2_fill_1 FILLER_48_148 ();
 sg13g2_fill_1 FILLER_48_163 ();
 sg13g2_fill_1 FILLER_48_175 ();
 sg13g2_decap_8 FILLER_48_221 ();
 sg13g2_decap_8 FILLER_48_228 ();
 sg13g2_decap_8 FILLER_48_235 ();
 sg13g2_decap_4 FILLER_48_242 ();
 sg13g2_fill_1 FILLER_48_246 ();
 sg13g2_decap_8 FILLER_48_251 ();
 sg13g2_decap_4 FILLER_48_258 ();
 sg13g2_fill_2 FILLER_48_262 ();
 sg13g2_decap_4 FILLER_48_268 ();
 sg13g2_fill_2 FILLER_48_272 ();
 sg13g2_decap_8 FILLER_48_291 ();
 sg13g2_decap_8 FILLER_48_298 ();
 sg13g2_decap_8 FILLER_48_305 ();
 sg13g2_decap_4 FILLER_48_312 ();
 sg13g2_fill_2 FILLER_48_316 ();
 sg13g2_decap_8 FILLER_48_356 ();
 sg13g2_decap_8 FILLER_48_363 ();
 sg13g2_decap_8 FILLER_48_370 ();
 sg13g2_decap_4 FILLER_48_377 ();
 sg13g2_decap_8 FILLER_48_395 ();
 sg13g2_decap_8 FILLER_48_402 ();
 sg13g2_decap_8 FILLER_48_409 ();
 sg13g2_decap_8 FILLER_48_416 ();
 sg13g2_decap_8 FILLER_48_423 ();
 sg13g2_decap_4 FILLER_48_430 ();
 sg13g2_decap_8 FILLER_48_458 ();
 sg13g2_decap_8 FILLER_48_465 ();
 sg13g2_decap_4 FILLER_48_478 ();
 sg13g2_decap_8 FILLER_48_499 ();
 sg13g2_decap_8 FILLER_48_506 ();
 sg13g2_decap_4 FILLER_48_513 ();
 sg13g2_fill_2 FILLER_48_517 ();
 sg13g2_decap_4 FILLER_48_548 ();
 sg13g2_fill_2 FILLER_48_552 ();
 sg13g2_decap_8 FILLER_48_557 ();
 sg13g2_decap_8 FILLER_48_564 ();
 sg13g2_decap_8 FILLER_48_577 ();
 sg13g2_decap_8 FILLER_48_584 ();
 sg13g2_decap_8 FILLER_48_591 ();
 sg13g2_decap_8 FILLER_48_598 ();
 sg13g2_fill_2 FILLER_48_605 ();
 sg13g2_decap_8 FILLER_48_622 ();
 sg13g2_decap_4 FILLER_48_629 ();
 sg13g2_fill_2 FILLER_48_633 ();
 sg13g2_decap_8 FILLER_48_654 ();
 sg13g2_decap_4 FILLER_48_664 ();
 sg13g2_decap_8 FILLER_48_694 ();
 sg13g2_decap_8 FILLER_48_701 ();
 sg13g2_decap_8 FILLER_48_708 ();
 sg13g2_decap_4 FILLER_48_715 ();
 sg13g2_fill_2 FILLER_48_723 ();
 sg13g2_decap_8 FILLER_48_729 ();
 sg13g2_fill_2 FILLER_48_736 ();
 sg13g2_decap_8 FILLER_48_764 ();
 sg13g2_decap_8 FILLER_48_771 ();
 sg13g2_decap_8 FILLER_48_778 ();
 sg13g2_decap_8 FILLER_48_785 ();
 sg13g2_decap_8 FILLER_48_792 ();
 sg13g2_decap_8 FILLER_48_799 ();
 sg13g2_decap_8 FILLER_48_806 ();
 sg13g2_decap_4 FILLER_48_813 ();
 sg13g2_fill_2 FILLER_48_817 ();
 sg13g2_decap_4 FILLER_48_824 ();
 sg13g2_fill_1 FILLER_48_828 ();
 sg13g2_fill_2 FILLER_48_834 ();
 sg13g2_fill_1 FILLER_48_836 ();
 sg13g2_decap_8 FILLER_48_858 ();
 sg13g2_decap_8 FILLER_48_865 ();
 sg13g2_decap_8 FILLER_48_872 ();
 sg13g2_decap_4 FILLER_48_879 ();
 sg13g2_decap_8 FILLER_48_899 ();
 sg13g2_decap_8 FILLER_48_906 ();
 sg13g2_fill_2 FILLER_48_913 ();
 sg13g2_fill_1 FILLER_48_915 ();
 sg13g2_fill_1 FILLER_48_936 ();
 sg13g2_decap_8 FILLER_48_951 ();
 sg13g2_decap_8 FILLER_48_958 ();
 sg13g2_decap_8 FILLER_48_965 ();
 sg13g2_decap_8 FILLER_48_972 ();
 sg13g2_decap_8 FILLER_48_979 ();
 sg13g2_fill_2 FILLER_48_986 ();
 sg13g2_fill_2 FILLER_48_1001 ();
 sg13g2_decap_8 FILLER_48_1025 ();
 sg13g2_decap_8 FILLER_48_1032 ();
 sg13g2_decap_8 FILLER_48_1039 ();
 sg13g2_fill_2 FILLER_48_1046 ();
 sg13g2_fill_1 FILLER_48_1048 ();
 sg13g2_fill_2 FILLER_48_1080 ();
 sg13g2_decap_8 FILLER_48_1090 ();
 sg13g2_decap_8 FILLER_48_1097 ();
 sg13g2_decap_8 FILLER_48_1104 ();
 sg13g2_decap_8 FILLER_48_1111 ();
 sg13g2_fill_2 FILLER_48_1147 ();
 sg13g2_decap_8 FILLER_48_1159 ();
 sg13g2_decap_8 FILLER_48_1166 ();
 sg13g2_decap_8 FILLER_48_1173 ();
 sg13g2_decap_8 FILLER_48_1180 ();
 sg13g2_decap_8 FILLER_48_1187 ();
 sg13g2_decap_8 FILLER_48_1194 ();
 sg13g2_decap_8 FILLER_48_1201 ();
 sg13g2_decap_8 FILLER_48_1208 ();
 sg13g2_decap_8 FILLER_48_1215 ();
 sg13g2_decap_8 FILLER_48_1222 ();
 sg13g2_fill_2 FILLER_48_1229 ();
 sg13g2_fill_1 FILLER_48_1231 ();
 sg13g2_decap_8 FILLER_48_1257 ();
 sg13g2_decap_8 FILLER_48_1264 ();
 sg13g2_decap_8 FILLER_48_1271 ();
 sg13g2_decap_8 FILLER_48_1278 ();
 sg13g2_decap_8 FILLER_48_1285 ();
 sg13g2_decap_8 FILLER_48_1292 ();
 sg13g2_decap_8 FILLER_48_1299 ();
 sg13g2_decap_8 FILLER_48_1306 ();
 sg13g2_decap_4 FILLER_48_1313 ();
 sg13g2_decap_8 FILLER_48_1343 ();
 sg13g2_decap_8 FILLER_48_1350 ();
 sg13g2_fill_2 FILLER_48_1357 ();
 sg13g2_decap_8 FILLER_48_1385 ();
 sg13g2_decap_8 FILLER_48_1392 ();
 sg13g2_decap_8 FILLER_48_1409 ();
 sg13g2_decap_8 FILLER_48_1416 ();
 sg13g2_decap_8 FILLER_48_1423 ();
 sg13g2_decap_8 FILLER_48_1430 ();
 sg13g2_decap_8 FILLER_48_1437 ();
 sg13g2_decap_8 FILLER_48_1444 ();
 sg13g2_fill_1 FILLER_48_1451 ();
 sg13g2_fill_2 FILLER_48_1455 ();
 sg13g2_fill_1 FILLER_48_1457 ();
 sg13g2_decap_8 FILLER_48_1494 ();
 sg13g2_decap_8 FILLER_48_1501 ();
 sg13g2_decap_8 FILLER_48_1508 ();
 sg13g2_decap_8 FILLER_48_1515 ();
 sg13g2_decap_8 FILLER_48_1522 ();
 sg13g2_decap_8 FILLER_48_1529 ();
 sg13g2_decap_4 FILLER_48_1536 ();
 sg13g2_decap_8 FILLER_48_1576 ();
 sg13g2_decap_8 FILLER_48_1583 ();
 sg13g2_decap_8 FILLER_48_1590 ();
 sg13g2_decap_8 FILLER_48_1597 ();
 sg13g2_fill_1 FILLER_48_1604 ();
 sg13g2_decap_8 FILLER_48_1621 ();
 sg13g2_decap_8 FILLER_48_1628 ();
 sg13g2_decap_4 FILLER_48_1635 ();
 sg13g2_decap_8 FILLER_48_1665 ();
 sg13g2_decap_8 FILLER_48_1672 ();
 sg13g2_decap_8 FILLER_48_1679 ();
 sg13g2_decap_8 FILLER_48_1686 ();
 sg13g2_decap_8 FILLER_48_1693 ();
 sg13g2_decap_8 FILLER_48_1700 ();
 sg13g2_decap_4 FILLER_48_1707 ();
 sg13g2_fill_2 FILLER_48_1711 ();
 sg13g2_decap_8 FILLER_48_1739 ();
 sg13g2_decap_8 FILLER_48_1746 ();
 sg13g2_decap_8 FILLER_48_1753 ();
 sg13g2_decap_4 FILLER_48_1760 ();
 sg13g2_decap_8 FILLER_48_1788 ();
 sg13g2_decap_8 FILLER_48_1795 ();
 sg13g2_decap_8 FILLER_48_1802 ();
 sg13g2_decap_4 FILLER_48_1809 ();
 sg13g2_decap_8 FILLER_48_1822 ();
 sg13g2_decap_8 FILLER_48_1829 ();
 sg13g2_decap_8 FILLER_48_1836 ();
 sg13g2_decap_8 FILLER_48_1843 ();
 sg13g2_decap_8 FILLER_48_1850 ();
 sg13g2_decap_8 FILLER_48_1857 ();
 sg13g2_decap_8 FILLER_48_1864 ();
 sg13g2_decap_8 FILLER_48_1871 ();
 sg13g2_decap_8 FILLER_48_1878 ();
 sg13g2_decap_8 FILLER_48_1885 ();
 sg13g2_decap_8 FILLER_48_1892 ();
 sg13g2_decap_8 FILLER_48_1899 ();
 sg13g2_decap_8 FILLER_48_1906 ();
 sg13g2_decap_8 FILLER_48_1913 ();
 sg13g2_decap_8 FILLER_48_1920 ();
 sg13g2_decap_8 FILLER_48_1927 ();
 sg13g2_decap_8 FILLER_48_1934 ();
 sg13g2_decap_4 FILLER_48_1941 ();
 sg13g2_decap_8 FILLER_48_1949 ();
 sg13g2_decap_8 FILLER_48_1956 ();
 sg13g2_decap_4 FILLER_48_1963 ();
 sg13g2_decap_8 FILLER_48_1997 ();
 sg13g2_decap_8 FILLER_48_2004 ();
 sg13g2_decap_8 FILLER_48_2011 ();
 sg13g2_decap_8 FILLER_48_2018 ();
 sg13g2_decap_8 FILLER_48_2025 ();
 sg13g2_fill_1 FILLER_48_2032 ();
 sg13g2_decap_8 FILLER_48_2039 ();
 sg13g2_decap_8 FILLER_48_2046 ();
 sg13g2_decap_8 FILLER_48_2053 ();
 sg13g2_decap_8 FILLER_48_2060 ();
 sg13g2_decap_8 FILLER_48_2067 ();
 sg13g2_decap_8 FILLER_48_2074 ();
 sg13g2_decap_8 FILLER_48_2081 ();
 sg13g2_decap_8 FILLER_48_2088 ();
 sg13g2_decap_8 FILLER_48_2095 ();
 sg13g2_decap_8 FILLER_48_2102 ();
 sg13g2_decap_8 FILLER_48_2109 ();
 sg13g2_decap_8 FILLER_48_2116 ();
 sg13g2_fill_2 FILLER_48_2123 ();
 sg13g2_fill_1 FILLER_48_2125 ();
 sg13g2_decap_8 FILLER_48_2132 ();
 sg13g2_fill_2 FILLER_48_2139 ();
 sg13g2_fill_1 FILLER_48_2141 ();
 sg13g2_fill_1 FILLER_48_2146 ();
 sg13g2_fill_2 FILLER_48_2157 ();
 sg13g2_decap_8 FILLER_48_2165 ();
 sg13g2_decap_8 FILLER_48_2172 ();
 sg13g2_decap_8 FILLER_48_2179 ();
 sg13g2_decap_8 FILLER_48_2186 ();
 sg13g2_fill_2 FILLER_48_2193 ();
 sg13g2_decap_4 FILLER_48_2201 ();
 sg13g2_fill_1 FILLER_48_2205 ();
 sg13g2_decap_8 FILLER_48_2226 ();
 sg13g2_decap_8 FILLER_48_2233 ();
 sg13g2_decap_8 FILLER_48_2240 ();
 sg13g2_decap_8 FILLER_48_2247 ();
 sg13g2_decap_8 FILLER_48_2254 ();
 sg13g2_decap_8 FILLER_48_2261 ();
 sg13g2_decap_8 FILLER_48_2268 ();
 sg13g2_decap_8 FILLER_48_2288 ();
 sg13g2_decap_4 FILLER_48_2295 ();
 sg13g2_fill_2 FILLER_48_2299 ();
 sg13g2_decap_8 FILLER_48_2327 ();
 sg13g2_decap_4 FILLER_48_2334 ();
 sg13g2_decap_8 FILLER_48_2348 ();
 sg13g2_decap_8 FILLER_48_2355 ();
 sg13g2_fill_2 FILLER_48_2362 ();
 sg13g2_decap_8 FILLER_48_2373 ();
 sg13g2_fill_2 FILLER_48_2380 ();
 sg13g2_decap_8 FILLER_48_2414 ();
 sg13g2_fill_1 FILLER_48_2421 ();
 sg13g2_decap_8 FILLER_48_2428 ();
 sg13g2_decap_4 FILLER_48_2435 ();
 sg13g2_fill_1 FILLER_48_2439 ();
 sg13g2_decap_8 FILLER_48_2466 ();
 sg13g2_decap_8 FILLER_48_2473 ();
 sg13g2_decap_8 FILLER_48_2480 ();
 sg13g2_decap_8 FILLER_48_2487 ();
 sg13g2_fill_2 FILLER_48_2494 ();
 sg13g2_decap_4 FILLER_48_2521 ();
 sg13g2_decap_8 FILLER_48_2530 ();
 sg13g2_decap_8 FILLER_48_2537 ();
 sg13g2_decap_8 FILLER_48_2544 ();
 sg13g2_decap_8 FILLER_48_2551 ();
 sg13g2_fill_2 FILLER_48_2558 ();
 sg13g2_decap_8 FILLER_48_2568 ();
 sg13g2_decap_8 FILLER_48_2575 ();
 sg13g2_decap_8 FILLER_48_2582 ();
 sg13g2_decap_8 FILLER_48_2589 ();
 sg13g2_decap_8 FILLER_48_2596 ();
 sg13g2_decap_8 FILLER_48_2603 ();
 sg13g2_decap_8 FILLER_48_2610 ();
 sg13g2_decap_8 FILLER_48_2617 ();
 sg13g2_decap_8 FILLER_48_2624 ();
 sg13g2_decap_8 FILLER_48_2631 ();
 sg13g2_decap_8 FILLER_48_2638 ();
 sg13g2_decap_8 FILLER_48_2645 ();
 sg13g2_fill_1 FILLER_48_2652 ();
 sg13g2_decap_8 FILLER_48_2677 ();
 sg13g2_fill_1 FILLER_48_2684 ();
 sg13g2_decap_4 FILLER_48_2696 ();
 sg13g2_decap_4 FILLER_48_2704 ();
 sg13g2_fill_1 FILLER_48_2708 ();
 sg13g2_decap_8 FILLER_48_2713 ();
 sg13g2_decap_8 FILLER_48_2720 ();
 sg13g2_decap_4 FILLER_48_2727 ();
 sg13g2_decap_8 FILLER_48_2737 ();
 sg13g2_decap_8 FILLER_48_2744 ();
 sg13g2_decap_8 FILLER_48_2751 ();
 sg13g2_decap_8 FILLER_48_2758 ();
 sg13g2_decap_8 FILLER_48_2765 ();
 sg13g2_decap_8 FILLER_48_2772 ();
 sg13g2_fill_2 FILLER_48_2779 ();
 sg13g2_decap_8 FILLER_48_2807 ();
 sg13g2_decap_8 FILLER_48_2814 ();
 sg13g2_decap_8 FILLER_48_2821 ();
 sg13g2_decap_8 FILLER_48_2828 ();
 sg13g2_decap_8 FILLER_48_2835 ();
 sg13g2_decap_8 FILLER_48_2842 ();
 sg13g2_decap_8 FILLER_48_2849 ();
 sg13g2_decap_8 FILLER_48_2856 ();
 sg13g2_decap_8 FILLER_48_2863 ();
 sg13g2_decap_8 FILLER_48_2870 ();
 sg13g2_decap_8 FILLER_48_2877 ();
 sg13g2_decap_8 FILLER_48_2884 ();
 sg13g2_decap_8 FILLER_48_2891 ();
 sg13g2_decap_8 FILLER_48_2898 ();
 sg13g2_decap_8 FILLER_48_2905 ();
 sg13g2_decap_8 FILLER_48_2912 ();
 sg13g2_decap_8 FILLER_48_2919 ();
 sg13g2_fill_1 FILLER_48_2926 ();
 sg13g2_decap_8 FILLER_48_2953 ();
 sg13g2_decap_8 FILLER_48_2960 ();
 sg13g2_decap_8 FILLER_48_2967 ();
 sg13g2_decap_8 FILLER_48_2974 ();
 sg13g2_decap_4 FILLER_48_2981 ();
 sg13g2_decap_8 FILLER_48_2993 ();
 sg13g2_decap_8 FILLER_48_3000 ();
 sg13g2_decap_8 FILLER_48_3007 ();
 sg13g2_decap_8 FILLER_48_3014 ();
 sg13g2_decap_8 FILLER_48_3021 ();
 sg13g2_decap_4 FILLER_48_3033 ();
 sg13g2_fill_1 FILLER_48_3037 ();
 sg13g2_decap_8 FILLER_48_3046 ();
 sg13g2_decap_8 FILLER_48_3053 ();
 sg13g2_decap_8 FILLER_48_3060 ();
 sg13g2_decap_8 FILLER_48_3067 ();
 sg13g2_decap_8 FILLER_48_3074 ();
 sg13g2_decap_8 FILLER_48_3081 ();
 sg13g2_decap_8 FILLER_48_3088 ();
 sg13g2_decap_4 FILLER_48_3095 ();
 sg13g2_decap_8 FILLER_48_3135 ();
 sg13g2_decap_8 FILLER_48_3142 ();
 sg13g2_decap_8 FILLER_48_3149 ();
 sg13g2_decap_4 FILLER_48_3156 ();
 sg13g2_decap_8 FILLER_48_3170 ();
 sg13g2_decap_8 FILLER_48_3177 ();
 sg13g2_decap_8 FILLER_48_3184 ();
 sg13g2_decap_8 FILLER_48_3239 ();
 sg13g2_decap_8 FILLER_48_3246 ();
 sg13g2_decap_8 FILLER_48_3253 ();
 sg13g2_decap_4 FILLER_48_3260 ();
 sg13g2_fill_1 FILLER_48_3264 ();
 sg13g2_decap_8 FILLER_48_3275 ();
 sg13g2_decap_8 FILLER_48_3282 ();
 sg13g2_decap_8 FILLER_48_3289 ();
 sg13g2_decap_8 FILLER_48_3296 ();
 sg13g2_decap_8 FILLER_48_3303 ();
 sg13g2_decap_8 FILLER_48_3310 ();
 sg13g2_decap_8 FILLER_48_3317 ();
 sg13g2_decap_8 FILLER_48_3324 ();
 sg13g2_decap_4 FILLER_48_3331 ();
 sg13g2_fill_1 FILLER_48_3335 ();
 sg13g2_fill_2 FILLER_48_3342 ();
 sg13g2_decap_8 FILLER_48_3354 ();
 sg13g2_decap_8 FILLER_48_3361 ();
 sg13g2_decap_8 FILLER_48_3368 ();
 sg13g2_decap_8 FILLER_48_3375 ();
 sg13g2_decap_8 FILLER_48_3382 ();
 sg13g2_decap_8 FILLER_48_3389 ();
 sg13g2_fill_2 FILLER_48_3396 ();
 sg13g2_fill_1 FILLER_48_3398 ();
 sg13g2_decap_8 FILLER_48_3434 ();
 sg13g2_decap_8 FILLER_48_3441 ();
 sg13g2_decap_8 FILLER_48_3448 ();
 sg13g2_decap_8 FILLER_48_3455 ();
 sg13g2_decap_8 FILLER_48_3462 ();
 sg13g2_decap_8 FILLER_48_3469 ();
 sg13g2_decap_4 FILLER_48_3476 ();
 sg13g2_fill_1 FILLER_48_3480 ();
 sg13g2_fill_1 FILLER_48_3491 ();
 sg13g2_decap_8 FILLER_48_3497 ();
 sg13g2_decap_8 FILLER_48_3504 ();
 sg13g2_decap_8 FILLER_48_3511 ();
 sg13g2_decap_8 FILLER_48_3518 ();
 sg13g2_fill_1 FILLER_48_3525 ();
 sg13g2_decap_8 FILLER_48_3536 ();
 sg13g2_decap_8 FILLER_48_3543 ();
 sg13g2_decap_8 FILLER_48_3550 ();
 sg13g2_decap_8 FILLER_48_3557 ();
 sg13g2_decap_8 FILLER_48_3564 ();
 sg13g2_decap_8 FILLER_48_3571 ();
 sg13g2_fill_2 FILLER_48_3578 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_4 FILLER_49_7 ();
 sg13g2_fill_2 FILLER_49_11 ();
 sg13g2_decap_8 FILLER_49_39 ();
 sg13g2_decap_8 FILLER_49_46 ();
 sg13g2_decap_8 FILLER_49_53 ();
 sg13g2_decap_8 FILLER_49_60 ();
 sg13g2_decap_4 FILLER_49_67 ();
 sg13g2_fill_1 FILLER_49_71 ();
 sg13g2_decap_8 FILLER_49_94 ();
 sg13g2_decap_8 FILLER_49_101 ();
 sg13g2_decap_8 FILLER_49_108 ();
 sg13g2_decap_8 FILLER_49_115 ();
 sg13g2_decap_8 FILLER_49_122 ();
 sg13g2_decap_4 FILLER_49_129 ();
 sg13g2_fill_2 FILLER_49_145 ();
 sg13g2_fill_1 FILLER_49_147 ();
 sg13g2_decap_8 FILLER_49_158 ();
 sg13g2_decap_8 FILLER_49_165 ();
 sg13g2_decap_8 FILLER_49_172 ();
 sg13g2_decap_8 FILLER_49_179 ();
 sg13g2_fill_2 FILLER_49_186 ();
 sg13g2_fill_2 FILLER_49_193 ();
 sg13g2_fill_1 FILLER_49_195 ();
 sg13g2_decap_8 FILLER_49_202 ();
 sg13g2_decap_8 FILLER_49_209 ();
 sg13g2_decap_8 FILLER_49_216 ();
 sg13g2_decap_8 FILLER_49_223 ();
 sg13g2_decap_8 FILLER_49_230 ();
 sg13g2_decap_8 FILLER_49_237 ();
 sg13g2_decap_8 FILLER_49_244 ();
 sg13g2_decap_8 FILLER_49_251 ();
 sg13g2_decap_8 FILLER_49_258 ();
 sg13g2_fill_2 FILLER_49_265 ();
 sg13g2_decap_8 FILLER_49_272 ();
 sg13g2_decap_8 FILLER_49_279 ();
 sg13g2_decap_8 FILLER_49_289 ();
 sg13g2_decap_8 FILLER_49_296 ();
 sg13g2_decap_8 FILLER_49_303 ();
 sg13g2_decap_8 FILLER_49_310 ();
 sg13g2_decap_4 FILLER_49_325 ();
 sg13g2_fill_2 FILLER_49_337 ();
 sg13g2_decap_4 FILLER_49_342 ();
 sg13g2_fill_1 FILLER_49_346 ();
 sg13g2_decap_8 FILLER_49_358 ();
 sg13g2_fill_2 FILLER_49_365 ();
 sg13g2_decap_8 FILLER_49_393 ();
 sg13g2_decap_8 FILLER_49_400 ();
 sg13g2_decap_8 FILLER_49_407 ();
 sg13g2_decap_8 FILLER_49_414 ();
 sg13g2_decap_8 FILLER_49_421 ();
 sg13g2_decap_4 FILLER_49_428 ();
 sg13g2_decap_8 FILLER_49_465 ();
 sg13g2_decap_8 FILLER_49_472 ();
 sg13g2_fill_1 FILLER_49_479 ();
 sg13g2_decap_8 FILLER_49_492 ();
 sg13g2_decap_4 FILLER_49_499 ();
 sg13g2_decap_8 FILLER_49_515 ();
 sg13g2_decap_8 FILLER_49_522 ();
 sg13g2_decap_8 FILLER_49_529 ();
 sg13g2_decap_8 FILLER_49_536 ();
 sg13g2_fill_2 FILLER_49_543 ();
 sg13g2_fill_1 FILLER_49_553 ();
 sg13g2_decap_4 FILLER_49_583 ();
 sg13g2_decap_8 FILLER_49_595 ();
 sg13g2_decap_8 FILLER_49_602 ();
 sg13g2_fill_2 FILLER_49_609 ();
 sg13g2_fill_1 FILLER_49_611 ();
 sg13g2_decap_8 FILLER_49_616 ();
 sg13g2_fill_1 FILLER_49_623 ();
 sg13g2_decap_8 FILLER_49_653 ();
 sg13g2_decap_8 FILLER_49_660 ();
 sg13g2_decap_4 FILLER_49_667 ();
 sg13g2_fill_1 FILLER_49_671 ();
 sg13g2_fill_2 FILLER_49_698 ();
 sg13g2_decap_8 FILLER_49_705 ();
 sg13g2_decap_8 FILLER_49_734 ();
 sg13g2_fill_2 FILLER_49_741 ();
 sg13g2_fill_1 FILLER_49_743 ();
 sg13g2_decap_8 FILLER_49_749 ();
 sg13g2_decap_8 FILLER_49_756 ();
 sg13g2_decap_8 FILLER_49_763 ();
 sg13g2_decap_8 FILLER_49_770 ();
 sg13g2_decap_8 FILLER_49_777 ();
 sg13g2_decap_4 FILLER_49_784 ();
 sg13g2_fill_1 FILLER_49_788 ();
 sg13g2_decap_4 FILLER_49_808 ();
 sg13g2_fill_2 FILLER_49_812 ();
 sg13g2_decap_8 FILLER_49_818 ();
 sg13g2_decap_8 FILLER_49_825 ();
 sg13g2_decap_8 FILLER_49_832 ();
 sg13g2_decap_4 FILLER_49_839 ();
 sg13g2_fill_1 FILLER_49_843 ();
 sg13g2_decap_8 FILLER_49_852 ();
 sg13g2_decap_4 FILLER_49_859 ();
 sg13g2_fill_1 FILLER_49_863 ();
 sg13g2_decap_8 FILLER_49_873 ();
 sg13g2_decap_4 FILLER_49_880 ();
 sg13g2_decap_8 FILLER_49_895 ();
 sg13g2_decap_8 FILLER_49_902 ();
 sg13g2_decap_8 FILLER_49_909 ();
 sg13g2_decap_4 FILLER_49_916 ();
 sg13g2_fill_2 FILLER_49_934 ();
 sg13g2_fill_1 FILLER_49_936 ();
 sg13g2_fill_1 FILLER_49_942 ();
 sg13g2_decap_8 FILLER_49_947 ();
 sg13g2_decap_8 FILLER_49_954 ();
 sg13g2_decap_8 FILLER_49_961 ();
 sg13g2_fill_2 FILLER_49_968 ();
 sg13g2_fill_1 FILLER_49_970 ();
 sg13g2_fill_2 FILLER_49_992 ();
 sg13g2_fill_1 FILLER_49_1006 ();
 sg13g2_fill_1 FILLER_49_1012 ();
 sg13g2_decap_8 FILLER_49_1016 ();
 sg13g2_decap_8 FILLER_49_1023 ();
 sg13g2_decap_8 FILLER_49_1030 ();
 sg13g2_decap_8 FILLER_49_1037 ();
 sg13g2_decap_8 FILLER_49_1044 ();
 sg13g2_decap_8 FILLER_49_1051 ();
 sg13g2_decap_8 FILLER_49_1058 ();
 sg13g2_fill_2 FILLER_49_1065 ();
 sg13g2_decap_8 FILLER_49_1071 ();
 sg13g2_fill_1 FILLER_49_1078 ();
 sg13g2_decap_8 FILLER_49_1084 ();
 sg13g2_decap_8 FILLER_49_1091 ();
 sg13g2_decap_8 FILLER_49_1098 ();
 sg13g2_decap_8 FILLER_49_1105 ();
 sg13g2_decap_8 FILLER_49_1112 ();
 sg13g2_decap_8 FILLER_49_1119 ();
 sg13g2_decap_8 FILLER_49_1126 ();
 sg13g2_decap_8 FILLER_49_1133 ();
 sg13g2_decap_8 FILLER_49_1140 ();
 sg13g2_decap_8 FILLER_49_1147 ();
 sg13g2_decap_8 FILLER_49_1154 ();
 sg13g2_decap_8 FILLER_49_1161 ();
 sg13g2_decap_8 FILLER_49_1168 ();
 sg13g2_decap_8 FILLER_49_1175 ();
 sg13g2_decap_8 FILLER_49_1182 ();
 sg13g2_decap_8 FILLER_49_1189 ();
 sg13g2_decap_8 FILLER_49_1196 ();
 sg13g2_decap_8 FILLER_49_1203 ();
 sg13g2_decap_8 FILLER_49_1210 ();
 sg13g2_decap_8 FILLER_49_1217 ();
 sg13g2_fill_2 FILLER_49_1224 ();
 sg13g2_fill_1 FILLER_49_1240 ();
 sg13g2_fill_1 FILLER_49_1246 ();
 sg13g2_decap_8 FILLER_49_1252 ();
 sg13g2_decap_8 FILLER_49_1259 ();
 sg13g2_decap_8 FILLER_49_1266 ();
 sg13g2_decap_8 FILLER_49_1273 ();
 sg13g2_decap_8 FILLER_49_1280 ();
 sg13g2_decap_8 FILLER_49_1287 ();
 sg13g2_decap_8 FILLER_49_1294 ();
 sg13g2_fill_1 FILLER_49_1301 ();
 sg13g2_decap_8 FILLER_49_1348 ();
 sg13g2_decap_8 FILLER_49_1355 ();
 sg13g2_decap_8 FILLER_49_1362 ();
 sg13g2_decap_8 FILLER_49_1369 ();
 sg13g2_decap_8 FILLER_49_1376 ();
 sg13g2_decap_8 FILLER_49_1383 ();
 sg13g2_decap_8 FILLER_49_1390 ();
 sg13g2_fill_1 FILLER_49_1397 ();
 sg13g2_decap_8 FILLER_49_1402 ();
 sg13g2_decap_8 FILLER_49_1409 ();
 sg13g2_decap_8 FILLER_49_1416 ();
 sg13g2_decap_8 FILLER_49_1423 ();
 sg13g2_decap_8 FILLER_49_1430 ();
 sg13g2_decap_8 FILLER_49_1437 ();
 sg13g2_fill_2 FILLER_49_1444 ();
 sg13g2_fill_1 FILLER_49_1446 ();
 sg13g2_decap_8 FILLER_49_1465 ();
 sg13g2_decap_8 FILLER_49_1472 ();
 sg13g2_decap_8 FILLER_49_1479 ();
 sg13g2_decap_8 FILLER_49_1486 ();
 sg13g2_decap_8 FILLER_49_1493 ();
 sg13g2_decap_8 FILLER_49_1500 ();
 sg13g2_decap_8 FILLER_49_1507 ();
 sg13g2_decap_8 FILLER_49_1514 ();
 sg13g2_decap_8 FILLER_49_1521 ();
 sg13g2_decap_8 FILLER_49_1528 ();
 sg13g2_decap_8 FILLER_49_1535 ();
 sg13g2_decap_8 FILLER_49_1542 ();
 sg13g2_decap_8 FILLER_49_1549 ();
 sg13g2_decap_8 FILLER_49_1556 ();
 sg13g2_decap_8 FILLER_49_1563 ();
 sg13g2_decap_8 FILLER_49_1570 ();
 sg13g2_decap_8 FILLER_49_1577 ();
 sg13g2_decap_8 FILLER_49_1584 ();
 sg13g2_decap_4 FILLER_49_1591 ();
 sg13g2_decap_8 FILLER_49_1621 ();
 sg13g2_decap_8 FILLER_49_1638 ();
 sg13g2_decap_8 FILLER_49_1645 ();
 sg13g2_fill_1 FILLER_49_1652 ();
 sg13g2_decap_8 FILLER_49_1661 ();
 sg13g2_decap_8 FILLER_49_1668 ();
 sg13g2_decap_8 FILLER_49_1675 ();
 sg13g2_decap_8 FILLER_49_1682 ();
 sg13g2_decap_8 FILLER_49_1689 ();
 sg13g2_decap_8 FILLER_49_1696 ();
 sg13g2_fill_1 FILLER_49_1703 ();
 sg13g2_decap_8 FILLER_49_1712 ();
 sg13g2_decap_8 FILLER_49_1719 ();
 sg13g2_decap_8 FILLER_49_1726 ();
 sg13g2_decap_8 FILLER_49_1733 ();
 sg13g2_decap_8 FILLER_49_1740 ();
 sg13g2_decap_8 FILLER_49_1747 ();
 sg13g2_decap_8 FILLER_49_1754 ();
 sg13g2_fill_2 FILLER_49_1761 ();
 sg13g2_fill_1 FILLER_49_1763 ();
 sg13g2_decap_8 FILLER_49_1774 ();
 sg13g2_decap_8 FILLER_49_1794 ();
 sg13g2_decap_4 FILLER_49_1801 ();
 sg13g2_fill_2 FILLER_49_1811 ();
 sg13g2_decap_4 FILLER_49_1823 ();
 sg13g2_decap_8 FILLER_49_1853 ();
 sg13g2_decap_8 FILLER_49_1860 ();
 sg13g2_decap_8 FILLER_49_1867 ();
 sg13g2_decap_8 FILLER_49_1874 ();
 sg13g2_decap_8 FILLER_49_1881 ();
 sg13g2_decap_8 FILLER_49_1888 ();
 sg13g2_decap_8 FILLER_49_1895 ();
 sg13g2_decap_4 FILLER_49_1902 ();
 sg13g2_fill_1 FILLER_49_1906 ();
 sg13g2_decap_4 FILLER_49_1912 ();
 sg13g2_decap_8 FILLER_49_1921 ();
 sg13g2_decap_4 FILLER_49_1928 ();
 sg13g2_fill_2 FILLER_49_1932 ();
 sg13g2_decap_8 FILLER_49_1958 ();
 sg13g2_fill_1 FILLER_49_1965 ();
 sg13g2_decap_8 FILLER_49_1970 ();
 sg13g2_decap_8 FILLER_49_1977 ();
 sg13g2_decap_8 FILLER_49_1984 ();
 sg13g2_decap_8 FILLER_49_1991 ();
 sg13g2_decap_8 FILLER_49_1998 ();
 sg13g2_decap_8 FILLER_49_2005 ();
 sg13g2_decap_8 FILLER_49_2012 ();
 sg13g2_decap_8 FILLER_49_2019 ();
 sg13g2_decap_8 FILLER_49_2047 ();
 sg13g2_decap_8 FILLER_49_2054 ();
 sg13g2_decap_8 FILLER_49_2061 ();
 sg13g2_decap_8 FILLER_49_2073 ();
 sg13g2_fill_1 FILLER_49_2080 ();
 sg13g2_decap_8 FILLER_49_2089 ();
 sg13g2_decap_8 FILLER_49_2096 ();
 sg13g2_decap_8 FILLER_49_2103 ();
 sg13g2_decap_4 FILLER_49_2110 ();
 sg13g2_fill_2 FILLER_49_2114 ();
 sg13g2_fill_2 FILLER_49_2124 ();
 sg13g2_fill_2 FILLER_49_2146 ();
 sg13g2_fill_1 FILLER_49_2148 ();
 sg13g2_decap_8 FILLER_49_2175 ();
 sg13g2_decap_4 FILLER_49_2182 ();
 sg13g2_decap_8 FILLER_49_2192 ();
 sg13g2_decap_4 FILLER_49_2199 ();
 sg13g2_fill_2 FILLER_49_2203 ();
 sg13g2_decap_4 FILLER_49_2213 ();
 sg13g2_decap_8 FILLER_49_2225 ();
 sg13g2_decap_8 FILLER_49_2232 ();
 sg13g2_decap_8 FILLER_49_2239 ();
 sg13g2_fill_2 FILLER_49_2246 ();
 sg13g2_decap_8 FILLER_49_2304 ();
 sg13g2_decap_8 FILLER_49_2311 ();
 sg13g2_fill_2 FILLER_49_2376 ();
 sg13g2_decap_8 FILLER_49_2384 ();
 sg13g2_decap_8 FILLER_49_2391 ();
 sg13g2_decap_8 FILLER_49_2398 ();
 sg13g2_decap_8 FILLER_49_2405 ();
 sg13g2_decap_8 FILLER_49_2412 ();
 sg13g2_fill_2 FILLER_49_2419 ();
 sg13g2_fill_1 FILLER_49_2421 ();
 sg13g2_decap_8 FILLER_49_2432 ();
 sg13g2_fill_2 FILLER_49_2439 ();
 sg13g2_fill_2 FILLER_49_2444 ();
 sg13g2_fill_2 FILLER_49_2456 ();
 sg13g2_fill_1 FILLER_49_2458 ();
 sg13g2_decap_8 FILLER_49_2463 ();
 sg13g2_decap_8 FILLER_49_2470 ();
 sg13g2_decap_4 FILLER_49_2477 ();
 sg13g2_fill_2 FILLER_49_2481 ();
 sg13g2_fill_2 FILLER_49_2487 ();
 sg13g2_fill_1 FILLER_49_2489 ();
 sg13g2_decap_8 FILLER_49_2499 ();
 sg13g2_decap_8 FILLER_49_2506 ();
 sg13g2_decap_8 FILLER_49_2513 ();
 sg13g2_decap_8 FILLER_49_2520 ();
 sg13g2_decap_8 FILLER_49_2527 ();
 sg13g2_decap_8 FILLER_49_2534 ();
 sg13g2_decap_8 FILLER_49_2541 ();
 sg13g2_decap_8 FILLER_49_2548 ();
 sg13g2_decap_4 FILLER_49_2555 ();
 sg13g2_fill_2 FILLER_49_2559 ();
 sg13g2_decap_8 FILLER_49_2569 ();
 sg13g2_decap_8 FILLER_49_2576 ();
 sg13g2_decap_8 FILLER_49_2583 ();
 sg13g2_fill_1 FILLER_49_2590 ();
 sg13g2_decap_8 FILLER_49_2627 ();
 sg13g2_decap_8 FILLER_49_2634 ();
 sg13g2_decap_8 FILLER_49_2641 ();
 sg13g2_decap_8 FILLER_49_2648 ();
 sg13g2_decap_8 FILLER_49_2655 ();
 sg13g2_decap_8 FILLER_49_2662 ();
 sg13g2_decap_8 FILLER_49_2669 ();
 sg13g2_decap_4 FILLER_49_2676 ();
 sg13g2_fill_1 FILLER_49_2680 ();
 sg13g2_decap_8 FILLER_49_2694 ();
 sg13g2_decap_8 FILLER_49_2701 ();
 sg13g2_fill_1 FILLER_49_2708 ();
 sg13g2_fill_1 FILLER_49_2717 ();
 sg13g2_decap_8 FILLER_49_2726 ();
 sg13g2_decap_8 FILLER_49_2733 ();
 sg13g2_decap_8 FILLER_49_2740 ();
 sg13g2_decap_8 FILLER_49_2747 ();
 sg13g2_decap_8 FILLER_49_2754 ();
 sg13g2_decap_8 FILLER_49_2761 ();
 sg13g2_decap_8 FILLER_49_2768 ();
 sg13g2_decap_8 FILLER_49_2775 ();
 sg13g2_decap_8 FILLER_49_2782 ();
 sg13g2_decap_8 FILLER_49_2789 ();
 sg13g2_decap_8 FILLER_49_2822 ();
 sg13g2_decap_4 FILLER_49_2829 ();
 sg13g2_fill_1 FILLER_49_2833 ();
 sg13g2_fill_1 FILLER_49_2846 ();
 sg13g2_fill_2 FILLER_49_2883 ();
 sg13g2_fill_1 FILLER_49_2885 ();
 sg13g2_decap_8 FILLER_49_2890 ();
 sg13g2_fill_1 FILLER_49_2897 ();
 sg13g2_decap_4 FILLER_49_2903 ();
 sg13g2_decap_8 FILLER_49_2912 ();
 sg13g2_decap_8 FILLER_49_2919 ();
 sg13g2_decap_8 FILLER_49_2926 ();
 sg13g2_decap_8 FILLER_49_2933 ();
 sg13g2_decap_8 FILLER_49_2940 ();
 sg13g2_decap_8 FILLER_49_2947 ();
 sg13g2_decap_8 FILLER_49_2954 ();
 sg13g2_decap_8 FILLER_49_2961 ();
 sg13g2_decap_8 FILLER_49_2968 ();
 sg13g2_decap_8 FILLER_49_2975 ();
 sg13g2_decap_8 FILLER_49_2982 ();
 sg13g2_decap_8 FILLER_49_2989 ();
 sg13g2_decap_8 FILLER_49_2996 ();
 sg13g2_decap_8 FILLER_49_3003 ();
 sg13g2_fill_2 FILLER_49_3010 ();
 sg13g2_fill_1 FILLER_49_3012 ();
 sg13g2_decap_8 FILLER_49_3039 ();
 sg13g2_decap_8 FILLER_49_3046 ();
 sg13g2_fill_2 FILLER_49_3053 ();
 sg13g2_decap_8 FILLER_49_3060 ();
 sg13g2_decap_8 FILLER_49_3067 ();
 sg13g2_decap_8 FILLER_49_3074 ();
 sg13g2_decap_8 FILLER_49_3100 ();
 sg13g2_fill_2 FILLER_49_3107 ();
 sg13g2_fill_1 FILLER_49_3109 ();
 sg13g2_decap_4 FILLER_49_3120 ();
 sg13g2_fill_1 FILLER_49_3124 ();
 sg13g2_decap_8 FILLER_49_3161 ();
 sg13g2_decap_8 FILLER_49_3194 ();
 sg13g2_decap_8 FILLER_49_3201 ();
 sg13g2_fill_2 FILLER_49_3208 ();
 sg13g2_decap_8 FILLER_49_3216 ();
 sg13g2_decap_8 FILLER_49_3223 ();
 sg13g2_decap_8 FILLER_49_3230 ();
 sg13g2_decap_8 FILLER_49_3237 ();
 sg13g2_fill_2 FILLER_49_3244 ();
 sg13g2_decap_8 FILLER_49_3272 ();
 sg13g2_decap_8 FILLER_49_3279 ();
 sg13g2_decap_8 FILLER_49_3286 ();
 sg13g2_decap_8 FILLER_49_3293 ();
 sg13g2_decap_8 FILLER_49_3300 ();
 sg13g2_decap_8 FILLER_49_3307 ();
 sg13g2_decap_8 FILLER_49_3314 ();
 sg13g2_decap_4 FILLER_49_3321 ();
 sg13g2_decap_8 FILLER_49_3377 ();
 sg13g2_decap_8 FILLER_49_3384 ();
 sg13g2_decap_8 FILLER_49_3391 ();
 sg13g2_decap_8 FILLER_49_3398 ();
 sg13g2_fill_1 FILLER_49_3405 ();
 sg13g2_decap_8 FILLER_49_3432 ();
 sg13g2_decap_8 FILLER_49_3439 ();
 sg13g2_decap_8 FILLER_49_3446 ();
 sg13g2_decap_8 FILLER_49_3453 ();
 sg13g2_decap_8 FILLER_49_3460 ();
 sg13g2_decap_8 FILLER_49_3467 ();
 sg13g2_decap_8 FILLER_49_3479 ();
 sg13g2_decap_4 FILLER_49_3486 ();
 sg13g2_fill_1 FILLER_49_3490 ();
 sg13g2_decap_8 FILLER_49_3512 ();
 sg13g2_decap_8 FILLER_49_3519 ();
 sg13g2_decap_4 FILLER_49_3526 ();
 sg13g2_fill_2 FILLER_49_3530 ();
 sg13g2_fill_2 FILLER_49_3537 ();
 sg13g2_decap_8 FILLER_49_3567 ();
 sg13g2_decap_4 FILLER_49_3574 ();
 sg13g2_fill_2 FILLER_49_3578 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_8 FILLER_50_7 ();
 sg13g2_fill_1 FILLER_50_14 ();
 sg13g2_fill_2 FILLER_50_34 ();
 sg13g2_decap_8 FILLER_50_52 ();
 sg13g2_decap_8 FILLER_50_59 ();
 sg13g2_fill_2 FILLER_50_66 ();
 sg13g2_decap_8 FILLER_50_110 ();
 sg13g2_decap_8 FILLER_50_117 ();
 sg13g2_decap_8 FILLER_50_124 ();
 sg13g2_decap_4 FILLER_50_131 ();
 sg13g2_decap_8 FILLER_50_152 ();
 sg13g2_fill_2 FILLER_50_159 ();
 sg13g2_decap_8 FILLER_50_167 ();
 sg13g2_fill_2 FILLER_50_174 ();
 sg13g2_fill_1 FILLER_50_176 ();
 sg13g2_decap_4 FILLER_50_181 ();
 sg13g2_decap_8 FILLER_50_189 ();
 sg13g2_decap_8 FILLER_50_196 ();
 sg13g2_decap_8 FILLER_50_203 ();
 sg13g2_decap_8 FILLER_50_210 ();
 sg13g2_decap_8 FILLER_50_217 ();
 sg13g2_decap_4 FILLER_50_224 ();
 sg13g2_fill_1 FILLER_50_228 ();
 sg13g2_decap_8 FILLER_50_233 ();
 sg13g2_decap_8 FILLER_50_249 ();
 sg13g2_decap_8 FILLER_50_256 ();
 sg13g2_decap_8 FILLER_50_263 ();
 sg13g2_decap_8 FILLER_50_270 ();
 sg13g2_decap_8 FILLER_50_277 ();
 sg13g2_fill_2 FILLER_50_284 ();
 sg13g2_decap_4 FILLER_50_289 ();
 sg13g2_fill_2 FILLER_50_293 ();
 sg13g2_decap_8 FILLER_50_299 ();
 sg13g2_decap_8 FILLER_50_306 ();
 sg13g2_decap_4 FILLER_50_313 ();
 sg13g2_fill_1 FILLER_50_317 ();
 sg13g2_decap_4 FILLER_50_328 ();
 sg13g2_fill_2 FILLER_50_337 ();
 sg13g2_decap_8 FILLER_50_395 ();
 sg13g2_decap_8 FILLER_50_402 ();
 sg13g2_decap_8 FILLER_50_409 ();
 sg13g2_decap_4 FILLER_50_416 ();
 sg13g2_decap_8 FILLER_50_426 ();
 sg13g2_decap_4 FILLER_50_433 ();
 sg13g2_fill_1 FILLER_50_437 ();
 sg13g2_decap_4 FILLER_50_456 ();
 sg13g2_fill_2 FILLER_50_460 ();
 sg13g2_decap_8 FILLER_50_468 ();
 sg13g2_fill_2 FILLER_50_475 ();
 sg13g2_decap_8 FILLER_50_483 ();
 sg13g2_decap_8 FILLER_50_490 ();
 sg13g2_decap_8 FILLER_50_497 ();
 sg13g2_decap_8 FILLER_50_504 ();
 sg13g2_decap_8 FILLER_50_511 ();
 sg13g2_decap_8 FILLER_50_518 ();
 sg13g2_decap_8 FILLER_50_525 ();
 sg13g2_decap_8 FILLER_50_532 ();
 sg13g2_decap_4 FILLER_50_539 ();
 sg13g2_fill_2 FILLER_50_543 ();
 sg13g2_decap_4 FILLER_50_548 ();
 sg13g2_fill_2 FILLER_50_552 ();
 sg13g2_decap_4 FILLER_50_557 ();
 sg13g2_decap_8 FILLER_50_589 ();
 sg13g2_decap_8 FILLER_50_596 ();
 sg13g2_decap_8 FILLER_50_603 ();
 sg13g2_decap_8 FILLER_50_610 ();
 sg13g2_decap_4 FILLER_50_617 ();
 sg13g2_decap_8 FILLER_50_639 ();
 sg13g2_decap_8 FILLER_50_646 ();
 sg13g2_decap_8 FILLER_50_653 ();
 sg13g2_decap_8 FILLER_50_660 ();
 sg13g2_decap_8 FILLER_50_667 ();
 sg13g2_decap_4 FILLER_50_674 ();
 sg13g2_fill_2 FILLER_50_678 ();
 sg13g2_decap_8 FILLER_50_689 ();
 sg13g2_decap_8 FILLER_50_696 ();
 sg13g2_decap_8 FILLER_50_703 ();
 sg13g2_decap_8 FILLER_50_710 ();
 sg13g2_fill_1 FILLER_50_717 ();
 sg13g2_decap_4 FILLER_50_729 ();
 sg13g2_decap_8 FILLER_50_746 ();
 sg13g2_decap_4 FILLER_50_753 ();
 sg13g2_fill_2 FILLER_50_757 ();
 sg13g2_decap_8 FILLER_50_764 ();
 sg13g2_decap_8 FILLER_50_771 ();
 sg13g2_fill_2 FILLER_50_778 ();
 sg13g2_fill_1 FILLER_50_823 ();
 sg13g2_fill_1 FILLER_50_830 ();
 sg13g2_decap_8 FILLER_50_852 ();
 sg13g2_decap_8 FILLER_50_859 ();
 sg13g2_decap_8 FILLER_50_866 ();
 sg13g2_decap_8 FILLER_50_873 ();
 sg13g2_fill_1 FILLER_50_880 ();
 sg13g2_decap_4 FILLER_50_892 ();
 sg13g2_decap_8 FILLER_50_909 ();
 sg13g2_decap_4 FILLER_50_916 ();
 sg13g2_fill_1 FILLER_50_920 ();
 sg13g2_decap_8 FILLER_50_926 ();
 sg13g2_decap_8 FILLER_50_933 ();
 sg13g2_decap_8 FILLER_50_940 ();
 sg13g2_decap_8 FILLER_50_947 ();
 sg13g2_decap_8 FILLER_50_954 ();
 sg13g2_decap_8 FILLER_50_961 ();
 sg13g2_decap_8 FILLER_50_968 ();
 sg13g2_decap_8 FILLER_50_975 ();
 sg13g2_decap_8 FILLER_50_982 ();
 sg13g2_decap_8 FILLER_50_989 ();
 sg13g2_fill_2 FILLER_50_996 ();
 sg13g2_fill_1 FILLER_50_998 ();
 sg13g2_decap_8 FILLER_50_1004 ();
 sg13g2_decap_4 FILLER_50_1011 ();
 sg13g2_fill_1 FILLER_50_1015 ();
 sg13g2_decap_8 FILLER_50_1025 ();
 sg13g2_decap_8 FILLER_50_1032 ();
 sg13g2_decap_8 FILLER_50_1039 ();
 sg13g2_fill_2 FILLER_50_1046 ();
 sg13g2_fill_1 FILLER_50_1048 ();
 sg13g2_fill_1 FILLER_50_1068 ();
 sg13g2_fill_1 FILLER_50_1082 ();
 sg13g2_decap_8 FILLER_50_1091 ();
 sg13g2_decap_8 FILLER_50_1098 ();
 sg13g2_fill_2 FILLER_50_1105 ();
 sg13g2_fill_1 FILLER_50_1107 ();
 sg13g2_decap_8 FILLER_50_1113 ();
 sg13g2_decap_4 FILLER_50_1120 ();
 sg13g2_decap_8 FILLER_50_1150 ();
 sg13g2_decap_8 FILLER_50_1157 ();
 sg13g2_decap_8 FILLER_50_1164 ();
 sg13g2_decap_8 FILLER_50_1171 ();
 sg13g2_decap_8 FILLER_50_1178 ();
 sg13g2_decap_4 FILLER_50_1185 ();
 sg13g2_fill_2 FILLER_50_1205 ();
 sg13g2_decap_8 FILLER_50_1227 ();
 sg13g2_decap_4 FILLER_50_1234 ();
 sg13g2_fill_2 FILLER_50_1238 ();
 sg13g2_decap_8 FILLER_50_1245 ();
 sg13g2_fill_2 FILLER_50_1252 ();
 sg13g2_fill_1 FILLER_50_1254 ();
 sg13g2_decap_8 FILLER_50_1260 ();
 sg13g2_fill_1 FILLER_50_1267 ();
 sg13g2_fill_2 FILLER_50_1288 ();
 sg13g2_decap_8 FILLER_50_1316 ();
 sg13g2_decap_8 FILLER_50_1341 ();
 sg13g2_decap_4 FILLER_50_1348 ();
 sg13g2_fill_2 FILLER_50_1352 ();
 sg13g2_decap_8 FILLER_50_1359 ();
 sg13g2_decap_8 FILLER_50_1379 ();
 sg13g2_fill_2 FILLER_50_1386 ();
 sg13g2_fill_1 FILLER_50_1388 ();
 sg13g2_decap_8 FILLER_50_1420 ();
 sg13g2_decap_4 FILLER_50_1427 ();
 sg13g2_decap_4 FILLER_50_1434 ();
 sg13g2_fill_2 FILLER_50_1438 ();
 sg13g2_fill_2 FILLER_50_1446 ();
 sg13g2_fill_1 FILLER_50_1448 ();
 sg13g2_decap_8 FILLER_50_1461 ();
 sg13g2_decap_8 FILLER_50_1468 ();
 sg13g2_decap_8 FILLER_50_1475 ();
 sg13g2_decap_8 FILLER_50_1482 ();
 sg13g2_decap_8 FILLER_50_1489 ();
 sg13g2_decap_8 FILLER_50_1496 ();
 sg13g2_decap_8 FILLER_50_1503 ();
 sg13g2_decap_8 FILLER_50_1510 ();
 sg13g2_decap_8 FILLER_50_1517 ();
 sg13g2_fill_1 FILLER_50_1524 ();
 sg13g2_decap_8 FILLER_50_1535 ();
 sg13g2_fill_1 FILLER_50_1542 ();
 sg13g2_decap_8 FILLER_50_1589 ();
 sg13g2_decap_8 FILLER_50_1596 ();
 sg13g2_decap_8 FILLER_50_1603 ();
 sg13g2_decap_8 FILLER_50_1610 ();
 sg13g2_decap_8 FILLER_50_1617 ();
 sg13g2_decap_8 FILLER_50_1624 ();
 sg13g2_decap_8 FILLER_50_1631 ();
 sg13g2_decap_8 FILLER_50_1638 ();
 sg13g2_decap_8 FILLER_50_1650 ();
 sg13g2_decap_8 FILLER_50_1657 ();
 sg13g2_decap_8 FILLER_50_1664 ();
 sg13g2_decap_8 FILLER_50_1671 ();
 sg13g2_decap_8 FILLER_50_1678 ();
 sg13g2_decap_4 FILLER_50_1685 ();
 sg13g2_fill_1 FILLER_50_1689 ();
 sg13g2_decap_4 FILLER_50_1704 ();
 sg13g2_decap_4 FILLER_50_1721 ();
 sg13g2_fill_1 FILLER_50_1725 ();
 sg13g2_decap_8 FILLER_50_1736 ();
 sg13g2_decap_8 FILLER_50_1743 ();
 sg13g2_fill_1 FILLER_50_1750 ();
 sg13g2_decap_8 FILLER_50_1780 ();
 sg13g2_decap_4 FILLER_50_1794 ();
 sg13g2_fill_1 FILLER_50_1798 ();
 sg13g2_decap_8 FILLER_50_1841 ();
 sg13g2_decap_8 FILLER_50_1848 ();
 sg13g2_fill_1 FILLER_50_1855 ();
 sg13g2_decap_8 FILLER_50_1887 ();
 sg13g2_decap_4 FILLER_50_1894 ();
 sg13g2_fill_2 FILLER_50_1898 ();
 sg13g2_fill_2 FILLER_50_1913 ();
 sg13g2_decap_4 FILLER_50_1922 ();
 sg13g2_decap_8 FILLER_50_1943 ();
 sg13g2_decap_8 FILLER_50_1950 ();
 sg13g2_decap_4 FILLER_50_1957 ();
 sg13g2_fill_1 FILLER_50_1983 ();
 sg13g2_decap_8 FILLER_50_1990 ();
 sg13g2_decap_8 FILLER_50_1997 ();
 sg13g2_decap_8 FILLER_50_2004 ();
 sg13g2_decap_4 FILLER_50_2011 ();
 sg13g2_fill_2 FILLER_50_2015 ();
 sg13g2_decap_4 FILLER_50_2054 ();
 sg13g2_fill_1 FILLER_50_2058 ();
 sg13g2_decap_8 FILLER_50_2102 ();
 sg13g2_decap_8 FILLER_50_2109 ();
 sg13g2_decap_8 FILLER_50_2116 ();
 sg13g2_decap_4 FILLER_50_2123 ();
 sg13g2_fill_1 FILLER_50_2127 ();
 sg13g2_decap_8 FILLER_50_2132 ();
 sg13g2_decap_8 FILLER_50_2139 ();
 sg13g2_fill_2 FILLER_50_2146 ();
 sg13g2_fill_1 FILLER_50_2148 ();
 sg13g2_fill_1 FILLER_50_2153 ();
 sg13g2_decap_4 FILLER_50_2158 ();
 sg13g2_decap_8 FILLER_50_2172 ();
 sg13g2_decap_8 FILLER_50_2179 ();
 sg13g2_decap_8 FILLER_50_2186 ();
 sg13g2_decap_8 FILLER_50_2193 ();
 sg13g2_fill_2 FILLER_50_2200 ();
 sg13g2_fill_1 FILLER_50_2202 ();
 sg13g2_fill_1 FILLER_50_2211 ();
 sg13g2_decap_4 FILLER_50_2217 ();
 sg13g2_fill_2 FILLER_50_2221 ();
 sg13g2_decap_8 FILLER_50_2265 ();
 sg13g2_fill_2 FILLER_50_2272 ();
 sg13g2_decap_8 FILLER_50_2290 ();
 sg13g2_decap_8 FILLER_50_2297 ();
 sg13g2_decap_8 FILLER_50_2304 ();
 sg13g2_decap_8 FILLER_50_2311 ();
 sg13g2_decap_8 FILLER_50_2318 ();
 sg13g2_fill_2 FILLER_50_2325 ();
 sg13g2_fill_1 FILLER_50_2327 ();
 sg13g2_decap_8 FILLER_50_2336 ();
 sg13g2_decap_8 FILLER_50_2343 ();
 sg13g2_decap_8 FILLER_50_2350 ();
 sg13g2_decap_8 FILLER_50_2357 ();
 sg13g2_decap_8 FILLER_50_2373 ();
 sg13g2_fill_2 FILLER_50_2380 ();
 sg13g2_decap_8 FILLER_50_2408 ();
 sg13g2_decap_8 FILLER_50_2415 ();
 sg13g2_decap_8 FILLER_50_2422 ();
 sg13g2_decap_8 FILLER_50_2429 ();
 sg13g2_decap_8 FILLER_50_2436 ();
 sg13g2_fill_2 FILLER_50_2443 ();
 sg13g2_decap_8 FILLER_50_2451 ();
 sg13g2_decap_8 FILLER_50_2458 ();
 sg13g2_decap_8 FILLER_50_2465 ();
 sg13g2_decap_8 FILLER_50_2472 ();
 sg13g2_fill_2 FILLER_50_2479 ();
 sg13g2_decap_8 FILLER_50_2485 ();
 sg13g2_decap_8 FILLER_50_2492 ();
 sg13g2_decap_8 FILLER_50_2499 ();
 sg13g2_decap_4 FILLER_50_2506 ();
 sg13g2_fill_2 FILLER_50_2520 ();
 sg13g2_fill_1 FILLER_50_2522 ();
 sg13g2_decap_8 FILLER_50_2554 ();
 sg13g2_decap_8 FILLER_50_2561 ();
 sg13g2_decap_8 FILLER_50_2568 ();
 sg13g2_decap_8 FILLER_50_2575 ();
 sg13g2_decap_8 FILLER_50_2582 ();
 sg13g2_decap_8 FILLER_50_2625 ();
 sg13g2_decap_8 FILLER_50_2632 ();
 sg13g2_decap_8 FILLER_50_2639 ();
 sg13g2_decap_8 FILLER_50_2646 ();
 sg13g2_fill_1 FILLER_50_2653 ();
 sg13g2_decap_8 FILLER_50_2673 ();
 sg13g2_decap_8 FILLER_50_2680 ();
 sg13g2_decap_8 FILLER_50_2687 ();
 sg13g2_decap_8 FILLER_50_2694 ();
 sg13g2_decap_8 FILLER_50_2701 ();
 sg13g2_decap_8 FILLER_50_2708 ();
 sg13g2_decap_8 FILLER_50_2715 ();
 sg13g2_decap_8 FILLER_50_2722 ();
 sg13g2_decap_8 FILLER_50_2729 ();
 sg13g2_decap_8 FILLER_50_2736 ();
 sg13g2_decap_8 FILLER_50_2743 ();
 sg13g2_decap_8 FILLER_50_2769 ();
 sg13g2_decap_8 FILLER_50_2776 ();
 sg13g2_decap_8 FILLER_50_2783 ();
 sg13g2_decap_4 FILLER_50_2790 ();
 sg13g2_fill_2 FILLER_50_2794 ();
 sg13g2_decap_8 FILLER_50_2817 ();
 sg13g2_decap_8 FILLER_50_2824 ();
 sg13g2_decap_4 FILLER_50_2831 ();
 sg13g2_decap_8 FILLER_50_2841 ();
 sg13g2_decap_8 FILLER_50_2854 ();
 sg13g2_fill_2 FILLER_50_2861 ();
 sg13g2_decap_4 FILLER_50_2873 ();
 sg13g2_decap_8 FILLER_50_2903 ();
 sg13g2_decap_8 FILLER_50_2910 ();
 sg13g2_decap_8 FILLER_50_2917 ();
 sg13g2_fill_1 FILLER_50_2924 ();
 sg13g2_decap_8 FILLER_50_2951 ();
 sg13g2_decap_8 FILLER_50_2958 ();
 sg13g2_decap_8 FILLER_50_2965 ();
 sg13g2_decap_8 FILLER_50_2972 ();
 sg13g2_decap_8 FILLER_50_2979 ();
 sg13g2_decap_8 FILLER_50_2986 ();
 sg13g2_decap_8 FILLER_50_2993 ();
 sg13g2_decap_4 FILLER_50_3000 ();
 sg13g2_fill_1 FILLER_50_3004 ();
 sg13g2_fill_2 FILLER_50_3041 ();
 sg13g2_fill_2 FILLER_50_3069 ();
 sg13g2_decap_8 FILLER_50_3107 ();
 sg13g2_decap_8 FILLER_50_3114 ();
 sg13g2_decap_8 FILLER_50_3121 ();
 sg13g2_decap_8 FILLER_50_3128 ();
 sg13g2_decap_8 FILLER_50_3135 ();
 sg13g2_decap_8 FILLER_50_3142 ();
 sg13g2_decap_4 FILLER_50_3149 ();
 sg13g2_fill_1 FILLER_50_3179 ();
 sg13g2_decap_8 FILLER_50_3195 ();
 sg13g2_decap_8 FILLER_50_3202 ();
 sg13g2_decap_8 FILLER_50_3209 ();
 sg13g2_decap_8 FILLER_50_3216 ();
 sg13g2_decap_8 FILLER_50_3223 ();
 sg13g2_decap_8 FILLER_50_3230 ();
 sg13g2_decap_8 FILLER_50_3237 ();
 sg13g2_fill_1 FILLER_50_3244 ();
 sg13g2_decap_8 FILLER_50_3271 ();
 sg13g2_decap_4 FILLER_50_3278 ();
 sg13g2_fill_1 FILLER_50_3282 ();
 sg13g2_decap_8 FILLER_50_3309 ();
 sg13g2_decap_4 FILLER_50_3316 ();
 sg13g2_fill_1 FILLER_50_3330 ();
 sg13g2_fill_1 FILLER_50_3336 ();
 sg13g2_decap_8 FILLER_50_3345 ();
 sg13g2_decap_8 FILLER_50_3352 ();
 sg13g2_decap_8 FILLER_50_3359 ();
 sg13g2_decap_8 FILLER_50_3366 ();
 sg13g2_decap_8 FILLER_50_3373 ();
 sg13g2_decap_8 FILLER_50_3380 ();
 sg13g2_decap_8 FILLER_50_3387 ();
 sg13g2_decap_4 FILLER_50_3394 ();
 sg13g2_fill_1 FILLER_50_3398 ();
 sg13g2_decap_8 FILLER_50_3425 ();
 sg13g2_decap_8 FILLER_50_3432 ();
 sg13g2_decap_8 FILLER_50_3439 ();
 sg13g2_decap_8 FILLER_50_3446 ();
 sg13g2_decap_4 FILLER_50_3453 ();
 sg13g2_decap_8 FILLER_50_3461 ();
 sg13g2_decap_8 FILLER_50_3468 ();
 sg13g2_decap_8 FILLER_50_3475 ();
 sg13g2_fill_1 FILLER_50_3482 ();
 sg13g2_fill_1 FILLER_50_3519 ();
 sg13g2_decap_8 FILLER_50_3525 ();
 sg13g2_decap_4 FILLER_50_3532 ();
 sg13g2_fill_2 FILLER_50_3536 ();
 sg13g2_decap_8 FILLER_50_3569 ();
 sg13g2_decap_4 FILLER_50_3576 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_decap_8 FILLER_51_7 ();
 sg13g2_decap_8 FILLER_51_14 ();
 sg13g2_decap_8 FILLER_51_21 ();
 sg13g2_decap_4 FILLER_51_28 ();
 sg13g2_fill_2 FILLER_51_32 ();
 sg13g2_decap_4 FILLER_51_47 ();
 sg13g2_fill_2 FILLER_51_51 ();
 sg13g2_decap_8 FILLER_51_57 ();
 sg13g2_decap_8 FILLER_51_64 ();
 sg13g2_decap_4 FILLER_51_71 ();
 sg13g2_decap_8 FILLER_51_90 ();
 sg13g2_decap_8 FILLER_51_97 ();
 sg13g2_decap_8 FILLER_51_104 ();
 sg13g2_fill_2 FILLER_51_111 ();
 sg13g2_fill_1 FILLER_51_113 ();
 sg13g2_fill_2 FILLER_51_140 ();
 sg13g2_decap_8 FILLER_51_159 ();
 sg13g2_fill_2 FILLER_51_166 ();
 sg13g2_fill_1 FILLER_51_168 ();
 sg13g2_decap_8 FILLER_51_174 ();
 sg13g2_decap_4 FILLER_51_181 ();
 sg13g2_decap_8 FILLER_51_195 ();
 sg13g2_decap_8 FILLER_51_202 ();
 sg13g2_decap_8 FILLER_51_209 ();
 sg13g2_decap_4 FILLER_51_216 ();
 sg13g2_fill_2 FILLER_51_220 ();
 sg13g2_fill_2 FILLER_51_246 ();
 sg13g2_fill_2 FILLER_51_258 ();
 sg13g2_decap_8 FILLER_51_266 ();
 sg13g2_decap_4 FILLER_51_273 ();
 sg13g2_fill_2 FILLER_51_281 ();
 sg13g2_fill_1 FILLER_51_283 ();
 sg13g2_decap_8 FILLER_51_289 ();
 sg13g2_fill_2 FILLER_51_296 ();
 sg13g2_fill_2 FILLER_51_322 ();
 sg13g2_fill_1 FILLER_51_324 ();
 sg13g2_decap_8 FILLER_51_342 ();
 sg13g2_decap_8 FILLER_51_349 ();
 sg13g2_decap_8 FILLER_51_356 ();
 sg13g2_decap_8 FILLER_51_363 ();
 sg13g2_decap_8 FILLER_51_370 ();
 sg13g2_decap_8 FILLER_51_389 ();
 sg13g2_decap_8 FILLER_51_396 ();
 sg13g2_decap_8 FILLER_51_403 ();
 sg13g2_fill_2 FILLER_51_410 ();
 sg13g2_decap_8 FILLER_51_416 ();
 sg13g2_decap_8 FILLER_51_423 ();
 sg13g2_decap_8 FILLER_51_430 ();
 sg13g2_decap_8 FILLER_51_437 ();
 sg13g2_fill_2 FILLER_51_444 ();
 sg13g2_fill_1 FILLER_51_453 ();
 sg13g2_decap_4 FILLER_51_465 ();
 sg13g2_fill_2 FILLER_51_481 ();
 sg13g2_fill_1 FILLER_51_483 ();
 sg13g2_decap_8 FILLER_51_490 ();
 sg13g2_decap_4 FILLER_51_497 ();
 sg13g2_fill_1 FILLER_51_501 ();
 sg13g2_decap_8 FILLER_51_510 ();
 sg13g2_fill_1 FILLER_51_517 ();
 sg13g2_decap_4 FILLER_51_524 ();
 sg13g2_decap_8 FILLER_51_536 ();
 sg13g2_decap_8 FILLER_51_543 ();
 sg13g2_decap_8 FILLER_51_550 ();
 sg13g2_decap_8 FILLER_51_557 ();
 sg13g2_decap_8 FILLER_51_564 ();
 sg13g2_decap_8 FILLER_51_571 ();
 sg13g2_decap_8 FILLER_51_578 ();
 sg13g2_decap_8 FILLER_51_585 ();
 sg13g2_decap_4 FILLER_51_592 ();
 sg13g2_decap_8 FILLER_51_608 ();
 sg13g2_decap_8 FILLER_51_615 ();
 sg13g2_fill_2 FILLER_51_622 ();
 sg13g2_decap_8 FILLER_51_627 ();
 sg13g2_decap_8 FILLER_51_634 ();
 sg13g2_decap_8 FILLER_51_641 ();
 sg13g2_decap_8 FILLER_51_648 ();
 sg13g2_decap_8 FILLER_51_655 ();
 sg13g2_decap_8 FILLER_51_662 ();
 sg13g2_decap_4 FILLER_51_669 ();
 sg13g2_fill_2 FILLER_51_673 ();
 sg13g2_decap_8 FILLER_51_689 ();
 sg13g2_decap_8 FILLER_51_696 ();
 sg13g2_decap_8 FILLER_51_703 ();
 sg13g2_decap_4 FILLER_51_710 ();
 sg13g2_fill_2 FILLER_51_714 ();
 sg13g2_decap_8 FILLER_51_736 ();
 sg13g2_decap_8 FILLER_51_743 ();
 sg13g2_fill_1 FILLER_51_750 ();
 sg13g2_fill_2 FILLER_51_767 ();
 sg13g2_decap_8 FILLER_51_790 ();
 sg13g2_decap_8 FILLER_51_797 ();
 sg13g2_decap_4 FILLER_51_804 ();
 sg13g2_fill_1 FILLER_51_808 ();
 sg13g2_fill_2 FILLER_51_812 ();
 sg13g2_fill_1 FILLER_51_814 ();
 sg13g2_fill_1 FILLER_51_831 ();
 sg13g2_fill_2 FILLER_51_844 ();
 sg13g2_decap_8 FILLER_51_855 ();
 sg13g2_decap_8 FILLER_51_862 ();
 sg13g2_fill_1 FILLER_51_869 ();
 sg13g2_decap_4 FILLER_51_879 ();
 sg13g2_fill_1 FILLER_51_883 ();
 sg13g2_decap_8 FILLER_51_902 ();
 sg13g2_decap_8 FILLER_51_909 ();
 sg13g2_decap_8 FILLER_51_916 ();
 sg13g2_fill_2 FILLER_51_923 ();
 sg13g2_fill_2 FILLER_51_930 ();
 sg13g2_fill_1 FILLER_51_932 ();
 sg13g2_decap_8 FILLER_51_949 ();
 sg13g2_decap_8 FILLER_51_956 ();
 sg13g2_decap_8 FILLER_51_963 ();
 sg13g2_decap_8 FILLER_51_970 ();
 sg13g2_fill_2 FILLER_51_977 ();
 sg13g2_fill_1 FILLER_51_979 ();
 sg13g2_decap_4 FILLER_51_1006 ();
 sg13g2_decap_8 FILLER_51_1024 ();
 sg13g2_fill_2 FILLER_51_1031 ();
 sg13g2_decap_8 FILLER_51_1085 ();
 sg13g2_fill_2 FILLER_51_1092 ();
 sg13g2_decap_8 FILLER_51_1138 ();
 sg13g2_decap_4 FILLER_51_1145 ();
 sg13g2_fill_2 FILLER_51_1149 ();
 sg13g2_decap_8 FILLER_51_1187 ();
 sg13g2_decap_8 FILLER_51_1194 ();
 sg13g2_decap_8 FILLER_51_1201 ();
 sg13g2_decap_8 FILLER_51_1208 ();
 sg13g2_decap_8 FILLER_51_1215 ();
 sg13g2_fill_2 FILLER_51_1253 ();
 sg13g2_fill_1 FILLER_51_1255 ();
 sg13g2_decap_8 FILLER_51_1269 ();
 sg13g2_fill_2 FILLER_51_1311 ();
 sg13g2_decap_8 FILLER_51_1322 ();
 sg13g2_decap_8 FILLER_51_1329 ();
 sg13g2_decap_8 FILLER_51_1336 ();
 sg13g2_fill_1 FILLER_51_1343 ();
 sg13g2_decap_8 FILLER_51_1354 ();
 sg13g2_decap_8 FILLER_51_1361 ();
 sg13g2_decap_4 FILLER_51_1368 ();
 sg13g2_fill_2 FILLER_51_1372 ();
 sg13g2_decap_8 FILLER_51_1382 ();
 sg13g2_fill_2 FILLER_51_1389 ();
 sg13g2_fill_1 FILLER_51_1391 ();
 sg13g2_decap_8 FILLER_51_1428 ();
 sg13g2_decap_8 FILLER_51_1435 ();
 sg13g2_decap_8 FILLER_51_1442 ();
 sg13g2_fill_2 FILLER_51_1449 ();
 sg13g2_fill_1 FILLER_51_1451 ();
 sg13g2_fill_2 FILLER_51_1458 ();
 sg13g2_fill_2 FILLER_51_1486 ();
 sg13g2_decap_8 FILLER_51_1496 ();
 sg13g2_decap_8 FILLER_51_1503 ();
 sg13g2_decap_8 FILLER_51_1510 ();
 sg13g2_fill_1 FILLER_51_1517 ();
 sg13g2_fill_2 FILLER_51_1528 ();
 sg13g2_fill_1 FILLER_51_1530 ();
 sg13g2_decap_8 FILLER_51_1557 ();
 sg13g2_decap_8 FILLER_51_1564 ();
 sg13g2_decap_8 FILLER_51_1571 ();
 sg13g2_decap_8 FILLER_51_1578 ();
 sg13g2_decap_8 FILLER_51_1598 ();
 sg13g2_decap_8 FILLER_51_1605 ();
 sg13g2_decap_8 FILLER_51_1612 ();
 sg13g2_decap_8 FILLER_51_1619 ();
 sg13g2_decap_8 FILLER_51_1626 ();
 sg13g2_decap_8 FILLER_51_1633 ();
 sg13g2_decap_8 FILLER_51_1640 ();
 sg13g2_decap_8 FILLER_51_1647 ();
 sg13g2_decap_4 FILLER_51_1654 ();
 sg13g2_decap_8 FILLER_51_1674 ();
 sg13g2_decap_8 FILLER_51_1681 ();
 sg13g2_decap_8 FILLER_51_1688 ();
 sg13g2_decap_4 FILLER_51_1695 ();
 sg13g2_fill_1 FILLER_51_1699 ();
 sg13g2_decap_4 FILLER_51_1705 ();
 sg13g2_decap_8 FILLER_51_1717 ();
 sg13g2_fill_2 FILLER_51_1724 ();
 sg13g2_decap_8 FILLER_51_1752 ();
 sg13g2_decap_8 FILLER_51_1759 ();
 sg13g2_decap_8 FILLER_51_1766 ();
 sg13g2_decap_4 FILLER_51_1773 ();
 sg13g2_decap_8 FILLER_51_1780 ();
 sg13g2_fill_2 FILLER_51_1796 ();
 sg13g2_fill_1 FILLER_51_1804 ();
 sg13g2_decap_8 FILLER_51_1844 ();
 sg13g2_decap_8 FILLER_51_1851 ();
 sg13g2_fill_2 FILLER_51_1858 ();
 sg13g2_fill_1 FILLER_51_1860 ();
 sg13g2_decap_8 FILLER_51_1871 ();
 sg13g2_decap_8 FILLER_51_1878 ();
 sg13g2_decap_8 FILLER_51_1885 ();
 sg13g2_decap_8 FILLER_51_1892 ();
 sg13g2_decap_8 FILLER_51_1899 ();
 sg13g2_fill_1 FILLER_51_1906 ();
 sg13g2_fill_1 FILLER_51_1920 ();
 sg13g2_decap_8 FILLER_51_1935 ();
 sg13g2_decap_8 FILLER_51_1942 ();
 sg13g2_decap_8 FILLER_51_1949 ();
 sg13g2_decap_8 FILLER_51_1956 ();
 sg13g2_decap_4 FILLER_51_1963 ();
 sg13g2_fill_2 FILLER_51_1967 ();
 sg13g2_decap_8 FILLER_51_1995 ();
 sg13g2_decap_8 FILLER_51_2002 ();
 sg13g2_decap_8 FILLER_51_2009 ();
 sg13g2_decap_8 FILLER_51_2016 ();
 sg13g2_decap_8 FILLER_51_2045 ();
 sg13g2_decap_8 FILLER_51_2052 ();
 sg13g2_decap_4 FILLER_51_2059 ();
 sg13g2_fill_2 FILLER_51_2063 ();
 sg13g2_decap_8 FILLER_51_2090 ();
 sg13g2_decap_8 FILLER_51_2097 ();
 sg13g2_fill_2 FILLER_51_2104 ();
 sg13g2_fill_1 FILLER_51_2106 ();
 sg13g2_decap_8 FILLER_51_2122 ();
 sg13g2_decap_8 FILLER_51_2129 ();
 sg13g2_decap_8 FILLER_51_2136 ();
 sg13g2_decap_8 FILLER_51_2143 ();
 sg13g2_decap_8 FILLER_51_2150 ();
 sg13g2_decap_4 FILLER_51_2157 ();
 sg13g2_decap_8 FILLER_51_2195 ();
 sg13g2_decap_8 FILLER_51_2202 ();
 sg13g2_decap_8 FILLER_51_2209 ();
 sg13g2_decap_8 FILLER_51_2216 ();
 sg13g2_fill_1 FILLER_51_2223 ();
 sg13g2_fill_1 FILLER_51_2234 ();
 sg13g2_decap_8 FILLER_51_2264 ();
 sg13g2_decap_8 FILLER_51_2271 ();
 sg13g2_decap_8 FILLER_51_2278 ();
 sg13g2_decap_8 FILLER_51_2285 ();
 sg13g2_decap_8 FILLER_51_2292 ();
 sg13g2_decap_8 FILLER_51_2299 ();
 sg13g2_decap_4 FILLER_51_2306 ();
 sg13g2_decap_8 FILLER_51_2341 ();
 sg13g2_decap_8 FILLER_51_2348 ();
 sg13g2_decap_8 FILLER_51_2355 ();
 sg13g2_decap_8 FILLER_51_2362 ();
 sg13g2_decap_4 FILLER_51_2369 ();
 sg13g2_fill_2 FILLER_51_2373 ();
 sg13g2_decap_8 FILLER_51_2401 ();
 sg13g2_decap_8 FILLER_51_2408 ();
 sg13g2_fill_2 FILLER_51_2415 ();
 sg13g2_decap_8 FILLER_51_2422 ();
 sg13g2_fill_1 FILLER_51_2429 ();
 sg13g2_decap_8 FILLER_51_2436 ();
 sg13g2_fill_2 FILLER_51_2443 ();
 sg13g2_fill_1 FILLER_51_2445 ();
 sg13g2_decap_8 FILLER_51_2461 ();
 sg13g2_decap_8 FILLER_51_2482 ();
 sg13g2_decap_8 FILLER_51_2489 ();
 sg13g2_decap_8 FILLER_51_2496 ();
 sg13g2_decap_8 FILLER_51_2503 ();
 sg13g2_decap_8 FILLER_51_2510 ();
 sg13g2_fill_2 FILLER_51_2517 ();
 sg13g2_fill_2 FILLER_51_2529 ();
 sg13g2_decap_8 FILLER_51_2557 ();
 sg13g2_decap_8 FILLER_51_2564 ();
 sg13g2_decap_8 FILLER_51_2571 ();
 sg13g2_decap_8 FILLER_51_2578 ();
 sg13g2_decap_4 FILLER_51_2585 ();
 sg13g2_fill_2 FILLER_51_2589 ();
 sg13g2_decap_8 FILLER_51_2627 ();
 sg13g2_decap_8 FILLER_51_2634 ();
 sg13g2_decap_8 FILLER_51_2641 ();
 sg13g2_decap_8 FILLER_51_2648 ();
 sg13g2_decap_8 FILLER_51_2655 ();
 sg13g2_decap_8 FILLER_51_2680 ();
 sg13g2_decap_8 FILLER_51_2687 ();
 sg13g2_decap_8 FILLER_51_2723 ();
 sg13g2_decap_8 FILLER_51_2730 ();
 sg13g2_fill_2 FILLER_51_2737 ();
 sg13g2_fill_1 FILLER_51_2739 ();
 sg13g2_decap_8 FILLER_51_2746 ();
 sg13g2_fill_2 FILLER_51_2753 ();
 sg13g2_decap_8 FILLER_51_2771 ();
 sg13g2_decap_8 FILLER_51_2778 ();
 sg13g2_decap_8 FILLER_51_2785 ();
 sg13g2_decap_8 FILLER_51_2792 ();
 sg13g2_decap_8 FILLER_51_2799 ();
 sg13g2_decap_8 FILLER_51_2806 ();
 sg13g2_fill_1 FILLER_51_2813 ();
 sg13g2_fill_1 FILLER_51_2820 ();
 sg13g2_fill_2 FILLER_51_2833 ();
 sg13g2_decap_8 FILLER_51_2841 ();
 sg13g2_decap_8 FILLER_51_2848 ();
 sg13g2_decap_8 FILLER_51_2855 ();
 sg13g2_decap_8 FILLER_51_2898 ();
 sg13g2_decap_8 FILLER_51_2905 ();
 sg13g2_fill_1 FILLER_51_2912 ();
 sg13g2_decap_8 FILLER_51_2949 ();
 sg13g2_decap_8 FILLER_51_2956 ();
 sg13g2_decap_8 FILLER_51_2963 ();
 sg13g2_decap_4 FILLER_51_2970 ();
 sg13g2_fill_1 FILLER_51_2974 ();
 sg13g2_decap_8 FILLER_51_3001 ();
 sg13g2_decap_8 FILLER_51_3008 ();
 sg13g2_decap_8 FILLER_51_3015 ();
 sg13g2_decap_4 FILLER_51_3022 ();
 sg13g2_fill_2 FILLER_51_3026 ();
 sg13g2_decap_8 FILLER_51_3038 ();
 sg13g2_decap_8 FILLER_51_3045 ();
 sg13g2_fill_2 FILLER_51_3052 ();
 sg13g2_decap_8 FILLER_51_3058 ();
 sg13g2_decap_8 FILLER_51_3065 ();
 sg13g2_decap_8 FILLER_51_3072 ();
 sg13g2_fill_2 FILLER_51_3079 ();
 sg13g2_fill_1 FILLER_51_3081 ();
 sg13g2_decap_8 FILLER_51_3103 ();
 sg13g2_decap_8 FILLER_51_3110 ();
 sg13g2_decap_8 FILLER_51_3117 ();
 sg13g2_decap_8 FILLER_51_3124 ();
 sg13g2_decap_8 FILLER_51_3131 ();
 sg13g2_decap_8 FILLER_51_3138 ();
 sg13g2_fill_1 FILLER_51_3145 ();
 sg13g2_decap_8 FILLER_51_3151 ();
 sg13g2_fill_1 FILLER_51_3158 ();
 sg13g2_decap_8 FILLER_51_3164 ();
 sg13g2_decap_8 FILLER_51_3171 ();
 sg13g2_decap_4 FILLER_51_3178 ();
 sg13g2_fill_2 FILLER_51_3197 ();
 sg13g2_fill_1 FILLER_51_3199 ();
 sg13g2_decap_8 FILLER_51_3226 ();
 sg13g2_decap_4 FILLER_51_3233 ();
 sg13g2_fill_1 FILLER_51_3237 ();
 sg13g2_decap_8 FILLER_51_3264 ();
 sg13g2_decap_8 FILLER_51_3271 ();
 sg13g2_decap_4 FILLER_51_3278 ();
 sg13g2_fill_1 FILLER_51_3282 ();
 sg13g2_decap_8 FILLER_51_3293 ();
 sg13g2_decap_8 FILLER_51_3300 ();
 sg13g2_decap_8 FILLER_51_3307 ();
 sg13g2_decap_8 FILLER_51_3314 ();
 sg13g2_decap_8 FILLER_51_3321 ();
 sg13g2_fill_2 FILLER_51_3328 ();
 sg13g2_decap_8 FILLER_51_3345 ();
 sg13g2_decap_8 FILLER_51_3352 ();
 sg13g2_decap_8 FILLER_51_3359 ();
 sg13g2_decap_8 FILLER_51_3366 ();
 sg13g2_decap_8 FILLER_51_3373 ();
 sg13g2_decap_8 FILLER_51_3380 ();
 sg13g2_decap_4 FILLER_51_3387 ();
 sg13g2_fill_2 FILLER_51_3391 ();
 sg13g2_fill_2 FILLER_51_3403 ();
 sg13g2_decap_8 FILLER_51_3431 ();
 sg13g2_decap_8 FILLER_51_3438 ();
 sg13g2_decap_4 FILLER_51_3445 ();
 sg13g2_decap_4 FILLER_51_3454 ();
 sg13g2_fill_2 FILLER_51_3458 ();
 sg13g2_decap_8 FILLER_51_3496 ();
 sg13g2_decap_8 FILLER_51_3513 ();
 sg13g2_decap_8 FILLER_51_3520 ();
 sg13g2_decap_4 FILLER_51_3527 ();
 sg13g2_fill_2 FILLER_51_3531 ();
 sg13g2_decap_8 FILLER_51_3569 ();
 sg13g2_decap_4 FILLER_51_3576 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_decap_8 FILLER_52_7 ();
 sg13g2_decap_8 FILLER_52_14 ();
 sg13g2_decap_4 FILLER_52_21 ();
 sg13g2_fill_1 FILLER_52_25 ();
 sg13g2_fill_2 FILLER_52_31 ();
 sg13g2_fill_1 FILLER_52_33 ();
 sg13g2_decap_4 FILLER_52_43 ();
 sg13g2_decap_8 FILLER_52_51 ();
 sg13g2_decap_8 FILLER_52_58 ();
 sg13g2_decap_8 FILLER_52_65 ();
 sg13g2_decap_8 FILLER_52_72 ();
 sg13g2_decap_8 FILLER_52_79 ();
 sg13g2_decap_8 FILLER_52_86 ();
 sg13g2_decap_8 FILLER_52_93 ();
 sg13g2_decap_8 FILLER_52_100 ();
 sg13g2_decap_8 FILLER_52_107 ();
 sg13g2_decap_8 FILLER_52_114 ();
 sg13g2_fill_2 FILLER_52_121 ();
 sg13g2_fill_1 FILLER_52_123 ();
 sg13g2_decap_8 FILLER_52_132 ();
 sg13g2_fill_1 FILLER_52_139 ();
 sg13g2_decap_8 FILLER_52_143 ();
 sg13g2_decap_8 FILLER_52_150 ();
 sg13g2_fill_2 FILLER_52_157 ();
 sg13g2_fill_1 FILLER_52_159 ();
 sg13g2_decap_8 FILLER_52_171 ();
 sg13g2_decap_8 FILLER_52_178 ();
 sg13g2_fill_2 FILLER_52_185 ();
 sg13g2_decap_8 FILLER_52_204 ();
 sg13g2_decap_8 FILLER_52_211 ();
 sg13g2_fill_1 FILLER_52_230 ();
 sg13g2_fill_2 FILLER_52_247 ();
 sg13g2_decap_8 FILLER_52_265 ();
 sg13g2_decap_8 FILLER_52_280 ();
 sg13g2_fill_2 FILLER_52_287 ();
 sg13g2_decap_8 FILLER_52_299 ();
 sg13g2_decap_4 FILLER_52_306 ();
 sg13g2_fill_2 FILLER_52_310 ();
 sg13g2_decap_8 FILLER_52_317 ();
 sg13g2_fill_2 FILLER_52_324 ();
 sg13g2_decap_8 FILLER_52_334 ();
 sg13g2_decap_8 FILLER_52_341 ();
 sg13g2_decap_8 FILLER_52_348 ();
 sg13g2_decap_8 FILLER_52_355 ();
 sg13g2_decap_8 FILLER_52_362 ();
 sg13g2_decap_8 FILLER_52_369 ();
 sg13g2_decap_8 FILLER_52_376 ();
 sg13g2_decap_8 FILLER_52_383 ();
 sg13g2_decap_8 FILLER_52_390 ();
 sg13g2_decap_8 FILLER_52_397 ();
 sg13g2_decap_8 FILLER_52_404 ();
 sg13g2_decap_8 FILLER_52_411 ();
 sg13g2_decap_8 FILLER_52_418 ();
 sg13g2_decap_8 FILLER_52_425 ();
 sg13g2_decap_4 FILLER_52_432 ();
 sg13g2_fill_1 FILLER_52_436 ();
 sg13g2_decap_8 FILLER_52_452 ();
 sg13g2_decap_8 FILLER_52_459 ();
 sg13g2_decap_8 FILLER_52_466 ();
 sg13g2_decap_8 FILLER_52_479 ();
 sg13g2_decap_8 FILLER_52_486 ();
 sg13g2_decap_8 FILLER_52_493 ();
 sg13g2_decap_8 FILLER_52_500 ();
 sg13g2_decap_8 FILLER_52_507 ();
 sg13g2_fill_1 FILLER_52_514 ();
 sg13g2_decap_8 FILLER_52_544 ();
 sg13g2_decap_8 FILLER_52_551 ();
 sg13g2_decap_8 FILLER_52_558 ();
 sg13g2_decap_8 FILLER_52_565 ();
 sg13g2_decap_8 FILLER_52_572 ();
 sg13g2_decap_4 FILLER_52_579 ();
 sg13g2_fill_2 FILLER_52_583 ();
 sg13g2_decap_4 FILLER_52_593 ();
 sg13g2_fill_2 FILLER_52_597 ();
 sg13g2_decap_8 FILLER_52_607 ();
 sg13g2_decap_8 FILLER_52_614 ();
 sg13g2_fill_2 FILLER_52_621 ();
 sg13g2_decap_8 FILLER_52_637 ();
 sg13g2_fill_1 FILLER_52_644 ();
 sg13g2_decap_8 FILLER_52_666 ();
 sg13g2_fill_1 FILLER_52_673 ();
 sg13g2_decap_8 FILLER_52_686 ();
 sg13g2_decap_8 FILLER_52_693 ();
 sg13g2_decap_8 FILLER_52_700 ();
 sg13g2_decap_8 FILLER_52_707 ();
 sg13g2_decap_8 FILLER_52_714 ();
 sg13g2_decap_4 FILLER_52_721 ();
 sg13g2_fill_1 FILLER_52_725 ();
 sg13g2_decap_8 FILLER_52_730 ();
 sg13g2_decap_8 FILLER_52_737 ();
 sg13g2_decap_8 FILLER_52_744 ();
 sg13g2_decap_8 FILLER_52_751 ();
 sg13g2_decap_8 FILLER_52_758 ();
 sg13g2_decap_8 FILLER_52_765 ();
 sg13g2_decap_8 FILLER_52_772 ();
 sg13g2_decap_8 FILLER_52_779 ();
 sg13g2_decap_8 FILLER_52_786 ();
 sg13g2_decap_8 FILLER_52_793 ();
 sg13g2_decap_8 FILLER_52_800 ();
 sg13g2_fill_1 FILLER_52_807 ();
 sg13g2_decap_4 FILLER_52_824 ();
 sg13g2_decap_8 FILLER_52_848 ();
 sg13g2_decap_8 FILLER_52_855 ();
 sg13g2_decap_4 FILLER_52_862 ();
 sg13g2_fill_1 FILLER_52_866 ();
 sg13g2_fill_2 FILLER_52_893 ();
 sg13g2_decap_8 FILLER_52_902 ();
 sg13g2_decap_8 FILLER_52_909 ();
 sg13g2_fill_2 FILLER_52_916 ();
 sg13g2_fill_1 FILLER_52_918 ();
 sg13g2_decap_8 FILLER_52_961 ();
 sg13g2_decap_8 FILLER_52_968 ();
 sg13g2_fill_1 FILLER_52_989 ();
 sg13g2_decap_8 FILLER_52_1039 ();
 sg13g2_decap_4 FILLER_52_1046 ();
 sg13g2_fill_1 FILLER_52_1050 ();
 sg13g2_fill_2 FILLER_52_1060 ();
 sg13g2_fill_1 FILLER_52_1062 ();
 sg13g2_decap_8 FILLER_52_1068 ();
 sg13g2_decap_8 FILLER_52_1075 ();
 sg13g2_decap_8 FILLER_52_1082 ();
 sg13g2_decap_8 FILLER_52_1089 ();
 sg13g2_decap_8 FILLER_52_1096 ();
 sg13g2_decap_8 FILLER_52_1103 ();
 sg13g2_decap_8 FILLER_52_1110 ();
 sg13g2_decap_8 FILLER_52_1125 ();
 sg13g2_decap_8 FILLER_52_1132 ();
 sg13g2_decap_8 FILLER_52_1139 ();
 sg13g2_decap_4 FILLER_52_1146 ();
 sg13g2_fill_1 FILLER_52_1150 ();
 sg13g2_decap_8 FILLER_52_1182 ();
 sg13g2_decap_8 FILLER_52_1189 ();
 sg13g2_decap_8 FILLER_52_1196 ();
 sg13g2_decap_8 FILLER_52_1203 ();
 sg13g2_decap_8 FILLER_52_1210 ();
 sg13g2_decap_8 FILLER_52_1217 ();
 sg13g2_decap_8 FILLER_52_1224 ();
 sg13g2_decap_8 FILLER_52_1231 ();
 sg13g2_decap_8 FILLER_52_1238 ();
 sg13g2_decap_8 FILLER_52_1245 ();
 sg13g2_decap_4 FILLER_52_1252 ();
 sg13g2_fill_2 FILLER_52_1260 ();
 sg13g2_decap_4 FILLER_52_1270 ();
 sg13g2_fill_2 FILLER_52_1274 ();
 sg13g2_decap_8 FILLER_52_1281 ();
 sg13g2_fill_2 FILLER_52_1288 ();
 sg13g2_fill_1 FILLER_52_1290 ();
 sg13g2_decap_4 FILLER_52_1298 ();
 sg13g2_decap_8 FILLER_52_1311 ();
 sg13g2_decap_8 FILLER_52_1318 ();
 sg13g2_decap_8 FILLER_52_1325 ();
 sg13g2_decap_8 FILLER_52_1332 ();
 sg13g2_decap_8 FILLER_52_1339 ();
 sg13g2_decap_8 FILLER_52_1372 ();
 sg13g2_decap_8 FILLER_52_1379 ();
 sg13g2_decap_4 FILLER_52_1386 ();
 sg13g2_fill_1 FILLER_52_1390 ();
 sg13g2_decap_8 FILLER_52_1394 ();
 sg13g2_decap_8 FILLER_52_1401 ();
 sg13g2_decap_8 FILLER_52_1408 ();
 sg13g2_decap_8 FILLER_52_1415 ();
 sg13g2_decap_8 FILLER_52_1422 ();
 sg13g2_decap_8 FILLER_52_1429 ();
 sg13g2_decap_8 FILLER_52_1436 ();
 sg13g2_decap_8 FILLER_52_1443 ();
 sg13g2_decap_8 FILLER_52_1470 ();
 sg13g2_decap_8 FILLER_52_1477 ();
 sg13g2_decap_8 FILLER_52_1484 ();
 sg13g2_decap_8 FILLER_52_1491 ();
 sg13g2_decap_8 FILLER_52_1498 ();
 sg13g2_decap_8 FILLER_52_1505 ();
 sg13g2_fill_2 FILLER_52_1512 ();
 sg13g2_decap_8 FILLER_52_1520 ();
 sg13g2_decap_8 FILLER_52_1527 ();
 sg13g2_fill_2 FILLER_52_1534 ();
 sg13g2_decap_8 FILLER_52_1562 ();
 sg13g2_decap_8 FILLER_52_1569 ();
 sg13g2_decap_8 FILLER_52_1576 ();
 sg13g2_fill_1 FILLER_52_1583 ();
 sg13g2_fill_2 FILLER_52_1603 ();
 sg13g2_fill_1 FILLER_52_1605 ();
 sg13g2_decap_8 FILLER_52_1637 ();
 sg13g2_decap_8 FILLER_52_1644 ();
 sg13g2_fill_2 FILLER_52_1651 ();
 sg13g2_fill_1 FILLER_52_1653 ();
 sg13g2_decap_8 FILLER_52_1686 ();
 sg13g2_decap_8 FILLER_52_1693 ();
 sg13g2_decap_8 FILLER_52_1700 ();
 sg13g2_decap_8 FILLER_52_1707 ();
 sg13g2_decap_8 FILLER_52_1714 ();
 sg13g2_decap_8 FILLER_52_1721 ();
 sg13g2_fill_2 FILLER_52_1728 ();
 sg13g2_decap_8 FILLER_52_1740 ();
 sg13g2_decap_8 FILLER_52_1747 ();
 sg13g2_decap_8 FILLER_52_1754 ();
 sg13g2_decap_8 FILLER_52_1761 ();
 sg13g2_decap_4 FILLER_52_1768 ();
 sg13g2_fill_2 FILLER_52_1772 ();
 sg13g2_fill_1 FILLER_52_1786 ();
 sg13g2_fill_2 FILLER_52_1799 ();
 sg13g2_fill_1 FILLER_52_1804 ();
 sg13g2_decap_8 FILLER_52_1811 ();
 sg13g2_decap_8 FILLER_52_1818 ();
 sg13g2_decap_8 FILLER_52_1825 ();
 sg13g2_decap_8 FILLER_52_1832 ();
 sg13g2_decap_8 FILLER_52_1839 ();
 sg13g2_decap_8 FILLER_52_1846 ();
 sg13g2_decap_8 FILLER_52_1853 ();
 sg13g2_decap_4 FILLER_52_1860 ();
 sg13g2_fill_1 FILLER_52_1864 ();
 sg13g2_decap_8 FILLER_52_1876 ();
 sg13g2_decap_8 FILLER_52_1883 ();
 sg13g2_decap_8 FILLER_52_1890 ();
 sg13g2_decap_8 FILLER_52_1897 ();
 sg13g2_decap_8 FILLER_52_1904 ();
 sg13g2_decap_8 FILLER_52_1911 ();
 sg13g2_fill_2 FILLER_52_1918 ();
 sg13g2_decap_8 FILLER_52_1928 ();
 sg13g2_decap_8 FILLER_52_1935 ();
 sg13g2_decap_8 FILLER_52_1942 ();
 sg13g2_decap_8 FILLER_52_1949 ();
 sg13g2_decap_8 FILLER_52_1956 ();
 sg13g2_decap_4 FILLER_52_1963 ();
 sg13g2_fill_1 FILLER_52_1967 ();
 sg13g2_decap_8 FILLER_52_1978 ();
 sg13g2_decap_8 FILLER_52_1985 ();
 sg13g2_decap_8 FILLER_52_1992 ();
 sg13g2_decap_8 FILLER_52_1999 ();
 sg13g2_decap_8 FILLER_52_2006 ();
 sg13g2_decap_8 FILLER_52_2013 ();
 sg13g2_decap_8 FILLER_52_2020 ();
 sg13g2_decap_4 FILLER_52_2027 ();
 sg13g2_decap_8 FILLER_52_2041 ();
 sg13g2_decap_8 FILLER_52_2048 ();
 sg13g2_decap_8 FILLER_52_2055 ();
 sg13g2_decap_8 FILLER_52_2062 ();
 sg13g2_decap_4 FILLER_52_2069 ();
 sg13g2_decap_8 FILLER_52_2079 ();
 sg13g2_decap_8 FILLER_52_2086 ();
 sg13g2_decap_8 FILLER_52_2093 ();
 sg13g2_decap_8 FILLER_52_2100 ();
 sg13g2_decap_8 FILLER_52_2107 ();
 sg13g2_decap_8 FILLER_52_2114 ();
 sg13g2_decap_8 FILLER_52_2121 ();
 sg13g2_fill_1 FILLER_52_2128 ();
 sg13g2_decap_8 FILLER_52_2139 ();
 sg13g2_decap_8 FILLER_52_2146 ();
 sg13g2_decap_8 FILLER_52_2153 ();
 sg13g2_decap_8 FILLER_52_2160 ();
 sg13g2_decap_8 FILLER_52_2167 ();
 sg13g2_decap_8 FILLER_52_2174 ();
 sg13g2_decap_8 FILLER_52_2181 ();
 sg13g2_decap_8 FILLER_52_2188 ();
 sg13g2_decap_4 FILLER_52_2195 ();
 sg13g2_fill_2 FILLER_52_2199 ();
 sg13g2_decap_8 FILLER_52_2211 ();
 sg13g2_decap_8 FILLER_52_2218 ();
 sg13g2_fill_1 FILLER_52_2225 ();
 sg13g2_fill_1 FILLER_52_2244 ();
 sg13g2_decap_8 FILLER_52_2253 ();
 sg13g2_decap_8 FILLER_52_2260 ();
 sg13g2_decap_8 FILLER_52_2267 ();
 sg13g2_decap_8 FILLER_52_2274 ();
 sg13g2_decap_8 FILLER_52_2281 ();
 sg13g2_decap_8 FILLER_52_2288 ();
 sg13g2_decap_8 FILLER_52_2295 ();
 sg13g2_decap_4 FILLER_52_2302 ();
 sg13g2_decap_8 FILLER_52_2316 ();
 sg13g2_decap_8 FILLER_52_2323 ();
 sg13g2_decap_8 FILLER_52_2330 ();
 sg13g2_decap_8 FILLER_52_2337 ();
 sg13g2_decap_8 FILLER_52_2344 ();
 sg13g2_decap_8 FILLER_52_2351 ();
 sg13g2_decap_8 FILLER_52_2358 ();
 sg13g2_decap_8 FILLER_52_2365 ();
 sg13g2_fill_2 FILLER_52_2372 ();
 sg13g2_decap_8 FILLER_52_2394 ();
 sg13g2_decap_8 FILLER_52_2401 ();
 sg13g2_decap_8 FILLER_52_2408 ();
 sg13g2_decap_8 FILLER_52_2415 ();
 sg13g2_decap_8 FILLER_52_2422 ();
 sg13g2_decap_8 FILLER_52_2429 ();
 sg13g2_fill_2 FILLER_52_2436 ();
 sg13g2_fill_1 FILLER_52_2452 ();
 sg13g2_decap_8 FILLER_52_2470 ();
 sg13g2_decap_8 FILLER_52_2477 ();
 sg13g2_fill_1 FILLER_52_2484 ();
 sg13g2_decap_8 FILLER_52_2495 ();
 sg13g2_decap_8 FILLER_52_2502 ();
 sg13g2_decap_8 FILLER_52_2509 ();
 sg13g2_decap_8 FILLER_52_2516 ();
 sg13g2_decap_8 FILLER_52_2523 ();
 sg13g2_fill_1 FILLER_52_2530 ();
 sg13g2_decap_8 FILLER_52_2536 ();
 sg13g2_decap_8 FILLER_52_2543 ();
 sg13g2_decap_8 FILLER_52_2550 ();
 sg13g2_decap_4 FILLER_52_2557 ();
 sg13g2_fill_1 FILLER_52_2561 ();
 sg13g2_decap_8 FILLER_52_2570 ();
 sg13g2_decap_8 FILLER_52_2577 ();
 sg13g2_decap_8 FILLER_52_2584 ();
 sg13g2_decap_8 FILLER_52_2591 ();
 sg13g2_decap_8 FILLER_52_2598 ();
 sg13g2_decap_8 FILLER_52_2605 ();
 sg13g2_decap_8 FILLER_52_2612 ();
 sg13g2_decap_8 FILLER_52_2619 ();
 sg13g2_decap_8 FILLER_52_2626 ();
 sg13g2_fill_2 FILLER_52_2633 ();
 sg13g2_fill_1 FILLER_52_2635 ();
 sg13g2_decap_8 FILLER_52_2640 ();
 sg13g2_decap_8 FILLER_52_2647 ();
 sg13g2_fill_2 FILLER_52_2654 ();
 sg13g2_decap_4 FILLER_52_2675 ();
 sg13g2_decap_4 FILLER_52_2687 ();
 sg13g2_fill_2 FILLER_52_2691 ();
 sg13g2_decap_8 FILLER_52_2699 ();
 sg13g2_fill_2 FILLER_52_2706 ();
 sg13g2_fill_1 FILLER_52_2708 ();
 sg13g2_decap_8 FILLER_52_2735 ();
 sg13g2_decap_8 FILLER_52_2742 ();
 sg13g2_decap_8 FILLER_52_2749 ();
 sg13g2_decap_8 FILLER_52_2756 ();
 sg13g2_decap_8 FILLER_52_2763 ();
 sg13g2_fill_2 FILLER_52_2770 ();
 sg13g2_decap_8 FILLER_52_2780 ();
 sg13g2_decap_8 FILLER_52_2787 ();
 sg13g2_decap_4 FILLER_52_2794 ();
 sg13g2_fill_1 FILLER_52_2798 ();
 sg13g2_decap_8 FILLER_52_2812 ();
 sg13g2_decap_8 FILLER_52_2819 ();
 sg13g2_fill_1 FILLER_52_2826 ();
 sg13g2_fill_2 FILLER_52_2833 ();
 sg13g2_fill_1 FILLER_52_2838 ();
 sg13g2_decap_8 FILLER_52_2847 ();
 sg13g2_decap_8 FILLER_52_2854 ();
 sg13g2_decap_8 FILLER_52_2861 ();
 sg13g2_decap_8 FILLER_52_2868 ();
 sg13g2_decap_8 FILLER_52_2875 ();
 sg13g2_decap_8 FILLER_52_2882 ();
 sg13g2_decap_8 FILLER_52_2889 ();
 sg13g2_decap_8 FILLER_52_2896 ();
 sg13g2_decap_8 FILLER_52_2903 ();
 sg13g2_decap_8 FILLER_52_2910 ();
 sg13g2_fill_2 FILLER_52_2917 ();
 sg13g2_decap_8 FILLER_52_2929 ();
 sg13g2_decap_8 FILLER_52_2936 ();
 sg13g2_decap_8 FILLER_52_2943 ();
 sg13g2_decap_4 FILLER_52_2950 ();
 sg13g2_fill_1 FILLER_52_2954 ();
 sg13g2_decap_8 FILLER_52_2969 ();
 sg13g2_decap_8 FILLER_52_3002 ();
 sg13g2_decap_8 FILLER_52_3009 ();
 sg13g2_decap_8 FILLER_52_3016 ();
 sg13g2_decap_8 FILLER_52_3023 ();
 sg13g2_decap_8 FILLER_52_3030 ();
 sg13g2_decap_8 FILLER_52_3037 ();
 sg13g2_decap_8 FILLER_52_3044 ();
 sg13g2_decap_8 FILLER_52_3051 ();
 sg13g2_decap_8 FILLER_52_3058 ();
 sg13g2_decap_8 FILLER_52_3065 ();
 sg13g2_decap_8 FILLER_52_3072 ();
 sg13g2_fill_2 FILLER_52_3079 ();
 sg13g2_decap_8 FILLER_52_3111 ();
 sg13g2_decap_8 FILLER_52_3118 ();
 sg13g2_decap_8 FILLER_52_3125 ();
 sg13g2_decap_8 FILLER_52_3132 ();
 sg13g2_decap_8 FILLER_52_3139 ();
 sg13g2_decap_4 FILLER_52_3146 ();
 sg13g2_decap_4 FILLER_52_3155 ();
 sg13g2_fill_1 FILLER_52_3159 ();
 sg13g2_decap_8 FILLER_52_3170 ();
 sg13g2_decap_8 FILLER_52_3177 ();
 sg13g2_decap_8 FILLER_52_3184 ();
 sg13g2_decap_8 FILLER_52_3217 ();
 sg13g2_decap_8 FILLER_52_3224 ();
 sg13g2_decap_8 FILLER_52_3231 ();
 sg13g2_decap_4 FILLER_52_3238 ();
 sg13g2_decap_8 FILLER_52_3252 ();
 sg13g2_decap_8 FILLER_52_3259 ();
 sg13g2_decap_8 FILLER_52_3266 ();
 sg13g2_decap_8 FILLER_52_3273 ();
 sg13g2_fill_1 FILLER_52_3280 ();
 sg13g2_decap_8 FILLER_52_3307 ();
 sg13g2_decap_8 FILLER_52_3314 ();
 sg13g2_decap_8 FILLER_52_3321 ();
 sg13g2_decap_8 FILLER_52_3354 ();
 sg13g2_decap_8 FILLER_52_3361 ();
 sg13g2_decap_8 FILLER_52_3368 ();
 sg13g2_decap_8 FILLER_52_3375 ();
 sg13g2_decap_8 FILLER_52_3382 ();
 sg13g2_decap_8 FILLER_52_3389 ();
 sg13g2_fill_1 FILLER_52_3396 ();
 sg13g2_fill_1 FILLER_52_3407 ();
 sg13g2_decap_8 FILLER_52_3433 ();
 sg13g2_decap_8 FILLER_52_3440 ();
 sg13g2_decap_8 FILLER_52_3447 ();
 sg13g2_decap_8 FILLER_52_3454 ();
 sg13g2_fill_2 FILLER_52_3461 ();
 sg13g2_fill_1 FILLER_52_3463 ();
 sg13g2_decap_8 FILLER_52_3468 ();
 sg13g2_decap_8 FILLER_52_3475 ();
 sg13g2_decap_8 FILLER_52_3482 ();
 sg13g2_decap_8 FILLER_52_3489 ();
 sg13g2_fill_2 FILLER_52_3496 ();
 sg13g2_fill_1 FILLER_52_3513 ();
 sg13g2_decap_8 FILLER_52_3518 ();
 sg13g2_decap_8 FILLER_52_3525 ();
 sg13g2_fill_2 FILLER_52_3532 ();
 sg13g2_fill_1 FILLER_52_3534 ();
 sg13g2_decap_8 FILLER_52_3545 ();
 sg13g2_decap_8 FILLER_52_3552 ();
 sg13g2_decap_8 FILLER_52_3559 ();
 sg13g2_decap_8 FILLER_52_3566 ();
 sg13g2_decap_8 FILLER_52_3573 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_decap_4 FILLER_53_7 ();
 sg13g2_fill_1 FILLER_53_11 ();
 sg13g2_fill_2 FILLER_53_59 ();
 sg13g2_fill_1 FILLER_53_61 ();
 sg13g2_decap_4 FILLER_53_67 ();
 sg13g2_decap_8 FILLER_53_81 ();
 sg13g2_fill_1 FILLER_53_88 ();
 sg13g2_decap_8 FILLER_53_93 ();
 sg13g2_decap_8 FILLER_53_100 ();
 sg13g2_decap_8 FILLER_53_107 ();
 sg13g2_decap_8 FILLER_53_114 ();
 sg13g2_decap_8 FILLER_53_121 ();
 sg13g2_decap_4 FILLER_53_128 ();
 sg13g2_fill_1 FILLER_53_132 ();
 sg13g2_fill_2 FILLER_53_164 ();
 sg13g2_fill_1 FILLER_53_166 ();
 sg13g2_fill_1 FILLER_53_181 ();
 sg13g2_decap_4 FILLER_53_226 ();
 sg13g2_fill_2 FILLER_53_243 ();
 sg13g2_fill_1 FILLER_53_245 ();
 sg13g2_decap_8 FILLER_53_258 ();
 sg13g2_decap_8 FILLER_53_265 ();
 sg13g2_decap_8 FILLER_53_272 ();
 sg13g2_decap_8 FILLER_53_279 ();
 sg13g2_decap_8 FILLER_53_286 ();
 sg13g2_decap_8 FILLER_53_293 ();
 sg13g2_decap_8 FILLER_53_300 ();
 sg13g2_decap_8 FILLER_53_307 ();
 sg13g2_decap_8 FILLER_53_314 ();
 sg13g2_decap_8 FILLER_53_321 ();
 sg13g2_decap_8 FILLER_53_328 ();
 sg13g2_decap_8 FILLER_53_335 ();
 sg13g2_fill_2 FILLER_53_350 ();
 sg13g2_decap_8 FILLER_53_361 ();
 sg13g2_decap_8 FILLER_53_368 ();
 sg13g2_decap_8 FILLER_53_375 ();
 sg13g2_decap_8 FILLER_53_382 ();
 sg13g2_decap_8 FILLER_53_389 ();
 sg13g2_decap_8 FILLER_53_396 ();
 sg13g2_fill_2 FILLER_53_403 ();
 sg13g2_fill_1 FILLER_53_405 ();
 sg13g2_decap_8 FILLER_53_436 ();
 sg13g2_fill_2 FILLER_53_443 ();
 sg13g2_fill_1 FILLER_53_445 ();
 sg13g2_decap_4 FILLER_53_449 ();
 sg13g2_fill_1 FILLER_53_453 ();
 sg13g2_decap_8 FILLER_53_460 ();
 sg13g2_decap_8 FILLER_53_467 ();
 sg13g2_decap_8 FILLER_53_474 ();
 sg13g2_decap_8 FILLER_53_486 ();
 sg13g2_decap_8 FILLER_53_493 ();
 sg13g2_decap_8 FILLER_53_500 ();
 sg13g2_decap_8 FILLER_53_507 ();
 sg13g2_decap_4 FILLER_53_514 ();
 sg13g2_decap_8 FILLER_53_521 ();
 sg13g2_fill_2 FILLER_53_528 ();
 sg13g2_decap_8 FILLER_53_556 ();
 sg13g2_decap_8 FILLER_53_563 ();
 sg13g2_decap_8 FILLER_53_570 ();
 sg13g2_decap_8 FILLER_53_577 ();
 sg13g2_decap_8 FILLER_53_584 ();
 sg13g2_fill_2 FILLER_53_591 ();
 sg13g2_fill_1 FILLER_53_593 ();
 sg13g2_decap_8 FILLER_53_615 ();
 sg13g2_decap_8 FILLER_53_622 ();
 sg13g2_fill_2 FILLER_53_629 ();
 sg13g2_fill_1 FILLER_53_631 ();
 sg13g2_decap_8 FILLER_53_640 ();
 sg13g2_decap_8 FILLER_53_647 ();
 sg13g2_decap_8 FILLER_53_654 ();
 sg13g2_fill_2 FILLER_53_661 ();
 sg13g2_decap_4 FILLER_53_671 ();
 sg13g2_fill_1 FILLER_53_675 ();
 sg13g2_decap_8 FILLER_53_681 ();
 sg13g2_decap_8 FILLER_53_688 ();
 sg13g2_decap_8 FILLER_53_695 ();
 sg13g2_decap_4 FILLER_53_702 ();
 sg13g2_fill_1 FILLER_53_706 ();
 sg13g2_decap_8 FILLER_53_733 ();
 sg13g2_decap_8 FILLER_53_740 ();
 sg13g2_decap_8 FILLER_53_747 ();
 sg13g2_decap_8 FILLER_53_754 ();
 sg13g2_decap_8 FILLER_53_761 ();
 sg13g2_decap_8 FILLER_53_768 ();
 sg13g2_decap_8 FILLER_53_775 ();
 sg13g2_decap_8 FILLER_53_782 ();
 sg13g2_decap_8 FILLER_53_789 ();
 sg13g2_decap_8 FILLER_53_796 ();
 sg13g2_decap_8 FILLER_53_803 ();
 sg13g2_decap_4 FILLER_53_810 ();
 sg13g2_fill_2 FILLER_53_814 ();
 sg13g2_fill_2 FILLER_53_821 ();
 sg13g2_fill_1 FILLER_53_823 ();
 sg13g2_decap_8 FILLER_53_829 ();
 sg13g2_decap_8 FILLER_53_836 ();
 sg13g2_decap_8 FILLER_53_848 ();
 sg13g2_decap_8 FILLER_53_881 ();
 sg13g2_decap_8 FILLER_53_888 ();
 sg13g2_decap_4 FILLER_53_927 ();
 sg13g2_decap_8 FILLER_53_954 ();
 sg13g2_decap_8 FILLER_53_961 ();
 sg13g2_decap_8 FILLER_53_968 ();
 sg13g2_decap_8 FILLER_53_975 ();
 sg13g2_fill_1 FILLER_53_982 ();
 sg13g2_decap_8 FILLER_53_988 ();
 sg13g2_decap_8 FILLER_53_995 ();
 sg13g2_fill_2 FILLER_53_1002 ();
 sg13g2_fill_1 FILLER_53_1004 ();
 sg13g2_decap_8 FILLER_53_1021 ();
 sg13g2_decap_8 FILLER_53_1028 ();
 sg13g2_fill_2 FILLER_53_1035 ();
 sg13g2_fill_2 FILLER_53_1063 ();
 sg13g2_fill_1 FILLER_53_1065 ();
 sg13g2_decap_8 FILLER_53_1078 ();
 sg13g2_decap_8 FILLER_53_1085 ();
 sg13g2_decap_8 FILLER_53_1092 ();
 sg13g2_decap_8 FILLER_53_1099 ();
 sg13g2_decap_8 FILLER_53_1106 ();
 sg13g2_decap_8 FILLER_53_1113 ();
 sg13g2_decap_8 FILLER_53_1120 ();
 sg13g2_decap_8 FILLER_53_1127 ();
 sg13g2_decap_8 FILLER_53_1134 ();
 sg13g2_decap_8 FILLER_53_1141 ();
 sg13g2_decap_8 FILLER_53_1148 ();
 sg13g2_fill_1 FILLER_53_1155 ();
 sg13g2_decap_8 FILLER_53_1160 ();
 sg13g2_decap_8 FILLER_53_1167 ();
 sg13g2_decap_8 FILLER_53_1174 ();
 sg13g2_decap_8 FILLER_53_1181 ();
 sg13g2_decap_8 FILLER_53_1188 ();
 sg13g2_decap_8 FILLER_53_1195 ();
 sg13g2_decap_8 FILLER_53_1202 ();
 sg13g2_decap_8 FILLER_53_1209 ();
 sg13g2_fill_1 FILLER_53_1216 ();
 sg13g2_decap_8 FILLER_53_1238 ();
 sg13g2_decap_8 FILLER_53_1245 ();
 sg13g2_decap_8 FILLER_53_1252 ();
 sg13g2_decap_8 FILLER_53_1259 ();
 sg13g2_decap_8 FILLER_53_1266 ();
 sg13g2_decap_8 FILLER_53_1273 ();
 sg13g2_decap_8 FILLER_53_1280 ();
 sg13g2_decap_8 FILLER_53_1287 ();
 sg13g2_decap_8 FILLER_53_1294 ();
 sg13g2_decap_8 FILLER_53_1306 ();
 sg13g2_decap_8 FILLER_53_1313 ();
 sg13g2_decap_8 FILLER_53_1320 ();
 sg13g2_decap_8 FILLER_53_1327 ();
 sg13g2_decap_8 FILLER_53_1334 ();
 sg13g2_decap_8 FILLER_53_1341 ();
 sg13g2_decap_8 FILLER_53_1348 ();
 sg13g2_decap_8 FILLER_53_1355 ();
 sg13g2_decap_8 FILLER_53_1362 ();
 sg13g2_decap_8 FILLER_53_1369 ();
 sg13g2_decap_8 FILLER_53_1376 ();
 sg13g2_decap_8 FILLER_53_1383 ();
 sg13g2_decap_8 FILLER_53_1390 ();
 sg13g2_decap_8 FILLER_53_1397 ();
 sg13g2_decap_4 FILLER_53_1404 ();
 sg13g2_decap_8 FILLER_53_1418 ();
 sg13g2_decap_8 FILLER_53_1425 ();
 sg13g2_decap_8 FILLER_53_1432 ();
 sg13g2_decap_8 FILLER_53_1439 ();
 sg13g2_fill_2 FILLER_53_1446 ();
 sg13g2_fill_1 FILLER_53_1448 ();
 sg13g2_decap_8 FILLER_53_1487 ();
 sg13g2_decap_8 FILLER_53_1494 ();
 sg13g2_decap_4 FILLER_53_1501 ();
 sg13g2_fill_1 FILLER_53_1505 ();
 sg13g2_fill_2 FILLER_53_1520 ();
 sg13g2_decap_8 FILLER_53_1537 ();
 sg13g2_decap_8 FILLER_53_1544 ();
 sg13g2_decap_8 FILLER_53_1551 ();
 sg13g2_decap_8 FILLER_53_1558 ();
 sg13g2_decap_8 FILLER_53_1565 ();
 sg13g2_decap_8 FILLER_53_1572 ();
 sg13g2_decap_8 FILLER_53_1579 ();
 sg13g2_fill_2 FILLER_53_1586 ();
 sg13g2_decap_8 FILLER_53_1599 ();
 sg13g2_decap_8 FILLER_53_1606 ();
 sg13g2_decap_4 FILLER_53_1613 ();
 sg13g2_decap_8 FILLER_53_1622 ();
 sg13g2_decap_8 FILLER_53_1629 ();
 sg13g2_decap_4 FILLER_53_1636 ();
 sg13g2_decap_8 FILLER_53_1687 ();
 sg13g2_decap_8 FILLER_53_1694 ();
 sg13g2_decap_4 FILLER_53_1701 ();
 sg13g2_fill_1 FILLER_53_1705 ();
 sg13g2_decap_8 FILLER_53_1711 ();
 sg13g2_decap_4 FILLER_53_1718 ();
 sg13g2_decap_8 FILLER_53_1752 ();
 sg13g2_decap_4 FILLER_53_1759 ();
 sg13g2_fill_2 FILLER_53_1763 ();
 sg13g2_fill_2 FILLER_53_1797 ();
 sg13g2_fill_2 FILLER_53_1805 ();
 sg13g2_decap_8 FILLER_53_1813 ();
 sg13g2_decap_8 FILLER_53_1820 ();
 sg13g2_decap_8 FILLER_53_1827 ();
 sg13g2_decap_8 FILLER_53_1834 ();
 sg13g2_decap_8 FILLER_53_1841 ();
 sg13g2_decap_8 FILLER_53_1848 ();
 sg13g2_decap_8 FILLER_53_1855 ();
 sg13g2_fill_1 FILLER_53_1862 ();
 sg13g2_decap_8 FILLER_53_1873 ();
 sg13g2_decap_8 FILLER_53_1880 ();
 sg13g2_decap_8 FILLER_53_1887 ();
 sg13g2_decap_8 FILLER_53_1894 ();
 sg13g2_decap_8 FILLER_53_1901 ();
 sg13g2_decap_8 FILLER_53_1908 ();
 sg13g2_decap_4 FILLER_53_1915 ();
 sg13g2_fill_1 FILLER_53_1919 ();
 sg13g2_decap_8 FILLER_53_1930 ();
 sg13g2_decap_8 FILLER_53_1937 ();
 sg13g2_decap_8 FILLER_53_1944 ();
 sg13g2_decap_8 FILLER_53_1951 ();
 sg13g2_decap_4 FILLER_53_1964 ();
 sg13g2_fill_2 FILLER_53_1968 ();
 sg13g2_decap_8 FILLER_53_1996 ();
 sg13g2_decap_8 FILLER_53_2003 ();
 sg13g2_decap_4 FILLER_53_2010 ();
 sg13g2_decap_8 FILLER_53_2024 ();
 sg13g2_decap_8 FILLER_53_2031 ();
 sg13g2_decap_8 FILLER_53_2038 ();
 sg13g2_decap_8 FILLER_53_2045 ();
 sg13g2_decap_8 FILLER_53_2052 ();
 sg13g2_decap_4 FILLER_53_2059 ();
 sg13g2_fill_2 FILLER_53_2063 ();
 sg13g2_decap_8 FILLER_53_2075 ();
 sg13g2_decap_8 FILLER_53_2082 ();
 sg13g2_decap_8 FILLER_53_2089 ();
 sg13g2_decap_4 FILLER_53_2096 ();
 sg13g2_fill_1 FILLER_53_2100 ();
 sg13g2_fill_1 FILLER_53_2127 ();
 sg13g2_decap_8 FILLER_53_2167 ();
 sg13g2_decap_8 FILLER_53_2174 ();
 sg13g2_decap_8 FILLER_53_2181 ();
 sg13g2_decap_8 FILLER_53_2188 ();
 sg13g2_fill_2 FILLER_53_2195 ();
 sg13g2_fill_1 FILLER_53_2197 ();
 sg13g2_decap_8 FILLER_53_2211 ();
 sg13g2_decap_8 FILLER_53_2218 ();
 sg13g2_decap_4 FILLER_53_2225 ();
 sg13g2_decap_8 FILLER_53_2264 ();
 sg13g2_decap_8 FILLER_53_2271 ();
 sg13g2_decap_8 FILLER_53_2278 ();
 sg13g2_decap_4 FILLER_53_2285 ();
 sg13g2_fill_1 FILLER_53_2289 ();
 sg13g2_decap_8 FILLER_53_2296 ();
 sg13g2_decap_8 FILLER_53_2329 ();
 sg13g2_decap_8 FILLER_53_2336 ();
 sg13g2_decap_8 FILLER_53_2343 ();
 sg13g2_decap_4 FILLER_53_2350 ();
 sg13g2_fill_1 FILLER_53_2354 ();
 sg13g2_decap_8 FILLER_53_2401 ();
 sg13g2_decap_8 FILLER_53_2408 ();
 sg13g2_decap_8 FILLER_53_2421 ();
 sg13g2_decap_8 FILLER_53_2444 ();
 sg13g2_decap_8 FILLER_53_2451 ();
 sg13g2_decap_8 FILLER_53_2458 ();
 sg13g2_fill_2 FILLER_53_2465 ();
 sg13g2_fill_1 FILLER_53_2467 ();
 sg13g2_decap_8 FILLER_53_2474 ();
 sg13g2_decap_8 FILLER_53_2481 ();
 sg13g2_decap_4 FILLER_53_2488 ();
 sg13g2_fill_1 FILLER_53_2492 ();
 sg13g2_fill_1 FILLER_53_2519 ();
 sg13g2_decap_4 FILLER_53_2524 ();
 sg13g2_decap_8 FILLER_53_2532 ();
 sg13g2_decap_8 FILLER_53_2539 ();
 sg13g2_decap_8 FILLER_53_2546 ();
 sg13g2_decap_8 FILLER_53_2553 ();
 sg13g2_decap_8 FILLER_53_2560 ();
 sg13g2_decap_4 FILLER_53_2567 ();
 sg13g2_decap_8 FILLER_53_2597 ();
 sg13g2_decap_8 FILLER_53_2604 ();
 sg13g2_decap_8 FILLER_53_2611 ();
 sg13g2_decap_4 FILLER_53_2618 ();
 sg13g2_fill_2 FILLER_53_2622 ();
 sg13g2_decap_8 FILLER_53_2650 ();
 sg13g2_decap_8 FILLER_53_2657 ();
 sg13g2_decap_8 FILLER_53_2664 ();
 sg13g2_decap_8 FILLER_53_2671 ();
 sg13g2_decap_8 FILLER_53_2678 ();
 sg13g2_decap_8 FILLER_53_2685 ();
 sg13g2_fill_2 FILLER_53_2692 ();
 sg13g2_fill_1 FILLER_53_2694 ();
 sg13g2_decap_4 FILLER_53_2705 ();
 sg13g2_fill_2 FILLER_53_2709 ();
 sg13g2_decap_8 FILLER_53_2737 ();
 sg13g2_decap_8 FILLER_53_2744 ();
 sg13g2_decap_4 FILLER_53_2751 ();
 sg13g2_fill_2 FILLER_53_2755 ();
 sg13g2_decap_8 FILLER_53_2765 ();
 sg13g2_decap_4 FILLER_53_2772 ();
 sg13g2_decap_8 FILLER_53_2795 ();
 sg13g2_decap_8 FILLER_53_2802 ();
 sg13g2_decap_8 FILLER_53_2809 ();
 sg13g2_decap_4 FILLER_53_2816 ();
 sg13g2_fill_2 FILLER_53_2820 ();
 sg13g2_decap_8 FILLER_53_2846 ();
 sg13g2_decap_8 FILLER_53_2853 ();
 sg13g2_decap_8 FILLER_53_2860 ();
 sg13g2_decap_8 FILLER_53_2867 ();
 sg13g2_decap_8 FILLER_53_2874 ();
 sg13g2_decap_8 FILLER_53_2881 ();
 sg13g2_decap_8 FILLER_53_2888 ();
 sg13g2_decap_8 FILLER_53_2895 ();
 sg13g2_decap_8 FILLER_53_2902 ();
 sg13g2_decap_8 FILLER_53_2909 ();
 sg13g2_decap_8 FILLER_53_2916 ();
 sg13g2_decap_8 FILLER_53_2931 ();
 sg13g2_fill_2 FILLER_53_2938 ();
 sg13g2_decap_8 FILLER_53_2946 ();
 sg13g2_decap_8 FILLER_53_2953 ();
 sg13g2_decap_4 FILLER_53_2960 ();
 sg13g2_fill_2 FILLER_53_2964 ();
 sg13g2_decap_8 FILLER_53_2986 ();
 sg13g2_decap_8 FILLER_53_2993 ();
 sg13g2_decap_8 FILLER_53_3000 ();
 sg13g2_decap_8 FILLER_53_3007 ();
 sg13g2_decap_8 FILLER_53_3014 ();
 sg13g2_decap_8 FILLER_53_3021 ();
 sg13g2_fill_2 FILLER_53_3028 ();
 sg13g2_fill_1 FILLER_53_3030 ();
 sg13g2_decap_8 FILLER_53_3057 ();
 sg13g2_decap_8 FILLER_53_3064 ();
 sg13g2_decap_8 FILLER_53_3071 ();
 sg13g2_decap_8 FILLER_53_3078 ();
 sg13g2_decap_4 FILLER_53_3085 ();
 sg13g2_fill_1 FILLER_53_3089 ();
 sg13g2_decap_8 FILLER_53_3109 ();
 sg13g2_decap_8 FILLER_53_3116 ();
 sg13g2_decap_8 FILLER_53_3123 ();
 sg13g2_decap_8 FILLER_53_3130 ();
 sg13g2_decap_8 FILLER_53_3137 ();
 sg13g2_decap_4 FILLER_53_3154 ();
 sg13g2_decap_8 FILLER_53_3179 ();
 sg13g2_decap_8 FILLER_53_3186 ();
 sg13g2_decap_8 FILLER_53_3193 ();
 sg13g2_fill_2 FILLER_53_3200 ();
 sg13g2_fill_2 FILLER_53_3210 ();
 sg13g2_decap_8 FILLER_53_3225 ();
 sg13g2_fill_2 FILLER_53_3232 ();
 sg13g2_decap_8 FILLER_53_3248 ();
 sg13g2_decap_8 FILLER_53_3255 ();
 sg13g2_decap_8 FILLER_53_3262 ();
 sg13g2_decap_8 FILLER_53_3269 ();
 sg13g2_fill_2 FILLER_53_3276 ();
 sg13g2_fill_1 FILLER_53_3278 ();
 sg13g2_fill_1 FILLER_53_3315 ();
 sg13g2_decap_4 FILLER_53_3326 ();
 sg13g2_decap_8 FILLER_53_3382 ();
 sg13g2_decap_8 FILLER_53_3389 ();
 sg13g2_decap_8 FILLER_53_3396 ();
 sg13g2_decap_4 FILLER_53_3403 ();
 sg13g2_fill_1 FILLER_53_3407 ();
 sg13g2_decap_8 FILLER_53_3428 ();
 sg13g2_decap_8 FILLER_53_3435 ();
 sg13g2_decap_8 FILLER_53_3485 ();
 sg13g2_decap_8 FILLER_53_3492 ();
 sg13g2_decap_8 FILLER_53_3499 ();
 sg13g2_decap_8 FILLER_53_3506 ();
 sg13g2_decap_8 FILLER_53_3513 ();
 sg13g2_decap_8 FILLER_53_3520 ();
 sg13g2_decap_8 FILLER_53_3532 ();
 sg13g2_decap_8 FILLER_53_3539 ();
 sg13g2_decap_8 FILLER_53_3546 ();
 sg13g2_decap_8 FILLER_53_3553 ();
 sg13g2_decap_8 FILLER_53_3560 ();
 sg13g2_decap_8 FILLER_53_3567 ();
 sg13g2_decap_4 FILLER_53_3574 ();
 sg13g2_fill_2 FILLER_53_3578 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_fill_2 FILLER_54_7 ();
 sg13g2_fill_1 FILLER_54_40 ();
 sg13g2_fill_1 FILLER_54_54 ();
 sg13g2_decap_8 FILLER_54_95 ();
 sg13g2_fill_2 FILLER_54_102 ();
 sg13g2_fill_2 FILLER_54_110 ();
 sg13g2_decap_8 FILLER_54_118 ();
 sg13g2_decap_8 FILLER_54_125 ();
 sg13g2_decap_8 FILLER_54_132 ();
 sg13g2_decap_8 FILLER_54_139 ();
 sg13g2_decap_8 FILLER_54_146 ();
 sg13g2_fill_2 FILLER_54_153 ();
 sg13g2_fill_2 FILLER_54_161 ();
 sg13g2_fill_1 FILLER_54_163 ();
 sg13g2_decap_8 FILLER_54_176 ();
 sg13g2_decap_8 FILLER_54_183 ();
 sg13g2_decap_8 FILLER_54_190 ();
 sg13g2_decap_8 FILLER_54_197 ();
 sg13g2_decap_8 FILLER_54_204 ();
 sg13g2_decap_8 FILLER_54_211 ();
 sg13g2_decap_8 FILLER_54_218 ();
 sg13g2_decap_8 FILLER_54_230 ();
 sg13g2_decap_8 FILLER_54_237 ();
 sg13g2_decap_8 FILLER_54_244 ();
 sg13g2_fill_1 FILLER_54_251 ();
 sg13g2_decap_8 FILLER_54_260 ();
 sg13g2_decap_8 FILLER_54_267 ();
 sg13g2_decap_8 FILLER_54_274 ();
 sg13g2_fill_2 FILLER_54_281 ();
 sg13g2_fill_1 FILLER_54_283 ();
 sg13g2_decap_8 FILLER_54_289 ();
 sg13g2_decap_4 FILLER_54_296 ();
 sg13g2_decap_8 FILLER_54_313 ();
 sg13g2_decap_8 FILLER_54_320 ();
 sg13g2_decap_8 FILLER_54_327 ();
 sg13g2_fill_2 FILLER_54_334 ();
 sg13g2_decap_4 FILLER_54_362 ();
 sg13g2_fill_1 FILLER_54_366 ();
 sg13g2_decap_4 FILLER_54_386 ();
 sg13g2_fill_1 FILLER_54_390 ();
 sg13g2_decap_8 FILLER_54_417 ();
 sg13g2_decap_8 FILLER_54_424 ();
 sg13g2_decap_8 FILLER_54_431 ();
 sg13g2_fill_2 FILLER_54_438 ();
 sg13g2_decap_8 FILLER_54_448 ();
 sg13g2_decap_4 FILLER_54_455 ();
 sg13g2_fill_2 FILLER_54_459 ();
 sg13g2_decap_4 FILLER_54_469 ();
 sg13g2_decap_4 FILLER_54_481 ();
 sg13g2_decap_8 FILLER_54_498 ();
 sg13g2_decap_8 FILLER_54_505 ();
 sg13g2_decap_4 FILLER_54_512 ();
 sg13g2_fill_2 FILLER_54_516 ();
 sg13g2_decap_4 FILLER_54_524 ();
 sg13g2_fill_1 FILLER_54_528 ();
 sg13g2_fill_1 FILLER_54_539 ();
 sg13g2_decap_8 FILLER_54_566 ();
 sg13g2_decap_8 FILLER_54_573 ();
 sg13g2_decap_8 FILLER_54_580 ();
 sg13g2_decap_8 FILLER_54_587 ();
 sg13g2_decap_8 FILLER_54_594 ();
 sg13g2_fill_2 FILLER_54_601 ();
 sg13g2_fill_1 FILLER_54_603 ();
 sg13g2_decap_8 FILLER_54_609 ();
 sg13g2_decap_8 FILLER_54_616 ();
 sg13g2_decap_8 FILLER_54_623 ();
 sg13g2_fill_1 FILLER_54_630 ();
 sg13g2_decap_8 FILLER_54_639 ();
 sg13g2_decap_8 FILLER_54_646 ();
 sg13g2_decap_4 FILLER_54_653 ();
 sg13g2_fill_2 FILLER_54_657 ();
 sg13g2_fill_2 FILLER_54_679 ();
 sg13g2_decap_8 FILLER_54_689 ();
 sg13g2_decap_8 FILLER_54_696 ();
 sg13g2_decap_8 FILLER_54_703 ();
 sg13g2_decap_8 FILLER_54_736 ();
 sg13g2_fill_2 FILLER_54_743 ();
 sg13g2_decap_8 FILLER_54_755 ();
 sg13g2_decap_4 FILLER_54_762 ();
 sg13g2_fill_1 FILLER_54_766 ();
 sg13g2_decap_8 FILLER_54_778 ();
 sg13g2_decap_8 FILLER_54_785 ();
 sg13g2_decap_8 FILLER_54_792 ();
 sg13g2_decap_8 FILLER_54_799 ();
 sg13g2_decap_8 FILLER_54_806 ();
 sg13g2_decap_8 FILLER_54_813 ();
 sg13g2_decap_4 FILLER_54_820 ();
 sg13g2_decap_8 FILLER_54_829 ();
 sg13g2_decap_8 FILLER_54_836 ();
 sg13g2_decap_4 FILLER_54_843 ();
 sg13g2_fill_1 FILLER_54_847 ();
 sg13g2_decap_8 FILLER_54_853 ();
 sg13g2_decap_8 FILLER_54_860 ();
 sg13g2_decap_8 FILLER_54_876 ();
 sg13g2_decap_4 FILLER_54_883 ();
 sg13g2_decap_8 FILLER_54_893 ();
 sg13g2_decap_8 FILLER_54_900 ();
 sg13g2_decap_8 FILLER_54_907 ();
 sg13g2_decap_4 FILLER_54_914 ();
 sg13g2_fill_1 FILLER_54_918 ();
 sg13g2_decap_8 FILLER_54_931 ();
 sg13g2_decap_8 FILLER_54_938 ();
 sg13g2_decap_8 FILLER_54_945 ();
 sg13g2_decap_8 FILLER_54_952 ();
 sg13g2_decap_8 FILLER_54_959 ();
 sg13g2_decap_8 FILLER_54_966 ();
 sg13g2_decap_8 FILLER_54_973 ();
 sg13g2_decap_8 FILLER_54_980 ();
 sg13g2_decap_8 FILLER_54_987 ();
 sg13g2_decap_8 FILLER_54_994 ();
 sg13g2_decap_8 FILLER_54_1001 ();
 sg13g2_fill_2 FILLER_54_1008 ();
 sg13g2_fill_1 FILLER_54_1010 ();
 sg13g2_decap_8 FILLER_54_1019 ();
 sg13g2_decap_8 FILLER_54_1026 ();
 sg13g2_decap_8 FILLER_54_1033 ();
 sg13g2_decap_8 FILLER_54_1040 ();
 sg13g2_decap_8 FILLER_54_1047 ();
 sg13g2_fill_2 FILLER_54_1080 ();
 sg13g2_fill_1 FILLER_54_1082 ();
 sg13g2_decap_8 FILLER_54_1093 ();
 sg13g2_decap_8 FILLER_54_1100 ();
 sg13g2_fill_1 FILLER_54_1107 ();
 sg13g2_decap_8 FILLER_54_1116 ();
 sg13g2_decap_8 FILLER_54_1123 ();
 sg13g2_decap_8 FILLER_54_1130 ();
 sg13g2_decap_8 FILLER_54_1147 ();
 sg13g2_decap_8 FILLER_54_1154 ();
 sg13g2_decap_8 FILLER_54_1161 ();
 sg13g2_decap_8 FILLER_54_1168 ();
 sg13g2_decap_8 FILLER_54_1175 ();
 sg13g2_decap_8 FILLER_54_1182 ();
 sg13g2_fill_2 FILLER_54_1189 ();
 sg13g2_fill_1 FILLER_54_1201 ();
 sg13g2_fill_2 FILLER_54_1207 ();
 sg13g2_fill_1 FILLER_54_1209 ();
 sg13g2_decap_8 FILLER_54_1214 ();
 sg13g2_decap_8 FILLER_54_1221 ();
 sg13g2_fill_1 FILLER_54_1228 ();
 sg13g2_decap_8 FILLER_54_1271 ();
 sg13g2_decap_8 FILLER_54_1278 ();
 sg13g2_decap_4 FILLER_54_1285 ();
 sg13g2_decap_4 FILLER_54_1297 ();
 sg13g2_decap_8 FILLER_54_1311 ();
 sg13g2_fill_2 FILLER_54_1318 ();
 sg13g2_decap_8 FILLER_54_1335 ();
 sg13g2_decap_8 FILLER_54_1342 ();
 sg13g2_decap_4 FILLER_54_1385 ();
 sg13g2_fill_1 FILLER_54_1389 ();
 sg13g2_decap_8 FILLER_54_1400 ();
 sg13g2_decap_8 FILLER_54_1433 ();
 sg13g2_decap_8 FILLER_54_1440 ();
 sg13g2_decap_4 FILLER_54_1447 ();
 sg13g2_fill_2 FILLER_54_1451 ();
 sg13g2_decap_8 FILLER_54_1459 ();
 sg13g2_decap_8 FILLER_54_1495 ();
 sg13g2_decap_8 FILLER_54_1502 ();
 sg13g2_fill_1 FILLER_54_1509 ();
 sg13g2_decap_8 FILLER_54_1515 ();
 sg13g2_decap_8 FILLER_54_1522 ();
 sg13g2_decap_8 FILLER_54_1529 ();
 sg13g2_decap_8 FILLER_54_1536 ();
 sg13g2_fill_1 FILLER_54_1543 ();
 sg13g2_decap_4 FILLER_54_1549 ();
 sg13g2_decap_8 FILLER_54_1563 ();
 sg13g2_decap_8 FILLER_54_1570 ();
 sg13g2_decap_8 FILLER_54_1577 ();
 sg13g2_decap_8 FILLER_54_1584 ();
 sg13g2_decap_8 FILLER_54_1591 ();
 sg13g2_fill_1 FILLER_54_1598 ();
 sg13g2_decap_8 FILLER_54_1618 ();
 sg13g2_decap_8 FILLER_54_1625 ();
 sg13g2_decap_8 FILLER_54_1632 ();
 sg13g2_decap_8 FILLER_54_1639 ();
 sg13g2_decap_8 FILLER_54_1646 ();
 sg13g2_fill_1 FILLER_54_1653 ();
 sg13g2_decap_8 FILLER_54_1664 ();
 sg13g2_decap_8 FILLER_54_1671 ();
 sg13g2_decap_8 FILLER_54_1678 ();
 sg13g2_decap_8 FILLER_54_1685 ();
 sg13g2_decap_8 FILLER_54_1692 ();
 sg13g2_decap_8 FILLER_54_1699 ();
 sg13g2_decap_8 FILLER_54_1706 ();
 sg13g2_decap_8 FILLER_54_1713 ();
 sg13g2_fill_1 FILLER_54_1720 ();
 sg13g2_fill_1 FILLER_54_1725 ();
 sg13g2_decap_8 FILLER_54_1752 ();
 sg13g2_fill_1 FILLER_54_1759 ();
 sg13g2_fill_2 FILLER_54_1773 ();
 sg13g2_fill_2 FILLER_54_1785 ();
 sg13g2_fill_2 FILLER_54_1808 ();
 sg13g2_decap_8 FILLER_54_1846 ();
 sg13g2_decap_8 FILLER_54_1853 ();
 sg13g2_decap_4 FILLER_54_1860 ();
 sg13g2_fill_1 FILLER_54_1864 ();
 sg13g2_decap_8 FILLER_54_1897 ();
 sg13g2_decap_8 FILLER_54_1904 ();
 sg13g2_fill_2 FILLER_54_1911 ();
 sg13g2_fill_1 FILLER_54_1913 ();
 sg13g2_decap_8 FILLER_54_1940 ();
 sg13g2_decap_8 FILLER_54_1947 ();
 sg13g2_decap_8 FILLER_54_1954 ();
 sg13g2_decap_8 FILLER_54_1961 ();
 sg13g2_decap_8 FILLER_54_1968 ();
 sg13g2_decap_8 FILLER_54_1975 ();
 sg13g2_decap_8 FILLER_54_1982 ();
 sg13g2_fill_2 FILLER_54_1989 ();
 sg13g2_fill_1 FILLER_54_1991 ();
 sg13g2_decap_8 FILLER_54_1998 ();
 sg13g2_decap_8 FILLER_54_2005 ();
 sg13g2_decap_8 FILLER_54_2038 ();
 sg13g2_decap_8 FILLER_54_2045 ();
 sg13g2_decap_8 FILLER_54_2052 ();
 sg13g2_decap_8 FILLER_54_2085 ();
 sg13g2_fill_2 FILLER_54_2092 ();
 sg13g2_fill_1 FILLER_54_2094 ();
 sg13g2_decap_8 FILLER_54_2111 ();
 sg13g2_decap_8 FILLER_54_2118 ();
 sg13g2_fill_2 FILLER_54_2125 ();
 sg13g2_fill_1 FILLER_54_2127 ();
 sg13g2_decap_8 FILLER_54_2136 ();
 sg13g2_decap_8 FILLER_54_2143 ();
 sg13g2_decap_8 FILLER_54_2150 ();
 sg13g2_decap_8 FILLER_54_2157 ();
 sg13g2_decap_8 FILLER_54_2190 ();
 sg13g2_decap_8 FILLER_54_2197 ();
 sg13g2_decap_8 FILLER_54_2204 ();
 sg13g2_decap_8 FILLER_54_2211 ();
 sg13g2_decap_8 FILLER_54_2218 ();
 sg13g2_decap_4 FILLER_54_2225 ();
 sg13g2_fill_2 FILLER_54_2229 ();
 sg13g2_decap_8 FILLER_54_2243 ();
 sg13g2_decap_8 FILLER_54_2250 ();
 sg13g2_decap_4 FILLER_54_2257 ();
 sg13g2_fill_2 FILLER_54_2261 ();
 sg13g2_decap_8 FILLER_54_2280 ();
 sg13g2_decap_8 FILLER_54_2287 ();
 sg13g2_decap_8 FILLER_54_2294 ();
 sg13g2_fill_1 FILLER_54_2301 ();
 sg13g2_decap_8 FILLER_54_2312 ();
 sg13g2_decap_8 FILLER_54_2319 ();
 sg13g2_decap_8 FILLER_54_2326 ();
 sg13g2_decap_8 FILLER_54_2333 ();
 sg13g2_fill_1 FILLER_54_2340 ();
 sg13g2_decap_8 FILLER_54_2346 ();
 sg13g2_decap_8 FILLER_54_2353 ();
 sg13g2_fill_1 FILLER_54_2360 ();
 sg13g2_fill_1 FILLER_54_2371 ();
 sg13g2_decap_8 FILLER_54_2375 ();
 sg13g2_decap_8 FILLER_54_2382 ();
 sg13g2_decap_8 FILLER_54_2389 ();
 sg13g2_decap_8 FILLER_54_2396 ();
 sg13g2_fill_2 FILLER_54_2403 ();
 sg13g2_fill_1 FILLER_54_2405 ();
 sg13g2_decap_8 FILLER_54_2412 ();
 sg13g2_decap_8 FILLER_54_2419 ();
 sg13g2_decap_8 FILLER_54_2426 ();
 sg13g2_decap_8 FILLER_54_2433 ();
 sg13g2_decap_8 FILLER_54_2440 ();
 sg13g2_decap_8 FILLER_54_2447 ();
 sg13g2_fill_2 FILLER_54_2454 ();
 sg13g2_decap_8 FILLER_54_2470 ();
 sg13g2_decap_8 FILLER_54_2477 ();
 sg13g2_decap_8 FILLER_54_2484 ();
 sg13g2_decap_8 FILLER_54_2491 ();
 sg13g2_decap_8 FILLER_54_2498 ();
 sg13g2_decap_4 FILLER_54_2505 ();
 sg13g2_fill_1 FILLER_54_2509 ();
 sg13g2_decap_8 FILLER_54_2520 ();
 sg13g2_decap_8 FILLER_54_2527 ();
 sg13g2_decap_8 FILLER_54_2534 ();
 sg13g2_fill_2 FILLER_54_2541 ();
 sg13g2_decap_4 FILLER_54_2548 ();
 sg13g2_fill_1 FILLER_54_2552 ();
 sg13g2_decap_8 FILLER_54_2589 ();
 sg13g2_decap_8 FILLER_54_2596 ();
 sg13g2_decap_8 FILLER_54_2603 ();
 sg13g2_fill_2 FILLER_54_2610 ();
 sg13g2_fill_1 FILLER_54_2612 ();
 sg13g2_decap_8 FILLER_54_2649 ();
 sg13g2_decap_8 FILLER_54_2656 ();
 sg13g2_decap_8 FILLER_54_2663 ();
 sg13g2_fill_2 FILLER_54_2670 ();
 sg13g2_fill_1 FILLER_54_2672 ();
 sg13g2_decap_8 FILLER_54_2682 ();
 sg13g2_decap_8 FILLER_54_2689 ();
 sg13g2_decap_8 FILLER_54_2696 ();
 sg13g2_decap_8 FILLER_54_2723 ();
 sg13g2_decap_8 FILLER_54_2730 ();
 sg13g2_decap_8 FILLER_54_2737 ();
 sg13g2_decap_8 FILLER_54_2744 ();
 sg13g2_decap_8 FILLER_54_2751 ();
 sg13g2_decap_8 FILLER_54_2758 ();
 sg13g2_fill_1 FILLER_54_2765 ();
 sg13g2_decap_8 FILLER_54_2771 ();
 sg13g2_decap_8 FILLER_54_2778 ();
 sg13g2_decap_8 FILLER_54_2785 ();
 sg13g2_decap_8 FILLER_54_2792 ();
 sg13g2_decap_8 FILLER_54_2799 ();
 sg13g2_decap_8 FILLER_54_2806 ();
 sg13g2_decap_8 FILLER_54_2813 ();
 sg13g2_decap_8 FILLER_54_2820 ();
 sg13g2_decap_8 FILLER_54_2827 ();
 sg13g2_fill_1 FILLER_54_2834 ();
 sg13g2_decap_8 FILLER_54_2844 ();
 sg13g2_decap_8 FILLER_54_2851 ();
 sg13g2_decap_8 FILLER_54_2858 ();
 sg13g2_decap_4 FILLER_54_2865 ();
 sg13g2_fill_2 FILLER_54_2869 ();
 sg13g2_decap_8 FILLER_54_2876 ();
 sg13g2_fill_2 FILLER_54_2888 ();
 sg13g2_decap_8 FILLER_54_2898 ();
 sg13g2_decap_8 FILLER_54_2905 ();
 sg13g2_decap_8 FILLER_54_2912 ();
 sg13g2_decap_4 FILLER_54_2919 ();
 sg13g2_decap_8 FILLER_54_2949 ();
 sg13g2_decap_8 FILLER_54_2956 ();
 sg13g2_decap_8 FILLER_54_2963 ();
 sg13g2_decap_8 FILLER_54_2970 ();
 sg13g2_decap_8 FILLER_54_2977 ();
 sg13g2_decap_4 FILLER_54_2984 ();
 sg13g2_fill_2 FILLER_54_2988 ();
 sg13g2_decap_8 FILLER_54_3003 ();
 sg13g2_decap_4 FILLER_54_3010 ();
 sg13g2_fill_2 FILLER_54_3014 ();
 sg13g2_decap_8 FILLER_54_3052 ();
 sg13g2_decap_8 FILLER_54_3059 ();
 sg13g2_decap_8 FILLER_54_3066 ();
 sg13g2_decap_8 FILLER_54_3073 ();
 sg13g2_decap_8 FILLER_54_3080 ();
 sg13g2_fill_2 FILLER_54_3087 ();
 sg13g2_fill_1 FILLER_54_3089 ();
 sg13g2_decap_8 FILLER_54_3116 ();
 sg13g2_decap_8 FILLER_54_3123 ();
 sg13g2_decap_8 FILLER_54_3130 ();
 sg13g2_decap_8 FILLER_54_3137 ();
 sg13g2_decap_8 FILLER_54_3144 ();
 sg13g2_decap_4 FILLER_54_3156 ();
 sg13g2_fill_2 FILLER_54_3160 ();
 sg13g2_decap_8 FILLER_54_3182 ();
 sg13g2_decap_8 FILLER_54_3189 ();
 sg13g2_decap_8 FILLER_54_3196 ();
 sg13g2_fill_2 FILLER_54_3203 ();
 sg13g2_fill_2 FILLER_54_3215 ();
 sg13g2_fill_1 FILLER_54_3217 ();
 sg13g2_decap_8 FILLER_54_3244 ();
 sg13g2_decap_8 FILLER_54_3251 ();
 sg13g2_decap_8 FILLER_54_3258 ();
 sg13g2_decap_8 FILLER_54_3265 ();
 sg13g2_decap_8 FILLER_54_3272 ();
 sg13g2_decap_8 FILLER_54_3289 ();
 sg13g2_decap_8 FILLER_54_3296 ();
 sg13g2_decap_8 FILLER_54_3303 ();
 sg13g2_decap_8 FILLER_54_3310 ();
 sg13g2_decap_8 FILLER_54_3317 ();
 sg13g2_decap_4 FILLER_54_3324 ();
 sg13g2_fill_2 FILLER_54_3328 ();
 sg13g2_decap_8 FILLER_54_3340 ();
 sg13g2_decap_8 FILLER_54_3347 ();
 sg13g2_decap_8 FILLER_54_3354 ();
 sg13g2_fill_2 FILLER_54_3361 ();
 sg13g2_fill_1 FILLER_54_3363 ();
 sg13g2_decap_8 FILLER_54_3372 ();
 sg13g2_decap_8 FILLER_54_3379 ();
 sg13g2_decap_8 FILLER_54_3386 ();
 sg13g2_decap_8 FILLER_54_3393 ();
 sg13g2_decap_8 FILLER_54_3400 ();
 sg13g2_decap_8 FILLER_54_3407 ();
 sg13g2_decap_8 FILLER_54_3414 ();
 sg13g2_decap_4 FILLER_54_3421 ();
 sg13g2_decap_8 FILLER_54_3430 ();
 sg13g2_decap_8 FILLER_54_3437 ();
 sg13g2_decap_8 FILLER_54_3444 ();
 sg13g2_decap_8 FILLER_54_3451 ();
 sg13g2_decap_4 FILLER_54_3458 ();
 sg13g2_decap_8 FILLER_54_3484 ();
 sg13g2_decap_8 FILLER_54_3491 ();
 sg13g2_decap_8 FILLER_54_3498 ();
 sg13g2_decap_8 FILLER_54_3505 ();
 sg13g2_decap_8 FILLER_54_3512 ();
 sg13g2_decap_8 FILLER_54_3519 ();
 sg13g2_fill_1 FILLER_54_3526 ();
 sg13g2_decap_8 FILLER_54_3536 ();
 sg13g2_fill_1 FILLER_54_3543 ();
 sg13g2_decap_8 FILLER_54_3553 ();
 sg13g2_decap_8 FILLER_54_3560 ();
 sg13g2_decap_8 FILLER_54_3567 ();
 sg13g2_decap_4 FILLER_54_3574 ();
 sg13g2_fill_2 FILLER_54_3578 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_decap_8 FILLER_55_7 ();
 sg13g2_decap_8 FILLER_55_14 ();
 sg13g2_decap_8 FILLER_55_21 ();
 sg13g2_fill_1 FILLER_55_28 ();
 sg13g2_fill_2 FILLER_55_53 ();
 sg13g2_fill_1 FILLER_55_55 ();
 sg13g2_fill_2 FILLER_55_74 ();
 sg13g2_fill_1 FILLER_55_76 ();
 sg13g2_fill_2 FILLER_55_85 ();
 sg13g2_fill_1 FILLER_55_87 ();
 sg13g2_decap_4 FILLER_55_96 ();
 sg13g2_fill_1 FILLER_55_100 ();
 sg13g2_decap_8 FILLER_55_128 ();
 sg13g2_decap_8 FILLER_55_135 ();
 sg13g2_decap_8 FILLER_55_142 ();
 sg13g2_decap_8 FILLER_55_149 ();
 sg13g2_decap_4 FILLER_55_156 ();
 sg13g2_fill_1 FILLER_55_160 ();
 sg13g2_decap_8 FILLER_55_166 ();
 sg13g2_decap_8 FILLER_55_173 ();
 sg13g2_decap_8 FILLER_55_180 ();
 sg13g2_decap_8 FILLER_55_187 ();
 sg13g2_decap_8 FILLER_55_194 ();
 sg13g2_decap_8 FILLER_55_201 ();
 sg13g2_decap_8 FILLER_55_208 ();
 sg13g2_decap_8 FILLER_55_215 ();
 sg13g2_decap_8 FILLER_55_222 ();
 sg13g2_decap_8 FILLER_55_229 ();
 sg13g2_decap_8 FILLER_55_236 ();
 sg13g2_decap_8 FILLER_55_243 ();
 sg13g2_decap_8 FILLER_55_250 ();
 sg13g2_decap_8 FILLER_55_262 ();
 sg13g2_decap_8 FILLER_55_269 ();
 sg13g2_decap_8 FILLER_55_276 ();
 sg13g2_decap_8 FILLER_55_283 ();
 sg13g2_decap_8 FILLER_55_321 ();
 sg13g2_decap_4 FILLER_55_328 ();
 sg13g2_decap_8 FILLER_55_346 ();
 sg13g2_decap_8 FILLER_55_353 ();
 sg13g2_fill_1 FILLER_55_372 ();
 sg13g2_fill_1 FILLER_55_403 ();
 sg13g2_fill_2 FILLER_55_412 ();
 sg13g2_decap_8 FILLER_55_423 ();
 sg13g2_decap_4 FILLER_55_430 ();
 sg13g2_decap_8 FILLER_55_445 ();
 sg13g2_decap_8 FILLER_55_452 ();
 sg13g2_decap_8 FILLER_55_459 ();
 sg13g2_fill_1 FILLER_55_466 ();
 sg13g2_fill_1 FILLER_55_476 ();
 sg13g2_decap_8 FILLER_55_509 ();
 sg13g2_decap_8 FILLER_55_516 ();
 sg13g2_fill_1 FILLER_55_523 ();
 sg13g2_decap_8 FILLER_55_527 ();
 sg13g2_fill_1 FILLER_55_542 ();
 sg13g2_decap_8 FILLER_55_565 ();
 sg13g2_decap_8 FILLER_55_572 ();
 sg13g2_decap_8 FILLER_55_579 ();
 sg13g2_decap_8 FILLER_55_586 ();
 sg13g2_decap_4 FILLER_55_593 ();
 sg13g2_fill_1 FILLER_55_597 ();
 sg13g2_decap_8 FILLER_55_602 ();
 sg13g2_fill_2 FILLER_55_609 ();
 sg13g2_decap_4 FILLER_55_645 ();
 sg13g2_decap_8 FILLER_55_655 ();
 sg13g2_decap_4 FILLER_55_662 ();
 sg13g2_fill_2 FILLER_55_666 ();
 sg13g2_fill_2 FILLER_55_678 ();
 sg13g2_fill_1 FILLER_55_680 ();
 sg13g2_decap_4 FILLER_55_687 ();
 sg13g2_fill_2 FILLER_55_691 ();
 sg13g2_decap_4 FILLER_55_699 ();
 sg13g2_fill_1 FILLER_55_703 ();
 sg13g2_decap_8 FILLER_55_722 ();
 sg13g2_fill_1 FILLER_55_729 ();
 sg13g2_fill_1 FILLER_55_755 ();
 sg13g2_fill_1 FILLER_55_779 ();
 sg13g2_decap_8 FILLER_55_796 ();
 sg13g2_decap_8 FILLER_55_803 ();
 sg13g2_decap_8 FILLER_55_810 ();
 sg13g2_decap_4 FILLER_55_817 ();
 sg13g2_fill_2 FILLER_55_821 ();
 sg13g2_decap_8 FILLER_55_831 ();
 sg13g2_decap_8 FILLER_55_838 ();
 sg13g2_decap_8 FILLER_55_845 ();
 sg13g2_decap_8 FILLER_55_852 ();
 sg13g2_decap_8 FILLER_55_859 ();
 sg13g2_decap_8 FILLER_55_866 ();
 sg13g2_decap_8 FILLER_55_873 ();
 sg13g2_decap_8 FILLER_55_880 ();
 sg13g2_decap_8 FILLER_55_887 ();
 sg13g2_decap_8 FILLER_55_894 ();
 sg13g2_decap_8 FILLER_55_901 ();
 sg13g2_decap_8 FILLER_55_908 ();
 sg13g2_decap_8 FILLER_55_915 ();
 sg13g2_decap_8 FILLER_55_922 ();
 sg13g2_decap_4 FILLER_55_929 ();
 sg13g2_fill_1 FILLER_55_933 ();
 sg13g2_decap_8 FILLER_55_941 ();
 sg13g2_decap_8 FILLER_55_948 ();
 sg13g2_decap_8 FILLER_55_955 ();
 sg13g2_decap_8 FILLER_55_962 ();
 sg13g2_decap_8 FILLER_55_969 ();
 sg13g2_decap_8 FILLER_55_976 ();
 sg13g2_decap_8 FILLER_55_983 ();
 sg13g2_decap_8 FILLER_55_990 ();
 sg13g2_decap_8 FILLER_55_997 ();
 sg13g2_decap_8 FILLER_55_1004 ();
 sg13g2_decap_8 FILLER_55_1011 ();
 sg13g2_decap_8 FILLER_55_1018 ();
 sg13g2_decap_8 FILLER_55_1025 ();
 sg13g2_decap_8 FILLER_55_1032 ();
 sg13g2_decap_8 FILLER_55_1039 ();
 sg13g2_decap_8 FILLER_55_1046 ();
 sg13g2_decap_4 FILLER_55_1053 ();
 sg13g2_fill_1 FILLER_55_1057 ();
 sg13g2_fill_2 FILLER_55_1068 ();
 sg13g2_fill_1 FILLER_55_1070 ();
 sg13g2_decap_4 FILLER_55_1080 ();
 sg13g2_fill_1 FILLER_55_1084 ();
 sg13g2_fill_2 FILLER_55_1111 ();
 sg13g2_decap_8 FILLER_55_1123 ();
 sg13g2_fill_1 FILLER_55_1130 ();
 sg13g2_fill_2 FILLER_55_1173 ();
 sg13g2_fill_1 FILLER_55_1183 ();
 sg13g2_fill_2 FILLER_55_1213 ();
 sg13g2_fill_1 FILLER_55_1215 ();
 sg13g2_fill_2 FILLER_55_1221 ();
 sg13g2_fill_2 FILLER_55_1249 ();
 sg13g2_fill_2 FILLER_55_1261 ();
 sg13g2_decap_4 FILLER_55_1273 ();
 sg13g2_fill_1 FILLER_55_1282 ();
 sg13g2_decap_4 FILLER_55_1287 ();
 sg13g2_fill_1 FILLER_55_1291 ();
 sg13g2_decap_8 FILLER_55_1301 ();
 sg13g2_decap_4 FILLER_55_1308 ();
 sg13g2_decap_8 FILLER_55_1347 ();
 sg13g2_decap_4 FILLER_55_1354 ();
 sg13g2_fill_2 FILLER_55_1358 ();
 sg13g2_decap_4 FILLER_55_1372 ();
 sg13g2_fill_2 FILLER_55_1376 ();
 sg13g2_decap_8 FILLER_55_1383 ();
 sg13g2_fill_2 FILLER_55_1390 ();
 sg13g2_fill_1 FILLER_55_1392 ();
 sg13g2_decap_8 FILLER_55_1419 ();
 sg13g2_decap_8 FILLER_55_1426 ();
 sg13g2_decap_8 FILLER_55_1433 ();
 sg13g2_decap_8 FILLER_55_1440 ();
 sg13g2_decap_8 FILLER_55_1447 ();
 sg13g2_decap_8 FILLER_55_1454 ();
 sg13g2_fill_1 FILLER_55_1461 ();
 sg13g2_decap_4 FILLER_55_1466 ();
 sg13g2_fill_1 FILLER_55_1476 ();
 sg13g2_decap_8 FILLER_55_1488 ();
 sg13g2_decap_8 FILLER_55_1495 ();
 sg13g2_decap_8 FILLER_55_1521 ();
 sg13g2_decap_8 FILLER_55_1533 ();
 sg13g2_decap_8 FILLER_55_1540 ();
 sg13g2_fill_1 FILLER_55_1547 ();
 sg13g2_decap_8 FILLER_55_1574 ();
 sg13g2_decap_8 FILLER_55_1581 ();
 sg13g2_decap_8 FILLER_55_1588 ();
 sg13g2_decap_8 FILLER_55_1595 ();
 sg13g2_decap_8 FILLER_55_1602 ();
 sg13g2_decap_8 FILLER_55_1609 ();
 sg13g2_decap_8 FILLER_55_1616 ();
 sg13g2_fill_2 FILLER_55_1623 ();
 sg13g2_fill_1 FILLER_55_1625 ();
 sg13g2_decap_8 FILLER_55_1662 ();
 sg13g2_decap_8 FILLER_55_1669 ();
 sg13g2_decap_8 FILLER_55_1676 ();
 sg13g2_fill_1 FILLER_55_1683 ();
 sg13g2_decap_8 FILLER_55_1698 ();
 sg13g2_fill_2 FILLER_55_1705 ();
 sg13g2_fill_1 FILLER_55_1707 ();
 sg13g2_decap_8 FILLER_55_1720 ();
 sg13g2_decap_8 FILLER_55_1727 ();
 sg13g2_fill_1 FILLER_55_1734 ();
 sg13g2_decap_8 FILLER_55_1745 ();
 sg13g2_decap_8 FILLER_55_1752 ();
 sg13g2_fill_2 FILLER_55_1759 ();
 sg13g2_decap_8 FILLER_55_1821 ();
 sg13g2_decap_8 FILLER_55_1828 ();
 sg13g2_decap_8 FILLER_55_1835 ();
 sg13g2_decap_8 FILLER_55_1842 ();
 sg13g2_fill_2 FILLER_55_1849 ();
 sg13g2_fill_1 FILLER_55_1851 ();
 sg13g2_decap_8 FILLER_55_1860 ();
 sg13g2_decap_8 FILLER_55_1867 ();
 sg13g2_decap_4 FILLER_55_1874 ();
 sg13g2_fill_1 FILLER_55_1878 ();
 sg13g2_fill_2 FILLER_55_1887 ();
 sg13g2_fill_1 FILLER_55_1889 ();
 sg13g2_decap_8 FILLER_55_1896 ();
 sg13g2_decap_4 FILLER_55_1903 ();
 sg13g2_fill_2 FILLER_55_1907 ();
 sg13g2_decap_4 FILLER_55_1924 ();
 sg13g2_fill_1 FILLER_55_1928 ();
 sg13g2_decap_8 FILLER_55_1960 ();
 sg13g2_decap_8 FILLER_55_1967 ();
 sg13g2_decap_8 FILLER_55_1974 ();
 sg13g2_decap_8 FILLER_55_1981 ();
 sg13g2_decap_4 FILLER_55_1988 ();
 sg13g2_fill_2 FILLER_55_1992 ();
 sg13g2_decap_8 FILLER_55_2010 ();
 sg13g2_decap_8 FILLER_55_2017 ();
 sg13g2_fill_1 FILLER_55_2024 ();
 sg13g2_decap_8 FILLER_55_2061 ();
 sg13g2_decap_8 FILLER_55_2068 ();
 sg13g2_decap_8 FILLER_55_2075 ();
 sg13g2_decap_8 FILLER_55_2082 ();
 sg13g2_decap_8 FILLER_55_2089 ();
 sg13g2_decap_8 FILLER_55_2096 ();
 sg13g2_decap_4 FILLER_55_2103 ();
 sg13g2_fill_2 FILLER_55_2125 ();
 sg13g2_decap_8 FILLER_55_2137 ();
 sg13g2_decap_8 FILLER_55_2144 ();
 sg13g2_decap_8 FILLER_55_2151 ();
 sg13g2_decap_8 FILLER_55_2158 ();
 sg13g2_decap_8 FILLER_55_2165 ();
 sg13g2_fill_2 FILLER_55_2172 ();
 sg13g2_decap_8 FILLER_55_2184 ();
 sg13g2_decap_8 FILLER_55_2191 ();
 sg13g2_decap_8 FILLER_55_2198 ();
 sg13g2_decap_8 FILLER_55_2205 ();
 sg13g2_decap_8 FILLER_55_2212 ();
 sg13g2_fill_2 FILLER_55_2219 ();
 sg13g2_decap_8 FILLER_55_2255 ();
 sg13g2_fill_1 FILLER_55_2262 ();
 sg13g2_fill_2 FILLER_55_2299 ();
 sg13g2_decap_8 FILLER_55_2327 ();
 sg13g2_fill_2 FILLER_55_2334 ();
 sg13g2_fill_1 FILLER_55_2336 ();
 sg13g2_decap_8 FILLER_55_2350 ();
 sg13g2_decap_8 FILLER_55_2357 ();
 sg13g2_decap_8 FILLER_55_2364 ();
 sg13g2_decap_8 FILLER_55_2371 ();
 sg13g2_decap_8 FILLER_55_2378 ();
 sg13g2_decap_8 FILLER_55_2385 ();
 sg13g2_fill_2 FILLER_55_2392 ();
 sg13g2_fill_1 FILLER_55_2394 ();
 sg13g2_decap_8 FILLER_55_2401 ();
 sg13g2_decap_8 FILLER_55_2408 ();
 sg13g2_decap_8 FILLER_55_2415 ();
 sg13g2_decap_8 FILLER_55_2422 ();
 sg13g2_decap_8 FILLER_55_2429 ();
 sg13g2_decap_8 FILLER_55_2436 ();
 sg13g2_decap_8 FILLER_55_2443 ();
 sg13g2_fill_2 FILLER_55_2450 ();
 sg13g2_decap_8 FILLER_55_2476 ();
 sg13g2_decap_4 FILLER_55_2483 ();
 sg13g2_decap_4 FILLER_55_2549 ();
 sg13g2_fill_1 FILLER_55_2553 ();
 sg13g2_decap_8 FILLER_55_2559 ();
 sg13g2_decap_4 FILLER_55_2566 ();
 sg13g2_decap_8 FILLER_55_2580 ();
 sg13g2_decap_8 FILLER_55_2587 ();
 sg13g2_decap_8 FILLER_55_2594 ();
 sg13g2_decap_4 FILLER_55_2601 ();
 sg13g2_fill_1 FILLER_55_2605 ();
 sg13g2_decap_8 FILLER_55_2616 ();
 sg13g2_decap_4 FILLER_55_2623 ();
 sg13g2_decap_8 FILLER_55_2635 ();
 sg13g2_decap_8 FILLER_55_2642 ();
 sg13g2_decap_8 FILLER_55_2649 ();
 sg13g2_decap_8 FILLER_55_2656 ();
 sg13g2_decap_8 FILLER_55_2663 ();
 sg13g2_decap_8 FILLER_55_2670 ();
 sg13g2_decap_4 FILLER_55_2677 ();
 sg13g2_fill_1 FILLER_55_2681 ();
 sg13g2_decap_8 FILLER_55_2690 ();
 sg13g2_decap_8 FILLER_55_2697 ();
 sg13g2_decap_8 FILLER_55_2704 ();
 sg13g2_decap_8 FILLER_55_2711 ();
 sg13g2_decap_8 FILLER_55_2718 ();
 sg13g2_decap_8 FILLER_55_2725 ();
 sg13g2_decap_8 FILLER_55_2732 ();
 sg13g2_decap_8 FILLER_55_2739 ();
 sg13g2_decap_8 FILLER_55_2746 ();
 sg13g2_fill_2 FILLER_55_2753 ();
 sg13g2_decap_8 FILLER_55_2791 ();
 sg13g2_decap_8 FILLER_55_2798 ();
 sg13g2_decap_8 FILLER_55_2805 ();
 sg13g2_decap_8 FILLER_55_2812 ();
 sg13g2_fill_1 FILLER_55_2819 ();
 sg13g2_decap_8 FILLER_55_2846 ();
 sg13g2_fill_2 FILLER_55_2853 ();
 sg13g2_fill_1 FILLER_55_2855 ();
 sg13g2_decap_8 FILLER_55_2900 ();
 sg13g2_decap_8 FILLER_55_2907 ();
 sg13g2_decap_8 FILLER_55_2924 ();
 sg13g2_decap_8 FILLER_55_2931 ();
 sg13g2_decap_8 FILLER_55_2938 ();
 sg13g2_decap_8 FILLER_55_2945 ();
 sg13g2_decap_8 FILLER_55_2952 ();
 sg13g2_decap_8 FILLER_55_2959 ();
 sg13g2_fill_2 FILLER_55_2966 ();
 sg13g2_decap_8 FILLER_55_2976 ();
 sg13g2_decap_8 FILLER_55_2983 ();
 sg13g2_decap_8 FILLER_55_2990 ();
 sg13g2_decap_8 FILLER_55_2997 ();
 sg13g2_decap_8 FILLER_55_3004 ();
 sg13g2_decap_8 FILLER_55_3011 ();
 sg13g2_decap_8 FILLER_55_3018 ();
 sg13g2_decap_4 FILLER_55_3025 ();
 sg13g2_decap_8 FILLER_55_3039 ();
 sg13g2_decap_8 FILLER_55_3046 ();
 sg13g2_decap_4 FILLER_55_3053 ();
 sg13g2_fill_2 FILLER_55_3057 ();
 sg13g2_decap_8 FILLER_55_3062 ();
 sg13g2_decap_8 FILLER_55_3069 ();
 sg13g2_decap_8 FILLER_55_3076 ();
 sg13g2_fill_2 FILLER_55_3083 ();
 sg13g2_fill_1 FILLER_55_3085 ();
 sg13g2_decap_8 FILLER_55_3120 ();
 sg13g2_decap_4 FILLER_55_3127 ();
 sg13g2_fill_2 FILLER_55_3131 ();
 sg13g2_decap_8 FILLER_55_3138 ();
 sg13g2_fill_1 FILLER_55_3149 ();
 sg13g2_fill_2 FILLER_55_3155 ();
 sg13g2_fill_1 FILLER_55_3157 ();
 sg13g2_fill_2 FILLER_55_3168 ();
 sg13g2_decap_8 FILLER_55_3180 ();
 sg13g2_decap_8 FILLER_55_3187 ();
 sg13g2_decap_8 FILLER_55_3194 ();
 sg13g2_decap_8 FILLER_55_3201 ();
 sg13g2_decap_8 FILLER_55_3216 ();
 sg13g2_decap_8 FILLER_55_3223 ();
 sg13g2_decap_8 FILLER_55_3230 ();
 sg13g2_decap_8 FILLER_55_3237 ();
 sg13g2_decap_8 FILLER_55_3244 ();
 sg13g2_decap_8 FILLER_55_3251 ();
 sg13g2_decap_8 FILLER_55_3258 ();
 sg13g2_decap_8 FILLER_55_3265 ();
 sg13g2_decap_4 FILLER_55_3272 ();
 sg13g2_decap_8 FILLER_55_3282 ();
 sg13g2_decap_8 FILLER_55_3289 ();
 sg13g2_decap_8 FILLER_55_3296 ();
 sg13g2_decap_8 FILLER_55_3303 ();
 sg13g2_decap_8 FILLER_55_3310 ();
 sg13g2_decap_8 FILLER_55_3317 ();
 sg13g2_decap_8 FILLER_55_3324 ();
 sg13g2_decap_8 FILLER_55_3331 ();
 sg13g2_decap_8 FILLER_55_3338 ();
 sg13g2_decap_8 FILLER_55_3345 ();
 sg13g2_decap_8 FILLER_55_3352 ();
 sg13g2_decap_8 FILLER_55_3359 ();
 sg13g2_decap_8 FILLER_55_3366 ();
 sg13g2_decap_8 FILLER_55_3373 ();
 sg13g2_decap_4 FILLER_55_3380 ();
 sg13g2_fill_1 FILLER_55_3384 ();
 sg13g2_decap_8 FILLER_55_3391 ();
 sg13g2_decap_8 FILLER_55_3398 ();
 sg13g2_decap_8 FILLER_55_3405 ();
 sg13g2_decap_8 FILLER_55_3412 ();
 sg13g2_fill_2 FILLER_55_3419 ();
 sg13g2_fill_1 FILLER_55_3421 ();
 sg13g2_decap_8 FILLER_55_3426 ();
 sg13g2_fill_1 FILLER_55_3433 ();
 sg13g2_decap_8 FILLER_55_3449 ();
 sg13g2_decap_8 FILLER_55_3456 ();
 sg13g2_decap_8 FILLER_55_3463 ();
 sg13g2_decap_8 FILLER_55_3470 ();
 sg13g2_decap_8 FILLER_55_3503 ();
 sg13g2_decap_8 FILLER_55_3510 ();
 sg13g2_decap_8 FILLER_55_3517 ();
 sg13g2_decap_8 FILLER_55_3554 ();
 sg13g2_decap_8 FILLER_55_3561 ();
 sg13g2_decap_8 FILLER_55_3568 ();
 sg13g2_decap_4 FILLER_55_3575 ();
 sg13g2_fill_1 FILLER_55_3579 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_decap_8 FILLER_56_7 ();
 sg13g2_decap_8 FILLER_56_14 ();
 sg13g2_decap_8 FILLER_56_21 ();
 sg13g2_decap_8 FILLER_56_28 ();
 sg13g2_decap_8 FILLER_56_35 ();
 sg13g2_decap_8 FILLER_56_42 ();
 sg13g2_decap_8 FILLER_56_49 ();
 sg13g2_decap_8 FILLER_56_56 ();
 sg13g2_decap_8 FILLER_56_63 ();
 sg13g2_decap_8 FILLER_56_70 ();
 sg13g2_decap_8 FILLER_56_77 ();
 sg13g2_decap_8 FILLER_56_84 ();
 sg13g2_decap_8 FILLER_56_91 ();
 sg13g2_decap_4 FILLER_56_98 ();
 sg13g2_fill_2 FILLER_56_102 ();
 sg13g2_decap_4 FILLER_56_107 ();
 sg13g2_fill_1 FILLER_56_111 ();
 sg13g2_decap_8 FILLER_56_115 ();
 sg13g2_decap_4 FILLER_56_122 ();
 sg13g2_decap_8 FILLER_56_152 ();
 sg13g2_decap_8 FILLER_56_159 ();
 sg13g2_decap_8 FILLER_56_166 ();
 sg13g2_decap_8 FILLER_56_173 ();
 sg13g2_decap_4 FILLER_56_180 ();
 sg13g2_fill_2 FILLER_56_184 ();
 sg13g2_decap_8 FILLER_56_203 ();
 sg13g2_decap_8 FILLER_56_210 ();
 sg13g2_decap_8 FILLER_56_217 ();
 sg13g2_decap_8 FILLER_56_224 ();
 sg13g2_decap_8 FILLER_56_231 ();
 sg13g2_decap_8 FILLER_56_238 ();
 sg13g2_fill_2 FILLER_56_245 ();
 sg13g2_fill_2 FILLER_56_266 ();
 sg13g2_decap_8 FILLER_56_278 ();
 sg13g2_decap_8 FILLER_56_285 ();
 sg13g2_decap_8 FILLER_56_292 ();
 sg13g2_decap_4 FILLER_56_299 ();
 sg13g2_fill_1 FILLER_56_303 ();
 sg13g2_decap_8 FILLER_56_334 ();
 sg13g2_decap_4 FILLER_56_341 ();
 sg13g2_fill_1 FILLER_56_345 ();
 sg13g2_decap_8 FILLER_56_351 ();
 sg13g2_decap_8 FILLER_56_358 ();
 sg13g2_fill_2 FILLER_56_365 ();
 sg13g2_decap_4 FILLER_56_372 ();
 sg13g2_fill_1 FILLER_56_376 ();
 sg13g2_fill_1 FILLER_56_387 ();
 sg13g2_decap_4 FILLER_56_400 ();
 sg13g2_fill_1 FILLER_56_404 ();
 sg13g2_decap_8 FILLER_56_413 ();
 sg13g2_decap_8 FILLER_56_420 ();
 sg13g2_decap_8 FILLER_56_427 ();
 sg13g2_decap_8 FILLER_56_434 ();
 sg13g2_decap_8 FILLER_56_441 ();
 sg13g2_fill_2 FILLER_56_448 ();
 sg13g2_fill_1 FILLER_56_450 ();
 sg13g2_decap_4 FILLER_56_477 ();
 sg13g2_fill_2 FILLER_56_487 ();
 sg13g2_fill_2 FILLER_56_494 ();
 sg13g2_fill_1 FILLER_56_504 ();
 sg13g2_decap_4 FILLER_56_510 ();
 sg13g2_fill_2 FILLER_56_514 ();
 sg13g2_decap_8 FILLER_56_522 ();
 sg13g2_decap_8 FILLER_56_529 ();
 sg13g2_decap_4 FILLER_56_549 ();
 sg13g2_fill_2 FILLER_56_558 ();
 sg13g2_decap_8 FILLER_56_573 ();
 sg13g2_decap_8 FILLER_56_580 ();
 sg13g2_decap_8 FILLER_56_587 ();
 sg13g2_decap_4 FILLER_56_594 ();
 sg13g2_fill_1 FILLER_56_598 ();
 sg13g2_fill_2 FILLER_56_623 ();
 sg13g2_decap_4 FILLER_56_639 ();
 sg13g2_decap_8 FILLER_56_648 ();
 sg13g2_decap_8 FILLER_56_655 ();
 sg13g2_fill_2 FILLER_56_662 ();
 sg13g2_decap_8 FILLER_56_675 ();
 sg13g2_decap_4 FILLER_56_682 ();
 sg13g2_decap_8 FILLER_56_691 ();
 sg13g2_decap_8 FILLER_56_698 ();
 sg13g2_decap_4 FILLER_56_705 ();
 sg13g2_decap_8 FILLER_56_719 ();
 sg13g2_decap_4 FILLER_56_726 ();
 sg13g2_fill_2 FILLER_56_730 ();
 sg13g2_decap_4 FILLER_56_740 ();
 sg13g2_fill_1 FILLER_56_744 ();
 sg13g2_decap_8 FILLER_56_753 ();
 sg13g2_decap_4 FILLER_56_760 ();
 sg13g2_fill_1 FILLER_56_764 ();
 sg13g2_decap_8 FILLER_56_780 ();
 sg13g2_decap_8 FILLER_56_787 ();
 sg13g2_decap_8 FILLER_56_794 ();
 sg13g2_decap_8 FILLER_56_801 ();
 sg13g2_fill_2 FILLER_56_808 ();
 sg13g2_decap_8 FILLER_56_818 ();
 sg13g2_fill_2 FILLER_56_825 ();
 sg13g2_decap_8 FILLER_56_839 ();
 sg13g2_decap_8 FILLER_56_846 ();
 sg13g2_decap_8 FILLER_56_853 ();
 sg13g2_decap_4 FILLER_56_860 ();
 sg13g2_decap_8 FILLER_56_872 ();
 sg13g2_decap_8 FILLER_56_879 ();
 sg13g2_fill_2 FILLER_56_886 ();
 sg13g2_fill_1 FILLER_56_888 ();
 sg13g2_decap_8 FILLER_56_896 ();
 sg13g2_decap_8 FILLER_56_903 ();
 sg13g2_decap_8 FILLER_56_910 ();
 sg13g2_decap_8 FILLER_56_917 ();
 sg13g2_decap_8 FILLER_56_924 ();
 sg13g2_decap_8 FILLER_56_931 ();
 sg13g2_decap_4 FILLER_56_938 ();
 sg13g2_fill_1 FILLER_56_942 ();
 sg13g2_fill_1 FILLER_56_956 ();
 sg13g2_decap_8 FILLER_56_973 ();
 sg13g2_decap_8 FILLER_56_980 ();
 sg13g2_decap_8 FILLER_56_987 ();
 sg13g2_decap_8 FILLER_56_994 ();
 sg13g2_fill_2 FILLER_56_1001 ();
 sg13g2_fill_1 FILLER_56_1003 ();
 sg13g2_decap_8 FILLER_56_1008 ();
 sg13g2_decap_8 FILLER_56_1015 ();
 sg13g2_decap_4 FILLER_56_1022 ();
 sg13g2_fill_2 FILLER_56_1026 ();
 sg13g2_decap_8 FILLER_56_1036 ();
 sg13g2_decap_8 FILLER_56_1043 ();
 sg13g2_decap_8 FILLER_56_1050 ();
 sg13g2_decap_8 FILLER_56_1057 ();
 sg13g2_decap_8 FILLER_56_1064 ();
 sg13g2_decap_8 FILLER_56_1071 ();
 sg13g2_decap_8 FILLER_56_1078 ();
 sg13g2_decap_8 FILLER_56_1085 ();
 sg13g2_decap_8 FILLER_56_1092 ();
 sg13g2_decap_8 FILLER_56_1099 ();
 sg13g2_fill_1 FILLER_56_1106 ();
 sg13g2_decap_8 FILLER_56_1169 ();
 sg13g2_decap_8 FILLER_56_1176 ();
 sg13g2_decap_4 FILLER_56_1183 ();
 sg13g2_fill_1 FILLER_56_1187 ();
 sg13g2_fill_2 FILLER_56_1198 ();
 sg13g2_decap_8 FILLER_56_1210 ();
 sg13g2_decap_8 FILLER_56_1217 ();
 sg13g2_decap_8 FILLER_56_1224 ();
 sg13g2_decap_8 FILLER_56_1231 ();
 sg13g2_decap_8 FILLER_56_1238 ();
 sg13g2_decap_8 FILLER_56_1245 ();
 sg13g2_decap_8 FILLER_56_1252 ();
 sg13g2_fill_2 FILLER_56_1259 ();
 sg13g2_decap_4 FILLER_56_1266 ();
 sg13g2_fill_2 FILLER_56_1270 ();
 sg13g2_decap_4 FILLER_56_1311 ();
 sg13g2_fill_2 FILLER_56_1315 ();
 sg13g2_decap_8 FILLER_56_1326 ();
 sg13g2_decap_8 FILLER_56_1333 ();
 sg13g2_decap_8 FILLER_56_1340 ();
 sg13g2_decap_4 FILLER_56_1347 ();
 sg13g2_fill_2 FILLER_56_1351 ();
 sg13g2_fill_2 FILLER_56_1363 ();
 sg13g2_fill_1 FILLER_56_1365 ();
 sg13g2_decap_8 FILLER_56_1392 ();
 sg13g2_decap_8 FILLER_56_1399 ();
 sg13g2_decap_8 FILLER_56_1406 ();
 sg13g2_decap_8 FILLER_56_1413 ();
 sg13g2_decap_8 FILLER_56_1420 ();
 sg13g2_decap_8 FILLER_56_1427 ();
 sg13g2_decap_8 FILLER_56_1434 ();
 sg13g2_decap_8 FILLER_56_1441 ();
 sg13g2_decap_8 FILLER_56_1448 ();
 sg13g2_decap_8 FILLER_56_1455 ();
 sg13g2_fill_2 FILLER_56_1462 ();
 sg13g2_fill_1 FILLER_56_1464 ();
 sg13g2_fill_1 FILLER_56_1473 ();
 sg13g2_decap_8 FILLER_56_1499 ();
 sg13g2_decap_8 FILLER_56_1506 ();
 sg13g2_decap_8 FILLER_56_1513 ();
 sg13g2_decap_8 FILLER_56_1520 ();
 sg13g2_decap_8 FILLER_56_1527 ();
 sg13g2_decap_8 FILLER_56_1534 ();
 sg13g2_fill_2 FILLER_56_1541 ();
 sg13g2_decap_8 FILLER_56_1569 ();
 sg13g2_decap_4 FILLER_56_1576 ();
 sg13g2_fill_1 FILLER_56_1580 ();
 sg13g2_fill_2 FILLER_56_1587 ();
 sg13g2_decap_8 FILLER_56_1603 ();
 sg13g2_decap_8 FILLER_56_1610 ();
 sg13g2_decap_8 FILLER_56_1617 ();
 sg13g2_decap_8 FILLER_56_1624 ();
 sg13g2_decap_8 FILLER_56_1631 ();
 sg13g2_decap_8 FILLER_56_1638 ();
 sg13g2_decap_8 FILLER_56_1645 ();
 sg13g2_decap_8 FILLER_56_1652 ();
 sg13g2_decap_8 FILLER_56_1659 ();
 sg13g2_decap_8 FILLER_56_1666 ();
 sg13g2_decap_8 FILLER_56_1673 ();
 sg13g2_decap_8 FILLER_56_1680 ();
 sg13g2_decap_8 FILLER_56_1687 ();
 sg13g2_decap_8 FILLER_56_1702 ();
 sg13g2_decap_8 FILLER_56_1709 ();
 sg13g2_decap_8 FILLER_56_1716 ();
 sg13g2_decap_8 FILLER_56_1733 ();
 sg13g2_decap_8 FILLER_56_1740 ();
 sg13g2_decap_8 FILLER_56_1747 ();
 sg13g2_decap_8 FILLER_56_1754 ();
 sg13g2_fill_1 FILLER_56_1761 ();
 sg13g2_decap_8 FILLER_56_1770 ();
 sg13g2_decap_8 FILLER_56_1816 ();
 sg13g2_decap_4 FILLER_56_1823 ();
 sg13g2_fill_2 FILLER_56_1827 ();
 sg13g2_decap_8 FILLER_56_1865 ();
 sg13g2_fill_2 FILLER_56_1872 ();
 sg13g2_decap_8 FILLER_56_1890 ();
 sg13g2_fill_2 FILLER_56_1897 ();
 sg13g2_decap_8 FILLER_56_1925 ();
 sg13g2_decap_4 FILLER_56_1932 ();
 sg13g2_fill_2 FILLER_56_1936 ();
 sg13g2_decap_8 FILLER_56_1948 ();
 sg13g2_fill_2 FILLER_56_1955 ();
 sg13g2_fill_1 FILLER_56_1957 ();
 sg13g2_decap_8 FILLER_56_1984 ();
 sg13g2_decap_8 FILLER_56_1991 ();
 sg13g2_decap_8 FILLER_56_1998 ();
 sg13g2_decap_8 FILLER_56_2005 ();
 sg13g2_decap_8 FILLER_56_2012 ();
 sg13g2_decap_4 FILLER_56_2019 ();
 sg13g2_fill_2 FILLER_56_2023 ();
 sg13g2_decap_8 FILLER_56_2033 ();
 sg13g2_decap_8 FILLER_56_2040 ();
 sg13g2_decap_8 FILLER_56_2047 ();
 sg13g2_fill_2 FILLER_56_2054 ();
 sg13g2_fill_1 FILLER_56_2056 ();
 sg13g2_decap_8 FILLER_56_2083 ();
 sg13g2_decap_8 FILLER_56_2090 ();
 sg13g2_decap_8 FILLER_56_2097 ();
 sg13g2_decap_8 FILLER_56_2104 ();
 sg13g2_decap_4 FILLER_56_2111 ();
 sg13g2_decap_4 FILLER_56_2127 ();
 sg13g2_fill_1 FILLER_56_2131 ();
 sg13g2_decap_8 FILLER_56_2158 ();
 sg13g2_decap_8 FILLER_56_2165 ();
 sg13g2_decap_4 FILLER_56_2172 ();
 sg13g2_fill_1 FILLER_56_2176 ();
 sg13g2_fill_2 FILLER_56_2183 ();
 sg13g2_decap_8 FILLER_56_2191 ();
 sg13g2_decap_4 FILLER_56_2198 ();
 sg13g2_fill_1 FILLER_56_2202 ();
 sg13g2_decap_8 FILLER_56_2209 ();
 sg13g2_decap_8 FILLER_56_2216 ();
 sg13g2_fill_2 FILLER_56_2223 ();
 sg13g2_decap_4 FILLER_56_2263 ();
 sg13g2_fill_2 FILLER_56_2267 ();
 sg13g2_decap_8 FILLER_56_2275 ();
 sg13g2_decap_8 FILLER_56_2282 ();
 sg13g2_decap_8 FILLER_56_2289 ();
 sg13g2_fill_1 FILLER_56_2296 ();
 sg13g2_decap_8 FILLER_56_2307 ();
 sg13g2_decap_8 FILLER_56_2314 ();
 sg13g2_decap_8 FILLER_56_2321 ();
 sg13g2_decap_8 FILLER_56_2328 ();
 sg13g2_decap_4 FILLER_56_2335 ();
 sg13g2_decap_8 FILLER_56_2375 ();
 sg13g2_decap_8 FILLER_56_2382 ();
 sg13g2_decap_8 FILLER_56_2389 ();
 sg13g2_decap_8 FILLER_56_2396 ();
 sg13g2_decap_8 FILLER_56_2407 ();
 sg13g2_decap_8 FILLER_56_2414 ();
 sg13g2_decap_8 FILLER_56_2421 ();
 sg13g2_decap_8 FILLER_56_2428 ();
 sg13g2_decap_8 FILLER_56_2435 ();
 sg13g2_fill_1 FILLER_56_2442 ();
 sg13g2_fill_1 FILLER_56_2456 ();
 sg13g2_decap_8 FILLER_56_2476 ();
 sg13g2_decap_8 FILLER_56_2483 ();
 sg13g2_decap_8 FILLER_56_2490 ();
 sg13g2_decap_8 FILLER_56_2497 ();
 sg13g2_decap_8 FILLER_56_2504 ();
 sg13g2_decap_4 FILLER_56_2511 ();
 sg13g2_decap_8 FILLER_56_2541 ();
 sg13g2_decap_8 FILLER_56_2548 ();
 sg13g2_decap_8 FILLER_56_2555 ();
 sg13g2_decap_8 FILLER_56_2562 ();
 sg13g2_decap_8 FILLER_56_2569 ();
 sg13g2_decap_8 FILLER_56_2576 ();
 sg13g2_decap_8 FILLER_56_2583 ();
 sg13g2_decap_8 FILLER_56_2590 ();
 sg13g2_decap_8 FILLER_56_2597 ();
 sg13g2_decap_8 FILLER_56_2604 ();
 sg13g2_decap_8 FILLER_56_2611 ();
 sg13g2_decap_8 FILLER_56_2618 ();
 sg13g2_decap_8 FILLER_56_2625 ();
 sg13g2_decap_8 FILLER_56_2632 ();
 sg13g2_decap_8 FILLER_56_2639 ();
 sg13g2_decap_8 FILLER_56_2646 ();
 sg13g2_decap_8 FILLER_56_2653 ();
 sg13g2_fill_2 FILLER_56_2660 ();
 sg13g2_fill_1 FILLER_56_2662 ();
 sg13g2_decap_8 FILLER_56_2689 ();
 sg13g2_fill_2 FILLER_56_2696 ();
 sg13g2_decap_8 FILLER_56_2714 ();
 sg13g2_decap_8 FILLER_56_2721 ();
 sg13g2_decap_8 FILLER_56_2728 ();
 sg13g2_fill_2 FILLER_56_2735 ();
 sg13g2_fill_1 FILLER_56_2737 ();
 sg13g2_decap_8 FILLER_56_2748 ();
 sg13g2_decap_8 FILLER_56_2755 ();
 sg13g2_decap_4 FILLER_56_2762 ();
 sg13g2_fill_1 FILLER_56_2766 ();
 sg13g2_decap_8 FILLER_56_2772 ();
 sg13g2_decap_8 FILLER_56_2779 ();
 sg13g2_decap_8 FILLER_56_2786 ();
 sg13g2_decap_8 FILLER_56_2793 ();
 sg13g2_decap_4 FILLER_56_2800 ();
 sg13g2_fill_1 FILLER_56_2804 ();
 sg13g2_decap_8 FILLER_56_2841 ();
 sg13g2_decap_8 FILLER_56_2848 ();
 sg13g2_decap_8 FILLER_56_2855 ();
 sg13g2_decap_8 FILLER_56_2862 ();
 sg13g2_decap_8 FILLER_56_2869 ();
 sg13g2_decap_4 FILLER_56_2876 ();
 sg13g2_fill_2 FILLER_56_2880 ();
 sg13g2_decap_4 FILLER_56_2887 ();
 sg13g2_fill_1 FILLER_56_2891 ();
 sg13g2_decap_8 FILLER_56_2897 ();
 sg13g2_decap_8 FILLER_56_2904 ();
 sg13g2_decap_8 FILLER_56_2911 ();
 sg13g2_decap_8 FILLER_56_2918 ();
 sg13g2_decap_4 FILLER_56_2925 ();
 sg13g2_fill_2 FILLER_56_2929 ();
 sg13g2_decap_8 FILLER_56_2957 ();
 sg13g2_decap_8 FILLER_56_2964 ();
 sg13g2_decap_8 FILLER_56_2971 ();
 sg13g2_decap_4 FILLER_56_2978 ();
 sg13g2_fill_1 FILLER_56_2982 ();
 sg13g2_decap_8 FILLER_56_2996 ();
 sg13g2_decap_8 FILLER_56_3003 ();
 sg13g2_decap_4 FILLER_56_3010 ();
 sg13g2_fill_1 FILLER_56_3014 ();
 sg13g2_decap_4 FILLER_56_3025 ();
 sg13g2_fill_1 FILLER_56_3029 ();
 sg13g2_decap_8 FILLER_56_3035 ();
 sg13g2_decap_8 FILLER_56_3050 ();
 sg13g2_decap_8 FILLER_56_3057 ();
 sg13g2_decap_8 FILLER_56_3064 ();
 sg13g2_decap_8 FILLER_56_3071 ();
 sg13g2_decap_8 FILLER_56_3078 ();
 sg13g2_decap_8 FILLER_56_3085 ();
 sg13g2_decap_8 FILLER_56_3124 ();
 sg13g2_decap_8 FILLER_56_3131 ();
 sg13g2_decap_8 FILLER_56_3138 ();
 sg13g2_decap_8 FILLER_56_3145 ();
 sg13g2_decap_8 FILLER_56_3152 ();
 sg13g2_decap_8 FILLER_56_3159 ();
 sg13g2_decap_8 FILLER_56_3166 ();
 sg13g2_fill_2 FILLER_56_3173 ();
 sg13g2_fill_1 FILLER_56_3175 ();
 sg13g2_decap_8 FILLER_56_3181 ();
 sg13g2_decap_8 FILLER_56_3188 ();
 sg13g2_fill_2 FILLER_56_3195 ();
 sg13g2_decap_8 FILLER_56_3220 ();
 sg13g2_decap_8 FILLER_56_3227 ();
 sg13g2_decap_8 FILLER_56_3234 ();
 sg13g2_decap_8 FILLER_56_3241 ();
 sg13g2_decap_8 FILLER_56_3248 ();
 sg13g2_decap_8 FILLER_56_3255 ();
 sg13g2_decap_8 FILLER_56_3262 ();
 sg13g2_fill_2 FILLER_56_3269 ();
 sg13g2_decap_8 FILLER_56_3297 ();
 sg13g2_decap_8 FILLER_56_3304 ();
 sg13g2_decap_8 FILLER_56_3311 ();
 sg13g2_decap_8 FILLER_56_3318 ();
 sg13g2_decap_8 FILLER_56_3325 ();
 sg13g2_decap_8 FILLER_56_3332 ();
 sg13g2_decap_8 FILLER_56_3339 ();
 sg13g2_decap_8 FILLER_56_3346 ();
 sg13g2_decap_8 FILLER_56_3353 ();
 sg13g2_decap_8 FILLER_56_3360 ();
 sg13g2_decap_8 FILLER_56_3367 ();
 sg13g2_decap_4 FILLER_56_3374 ();
 sg13g2_fill_1 FILLER_56_3378 ();
 sg13g2_decap_8 FILLER_56_3405 ();
 sg13g2_decap_8 FILLER_56_3412 ();
 sg13g2_fill_1 FILLER_56_3419 ();
 sg13g2_decap_8 FILLER_56_3451 ();
 sg13g2_decap_8 FILLER_56_3458 ();
 sg13g2_fill_2 FILLER_56_3465 ();
 sg13g2_fill_1 FILLER_56_3467 ();
 sg13g2_fill_1 FILLER_56_3494 ();
 sg13g2_decap_8 FILLER_56_3508 ();
 sg13g2_decap_8 FILLER_56_3515 ();
 sg13g2_decap_4 FILLER_56_3522 ();
 sg13g2_fill_1 FILLER_56_3526 ();
 sg13g2_fill_1 FILLER_56_3579 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_decap_8 FILLER_57_7 ();
 sg13g2_decap_8 FILLER_57_14 ();
 sg13g2_decap_8 FILLER_57_21 ();
 sg13g2_fill_1 FILLER_57_28 ();
 sg13g2_decap_8 FILLER_57_33 ();
 sg13g2_decap_8 FILLER_57_40 ();
 sg13g2_decap_8 FILLER_57_47 ();
 sg13g2_decap_8 FILLER_57_54 ();
 sg13g2_decap_8 FILLER_57_61 ();
 sg13g2_decap_8 FILLER_57_68 ();
 sg13g2_decap_8 FILLER_57_75 ();
 sg13g2_decap_8 FILLER_57_82 ();
 sg13g2_decap_8 FILLER_57_89 ();
 sg13g2_fill_2 FILLER_57_96 ();
 sg13g2_decap_8 FILLER_57_103 ();
 sg13g2_decap_8 FILLER_57_110 ();
 sg13g2_decap_8 FILLER_57_117 ();
 sg13g2_fill_2 FILLER_57_124 ();
 sg13g2_fill_1 FILLER_57_126 ();
 sg13g2_decap_8 FILLER_57_170 ();
 sg13g2_fill_1 FILLER_57_177 ();
 sg13g2_decap_8 FILLER_57_230 ();
 sg13g2_fill_2 FILLER_57_237 ();
 sg13g2_fill_1 FILLER_57_239 ();
 sg13g2_decap_8 FILLER_57_274 ();
 sg13g2_decap_8 FILLER_57_281 ();
 sg13g2_decap_8 FILLER_57_288 ();
 sg13g2_decap_8 FILLER_57_295 ();
 sg13g2_decap_8 FILLER_57_302 ();
 sg13g2_fill_1 FILLER_57_309 ();
 sg13g2_decap_8 FILLER_57_316 ();
 sg13g2_fill_2 FILLER_57_323 ();
 sg13g2_decap_8 FILLER_57_332 ();
 sg13g2_decap_8 FILLER_57_339 ();
 sg13g2_decap_8 FILLER_57_346 ();
 sg13g2_decap_8 FILLER_57_353 ();
 sg13g2_decap_8 FILLER_57_360 ();
 sg13g2_decap_8 FILLER_57_367 ();
 sg13g2_decap_8 FILLER_57_374 ();
 sg13g2_decap_8 FILLER_57_381 ();
 sg13g2_decap_8 FILLER_57_388 ();
 sg13g2_decap_8 FILLER_57_395 ();
 sg13g2_decap_8 FILLER_57_402 ();
 sg13g2_decap_8 FILLER_57_409 ();
 sg13g2_decap_8 FILLER_57_416 ();
 sg13g2_decap_8 FILLER_57_423 ();
 sg13g2_decap_8 FILLER_57_430 ();
 sg13g2_decap_8 FILLER_57_443 ();
 sg13g2_decap_8 FILLER_57_450 ();
 sg13g2_decap_8 FILLER_57_457 ();
 sg13g2_decap_8 FILLER_57_464 ();
 sg13g2_decap_4 FILLER_57_471 ();
 sg13g2_decap_8 FILLER_57_480 ();
 sg13g2_fill_2 FILLER_57_490 ();
 sg13g2_fill_1 FILLER_57_492 ();
 sg13g2_fill_2 FILLER_57_498 ();
 sg13g2_fill_1 FILLER_57_500 ();
 sg13g2_decap_8 FILLER_57_507 ();
 sg13g2_decap_8 FILLER_57_514 ();
 sg13g2_decap_4 FILLER_57_521 ();
 sg13g2_decap_8 FILLER_57_551 ();
 sg13g2_decap_8 FILLER_57_558 ();
 sg13g2_fill_2 FILLER_57_565 ();
 sg13g2_decap_8 FILLER_57_572 ();
 sg13g2_decap_8 FILLER_57_579 ();
 sg13g2_decap_8 FILLER_57_586 ();
 sg13g2_decap_8 FILLER_57_593 ();
 sg13g2_decap_8 FILLER_57_600 ();
 sg13g2_decap_8 FILLER_57_607 ();
 sg13g2_decap_4 FILLER_57_614 ();
 sg13g2_decap_8 FILLER_57_633 ();
 sg13g2_decap_8 FILLER_57_640 ();
 sg13g2_decap_8 FILLER_57_647 ();
 sg13g2_decap_4 FILLER_57_654 ();
 sg13g2_fill_2 FILLER_57_658 ();
 sg13g2_decap_8 FILLER_57_704 ();
 sg13g2_decap_8 FILLER_57_711 ();
 sg13g2_decap_8 FILLER_57_718 ();
 sg13g2_decap_8 FILLER_57_725 ();
 sg13g2_decap_8 FILLER_57_732 ();
 sg13g2_decap_8 FILLER_57_739 ();
 sg13g2_decap_8 FILLER_57_746 ();
 sg13g2_decap_4 FILLER_57_753 ();
 sg13g2_fill_2 FILLER_57_757 ();
 sg13g2_decap_4 FILLER_57_764 ();
 sg13g2_fill_2 FILLER_57_768 ();
 sg13g2_decap_8 FILLER_57_778 ();
 sg13g2_decap_4 FILLER_57_785 ();
 sg13g2_fill_1 FILLER_57_789 ();
 sg13g2_decap_8 FILLER_57_795 ();
 sg13g2_decap_8 FILLER_57_802 ();
 sg13g2_fill_1 FILLER_57_809 ();
 sg13g2_decap_8 FILLER_57_814 ();
 sg13g2_decap_8 FILLER_57_821 ();
 sg13g2_decap_8 FILLER_57_828 ();
 sg13g2_fill_2 FILLER_57_835 ();
 sg13g2_decap_8 FILLER_57_843 ();
 sg13g2_fill_2 FILLER_57_850 ();
 sg13g2_decap_4 FILLER_57_856 ();
 sg13g2_decap_8 FILLER_57_878 ();
 sg13g2_fill_1 FILLER_57_885 ();
 sg13g2_fill_1 FILLER_57_907 ();
 sg13g2_decap_8 FILLER_57_920 ();
 sg13g2_decap_4 FILLER_57_927 ();
 sg13g2_fill_1 FILLER_57_931 ();
 sg13g2_fill_1 FILLER_57_940 ();
 sg13g2_decap_8 FILLER_57_977 ();
 sg13g2_decap_8 FILLER_57_984 ();
 sg13g2_decap_4 FILLER_57_991 ();
 sg13g2_fill_1 FILLER_57_995 ();
 sg13g2_decap_8 FILLER_57_1027 ();
 sg13g2_fill_1 FILLER_57_1034 ();
 sg13g2_decap_8 FILLER_57_1043 ();
 sg13g2_decap_8 FILLER_57_1054 ();
 sg13g2_decap_8 FILLER_57_1061 ();
 sg13g2_decap_8 FILLER_57_1068 ();
 sg13g2_decap_8 FILLER_57_1075 ();
 sg13g2_decap_8 FILLER_57_1082 ();
 sg13g2_fill_2 FILLER_57_1089 ();
 sg13g2_fill_1 FILLER_57_1091 ();
 sg13g2_decap_8 FILLER_57_1101 ();
 sg13g2_decap_8 FILLER_57_1108 ();
 sg13g2_decap_8 FILLER_57_1115 ();
 sg13g2_decap_8 FILLER_57_1122 ();
 sg13g2_decap_8 FILLER_57_1129 ();
 sg13g2_decap_8 FILLER_57_1136 ();
 sg13g2_decap_4 FILLER_57_1143 ();
 sg13g2_fill_1 FILLER_57_1147 ();
 sg13g2_decap_8 FILLER_57_1156 ();
 sg13g2_decap_8 FILLER_57_1163 ();
 sg13g2_decap_8 FILLER_57_1170 ();
 sg13g2_decap_8 FILLER_57_1177 ();
 sg13g2_decap_8 FILLER_57_1184 ();
 sg13g2_decap_8 FILLER_57_1191 ();
 sg13g2_decap_8 FILLER_57_1198 ();
 sg13g2_decap_8 FILLER_57_1205 ();
 sg13g2_decap_8 FILLER_57_1212 ();
 sg13g2_decap_8 FILLER_57_1219 ();
 sg13g2_decap_8 FILLER_57_1226 ();
 sg13g2_decap_8 FILLER_57_1233 ();
 sg13g2_decap_8 FILLER_57_1240 ();
 sg13g2_decap_8 FILLER_57_1247 ();
 sg13g2_decap_8 FILLER_57_1254 ();
 sg13g2_decap_8 FILLER_57_1261 ();
 sg13g2_decap_8 FILLER_57_1268 ();
 sg13g2_decap_8 FILLER_57_1275 ();
 sg13g2_decap_4 FILLER_57_1282 ();
 sg13g2_decap_8 FILLER_57_1296 ();
 sg13g2_decap_8 FILLER_57_1312 ();
 sg13g2_decap_8 FILLER_57_1319 ();
 sg13g2_fill_1 FILLER_57_1326 ();
 sg13g2_decap_8 FILLER_57_1337 ();
 sg13g2_decap_8 FILLER_57_1344 ();
 sg13g2_decap_8 FILLER_57_1351 ();
 sg13g2_decap_8 FILLER_57_1358 ();
 sg13g2_decap_8 FILLER_57_1365 ();
 sg13g2_decap_8 FILLER_57_1372 ();
 sg13g2_decap_8 FILLER_57_1379 ();
 sg13g2_decap_8 FILLER_57_1386 ();
 sg13g2_decap_8 FILLER_57_1393 ();
 sg13g2_fill_1 FILLER_57_1400 ();
 sg13g2_decap_8 FILLER_57_1419 ();
 sg13g2_decap_8 FILLER_57_1426 ();
 sg13g2_fill_2 FILLER_57_1433 ();
 sg13g2_fill_1 FILLER_57_1435 ();
 sg13g2_decap_8 FILLER_57_1449 ();
 sg13g2_decap_8 FILLER_57_1456 ();
 sg13g2_decap_8 FILLER_57_1463 ();
 sg13g2_fill_2 FILLER_57_1470 ();
 sg13g2_fill_1 FILLER_57_1472 ();
 sg13g2_decap_8 FILLER_57_1501 ();
 sg13g2_decap_8 FILLER_57_1508 ();
 sg13g2_decap_8 FILLER_57_1515 ();
 sg13g2_decap_8 FILLER_57_1522 ();
 sg13g2_decap_8 FILLER_57_1529 ();
 sg13g2_decap_4 FILLER_57_1536 ();
 sg13g2_fill_1 FILLER_57_1540 ();
 sg13g2_decap_8 FILLER_57_1551 ();
 sg13g2_decap_8 FILLER_57_1558 ();
 sg13g2_decap_8 FILLER_57_1565 ();
 sg13g2_decap_8 FILLER_57_1572 ();
 sg13g2_decap_8 FILLER_57_1579 ();
 sg13g2_fill_2 FILLER_57_1586 ();
 sg13g2_decap_8 FILLER_57_1608 ();
 sg13g2_fill_1 FILLER_57_1615 ();
 sg13g2_fill_2 FILLER_57_1634 ();
 sg13g2_decap_8 FILLER_57_1662 ();
 sg13g2_decap_8 FILLER_57_1669 ();
 sg13g2_fill_2 FILLER_57_1676 ();
 sg13g2_fill_1 FILLER_57_1678 ();
 sg13g2_decap_8 FILLER_57_1695 ();
 sg13g2_decap_8 FILLER_57_1702 ();
 sg13g2_decap_4 FILLER_57_1709 ();
 sg13g2_fill_2 FILLER_57_1713 ();
 sg13g2_decap_8 FILLER_57_1741 ();
 sg13g2_decap_8 FILLER_57_1748 ();
 sg13g2_decap_8 FILLER_57_1755 ();
 sg13g2_fill_2 FILLER_57_1762 ();
 sg13g2_fill_1 FILLER_57_1785 ();
 sg13g2_decap_4 FILLER_57_1789 ();
 sg13g2_fill_2 FILLER_57_1793 ();
 sg13g2_decap_8 FILLER_57_1817 ();
 sg13g2_decap_8 FILLER_57_1824 ();
 sg13g2_decap_8 FILLER_57_1831 ();
 sg13g2_decap_8 FILLER_57_1838 ();
 sg13g2_decap_8 FILLER_57_1845 ();
 sg13g2_decap_8 FILLER_57_1852 ();
 sg13g2_decap_8 FILLER_57_1859 ();
 sg13g2_decap_8 FILLER_57_1866 ();
 sg13g2_decap_8 FILLER_57_1873 ();
 sg13g2_decap_8 FILLER_57_1880 ();
 sg13g2_decap_8 FILLER_57_1887 ();
 sg13g2_decap_8 FILLER_57_1894 ();
 sg13g2_decap_8 FILLER_57_1901 ();
 sg13g2_decap_8 FILLER_57_1908 ();
 sg13g2_decap_8 FILLER_57_1915 ();
 sg13g2_decap_8 FILLER_57_1922 ();
 sg13g2_decap_8 FILLER_57_1929 ();
 sg13g2_decap_8 FILLER_57_1936 ();
 sg13g2_decap_8 FILLER_57_1943 ();
 sg13g2_fill_2 FILLER_57_1950 ();
 sg13g2_decap_8 FILLER_57_1984 ();
 sg13g2_decap_8 FILLER_57_1991 ();
 sg13g2_decap_8 FILLER_57_2004 ();
 sg13g2_decap_8 FILLER_57_2011 ();
 sg13g2_decap_8 FILLER_57_2018 ();
 sg13g2_decap_4 FILLER_57_2025 ();
 sg13g2_decap_8 FILLER_57_2034 ();
 sg13g2_decap_8 FILLER_57_2041 ();
 sg13g2_decap_8 FILLER_57_2048 ();
 sg13g2_decap_8 FILLER_57_2055 ();
 sg13g2_decap_8 FILLER_57_2072 ();
 sg13g2_decap_8 FILLER_57_2079 ();
 sg13g2_decap_8 FILLER_57_2086 ();
 sg13g2_decap_8 FILLER_57_2093 ();
 sg13g2_decap_8 FILLER_57_2100 ();
 sg13g2_decap_8 FILLER_57_2107 ();
 sg13g2_decap_8 FILLER_57_2114 ();
 sg13g2_decap_4 FILLER_57_2121 ();
 sg13g2_fill_1 FILLER_57_2125 ();
 sg13g2_decap_8 FILLER_57_2134 ();
 sg13g2_decap_8 FILLER_57_2141 ();
 sg13g2_decap_8 FILLER_57_2148 ();
 sg13g2_decap_8 FILLER_57_2155 ();
 sg13g2_decap_8 FILLER_57_2162 ();
 sg13g2_decap_4 FILLER_57_2169 ();
 sg13g2_fill_1 FILLER_57_2173 ();
 sg13g2_decap_8 FILLER_57_2206 ();
 sg13g2_decap_8 FILLER_57_2213 ();
 sg13g2_decap_4 FILLER_57_2220 ();
 sg13g2_fill_2 FILLER_57_2224 ();
 sg13g2_decap_8 FILLER_57_2243 ();
 sg13g2_decap_8 FILLER_57_2250 ();
 sg13g2_decap_8 FILLER_57_2257 ();
 sg13g2_decap_8 FILLER_57_2264 ();
 sg13g2_decap_8 FILLER_57_2271 ();
 sg13g2_decap_8 FILLER_57_2278 ();
 sg13g2_decap_4 FILLER_57_2285 ();
 sg13g2_fill_1 FILLER_57_2297 ();
 sg13g2_decap_8 FILLER_57_2310 ();
 sg13g2_decap_8 FILLER_57_2317 ();
 sg13g2_decap_8 FILLER_57_2324 ();
 sg13g2_decap_8 FILLER_57_2331 ();
 sg13g2_decap_8 FILLER_57_2338 ();
 sg13g2_decap_4 FILLER_57_2345 ();
 sg13g2_decap_8 FILLER_57_2354 ();
 sg13g2_decap_8 FILLER_57_2361 ();
 sg13g2_decap_8 FILLER_57_2368 ();
 sg13g2_decap_8 FILLER_57_2375 ();
 sg13g2_decap_4 FILLER_57_2382 ();
 sg13g2_fill_2 FILLER_57_2386 ();
 sg13g2_fill_1 FILLER_57_2394 ();
 sg13g2_decap_4 FILLER_57_2413 ();
 sg13g2_decap_8 FILLER_57_2431 ();
 sg13g2_decap_8 FILLER_57_2438 ();
 sg13g2_decap_4 FILLER_57_2445 ();
 sg13g2_fill_1 FILLER_57_2462 ();
 sg13g2_decap_8 FILLER_57_2477 ();
 sg13g2_decap_4 FILLER_57_2484 ();
 sg13g2_fill_1 FILLER_57_2488 ();
 sg13g2_decap_8 FILLER_57_2495 ();
 sg13g2_decap_8 FILLER_57_2502 ();
 sg13g2_decap_4 FILLER_57_2509 ();
 sg13g2_decap_8 FILLER_57_2523 ();
 sg13g2_decap_8 FILLER_57_2530 ();
 sg13g2_decap_8 FILLER_57_2537 ();
 sg13g2_decap_8 FILLER_57_2544 ();
 sg13g2_decap_4 FILLER_57_2551 ();
 sg13g2_fill_1 FILLER_57_2555 ();
 sg13g2_decap_8 FILLER_57_2566 ();
 sg13g2_decap_4 FILLER_57_2573 ();
 sg13g2_fill_2 FILLER_57_2577 ();
 sg13g2_decap_8 FILLER_57_2589 ();
 sg13g2_fill_2 FILLER_57_2596 ();
 sg13g2_fill_1 FILLER_57_2598 ();
 sg13g2_fill_2 FILLER_57_2605 ();
 sg13g2_decap_8 FILLER_57_2613 ();
 sg13g2_fill_2 FILLER_57_2620 ();
 sg13g2_fill_1 FILLER_57_2622 ();
 sg13g2_decap_4 FILLER_57_2644 ();
 sg13g2_fill_2 FILLER_57_2648 ();
 sg13g2_decap_8 FILLER_57_2658 ();
 sg13g2_decap_8 FILLER_57_2665 ();
 sg13g2_fill_1 FILLER_57_2672 ();
 sg13g2_decap_8 FILLER_57_2683 ();
 sg13g2_decap_8 FILLER_57_2690 ();
 sg13g2_fill_1 FILLER_57_2697 ();
 sg13g2_decap_8 FILLER_57_2724 ();
 sg13g2_fill_2 FILLER_57_2731 ();
 sg13g2_fill_1 FILLER_57_2733 ();
 sg13g2_decap_8 FILLER_57_2766 ();
 sg13g2_decap_8 FILLER_57_2773 ();
 sg13g2_decap_8 FILLER_57_2780 ();
 sg13g2_fill_2 FILLER_57_2787 ();
 sg13g2_fill_1 FILLER_57_2789 ();
 sg13g2_decap_8 FILLER_57_2798 ();
 sg13g2_decap_8 FILLER_57_2805 ();
 sg13g2_decap_8 FILLER_57_2812 ();
 sg13g2_fill_2 FILLER_57_2819 ();
 sg13g2_decap_8 FILLER_57_2847 ();
 sg13g2_decap_8 FILLER_57_2854 ();
 sg13g2_decap_8 FILLER_57_2861 ();
 sg13g2_decap_8 FILLER_57_2868 ();
 sg13g2_decap_8 FILLER_57_2875 ();
 sg13g2_decap_8 FILLER_57_2882 ();
 sg13g2_decap_8 FILLER_57_2899 ();
 sg13g2_decap_8 FILLER_57_2906 ();
 sg13g2_decap_8 FILLER_57_2913 ();
 sg13g2_decap_8 FILLER_57_2920 ();
 sg13g2_decap_8 FILLER_57_2927 ();
 sg13g2_decap_4 FILLER_57_2934 ();
 sg13g2_fill_1 FILLER_57_2938 ();
 sg13g2_fill_1 FILLER_57_2949 ();
 sg13g2_decap_8 FILLER_57_2960 ();
 sg13g2_decap_8 FILLER_57_2967 ();
 sg13g2_decap_8 FILLER_57_2974 ();
 sg13g2_decap_8 FILLER_57_2981 ();
 sg13g2_decap_8 FILLER_57_3014 ();
 sg13g2_decap_8 FILLER_57_3021 ();
 sg13g2_decap_8 FILLER_57_3028 ();
 sg13g2_decap_8 FILLER_57_3035 ();
 sg13g2_decap_4 FILLER_57_3042 ();
 sg13g2_decap_8 FILLER_57_3072 ();
 sg13g2_decap_8 FILLER_57_3079 ();
 sg13g2_decap_8 FILLER_57_3086 ();
 sg13g2_decap_4 FILLER_57_3093 ();
 sg13g2_decap_8 FILLER_57_3132 ();
 sg13g2_fill_2 FILLER_57_3139 ();
 sg13g2_fill_1 FILLER_57_3141 ();
 sg13g2_decap_8 FILLER_57_3160 ();
 sg13g2_decap_4 FILLER_57_3167 ();
 sg13g2_fill_1 FILLER_57_3171 ();
 sg13g2_fill_2 FILLER_57_3200 ();
 sg13g2_fill_2 FILLER_57_3208 ();
 sg13g2_decap_8 FILLER_57_3236 ();
 sg13g2_decap_8 FILLER_57_3243 ();
 sg13g2_fill_2 FILLER_57_3250 ();
 sg13g2_fill_1 FILLER_57_3252 ();
 sg13g2_decap_8 FILLER_57_3289 ();
 sg13g2_decap_8 FILLER_57_3296 ();
 sg13g2_decap_8 FILLER_57_3303 ();
 sg13g2_fill_2 FILLER_57_3310 ();
 sg13g2_fill_2 FILLER_57_3322 ();
 sg13g2_decap_8 FILLER_57_3350 ();
 sg13g2_decap_8 FILLER_57_3357 ();
 sg13g2_decap_4 FILLER_57_3364 ();
 sg13g2_fill_2 FILLER_57_3368 ();
 sg13g2_decap_8 FILLER_57_3402 ();
 sg13g2_decap_8 FILLER_57_3409 ();
 sg13g2_decap_8 FILLER_57_3416 ();
 sg13g2_decap_8 FILLER_57_3423 ();
 sg13g2_fill_2 FILLER_57_3430 ();
 sg13g2_fill_1 FILLER_57_3432 ();
 sg13g2_decap_8 FILLER_57_3437 ();
 sg13g2_decap_8 FILLER_57_3444 ();
 sg13g2_decap_8 FILLER_57_3451 ();
 sg13g2_decap_8 FILLER_57_3458 ();
 sg13g2_decap_8 FILLER_57_3465 ();
 sg13g2_fill_2 FILLER_57_3472 ();
 sg13g2_decap_4 FILLER_57_3504 ();
 sg13g2_fill_1 FILLER_57_3508 ();
 sg13g2_decap_8 FILLER_57_3514 ();
 sg13g2_decap_8 FILLER_57_3521 ();
 sg13g2_decap_8 FILLER_57_3557 ();
 sg13g2_decap_8 FILLER_57_3564 ();
 sg13g2_decap_8 FILLER_57_3571 ();
 sg13g2_fill_2 FILLER_57_3578 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_fill_2 FILLER_58_7 ();
 sg13g2_fill_2 FILLER_58_40 ();
 sg13g2_decap_8 FILLER_58_68 ();
 sg13g2_decap_8 FILLER_58_75 ();
 sg13g2_decap_8 FILLER_58_82 ();
 sg13g2_decap_8 FILLER_58_115 ();
 sg13g2_decap_8 FILLER_58_122 ();
 sg13g2_decap_8 FILLER_58_129 ();
 sg13g2_decap_4 FILLER_58_136 ();
 sg13g2_fill_2 FILLER_58_140 ();
 sg13g2_decap_8 FILLER_58_173 ();
 sg13g2_fill_2 FILLER_58_195 ();
 sg13g2_decap_8 FILLER_58_202 ();
 sg13g2_decap_8 FILLER_58_209 ();
 sg13g2_decap_8 FILLER_58_216 ();
 sg13g2_decap_8 FILLER_58_223 ();
 sg13g2_decap_8 FILLER_58_230 ();
 sg13g2_decap_4 FILLER_58_237 ();
 sg13g2_decap_8 FILLER_58_271 ();
 sg13g2_decap_8 FILLER_58_278 ();
 sg13g2_decap_8 FILLER_58_285 ();
 sg13g2_decap_8 FILLER_58_292 ();
 sg13g2_decap_8 FILLER_58_299 ();
 sg13g2_decap_8 FILLER_58_306 ();
 sg13g2_decap_8 FILLER_58_322 ();
 sg13g2_fill_1 FILLER_58_338 ();
 sg13g2_decap_4 FILLER_58_344 ();
 sg13g2_fill_1 FILLER_58_348 ();
 sg13g2_decap_8 FILLER_58_354 ();
 sg13g2_decap_4 FILLER_58_361 ();
 sg13g2_decap_8 FILLER_58_370 ();
 sg13g2_decap_4 FILLER_58_377 ();
 sg13g2_fill_1 FILLER_58_381 ();
 sg13g2_fill_1 FILLER_58_387 ();
 sg13g2_decap_8 FILLER_58_415 ();
 sg13g2_decap_8 FILLER_58_422 ();
 sg13g2_decap_8 FILLER_58_429 ();
 sg13g2_decap_8 FILLER_58_436 ();
 sg13g2_decap_8 FILLER_58_443 ();
 sg13g2_decap_8 FILLER_58_450 ();
 sg13g2_decap_8 FILLER_58_457 ();
 sg13g2_decap_8 FILLER_58_464 ();
 sg13g2_decap_8 FILLER_58_471 ();
 sg13g2_decap_4 FILLER_58_478 ();
 sg13g2_fill_2 FILLER_58_482 ();
 sg13g2_decap_8 FILLER_58_490 ();
 sg13g2_decap_8 FILLER_58_497 ();
 sg13g2_decap_8 FILLER_58_504 ();
 sg13g2_fill_1 FILLER_58_511 ();
 sg13g2_decap_8 FILLER_58_525 ();
 sg13g2_decap_8 FILLER_58_532 ();
 sg13g2_decap_8 FILLER_58_539 ();
 sg13g2_decap_8 FILLER_58_546 ();
 sg13g2_fill_2 FILLER_58_553 ();
 sg13g2_decap_8 FILLER_58_577 ();
 sg13g2_decap_8 FILLER_58_584 ();
 sg13g2_decap_8 FILLER_58_591 ();
 sg13g2_decap_8 FILLER_58_598 ();
 sg13g2_decap_8 FILLER_58_605 ();
 sg13g2_decap_8 FILLER_58_612 ();
 sg13g2_decap_8 FILLER_58_619 ();
 sg13g2_decap_8 FILLER_58_639 ();
 sg13g2_decap_8 FILLER_58_646 ();
 sg13g2_decap_8 FILLER_58_653 ();
 sg13g2_decap_8 FILLER_58_660 ();
 sg13g2_fill_1 FILLER_58_667 ();
 sg13g2_fill_1 FILLER_58_679 ();
 sg13g2_decap_4 FILLER_58_696 ();
 sg13g2_decap_8 FILLER_58_706 ();
 sg13g2_decap_8 FILLER_58_713 ();
 sg13g2_decap_4 FILLER_58_720 ();
 sg13g2_fill_1 FILLER_58_724 ();
 sg13g2_fill_2 FILLER_58_738 ();
 sg13g2_fill_1 FILLER_58_740 ();
 sg13g2_decap_4 FILLER_58_744 ();
 sg13g2_fill_1 FILLER_58_748 ();
 sg13g2_decap_8 FILLER_58_775 ();
 sg13g2_decap_8 FILLER_58_782 ();
 sg13g2_decap_8 FILLER_58_789 ();
 sg13g2_fill_2 FILLER_58_796 ();
 sg13g2_fill_1 FILLER_58_798 ();
 sg13g2_fill_2 FILLER_58_812 ();
 sg13g2_decap_4 FILLER_58_818 ();
 sg13g2_decap_8 FILLER_58_831 ();
 sg13g2_fill_1 FILLER_58_838 ();
 sg13g2_decap_4 FILLER_58_847 ();
 sg13g2_fill_1 FILLER_58_851 ();
 sg13g2_decap_8 FILLER_58_856 ();
 sg13g2_fill_1 FILLER_58_863 ();
 sg13g2_fill_1 FILLER_58_872 ();
 sg13g2_decap_8 FILLER_58_878 ();
 sg13g2_decap_4 FILLER_58_885 ();
 sg13g2_fill_2 FILLER_58_889 ();
 sg13g2_decap_4 FILLER_58_899 ();
 sg13g2_decap_8 FILLER_58_924 ();
 sg13g2_decap_8 FILLER_58_931 ();
 sg13g2_decap_8 FILLER_58_938 ();
 sg13g2_fill_1 FILLER_58_945 ();
 sg13g2_decap_8 FILLER_58_970 ();
 sg13g2_decap_8 FILLER_58_977 ();
 sg13g2_decap_8 FILLER_58_984 ();
 sg13g2_decap_4 FILLER_58_991 ();
 sg13g2_fill_1 FILLER_58_995 ();
 sg13g2_fill_1 FILLER_58_1007 ();
 sg13g2_fill_2 FILLER_58_1029 ();
 sg13g2_fill_1 FILLER_58_1039 ();
 sg13g2_fill_2 FILLER_58_1063 ();
 sg13g2_decap_4 FILLER_58_1073 ();
 sg13g2_fill_2 FILLER_58_1077 ();
 sg13g2_fill_1 FILLER_58_1083 ();
 sg13g2_decap_8 FILLER_58_1107 ();
 sg13g2_decap_8 FILLER_58_1114 ();
 sg13g2_decap_8 FILLER_58_1121 ();
 sg13g2_decap_8 FILLER_58_1128 ();
 sg13g2_decap_8 FILLER_58_1135 ();
 sg13g2_decap_8 FILLER_58_1142 ();
 sg13g2_decap_8 FILLER_58_1149 ();
 sg13g2_decap_8 FILLER_58_1156 ();
 sg13g2_decap_8 FILLER_58_1163 ();
 sg13g2_decap_8 FILLER_58_1170 ();
 sg13g2_decap_8 FILLER_58_1177 ();
 sg13g2_decap_8 FILLER_58_1184 ();
 sg13g2_fill_2 FILLER_58_1196 ();
 sg13g2_fill_1 FILLER_58_1198 ();
 sg13g2_decap_8 FILLER_58_1209 ();
 sg13g2_fill_1 FILLER_58_1216 ();
 sg13g2_decap_8 FILLER_58_1226 ();
 sg13g2_decap_8 FILLER_58_1233 ();
 sg13g2_decap_8 FILLER_58_1240 ();
 sg13g2_decap_8 FILLER_58_1247 ();
 sg13g2_fill_1 FILLER_58_1254 ();
 sg13g2_decap_8 FILLER_58_1265 ();
 sg13g2_decap_8 FILLER_58_1272 ();
 sg13g2_decap_8 FILLER_58_1279 ();
 sg13g2_decap_4 FILLER_58_1286 ();
 sg13g2_fill_2 FILLER_58_1326 ();
 sg13g2_decap_8 FILLER_58_1338 ();
 sg13g2_decap_8 FILLER_58_1345 ();
 sg13g2_decap_8 FILLER_58_1352 ();
 sg13g2_decap_8 FILLER_58_1359 ();
 sg13g2_decap_8 FILLER_58_1366 ();
 sg13g2_decap_8 FILLER_58_1373 ();
 sg13g2_decap_8 FILLER_58_1388 ();
 sg13g2_decap_8 FILLER_58_1395 ();
 sg13g2_decap_8 FILLER_58_1402 ();
 sg13g2_fill_2 FILLER_58_1409 ();
 sg13g2_decap_8 FILLER_58_1445 ();
 sg13g2_decap_8 FILLER_58_1452 ();
 sg13g2_decap_8 FILLER_58_1459 ();
 sg13g2_decap_8 FILLER_58_1466 ();
 sg13g2_decap_8 FILLER_58_1491 ();
 sg13g2_decap_8 FILLER_58_1498 ();
 sg13g2_decap_8 FILLER_58_1505 ();
 sg13g2_decap_8 FILLER_58_1512 ();
 sg13g2_decap_8 FILLER_58_1519 ();
 sg13g2_decap_8 FILLER_58_1526 ();
 sg13g2_fill_2 FILLER_58_1533 ();
 sg13g2_decap_8 FILLER_58_1545 ();
 sg13g2_decap_8 FILLER_58_1552 ();
 sg13g2_decap_8 FILLER_58_1559 ();
 sg13g2_decap_8 FILLER_58_1566 ();
 sg13g2_decap_8 FILLER_58_1573 ();
 sg13g2_decap_8 FILLER_58_1580 ();
 sg13g2_decap_4 FILLER_58_1587 ();
 sg13g2_decap_8 FILLER_58_1600 ();
 sg13g2_decap_8 FILLER_58_1607 ();
 sg13g2_decap_8 FILLER_58_1614 ();
 sg13g2_decap_4 FILLER_58_1621 ();
 sg13g2_fill_2 FILLER_58_1635 ();
 sg13g2_decap_8 FILLER_58_1663 ();
 sg13g2_decap_8 FILLER_58_1670 ();
 sg13g2_decap_4 FILLER_58_1677 ();
 sg13g2_fill_2 FILLER_58_1681 ();
 sg13g2_fill_2 FILLER_58_1688 ();
 sg13g2_fill_1 FILLER_58_1690 ();
 sg13g2_decap_8 FILLER_58_1696 ();
 sg13g2_decap_8 FILLER_58_1703 ();
 sg13g2_decap_8 FILLER_58_1710 ();
 sg13g2_decap_8 FILLER_58_1717 ();
 sg13g2_decap_8 FILLER_58_1724 ();
 sg13g2_decap_8 FILLER_58_1731 ();
 sg13g2_decap_8 FILLER_58_1738 ();
 sg13g2_decap_8 FILLER_58_1745 ();
 sg13g2_decap_8 FILLER_58_1752 ();
 sg13g2_decap_8 FILLER_58_1789 ();
 sg13g2_decap_4 FILLER_58_1796 ();
 sg13g2_fill_1 FILLER_58_1800 ();
 sg13g2_decap_8 FILLER_58_1807 ();
 sg13g2_decap_8 FILLER_58_1814 ();
 sg13g2_decap_8 FILLER_58_1821 ();
 sg13g2_decap_4 FILLER_58_1828 ();
 sg13g2_fill_2 FILLER_58_1832 ();
 sg13g2_fill_2 FILLER_58_1844 ();
 sg13g2_decap_4 FILLER_58_1856 ();
 sg13g2_fill_2 FILLER_58_1860 ();
 sg13g2_decap_8 FILLER_58_1888 ();
 sg13g2_decap_8 FILLER_58_1895 ();
 sg13g2_decap_8 FILLER_58_1902 ();
 sg13g2_decap_8 FILLER_58_1909 ();
 sg13g2_decap_8 FILLER_58_1925 ();
 sg13g2_decap_8 FILLER_58_1932 ();
 sg13g2_decap_8 FILLER_58_1939 ();
 sg13g2_decap_8 FILLER_58_1946 ();
 sg13g2_decap_8 FILLER_58_1953 ();
 sg13g2_decap_8 FILLER_58_1960 ();
 sg13g2_fill_1 FILLER_58_1967 ();
 sg13g2_decap_8 FILLER_58_1978 ();
 sg13g2_decap_8 FILLER_58_1985 ();
 sg13g2_decap_8 FILLER_58_1992 ();
 sg13g2_decap_8 FILLER_58_1999 ();
 sg13g2_decap_8 FILLER_58_2006 ();
 sg13g2_decap_8 FILLER_58_2047 ();
 sg13g2_decap_8 FILLER_58_2054 ();
 sg13g2_fill_2 FILLER_58_2061 ();
 sg13g2_fill_1 FILLER_58_2067 ();
 sg13g2_decap_8 FILLER_58_2108 ();
 sg13g2_fill_1 FILLER_58_2121 ();
 sg13g2_fill_2 FILLER_58_2135 ();
 sg13g2_fill_1 FILLER_58_2137 ();
 sg13g2_decap_8 FILLER_58_2164 ();
 sg13g2_decap_8 FILLER_58_2171 ();
 sg13g2_fill_2 FILLER_58_2178 ();
 sg13g2_decap_8 FILLER_58_2189 ();
 sg13g2_fill_2 FILLER_58_2196 ();
 sg13g2_decap_8 FILLER_58_2204 ();
 sg13g2_decap_8 FILLER_58_2211 ();
 sg13g2_decap_8 FILLER_58_2218 ();
 sg13g2_decap_8 FILLER_58_2225 ();
 sg13g2_decap_8 FILLER_58_2232 ();
 sg13g2_decap_8 FILLER_58_2239 ();
 sg13g2_decap_8 FILLER_58_2246 ();
 sg13g2_decap_8 FILLER_58_2253 ();
 sg13g2_decap_8 FILLER_58_2260 ();
 sg13g2_decap_8 FILLER_58_2267 ();
 sg13g2_decap_8 FILLER_58_2274 ();
 sg13g2_fill_2 FILLER_58_2281 ();
 sg13g2_decap_8 FILLER_58_2298 ();
 sg13g2_decap_8 FILLER_58_2305 ();
 sg13g2_decap_8 FILLER_58_2312 ();
 sg13g2_fill_1 FILLER_58_2319 ();
 sg13g2_decap_8 FILLER_58_2326 ();
 sg13g2_fill_1 FILLER_58_2333 ();
 sg13g2_decap_8 FILLER_58_2349 ();
 sg13g2_decap_8 FILLER_58_2356 ();
 sg13g2_decap_8 FILLER_58_2363 ();
 sg13g2_decap_8 FILLER_58_2370 ();
 sg13g2_decap_4 FILLER_58_2377 ();
 sg13g2_fill_1 FILLER_58_2381 ();
 sg13g2_fill_2 FILLER_58_2411 ();
 sg13g2_decap_8 FILLER_58_2441 ();
 sg13g2_decap_4 FILLER_58_2448 ();
 sg13g2_fill_1 FILLER_58_2452 ();
 sg13g2_decap_4 FILLER_58_2474 ();
 sg13g2_fill_2 FILLER_58_2478 ();
 sg13g2_decap_8 FILLER_58_2490 ();
 sg13g2_decap_8 FILLER_58_2497 ();
 sg13g2_decap_8 FILLER_58_2504 ();
 sg13g2_decap_8 FILLER_58_2511 ();
 sg13g2_decap_8 FILLER_58_2518 ();
 sg13g2_decap_8 FILLER_58_2525 ();
 sg13g2_decap_8 FILLER_58_2532 ();
 sg13g2_decap_8 FILLER_58_2539 ();
 sg13g2_decap_8 FILLER_58_2546 ();
 sg13g2_fill_2 FILLER_58_2553 ();
 sg13g2_decap_4 FILLER_58_2581 ();
 sg13g2_fill_2 FILLER_58_2585 ();
 sg13g2_decap_8 FILLER_58_2621 ();
 sg13g2_decap_8 FILLER_58_2628 ();
 sg13g2_decap_8 FILLER_58_2635 ();
 sg13g2_fill_1 FILLER_58_2642 ();
 sg13g2_decap_8 FILLER_58_2669 ();
 sg13g2_decap_8 FILLER_58_2676 ();
 sg13g2_decap_8 FILLER_58_2683 ();
 sg13g2_decap_8 FILLER_58_2690 ();
 sg13g2_decap_4 FILLER_58_2697 ();
 sg13g2_decap_8 FILLER_58_2727 ();
 sg13g2_decap_8 FILLER_58_2734 ();
 sg13g2_decap_8 FILLER_58_2741 ();
 sg13g2_decap_8 FILLER_58_2748 ();
 sg13g2_decap_8 FILLER_58_2760 ();
 sg13g2_decap_8 FILLER_58_2767 ();
 sg13g2_decap_8 FILLER_58_2774 ();
 sg13g2_decap_8 FILLER_58_2781 ();
 sg13g2_decap_8 FILLER_58_2799 ();
 sg13g2_decap_8 FILLER_58_2806 ();
 sg13g2_decap_8 FILLER_58_2813 ();
 sg13g2_fill_1 FILLER_58_2820 ();
 sg13g2_fill_2 FILLER_58_2831 ();
 sg13g2_fill_1 FILLER_58_2833 ();
 sg13g2_decap_8 FILLER_58_2854 ();
 sg13g2_decap_8 FILLER_58_2861 ();
 sg13g2_decap_8 FILLER_58_2868 ();
 sg13g2_decap_8 FILLER_58_2875 ();
 sg13g2_decap_4 FILLER_58_2882 ();
 sg13g2_fill_2 FILLER_58_2886 ();
 sg13g2_decap_8 FILLER_58_2914 ();
 sg13g2_fill_2 FILLER_58_2921 ();
 sg13g2_fill_1 FILLER_58_2923 ();
 sg13g2_decap_8 FILLER_58_2950 ();
 sg13g2_decap_8 FILLER_58_2957 ();
 sg13g2_fill_2 FILLER_58_2964 ();
 sg13g2_fill_1 FILLER_58_2966 ();
 sg13g2_decap_4 FILLER_58_2986 ();
 sg13g2_fill_2 FILLER_58_2990 ();
 sg13g2_decap_8 FILLER_58_3002 ();
 sg13g2_decap_8 FILLER_58_3009 ();
 sg13g2_decap_8 FILLER_58_3016 ();
 sg13g2_fill_1 FILLER_58_3023 ();
 sg13g2_fill_2 FILLER_58_3055 ();
 sg13g2_fill_1 FILLER_58_3062 ();
 sg13g2_decap_8 FILLER_58_3073 ();
 sg13g2_decap_8 FILLER_58_3080 ();
 sg13g2_decap_8 FILLER_58_3087 ();
 sg13g2_decap_8 FILLER_58_3094 ();
 sg13g2_decap_8 FILLER_58_3101 ();
 sg13g2_decap_8 FILLER_58_3108 ();
 sg13g2_decap_8 FILLER_58_3115 ();
 sg13g2_decap_8 FILLER_58_3122 ();
 sg13g2_decap_8 FILLER_58_3129 ();
 sg13g2_decap_4 FILLER_58_3136 ();
 sg13g2_fill_1 FILLER_58_3140 ();
 sg13g2_decap_8 FILLER_58_3167 ();
 sg13g2_decap_4 FILLER_58_3174 ();
 sg13g2_decap_4 FILLER_58_3209 ();
 sg13g2_decap_8 FILLER_58_3239 ();
 sg13g2_decap_8 FILLER_58_3246 ();
 sg13g2_decap_8 FILLER_58_3253 ();
 sg13g2_decap_8 FILLER_58_3260 ();
 sg13g2_decap_8 FILLER_58_3267 ();
 sg13g2_decap_4 FILLER_58_3274 ();
 sg13g2_decap_8 FILLER_58_3288 ();
 sg13g2_decap_8 FILLER_58_3295 ();
 sg13g2_decap_8 FILLER_58_3302 ();
 sg13g2_decap_4 FILLER_58_3309 ();
 sg13g2_decap_4 FILLER_58_3349 ();
 sg13g2_decap_8 FILLER_58_3361 ();
 sg13g2_decap_4 FILLER_58_3368 ();
 sg13g2_fill_2 FILLER_58_3372 ();
 sg13g2_decap_8 FILLER_58_3394 ();
 sg13g2_decap_8 FILLER_58_3401 ();
 sg13g2_decap_8 FILLER_58_3408 ();
 sg13g2_decap_8 FILLER_58_3415 ();
 sg13g2_decap_8 FILLER_58_3422 ();
 sg13g2_fill_1 FILLER_58_3429 ();
 sg13g2_decap_8 FILLER_58_3443 ();
 sg13g2_decap_8 FILLER_58_3450 ();
 sg13g2_decap_8 FILLER_58_3457 ();
 sg13g2_decap_8 FILLER_58_3464 ();
 sg13g2_fill_1 FILLER_58_3471 ();
 sg13g2_decap_8 FILLER_58_3477 ();
 sg13g2_decap_8 FILLER_58_3484 ();
 sg13g2_decap_8 FILLER_58_3491 ();
 sg13g2_decap_8 FILLER_58_3498 ();
 sg13g2_decap_8 FILLER_58_3505 ();
 sg13g2_decap_8 FILLER_58_3512 ();
 sg13g2_decap_8 FILLER_58_3519 ();
 sg13g2_decap_8 FILLER_58_3526 ();
 sg13g2_decap_8 FILLER_58_3533 ();
 sg13g2_decap_4 FILLER_58_3540 ();
 sg13g2_fill_2 FILLER_58_3544 ();
 sg13g2_decap_8 FILLER_58_3572 ();
 sg13g2_fill_1 FILLER_58_3579 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_fill_2 FILLER_59_7 ();
 sg13g2_decap_8 FILLER_59_71 ();
 sg13g2_decap_8 FILLER_59_78 ();
 sg13g2_decap_8 FILLER_59_85 ();
 sg13g2_fill_2 FILLER_59_92 ();
 sg13g2_fill_1 FILLER_59_99 ();
 sg13g2_decap_4 FILLER_59_104 ();
 sg13g2_decap_8 FILLER_59_117 ();
 sg13g2_decap_8 FILLER_59_124 ();
 sg13g2_decap_8 FILLER_59_131 ();
 sg13g2_fill_1 FILLER_59_151 ();
 sg13g2_decap_8 FILLER_59_170 ();
 sg13g2_decap_8 FILLER_59_177 ();
 sg13g2_decap_8 FILLER_59_184 ();
 sg13g2_decap_4 FILLER_59_191 ();
 sg13g2_fill_2 FILLER_59_195 ();
 sg13g2_decap_8 FILLER_59_205 ();
 sg13g2_decap_8 FILLER_59_212 ();
 sg13g2_decap_4 FILLER_59_219 ();
 sg13g2_fill_2 FILLER_59_223 ();
 sg13g2_fill_2 FILLER_59_234 ();
 sg13g2_fill_1 FILLER_59_236 ();
 sg13g2_decap_4 FILLER_59_245 ();
 sg13g2_fill_2 FILLER_59_249 ();
 sg13g2_decap_8 FILLER_59_259 ();
 sg13g2_decap_8 FILLER_59_266 ();
 sg13g2_decap_8 FILLER_59_273 ();
 sg13g2_decap_8 FILLER_59_280 ();
 sg13g2_decap_8 FILLER_59_287 ();
 sg13g2_decap_8 FILLER_59_294 ();
 sg13g2_decap_4 FILLER_59_301 ();
 sg13g2_fill_1 FILLER_59_355 ();
 sg13g2_decap_4 FILLER_59_376 ();
 sg13g2_fill_2 FILLER_59_380 ();
 sg13g2_fill_2 FILLER_59_406 ();
 sg13g2_decap_8 FILLER_59_434 ();
 sg13g2_fill_2 FILLER_59_441 ();
 sg13g2_fill_1 FILLER_59_443 ();
 sg13g2_fill_1 FILLER_59_457 ();
 sg13g2_fill_1 FILLER_59_484 ();
 sg13g2_decap_8 FILLER_59_497 ();
 sg13g2_fill_1 FILLER_59_504 ();
 sg13g2_decap_8 FILLER_59_524 ();
 sg13g2_decap_8 FILLER_59_531 ();
 sg13g2_decap_8 FILLER_59_538 ();
 sg13g2_fill_1 FILLER_59_545 ();
 sg13g2_fill_1 FILLER_59_560 ();
 sg13g2_decap_8 FILLER_59_578 ();
 sg13g2_decap_8 FILLER_59_585 ();
 sg13g2_decap_8 FILLER_59_592 ();
 sg13g2_decap_8 FILLER_59_599 ();
 sg13g2_decap_8 FILLER_59_606 ();
 sg13g2_decap_8 FILLER_59_613 ();
 sg13g2_fill_2 FILLER_59_620 ();
 sg13g2_fill_1 FILLER_59_635 ();
 sg13g2_decap_8 FILLER_59_644 ();
 sg13g2_decap_8 FILLER_59_651 ();
 sg13g2_decap_8 FILLER_59_658 ();
 sg13g2_decap_8 FILLER_59_665 ();
 sg13g2_decap_8 FILLER_59_672 ();
 sg13g2_decap_8 FILLER_59_679 ();
 sg13g2_decap_8 FILLER_59_686 ();
 sg13g2_decap_8 FILLER_59_693 ();
 sg13g2_decap_4 FILLER_59_700 ();
 sg13g2_fill_1 FILLER_59_704 ();
 sg13g2_decap_8 FILLER_59_711 ();
 sg13g2_fill_1 FILLER_59_718 ();
 sg13g2_decap_8 FILLER_59_755 ();
 sg13g2_decap_8 FILLER_59_762 ();
 sg13g2_decap_8 FILLER_59_769 ();
 sg13g2_decap_8 FILLER_59_776 ();
 sg13g2_decap_8 FILLER_59_783 ();
 sg13g2_fill_2 FILLER_59_790 ();
 sg13g2_fill_1 FILLER_59_797 ();
 sg13g2_fill_1 FILLER_59_814 ();
 sg13g2_decap_8 FILLER_59_849 ();
 sg13g2_decap_4 FILLER_59_856 ();
 sg13g2_fill_2 FILLER_59_865 ();
 sg13g2_fill_1 FILLER_59_867 ();
 sg13g2_decap_8 FILLER_59_883 ();
 sg13g2_fill_1 FILLER_59_890 ();
 sg13g2_fill_2 FILLER_59_913 ();
 sg13g2_decap_8 FILLER_59_922 ();
 sg13g2_decap_8 FILLER_59_929 ();
 sg13g2_decap_8 FILLER_59_936 ();
 sg13g2_decap_8 FILLER_59_943 ();
 sg13g2_decap_4 FILLER_59_950 ();
 sg13g2_fill_2 FILLER_59_954 ();
 sg13g2_decap_8 FILLER_59_961 ();
 sg13g2_decap_8 FILLER_59_968 ();
 sg13g2_decap_8 FILLER_59_975 ();
 sg13g2_decap_8 FILLER_59_982 ();
 sg13g2_decap_8 FILLER_59_989 ();
 sg13g2_decap_8 FILLER_59_996 ();
 sg13g2_decap_8 FILLER_59_1003 ();
 sg13g2_decap_4 FILLER_59_1010 ();
 sg13g2_fill_2 FILLER_59_1014 ();
 sg13g2_decap_8 FILLER_59_1024 ();
 sg13g2_decap_4 FILLER_59_1031 ();
 sg13g2_fill_2 FILLER_59_1043 ();
 sg13g2_decap_8 FILLER_59_1050 ();
 sg13g2_decap_8 FILLER_59_1057 ();
 sg13g2_decap_8 FILLER_59_1064 ();
 sg13g2_decap_4 FILLER_59_1071 ();
 sg13g2_fill_2 FILLER_59_1075 ();
 sg13g2_decap_4 FILLER_59_1082 ();
 sg13g2_fill_1 FILLER_59_1086 ();
 sg13g2_decap_4 FILLER_59_1092 ();
 sg13g2_decap_8 FILLER_59_1104 ();
 sg13g2_decap_8 FILLER_59_1111 ();
 sg13g2_decap_8 FILLER_59_1118 ();
 sg13g2_decap_8 FILLER_59_1125 ();
 sg13g2_decap_8 FILLER_59_1132 ();
 sg13g2_fill_2 FILLER_59_1139 ();
 sg13g2_fill_1 FILLER_59_1141 ();
 sg13g2_decap_8 FILLER_59_1154 ();
 sg13g2_decap_8 FILLER_59_1161 ();
 sg13g2_decap_8 FILLER_59_1168 ();
 sg13g2_decap_4 FILLER_59_1175 ();
 sg13g2_fill_1 FILLER_59_1179 ();
 sg13g2_decap_8 FILLER_59_1232 ();
 sg13g2_decap_8 FILLER_59_1239 ();
 sg13g2_decap_8 FILLER_59_1246 ();
 sg13g2_decap_8 FILLER_59_1253 ();
 sg13g2_decap_8 FILLER_59_1260 ();
 sg13g2_decap_8 FILLER_59_1267 ();
 sg13g2_decap_8 FILLER_59_1274 ();
 sg13g2_decap_8 FILLER_59_1281 ();
 sg13g2_decap_8 FILLER_59_1288 ();
 sg13g2_decap_8 FILLER_59_1295 ();
 sg13g2_decap_8 FILLER_59_1302 ();
 sg13g2_decap_8 FILLER_59_1309 ();
 sg13g2_decap_8 FILLER_59_1316 ();
 sg13g2_decap_8 FILLER_59_1323 ();
 sg13g2_decap_8 FILLER_59_1330 ();
 sg13g2_fill_1 FILLER_59_1337 ();
 sg13g2_decap_8 FILLER_59_1364 ();
 sg13g2_decap_8 FILLER_59_1371 ();
 sg13g2_decap_4 FILLER_59_1378 ();
 sg13g2_decap_8 FILLER_59_1387 ();
 sg13g2_decap_8 FILLER_59_1394 ();
 sg13g2_decap_8 FILLER_59_1401 ();
 sg13g2_decap_8 FILLER_59_1408 ();
 sg13g2_decap_8 FILLER_59_1415 ();
 sg13g2_decap_4 FILLER_59_1422 ();
 sg13g2_fill_1 FILLER_59_1426 ();
 sg13g2_decap_8 FILLER_59_1435 ();
 sg13g2_fill_2 FILLER_59_1442 ();
 sg13g2_decap_8 FILLER_59_1454 ();
 sg13g2_decap_8 FILLER_59_1461 ();
 sg13g2_decap_8 FILLER_59_1468 ();
 sg13g2_decap_4 FILLER_59_1475 ();
 sg13g2_decap_8 FILLER_59_1487 ();
 sg13g2_decap_8 FILLER_59_1494 ();
 sg13g2_decap_8 FILLER_59_1501 ();
 sg13g2_fill_1 FILLER_59_1534 ();
 sg13g2_decap_8 FILLER_59_1561 ();
 sg13g2_decap_8 FILLER_59_1568 ();
 sg13g2_decap_8 FILLER_59_1575 ();
 sg13g2_decap_8 FILLER_59_1582 ();
 sg13g2_decap_8 FILLER_59_1601 ();
 sg13g2_decap_4 FILLER_59_1608 ();
 sg13g2_fill_1 FILLER_59_1612 ();
 sg13g2_decap_8 FILLER_59_1628 ();
 sg13g2_decap_8 FILLER_59_1635 ();
 sg13g2_decap_8 FILLER_59_1642 ();
 sg13g2_decap_8 FILLER_59_1649 ();
 sg13g2_decap_8 FILLER_59_1656 ();
 sg13g2_decap_8 FILLER_59_1663 ();
 sg13g2_decap_4 FILLER_59_1670 ();
 sg13g2_fill_1 FILLER_59_1690 ();
 sg13g2_decap_8 FILLER_59_1703 ();
 sg13g2_decap_8 FILLER_59_1710 ();
 sg13g2_decap_8 FILLER_59_1717 ();
 sg13g2_decap_4 FILLER_59_1724 ();
 sg13g2_fill_2 FILLER_59_1728 ();
 sg13g2_decap_8 FILLER_59_1744 ();
 sg13g2_decap_8 FILLER_59_1751 ();
 sg13g2_fill_2 FILLER_59_1758 ();
 sg13g2_decap_8 FILLER_59_1792 ();
 sg13g2_decap_8 FILLER_59_1799 ();
 sg13g2_decap_8 FILLER_59_1806 ();
 sg13g2_decap_8 FILLER_59_1813 ();
 sg13g2_fill_2 FILLER_59_1820 ();
 sg13g2_fill_1 FILLER_59_1822 ();
 sg13g2_fill_2 FILLER_59_1849 ();
 sg13g2_decap_8 FILLER_59_1877 ();
 sg13g2_decap_8 FILLER_59_1884 ();
 sg13g2_decap_8 FILLER_59_1891 ();
 sg13g2_decap_8 FILLER_59_1898 ();
 sg13g2_decap_8 FILLER_59_1905 ();
 sg13g2_decap_8 FILLER_59_1912 ();
 sg13g2_fill_2 FILLER_59_1919 ();
 sg13g2_fill_1 FILLER_59_1927 ();
 sg13g2_decap_8 FILLER_59_1938 ();
 sg13g2_decap_8 FILLER_59_1945 ();
 sg13g2_decap_8 FILLER_59_1952 ();
 sg13g2_decap_8 FILLER_59_1959 ();
 sg13g2_fill_1 FILLER_59_1966 ();
 sg13g2_decap_8 FILLER_59_1977 ();
 sg13g2_decap_8 FILLER_59_1996 ();
 sg13g2_decap_8 FILLER_59_2003 ();
 sg13g2_decap_4 FILLER_59_2010 ();
 sg13g2_decap_8 FILLER_59_2029 ();
 sg13g2_decap_8 FILLER_59_2036 ();
 sg13g2_fill_2 FILLER_59_2043 ();
 sg13g2_decap_8 FILLER_59_2053 ();
 sg13g2_decap_4 FILLER_59_2086 ();
 sg13g2_fill_2 FILLER_59_2090 ();
 sg13g2_decap_8 FILLER_59_2098 ();
 sg13g2_decap_8 FILLER_59_2105 ();
 sg13g2_decap_8 FILLER_59_2112 ();
 sg13g2_fill_1 FILLER_59_2119 ();
 sg13g2_decap_8 FILLER_59_2159 ();
 sg13g2_decap_8 FILLER_59_2166 ();
 sg13g2_decap_4 FILLER_59_2173 ();
 sg13g2_fill_1 FILLER_59_2177 ();
 sg13g2_fill_1 FILLER_59_2184 ();
 sg13g2_decap_4 FILLER_59_2193 ();
 sg13g2_fill_2 FILLER_59_2197 ();
 sg13g2_decap_8 FILLER_59_2218 ();
 sg13g2_decap_4 FILLER_59_2225 ();
 sg13g2_fill_1 FILLER_59_2229 ();
 sg13g2_decap_8 FILLER_59_2236 ();
 sg13g2_decap_8 FILLER_59_2243 ();
 sg13g2_decap_8 FILLER_59_2250 ();
 sg13g2_fill_2 FILLER_59_2263 ();
 sg13g2_decap_4 FILLER_59_2268 ();
 sg13g2_fill_2 FILLER_59_2272 ();
 sg13g2_fill_2 FILLER_59_2304 ();
 sg13g2_fill_1 FILLER_59_2306 ();
 sg13g2_fill_1 FILLER_59_2340 ();
 sg13g2_decap_8 FILLER_59_2367 ();
 sg13g2_decap_8 FILLER_59_2374 ();
 sg13g2_decap_8 FILLER_59_2381 ();
 sg13g2_fill_2 FILLER_59_2388 ();
 sg13g2_fill_1 FILLER_59_2390 ();
 sg13g2_decap_8 FILLER_59_2431 ();
 sg13g2_decap_8 FILLER_59_2438 ();
 sg13g2_decap_8 FILLER_59_2445 ();
 sg13g2_decap_8 FILLER_59_2452 ();
 sg13g2_decap_8 FILLER_59_2459 ();
 sg13g2_decap_8 FILLER_59_2466 ();
 sg13g2_decap_8 FILLER_59_2509 ();
 sg13g2_decap_8 FILLER_59_2516 ();
 sg13g2_decap_8 FILLER_59_2523 ();
 sg13g2_decap_8 FILLER_59_2530 ();
 sg13g2_fill_2 FILLER_59_2537 ();
 sg13g2_fill_1 FILLER_59_2539 ();
 sg13g2_fill_1 FILLER_59_2545 ();
 sg13g2_decap_8 FILLER_59_2564 ();
 sg13g2_decap_8 FILLER_59_2571 ();
 sg13g2_decap_8 FILLER_59_2578 ();
 sg13g2_decap_8 FILLER_59_2585 ();
 sg13g2_decap_8 FILLER_59_2592 ();
 sg13g2_decap_8 FILLER_59_2599 ();
 sg13g2_decap_8 FILLER_59_2616 ();
 sg13g2_decap_8 FILLER_59_2623 ();
 sg13g2_decap_8 FILLER_59_2630 ();
 sg13g2_decap_8 FILLER_59_2637 ();
 sg13g2_decap_8 FILLER_59_2644 ();
 sg13g2_decap_8 FILLER_59_2655 ();
 sg13g2_decap_4 FILLER_59_2662 ();
 sg13g2_fill_2 FILLER_59_2666 ();
 sg13g2_decap_8 FILLER_59_2673 ();
 sg13g2_decap_8 FILLER_59_2680 ();
 sg13g2_decap_8 FILLER_59_2687 ();
 sg13g2_decap_8 FILLER_59_2694 ();
 sg13g2_fill_2 FILLER_59_2701 ();
 sg13g2_decap_8 FILLER_59_2717 ();
 sg13g2_decap_8 FILLER_59_2724 ();
 sg13g2_decap_8 FILLER_59_2731 ();
 sg13g2_decap_8 FILLER_59_2738 ();
 sg13g2_fill_2 FILLER_59_2745 ();
 sg13g2_decap_8 FILLER_59_2773 ();
 sg13g2_decap_8 FILLER_59_2780 ();
 sg13g2_decap_8 FILLER_59_2787 ();
 sg13g2_decap_4 FILLER_59_2794 ();
 sg13g2_decap_8 FILLER_59_2804 ();
 sg13g2_decap_8 FILLER_59_2811 ();
 sg13g2_decap_8 FILLER_59_2818 ();
 sg13g2_decap_8 FILLER_59_2825 ();
 sg13g2_decap_8 FILLER_59_2832 ();
 sg13g2_decap_8 FILLER_59_2839 ();
 sg13g2_fill_2 FILLER_59_2846 ();
 sg13g2_decap_8 FILLER_59_2874 ();
 sg13g2_decap_8 FILLER_59_2881 ();
 sg13g2_decap_8 FILLER_59_2888 ();
 sg13g2_decap_8 FILLER_59_2895 ();
 sg13g2_decap_8 FILLER_59_2902 ();
 sg13g2_decap_8 FILLER_59_2909 ();
 sg13g2_decap_8 FILLER_59_2916 ();
 sg13g2_decap_8 FILLER_59_2923 ();
 sg13g2_decap_8 FILLER_59_2930 ();
 sg13g2_decap_8 FILLER_59_2937 ();
 sg13g2_decap_8 FILLER_59_2944 ();
 sg13g2_decap_8 FILLER_59_2951 ();
 sg13g2_decap_8 FILLER_59_2958 ();
 sg13g2_decap_8 FILLER_59_2965 ();
 sg13g2_fill_2 FILLER_59_2972 ();
 sg13g2_decap_8 FILLER_59_2980 ();
 sg13g2_decap_8 FILLER_59_2987 ();
 sg13g2_decap_8 FILLER_59_2994 ();
 sg13g2_fill_1 FILLER_59_3001 ();
 sg13g2_decap_8 FILLER_59_3012 ();
 sg13g2_decap_8 FILLER_59_3019 ();
 sg13g2_decap_8 FILLER_59_3026 ();
 sg13g2_decap_8 FILLER_59_3033 ();
 sg13g2_decap_8 FILLER_59_3040 ();
 sg13g2_decap_8 FILLER_59_3047 ();
 sg13g2_decap_4 FILLER_59_3054 ();
 sg13g2_fill_1 FILLER_59_3058 ();
 sg13g2_decap_8 FILLER_59_3063 ();
 sg13g2_decap_8 FILLER_59_3070 ();
 sg13g2_fill_1 FILLER_59_3077 ();
 sg13g2_decap_8 FILLER_59_3084 ();
 sg13g2_decap_8 FILLER_59_3091 ();
 sg13g2_decap_8 FILLER_59_3098 ();
 sg13g2_fill_2 FILLER_59_3105 ();
 sg13g2_fill_1 FILLER_59_3107 ();
 sg13g2_decap_8 FILLER_59_3113 ();
 sg13g2_decap_8 FILLER_59_3120 ();
 sg13g2_decap_8 FILLER_59_3127 ();
 sg13g2_decap_8 FILLER_59_3134 ();
 sg13g2_decap_8 FILLER_59_3141 ();
 sg13g2_decap_8 FILLER_59_3157 ();
 sg13g2_decap_8 FILLER_59_3164 ();
 sg13g2_decap_8 FILLER_59_3171 ();
 sg13g2_decap_8 FILLER_59_3178 ();
 sg13g2_decap_8 FILLER_59_3185 ();
 sg13g2_decap_4 FILLER_59_3192 ();
 sg13g2_fill_1 FILLER_59_3196 ();
 sg13g2_decap_8 FILLER_59_3202 ();
 sg13g2_decap_8 FILLER_59_3209 ();
 sg13g2_decap_8 FILLER_59_3216 ();
 sg13g2_fill_2 FILLER_59_3223 ();
 sg13g2_fill_1 FILLER_59_3225 ();
 sg13g2_decap_8 FILLER_59_3234 ();
 sg13g2_decap_8 FILLER_59_3241 ();
 sg13g2_decap_4 FILLER_59_3248 ();
 sg13g2_fill_1 FILLER_59_3252 ();
 sg13g2_decap_8 FILLER_59_3289 ();
 sg13g2_decap_8 FILLER_59_3296 ();
 sg13g2_decap_8 FILLER_59_3303 ();
 sg13g2_fill_2 FILLER_59_3310 ();
 sg13g2_fill_1 FILLER_59_3312 ();
 sg13g2_decap_8 FILLER_59_3336 ();
 sg13g2_decap_8 FILLER_59_3343 ();
 sg13g2_decap_8 FILLER_59_3350 ();
 sg13g2_decap_4 FILLER_59_3357 ();
 sg13g2_fill_2 FILLER_59_3361 ();
 sg13g2_decap_8 FILLER_59_3389 ();
 sg13g2_decap_8 FILLER_59_3396 ();
 sg13g2_decap_8 FILLER_59_3403 ();
 sg13g2_decap_8 FILLER_59_3410 ();
 sg13g2_decap_8 FILLER_59_3417 ();
 sg13g2_decap_4 FILLER_59_3424 ();
 sg13g2_decap_8 FILLER_59_3463 ();
 sg13g2_decap_4 FILLER_59_3470 ();
 sg13g2_fill_1 FILLER_59_3474 ();
 sg13g2_decap_8 FILLER_59_3483 ();
 sg13g2_decap_8 FILLER_59_3490 ();
 sg13g2_decap_8 FILLER_59_3497 ();
 sg13g2_decap_4 FILLER_59_3504 ();
 sg13g2_fill_1 FILLER_59_3512 ();
 sg13g2_decap_8 FILLER_59_3542 ();
 sg13g2_fill_2 FILLER_59_3549 ();
 sg13g2_fill_1 FILLER_59_3551 ();
 sg13g2_decap_8 FILLER_59_3561 ();
 sg13g2_decap_8 FILLER_59_3568 ();
 sg13g2_decap_4 FILLER_59_3575 ();
 sg13g2_fill_1 FILLER_59_3579 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_decap_4 FILLER_60_7 ();
 sg13g2_fill_2 FILLER_60_29 ();
 sg13g2_decap_8 FILLER_60_67 ();
 sg13g2_decap_4 FILLER_60_74 ();
 sg13g2_fill_2 FILLER_60_92 ();
 sg13g2_fill_2 FILLER_60_103 ();
 sg13g2_decap_8 FILLER_60_110 ();
 sg13g2_decap_8 FILLER_60_117 ();
 sg13g2_decap_8 FILLER_60_124 ();
 sg13g2_decap_8 FILLER_60_131 ();
 sg13g2_decap_4 FILLER_60_138 ();
 sg13g2_fill_1 FILLER_60_142 ();
 sg13g2_decap_8 FILLER_60_163 ();
 sg13g2_decap_8 FILLER_60_170 ();
 sg13g2_decap_8 FILLER_60_177 ();
 sg13g2_decap_8 FILLER_60_184 ();
 sg13g2_fill_1 FILLER_60_191 ();
 sg13g2_decap_8 FILLER_60_229 ();
 sg13g2_decap_8 FILLER_60_236 ();
 sg13g2_decap_8 FILLER_60_243 ();
 sg13g2_fill_2 FILLER_60_253 ();
 sg13g2_decap_8 FILLER_60_260 ();
 sg13g2_decap_8 FILLER_60_267 ();
 sg13g2_decap_8 FILLER_60_274 ();
 sg13g2_decap_8 FILLER_60_281 ();
 sg13g2_decap_8 FILLER_60_288 ();
 sg13g2_decap_8 FILLER_60_295 ();
 sg13g2_fill_2 FILLER_60_302 ();
 sg13g2_fill_1 FILLER_60_304 ();
 sg13g2_decap_4 FILLER_60_318 ();
 sg13g2_decap_4 FILLER_60_336 ();
 sg13g2_decap_8 FILLER_60_345 ();
 sg13g2_decap_8 FILLER_60_352 ();
 sg13g2_decap_8 FILLER_60_359 ();
 sg13g2_decap_8 FILLER_60_366 ();
 sg13g2_decap_8 FILLER_60_373 ();
 sg13g2_decap_8 FILLER_60_380 ();
 sg13g2_decap_8 FILLER_60_387 ();
 sg13g2_decap_4 FILLER_60_410 ();
 sg13g2_fill_1 FILLER_60_414 ();
 sg13g2_decap_8 FILLER_60_424 ();
 sg13g2_decap_8 FILLER_60_431 ();
 sg13g2_decap_8 FILLER_60_438 ();
 sg13g2_decap_8 FILLER_60_445 ();
 sg13g2_decap_8 FILLER_60_452 ();
 sg13g2_decap_8 FILLER_60_459 ();
 sg13g2_decap_8 FILLER_60_466 ();
 sg13g2_decap_8 FILLER_60_473 ();
 sg13g2_fill_2 FILLER_60_480 ();
 sg13g2_decap_8 FILLER_60_487 ();
 sg13g2_decap_4 FILLER_60_494 ();
 sg13g2_fill_1 FILLER_60_498 ();
 sg13g2_decap_8 FILLER_60_529 ();
 sg13g2_decap_4 FILLER_60_536 ();
 sg13g2_fill_1 FILLER_60_540 ();
 sg13g2_decap_8 FILLER_60_582 ();
 sg13g2_decap_8 FILLER_60_589 ();
 sg13g2_decap_8 FILLER_60_596 ();
 sg13g2_decap_8 FILLER_60_603 ();
 sg13g2_decap_4 FILLER_60_610 ();
 sg13g2_fill_1 FILLER_60_614 ();
 sg13g2_decap_8 FILLER_60_628 ();
 sg13g2_decap_8 FILLER_60_635 ();
 sg13g2_decap_8 FILLER_60_642 ();
 sg13g2_decap_8 FILLER_60_649 ();
 sg13g2_decap_8 FILLER_60_656 ();
 sg13g2_decap_4 FILLER_60_663 ();
 sg13g2_fill_2 FILLER_60_667 ();
 sg13g2_decap_8 FILLER_60_674 ();
 sg13g2_fill_1 FILLER_60_681 ();
 sg13g2_decap_8 FILLER_60_687 ();
 sg13g2_decap_8 FILLER_60_694 ();
 sg13g2_decap_8 FILLER_60_701 ();
 sg13g2_decap_8 FILLER_60_708 ();
 sg13g2_decap_8 FILLER_60_715 ();
 sg13g2_decap_8 FILLER_60_722 ();
 sg13g2_decap_8 FILLER_60_729 ();
 sg13g2_decap_8 FILLER_60_736 ();
 sg13g2_decap_8 FILLER_60_743 ();
 sg13g2_decap_8 FILLER_60_750 ();
 sg13g2_decap_8 FILLER_60_757 ();
 sg13g2_decap_8 FILLER_60_764 ();
 sg13g2_decap_8 FILLER_60_779 ();
 sg13g2_decap_8 FILLER_60_786 ();
 sg13g2_decap_8 FILLER_60_793 ();
 sg13g2_decap_8 FILLER_60_800 ();
 sg13g2_decap_8 FILLER_60_807 ();
 sg13g2_decap_8 FILLER_60_814 ();
 sg13g2_fill_2 FILLER_60_821 ();
 sg13g2_fill_1 FILLER_60_823 ();
 sg13g2_decap_8 FILLER_60_828 ();
 sg13g2_fill_2 FILLER_60_835 ();
 sg13g2_decap_8 FILLER_60_842 ();
 sg13g2_decap_8 FILLER_60_849 ();
 sg13g2_decap_8 FILLER_60_856 ();
 sg13g2_decap_8 FILLER_60_863 ();
 sg13g2_decap_8 FILLER_60_870 ();
 sg13g2_decap_8 FILLER_60_877 ();
 sg13g2_decap_8 FILLER_60_884 ();
 sg13g2_decap_8 FILLER_60_891 ();
 sg13g2_decap_8 FILLER_60_898 ();
 sg13g2_decap_8 FILLER_60_905 ();
 sg13g2_decap_8 FILLER_60_912 ();
 sg13g2_decap_8 FILLER_60_919 ();
 sg13g2_decap_8 FILLER_60_926 ();
 sg13g2_decap_8 FILLER_60_933 ();
 sg13g2_fill_2 FILLER_60_940 ();
 sg13g2_fill_1 FILLER_60_942 ();
 sg13g2_decap_8 FILLER_60_956 ();
 sg13g2_decap_8 FILLER_60_963 ();
 sg13g2_decap_8 FILLER_60_970 ();
 sg13g2_decap_8 FILLER_60_977 ();
 sg13g2_decap_8 FILLER_60_984 ();
 sg13g2_decap_8 FILLER_60_991 ();
 sg13g2_decap_8 FILLER_60_998 ();
 sg13g2_decap_8 FILLER_60_1005 ();
 sg13g2_decap_8 FILLER_60_1012 ();
 sg13g2_decap_8 FILLER_60_1019 ();
 sg13g2_decap_8 FILLER_60_1026 ();
 sg13g2_decap_8 FILLER_60_1033 ();
 sg13g2_decap_8 FILLER_60_1040 ();
 sg13g2_decap_8 FILLER_60_1047 ();
 sg13g2_decap_8 FILLER_60_1054 ();
 sg13g2_decap_8 FILLER_60_1061 ();
 sg13g2_decap_8 FILLER_60_1068 ();
 sg13g2_decap_8 FILLER_60_1075 ();
 sg13g2_decap_8 FILLER_60_1082 ();
 sg13g2_decap_8 FILLER_60_1089 ();
 sg13g2_decap_8 FILLER_60_1096 ();
 sg13g2_decap_8 FILLER_60_1103 ();
 sg13g2_decap_8 FILLER_60_1110 ();
 sg13g2_decap_8 FILLER_60_1117 ();
 sg13g2_decap_8 FILLER_60_1124 ();
 sg13g2_fill_2 FILLER_60_1131 ();
 sg13g2_fill_1 FILLER_60_1133 ();
 sg13g2_decap_4 FILLER_60_1160 ();
 sg13g2_fill_1 FILLER_60_1164 ();
 sg13g2_decap_8 FILLER_60_1178 ();
 sg13g2_decap_8 FILLER_60_1185 ();
 sg13g2_fill_2 FILLER_60_1192 ();
 sg13g2_decap_4 FILLER_60_1197 ();
 sg13g2_fill_2 FILLER_60_1210 ();
 sg13g2_decap_4 FILLER_60_1243 ();
 sg13g2_fill_1 FILLER_60_1247 ();
 sg13g2_fill_2 FILLER_60_1263 ();
 sg13g2_decap_8 FILLER_60_1281 ();
 sg13g2_decap_8 FILLER_60_1288 ();
 sg13g2_decap_8 FILLER_60_1295 ();
 sg13g2_decap_8 FILLER_60_1302 ();
 sg13g2_decap_8 FILLER_60_1309 ();
 sg13g2_decap_8 FILLER_60_1316 ();
 sg13g2_decap_8 FILLER_60_1323 ();
 sg13g2_fill_2 FILLER_60_1330 ();
 sg13g2_fill_1 FILLER_60_1332 ();
 sg13g2_decap_4 FILLER_60_1369 ();
 sg13g2_decap_8 FILLER_60_1409 ();
 sg13g2_decap_8 FILLER_60_1416 ();
 sg13g2_decap_8 FILLER_60_1423 ();
 sg13g2_decap_8 FILLER_60_1430 ();
 sg13g2_decap_4 FILLER_60_1437 ();
 sg13g2_fill_2 FILLER_60_1441 ();
 sg13g2_fill_2 FILLER_60_1453 ();
 sg13g2_fill_1 FILLER_60_1455 ();
 sg13g2_decap_8 FILLER_60_1482 ();
 sg13g2_decap_8 FILLER_60_1489 ();
 sg13g2_decap_4 FILLER_60_1496 ();
 sg13g2_fill_1 FILLER_60_1500 ();
 sg13g2_fill_1 FILLER_60_1509 ();
 sg13g2_fill_2 FILLER_60_1520 ();
 sg13g2_fill_1 FILLER_60_1522 ();
 sg13g2_decap_8 FILLER_60_1549 ();
 sg13g2_decap_8 FILLER_60_1556 ();
 sg13g2_decap_4 FILLER_60_1563 ();
 sg13g2_decap_8 FILLER_60_1587 ();
 sg13g2_decap_8 FILLER_60_1594 ();
 sg13g2_decap_4 FILLER_60_1601 ();
 sg13g2_fill_1 FILLER_60_1605 ();
 sg13g2_decap_8 FILLER_60_1610 ();
 sg13g2_decap_8 FILLER_60_1617 ();
 sg13g2_decap_8 FILLER_60_1624 ();
 sg13g2_decap_8 FILLER_60_1631 ();
 sg13g2_decap_8 FILLER_60_1638 ();
 sg13g2_decap_8 FILLER_60_1645 ();
 sg13g2_decap_8 FILLER_60_1652 ();
 sg13g2_fill_1 FILLER_60_1659 ();
 sg13g2_decap_8 FILLER_60_1686 ();
 sg13g2_decap_8 FILLER_60_1693 ();
 sg13g2_fill_2 FILLER_60_1700 ();
 sg13g2_decap_8 FILLER_60_1733 ();
 sg13g2_decap_8 FILLER_60_1740 ();
 sg13g2_decap_8 FILLER_60_1747 ();
 sg13g2_decap_8 FILLER_60_1754 ();
 sg13g2_decap_4 FILLER_60_1761 ();
 sg13g2_fill_1 FILLER_60_1765 ();
 sg13g2_decap_8 FILLER_60_1798 ();
 sg13g2_decap_8 FILLER_60_1805 ();
 sg13g2_fill_2 FILLER_60_1812 ();
 sg13g2_fill_1 FILLER_60_1830 ();
 sg13g2_decap_8 FILLER_60_1849 ();
 sg13g2_decap_8 FILLER_60_1856 ();
 sg13g2_decap_8 FILLER_60_1863 ();
 sg13g2_decap_8 FILLER_60_1870 ();
 sg13g2_decap_8 FILLER_60_1877 ();
 sg13g2_decap_8 FILLER_60_1884 ();
 sg13g2_decap_8 FILLER_60_1891 ();
 sg13g2_decap_8 FILLER_60_1898 ();
 sg13g2_decap_4 FILLER_60_1905 ();
 sg13g2_fill_1 FILLER_60_1909 ();
 sg13g2_decap_8 FILLER_60_1936 ();
 sg13g2_decap_8 FILLER_60_1943 ();
 sg13g2_decap_8 FILLER_60_1950 ();
 sg13g2_decap_8 FILLER_60_1957 ();
 sg13g2_decap_8 FILLER_60_1964 ();
 sg13g2_decap_8 FILLER_60_1971 ();
 sg13g2_decap_4 FILLER_60_1992 ();
 sg13g2_fill_1 FILLER_60_1996 ();
 sg13g2_decap_8 FILLER_60_2011 ();
 sg13g2_decap_8 FILLER_60_2018 ();
 sg13g2_fill_2 FILLER_60_2025 ();
 sg13g2_decap_8 FILLER_60_2033 ();
 sg13g2_decap_4 FILLER_60_2040 ();
 sg13g2_decap_8 FILLER_60_2094 ();
 sg13g2_decap_8 FILLER_60_2101 ();
 sg13g2_decap_4 FILLER_60_2108 ();
 sg13g2_fill_2 FILLER_60_2112 ();
 sg13g2_decap_8 FILLER_60_2120 ();
 sg13g2_fill_2 FILLER_60_2127 ();
 sg13g2_fill_1 FILLER_60_2129 ();
 sg13g2_decap_8 FILLER_60_2136 ();
 sg13g2_decap_8 FILLER_60_2143 ();
 sg13g2_decap_8 FILLER_60_2150 ();
 sg13g2_decap_8 FILLER_60_2157 ();
 sg13g2_decap_8 FILLER_60_2164 ();
 sg13g2_decap_8 FILLER_60_2171 ();
 sg13g2_decap_8 FILLER_60_2178 ();
 sg13g2_decap_4 FILLER_60_2185 ();
 sg13g2_fill_1 FILLER_60_2189 ();
 sg13g2_decap_8 FILLER_60_2196 ();
 sg13g2_decap_8 FILLER_60_2203 ();
 sg13g2_decap_4 FILLER_60_2210 ();
 sg13g2_fill_2 FILLER_60_2214 ();
 sg13g2_decap_8 FILLER_60_2224 ();
 sg13g2_decap_8 FILLER_60_2231 ();
 sg13g2_decap_8 FILLER_60_2238 ();
 sg13g2_fill_1 FILLER_60_2245 ();
 sg13g2_fill_1 FILLER_60_2254 ();
 sg13g2_fill_2 FILLER_60_2284 ();
 sg13g2_decap_4 FILLER_60_2307 ();
 sg13g2_fill_1 FILLER_60_2311 ();
 sg13g2_decap_8 FILLER_60_2323 ();
 sg13g2_decap_8 FILLER_60_2330 ();
 sg13g2_decap_8 FILLER_60_2340 ();
 sg13g2_fill_1 FILLER_60_2347 ();
 sg13g2_decap_8 FILLER_60_2353 ();
 sg13g2_fill_2 FILLER_60_2360 ();
 sg13g2_fill_1 FILLER_60_2362 ();
 sg13g2_decap_8 FILLER_60_2380 ();
 sg13g2_decap_8 FILLER_60_2387 ();
 sg13g2_decap_8 FILLER_60_2394 ();
 sg13g2_decap_8 FILLER_60_2401 ();
 sg13g2_fill_2 FILLER_60_2408 ();
 sg13g2_decap_8 FILLER_60_2420 ();
 sg13g2_decap_8 FILLER_60_2427 ();
 sg13g2_decap_8 FILLER_60_2434 ();
 sg13g2_decap_8 FILLER_60_2441 ();
 sg13g2_decap_8 FILLER_60_2448 ();
 sg13g2_decap_8 FILLER_60_2455 ();
 sg13g2_decap_8 FILLER_60_2462 ();
 sg13g2_decap_8 FILLER_60_2469 ();
 sg13g2_fill_2 FILLER_60_2476 ();
 sg13g2_fill_1 FILLER_60_2478 ();
 sg13g2_decap_8 FILLER_60_2505 ();
 sg13g2_decap_8 FILLER_60_2512 ();
 sg13g2_decap_8 FILLER_60_2519 ();
 sg13g2_decap_8 FILLER_60_2526 ();
 sg13g2_decap_8 FILLER_60_2533 ();
 sg13g2_decap_8 FILLER_60_2540 ();
 sg13g2_decap_8 FILLER_60_2547 ();
 sg13g2_decap_8 FILLER_60_2554 ();
 sg13g2_decap_8 FILLER_60_2561 ();
 sg13g2_decap_8 FILLER_60_2568 ();
 sg13g2_decap_8 FILLER_60_2575 ();
 sg13g2_decap_8 FILLER_60_2582 ();
 sg13g2_decap_8 FILLER_60_2589 ();
 sg13g2_fill_1 FILLER_60_2596 ();
 sg13g2_decap_8 FILLER_60_2623 ();
 sg13g2_decap_8 FILLER_60_2630 ();
 sg13g2_decap_4 FILLER_60_2637 ();
 sg13g2_fill_2 FILLER_60_2641 ();
 sg13g2_decap_8 FILLER_60_2669 ();
 sg13g2_decap_8 FILLER_60_2676 ();
 sg13g2_decap_8 FILLER_60_2683 ();
 sg13g2_decap_8 FILLER_60_2690 ();
 sg13g2_decap_8 FILLER_60_2697 ();
 sg13g2_decap_4 FILLER_60_2704 ();
 sg13g2_fill_2 FILLER_60_2708 ();
 sg13g2_decap_4 FILLER_60_2722 ();
 sg13g2_fill_1 FILLER_60_2726 ();
 sg13g2_decap_8 FILLER_60_2748 ();
 sg13g2_decap_8 FILLER_60_2755 ();
 sg13g2_decap_8 FILLER_60_2762 ();
 sg13g2_fill_1 FILLER_60_2769 ();
 sg13g2_decap_8 FILLER_60_2778 ();
 sg13g2_fill_2 FILLER_60_2795 ();
 sg13g2_fill_1 FILLER_60_2797 ();
 sg13g2_decap_8 FILLER_60_2824 ();
 sg13g2_decap_8 FILLER_60_2831 ();
 sg13g2_decap_8 FILLER_60_2838 ();
 sg13g2_decap_8 FILLER_60_2871 ();
 sg13g2_decap_8 FILLER_60_2878 ();
 sg13g2_decap_4 FILLER_60_2885 ();
 sg13g2_fill_1 FILLER_60_2897 ();
 sg13g2_fill_2 FILLER_60_2903 ();
 sg13g2_fill_1 FILLER_60_2905 ();
 sg13g2_fill_2 FILLER_60_2916 ();
 sg13g2_decap_4 FILLER_60_2939 ();
 sg13g2_fill_1 FILLER_60_2943 ();
 sg13g2_decap_8 FILLER_60_2962 ();
 sg13g2_decap_8 FILLER_60_2969 ();
 sg13g2_decap_8 FILLER_60_2976 ();
 sg13g2_decap_8 FILLER_60_2983 ();
 sg13g2_decap_8 FILLER_60_2990 ();
 sg13g2_decap_4 FILLER_60_2997 ();
 sg13g2_fill_1 FILLER_60_3001 ();
 sg13g2_decap_8 FILLER_60_3015 ();
 sg13g2_fill_2 FILLER_60_3022 ();
 sg13g2_fill_1 FILLER_60_3024 ();
 sg13g2_decap_8 FILLER_60_3038 ();
 sg13g2_decap_8 FILLER_60_3045 ();
 sg13g2_decap_8 FILLER_60_3052 ();
 sg13g2_fill_2 FILLER_60_3059 ();
 sg13g2_decap_8 FILLER_60_3087 ();
 sg13g2_decap_4 FILLER_60_3094 ();
 sg13g2_decap_8 FILLER_60_3116 ();
 sg13g2_decap_8 FILLER_60_3123 ();
 sg13g2_decap_8 FILLER_60_3130 ();
 sg13g2_decap_4 FILLER_60_3137 ();
 sg13g2_fill_2 FILLER_60_3141 ();
 sg13g2_decap_8 FILLER_60_3159 ();
 sg13g2_decap_8 FILLER_60_3166 ();
 sg13g2_decap_8 FILLER_60_3173 ();
 sg13g2_decap_8 FILLER_60_3180 ();
 sg13g2_decap_8 FILLER_60_3187 ();
 sg13g2_decap_8 FILLER_60_3194 ();
 sg13g2_decap_8 FILLER_60_3201 ();
 sg13g2_decap_8 FILLER_60_3208 ();
 sg13g2_decap_8 FILLER_60_3215 ();
 sg13g2_decap_8 FILLER_60_3222 ();
 sg13g2_decap_8 FILLER_60_3229 ();
 sg13g2_decap_8 FILLER_60_3236 ();
 sg13g2_decap_8 FILLER_60_3243 ();
 sg13g2_decap_8 FILLER_60_3250 ();
 sg13g2_decap_8 FILLER_60_3257 ();
 sg13g2_decap_8 FILLER_60_3264 ();
 sg13g2_decap_8 FILLER_60_3271 ();
 sg13g2_fill_2 FILLER_60_3278 ();
 sg13g2_fill_1 FILLER_60_3280 ();
 sg13g2_decap_8 FILLER_60_3291 ();
 sg13g2_decap_8 FILLER_60_3298 ();
 sg13g2_decap_8 FILLER_60_3305 ();
 sg13g2_decap_8 FILLER_60_3312 ();
 sg13g2_decap_8 FILLER_60_3319 ();
 sg13g2_decap_8 FILLER_60_3326 ();
 sg13g2_decap_8 FILLER_60_3333 ();
 sg13g2_decap_8 FILLER_60_3340 ();
 sg13g2_decap_8 FILLER_60_3347 ();
 sg13g2_decap_8 FILLER_60_3354 ();
 sg13g2_decap_8 FILLER_60_3361 ();
 sg13g2_decap_8 FILLER_60_3368 ();
 sg13g2_decap_8 FILLER_60_3375 ();
 sg13g2_decap_8 FILLER_60_3382 ();
 sg13g2_decap_8 FILLER_60_3389 ();
 sg13g2_decap_8 FILLER_60_3396 ();
 sg13g2_decap_8 FILLER_60_3403 ();
 sg13g2_decap_8 FILLER_60_3410 ();
 sg13g2_decap_8 FILLER_60_3417 ();
 sg13g2_fill_2 FILLER_60_3424 ();
 sg13g2_fill_1 FILLER_60_3426 ();
 sg13g2_decap_8 FILLER_60_3456 ();
 sg13g2_decap_8 FILLER_60_3463 ();
 sg13g2_decap_8 FILLER_60_3470 ();
 sg13g2_decap_8 FILLER_60_3477 ();
 sg13g2_decap_8 FILLER_60_3484 ();
 sg13g2_decap_8 FILLER_60_3491 ();
 sg13g2_decap_4 FILLER_60_3498 ();
 sg13g2_fill_1 FILLER_60_3502 ();
 sg13g2_decap_8 FILLER_60_3538 ();
 sg13g2_fill_1 FILLER_60_3545 ();
 sg13g2_decap_8 FILLER_60_3572 ();
 sg13g2_fill_1 FILLER_60_3579 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_decap_8 FILLER_61_7 ();
 sg13g2_decap_4 FILLER_61_14 ();
 sg13g2_fill_2 FILLER_61_18 ();
 sg13g2_fill_2 FILLER_61_30 ();
 sg13g2_fill_1 FILLER_61_32 ();
 sg13g2_decap_8 FILLER_61_42 ();
 sg13g2_decap_8 FILLER_61_54 ();
 sg13g2_decap_8 FILLER_61_61 ();
 sg13g2_decap_4 FILLER_61_68 ();
 sg13g2_fill_2 FILLER_61_72 ();
 sg13g2_decap_8 FILLER_61_110 ();
 sg13g2_decap_8 FILLER_61_117 ();
 sg13g2_decap_8 FILLER_61_124 ();
 sg13g2_decap_8 FILLER_61_131 ();
 sg13g2_decap_8 FILLER_61_138 ();
 sg13g2_fill_2 FILLER_61_145 ();
 sg13g2_fill_1 FILLER_61_147 ();
 sg13g2_decap_8 FILLER_61_163 ();
 sg13g2_decap_8 FILLER_61_170 ();
 sg13g2_decap_8 FILLER_61_177 ();
 sg13g2_decap_8 FILLER_61_184 ();
 sg13g2_decap_4 FILLER_61_191 ();
 sg13g2_fill_2 FILLER_61_195 ();
 sg13g2_decap_8 FILLER_61_203 ();
 sg13g2_decap_8 FILLER_61_219 ();
 sg13g2_decap_8 FILLER_61_226 ();
 sg13g2_decap_4 FILLER_61_236 ();
 sg13g2_fill_1 FILLER_61_252 ();
 sg13g2_decap_8 FILLER_61_269 ();
 sg13g2_decap_8 FILLER_61_276 ();
 sg13g2_decap_8 FILLER_61_283 ();
 sg13g2_decap_8 FILLER_61_290 ();
 sg13g2_decap_8 FILLER_61_297 ();
 sg13g2_fill_1 FILLER_61_304 ();
 sg13g2_fill_2 FILLER_61_318 ();
 sg13g2_fill_1 FILLER_61_320 ();
 sg13g2_decap_8 FILLER_61_337 ();
 sg13g2_decap_8 FILLER_61_344 ();
 sg13g2_decap_4 FILLER_61_351 ();
 sg13g2_fill_1 FILLER_61_355 ();
 sg13g2_decap_8 FILLER_61_364 ();
 sg13g2_decap_8 FILLER_61_371 ();
 sg13g2_decap_8 FILLER_61_378 ();
 sg13g2_decap_8 FILLER_61_385 ();
 sg13g2_decap_8 FILLER_61_392 ();
 sg13g2_fill_2 FILLER_61_399 ();
 sg13g2_fill_1 FILLER_61_401 ();
 sg13g2_decap_8 FILLER_61_407 ();
 sg13g2_decap_8 FILLER_61_414 ();
 sg13g2_decap_8 FILLER_61_421 ();
 sg13g2_decap_8 FILLER_61_428 ();
 sg13g2_decap_8 FILLER_61_435 ();
 sg13g2_decap_8 FILLER_61_442 ();
 sg13g2_decap_8 FILLER_61_449 ();
 sg13g2_decap_8 FILLER_61_456 ();
 sg13g2_decap_4 FILLER_61_463 ();
 sg13g2_decap_8 FILLER_61_479 ();
 sg13g2_fill_1 FILLER_61_486 ();
 sg13g2_decap_8 FILLER_61_509 ();
 sg13g2_decap_8 FILLER_61_516 ();
 sg13g2_decap_8 FILLER_61_523 ();
 sg13g2_decap_8 FILLER_61_530 ();
 sg13g2_decap_8 FILLER_61_537 ();
 sg13g2_fill_2 FILLER_61_544 ();
 sg13g2_fill_1 FILLER_61_546 ();
 sg13g2_fill_1 FILLER_61_571 ();
 sg13g2_decap_8 FILLER_61_580 ();
 sg13g2_decap_8 FILLER_61_587 ();
 sg13g2_decap_8 FILLER_61_594 ();
 sg13g2_fill_2 FILLER_61_601 ();
 sg13g2_fill_1 FILLER_61_603 ();
 sg13g2_decap_4 FILLER_61_625 ();
 sg13g2_fill_1 FILLER_61_629 ();
 sg13g2_decap_8 FILLER_61_638 ();
 sg13g2_decap_8 FILLER_61_645 ();
 sg13g2_decap_8 FILLER_61_652 ();
 sg13g2_decap_8 FILLER_61_659 ();
 sg13g2_decap_4 FILLER_61_666 ();
 sg13g2_fill_2 FILLER_61_684 ();
 sg13g2_decap_4 FILLER_61_702 ();
 sg13g2_fill_2 FILLER_61_706 ();
 sg13g2_decap_8 FILLER_61_735 ();
 sg13g2_decap_4 FILLER_61_742 ();
 sg13g2_fill_2 FILLER_61_746 ();
 sg13g2_decap_8 FILLER_61_783 ();
 sg13g2_decap_8 FILLER_61_790 ();
 sg13g2_fill_1 FILLER_61_797 ();
 sg13g2_decap_8 FILLER_61_806 ();
 sg13g2_decap_8 FILLER_61_813 ();
 sg13g2_decap_8 FILLER_61_820 ();
 sg13g2_decap_8 FILLER_61_827 ();
 sg13g2_decap_8 FILLER_61_834 ();
 sg13g2_decap_8 FILLER_61_841 ();
 sg13g2_fill_1 FILLER_61_848 ();
 sg13g2_decap_8 FILLER_61_857 ();
 sg13g2_decap_4 FILLER_61_864 ();
 sg13g2_fill_2 FILLER_61_868 ();
 sg13g2_decap_8 FILLER_61_877 ();
 sg13g2_decap_8 FILLER_61_884 ();
 sg13g2_decap_8 FILLER_61_891 ();
 sg13g2_decap_8 FILLER_61_898 ();
 sg13g2_decap_8 FILLER_61_905 ();
 sg13g2_decap_8 FILLER_61_912 ();
 sg13g2_fill_2 FILLER_61_919 ();
 sg13g2_decap_8 FILLER_61_935 ();
 sg13g2_decap_8 FILLER_61_942 ();
 sg13g2_decap_8 FILLER_61_949 ();
 sg13g2_fill_1 FILLER_61_956 ();
 sg13g2_decap_4 FILLER_61_983 ();
 sg13g2_fill_1 FILLER_61_987 ();
 sg13g2_decap_8 FILLER_61_991 ();
 sg13g2_decap_8 FILLER_61_998 ();
 sg13g2_decap_8 FILLER_61_1005 ();
 sg13g2_decap_8 FILLER_61_1012 ();
 sg13g2_decap_8 FILLER_61_1019 ();
 sg13g2_decap_4 FILLER_61_1035 ();
 sg13g2_decap_8 FILLER_61_1047 ();
 sg13g2_decap_8 FILLER_61_1054 ();
 sg13g2_decap_4 FILLER_61_1061 ();
 sg13g2_fill_1 FILLER_61_1065 ();
 sg13g2_fill_2 FILLER_61_1083 ();
 sg13g2_decap_8 FILLER_61_1102 ();
 sg13g2_decap_8 FILLER_61_1109 ();
 sg13g2_fill_2 FILLER_61_1124 ();
 sg13g2_fill_1 FILLER_61_1126 ();
 sg13g2_fill_2 FILLER_61_1153 ();
 sg13g2_fill_2 FILLER_61_1163 ();
 sg13g2_decap_8 FILLER_61_1191 ();
 sg13g2_decap_8 FILLER_61_1198 ();
 sg13g2_decap_8 FILLER_61_1205 ();
 sg13g2_decap_8 FILLER_61_1212 ();
 sg13g2_decap_8 FILLER_61_1219 ();
 sg13g2_decap_8 FILLER_61_1226 ();
 sg13g2_decap_8 FILLER_61_1233 ();
 sg13g2_fill_2 FILLER_61_1252 ();
 sg13g2_decap_8 FILLER_61_1271 ();
 sg13g2_decap_4 FILLER_61_1278 ();
 sg13g2_decap_8 FILLER_61_1286 ();
 sg13g2_decap_8 FILLER_61_1293 ();
 sg13g2_fill_2 FILLER_61_1308 ();
 sg13g2_decap_4 FILLER_61_1314 ();
 sg13g2_decap_8 FILLER_61_1338 ();
 sg13g2_decap_8 FILLER_61_1345 ();
 sg13g2_decap_8 FILLER_61_1352 ();
 sg13g2_decap_8 FILLER_61_1359 ();
 sg13g2_decap_8 FILLER_61_1366 ();
 sg13g2_decap_8 FILLER_61_1373 ();
 sg13g2_decap_8 FILLER_61_1380 ();
 sg13g2_decap_8 FILLER_61_1387 ();
 sg13g2_decap_8 FILLER_61_1394 ();
 sg13g2_decap_8 FILLER_61_1401 ();
 sg13g2_decap_8 FILLER_61_1408 ();
 sg13g2_decap_8 FILLER_61_1415 ();
 sg13g2_decap_8 FILLER_61_1422 ();
 sg13g2_decap_8 FILLER_61_1429 ();
 sg13g2_decap_8 FILLER_61_1436 ();
 sg13g2_decap_8 FILLER_61_1443 ();
 sg13g2_decap_8 FILLER_61_1450 ();
 sg13g2_fill_2 FILLER_61_1457 ();
 sg13g2_decap_8 FILLER_61_1485 ();
 sg13g2_decap_8 FILLER_61_1492 ();
 sg13g2_decap_8 FILLER_61_1499 ();
 sg13g2_decap_8 FILLER_61_1506 ();
 sg13g2_decap_8 FILLER_61_1513 ();
 sg13g2_decap_4 FILLER_61_1520 ();
 sg13g2_fill_1 FILLER_61_1524 ();
 sg13g2_decap_8 FILLER_61_1535 ();
 sg13g2_decap_8 FILLER_61_1542 ();
 sg13g2_decap_8 FILLER_61_1549 ();
 sg13g2_decap_8 FILLER_61_1556 ();
 sg13g2_decap_8 FILLER_61_1563 ();
 sg13g2_fill_2 FILLER_61_1570 ();
 sg13g2_decap_8 FILLER_61_1599 ();
 sg13g2_decap_8 FILLER_61_1606 ();
 sg13g2_decap_8 FILLER_61_1613 ();
 sg13g2_decap_8 FILLER_61_1620 ();
 sg13g2_decap_4 FILLER_61_1627 ();
 sg13g2_fill_2 FILLER_61_1631 ();
 sg13g2_decap_8 FILLER_61_1642 ();
 sg13g2_fill_2 FILLER_61_1649 ();
 sg13g2_fill_1 FILLER_61_1651 ();
 sg13g2_decap_8 FILLER_61_1666 ();
 sg13g2_decap_8 FILLER_61_1673 ();
 sg13g2_decap_8 FILLER_61_1680 ();
 sg13g2_decap_8 FILLER_61_1687 ();
 sg13g2_decap_8 FILLER_61_1694 ();
 sg13g2_decap_8 FILLER_61_1701 ();
 sg13g2_decap_8 FILLER_61_1708 ();
 sg13g2_decap_8 FILLER_61_1715 ();
 sg13g2_decap_8 FILLER_61_1722 ();
 sg13g2_decap_8 FILLER_61_1729 ();
 sg13g2_decap_8 FILLER_61_1736 ();
 sg13g2_decap_8 FILLER_61_1743 ();
 sg13g2_decap_8 FILLER_61_1750 ();
 sg13g2_decap_8 FILLER_61_1757 ();
 sg13g2_decap_8 FILLER_61_1764 ();
 sg13g2_decap_8 FILLER_61_1804 ();
 sg13g2_decap_8 FILLER_61_1811 ();
 sg13g2_decap_8 FILLER_61_1818 ();
 sg13g2_decap_8 FILLER_61_1825 ();
 sg13g2_decap_8 FILLER_61_1832 ();
 sg13g2_decap_8 FILLER_61_1839 ();
 sg13g2_decap_8 FILLER_61_1846 ();
 sg13g2_decap_8 FILLER_61_1853 ();
 sg13g2_decap_8 FILLER_61_1860 ();
 sg13g2_decap_8 FILLER_61_1867 ();
 sg13g2_decap_8 FILLER_61_1874 ();
 sg13g2_decap_8 FILLER_61_1881 ();
 sg13g2_decap_8 FILLER_61_1888 ();
 sg13g2_fill_2 FILLER_61_1895 ();
 sg13g2_fill_2 FILLER_61_1928 ();
 sg13g2_decap_8 FILLER_61_1946 ();
 sg13g2_decap_4 FILLER_61_1953 ();
 sg13g2_fill_1 FILLER_61_1957 ();
 sg13g2_decap_8 FILLER_61_1966 ();
 sg13g2_decap_8 FILLER_61_1973 ();
 sg13g2_decap_8 FILLER_61_1998 ();
 sg13g2_decap_8 FILLER_61_2005 ();
 sg13g2_decap_8 FILLER_61_2012 ();
 sg13g2_decap_8 FILLER_61_2019 ();
 sg13g2_decap_8 FILLER_61_2026 ();
 sg13g2_decap_8 FILLER_61_2033 ();
 sg13g2_decap_4 FILLER_61_2040 ();
 sg13g2_fill_2 FILLER_61_2044 ();
 sg13g2_decap_4 FILLER_61_2061 ();
 sg13g2_decap_8 FILLER_61_2068 ();
 sg13g2_decap_8 FILLER_61_2075 ();
 sg13g2_decap_8 FILLER_61_2082 ();
 sg13g2_decap_8 FILLER_61_2089 ();
 sg13g2_decap_8 FILLER_61_2096 ();
 sg13g2_decap_8 FILLER_61_2103 ();
 sg13g2_decap_8 FILLER_61_2110 ();
 sg13g2_decap_8 FILLER_61_2117 ();
 sg13g2_decap_8 FILLER_61_2124 ();
 sg13g2_decap_8 FILLER_61_2131 ();
 sg13g2_decap_8 FILLER_61_2138 ();
 sg13g2_decap_8 FILLER_61_2145 ();
 sg13g2_decap_8 FILLER_61_2152 ();
 sg13g2_decap_8 FILLER_61_2159 ();
 sg13g2_decap_8 FILLER_61_2166 ();
 sg13g2_decap_8 FILLER_61_2173 ();
 sg13g2_decap_4 FILLER_61_2180 ();
 sg13g2_fill_2 FILLER_61_2184 ();
 sg13g2_decap_8 FILLER_61_2211 ();
 sg13g2_decap_8 FILLER_61_2218 ();
 sg13g2_decap_8 FILLER_61_2225 ();
 sg13g2_fill_1 FILLER_61_2249 ();
 sg13g2_decap_8 FILLER_61_2273 ();
 sg13g2_fill_1 FILLER_61_2280 ();
 sg13g2_decap_8 FILLER_61_2284 ();
 sg13g2_decap_8 FILLER_61_2291 ();
 sg13g2_decap_8 FILLER_61_2298 ();
 sg13g2_decap_8 FILLER_61_2305 ();
 sg13g2_decap_8 FILLER_61_2312 ();
 sg13g2_decap_8 FILLER_61_2319 ();
 sg13g2_decap_8 FILLER_61_2326 ();
 sg13g2_decap_8 FILLER_61_2333 ();
 sg13g2_decap_8 FILLER_61_2340 ();
 sg13g2_decap_4 FILLER_61_2347 ();
 sg13g2_fill_1 FILLER_61_2351 ();
 sg13g2_decap_8 FILLER_61_2357 ();
 sg13g2_decap_8 FILLER_61_2364 ();
 sg13g2_decap_8 FILLER_61_2371 ();
 sg13g2_decap_8 FILLER_61_2378 ();
 sg13g2_decap_8 FILLER_61_2385 ();
 sg13g2_decap_8 FILLER_61_2392 ();
 sg13g2_fill_1 FILLER_61_2399 ();
 sg13g2_decap_8 FILLER_61_2410 ();
 sg13g2_decap_8 FILLER_61_2417 ();
 sg13g2_decap_8 FILLER_61_2424 ();
 sg13g2_decap_8 FILLER_61_2431 ();
 sg13g2_decap_8 FILLER_61_2438 ();
 sg13g2_decap_8 FILLER_61_2445 ();
 sg13g2_decap_8 FILLER_61_2452 ();
 sg13g2_decap_8 FILLER_61_2459 ();
 sg13g2_decap_8 FILLER_61_2466 ();
 sg13g2_decap_8 FILLER_61_2473 ();
 sg13g2_decap_8 FILLER_61_2480 ();
 sg13g2_decap_8 FILLER_61_2487 ();
 sg13g2_decap_8 FILLER_61_2494 ();
 sg13g2_decap_8 FILLER_61_2501 ();
 sg13g2_decap_8 FILLER_61_2508 ();
 sg13g2_decap_8 FILLER_61_2515 ();
 sg13g2_decap_4 FILLER_61_2522 ();
 sg13g2_fill_1 FILLER_61_2531 ();
 sg13g2_decap_8 FILLER_61_2540 ();
 sg13g2_decap_8 FILLER_61_2573 ();
 sg13g2_decap_8 FILLER_61_2580 ();
 sg13g2_decap_8 FILLER_61_2587 ();
 sg13g2_decap_8 FILLER_61_2594 ();
 sg13g2_decap_8 FILLER_61_2601 ();
 sg13g2_decap_8 FILLER_61_2608 ();
 sg13g2_fill_2 FILLER_61_2629 ();
 sg13g2_decap_8 FILLER_61_2667 ();
 sg13g2_decap_4 FILLER_61_2674 ();
 sg13g2_fill_2 FILLER_61_2678 ();
 sg13g2_decap_8 FILLER_61_2686 ();
 sg13g2_decap_8 FILLER_61_2693 ();
 sg13g2_decap_4 FILLER_61_2700 ();
 sg13g2_fill_1 FILLER_61_2704 ();
 sg13g2_decap_8 FILLER_61_2715 ();
 sg13g2_fill_2 FILLER_61_2722 ();
 sg13g2_fill_1 FILLER_61_2724 ();
 sg13g2_decap_8 FILLER_61_2733 ();
 sg13g2_decap_8 FILLER_61_2740 ();
 sg13g2_decap_8 FILLER_61_2747 ();
 sg13g2_decap_8 FILLER_61_2754 ();
 sg13g2_fill_2 FILLER_61_2761 ();
 sg13g2_decap_8 FILLER_61_2768 ();
 sg13g2_decap_8 FILLER_61_2775 ();
 sg13g2_decap_8 FILLER_61_2818 ();
 sg13g2_decap_8 FILLER_61_2825 ();
 sg13g2_decap_4 FILLER_61_2832 ();
 sg13g2_fill_1 FILLER_61_2836 ();
 sg13g2_decap_8 FILLER_61_2873 ();
 sg13g2_decap_8 FILLER_61_2880 ();
 sg13g2_decap_8 FILLER_61_2887 ();
 sg13g2_decap_4 FILLER_61_2894 ();
 sg13g2_fill_1 FILLER_61_2898 ();
 sg13g2_decap_8 FILLER_61_2925 ();
 sg13g2_decap_8 FILLER_61_2932 ();
 sg13g2_decap_4 FILLER_61_2939 ();
 sg13g2_fill_2 FILLER_61_2943 ();
 sg13g2_decap_8 FILLER_61_2971 ();
 sg13g2_decap_8 FILLER_61_2978 ();
 sg13g2_decap_8 FILLER_61_2985 ();
 sg13g2_decap_8 FILLER_61_2992 ();
 sg13g2_decap_8 FILLER_61_2999 ();
 sg13g2_decap_8 FILLER_61_3006 ();
 sg13g2_fill_2 FILLER_61_3013 ();
 sg13g2_decap_8 FILLER_61_3041 ();
 sg13g2_fill_2 FILLER_61_3048 ();
 sg13g2_fill_1 FILLER_61_3050 ();
 sg13g2_decap_8 FILLER_61_3092 ();
 sg13g2_fill_1 FILLER_61_3099 ();
 sg13g2_decap_8 FILLER_61_3126 ();
 sg13g2_fill_2 FILLER_61_3133 ();
 sg13g2_decap_8 FILLER_61_3143 ();
 sg13g2_fill_2 FILLER_61_3150 ();
 sg13g2_decap_8 FILLER_61_3170 ();
 sg13g2_decap_8 FILLER_61_3177 ();
 sg13g2_decap_8 FILLER_61_3184 ();
 sg13g2_decap_8 FILLER_61_3191 ();
 sg13g2_decap_8 FILLER_61_3198 ();
 sg13g2_decap_8 FILLER_61_3205 ();
 sg13g2_decap_4 FILLER_61_3212 ();
 sg13g2_fill_1 FILLER_61_3216 ();
 sg13g2_fill_2 FILLER_61_3225 ();
 sg13g2_fill_1 FILLER_61_3227 ();
 sg13g2_decap_8 FILLER_61_3233 ();
 sg13g2_decap_8 FILLER_61_3240 ();
 sg13g2_decap_8 FILLER_61_3247 ();
 sg13g2_fill_2 FILLER_61_3254 ();
 sg13g2_fill_1 FILLER_61_3256 ();
 sg13g2_decap_4 FILLER_61_3261 ();
 sg13g2_fill_2 FILLER_61_3265 ();
 sg13g2_decap_8 FILLER_61_3293 ();
 sg13g2_decap_8 FILLER_61_3300 ();
 sg13g2_decap_8 FILLER_61_3307 ();
 sg13g2_fill_2 FILLER_61_3314 ();
 sg13g2_fill_1 FILLER_61_3316 ();
 sg13g2_decap_4 FILLER_61_3327 ();
 sg13g2_decap_8 FILLER_61_3336 ();
 sg13g2_decap_8 FILLER_61_3343 ();
 sg13g2_decap_8 FILLER_61_3350 ();
 sg13g2_fill_1 FILLER_61_3357 ();
 sg13g2_decap_4 FILLER_61_3362 ();
 sg13g2_decap_8 FILLER_61_3371 ();
 sg13g2_fill_2 FILLER_61_3378 ();
 sg13g2_decap_8 FILLER_61_3406 ();
 sg13g2_decap_4 FILLER_61_3413 ();
 sg13g2_fill_1 FILLER_61_3417 ();
 sg13g2_decap_8 FILLER_61_3451 ();
 sg13g2_fill_2 FILLER_61_3494 ();
 sg13g2_fill_1 FILLER_61_3496 ();
 sg13g2_fill_2 FILLER_61_3513 ();
 sg13g2_decap_8 FILLER_61_3541 ();
 sg13g2_decap_8 FILLER_61_3548 ();
 sg13g2_decap_8 FILLER_61_3555 ();
 sg13g2_decap_8 FILLER_61_3562 ();
 sg13g2_decap_8 FILLER_61_3569 ();
 sg13g2_decap_4 FILLER_61_3576 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_decap_8 FILLER_62_7 ();
 sg13g2_decap_8 FILLER_62_14 ();
 sg13g2_decap_8 FILLER_62_21 ();
 sg13g2_decap_8 FILLER_62_37 ();
 sg13g2_decap_8 FILLER_62_44 ();
 sg13g2_decap_8 FILLER_62_51 ();
 sg13g2_decap_8 FILLER_62_58 ();
 sg13g2_decap_8 FILLER_62_65 ();
 sg13g2_decap_8 FILLER_62_72 ();
 sg13g2_fill_1 FILLER_62_79 ();
 sg13g2_fill_1 FILLER_62_93 ();
 sg13g2_decap_4 FILLER_62_101 ();
 sg13g2_decap_8 FILLER_62_111 ();
 sg13g2_decap_8 FILLER_62_118 ();
 sg13g2_decap_8 FILLER_62_125 ();
 sg13g2_decap_8 FILLER_62_132 ();
 sg13g2_decap_8 FILLER_62_139 ();
 sg13g2_decap_4 FILLER_62_146 ();
 sg13g2_fill_1 FILLER_62_150 ();
 sg13g2_decap_4 FILLER_62_173 ();
 sg13g2_fill_1 FILLER_62_180 ();
 sg13g2_fill_1 FILLER_62_187 ();
 sg13g2_decap_4 FILLER_62_200 ();
 sg13g2_decap_4 FILLER_62_209 ();
 sg13g2_fill_2 FILLER_62_213 ();
 sg13g2_decap_4 FILLER_62_218 ();
 sg13g2_fill_1 FILLER_62_225 ();
 sg13g2_fill_1 FILLER_62_229 ();
 sg13g2_fill_2 FILLER_62_261 ();
 sg13g2_decap_8 FILLER_62_279 ();
 sg13g2_fill_2 FILLER_62_286 ();
 sg13g2_fill_2 FILLER_62_309 ();
 sg13g2_fill_1 FILLER_62_322 ();
 sg13g2_decap_8 FILLER_62_331 ();
 sg13g2_decap_8 FILLER_62_338 ();
 sg13g2_decap_8 FILLER_62_345 ();
 sg13g2_fill_1 FILLER_62_352 ();
 sg13g2_decap_8 FILLER_62_358 ();
 sg13g2_decap_8 FILLER_62_365 ();
 sg13g2_decap_8 FILLER_62_372 ();
 sg13g2_decap_8 FILLER_62_379 ();
 sg13g2_decap_8 FILLER_62_391 ();
 sg13g2_fill_2 FILLER_62_408 ();
 sg13g2_fill_2 FILLER_62_418 ();
 sg13g2_decap_8 FILLER_62_424 ();
 sg13g2_decap_8 FILLER_62_431 ();
 sg13g2_decap_4 FILLER_62_438 ();
 sg13g2_fill_2 FILLER_62_442 ();
 sg13g2_fill_1 FILLER_62_449 ();
 sg13g2_decap_4 FILLER_62_455 ();
 sg13g2_fill_2 FILLER_62_459 ();
 sg13g2_decap_8 FILLER_62_466 ();
 sg13g2_decap_8 FILLER_62_473 ();
 sg13g2_decap_8 FILLER_62_480 ();
 sg13g2_decap_8 FILLER_62_487 ();
 sg13g2_decap_4 FILLER_62_494 ();
 sg13g2_fill_2 FILLER_62_498 ();
 sg13g2_decap_8 FILLER_62_510 ();
 sg13g2_decap_8 FILLER_62_517 ();
 sg13g2_decap_8 FILLER_62_524 ();
 sg13g2_decap_8 FILLER_62_531 ();
 sg13g2_decap_8 FILLER_62_538 ();
 sg13g2_fill_1 FILLER_62_545 ();
 sg13g2_decap_8 FILLER_62_551 ();
 sg13g2_fill_1 FILLER_62_558 ();
 sg13g2_decap_8 FILLER_62_564 ();
 sg13g2_decap_8 FILLER_62_571 ();
 sg13g2_decap_8 FILLER_62_578 ();
 sg13g2_decap_8 FILLER_62_585 ();
 sg13g2_decap_8 FILLER_62_592 ();
 sg13g2_decap_8 FILLER_62_599 ();
 sg13g2_decap_4 FILLER_62_606 ();
 sg13g2_fill_1 FILLER_62_610 ();
 sg13g2_decap_8 FILLER_62_620 ();
 sg13g2_decap_8 FILLER_62_633 ();
 sg13g2_decap_8 FILLER_62_640 ();
 sg13g2_decap_8 FILLER_62_647 ();
 sg13g2_decap_8 FILLER_62_654 ();
 sg13g2_decap_4 FILLER_62_661 ();
 sg13g2_fill_1 FILLER_62_665 ();
 sg13g2_decap_4 FILLER_62_678 ();
 sg13g2_fill_1 FILLER_62_682 ();
 sg13g2_fill_2 FILLER_62_695 ();
 sg13g2_decap_4 FILLER_62_707 ();
 sg13g2_fill_1 FILLER_62_716 ();
 sg13g2_fill_2 FILLER_62_725 ();
 sg13g2_decap_8 FILLER_62_743 ();
 sg13g2_decap_8 FILLER_62_750 ();
 sg13g2_decap_4 FILLER_62_757 ();
 sg13g2_fill_1 FILLER_62_761 ();
 sg13g2_decap_8 FILLER_62_788 ();
 sg13g2_decap_8 FILLER_62_795 ();
 sg13g2_decap_8 FILLER_62_802 ();
 sg13g2_decap_8 FILLER_62_809 ();
 sg13g2_decap_8 FILLER_62_816 ();
 sg13g2_decap_8 FILLER_62_823 ();
 sg13g2_fill_2 FILLER_62_830 ();
 sg13g2_fill_1 FILLER_62_832 ();
 sg13g2_decap_8 FILLER_62_836 ();
 sg13g2_decap_8 FILLER_62_843 ();
 sg13g2_decap_8 FILLER_62_850 ();
 sg13g2_decap_8 FILLER_62_857 ();
 sg13g2_decap_8 FILLER_62_864 ();
 sg13g2_decap_4 FILLER_62_871 ();
 sg13g2_fill_1 FILLER_62_875 ();
 sg13g2_decap_8 FILLER_62_884 ();
 sg13g2_decap_8 FILLER_62_891 ();
 sg13g2_decap_8 FILLER_62_898 ();
 sg13g2_decap_4 FILLER_62_905 ();
 sg13g2_fill_1 FILLER_62_909 ();
 sg13g2_decap_8 FILLER_62_947 ();
 sg13g2_decap_8 FILLER_62_954 ();
 sg13g2_decap_8 FILLER_62_961 ();
 sg13g2_decap_4 FILLER_62_968 ();
 sg13g2_fill_2 FILLER_62_1021 ();
 sg13g2_fill_2 FILLER_62_1042 ();
 sg13g2_decap_8 FILLER_62_1061 ();
 sg13g2_decap_8 FILLER_62_1068 ();
 sg13g2_decap_4 FILLER_62_1075 ();
 sg13g2_decap_8 FILLER_62_1108 ();
 sg13g2_decap_8 FILLER_62_1115 ();
 sg13g2_decap_8 FILLER_62_1122 ();
 sg13g2_decap_8 FILLER_62_1129 ();
 sg13g2_decap_8 FILLER_62_1136 ();
 sg13g2_decap_8 FILLER_62_1143 ();
 sg13g2_decap_8 FILLER_62_1150 ();
 sg13g2_decap_8 FILLER_62_1157 ();
 sg13g2_decap_8 FILLER_62_1164 ();
 sg13g2_decap_8 FILLER_62_1171 ();
 sg13g2_decap_8 FILLER_62_1178 ();
 sg13g2_decap_8 FILLER_62_1185 ();
 sg13g2_decap_8 FILLER_62_1192 ();
 sg13g2_decap_8 FILLER_62_1199 ();
 sg13g2_decap_4 FILLER_62_1206 ();
 sg13g2_fill_1 FILLER_62_1210 ();
 sg13g2_fill_2 FILLER_62_1216 ();
 sg13g2_fill_1 FILLER_62_1218 ();
 sg13g2_decap_8 FILLER_62_1224 ();
 sg13g2_decap_8 FILLER_62_1231 ();
 sg13g2_fill_2 FILLER_62_1238 ();
 sg13g2_fill_1 FILLER_62_1240 ();
 sg13g2_fill_1 FILLER_62_1249 ();
 sg13g2_decap_4 FILLER_62_1261 ();
 sg13g2_fill_1 FILLER_62_1265 ();
 sg13g2_decap_4 FILLER_62_1283 ();
 sg13g2_fill_2 FILLER_62_1287 ();
 sg13g2_fill_1 FILLER_62_1297 ();
 sg13g2_decap_8 FILLER_62_1316 ();
 sg13g2_decap_8 FILLER_62_1323 ();
 sg13g2_decap_8 FILLER_62_1330 ();
 sg13g2_decap_8 FILLER_62_1337 ();
 sg13g2_decap_8 FILLER_62_1344 ();
 sg13g2_decap_8 FILLER_62_1351 ();
 sg13g2_decap_4 FILLER_62_1358 ();
 sg13g2_fill_1 FILLER_62_1362 ();
 sg13g2_decap_8 FILLER_62_1399 ();
 sg13g2_decap_8 FILLER_62_1406 ();
 sg13g2_decap_8 FILLER_62_1413 ();
 sg13g2_fill_2 FILLER_62_1420 ();
 sg13g2_decap_8 FILLER_62_1430 ();
 sg13g2_decap_8 FILLER_62_1445 ();
 sg13g2_decap_8 FILLER_62_1452 ();
 sg13g2_decap_8 FILLER_62_1459 ();
 sg13g2_decap_8 FILLER_62_1466 ();
 sg13g2_fill_2 FILLER_62_1473 ();
 sg13g2_decap_8 FILLER_62_1483 ();
 sg13g2_decap_8 FILLER_62_1490 ();
 sg13g2_decap_8 FILLER_62_1497 ();
 sg13g2_decap_8 FILLER_62_1504 ();
 sg13g2_fill_2 FILLER_62_1511 ();
 sg13g2_decap_8 FILLER_62_1525 ();
 sg13g2_decap_8 FILLER_62_1532 ();
 sg13g2_decap_8 FILLER_62_1539 ();
 sg13g2_decap_8 FILLER_62_1546 ();
 sg13g2_decap_8 FILLER_62_1553 ();
 sg13g2_decap_8 FILLER_62_1560 ();
 sg13g2_decap_8 FILLER_62_1567 ();
 sg13g2_decap_4 FILLER_62_1574 ();
 sg13g2_decap_4 FILLER_62_1591 ();
 sg13g2_decap_8 FILLER_62_1608 ();
 sg13g2_decap_8 FILLER_62_1615 ();
 sg13g2_decap_4 FILLER_62_1622 ();
 sg13g2_fill_2 FILLER_62_1626 ();
 sg13g2_fill_1 FILLER_62_1644 ();
 sg13g2_decap_8 FILLER_62_1649 ();
 sg13g2_decap_8 FILLER_62_1656 ();
 sg13g2_decap_8 FILLER_62_1663 ();
 sg13g2_decap_8 FILLER_62_1670 ();
 sg13g2_fill_2 FILLER_62_1677 ();
 sg13g2_fill_1 FILLER_62_1679 ();
 sg13g2_decap_8 FILLER_62_1699 ();
 sg13g2_decap_8 FILLER_62_1706 ();
 sg13g2_decap_8 FILLER_62_1749 ();
 sg13g2_decap_8 FILLER_62_1756 ();
 sg13g2_decap_8 FILLER_62_1763 ();
 sg13g2_decap_4 FILLER_62_1770 ();
 sg13g2_fill_1 FILLER_62_1774 ();
 sg13g2_decap_8 FILLER_62_1807 ();
 sg13g2_decap_8 FILLER_62_1814 ();
 sg13g2_decap_8 FILLER_62_1821 ();
 sg13g2_decap_8 FILLER_62_1828 ();
 sg13g2_decap_8 FILLER_62_1835 ();
 sg13g2_decap_4 FILLER_62_1842 ();
 sg13g2_fill_2 FILLER_62_1846 ();
 sg13g2_decap_8 FILLER_62_1865 ();
 sg13g2_decap_8 FILLER_62_1872 ();
 sg13g2_fill_1 FILLER_62_1879 ();
 sg13g2_decap_8 FILLER_62_1888 ();
 sg13g2_decap_8 FILLER_62_1895 ();
 sg13g2_fill_2 FILLER_62_1902 ();
 sg13g2_fill_1 FILLER_62_1904 ();
 sg13g2_fill_2 FILLER_62_1910 ();
 sg13g2_decap_8 FILLER_62_1922 ();
 sg13g2_decap_8 FILLER_62_1929 ();
 sg13g2_decap_8 FILLER_62_1936 ();
 sg13g2_decap_8 FILLER_62_1943 ();
 sg13g2_decap_8 FILLER_62_1950 ();
 sg13g2_decap_4 FILLER_62_1957 ();
 sg13g2_fill_1 FILLER_62_1961 ();
 sg13g2_fill_2 FILLER_62_1983 ();
 sg13g2_decap_8 FILLER_62_1989 ();
 sg13g2_decap_8 FILLER_62_1996 ();
 sg13g2_decap_8 FILLER_62_2003 ();
 sg13g2_decap_8 FILLER_62_2010 ();
 sg13g2_decap_8 FILLER_62_2017 ();
 sg13g2_decap_4 FILLER_62_2024 ();
 sg13g2_fill_1 FILLER_62_2028 ();
 sg13g2_decap_8 FILLER_62_2045 ();
 sg13g2_decap_8 FILLER_62_2052 ();
 sg13g2_decap_8 FILLER_62_2059 ();
 sg13g2_decap_8 FILLER_62_2066 ();
 sg13g2_decap_8 FILLER_62_2073 ();
 sg13g2_decap_8 FILLER_62_2080 ();
 sg13g2_decap_8 FILLER_62_2087 ();
 sg13g2_decap_8 FILLER_62_2094 ();
 sg13g2_decap_8 FILLER_62_2101 ();
 sg13g2_decap_4 FILLER_62_2108 ();
 sg13g2_fill_2 FILLER_62_2112 ();
 sg13g2_fill_1 FILLER_62_2124 ();
 sg13g2_decap_8 FILLER_62_2161 ();
 sg13g2_decap_8 FILLER_62_2168 ();
 sg13g2_decap_8 FILLER_62_2201 ();
 sg13g2_decap_8 FILLER_62_2208 ();
 sg13g2_decap_4 FILLER_62_2215 ();
 sg13g2_fill_2 FILLER_62_2219 ();
 sg13g2_decap_8 FILLER_62_2231 ();
 sg13g2_decap_8 FILLER_62_2238 ();
 sg13g2_decap_4 FILLER_62_2245 ();
 sg13g2_fill_1 FILLER_62_2249 ();
 sg13g2_decap_8 FILLER_62_2256 ();
 sg13g2_decap_8 FILLER_62_2263 ();
 sg13g2_decap_8 FILLER_62_2270 ();
 sg13g2_decap_8 FILLER_62_2277 ();
 sg13g2_decap_8 FILLER_62_2284 ();
 sg13g2_decap_8 FILLER_62_2291 ();
 sg13g2_decap_8 FILLER_62_2298 ();
 sg13g2_decap_8 FILLER_62_2305 ();
 sg13g2_decap_8 FILLER_62_2312 ();
 sg13g2_decap_8 FILLER_62_2319 ();
 sg13g2_decap_8 FILLER_62_2326 ();
 sg13g2_fill_2 FILLER_62_2333 ();
 sg13g2_fill_1 FILLER_62_2335 ();
 sg13g2_decap_8 FILLER_62_2349 ();
 sg13g2_decap_8 FILLER_62_2356 ();
 sg13g2_decap_8 FILLER_62_2363 ();
 sg13g2_decap_8 FILLER_62_2370 ();
 sg13g2_decap_8 FILLER_62_2377 ();
 sg13g2_fill_2 FILLER_62_2384 ();
 sg13g2_decap_8 FILLER_62_2412 ();
 sg13g2_decap_8 FILLER_62_2419 ();
 sg13g2_decap_8 FILLER_62_2426 ();
 sg13g2_decap_8 FILLER_62_2433 ();
 sg13g2_fill_1 FILLER_62_2440 ();
 sg13g2_decap_8 FILLER_62_2467 ();
 sg13g2_fill_2 FILLER_62_2474 ();
 sg13g2_fill_1 FILLER_62_2476 ();
 sg13g2_decap_8 FILLER_62_2503 ();
 sg13g2_decap_8 FILLER_62_2510 ();
 sg13g2_fill_2 FILLER_62_2517 ();
 sg13g2_decap_8 FILLER_62_2581 ();
 sg13g2_decap_8 FILLER_62_2588 ();
 sg13g2_decap_8 FILLER_62_2595 ();
 sg13g2_decap_8 FILLER_62_2602 ();
 sg13g2_decap_4 FILLER_62_2609 ();
 sg13g2_fill_2 FILLER_62_2613 ();
 sg13g2_decap_8 FILLER_62_2623 ();
 sg13g2_decap_8 FILLER_62_2630 ();
 sg13g2_decap_8 FILLER_62_2637 ();
 sg13g2_decap_8 FILLER_62_2644 ();
 sg13g2_decap_8 FILLER_62_2651 ();
 sg13g2_decap_8 FILLER_62_2658 ();
 sg13g2_decap_8 FILLER_62_2665 ();
 sg13g2_fill_2 FILLER_62_2672 ();
 sg13g2_decap_8 FILLER_62_2736 ();
 sg13g2_decap_8 FILLER_62_2743 ();
 sg13g2_decap_8 FILLER_62_2750 ();
 sg13g2_decap_8 FILLER_62_2757 ();
 sg13g2_decap_8 FILLER_62_2764 ();
 sg13g2_decap_8 FILLER_62_2771 ();
 sg13g2_decap_8 FILLER_62_2778 ();
 sg13g2_decap_8 FILLER_62_2785 ();
 sg13g2_decap_8 FILLER_62_2792 ();
 sg13g2_decap_8 FILLER_62_2799 ();
 sg13g2_decap_8 FILLER_62_2806 ();
 sg13g2_decap_8 FILLER_62_2813 ();
 sg13g2_decap_8 FILLER_62_2820 ();
 sg13g2_decap_8 FILLER_62_2827 ();
 sg13g2_decap_8 FILLER_62_2834 ();
 sg13g2_decap_8 FILLER_62_2841 ();
 sg13g2_decap_8 FILLER_62_2848 ();
 sg13g2_decap_8 FILLER_62_2855 ();
 sg13g2_decap_8 FILLER_62_2862 ();
 sg13g2_decap_8 FILLER_62_2869 ();
 sg13g2_decap_8 FILLER_62_2876 ();
 sg13g2_decap_8 FILLER_62_2883 ();
 sg13g2_decap_8 FILLER_62_2890 ();
 sg13g2_decap_8 FILLER_62_2897 ();
 sg13g2_decap_8 FILLER_62_2904 ();
 sg13g2_decap_8 FILLER_62_2911 ();
 sg13g2_decap_8 FILLER_62_2918 ();
 sg13g2_decap_8 FILLER_62_2925 ();
 sg13g2_decap_8 FILLER_62_2932 ();
 sg13g2_decap_8 FILLER_62_2939 ();
 sg13g2_decap_8 FILLER_62_2946 ();
 sg13g2_decap_8 FILLER_62_2953 ();
 sg13g2_decap_8 FILLER_62_2960 ();
 sg13g2_fill_1 FILLER_62_2967 ();
 sg13g2_decap_8 FILLER_62_3004 ();
 sg13g2_decap_8 FILLER_62_3011 ();
 sg13g2_decap_8 FILLER_62_3018 ();
 sg13g2_decap_8 FILLER_62_3025 ();
 sg13g2_decap_8 FILLER_62_3032 ();
 sg13g2_decap_8 FILLER_62_3039 ();
 sg13g2_decap_8 FILLER_62_3046 ();
 sg13g2_decap_8 FILLER_62_3053 ();
 sg13g2_decap_4 FILLER_62_3060 ();
 sg13g2_fill_2 FILLER_62_3064 ();
 sg13g2_decap_8 FILLER_62_3076 ();
 sg13g2_decap_8 FILLER_62_3083 ();
 sg13g2_decap_8 FILLER_62_3090 ();
 sg13g2_decap_8 FILLER_62_3097 ();
 sg13g2_fill_2 FILLER_62_3104 ();
 sg13g2_fill_1 FILLER_62_3106 ();
 sg13g2_decap_8 FILLER_62_3116 ();
 sg13g2_decap_8 FILLER_62_3123 ();
 sg13g2_decap_8 FILLER_62_3130 ();
 sg13g2_decap_8 FILLER_62_3137 ();
 sg13g2_decap_8 FILLER_62_3144 ();
 sg13g2_decap_8 FILLER_62_3151 ();
 sg13g2_fill_2 FILLER_62_3158 ();
 sg13g2_fill_1 FILLER_62_3160 ();
 sg13g2_decap_4 FILLER_62_3207 ();
 sg13g2_fill_1 FILLER_62_3211 ();
 sg13g2_decap_8 FILLER_62_3248 ();
 sg13g2_decap_8 FILLER_62_3265 ();
 sg13g2_decap_8 FILLER_62_3272 ();
 sg13g2_fill_2 FILLER_62_3279 ();
 sg13g2_decap_8 FILLER_62_3286 ();
 sg13g2_decap_8 FILLER_62_3293 ();
 sg13g2_decap_8 FILLER_62_3300 ();
 sg13g2_decap_8 FILLER_62_3307 ();
 sg13g2_decap_8 FILLER_62_3324 ();
 sg13g2_fill_1 FILLER_62_3331 ();
 sg13g2_decap_8 FILLER_62_3358 ();
 sg13g2_decap_8 FILLER_62_3365 ();
 sg13g2_decap_8 FILLER_62_3408 ();
 sg13g2_decap_8 FILLER_62_3415 ();
 sg13g2_decap_8 FILLER_62_3422 ();
 sg13g2_fill_2 FILLER_62_3434 ();
 sg13g2_fill_1 FILLER_62_3436 ();
 sg13g2_decap_8 FILLER_62_3485 ();
 sg13g2_decap_8 FILLER_62_3492 ();
 sg13g2_decap_8 FILLER_62_3499 ();
 sg13g2_decap_8 FILLER_62_3506 ();
 sg13g2_decap_8 FILLER_62_3513 ();
 sg13g2_fill_2 FILLER_62_3520 ();
 sg13g2_fill_1 FILLER_62_3522 ();
 sg13g2_decap_8 FILLER_62_3531 ();
 sg13g2_decap_8 FILLER_62_3538 ();
 sg13g2_decap_8 FILLER_62_3545 ();
 sg13g2_decap_8 FILLER_62_3552 ();
 sg13g2_decap_8 FILLER_62_3559 ();
 sg13g2_decap_8 FILLER_62_3566 ();
 sg13g2_decap_8 FILLER_62_3573 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_decap_8 FILLER_63_7 ();
 sg13g2_decap_8 FILLER_63_14 ();
 sg13g2_fill_1 FILLER_63_21 ();
 sg13g2_decap_4 FILLER_63_31 ();
 sg13g2_decap_8 FILLER_63_44 ();
 sg13g2_decap_8 FILLER_63_51 ();
 sg13g2_decap_8 FILLER_63_58 ();
 sg13g2_decap_8 FILLER_63_65 ();
 sg13g2_decap_8 FILLER_63_72 ();
 sg13g2_decap_8 FILLER_63_79 ();
 sg13g2_decap_4 FILLER_63_86 ();
 sg13g2_fill_2 FILLER_63_95 ();
 sg13g2_fill_1 FILLER_63_97 ();
 sg13g2_decap_8 FILLER_63_103 ();
 sg13g2_decap_8 FILLER_63_116 ();
 sg13g2_decap_8 FILLER_63_123 ();
 sg13g2_decap_8 FILLER_63_130 ();
 sg13g2_decap_8 FILLER_63_137 ();
 sg13g2_fill_2 FILLER_63_144 ();
 sg13g2_fill_2 FILLER_63_190 ();
 sg13g2_fill_1 FILLER_63_225 ();
 sg13g2_fill_1 FILLER_63_236 ();
 sg13g2_fill_1 FILLER_63_312 ();
 sg13g2_fill_1 FILLER_63_328 ();
 sg13g2_decap_8 FILLER_63_347 ();
 sg13g2_decap_8 FILLER_63_354 ();
 sg13g2_decap_8 FILLER_63_361 ();
 sg13g2_decap_8 FILLER_63_373 ();
 sg13g2_decap_4 FILLER_63_380 ();
 sg13g2_fill_2 FILLER_63_384 ();
 sg13g2_fill_1 FILLER_63_394 ();
 sg13g2_decap_4 FILLER_63_403 ();
 sg13g2_fill_1 FILLER_63_421 ();
 sg13g2_fill_1 FILLER_63_442 ();
 sg13g2_fill_1 FILLER_63_458 ();
 sg13g2_fill_1 FILLER_63_466 ();
 sg13g2_decap_8 FILLER_63_479 ();
 sg13g2_decap_8 FILLER_63_486 ();
 sg13g2_decap_8 FILLER_63_493 ();
 sg13g2_decap_4 FILLER_63_500 ();
 sg13g2_fill_2 FILLER_63_512 ();
 sg13g2_fill_2 FILLER_63_519 ();
 sg13g2_decap_8 FILLER_63_525 ();
 sg13g2_decap_8 FILLER_63_532 ();
 sg13g2_decap_4 FILLER_63_539 ();
 sg13g2_fill_1 FILLER_63_543 ();
 sg13g2_decap_8 FILLER_63_552 ();
 sg13g2_decap_8 FILLER_63_559 ();
 sg13g2_decap_8 FILLER_63_566 ();
 sg13g2_decap_8 FILLER_63_573 ();
 sg13g2_decap_8 FILLER_63_580 ();
 sg13g2_fill_2 FILLER_63_587 ();
 sg13g2_fill_1 FILLER_63_589 ();
 sg13g2_fill_2 FILLER_63_598 ();
 sg13g2_decap_8 FILLER_63_609 ();
 sg13g2_decap_8 FILLER_63_616 ();
 sg13g2_decap_8 FILLER_63_623 ();
 sg13g2_decap_4 FILLER_63_630 ();
 sg13g2_decap_8 FILLER_63_644 ();
 sg13g2_decap_8 FILLER_63_651 ();
 sg13g2_decap_8 FILLER_63_658 ();
 sg13g2_decap_8 FILLER_63_665 ();
 sg13g2_decap_8 FILLER_63_672 ();
 sg13g2_fill_1 FILLER_63_679 ();
 sg13g2_fill_2 FILLER_63_689 ();
 sg13g2_fill_1 FILLER_63_691 ();
 sg13g2_decap_8 FILLER_63_697 ();
 sg13g2_decap_8 FILLER_63_704 ();
 sg13g2_decap_8 FILLER_63_711 ();
 sg13g2_decap_8 FILLER_63_718 ();
 sg13g2_decap_8 FILLER_63_725 ();
 sg13g2_decap_4 FILLER_63_738 ();
 sg13g2_fill_2 FILLER_63_742 ();
 sg13g2_fill_2 FILLER_63_758 ();
 sg13g2_fill_1 FILLER_63_760 ();
 sg13g2_decap_8 FILLER_63_770 ();
 sg13g2_decap_8 FILLER_63_777 ();
 sg13g2_decap_8 FILLER_63_784 ();
 sg13g2_decap_8 FILLER_63_791 ();
 sg13g2_decap_4 FILLER_63_798 ();
 sg13g2_fill_1 FILLER_63_802 ();
 sg13g2_decap_8 FILLER_63_811 ();
 sg13g2_fill_2 FILLER_63_818 ();
 sg13g2_decap_8 FILLER_63_834 ();
 sg13g2_decap_8 FILLER_63_841 ();
 sg13g2_decap_8 FILLER_63_848 ();
 sg13g2_decap_4 FILLER_63_855 ();
 sg13g2_fill_1 FILLER_63_859 ();
 sg13g2_decap_4 FILLER_63_872 ();
 sg13g2_decap_8 FILLER_63_896 ();
 sg13g2_decap_8 FILLER_63_903 ();
 sg13g2_decap_4 FILLER_63_910 ();
 sg13g2_fill_1 FILLER_63_914 ();
 sg13g2_decap_8 FILLER_63_936 ();
 sg13g2_decap_8 FILLER_63_943 ();
 sg13g2_decap_8 FILLER_63_950 ();
 sg13g2_decap_8 FILLER_63_957 ();
 sg13g2_decap_4 FILLER_63_964 ();
 sg13g2_fill_1 FILLER_63_968 ();
 sg13g2_decap_4 FILLER_63_1010 ();
 sg13g2_decap_8 FILLER_63_1053 ();
 sg13g2_decap_8 FILLER_63_1060 ();
 sg13g2_decap_8 FILLER_63_1067 ();
 sg13g2_decap_8 FILLER_63_1074 ();
 sg13g2_decap_8 FILLER_63_1081 ();
 sg13g2_fill_2 FILLER_63_1088 ();
 sg13g2_decap_8 FILLER_63_1113 ();
 sg13g2_decap_8 FILLER_63_1120 ();
 sg13g2_decap_8 FILLER_63_1127 ();
 sg13g2_decap_8 FILLER_63_1134 ();
 sg13g2_decap_8 FILLER_63_1141 ();
 sg13g2_decap_8 FILLER_63_1148 ();
 sg13g2_decap_8 FILLER_63_1155 ();
 sg13g2_decap_8 FILLER_63_1162 ();
 sg13g2_decap_8 FILLER_63_1169 ();
 sg13g2_decap_8 FILLER_63_1176 ();
 sg13g2_decap_8 FILLER_63_1183 ();
 sg13g2_decap_8 FILLER_63_1190 ();
 sg13g2_fill_2 FILLER_63_1197 ();
 sg13g2_fill_2 FILLER_63_1207 ();
 sg13g2_decap_4 FILLER_63_1229 ();
 sg13g2_fill_2 FILLER_63_1233 ();
 sg13g2_decap_8 FILLER_63_1238 ();
 sg13g2_decap_8 FILLER_63_1245 ();
 sg13g2_decap_8 FILLER_63_1252 ();
 sg13g2_fill_2 FILLER_63_1294 ();
 sg13g2_decap_8 FILLER_63_1330 ();
 sg13g2_decap_8 FILLER_63_1337 ();
 sg13g2_fill_2 FILLER_63_1344 ();
 sg13g2_fill_2 FILLER_63_1349 ();
 sg13g2_fill_1 FILLER_63_1354 ();
 sg13g2_decap_4 FILLER_63_1361 ();
 sg13g2_fill_2 FILLER_63_1365 ();
 sg13g2_decap_8 FILLER_63_1403 ();
 sg13g2_decap_8 FILLER_63_1410 ();
 sg13g2_decap_4 FILLER_63_1417 ();
 sg13g2_decap_4 FILLER_63_1434 ();
 sg13g2_fill_2 FILLER_63_1438 ();
 sg13g2_decap_8 FILLER_63_1450 ();
 sg13g2_decap_8 FILLER_63_1457 ();
 sg13g2_decap_8 FILLER_63_1464 ();
 sg13g2_decap_8 FILLER_63_1471 ();
 sg13g2_decap_8 FILLER_63_1478 ();
 sg13g2_decap_8 FILLER_63_1485 ();
 sg13g2_decap_8 FILLER_63_1492 ();
 sg13g2_decap_8 FILLER_63_1499 ();
 sg13g2_decap_8 FILLER_63_1506 ();
 sg13g2_decap_8 FILLER_63_1513 ();
 sg13g2_decap_8 FILLER_63_1520 ();
 sg13g2_decap_8 FILLER_63_1527 ();
 sg13g2_decap_8 FILLER_63_1534 ();
 sg13g2_decap_8 FILLER_63_1541 ();
 sg13g2_decap_8 FILLER_63_1548 ();
 sg13g2_decap_8 FILLER_63_1555 ();
 sg13g2_decap_8 FILLER_63_1562 ();
 sg13g2_fill_2 FILLER_63_1569 ();
 sg13g2_fill_1 FILLER_63_1571 ();
 sg13g2_decap_4 FILLER_63_1600 ();
 sg13g2_fill_2 FILLER_63_1620 ();
 sg13g2_fill_1 FILLER_63_1622 ();
 sg13g2_decap_8 FILLER_63_1631 ();
 sg13g2_fill_1 FILLER_63_1638 ();
 sg13g2_decap_8 FILLER_63_1647 ();
 sg13g2_decap_4 FILLER_63_1654 ();
 sg13g2_fill_2 FILLER_63_1658 ();
 sg13g2_decap_8 FILLER_63_1668 ();
 sg13g2_decap_8 FILLER_63_1675 ();
 sg13g2_decap_8 FILLER_63_1682 ();
 sg13g2_decap_8 FILLER_63_1689 ();
 sg13g2_decap_8 FILLER_63_1696 ();
 sg13g2_decap_8 FILLER_63_1703 ();
 sg13g2_decap_4 FILLER_63_1710 ();
 sg13g2_fill_1 FILLER_63_1714 ();
 sg13g2_decap_8 FILLER_63_1751 ();
 sg13g2_decap_8 FILLER_63_1758 ();
 sg13g2_decap_8 FILLER_63_1765 ();
 sg13g2_decap_8 FILLER_63_1772 ();
 sg13g2_decap_4 FILLER_63_1779 ();
 sg13g2_fill_1 FILLER_63_1783 ();
 sg13g2_decap_8 FILLER_63_1795 ();
 sg13g2_decap_8 FILLER_63_1802 ();
 sg13g2_decap_8 FILLER_63_1809 ();
 sg13g2_decap_8 FILLER_63_1816 ();
 sg13g2_decap_8 FILLER_63_1823 ();
 sg13g2_decap_8 FILLER_63_1830 ();
 sg13g2_decap_4 FILLER_63_1837 ();
 sg13g2_fill_2 FILLER_63_1841 ();
 sg13g2_decap_8 FILLER_63_1851 ();
 sg13g2_decap_8 FILLER_63_1858 ();
 sg13g2_decap_8 FILLER_63_1865 ();
 sg13g2_decap_8 FILLER_63_1887 ();
 sg13g2_decap_8 FILLER_63_1894 ();
 sg13g2_fill_1 FILLER_63_1901 ();
 sg13g2_decap_4 FILLER_63_1930 ();
 sg13g2_fill_2 FILLER_63_1934 ();
 sg13g2_decap_8 FILLER_63_1965 ();
 sg13g2_decap_4 FILLER_63_1972 ();
 sg13g2_fill_2 FILLER_63_1976 ();
 sg13g2_decap_8 FILLER_63_1993 ();
 sg13g2_decap_8 FILLER_63_2000 ();
 sg13g2_decap_8 FILLER_63_2007 ();
 sg13g2_decap_8 FILLER_63_2014 ();
 sg13g2_decap_8 FILLER_63_2021 ();
 sg13g2_decap_8 FILLER_63_2036 ();
 sg13g2_decap_8 FILLER_63_2043 ();
 sg13g2_decap_8 FILLER_63_2050 ();
 sg13g2_decap_8 FILLER_63_2057 ();
 sg13g2_decap_8 FILLER_63_2064 ();
 sg13g2_fill_1 FILLER_63_2071 ();
 sg13g2_decap_8 FILLER_63_2108 ();
 sg13g2_decap_8 FILLER_63_2115 ();
 sg13g2_decap_4 FILLER_63_2122 ();
 sg13g2_fill_2 FILLER_63_2126 ();
 sg13g2_decap_8 FILLER_63_2154 ();
 sg13g2_decap_8 FILLER_63_2161 ();
 sg13g2_decap_8 FILLER_63_2168 ();
 sg13g2_decap_4 FILLER_63_2175 ();
 sg13g2_decap_8 FILLER_63_2189 ();
 sg13g2_decap_8 FILLER_63_2196 ();
 sg13g2_decap_8 FILLER_63_2203 ();
 sg13g2_decap_8 FILLER_63_2210 ();
 sg13g2_decap_4 FILLER_63_2217 ();
 sg13g2_fill_2 FILLER_63_2221 ();
 sg13g2_decap_8 FILLER_63_2243 ();
 sg13g2_decap_8 FILLER_63_2250 ();
 sg13g2_decap_8 FILLER_63_2257 ();
 sg13g2_fill_2 FILLER_63_2264 ();
 sg13g2_decap_8 FILLER_63_2276 ();
 sg13g2_decap_8 FILLER_63_2309 ();
 sg13g2_decap_8 FILLER_63_2316 ();
 sg13g2_decap_4 FILLER_63_2323 ();
 sg13g2_decap_8 FILLER_63_2363 ();
 sg13g2_decap_4 FILLER_63_2370 ();
 sg13g2_fill_2 FILLER_63_2374 ();
 sg13g2_decap_8 FILLER_63_2412 ();
 sg13g2_decap_8 FILLER_63_2419 ();
 sg13g2_decap_8 FILLER_63_2426 ();
 sg13g2_decap_4 FILLER_63_2433 ();
 sg13g2_fill_2 FILLER_63_2437 ();
 sg13g2_decap_8 FILLER_63_2465 ();
 sg13g2_decap_8 FILLER_63_2472 ();
 sg13g2_fill_2 FILLER_63_2479 ();
 sg13g2_fill_1 FILLER_63_2481 ();
 sg13g2_decap_8 FILLER_63_2492 ();
 sg13g2_decap_8 FILLER_63_2499 ();
 sg13g2_decap_8 FILLER_63_2506 ();
 sg13g2_decap_8 FILLER_63_2513 ();
 sg13g2_decap_8 FILLER_63_2520 ();
 sg13g2_decap_8 FILLER_63_2527 ();
 sg13g2_decap_8 FILLER_63_2534 ();
 sg13g2_fill_2 FILLER_63_2541 ();
 sg13g2_fill_1 FILLER_63_2543 ();
 sg13g2_decap_8 FILLER_63_2563 ();
 sg13g2_decap_8 FILLER_63_2570 ();
 sg13g2_decap_8 FILLER_63_2577 ();
 sg13g2_decap_8 FILLER_63_2584 ();
 sg13g2_fill_1 FILLER_63_2591 ();
 sg13g2_decap_8 FILLER_63_2602 ();
 sg13g2_decap_8 FILLER_63_2609 ();
 sg13g2_decap_8 FILLER_63_2616 ();
 sg13g2_decap_8 FILLER_63_2623 ();
 sg13g2_decap_8 FILLER_63_2630 ();
 sg13g2_decap_8 FILLER_63_2637 ();
 sg13g2_decap_8 FILLER_63_2644 ();
 sg13g2_fill_2 FILLER_63_2651 ();
 sg13g2_decap_8 FILLER_63_2661 ();
 sg13g2_decap_8 FILLER_63_2668 ();
 sg13g2_decap_8 FILLER_63_2675 ();
 sg13g2_decap_8 FILLER_63_2682 ();
 sg13g2_decap_8 FILLER_63_2689 ();
 sg13g2_decap_8 FILLER_63_2696 ();
 sg13g2_decap_8 FILLER_63_2703 ();
 sg13g2_decap_8 FILLER_63_2710 ();
 sg13g2_decap_8 FILLER_63_2717 ();
 sg13g2_decap_8 FILLER_63_2724 ();
 sg13g2_decap_8 FILLER_63_2731 ();
 sg13g2_decap_8 FILLER_63_2738 ();
 sg13g2_fill_1 FILLER_63_2745 ();
 sg13g2_decap_8 FILLER_63_2782 ();
 sg13g2_decap_8 FILLER_63_2789 ();
 sg13g2_decap_8 FILLER_63_2796 ();
 sg13g2_decap_8 FILLER_63_2803 ();
 sg13g2_decap_8 FILLER_63_2810 ();
 sg13g2_decap_8 FILLER_63_2817 ();
 sg13g2_decap_8 FILLER_63_2824 ();
 sg13g2_decap_8 FILLER_63_2831 ();
 sg13g2_decap_8 FILLER_63_2838 ();
 sg13g2_decap_8 FILLER_63_2855 ();
 sg13g2_decap_8 FILLER_63_2862 ();
 sg13g2_decap_8 FILLER_63_2869 ();
 sg13g2_decap_8 FILLER_63_2876 ();
 sg13g2_decap_8 FILLER_63_2883 ();
 sg13g2_decap_8 FILLER_63_2890 ();
 sg13g2_decap_8 FILLER_63_2897 ();
 sg13g2_decap_8 FILLER_63_2904 ();
 sg13g2_decap_8 FILLER_63_2911 ();
 sg13g2_decap_8 FILLER_63_2918 ();
 sg13g2_decap_8 FILLER_63_2925 ();
 sg13g2_decap_8 FILLER_63_2932 ();
 sg13g2_decap_8 FILLER_63_2939 ();
 sg13g2_decap_8 FILLER_63_2946 ();
 sg13g2_decap_8 FILLER_63_2953 ();
 sg13g2_decap_4 FILLER_63_2960 ();
 sg13g2_fill_1 FILLER_63_2964 ();
 sg13g2_decap_8 FILLER_63_2976 ();
 sg13g2_decap_8 FILLER_63_2983 ();
 sg13g2_decap_8 FILLER_63_2990 ();
 sg13g2_fill_2 FILLER_63_2997 ();
 sg13g2_decap_8 FILLER_63_3009 ();
 sg13g2_decap_8 FILLER_63_3016 ();
 sg13g2_decap_8 FILLER_63_3023 ();
 sg13g2_decap_8 FILLER_63_3030 ();
 sg13g2_decap_8 FILLER_63_3037 ();
 sg13g2_decap_8 FILLER_63_3044 ();
 sg13g2_decap_8 FILLER_63_3051 ();
 sg13g2_decap_8 FILLER_63_3058 ();
 sg13g2_decap_8 FILLER_63_3065 ();
 sg13g2_decap_8 FILLER_63_3072 ();
 sg13g2_decap_8 FILLER_63_3079 ();
 sg13g2_decap_8 FILLER_63_3086 ();
 sg13g2_decap_8 FILLER_63_3093 ();
 sg13g2_decap_8 FILLER_63_3100 ();
 sg13g2_fill_2 FILLER_63_3107 ();
 sg13g2_decap_8 FILLER_63_3115 ();
 sg13g2_decap_8 FILLER_63_3122 ();
 sg13g2_decap_8 FILLER_63_3129 ();
 sg13g2_decap_8 FILLER_63_3136 ();
 sg13g2_decap_8 FILLER_63_3143 ();
 sg13g2_decap_4 FILLER_63_3150 ();
 sg13g2_decap_8 FILLER_63_3159 ();
 sg13g2_decap_8 FILLER_63_3166 ();
 sg13g2_decap_8 FILLER_63_3173 ();
 sg13g2_decap_4 FILLER_63_3180 ();
 sg13g2_fill_1 FILLER_63_3184 ();
 sg13g2_decap_8 FILLER_63_3211 ();
 sg13g2_decap_8 FILLER_63_3218 ();
 sg13g2_decap_8 FILLER_63_3225 ();
 sg13g2_decap_8 FILLER_63_3232 ();
 sg13g2_decap_8 FILLER_63_3239 ();
 sg13g2_decap_4 FILLER_63_3246 ();
 sg13g2_fill_1 FILLER_63_3250 ();
 sg13g2_decap_8 FILLER_63_3277 ();
 sg13g2_decap_8 FILLER_63_3284 ();
 sg13g2_decap_8 FILLER_63_3291 ();
 sg13g2_fill_1 FILLER_63_3298 ();
 sg13g2_decap_8 FILLER_63_3361 ();
 sg13g2_fill_2 FILLER_63_3368 ();
 sg13g2_fill_1 FILLER_63_3370 ();
 sg13g2_decap_8 FILLER_63_3407 ();
 sg13g2_decap_8 FILLER_63_3414 ();
 sg13g2_decap_8 FILLER_63_3421 ();
 sg13g2_decap_8 FILLER_63_3428 ();
 sg13g2_decap_8 FILLER_63_3435 ();
 sg13g2_decap_4 FILLER_63_3442 ();
 sg13g2_decap_8 FILLER_63_3482 ();
 sg13g2_decap_8 FILLER_63_3489 ();
 sg13g2_decap_8 FILLER_63_3496 ();
 sg13g2_fill_2 FILLER_63_3503 ();
 sg13g2_decap_8 FILLER_63_3531 ();
 sg13g2_decap_8 FILLER_63_3538 ();
 sg13g2_decap_8 FILLER_63_3545 ();
 sg13g2_decap_8 FILLER_63_3552 ();
 sg13g2_decap_8 FILLER_63_3559 ();
 sg13g2_decap_8 FILLER_63_3566 ();
 sg13g2_decap_8 FILLER_63_3573 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_8 FILLER_64_7 ();
 sg13g2_decap_8 FILLER_64_48 ();
 sg13g2_decap_8 FILLER_64_55 ();
 sg13g2_decap_8 FILLER_64_62 ();
 sg13g2_decap_8 FILLER_64_69 ();
 sg13g2_fill_2 FILLER_64_76 ();
 sg13g2_fill_1 FILLER_64_78 ();
 sg13g2_fill_1 FILLER_64_94 ();
 sg13g2_decap_8 FILLER_64_100 ();
 sg13g2_decap_8 FILLER_64_107 ();
 sg13g2_decap_8 FILLER_64_114 ();
 sg13g2_fill_2 FILLER_64_121 ();
 sg13g2_decap_8 FILLER_64_132 ();
 sg13g2_decap_8 FILLER_64_139 ();
 sg13g2_decap_8 FILLER_64_146 ();
 sg13g2_fill_2 FILLER_64_153 ();
 sg13g2_fill_1 FILLER_64_155 ();
 sg13g2_fill_1 FILLER_64_161 ();
 sg13g2_decap_8 FILLER_64_180 ();
 sg13g2_decap_8 FILLER_64_187 ();
 sg13g2_decap_8 FILLER_64_194 ();
 sg13g2_fill_2 FILLER_64_201 ();
 sg13g2_fill_2 FILLER_64_207 ();
 sg13g2_fill_1 FILLER_64_214 ();
 sg13g2_fill_2 FILLER_64_218 ();
 sg13g2_fill_1 FILLER_64_220 ();
 sg13g2_fill_1 FILLER_64_241 ();
 sg13g2_fill_2 FILLER_64_260 ();
 sg13g2_fill_1 FILLER_64_268 ();
 sg13g2_fill_1 FILLER_64_316 ();
 sg13g2_fill_1 FILLER_64_329 ();
 sg13g2_decap_4 FILLER_64_340 ();
 sg13g2_decap_8 FILLER_64_354 ();
 sg13g2_decap_8 FILLER_64_361 ();
 sg13g2_decap_8 FILLER_64_368 ();
 sg13g2_fill_2 FILLER_64_382 ();
 sg13g2_decap_4 FILLER_64_409 ();
 sg13g2_fill_1 FILLER_64_413 ();
 sg13g2_fill_1 FILLER_64_435 ();
 sg13g2_fill_2 FILLER_64_444 ();
 sg13g2_decap_8 FILLER_64_454 ();
 sg13g2_decap_8 FILLER_64_466 ();
 sg13g2_decap_8 FILLER_64_473 ();
 sg13g2_decap_8 FILLER_64_480 ();
 sg13g2_decap_8 FILLER_64_487 ();
 sg13g2_decap_8 FILLER_64_494 ();
 sg13g2_fill_1 FILLER_64_501 ();
 sg13g2_decap_8 FILLER_64_531 ();
 sg13g2_decap_4 FILLER_64_538 ();
 sg13g2_fill_1 FILLER_64_542 ();
 sg13g2_decap_8 FILLER_64_547 ();
 sg13g2_decap_8 FILLER_64_554 ();
 sg13g2_decap_8 FILLER_64_561 ();
 sg13g2_decap_8 FILLER_64_568 ();
 sg13g2_decap_4 FILLER_64_575 ();
 sg13g2_fill_2 FILLER_64_610 ();
 sg13g2_fill_1 FILLER_64_612 ();
 sg13g2_decap_4 FILLER_64_628 ();
 sg13g2_fill_1 FILLER_64_632 ();
 sg13g2_decap_8 FILLER_64_640 ();
 sg13g2_decap_8 FILLER_64_647 ();
 sg13g2_fill_1 FILLER_64_654 ();
 sg13g2_decap_8 FILLER_64_658 ();
 sg13g2_fill_2 FILLER_64_665 ();
 sg13g2_fill_1 FILLER_64_667 ();
 sg13g2_decap_8 FILLER_64_708 ();
 sg13g2_decap_8 FILLER_64_715 ();
 sg13g2_decap_8 FILLER_64_722 ();
 sg13g2_fill_2 FILLER_64_729 ();
 sg13g2_fill_2 FILLER_64_740 ();
 sg13g2_decap_8 FILLER_64_768 ();
 sg13g2_decap_8 FILLER_64_775 ();
 sg13g2_decap_8 FILLER_64_782 ();
 sg13g2_fill_2 FILLER_64_789 ();
 sg13g2_fill_1 FILLER_64_791 ();
 sg13g2_decap_8 FILLER_64_816 ();
 sg13g2_decap_8 FILLER_64_823 ();
 sg13g2_decap_8 FILLER_64_830 ();
 sg13g2_decap_8 FILLER_64_837 ();
 sg13g2_decap_8 FILLER_64_844 ();
 sg13g2_decap_4 FILLER_64_851 ();
 sg13g2_fill_2 FILLER_64_855 ();
 sg13g2_fill_1 FILLER_64_871 ();
 sg13g2_decap_4 FILLER_64_878 ();
 sg13g2_decap_8 FILLER_64_895 ();
 sg13g2_decap_8 FILLER_64_902 ();
 sg13g2_decap_8 FILLER_64_909 ();
 sg13g2_decap_8 FILLER_64_916 ();
 sg13g2_fill_2 FILLER_64_923 ();
 sg13g2_decap_8 FILLER_64_930 ();
 sg13g2_decap_8 FILLER_64_937 ();
 sg13g2_decap_8 FILLER_64_944 ();
 sg13g2_decap_8 FILLER_64_951 ();
 sg13g2_decap_8 FILLER_64_958 ();
 sg13g2_decap_8 FILLER_64_965 ();
 sg13g2_fill_2 FILLER_64_972 ();
 sg13g2_fill_1 FILLER_64_974 ();
 sg13g2_fill_1 FILLER_64_998 ();
 sg13g2_decap_8 FILLER_64_1004 ();
 sg13g2_decap_8 FILLER_64_1011 ();
 sg13g2_decap_8 FILLER_64_1018 ();
 sg13g2_decap_4 FILLER_64_1025 ();
 sg13g2_fill_1 FILLER_64_1029 ();
 sg13g2_fill_1 FILLER_64_1040 ();
 sg13g2_fill_2 FILLER_64_1044 ();
 sg13g2_decap_8 FILLER_64_1054 ();
 sg13g2_decap_8 FILLER_64_1061 ();
 sg13g2_decap_8 FILLER_64_1068 ();
 sg13g2_decap_8 FILLER_64_1075 ();
 sg13g2_decap_8 FILLER_64_1082 ();
 sg13g2_decap_4 FILLER_64_1089 ();
 sg13g2_fill_1 FILLER_64_1093 ();
 sg13g2_decap_8 FILLER_64_1111 ();
 sg13g2_decap_8 FILLER_64_1118 ();
 sg13g2_decap_8 FILLER_64_1125 ();
 sg13g2_decap_8 FILLER_64_1132 ();
 sg13g2_decap_8 FILLER_64_1139 ();
 sg13g2_decap_8 FILLER_64_1146 ();
 sg13g2_decap_4 FILLER_64_1153 ();
 sg13g2_fill_1 FILLER_64_1157 ();
 sg13g2_decap_4 FILLER_64_1162 ();
 sg13g2_fill_2 FILLER_64_1166 ();
 sg13g2_fill_1 FILLER_64_1182 ();
 sg13g2_decap_8 FILLER_64_1193 ();
 sg13g2_decap_8 FILLER_64_1200 ();
 sg13g2_fill_2 FILLER_64_1207 ();
 sg13g2_fill_1 FILLER_64_1209 ();
 sg13g2_decap_8 FILLER_64_1215 ();
 sg13g2_decap_8 FILLER_64_1222 ();
 sg13g2_decap_4 FILLER_64_1229 ();
 sg13g2_fill_2 FILLER_64_1233 ();
 sg13g2_decap_8 FILLER_64_1238 ();
 sg13g2_decap_8 FILLER_64_1245 ();
 sg13g2_decap_8 FILLER_64_1252 ();
 sg13g2_decap_8 FILLER_64_1259 ();
 sg13g2_decap_8 FILLER_64_1266 ();
 sg13g2_decap_8 FILLER_64_1273 ();
 sg13g2_decap_8 FILLER_64_1280 ();
 sg13g2_decap_8 FILLER_64_1287 ();
 sg13g2_decap_8 FILLER_64_1294 ();
 sg13g2_decap_8 FILLER_64_1301 ();
 sg13g2_fill_2 FILLER_64_1308 ();
 sg13g2_fill_1 FILLER_64_1310 ();
 sg13g2_decap_8 FILLER_64_1323 ();
 sg13g2_fill_1 FILLER_64_1330 ();
 sg13g2_fill_2 FILLER_64_1341 ();
 sg13g2_decap_8 FILLER_64_1391 ();
 sg13g2_decap_8 FILLER_64_1398 ();
 sg13g2_decap_8 FILLER_64_1405 ();
 sg13g2_decap_8 FILLER_64_1412 ();
 sg13g2_decap_8 FILLER_64_1419 ();
 sg13g2_fill_2 FILLER_64_1426 ();
 sg13g2_fill_1 FILLER_64_1428 ();
 sg13g2_decap_8 FILLER_64_1437 ();
 sg13g2_decap_8 FILLER_64_1444 ();
 sg13g2_fill_1 FILLER_64_1451 ();
 sg13g2_decap_8 FILLER_64_1478 ();
 sg13g2_decap_8 FILLER_64_1485 ();
 sg13g2_decap_8 FILLER_64_1492 ();
 sg13g2_decap_8 FILLER_64_1499 ();
 sg13g2_decap_8 FILLER_64_1506 ();
 sg13g2_fill_2 FILLER_64_1513 ();
 sg13g2_decap_8 FILLER_64_1525 ();
 sg13g2_decap_4 FILLER_64_1532 ();
 sg13g2_fill_2 FILLER_64_1536 ();
 sg13g2_decap_8 FILLER_64_1546 ();
 sg13g2_decap_8 FILLER_64_1553 ();
 sg13g2_decap_8 FILLER_64_1560 ();
 sg13g2_decap_8 FILLER_64_1567 ();
 sg13g2_decap_8 FILLER_64_1574 ();
 sg13g2_decap_8 FILLER_64_1581 ();
 sg13g2_decap_4 FILLER_64_1588 ();
 sg13g2_decap_8 FILLER_64_1600 ();
 sg13g2_decap_8 FILLER_64_1607 ();
 sg13g2_decap_8 FILLER_64_1614 ();
 sg13g2_decap_8 FILLER_64_1621 ();
 sg13g2_decap_8 FILLER_64_1628 ();
 sg13g2_decap_8 FILLER_64_1635 ();
 sg13g2_decap_4 FILLER_64_1642 ();
 sg13g2_fill_2 FILLER_64_1646 ();
 sg13g2_decap_8 FILLER_64_1656 ();
 sg13g2_decap_8 FILLER_64_1663 ();
 sg13g2_decap_8 FILLER_64_1670 ();
 sg13g2_decap_8 FILLER_64_1677 ();
 sg13g2_decap_8 FILLER_64_1684 ();
 sg13g2_decap_8 FILLER_64_1691 ();
 sg13g2_decap_8 FILLER_64_1698 ();
 sg13g2_decap_8 FILLER_64_1705 ();
 sg13g2_decap_8 FILLER_64_1712 ();
 sg13g2_decap_4 FILLER_64_1719 ();
 sg13g2_fill_1 FILLER_64_1723 ();
 sg13g2_decap_8 FILLER_64_1734 ();
 sg13g2_decap_8 FILLER_64_1741 ();
 sg13g2_decap_8 FILLER_64_1748 ();
 sg13g2_decap_8 FILLER_64_1755 ();
 sg13g2_decap_8 FILLER_64_1762 ();
 sg13g2_decap_8 FILLER_64_1769 ();
 sg13g2_decap_8 FILLER_64_1776 ();
 sg13g2_decap_8 FILLER_64_1783 ();
 sg13g2_decap_8 FILLER_64_1790 ();
 sg13g2_decap_8 FILLER_64_1797 ();
 sg13g2_decap_8 FILLER_64_1804 ();
 sg13g2_decap_8 FILLER_64_1811 ();
 sg13g2_fill_2 FILLER_64_1818 ();
 sg13g2_fill_1 FILLER_64_1820 ();
 sg13g2_fill_2 FILLER_64_1831 ();
 sg13g2_decap_8 FILLER_64_1885 ();
 sg13g2_decap_8 FILLER_64_1892 ();
 sg13g2_decap_8 FILLER_64_1899 ();
 sg13g2_decap_8 FILLER_64_1906 ();
 sg13g2_decap_8 FILLER_64_1913 ();
 sg13g2_decap_8 FILLER_64_1920 ();
 sg13g2_decap_8 FILLER_64_1927 ();
 sg13g2_decap_8 FILLER_64_1934 ();
 sg13g2_decap_8 FILLER_64_1941 ();
 sg13g2_decap_8 FILLER_64_1948 ();
 sg13g2_decap_8 FILLER_64_1955 ();
 sg13g2_decap_8 FILLER_64_1962 ();
 sg13g2_decap_4 FILLER_64_1969 ();
 sg13g2_decap_8 FILLER_64_2004 ();
 sg13g2_decap_8 FILLER_64_2011 ();
 sg13g2_decap_8 FILLER_64_2018 ();
 sg13g2_decap_8 FILLER_64_2025 ();
 sg13g2_fill_2 FILLER_64_2032 ();
 sg13g2_fill_1 FILLER_64_2034 ();
 sg13g2_decap_8 FILLER_64_2041 ();
 sg13g2_decap_8 FILLER_64_2048 ();
 sg13g2_decap_8 FILLER_64_2055 ();
 sg13g2_decap_8 FILLER_64_2062 ();
 sg13g2_decap_8 FILLER_64_2105 ();
 sg13g2_decap_8 FILLER_64_2112 ();
 sg13g2_decap_8 FILLER_64_2119 ();
 sg13g2_decap_8 FILLER_64_2126 ();
 sg13g2_decap_8 FILLER_64_2133 ();
 sg13g2_decap_8 FILLER_64_2140 ();
 sg13g2_decap_8 FILLER_64_2147 ();
 sg13g2_decap_8 FILLER_64_2154 ();
 sg13g2_decap_8 FILLER_64_2161 ();
 sg13g2_decap_4 FILLER_64_2168 ();
 sg13g2_fill_1 FILLER_64_2198 ();
 sg13g2_decap_8 FILLER_64_2205 ();
 sg13g2_decap_8 FILLER_64_2212 ();
 sg13g2_decap_4 FILLER_64_2219 ();
 sg13g2_fill_1 FILLER_64_2223 ();
 sg13g2_decap_8 FILLER_64_2250 ();
 sg13g2_decap_8 FILLER_64_2257 ();
 sg13g2_decap_8 FILLER_64_2308 ();
 sg13g2_decap_8 FILLER_64_2315 ();
 sg13g2_fill_2 FILLER_64_2322 ();
 sg13g2_fill_1 FILLER_64_2324 ();
 sg13g2_decap_8 FILLER_64_2351 ();
 sg13g2_decap_8 FILLER_64_2358 ();
 sg13g2_decap_8 FILLER_64_2365 ();
 sg13g2_decap_8 FILLER_64_2372 ();
 sg13g2_decap_4 FILLER_64_2379 ();
 sg13g2_decap_8 FILLER_64_2393 ();
 sg13g2_decap_8 FILLER_64_2400 ();
 sg13g2_decap_8 FILLER_64_2407 ();
 sg13g2_decap_8 FILLER_64_2414 ();
 sg13g2_decap_8 FILLER_64_2421 ();
 sg13g2_decap_8 FILLER_64_2428 ();
 sg13g2_fill_2 FILLER_64_2435 ();
 sg13g2_decap_8 FILLER_64_2457 ();
 sg13g2_decap_8 FILLER_64_2464 ();
 sg13g2_decap_8 FILLER_64_2471 ();
 sg13g2_decap_8 FILLER_64_2478 ();
 sg13g2_fill_2 FILLER_64_2485 ();
 sg13g2_fill_1 FILLER_64_2487 ();
 sg13g2_decap_8 FILLER_64_2502 ();
 sg13g2_decap_4 FILLER_64_2509 ();
 sg13g2_fill_1 FILLER_64_2513 ();
 sg13g2_decap_8 FILLER_64_2524 ();
 sg13g2_decap_8 FILLER_64_2531 ();
 sg13g2_decap_8 FILLER_64_2538 ();
 sg13g2_decap_8 FILLER_64_2545 ();
 sg13g2_decap_8 FILLER_64_2552 ();
 sg13g2_decap_8 FILLER_64_2559 ();
 sg13g2_decap_4 FILLER_64_2566 ();
 sg13g2_fill_1 FILLER_64_2570 ();
 sg13g2_decap_4 FILLER_64_2582 ();
 sg13g2_fill_2 FILLER_64_2586 ();
 sg13g2_decap_8 FILLER_64_2620 ();
 sg13g2_decap_8 FILLER_64_2627 ();
 sg13g2_decap_8 FILLER_64_2634 ();
 sg13g2_decap_4 FILLER_64_2641 ();
 sg13g2_fill_1 FILLER_64_2645 ();
 sg13g2_decap_8 FILLER_64_2672 ();
 sg13g2_decap_8 FILLER_64_2679 ();
 sg13g2_fill_1 FILLER_64_2686 ();
 sg13g2_decap_8 FILLER_64_2723 ();
 sg13g2_decap_8 FILLER_64_2730 ();
 sg13g2_decap_8 FILLER_64_2737 ();
 sg13g2_decap_8 FILLER_64_2744 ();
 sg13g2_fill_2 FILLER_64_2751 ();
 sg13g2_decap_8 FILLER_64_2779 ();
 sg13g2_decap_8 FILLER_64_2786 ();
 sg13g2_decap_8 FILLER_64_2793 ();
 sg13g2_decap_8 FILLER_64_2800 ();
 sg13g2_decap_8 FILLER_64_2807 ();
 sg13g2_decap_8 FILLER_64_2814 ();
 sg13g2_decap_8 FILLER_64_2821 ();
 sg13g2_decap_8 FILLER_64_2828 ();
 sg13g2_decap_4 FILLER_64_2835 ();
 sg13g2_fill_2 FILLER_64_2839 ();
 sg13g2_decap_8 FILLER_64_2877 ();
 sg13g2_decap_8 FILLER_64_2884 ();
 sg13g2_fill_2 FILLER_64_2927 ();
 sg13g2_decap_8 FILLER_64_2955 ();
 sg13g2_decap_8 FILLER_64_2962 ();
 sg13g2_decap_8 FILLER_64_2969 ();
 sg13g2_decap_4 FILLER_64_2976 ();
 sg13g2_decap_8 FILLER_64_2986 ();
 sg13g2_decap_8 FILLER_64_2993 ();
 sg13g2_decap_8 FILLER_64_3000 ();
 sg13g2_decap_4 FILLER_64_3007 ();
 sg13g2_decap_8 FILLER_64_3047 ();
 sg13g2_decap_8 FILLER_64_3054 ();
 sg13g2_fill_2 FILLER_64_3061 ();
 sg13g2_fill_1 FILLER_64_3063 ();
 sg13g2_fill_2 FILLER_64_3074 ();
 sg13g2_decap_8 FILLER_64_3082 ();
 sg13g2_decap_4 FILLER_64_3089 ();
 sg13g2_fill_1 FILLER_64_3093 ();
 sg13g2_decap_8 FILLER_64_3120 ();
 sg13g2_decap_8 FILLER_64_3127 ();
 sg13g2_decap_8 FILLER_64_3134 ();
 sg13g2_fill_2 FILLER_64_3141 ();
 sg13g2_decap_8 FILLER_64_3169 ();
 sg13g2_decap_8 FILLER_64_3176 ();
 sg13g2_decap_8 FILLER_64_3183 ();
 sg13g2_decap_8 FILLER_64_3190 ();
 sg13g2_decap_8 FILLER_64_3197 ();
 sg13g2_decap_8 FILLER_64_3204 ();
 sg13g2_decap_4 FILLER_64_3211 ();
 sg13g2_fill_1 FILLER_64_3215 ();
 sg13g2_decap_8 FILLER_64_3222 ();
 sg13g2_decap_8 FILLER_64_3229 ();
 sg13g2_decap_8 FILLER_64_3236 ();
 sg13g2_decap_8 FILLER_64_3243 ();
 sg13g2_decap_8 FILLER_64_3250 ();
 sg13g2_fill_1 FILLER_64_3257 ();
 sg13g2_decap_8 FILLER_64_3284 ();
 sg13g2_decap_8 FILLER_64_3291 ();
 sg13g2_decap_8 FILLER_64_3298 ();
 sg13g2_decap_8 FILLER_64_3305 ();
 sg13g2_decap_8 FILLER_64_3312 ();
 sg13g2_decap_8 FILLER_64_3319 ();
 sg13g2_decap_8 FILLER_64_3326 ();
 sg13g2_decap_8 FILLER_64_3333 ();
 sg13g2_decap_8 FILLER_64_3340 ();
 sg13g2_decap_8 FILLER_64_3347 ();
 sg13g2_decap_8 FILLER_64_3354 ();
 sg13g2_decap_8 FILLER_64_3361 ();
 sg13g2_decap_8 FILLER_64_3368 ();
 sg13g2_fill_1 FILLER_64_3375 ();
 sg13g2_decap_4 FILLER_64_3386 ();
 sg13g2_fill_2 FILLER_64_3390 ();
 sg13g2_decap_8 FILLER_64_3395 ();
 sg13g2_decap_8 FILLER_64_3402 ();
 sg13g2_decap_8 FILLER_64_3409 ();
 sg13g2_decap_8 FILLER_64_3416 ();
 sg13g2_decap_8 FILLER_64_3423 ();
 sg13g2_decap_8 FILLER_64_3430 ();
 sg13g2_decap_8 FILLER_64_3437 ();
 sg13g2_decap_8 FILLER_64_3444 ();
 sg13g2_fill_2 FILLER_64_3451 ();
 sg13g2_fill_1 FILLER_64_3453 ();
 sg13g2_decap_8 FILLER_64_3471 ();
 sg13g2_decap_8 FILLER_64_3478 ();
 sg13g2_decap_8 FILLER_64_3485 ();
 sg13g2_decap_8 FILLER_64_3492 ();
 sg13g2_fill_2 FILLER_64_3499 ();
 sg13g2_fill_1 FILLER_64_3501 ();
 sg13g2_decap_8 FILLER_64_3512 ();
 sg13g2_decap_8 FILLER_64_3519 ();
 sg13g2_decap_8 FILLER_64_3526 ();
 sg13g2_decap_8 FILLER_64_3533 ();
 sg13g2_decap_8 FILLER_64_3540 ();
 sg13g2_decap_8 FILLER_64_3547 ();
 sg13g2_decap_8 FILLER_64_3554 ();
 sg13g2_decap_8 FILLER_64_3561 ();
 sg13g2_decap_8 FILLER_64_3568 ();
 sg13g2_decap_4 FILLER_64_3575 ();
 sg13g2_fill_1 FILLER_64_3579 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_8 FILLER_65_59 ();
 sg13g2_decap_4 FILLER_65_66 ();
 sg13g2_fill_2 FILLER_65_70 ();
 sg13g2_decap_8 FILLER_65_102 ();
 sg13g2_decap_4 FILLER_65_109 ();
 sg13g2_fill_2 FILLER_65_113 ();
 sg13g2_decap_8 FILLER_65_150 ();
 sg13g2_decap_8 FILLER_65_157 ();
 sg13g2_decap_8 FILLER_65_164 ();
 sg13g2_decap_8 FILLER_65_176 ();
 sg13g2_decap_8 FILLER_65_183 ();
 sg13g2_decap_8 FILLER_65_190 ();
 sg13g2_decap_8 FILLER_65_197 ();
 sg13g2_decap_8 FILLER_65_204 ();
 sg13g2_decap_8 FILLER_65_211 ();
 sg13g2_decap_8 FILLER_65_218 ();
 sg13g2_decap_8 FILLER_65_225 ();
 sg13g2_fill_2 FILLER_65_232 ();
 sg13g2_fill_1 FILLER_65_239 ();
 sg13g2_fill_1 FILLER_65_254 ();
 sg13g2_fill_2 FILLER_65_275 ();
 sg13g2_fill_2 FILLER_65_283 ();
 sg13g2_fill_1 FILLER_65_285 ();
 sg13g2_fill_2 FILLER_65_289 ();
 sg13g2_fill_1 FILLER_65_306 ();
 sg13g2_decap_8 FILLER_65_358 ();
 sg13g2_decap_8 FILLER_65_365 ();
 sg13g2_decap_8 FILLER_65_372 ();
 sg13g2_decap_4 FILLER_65_379 ();
 sg13g2_fill_2 FILLER_65_383 ();
 sg13g2_decap_8 FILLER_65_398 ();
 sg13g2_decap_8 FILLER_65_405 ();
 sg13g2_decap_8 FILLER_65_412 ();
 sg13g2_decap_8 FILLER_65_419 ();
 sg13g2_decap_8 FILLER_65_426 ();
 sg13g2_decap_4 FILLER_65_433 ();
 sg13g2_decap_8 FILLER_65_442 ();
 sg13g2_decap_8 FILLER_65_449 ();
 sg13g2_decap_8 FILLER_65_456 ();
 sg13g2_decap_8 FILLER_65_463 ();
 sg13g2_decap_8 FILLER_65_470 ();
 sg13g2_decap_8 FILLER_65_477 ();
 sg13g2_decap_8 FILLER_65_484 ();
 sg13g2_decap_8 FILLER_65_491 ();
 sg13g2_decap_8 FILLER_65_498 ();
 sg13g2_decap_8 FILLER_65_505 ();
 sg13g2_fill_2 FILLER_65_512 ();
 sg13g2_fill_1 FILLER_65_514 ();
 sg13g2_decap_4 FILLER_65_519 ();
 sg13g2_decap_8 FILLER_65_528 ();
 sg13g2_decap_4 FILLER_65_535 ();
 sg13g2_decap_8 FILLER_65_553 ();
 sg13g2_decap_8 FILLER_65_560 ();
 sg13g2_fill_2 FILLER_65_567 ();
 sg13g2_decap_8 FILLER_65_577 ();
 sg13g2_fill_2 FILLER_65_584 ();
 sg13g2_fill_2 FILLER_65_596 ();
 sg13g2_decap_8 FILLER_65_610 ();
 sg13g2_decap_8 FILLER_65_617 ();
 sg13g2_decap_8 FILLER_65_624 ();
 sg13g2_fill_2 FILLER_65_631 ();
 sg13g2_fill_1 FILLER_65_633 ();
 sg13g2_decap_8 FILLER_65_638 ();
 sg13g2_fill_1 FILLER_65_645 ();
 sg13g2_decap_8 FILLER_65_663 ();
 sg13g2_decap_8 FILLER_65_670 ();
 sg13g2_decap_4 FILLER_65_677 ();
 sg13g2_fill_2 FILLER_65_681 ();
 sg13g2_fill_1 FILLER_65_693 ();
 sg13g2_decap_8 FILLER_65_700 ();
 sg13g2_decap_8 FILLER_65_707 ();
 sg13g2_fill_1 FILLER_65_714 ();
 sg13g2_decap_8 FILLER_65_724 ();
 sg13g2_decap_8 FILLER_65_731 ();
 sg13g2_decap_8 FILLER_65_738 ();
 sg13g2_decap_8 FILLER_65_745 ();
 sg13g2_decap_8 FILLER_65_752 ();
 sg13g2_decap_4 FILLER_65_759 ();
 sg13g2_fill_1 FILLER_65_763 ();
 sg13g2_decap_8 FILLER_65_768 ();
 sg13g2_decap_8 FILLER_65_775 ();
 sg13g2_decap_8 FILLER_65_782 ();
 sg13g2_decap_4 FILLER_65_789 ();
 sg13g2_fill_1 FILLER_65_793 ();
 sg13g2_fill_2 FILLER_65_820 ();
 sg13g2_fill_1 FILLER_65_822 ();
 sg13g2_decap_4 FILLER_65_831 ();
 sg13g2_fill_1 FILLER_65_835 ();
 sg13g2_decap_8 FILLER_65_848 ();
 sg13g2_decap_8 FILLER_65_855 ();
 sg13g2_decap_8 FILLER_65_862 ();
 sg13g2_decap_4 FILLER_65_869 ();
 sg13g2_decap_8 FILLER_65_883 ();
 sg13g2_decap_8 FILLER_65_890 ();
 sg13g2_decap_8 FILLER_65_897 ();
 sg13g2_decap_8 FILLER_65_904 ();
 sg13g2_decap_8 FILLER_65_911 ();
 sg13g2_decap_8 FILLER_65_918 ();
 sg13g2_decap_8 FILLER_65_930 ();
 sg13g2_decap_8 FILLER_65_937 ();
 sg13g2_decap_8 FILLER_65_944 ();
 sg13g2_decap_8 FILLER_65_951 ();
 sg13g2_decap_8 FILLER_65_958 ();
 sg13g2_decap_8 FILLER_65_970 ();
 sg13g2_decap_4 FILLER_65_977 ();
 sg13g2_fill_1 FILLER_65_981 ();
 sg13g2_decap_4 FILLER_65_987 ();
 sg13g2_fill_1 FILLER_65_991 ();
 sg13g2_decap_8 FILLER_65_997 ();
 sg13g2_decap_8 FILLER_65_1004 ();
 sg13g2_decap_8 FILLER_65_1011 ();
 sg13g2_decap_8 FILLER_65_1018 ();
 sg13g2_decap_8 FILLER_65_1025 ();
 sg13g2_decap_4 FILLER_65_1032 ();
 sg13g2_decap_8 FILLER_65_1065 ();
 sg13g2_decap_8 FILLER_65_1072 ();
 sg13g2_decap_8 FILLER_65_1079 ();
 sg13g2_decap_8 FILLER_65_1086 ();
 sg13g2_fill_1 FILLER_65_1093 ();
 sg13g2_fill_2 FILLER_65_1097 ();
 sg13g2_fill_1 FILLER_65_1099 ();
 sg13g2_decap_8 FILLER_65_1108 ();
 sg13g2_decap_8 FILLER_65_1115 ();
 sg13g2_decap_8 FILLER_65_1122 ();
 sg13g2_fill_2 FILLER_65_1129 ();
 sg13g2_fill_1 FILLER_65_1131 ();
 sg13g2_fill_2 FILLER_65_1153 ();
 sg13g2_fill_1 FILLER_65_1155 ();
 sg13g2_fill_1 FILLER_65_1167 ();
 sg13g2_decap_8 FILLER_65_1188 ();
 sg13g2_decap_8 FILLER_65_1195 ();
 sg13g2_decap_8 FILLER_65_1202 ();
 sg13g2_decap_8 FILLER_65_1209 ();
 sg13g2_decap_8 FILLER_65_1216 ();
 sg13g2_decap_8 FILLER_65_1223 ();
 sg13g2_decap_4 FILLER_65_1230 ();
 sg13g2_fill_1 FILLER_65_1234 ();
 sg13g2_decap_8 FILLER_65_1238 ();
 sg13g2_decap_8 FILLER_65_1245 ();
 sg13g2_decap_8 FILLER_65_1252 ();
 sg13g2_decap_8 FILLER_65_1259 ();
 sg13g2_decap_4 FILLER_65_1266 ();
 sg13g2_fill_1 FILLER_65_1270 ();
 sg13g2_decap_8 FILLER_65_1275 ();
 sg13g2_decap_8 FILLER_65_1282 ();
 sg13g2_decap_8 FILLER_65_1289 ();
 sg13g2_decap_8 FILLER_65_1296 ();
 sg13g2_decap_8 FILLER_65_1303 ();
 sg13g2_decap_8 FILLER_65_1310 ();
 sg13g2_decap_4 FILLER_65_1317 ();
 sg13g2_fill_1 FILLER_65_1321 ();
 sg13g2_decap_8 FILLER_65_1382 ();
 sg13g2_fill_1 FILLER_65_1389 ();
 sg13g2_decap_8 FILLER_65_1400 ();
 sg13g2_decap_8 FILLER_65_1407 ();
 sg13g2_decap_8 FILLER_65_1414 ();
 sg13g2_decap_8 FILLER_65_1421 ();
 sg13g2_decap_8 FILLER_65_1428 ();
 sg13g2_decap_8 FILLER_65_1435 ();
 sg13g2_fill_2 FILLER_65_1442 ();
 sg13g2_fill_1 FILLER_65_1444 ();
 sg13g2_decap_8 FILLER_65_1481 ();
 sg13g2_decap_8 FILLER_65_1488 ();
 sg13g2_decap_4 FILLER_65_1495 ();
 sg13g2_decap_4 FILLER_65_1509 ();
 sg13g2_decap_8 FILLER_65_1539 ();
 sg13g2_decap_8 FILLER_65_1546 ();
 sg13g2_fill_2 FILLER_65_1553 ();
 sg13g2_fill_1 FILLER_65_1555 ();
 sg13g2_decap_8 FILLER_65_1586 ();
 sg13g2_decap_8 FILLER_65_1593 ();
 sg13g2_decap_8 FILLER_65_1600 ();
 sg13g2_decap_8 FILLER_65_1607 ();
 sg13g2_decap_8 FILLER_65_1614 ();
 sg13g2_decap_8 FILLER_65_1621 ();
 sg13g2_fill_2 FILLER_65_1628 ();
 sg13g2_decap_4 FILLER_65_1638 ();
 sg13g2_fill_1 FILLER_65_1642 ();
 sg13g2_decap_8 FILLER_65_1662 ();
 sg13g2_decap_8 FILLER_65_1669 ();
 sg13g2_decap_8 FILLER_65_1676 ();
 sg13g2_decap_8 FILLER_65_1683 ();
 sg13g2_decap_8 FILLER_65_1690 ();
 sg13g2_decap_8 FILLER_65_1697 ();
 sg13g2_decap_8 FILLER_65_1704 ();
 sg13g2_decap_8 FILLER_65_1711 ();
 sg13g2_decap_4 FILLER_65_1718 ();
 sg13g2_fill_2 FILLER_65_1756 ();
 sg13g2_fill_1 FILLER_65_1758 ();
 sg13g2_decap_8 FILLER_65_1769 ();
 sg13g2_decap_8 FILLER_65_1776 ();
 sg13g2_decap_8 FILLER_65_1783 ();
 sg13g2_fill_2 FILLER_65_1790 ();
 sg13g2_decap_8 FILLER_65_1826 ();
 sg13g2_decap_8 FILLER_65_1833 ();
 sg13g2_decap_8 FILLER_65_1840 ();
 sg13g2_decap_8 FILLER_65_1847 ();
 sg13g2_decap_8 FILLER_65_1854 ();
 sg13g2_decap_8 FILLER_65_1861 ();
 sg13g2_decap_8 FILLER_65_1868 ();
 sg13g2_decap_8 FILLER_65_1875 ();
 sg13g2_fill_2 FILLER_65_1882 ();
 sg13g2_decap_8 FILLER_65_1888 ();
 sg13g2_fill_1 FILLER_65_1895 ();
 sg13g2_decap_8 FILLER_65_1901 ();
 sg13g2_decap_8 FILLER_65_1908 ();
 sg13g2_decap_8 FILLER_65_1915 ();
 sg13g2_decap_8 FILLER_65_1922 ();
 sg13g2_decap_4 FILLER_65_1929 ();
 sg13g2_fill_1 FILLER_65_1933 ();
 sg13g2_decap_4 FILLER_65_1944 ();
 sg13g2_decap_8 FILLER_65_1954 ();
 sg13g2_decap_8 FILLER_65_1961 ();
 sg13g2_fill_2 FILLER_65_1968 ();
 sg13g2_fill_1 FILLER_65_1970 ();
 sg13g2_decap_8 FILLER_65_2009 ();
 sg13g2_decap_8 FILLER_65_2016 ();
 sg13g2_decap_8 FILLER_65_2023 ();
 sg13g2_decap_4 FILLER_65_2030 ();
 sg13g2_fill_2 FILLER_65_2034 ();
 sg13g2_decap_8 FILLER_65_2072 ();
 sg13g2_decap_8 FILLER_65_2079 ();
 sg13g2_fill_2 FILLER_65_2086 ();
 sg13g2_fill_1 FILLER_65_2088 ();
 sg13g2_decap_8 FILLER_65_2101 ();
 sg13g2_decap_8 FILLER_65_2108 ();
 sg13g2_decap_8 FILLER_65_2115 ();
 sg13g2_decap_8 FILLER_65_2122 ();
 sg13g2_decap_4 FILLER_65_2129 ();
 sg13g2_decap_8 FILLER_65_2137 ();
 sg13g2_decap_8 FILLER_65_2144 ();
 sg13g2_fill_2 FILLER_65_2151 ();
 sg13g2_fill_1 FILLER_65_2153 ();
 sg13g2_decap_8 FILLER_65_2164 ();
 sg13g2_decap_8 FILLER_65_2171 ();
 sg13g2_decap_8 FILLER_65_2178 ();
 sg13g2_decap_8 FILLER_65_2185 ();
 sg13g2_decap_8 FILLER_65_2192 ();
 sg13g2_decap_8 FILLER_65_2199 ();
 sg13g2_decap_8 FILLER_65_2206 ();
 sg13g2_decap_8 FILLER_65_2213 ();
 sg13g2_decap_8 FILLER_65_2220 ();
 sg13g2_decap_8 FILLER_65_2253 ();
 sg13g2_decap_8 FILLER_65_2260 ();
 sg13g2_decap_8 FILLER_65_2267 ();
 sg13g2_decap_8 FILLER_65_2274 ();
 sg13g2_fill_2 FILLER_65_2281 ();
 sg13g2_decap_8 FILLER_65_2298 ();
 sg13g2_decap_8 FILLER_65_2305 ();
 sg13g2_decap_8 FILLER_65_2312 ();
 sg13g2_decap_8 FILLER_65_2319 ();
 sg13g2_fill_2 FILLER_65_2326 ();
 sg13g2_fill_1 FILLER_65_2328 ();
 sg13g2_fill_2 FILLER_65_2333 ();
 sg13g2_decap_8 FILLER_65_2361 ();
 sg13g2_decap_8 FILLER_65_2368 ();
 sg13g2_decap_8 FILLER_65_2375 ();
 sg13g2_fill_2 FILLER_65_2382 ();
 sg13g2_decap_8 FILLER_65_2410 ();
 sg13g2_decap_8 FILLER_65_2417 ();
 sg13g2_decap_8 FILLER_65_2424 ();
 sg13g2_decap_8 FILLER_65_2431 ();
 sg13g2_decap_4 FILLER_65_2438 ();
 sg13g2_fill_1 FILLER_65_2442 ();
 sg13g2_decap_8 FILLER_65_2469 ();
 sg13g2_decap_8 FILLER_65_2476 ();
 sg13g2_fill_1 FILLER_65_2483 ();
 sg13g2_decap_4 FILLER_65_2510 ();
 sg13g2_fill_2 FILLER_65_2514 ();
 sg13g2_decap_8 FILLER_65_2542 ();
 sg13g2_decap_4 FILLER_65_2549 ();
 sg13g2_fill_2 FILLER_65_2553 ();
 sg13g2_decap_8 FILLER_65_2565 ();
 sg13g2_decap_8 FILLER_65_2572 ();
 sg13g2_decap_8 FILLER_65_2579 ();
 sg13g2_decap_8 FILLER_65_2586 ();
 sg13g2_decap_8 FILLER_65_2593 ();
 sg13g2_decap_8 FILLER_65_2600 ();
 sg13g2_decap_4 FILLER_65_2607 ();
 sg13g2_fill_1 FILLER_65_2611 ();
 sg13g2_decap_8 FILLER_65_2622 ();
 sg13g2_decap_8 FILLER_65_2629 ();
 sg13g2_decap_8 FILLER_65_2636 ();
 sg13g2_fill_2 FILLER_65_2643 ();
 sg13g2_decap_8 FILLER_65_2681 ();
 sg13g2_decap_8 FILLER_65_2688 ();
 sg13g2_decap_8 FILLER_65_2695 ();
 sg13g2_decap_8 FILLER_65_2702 ();
 sg13g2_decap_8 FILLER_65_2709 ();
 sg13g2_decap_8 FILLER_65_2716 ();
 sg13g2_decap_8 FILLER_65_2723 ();
 sg13g2_decap_8 FILLER_65_2730 ();
 sg13g2_decap_8 FILLER_65_2737 ();
 sg13g2_decap_8 FILLER_65_2744 ();
 sg13g2_fill_2 FILLER_65_2751 ();
 sg13g2_decap_8 FILLER_65_2763 ();
 sg13g2_decap_8 FILLER_65_2770 ();
 sg13g2_decap_8 FILLER_65_2777 ();
 sg13g2_decap_8 FILLER_65_2784 ();
 sg13g2_decap_8 FILLER_65_2791 ();
 sg13g2_decap_8 FILLER_65_2798 ();
 sg13g2_fill_2 FILLER_65_2805 ();
 sg13g2_decap_8 FILLER_65_2833 ();
 sg13g2_decap_8 FILLER_65_2840 ();
 sg13g2_decap_4 FILLER_65_2847 ();
 sg13g2_fill_1 FILLER_65_2851 ();
 sg13g2_decap_8 FILLER_65_2878 ();
 sg13g2_decap_8 FILLER_65_2885 ();
 sg13g2_fill_1 FILLER_65_2892 ();
 sg13g2_decap_8 FILLER_65_2955 ();
 sg13g2_decap_8 FILLER_65_2962 ();
 sg13g2_fill_2 FILLER_65_2969 ();
 sg13g2_decap_4 FILLER_65_3007 ();
 sg13g2_fill_1 FILLER_65_3011 ();
 sg13g2_decap_8 FILLER_65_3126 ();
 sg13g2_fill_1 FILLER_65_3133 ();
 sg13g2_decap_8 FILLER_65_3168 ();
 sg13g2_decap_8 FILLER_65_3175 ();
 sg13g2_decap_8 FILLER_65_3182 ();
 sg13g2_decap_8 FILLER_65_3189 ();
 sg13g2_decap_8 FILLER_65_3196 ();
 sg13g2_fill_1 FILLER_65_3203 ();
 sg13g2_decap_8 FILLER_65_3230 ();
 sg13g2_decap_8 FILLER_65_3237 ();
 sg13g2_fill_2 FILLER_65_3244 ();
 sg13g2_decap_8 FILLER_65_3262 ();
 sg13g2_decap_4 FILLER_65_3269 ();
 sg13g2_fill_1 FILLER_65_3273 ();
 sg13g2_decap_8 FILLER_65_3284 ();
 sg13g2_decap_8 FILLER_65_3291 ();
 sg13g2_decap_8 FILLER_65_3298 ();
 sg13g2_decap_8 FILLER_65_3305 ();
 sg13g2_decap_8 FILLER_65_3312 ();
 sg13g2_decap_8 FILLER_65_3319 ();
 sg13g2_decap_8 FILLER_65_3326 ();
 sg13g2_decap_8 FILLER_65_3333 ();
 sg13g2_decap_8 FILLER_65_3340 ();
 sg13g2_decap_8 FILLER_65_3347 ();
 sg13g2_decap_8 FILLER_65_3354 ();
 sg13g2_decap_8 FILLER_65_3361 ();
 sg13g2_decap_8 FILLER_65_3368 ();
 sg13g2_decap_8 FILLER_65_3375 ();
 sg13g2_decap_8 FILLER_65_3382 ();
 sg13g2_decap_8 FILLER_65_3389 ();
 sg13g2_decap_8 FILLER_65_3396 ();
 sg13g2_decap_8 FILLER_65_3403 ();
 sg13g2_decap_8 FILLER_65_3410 ();
 sg13g2_decap_8 FILLER_65_3417 ();
 sg13g2_fill_1 FILLER_65_3424 ();
 sg13g2_fill_1 FILLER_65_3430 ();
 sg13g2_decap_8 FILLER_65_3435 ();
 sg13g2_decap_8 FILLER_65_3442 ();
 sg13g2_decap_8 FILLER_65_3449 ();
 sg13g2_decap_8 FILLER_65_3456 ();
 sg13g2_decap_8 FILLER_65_3463 ();
 sg13g2_decap_8 FILLER_65_3470 ();
 sg13g2_decap_8 FILLER_65_3477 ();
 sg13g2_decap_4 FILLER_65_3484 ();
 sg13g2_fill_2 FILLER_65_3488 ();
 sg13g2_decap_8 FILLER_65_3495 ();
 sg13g2_fill_2 FILLER_65_3502 ();
 sg13g2_decap_8 FILLER_65_3509 ();
 sg13g2_decap_8 FILLER_65_3516 ();
 sg13g2_decap_8 FILLER_65_3523 ();
 sg13g2_decap_8 FILLER_65_3530 ();
 sg13g2_decap_8 FILLER_65_3537 ();
 sg13g2_decap_8 FILLER_65_3544 ();
 sg13g2_decap_8 FILLER_65_3551 ();
 sg13g2_decap_8 FILLER_65_3558 ();
 sg13g2_decap_8 FILLER_65_3565 ();
 sg13g2_decap_8 FILLER_65_3572 ();
 sg13g2_fill_1 FILLER_65_3579 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_8 FILLER_66_7 ();
 sg13g2_fill_2 FILLER_66_14 ();
 sg13g2_decap_8 FILLER_66_56 ();
 sg13g2_decap_8 FILLER_66_63 ();
 sg13g2_decap_4 FILLER_66_70 ();
 sg13g2_fill_1 FILLER_66_74 ();
 sg13g2_decap_8 FILLER_66_102 ();
 sg13g2_decap_8 FILLER_66_109 ();
 sg13g2_decap_4 FILLER_66_116 ();
 sg13g2_fill_1 FILLER_66_120 ();
 sg13g2_fill_1 FILLER_66_131 ();
 sg13g2_decap_8 FILLER_66_139 ();
 sg13g2_decap_8 FILLER_66_146 ();
 sg13g2_decap_8 FILLER_66_153 ();
 sg13g2_decap_8 FILLER_66_160 ();
 sg13g2_decap_8 FILLER_66_167 ();
 sg13g2_decap_8 FILLER_66_174 ();
 sg13g2_decap_4 FILLER_66_188 ();
 sg13g2_fill_2 FILLER_66_192 ();
 sg13g2_decap_8 FILLER_66_203 ();
 sg13g2_decap_8 FILLER_66_210 ();
 sg13g2_decap_8 FILLER_66_217 ();
 sg13g2_decap_8 FILLER_66_224 ();
 sg13g2_decap_8 FILLER_66_231 ();
 sg13g2_decap_4 FILLER_66_238 ();
 sg13g2_fill_2 FILLER_66_242 ();
 sg13g2_decap_4 FILLER_66_248 ();
 sg13g2_fill_2 FILLER_66_252 ();
 sg13g2_fill_1 FILLER_66_268 ();
 sg13g2_fill_2 FILLER_66_307 ();
 sg13g2_fill_1 FILLER_66_309 ();
 sg13g2_decap_8 FILLER_66_313 ();
 sg13g2_fill_2 FILLER_66_336 ();
 sg13g2_fill_2 FILLER_66_346 ();
 sg13g2_fill_1 FILLER_66_348 ();
 sg13g2_decap_8 FILLER_66_366 ();
 sg13g2_decap_8 FILLER_66_373 ();
 sg13g2_decap_8 FILLER_66_380 ();
 sg13g2_decap_8 FILLER_66_387 ();
 sg13g2_decap_8 FILLER_66_394 ();
 sg13g2_decap_8 FILLER_66_401 ();
 sg13g2_decap_8 FILLER_66_408 ();
 sg13g2_decap_8 FILLER_66_415 ();
 sg13g2_decap_8 FILLER_66_422 ();
 sg13g2_decap_8 FILLER_66_429 ();
 sg13g2_decap_8 FILLER_66_436 ();
 sg13g2_decap_8 FILLER_66_443 ();
 sg13g2_decap_8 FILLER_66_450 ();
 sg13g2_decap_4 FILLER_66_457 ();
 sg13g2_decap_8 FILLER_66_476 ();
 sg13g2_decap_8 FILLER_66_483 ();
 sg13g2_decap_8 FILLER_66_490 ();
 sg13g2_decap_8 FILLER_66_497 ();
 sg13g2_decap_8 FILLER_66_504 ();
 sg13g2_decap_4 FILLER_66_511 ();
 sg13g2_fill_2 FILLER_66_515 ();
 sg13g2_decap_8 FILLER_66_536 ();
 sg13g2_decap_4 FILLER_66_543 ();
 sg13g2_fill_2 FILLER_66_547 ();
 sg13g2_decap_8 FILLER_66_553 ();
 sg13g2_decap_8 FILLER_66_560 ();
 sg13g2_fill_2 FILLER_66_567 ();
 sg13g2_decap_8 FILLER_66_592 ();
 sg13g2_decap_8 FILLER_66_604 ();
 sg13g2_decap_4 FILLER_66_611 ();
 sg13g2_fill_2 FILLER_66_615 ();
 sg13g2_decap_8 FILLER_66_623 ();
 sg13g2_decap_8 FILLER_66_630 ();
 sg13g2_decap_8 FILLER_66_637 ();
 sg13g2_fill_2 FILLER_66_644 ();
 sg13g2_decap_8 FILLER_66_658 ();
 sg13g2_decap_8 FILLER_66_665 ();
 sg13g2_decap_8 FILLER_66_672 ();
 sg13g2_decap_4 FILLER_66_679 ();
 sg13g2_fill_1 FILLER_66_683 ();
 sg13g2_decap_8 FILLER_66_688 ();
 sg13g2_decap_8 FILLER_66_695 ();
 sg13g2_decap_8 FILLER_66_702 ();
 sg13g2_fill_2 FILLER_66_709 ();
 sg13g2_fill_1 FILLER_66_711 ();
 sg13g2_decap_8 FILLER_66_766 ();
 sg13g2_decap_8 FILLER_66_773 ();
 sg13g2_fill_1 FILLER_66_813 ();
 sg13g2_decap_8 FILLER_66_819 ();
 sg13g2_decap_8 FILLER_66_826 ();
 sg13g2_decap_8 FILLER_66_833 ();
 sg13g2_decap_8 FILLER_66_840 ();
 sg13g2_decap_8 FILLER_66_847 ();
 sg13g2_decap_8 FILLER_66_858 ();
 sg13g2_decap_8 FILLER_66_865 ();
 sg13g2_decap_8 FILLER_66_872 ();
 sg13g2_decap_8 FILLER_66_879 ();
 sg13g2_decap_8 FILLER_66_886 ();
 sg13g2_decap_8 FILLER_66_893 ();
 sg13g2_decap_4 FILLER_66_900 ();
 sg13g2_decap_8 FILLER_66_935 ();
 sg13g2_decap_8 FILLER_66_942 ();
 sg13g2_decap_4 FILLER_66_949 ();
 sg13g2_fill_2 FILLER_66_958 ();
 sg13g2_fill_1 FILLER_66_960 ();
 sg13g2_fill_2 FILLER_66_969 ();
 sg13g2_decap_4 FILLER_66_979 ();
 sg13g2_fill_1 FILLER_66_983 ();
 sg13g2_decap_4 FILLER_66_992 ();
 sg13g2_decap_8 FILLER_66_1019 ();
 sg13g2_decap_8 FILLER_66_1026 ();
 sg13g2_decap_8 FILLER_66_1051 ();
 sg13g2_decap_8 FILLER_66_1058 ();
 sg13g2_decap_8 FILLER_66_1065 ();
 sg13g2_decap_8 FILLER_66_1072 ();
 sg13g2_decap_8 FILLER_66_1079 ();
 sg13g2_decap_8 FILLER_66_1086 ();
 sg13g2_decap_8 FILLER_66_1099 ();
 sg13g2_decap_8 FILLER_66_1106 ();
 sg13g2_fill_2 FILLER_66_1125 ();
 sg13g2_fill_1 FILLER_66_1127 ();
 sg13g2_fill_2 FILLER_66_1140 ();
 sg13g2_fill_2 FILLER_66_1169 ();
 sg13g2_fill_2 FILLER_66_1176 ();
 sg13g2_decap_8 FILLER_66_1204 ();
 sg13g2_decap_8 FILLER_66_1211 ();
 sg13g2_decap_8 FILLER_66_1218 ();
 sg13g2_decap_8 FILLER_66_1225 ();
 sg13g2_fill_2 FILLER_66_1232 ();
 sg13g2_fill_1 FILLER_66_1234 ();
 sg13g2_decap_8 FILLER_66_1243 ();
 sg13g2_fill_2 FILLER_66_1263 ();
 sg13g2_decap_8 FILLER_66_1280 ();
 sg13g2_decap_8 FILLER_66_1287 ();
 sg13g2_decap_8 FILLER_66_1294 ();
 sg13g2_decap_8 FILLER_66_1301 ();
 sg13g2_decap_8 FILLER_66_1308 ();
 sg13g2_decap_8 FILLER_66_1315 ();
 sg13g2_decap_8 FILLER_66_1322 ();
 sg13g2_fill_1 FILLER_66_1329 ();
 sg13g2_decap_8 FILLER_66_1366 ();
 sg13g2_decap_8 FILLER_66_1373 ();
 sg13g2_fill_1 FILLER_66_1380 ();
 sg13g2_decap_8 FILLER_66_1407 ();
 sg13g2_decap_8 FILLER_66_1414 ();
 sg13g2_decap_4 FILLER_66_1421 ();
 sg13g2_fill_2 FILLER_66_1425 ();
 sg13g2_decap_8 FILLER_66_1433 ();
 sg13g2_decap_4 FILLER_66_1440 ();
 sg13g2_fill_1 FILLER_66_1444 ();
 sg13g2_decap_4 FILLER_66_1455 ();
 sg13g2_decap_8 FILLER_66_1485 ();
 sg13g2_decap_8 FILLER_66_1492 ();
 sg13g2_decap_8 FILLER_66_1499 ();
 sg13g2_fill_1 FILLER_66_1506 ();
 sg13g2_decap_8 FILLER_66_1543 ();
 sg13g2_decap_4 FILLER_66_1570 ();
 sg13g2_decap_8 FILLER_66_1592 ();
 sg13g2_fill_1 FILLER_66_1599 ();
 sg13g2_decap_8 FILLER_66_1613 ();
 sg13g2_decap_8 FILLER_66_1620 ();
 sg13g2_decap_8 FILLER_66_1627 ();
 sg13g2_decap_8 FILLER_66_1634 ();
 sg13g2_fill_2 FILLER_66_1641 ();
 sg13g2_fill_1 FILLER_66_1643 ();
 sg13g2_decap_8 FILLER_66_1649 ();
 sg13g2_decap_8 FILLER_66_1656 ();
 sg13g2_fill_1 FILLER_66_1673 ();
 sg13g2_decap_8 FILLER_66_1713 ();
 sg13g2_decap_8 FILLER_66_1720 ();
 sg13g2_decap_8 FILLER_66_1727 ();
 sg13g2_decap_8 FILLER_66_1734 ();
 sg13g2_decap_8 FILLER_66_1741 ();
 sg13g2_decap_8 FILLER_66_1748 ();
 sg13g2_decap_4 FILLER_66_1755 ();
 sg13g2_decap_8 FILLER_66_1785 ();
 sg13g2_decap_8 FILLER_66_1792 ();
 sg13g2_decap_8 FILLER_66_1799 ();
 sg13g2_decap_8 FILLER_66_1806 ();
 sg13g2_fill_2 FILLER_66_1813 ();
 sg13g2_decap_8 FILLER_66_1823 ();
 sg13g2_decap_8 FILLER_66_1830 ();
 sg13g2_decap_8 FILLER_66_1837 ();
 sg13g2_fill_2 FILLER_66_1844 ();
 sg13g2_decap_4 FILLER_66_1850 ();
 sg13g2_fill_2 FILLER_66_1859 ();
 sg13g2_fill_1 FILLER_66_1866 ();
 sg13g2_fill_2 FILLER_66_1887 ();
 sg13g2_fill_1 FILLER_66_1889 ();
 sg13g2_decap_8 FILLER_66_1895 ();
 sg13g2_decap_8 FILLER_66_1902 ();
 sg13g2_fill_2 FILLER_66_1909 ();
 sg13g2_decap_8 FILLER_66_1942 ();
 sg13g2_decap_8 FILLER_66_1949 ();
 sg13g2_decap_8 FILLER_66_1956 ();
 sg13g2_decap_8 FILLER_66_1963 ();
 sg13g2_decap_8 FILLER_66_1970 ();
 sg13g2_fill_1 FILLER_66_1989 ();
 sg13g2_decap_8 FILLER_66_2013 ();
 sg13g2_decap_8 FILLER_66_2056 ();
 sg13g2_decap_8 FILLER_66_2063 ();
 sg13g2_decap_8 FILLER_66_2070 ();
 sg13g2_decap_8 FILLER_66_2077 ();
 sg13g2_decap_8 FILLER_66_2084 ();
 sg13g2_decap_8 FILLER_66_2091 ();
 sg13g2_decap_8 FILLER_66_2098 ();
 sg13g2_decap_8 FILLER_66_2105 ();
 sg13g2_decap_8 FILLER_66_2112 ();
 sg13g2_decap_8 FILLER_66_2119 ();
 sg13g2_decap_8 FILLER_66_2126 ();
 sg13g2_decap_8 FILLER_66_2133 ();
 sg13g2_decap_8 FILLER_66_2140 ();
 sg13g2_decap_8 FILLER_66_2147 ();
 sg13g2_decap_4 FILLER_66_2154 ();
 sg13g2_fill_1 FILLER_66_2158 ();
 sg13g2_decap_4 FILLER_66_2185 ();
 sg13g2_fill_2 FILLER_66_2189 ();
 sg13g2_decap_8 FILLER_66_2201 ();
 sg13g2_decap_8 FILLER_66_2208 ();
 sg13g2_decap_8 FILLER_66_2215 ();
 sg13g2_decap_8 FILLER_66_2222 ();
 sg13g2_decap_4 FILLER_66_2229 ();
 sg13g2_fill_1 FILLER_66_2233 ();
 sg13g2_decap_8 FILLER_66_2245 ();
 sg13g2_decap_8 FILLER_66_2252 ();
 sg13g2_decap_8 FILLER_66_2259 ();
 sg13g2_decap_8 FILLER_66_2266 ();
 sg13g2_decap_8 FILLER_66_2273 ();
 sg13g2_decap_8 FILLER_66_2280 ();
 sg13g2_decap_8 FILLER_66_2287 ();
 sg13g2_decap_8 FILLER_66_2294 ();
 sg13g2_decap_8 FILLER_66_2301 ();
 sg13g2_decap_8 FILLER_66_2308 ();
 sg13g2_decap_8 FILLER_66_2315 ();
 sg13g2_decap_8 FILLER_66_2322 ();
 sg13g2_decap_4 FILLER_66_2329 ();
 sg13g2_decap_8 FILLER_66_2338 ();
 sg13g2_decap_8 FILLER_66_2345 ();
 sg13g2_decap_8 FILLER_66_2352 ();
 sg13g2_decap_8 FILLER_66_2359 ();
 sg13g2_decap_8 FILLER_66_2366 ();
 sg13g2_decap_8 FILLER_66_2373 ();
 sg13g2_decap_8 FILLER_66_2380 ();
 sg13g2_decap_8 FILLER_66_2387 ();
 sg13g2_decap_8 FILLER_66_2420 ();
 sg13g2_decap_8 FILLER_66_2427 ();
 sg13g2_decap_4 FILLER_66_2434 ();
 sg13g2_decap_8 FILLER_66_2469 ();
 sg13g2_decap_8 FILLER_66_2476 ();
 sg13g2_decap_8 FILLER_66_2483 ();
 sg13g2_decap_8 FILLER_66_2490 ();
 sg13g2_decap_8 FILLER_66_2497 ();
 sg13g2_decap_8 FILLER_66_2504 ();
 sg13g2_fill_2 FILLER_66_2511 ();
 sg13g2_decap_8 FILLER_66_2539 ();
 sg13g2_decap_8 FILLER_66_2546 ();
 sg13g2_decap_4 FILLER_66_2553 ();
 sg13g2_fill_1 FILLER_66_2557 ();
 sg13g2_decap_4 FILLER_66_2584 ();
 sg13g2_fill_2 FILLER_66_2588 ();
 sg13g2_fill_1 FILLER_66_2600 ();
 sg13g2_decap_8 FILLER_66_2631 ();
 sg13g2_decap_8 FILLER_66_2638 ();
 sg13g2_decap_8 FILLER_66_2645 ();
 sg13g2_decap_8 FILLER_66_2652 ();
 sg13g2_decap_8 FILLER_66_2659 ();
 sg13g2_decap_4 FILLER_66_2666 ();
 sg13g2_decap_8 FILLER_66_2680 ();
 sg13g2_decap_8 FILLER_66_2687 ();
 sg13g2_decap_8 FILLER_66_2694 ();
 sg13g2_decap_8 FILLER_66_2701 ();
 sg13g2_decap_8 FILLER_66_2708 ();
 sg13g2_decap_8 FILLER_66_2715 ();
 sg13g2_decap_8 FILLER_66_2722 ();
 sg13g2_decap_8 FILLER_66_2729 ();
 sg13g2_decap_8 FILLER_66_2736 ();
 sg13g2_decap_4 FILLER_66_2743 ();
 sg13g2_fill_1 FILLER_66_2747 ();
 sg13g2_decap_8 FILLER_66_2779 ();
 sg13g2_decap_4 FILLER_66_2786 ();
 sg13g2_fill_1 FILLER_66_2800 ();
 sg13g2_decap_8 FILLER_66_2837 ();
 sg13g2_decap_8 FILLER_66_2844 ();
 sg13g2_decap_8 FILLER_66_2851 ();
 sg13g2_decap_8 FILLER_66_2858 ();
 sg13g2_decap_8 FILLER_66_2865 ();
 sg13g2_decap_8 FILLER_66_2883 ();
 sg13g2_decap_8 FILLER_66_2900 ();
 sg13g2_decap_8 FILLER_66_2907 ();
 sg13g2_fill_2 FILLER_66_2914 ();
 sg13g2_fill_1 FILLER_66_2916 ();
 sg13g2_decap_8 FILLER_66_2926 ();
 sg13g2_decap_8 FILLER_66_2933 ();
 sg13g2_decap_8 FILLER_66_2940 ();
 sg13g2_decap_8 FILLER_66_2947 ();
 sg13g2_decap_8 FILLER_66_2954 ();
 sg13g2_decap_8 FILLER_66_2961 ();
 sg13g2_decap_8 FILLER_66_2968 ();
 sg13g2_decap_8 FILLER_66_2975 ();
 sg13g2_decap_8 FILLER_66_2982 ();
 sg13g2_decap_8 FILLER_66_2989 ();
 sg13g2_decap_8 FILLER_66_2996 ();
 sg13g2_decap_8 FILLER_66_3003 ();
 sg13g2_decap_8 FILLER_66_3010 ();
 sg13g2_decap_8 FILLER_66_3017 ();
 sg13g2_decap_8 FILLER_66_3024 ();
 sg13g2_decap_8 FILLER_66_3031 ();
 sg13g2_decap_8 FILLER_66_3038 ();
 sg13g2_decap_8 FILLER_66_3045 ();
 sg13g2_decap_8 FILLER_66_3052 ();
 sg13g2_decap_8 FILLER_66_3059 ();
 sg13g2_decap_8 FILLER_66_3066 ();
 sg13g2_decap_8 FILLER_66_3073 ();
 sg13g2_decap_8 FILLER_66_3080 ();
 sg13g2_decap_8 FILLER_66_3087 ();
 sg13g2_fill_2 FILLER_66_3094 ();
 sg13g2_fill_1 FILLER_66_3096 ();
 sg13g2_decap_4 FILLER_66_3107 ();
 sg13g2_decap_8 FILLER_66_3124 ();
 sg13g2_decap_8 FILLER_66_3131 ();
 sg13g2_decap_8 FILLER_66_3138 ();
 sg13g2_fill_1 FILLER_66_3145 ();
 sg13g2_decap_8 FILLER_66_3181 ();
 sg13g2_decap_8 FILLER_66_3188 ();
 sg13g2_decap_8 FILLER_66_3231 ();
 sg13g2_decap_8 FILLER_66_3238 ();
 sg13g2_fill_2 FILLER_66_3245 ();
 sg13g2_decap_8 FILLER_66_3273 ();
 sg13g2_decap_8 FILLER_66_3280 ();
 sg13g2_decap_8 FILLER_66_3287 ();
 sg13g2_decap_8 FILLER_66_3294 ();
 sg13g2_decap_8 FILLER_66_3301 ();
 sg13g2_decap_8 FILLER_66_3308 ();
 sg13g2_decap_8 FILLER_66_3315 ();
 sg13g2_decap_8 FILLER_66_3322 ();
 sg13g2_decap_8 FILLER_66_3329 ();
 sg13g2_decap_8 FILLER_66_3336 ();
 sg13g2_decap_8 FILLER_66_3343 ();
 sg13g2_decap_4 FILLER_66_3355 ();
 sg13g2_fill_1 FILLER_66_3359 ();
 sg13g2_decap_8 FILLER_66_3381 ();
 sg13g2_decap_4 FILLER_66_3388 ();
 sg13g2_fill_2 FILLER_66_3392 ();
 sg13g2_fill_2 FILLER_66_3404 ();
 sg13g2_fill_1 FILLER_66_3406 ();
 sg13g2_fill_2 FILLER_66_3415 ();
 sg13g2_decap_4 FILLER_66_3422 ();
 sg13g2_fill_2 FILLER_66_3461 ();
 sg13g2_fill_1 FILLER_66_3463 ();
 sg13g2_decap_8 FILLER_66_3469 ();
 sg13g2_decap_4 FILLER_66_3476 ();
 sg13g2_fill_2 FILLER_66_3480 ();
 sg13g2_decap_8 FILLER_66_3524 ();
 sg13g2_decap_8 FILLER_66_3531 ();
 sg13g2_decap_8 FILLER_66_3538 ();
 sg13g2_decap_8 FILLER_66_3545 ();
 sg13g2_decap_8 FILLER_66_3552 ();
 sg13g2_decap_8 FILLER_66_3559 ();
 sg13g2_decap_8 FILLER_66_3566 ();
 sg13g2_decap_8 FILLER_66_3573 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_8 FILLER_67_7 ();
 sg13g2_fill_2 FILLER_67_14 ();
 sg13g2_fill_1 FILLER_67_16 ();
 sg13g2_fill_2 FILLER_67_39 ();
 sg13g2_fill_1 FILLER_67_41 ();
 sg13g2_decap_8 FILLER_67_51 ();
 sg13g2_decap_8 FILLER_67_58 ();
 sg13g2_decap_8 FILLER_67_65 ();
 sg13g2_decap_8 FILLER_67_72 ();
 sg13g2_decap_8 FILLER_67_79 ();
 sg13g2_decap_4 FILLER_67_86 ();
 sg13g2_fill_2 FILLER_67_90 ();
 sg13g2_decap_8 FILLER_67_96 ();
 sg13g2_decap_4 FILLER_67_103 ();
 sg13g2_decap_8 FILLER_67_115 ();
 sg13g2_decap_8 FILLER_67_122 ();
 sg13g2_fill_2 FILLER_67_129 ();
 sg13g2_fill_1 FILLER_67_131 ();
 sg13g2_decap_8 FILLER_67_140 ();
 sg13g2_decap_8 FILLER_67_147 ();
 sg13g2_decap_8 FILLER_67_154 ();
 sg13g2_decap_8 FILLER_67_161 ();
 sg13g2_decap_8 FILLER_67_168 ();
 sg13g2_decap_8 FILLER_67_175 ();
 sg13g2_decap_8 FILLER_67_182 ();
 sg13g2_fill_1 FILLER_67_189 ();
 sg13g2_decap_8 FILLER_67_214 ();
 sg13g2_decap_8 FILLER_67_221 ();
 sg13g2_decap_8 FILLER_67_228 ();
 sg13g2_fill_2 FILLER_67_235 ();
 sg13g2_fill_1 FILLER_67_237 ();
 sg13g2_fill_2 FILLER_67_246 ();
 sg13g2_decap_8 FILLER_67_253 ();
 sg13g2_decap_8 FILLER_67_260 ();
 sg13g2_decap_4 FILLER_67_267 ();
 sg13g2_fill_1 FILLER_67_277 ();
 sg13g2_fill_2 FILLER_67_289 ();
 sg13g2_fill_1 FILLER_67_291 ();
 sg13g2_decap_8 FILLER_67_300 ();
 sg13g2_decap_8 FILLER_67_307 ();
 sg13g2_decap_8 FILLER_67_314 ();
 sg13g2_fill_2 FILLER_67_321 ();
 sg13g2_fill_1 FILLER_67_323 ();
 sg13g2_decap_4 FILLER_67_341 ();
 sg13g2_fill_2 FILLER_67_345 ();
 sg13g2_decap_8 FILLER_67_356 ();
 sg13g2_decap_8 FILLER_67_368 ();
 sg13g2_decap_8 FILLER_67_375 ();
 sg13g2_decap_8 FILLER_67_382 ();
 sg13g2_decap_8 FILLER_67_389 ();
 sg13g2_decap_8 FILLER_67_396 ();
 sg13g2_decap_4 FILLER_67_403 ();
 sg13g2_fill_2 FILLER_67_407 ();
 sg13g2_decap_8 FILLER_67_414 ();
 sg13g2_decap_4 FILLER_67_421 ();
 sg13g2_fill_2 FILLER_67_425 ();
 sg13g2_decap_8 FILLER_67_432 ();
 sg13g2_decap_8 FILLER_67_439 ();
 sg13g2_decap_8 FILLER_67_446 ();
 sg13g2_fill_1 FILLER_67_453 ();
 sg13g2_decap_8 FILLER_67_494 ();
 sg13g2_decap_8 FILLER_67_501 ();
 sg13g2_decap_8 FILLER_67_508 ();
 sg13g2_decap_8 FILLER_67_515 ();
 sg13g2_decap_8 FILLER_67_522 ();
 sg13g2_decap_8 FILLER_67_529 ();
 sg13g2_fill_1 FILLER_67_541 ();
 sg13g2_fill_1 FILLER_67_547 ();
 sg13g2_fill_2 FILLER_67_558 ();
 sg13g2_decap_4 FILLER_67_568 ();
 sg13g2_fill_2 FILLER_67_572 ();
 sg13g2_fill_2 FILLER_67_579 ();
 sg13g2_fill_1 FILLER_67_581 ();
 sg13g2_decap_8 FILLER_67_587 ();
 sg13g2_decap_8 FILLER_67_594 ();
 sg13g2_decap_8 FILLER_67_601 ();
 sg13g2_decap_8 FILLER_67_608 ();
 sg13g2_decap_8 FILLER_67_615 ();
 sg13g2_decap_8 FILLER_67_622 ();
 sg13g2_decap_8 FILLER_67_629 ();
 sg13g2_decap_8 FILLER_67_636 ();
 sg13g2_decap_8 FILLER_67_643 ();
 sg13g2_decap_8 FILLER_67_650 ();
 sg13g2_decap_8 FILLER_67_657 ();
 sg13g2_decap_8 FILLER_67_664 ();
 sg13g2_decap_8 FILLER_67_671 ();
 sg13g2_fill_1 FILLER_67_683 ();
 sg13g2_decap_8 FILLER_67_692 ();
 sg13g2_decap_8 FILLER_67_699 ();
 sg13g2_decap_8 FILLER_67_706 ();
 sg13g2_decap_8 FILLER_67_713 ();
 sg13g2_decap_8 FILLER_67_720 ();
 sg13g2_decap_8 FILLER_67_727 ();
 sg13g2_decap_8 FILLER_67_734 ();
 sg13g2_fill_1 FILLER_67_741 ();
 sg13g2_decap_8 FILLER_67_773 ();
 sg13g2_decap_8 FILLER_67_780 ();
 sg13g2_decap_4 FILLER_67_787 ();
 sg13g2_fill_1 FILLER_67_791 ();
 sg13g2_decap_8 FILLER_67_812 ();
 sg13g2_decap_4 FILLER_67_819 ();
 sg13g2_fill_2 FILLER_67_823 ();
 sg13g2_decap_8 FILLER_67_833 ();
 sg13g2_decap_4 FILLER_67_840 ();
 sg13g2_fill_2 FILLER_67_844 ();
 sg13g2_fill_2 FILLER_67_860 ();
 sg13g2_fill_1 FILLER_67_870 ();
 sg13g2_fill_1 FILLER_67_879 ();
 sg13g2_decap_8 FILLER_67_885 ();
 sg13g2_decap_8 FILLER_67_892 ();
 sg13g2_decap_8 FILLER_67_899 ();
 sg13g2_decap_8 FILLER_67_906 ();
 sg13g2_decap_8 FILLER_67_913 ();
 sg13g2_decap_4 FILLER_67_920 ();
 sg13g2_decap_8 FILLER_67_929 ();
 sg13g2_decap_8 FILLER_67_936 ();
 sg13g2_decap_8 FILLER_67_943 ();
 sg13g2_decap_8 FILLER_67_950 ();
 sg13g2_fill_2 FILLER_67_957 ();
 sg13g2_decap_4 FILLER_67_962 ();
 sg13g2_fill_2 FILLER_67_966 ();
 sg13g2_decap_4 FILLER_67_977 ();
 sg13g2_fill_1 FILLER_67_981 ();
 sg13g2_fill_1 FILLER_67_1013 ();
 sg13g2_fill_1 FILLER_67_1023 ();
 sg13g2_fill_2 FILLER_67_1029 ();
 sg13g2_fill_1 FILLER_67_1031 ();
 sg13g2_decap_4 FILLER_67_1036 ();
 sg13g2_fill_1 FILLER_67_1040 ();
 sg13g2_decap_8 FILLER_67_1046 ();
 sg13g2_fill_2 FILLER_67_1053 ();
 sg13g2_fill_1 FILLER_67_1055 ();
 sg13g2_decap_8 FILLER_67_1061 ();
 sg13g2_decap_8 FILLER_67_1068 ();
 sg13g2_decap_4 FILLER_67_1075 ();
 sg13g2_fill_2 FILLER_67_1079 ();
 sg13g2_fill_2 FILLER_67_1116 ();
 sg13g2_fill_1 FILLER_67_1118 ();
 sg13g2_decap_8 FILLER_67_1151 ();
 sg13g2_fill_1 FILLER_67_1158 ();
 sg13g2_decap_8 FILLER_67_1169 ();
 sg13g2_decap_8 FILLER_67_1176 ();
 sg13g2_decap_4 FILLER_67_1183 ();
 sg13g2_fill_2 FILLER_67_1187 ();
 sg13g2_fill_2 FILLER_67_1192 ();
 sg13g2_decap_8 FILLER_67_1210 ();
 sg13g2_decap_8 FILLER_67_1217 ();
 sg13g2_decap_8 FILLER_67_1224 ();
 sg13g2_decap_4 FILLER_67_1231 ();
 sg13g2_fill_2 FILLER_67_1235 ();
 sg13g2_decap_8 FILLER_67_1272 ();
 sg13g2_decap_8 FILLER_67_1279 ();
 sg13g2_decap_8 FILLER_67_1286 ();
 sg13g2_decap_8 FILLER_67_1293 ();
 sg13g2_fill_2 FILLER_67_1300 ();
 sg13g2_decap_8 FILLER_67_1316 ();
 sg13g2_decap_8 FILLER_67_1323 ();
 sg13g2_decap_8 FILLER_67_1330 ();
 sg13g2_decap_8 FILLER_67_1337 ();
 sg13g2_decap_4 FILLER_67_1344 ();
 sg13g2_decap_8 FILLER_67_1351 ();
 sg13g2_decap_8 FILLER_67_1358 ();
 sg13g2_decap_8 FILLER_67_1365 ();
 sg13g2_fill_2 FILLER_67_1372 ();
 sg13g2_fill_1 FILLER_67_1374 ();
 sg13g2_decap_8 FILLER_67_1401 ();
 sg13g2_decap_8 FILLER_67_1408 ();
 sg13g2_decap_4 FILLER_67_1415 ();
 sg13g2_fill_1 FILLER_67_1419 ();
 sg13g2_decap_8 FILLER_67_1442 ();
 sg13g2_decap_8 FILLER_67_1449 ();
 sg13g2_decap_8 FILLER_67_1456 ();
 sg13g2_decap_8 FILLER_67_1463 ();
 sg13g2_decap_8 FILLER_67_1470 ();
 sg13g2_decap_8 FILLER_67_1477 ();
 sg13g2_decap_8 FILLER_67_1484 ();
 sg13g2_decap_8 FILLER_67_1491 ();
 sg13g2_fill_2 FILLER_67_1498 ();
 sg13g2_fill_1 FILLER_67_1500 ();
 sg13g2_decap_8 FILLER_67_1527 ();
 sg13g2_decap_8 FILLER_67_1534 ();
 sg13g2_decap_8 FILLER_67_1541 ();
 sg13g2_decap_8 FILLER_67_1548 ();
 sg13g2_decap_8 FILLER_67_1561 ();
 sg13g2_decap_8 FILLER_67_1568 ();
 sg13g2_decap_8 FILLER_67_1575 ();
 sg13g2_fill_2 FILLER_67_1582 ();
 sg13g2_fill_1 FILLER_67_1584 ();
 sg13g2_fill_1 FILLER_67_1594 ();
 sg13g2_decap_4 FILLER_67_1621 ();
 sg13g2_decap_8 FILLER_67_1637 ();
 sg13g2_decap_8 FILLER_67_1644 ();
 sg13g2_decap_8 FILLER_67_1651 ();
 sg13g2_decap_8 FILLER_67_1658 ();
 sg13g2_decap_8 FILLER_67_1697 ();
 sg13g2_decap_8 FILLER_67_1704 ();
 sg13g2_fill_1 FILLER_67_1711 ();
 sg13g2_decap_8 FILLER_67_1725 ();
 sg13g2_decap_8 FILLER_67_1732 ();
 sg13g2_decap_8 FILLER_67_1739 ();
 sg13g2_decap_8 FILLER_67_1746 ();
 sg13g2_decap_8 FILLER_67_1753 ();
 sg13g2_decap_8 FILLER_67_1760 ();
 sg13g2_decap_8 FILLER_67_1793 ();
 sg13g2_fill_2 FILLER_67_1800 ();
 sg13g2_fill_1 FILLER_67_1802 ();
 sg13g2_fill_2 FILLER_67_1813 ();
 sg13g2_decap_8 FILLER_67_1821 ();
 sg13g2_decap_8 FILLER_67_1828 ();
 sg13g2_decap_8 FILLER_67_1835 ();
 sg13g2_decap_4 FILLER_67_1842 ();
 sg13g2_fill_2 FILLER_67_1846 ();
 sg13g2_decap_4 FILLER_67_1866 ();
 sg13g2_fill_1 FILLER_67_1870 ();
 sg13g2_decap_8 FILLER_67_1876 ();
 sg13g2_decap_4 FILLER_67_1883 ();
 sg13g2_decap_8 FILLER_67_1897 ();
 sg13g2_fill_1 FILLER_67_1904 ();
 sg13g2_decap_8 FILLER_67_1913 ();
 sg13g2_decap_8 FILLER_67_1920 ();
 sg13g2_decap_8 FILLER_67_1927 ();
 sg13g2_decap_8 FILLER_67_1934 ();
 sg13g2_decap_8 FILLER_67_1941 ();
 sg13g2_decap_8 FILLER_67_1948 ();
 sg13g2_decap_8 FILLER_67_1955 ();
 sg13g2_decap_8 FILLER_67_1962 ();
 sg13g2_decap_8 FILLER_67_1969 ();
 sg13g2_decap_8 FILLER_67_1976 ();
 sg13g2_decap_8 FILLER_67_1983 ();
 sg13g2_decap_8 FILLER_67_2008 ();
 sg13g2_decap_8 FILLER_67_2015 ();
 sg13g2_decap_8 FILLER_67_2022 ();
 sg13g2_decap_8 FILLER_67_2029 ();
 sg13g2_decap_8 FILLER_67_2036 ();
 sg13g2_decap_8 FILLER_67_2043 ();
 sg13g2_decap_8 FILLER_67_2050 ();
 sg13g2_decap_8 FILLER_67_2057 ();
 sg13g2_fill_2 FILLER_67_2064 ();
 sg13g2_fill_1 FILLER_67_2066 ();
 sg13g2_decap_8 FILLER_67_2077 ();
 sg13g2_decap_8 FILLER_67_2084 ();
 sg13g2_decap_8 FILLER_67_2091 ();
 sg13g2_fill_2 FILLER_67_2098 ();
 sg13g2_decap_8 FILLER_67_2110 ();
 sg13g2_fill_1 FILLER_67_2117 ();
 sg13g2_decap_8 FILLER_67_2128 ();
 sg13g2_decap_8 FILLER_67_2135 ();
 sg13g2_decap_8 FILLER_67_2142 ();
 sg13g2_decap_8 FILLER_67_2149 ();
 sg13g2_decap_8 FILLER_67_2156 ();
 sg13g2_decap_4 FILLER_67_2163 ();
 sg13g2_decap_8 FILLER_67_2196 ();
 sg13g2_decap_8 FILLER_67_2203 ();
 sg13g2_decap_8 FILLER_67_2210 ();
 sg13g2_decap_8 FILLER_67_2217 ();
 sg13g2_decap_4 FILLER_67_2224 ();
 sg13g2_fill_1 FILLER_67_2228 ();
 sg13g2_decap_8 FILLER_67_2239 ();
 sg13g2_decap_8 FILLER_67_2246 ();
 sg13g2_decap_8 FILLER_67_2253 ();
 sg13g2_decap_8 FILLER_67_2260 ();
 sg13g2_fill_1 FILLER_67_2277 ();
 sg13g2_decap_8 FILLER_67_2308 ();
 sg13g2_decap_8 FILLER_67_2315 ();
 sg13g2_decap_8 FILLER_67_2322 ();
 sg13g2_decap_8 FILLER_67_2329 ();
 sg13g2_decap_4 FILLER_67_2336 ();
 sg13g2_fill_1 FILLER_67_2340 ();
 sg13g2_decap_8 FILLER_67_2353 ();
 sg13g2_decap_8 FILLER_67_2360 ();
 sg13g2_decap_8 FILLER_67_2367 ();
 sg13g2_decap_8 FILLER_67_2374 ();
 sg13g2_decap_8 FILLER_67_2381 ();
 sg13g2_decap_8 FILLER_67_2388 ();
 sg13g2_fill_2 FILLER_67_2395 ();
 sg13g2_fill_1 FILLER_67_2397 ();
 sg13g2_decap_8 FILLER_67_2408 ();
 sg13g2_decap_8 FILLER_67_2415 ();
 sg13g2_decap_8 FILLER_67_2422 ();
 sg13g2_decap_8 FILLER_67_2429 ();
 sg13g2_decap_8 FILLER_67_2436 ();
 sg13g2_decap_8 FILLER_67_2443 ();
 sg13g2_fill_1 FILLER_67_2450 ();
 sg13g2_decap_8 FILLER_67_2465 ();
 sg13g2_decap_8 FILLER_67_2472 ();
 sg13g2_decap_8 FILLER_67_2479 ();
 sg13g2_decap_8 FILLER_67_2486 ();
 sg13g2_decap_8 FILLER_67_2493 ();
 sg13g2_decap_8 FILLER_67_2500 ();
 sg13g2_decap_8 FILLER_67_2507 ();
 sg13g2_decap_4 FILLER_67_2514 ();
 sg13g2_decap_8 FILLER_67_2528 ();
 sg13g2_decap_8 FILLER_67_2535 ();
 sg13g2_decap_8 FILLER_67_2542 ();
 sg13g2_fill_2 FILLER_67_2549 ();
 sg13g2_fill_1 FILLER_67_2551 ();
 sg13g2_decap_8 FILLER_67_2563 ();
 sg13g2_decap_8 FILLER_67_2570 ();
 sg13g2_decap_8 FILLER_67_2577 ();
 sg13g2_decap_8 FILLER_67_2584 ();
 sg13g2_fill_1 FILLER_67_2591 ();
 sg13g2_decap_8 FILLER_67_2629 ();
 sg13g2_decap_8 FILLER_67_2636 ();
 sg13g2_decap_8 FILLER_67_2643 ();
 sg13g2_decap_8 FILLER_67_2650 ();
 sg13g2_decap_8 FILLER_67_2657 ();
 sg13g2_decap_8 FILLER_67_2664 ();
 sg13g2_decap_8 FILLER_67_2671 ();
 sg13g2_decap_8 FILLER_67_2678 ();
 sg13g2_decap_8 FILLER_67_2685 ();
 sg13g2_decap_4 FILLER_67_2692 ();
 sg13g2_fill_1 FILLER_67_2696 ();
 sg13g2_decap_8 FILLER_67_2707 ();
 sg13g2_decap_8 FILLER_67_2714 ();
 sg13g2_decap_8 FILLER_67_2736 ();
 sg13g2_decap_8 FILLER_67_2743 ();
 sg13g2_fill_2 FILLER_67_2750 ();
 sg13g2_fill_1 FILLER_67_2752 ();
 sg13g2_decap_8 FILLER_67_2757 ();
 sg13g2_decap_4 FILLER_67_2764 ();
 sg13g2_fill_2 FILLER_67_2768 ();
 sg13g2_decap_8 FILLER_67_2781 ();
 sg13g2_decap_8 FILLER_67_2788 ();
 sg13g2_decap_4 FILLER_67_2795 ();
 sg13g2_decap_8 FILLER_67_2835 ();
 sg13g2_decap_8 FILLER_67_2842 ();
 sg13g2_decap_8 FILLER_67_2849 ();
 sg13g2_decap_8 FILLER_67_2856 ();
 sg13g2_decap_4 FILLER_67_2863 ();
 sg13g2_fill_1 FILLER_67_2867 ();
 sg13g2_decap_8 FILLER_67_2879 ();
 sg13g2_decap_8 FILLER_67_2886 ();
 sg13g2_decap_8 FILLER_67_2893 ();
 sg13g2_decap_8 FILLER_67_2900 ();
 sg13g2_decap_8 FILLER_67_2907 ();
 sg13g2_decap_8 FILLER_67_2914 ();
 sg13g2_decap_8 FILLER_67_2921 ();
 sg13g2_decap_8 FILLER_67_2928 ();
 sg13g2_decap_8 FILLER_67_2938 ();
 sg13g2_fill_2 FILLER_67_2945 ();
 sg13g2_fill_1 FILLER_67_2947 ();
 sg13g2_fill_2 FILLER_67_2956 ();
 sg13g2_fill_1 FILLER_67_2958 ();
 sg13g2_decap_8 FILLER_67_2964 ();
 sg13g2_decap_8 FILLER_67_2971 ();
 sg13g2_decap_8 FILLER_67_2978 ();
 sg13g2_decap_8 FILLER_67_2985 ();
 sg13g2_decap_8 FILLER_67_2992 ();
 sg13g2_decap_8 FILLER_67_2999 ();
 sg13g2_decap_8 FILLER_67_3006 ();
 sg13g2_decap_8 FILLER_67_3013 ();
 sg13g2_decap_8 FILLER_67_3020 ();
 sg13g2_decap_8 FILLER_67_3027 ();
 sg13g2_decap_8 FILLER_67_3034 ();
 sg13g2_decap_8 FILLER_67_3041 ();
 sg13g2_decap_8 FILLER_67_3048 ();
 sg13g2_decap_8 FILLER_67_3055 ();
 sg13g2_decap_8 FILLER_67_3062 ();
 sg13g2_decap_8 FILLER_67_3069 ();
 sg13g2_decap_8 FILLER_67_3076 ();
 sg13g2_decap_8 FILLER_67_3083 ();
 sg13g2_decap_8 FILLER_67_3090 ();
 sg13g2_decap_8 FILLER_67_3097 ();
 sg13g2_decap_8 FILLER_67_3104 ();
 sg13g2_decap_8 FILLER_67_3147 ();
 sg13g2_decap_8 FILLER_67_3154 ();
 sg13g2_decap_8 FILLER_67_3161 ();
 sg13g2_decap_8 FILLER_67_3168 ();
 sg13g2_decap_4 FILLER_67_3175 ();
 sg13g2_fill_2 FILLER_67_3179 ();
 sg13g2_decap_8 FILLER_67_3186 ();
 sg13g2_decap_8 FILLER_67_3193 ();
 sg13g2_decap_8 FILLER_67_3200 ();
 sg13g2_fill_2 FILLER_67_3207 ();
 sg13g2_decap_8 FILLER_67_3219 ();
 sg13g2_decap_8 FILLER_67_3226 ();
 sg13g2_decap_8 FILLER_67_3233 ();
 sg13g2_decap_8 FILLER_67_3240 ();
 sg13g2_fill_2 FILLER_67_3247 ();
 sg13g2_fill_1 FILLER_67_3249 ();
 sg13g2_decap_8 FILLER_67_3276 ();
 sg13g2_decap_8 FILLER_67_3283 ();
 sg13g2_decap_8 FILLER_67_3290 ();
 sg13g2_decap_4 FILLER_67_3297 ();
 sg13g2_fill_2 FILLER_67_3301 ();
 sg13g2_fill_2 FILLER_67_3313 ();
 sg13g2_decap_8 FILLER_67_3320 ();
 sg13g2_decap_4 FILLER_67_3327 ();
 sg13g2_fill_2 FILLER_67_3331 ();
 sg13g2_decap_8 FILLER_67_3343 ();
 sg13g2_decap_4 FILLER_67_3350 ();
 sg13g2_fill_1 FILLER_67_3354 ();
 sg13g2_decap_8 FILLER_67_3381 ();
 sg13g2_decap_8 FILLER_67_3388 ();
 sg13g2_fill_1 FILLER_67_3395 ();
 sg13g2_decap_4 FILLER_67_3429 ();
 sg13g2_decap_8 FILLER_67_3437 ();
 sg13g2_decap_8 FILLER_67_3444 ();
 sg13g2_decap_4 FILLER_67_3451 ();
 sg13g2_decap_8 FILLER_67_3481 ();
 sg13g2_fill_1 FILLER_67_3488 ();
 sg13g2_decap_4 FILLER_67_3494 ();
 sg13g2_fill_1 FILLER_67_3498 ();
 sg13g2_decap_8 FILLER_67_3530 ();
 sg13g2_decap_8 FILLER_67_3537 ();
 sg13g2_decap_8 FILLER_67_3544 ();
 sg13g2_decap_8 FILLER_67_3551 ();
 sg13g2_decap_8 FILLER_67_3558 ();
 sg13g2_decap_8 FILLER_67_3565 ();
 sg13g2_decap_8 FILLER_67_3572 ();
 sg13g2_fill_1 FILLER_67_3579 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_8 FILLER_68_7 ();
 sg13g2_fill_2 FILLER_68_14 ();
 sg13g2_fill_1 FILLER_68_16 ();
 sg13g2_decap_8 FILLER_68_43 ();
 sg13g2_decap_8 FILLER_68_50 ();
 sg13g2_decap_8 FILLER_68_57 ();
 sg13g2_decap_8 FILLER_68_64 ();
 sg13g2_decap_8 FILLER_68_98 ();
 sg13g2_decap_8 FILLER_68_105 ();
 sg13g2_decap_8 FILLER_68_112 ();
 sg13g2_decap_8 FILLER_68_119 ();
 sg13g2_decap_8 FILLER_68_126 ();
 sg13g2_decap_8 FILLER_68_133 ();
 sg13g2_decap_8 FILLER_68_140 ();
 sg13g2_decap_8 FILLER_68_147 ();
 sg13g2_decap_4 FILLER_68_154 ();
 sg13g2_decap_8 FILLER_68_162 ();
 sg13g2_fill_2 FILLER_68_169 ();
 sg13g2_decap_4 FILLER_68_188 ();
 sg13g2_fill_1 FILLER_68_221 ();
 sg13g2_fill_2 FILLER_68_236 ();
 sg13g2_fill_1 FILLER_68_267 ();
 sg13g2_fill_2 FILLER_68_276 ();
 sg13g2_decap_8 FILLER_68_318 ();
 sg13g2_decap_8 FILLER_68_325 ();
 sg13g2_decap_8 FILLER_68_332 ();
 sg13g2_decap_8 FILLER_68_339 ();
 sg13g2_decap_8 FILLER_68_346 ();
 sg13g2_decap_8 FILLER_68_353 ();
 sg13g2_decap_8 FILLER_68_360 ();
 sg13g2_decap_8 FILLER_68_367 ();
 sg13g2_decap_8 FILLER_68_374 ();
 sg13g2_decap_8 FILLER_68_381 ();
 sg13g2_fill_1 FILLER_68_388 ();
 sg13g2_fill_2 FILLER_68_400 ();
 sg13g2_decap_8 FILLER_68_438 ();
 sg13g2_decap_4 FILLER_68_445 ();
 sg13g2_fill_2 FILLER_68_449 ();
 sg13g2_decap_8 FILLER_68_478 ();
 sg13g2_decap_8 FILLER_68_485 ();
 sg13g2_decap_8 FILLER_68_492 ();
 sg13g2_decap_8 FILLER_68_499 ();
 sg13g2_decap_4 FILLER_68_506 ();
 sg13g2_fill_2 FILLER_68_510 ();
 sg13g2_decap_8 FILLER_68_517 ();
 sg13g2_fill_2 FILLER_68_524 ();
 sg13g2_fill_1 FILLER_68_526 ();
 sg13g2_fill_2 FILLER_68_542 ();
 sg13g2_fill_1 FILLER_68_544 ();
 sg13g2_decap_8 FILLER_68_578 ();
 sg13g2_decap_8 FILLER_68_585 ();
 sg13g2_decap_8 FILLER_68_592 ();
 sg13g2_decap_8 FILLER_68_599 ();
 sg13g2_decap_8 FILLER_68_606 ();
 sg13g2_decap_8 FILLER_68_613 ();
 sg13g2_decap_8 FILLER_68_620 ();
 sg13g2_decap_8 FILLER_68_640 ();
 sg13g2_decap_8 FILLER_68_647 ();
 sg13g2_decap_8 FILLER_68_654 ();
 sg13g2_fill_2 FILLER_68_661 ();
 sg13g2_fill_1 FILLER_68_663 ();
 sg13g2_fill_2 FILLER_68_672 ();
 sg13g2_fill_1 FILLER_68_674 ();
 sg13g2_decap_8 FILLER_68_698 ();
 sg13g2_fill_2 FILLER_68_705 ();
 sg13g2_decap_8 FILLER_68_711 ();
 sg13g2_decap_4 FILLER_68_718 ();
 sg13g2_fill_1 FILLER_68_727 ();
 sg13g2_decap_8 FILLER_68_736 ();
 sg13g2_decap_8 FILLER_68_743 ();
 sg13g2_decap_8 FILLER_68_750 ();
 sg13g2_decap_8 FILLER_68_757 ();
 sg13g2_decap_8 FILLER_68_764 ();
 sg13g2_decap_8 FILLER_68_771 ();
 sg13g2_decap_4 FILLER_68_778 ();
 sg13g2_decap_8 FILLER_68_807 ();
 sg13g2_decap_8 FILLER_68_814 ();
 sg13g2_decap_8 FILLER_68_821 ();
 sg13g2_decap_8 FILLER_68_828 ();
 sg13g2_decap_8 FILLER_68_835 ();
 sg13g2_decap_8 FILLER_68_842 ();
 sg13g2_fill_2 FILLER_68_849 ();
 sg13g2_fill_2 FILLER_68_865 ();
 sg13g2_fill_1 FILLER_68_867 ();
 sg13g2_decap_4 FILLER_68_875 ();
 sg13g2_fill_2 FILLER_68_889 ();
 sg13g2_decap_8 FILLER_68_908 ();
 sg13g2_decap_8 FILLER_68_915 ();
 sg13g2_decap_8 FILLER_68_945 ();
 sg13g2_decap_8 FILLER_68_952 ();
 sg13g2_decap_8 FILLER_68_959 ();
 sg13g2_fill_2 FILLER_68_966 ();
 sg13g2_fill_1 FILLER_68_968 ();
 sg13g2_fill_2 FILLER_68_982 ();
 sg13g2_fill_1 FILLER_68_984 ();
 sg13g2_fill_1 FILLER_68_992 ();
 sg13g2_decap_8 FILLER_68_996 ();
 sg13g2_decap_8 FILLER_68_1003 ();
 sg13g2_decap_8 FILLER_68_1010 ();
 sg13g2_decap_8 FILLER_68_1017 ();
 sg13g2_decap_8 FILLER_68_1024 ();
 sg13g2_decap_4 FILLER_68_1031 ();
 sg13g2_fill_2 FILLER_68_1035 ();
 sg13g2_fill_1 FILLER_68_1044 ();
 sg13g2_fill_2 FILLER_68_1050 ();
 sg13g2_fill_2 FILLER_68_1064 ();
 sg13g2_decap_8 FILLER_68_1072 ();
 sg13g2_decap_8 FILLER_68_1079 ();
 sg13g2_fill_2 FILLER_68_1086 ();
 sg13g2_decap_8 FILLER_68_1119 ();
 sg13g2_decap_8 FILLER_68_1126 ();
 sg13g2_decap_8 FILLER_68_1133 ();
 sg13g2_decap_8 FILLER_68_1140 ();
 sg13g2_decap_8 FILLER_68_1147 ();
 sg13g2_decap_8 FILLER_68_1154 ();
 sg13g2_decap_8 FILLER_68_1161 ();
 sg13g2_decap_8 FILLER_68_1168 ();
 sg13g2_decap_8 FILLER_68_1175 ();
 sg13g2_decap_8 FILLER_68_1182 ();
 sg13g2_decap_8 FILLER_68_1220 ();
 sg13g2_decap_8 FILLER_68_1227 ();
 sg13g2_fill_2 FILLER_68_1234 ();
 sg13g2_fill_1 FILLER_68_1236 ();
 sg13g2_decap_8 FILLER_68_1240 ();
 sg13g2_decap_4 FILLER_68_1247 ();
 sg13g2_fill_2 FILLER_68_1251 ();
 sg13g2_fill_2 FILLER_68_1259 ();
 sg13g2_fill_2 FILLER_68_1264 ();
 sg13g2_decap_8 FILLER_68_1274 ();
 sg13g2_decap_8 FILLER_68_1281 ();
 sg13g2_decap_8 FILLER_68_1288 ();
 sg13g2_decap_8 FILLER_68_1295 ();
 sg13g2_fill_2 FILLER_68_1302 ();
 sg13g2_fill_1 FILLER_68_1304 ();
 sg13g2_decap_8 FILLER_68_1317 ();
 sg13g2_decap_8 FILLER_68_1324 ();
 sg13g2_decap_8 FILLER_68_1331 ();
 sg13g2_decap_8 FILLER_68_1338 ();
 sg13g2_decap_8 FILLER_68_1345 ();
 sg13g2_decap_8 FILLER_68_1352 ();
 sg13g2_decap_8 FILLER_68_1359 ();
 sg13g2_decap_8 FILLER_68_1366 ();
 sg13g2_decap_4 FILLER_68_1373 ();
 sg13g2_decap_8 FILLER_68_1387 ();
 sg13g2_decap_8 FILLER_68_1394 ();
 sg13g2_decap_8 FILLER_68_1401 ();
 sg13g2_decap_8 FILLER_68_1408 ();
 sg13g2_fill_2 FILLER_68_1415 ();
 sg13g2_fill_1 FILLER_68_1417 ();
 sg13g2_fill_2 FILLER_68_1424 ();
 sg13g2_decap_8 FILLER_68_1432 ();
 sg13g2_decap_8 FILLER_68_1439 ();
 sg13g2_decap_8 FILLER_68_1446 ();
 sg13g2_decap_8 FILLER_68_1453 ();
 sg13g2_decap_8 FILLER_68_1460 ();
 sg13g2_decap_8 FILLER_68_1467 ();
 sg13g2_decap_8 FILLER_68_1479 ();
 sg13g2_decap_8 FILLER_68_1486 ();
 sg13g2_decap_8 FILLER_68_1493 ();
 sg13g2_decap_8 FILLER_68_1500 ();
 sg13g2_decap_8 FILLER_68_1507 ();
 sg13g2_decap_8 FILLER_68_1514 ();
 sg13g2_decap_8 FILLER_68_1521 ();
 sg13g2_decap_8 FILLER_68_1528 ();
 sg13g2_decap_8 FILLER_68_1535 ();
 sg13g2_decap_8 FILLER_68_1542 ();
 sg13g2_decap_8 FILLER_68_1549 ();
 sg13g2_decap_8 FILLER_68_1556 ();
 sg13g2_decap_8 FILLER_68_1563 ();
 sg13g2_decap_8 FILLER_68_1570 ();
 sg13g2_decap_8 FILLER_68_1577 ();
 sg13g2_decap_8 FILLER_68_1584 ();
 sg13g2_decap_8 FILLER_68_1591 ();
 sg13g2_decap_8 FILLER_68_1598 ();
 sg13g2_fill_2 FILLER_68_1605 ();
 sg13g2_fill_1 FILLER_68_1607 ();
 sg13g2_decap_8 FILLER_68_1642 ();
 sg13g2_decap_8 FILLER_68_1649 ();
 sg13g2_decap_4 FILLER_68_1656 ();
 sg13g2_decap_8 FILLER_68_1699 ();
 sg13g2_decap_8 FILLER_68_1706 ();
 sg13g2_decap_8 FILLER_68_1713 ();
 sg13g2_decap_4 FILLER_68_1720 ();
 sg13g2_fill_2 FILLER_68_1724 ();
 sg13g2_decap_8 FILLER_68_1739 ();
 sg13g2_decap_8 FILLER_68_1746 ();
 sg13g2_decap_8 FILLER_68_1753 ();
 sg13g2_decap_8 FILLER_68_1760 ();
 sg13g2_decap_4 FILLER_68_1767 ();
 sg13g2_fill_1 FILLER_68_1771 ();
 sg13g2_decap_8 FILLER_68_1782 ();
 sg13g2_decap_8 FILLER_68_1789 ();
 sg13g2_decap_8 FILLER_68_1796 ();
 sg13g2_decap_8 FILLER_68_1803 ();
 sg13g2_decap_8 FILLER_68_1810 ();
 sg13g2_fill_1 FILLER_68_1817 ();
 sg13g2_decap_8 FILLER_68_1822 ();
 sg13g2_decap_4 FILLER_68_1829 ();
 sg13g2_fill_2 FILLER_68_1837 ();
 sg13g2_decap_8 FILLER_68_1843 ();
 sg13g2_decap_8 FILLER_68_1850 ();
 sg13g2_decap_8 FILLER_68_1857 ();
 sg13g2_decap_8 FILLER_68_1864 ();
 sg13g2_decap_8 FILLER_68_1871 ();
 sg13g2_decap_8 FILLER_68_1878 ();
 sg13g2_fill_2 FILLER_68_1885 ();
 sg13g2_fill_1 FILLER_68_1887 ();
 sg13g2_decap_4 FILLER_68_1914 ();
 sg13g2_fill_1 FILLER_68_1918 ();
 sg13g2_fill_1 FILLER_68_1929 ();
 sg13g2_decap_8 FILLER_68_1956 ();
 sg13g2_decap_8 FILLER_68_1963 ();
 sg13g2_decap_8 FILLER_68_1970 ();
 sg13g2_decap_4 FILLER_68_1977 ();
 sg13g2_decap_8 FILLER_68_2007 ();
 sg13g2_decap_8 FILLER_68_2014 ();
 sg13g2_decap_8 FILLER_68_2021 ();
 sg13g2_decap_8 FILLER_68_2028 ();
 sg13g2_decap_8 FILLER_68_2035 ();
 sg13g2_fill_2 FILLER_68_2042 ();
 sg13g2_fill_1 FILLER_68_2044 ();
 sg13g2_decap_8 FILLER_68_2053 ();
 sg13g2_decap_4 FILLER_68_2060 ();
 sg13g2_fill_2 FILLER_68_2064 ();
 sg13g2_decap_4 FILLER_68_2102 ();
 sg13g2_fill_1 FILLER_68_2106 ();
 sg13g2_decap_8 FILLER_68_2133 ();
 sg13g2_decap_8 FILLER_68_2140 ();
 sg13g2_decap_8 FILLER_68_2147 ();
 sg13g2_decap_8 FILLER_68_2154 ();
 sg13g2_decap_8 FILLER_68_2169 ();
 sg13g2_decap_8 FILLER_68_2176 ();
 sg13g2_decap_8 FILLER_68_2183 ();
 sg13g2_fill_2 FILLER_68_2190 ();
 sg13g2_fill_1 FILLER_68_2192 ();
 sg13g2_decap_8 FILLER_68_2204 ();
 sg13g2_decap_4 FILLER_68_2211 ();
 sg13g2_decap_8 FILLER_68_2251 ();
 sg13g2_fill_2 FILLER_68_2258 ();
 sg13g2_fill_1 FILLER_68_2260 ();
 sg13g2_decap_8 FILLER_68_2307 ();
 sg13g2_decap_8 FILLER_68_2314 ();
 sg13g2_decap_8 FILLER_68_2321 ();
 sg13g2_decap_8 FILLER_68_2328 ();
 sg13g2_fill_1 FILLER_68_2344 ();
 sg13g2_decap_8 FILLER_68_2364 ();
 sg13g2_decap_8 FILLER_68_2371 ();
 sg13g2_decap_8 FILLER_68_2378 ();
 sg13g2_decap_8 FILLER_68_2396 ();
 sg13g2_decap_8 FILLER_68_2403 ();
 sg13g2_decap_8 FILLER_68_2410 ();
 sg13g2_decap_8 FILLER_68_2417 ();
 sg13g2_decap_8 FILLER_68_2424 ();
 sg13g2_decap_8 FILLER_68_2431 ();
 sg13g2_decap_8 FILLER_68_2438 ();
 sg13g2_decap_8 FILLER_68_2445 ();
 sg13g2_decap_4 FILLER_68_2452 ();
 sg13g2_fill_1 FILLER_68_2456 ();
 sg13g2_decap_8 FILLER_68_2464 ();
 sg13g2_decap_8 FILLER_68_2471 ();
 sg13g2_decap_8 FILLER_68_2478 ();
 sg13g2_decap_8 FILLER_68_2485 ();
 sg13g2_decap_8 FILLER_68_2492 ();
 sg13g2_decap_8 FILLER_68_2499 ();
 sg13g2_decap_8 FILLER_68_2506 ();
 sg13g2_decap_8 FILLER_68_2513 ();
 sg13g2_decap_8 FILLER_68_2520 ();
 sg13g2_decap_8 FILLER_68_2527 ();
 sg13g2_decap_8 FILLER_68_2534 ();
 sg13g2_decap_8 FILLER_68_2541 ();
 sg13g2_decap_8 FILLER_68_2548 ();
 sg13g2_decap_8 FILLER_68_2555 ();
 sg13g2_decap_8 FILLER_68_2562 ();
 sg13g2_decap_8 FILLER_68_2569 ();
 sg13g2_decap_8 FILLER_68_2576 ();
 sg13g2_decap_8 FILLER_68_2583 ();
 sg13g2_decap_8 FILLER_68_2590 ();
 sg13g2_decap_8 FILLER_68_2597 ();
 sg13g2_decap_8 FILLER_68_2604 ();
 sg13g2_decap_8 FILLER_68_2611 ();
 sg13g2_decap_8 FILLER_68_2618 ();
 sg13g2_decap_8 FILLER_68_2625 ();
 sg13g2_decap_8 FILLER_68_2632 ();
 sg13g2_decap_8 FILLER_68_2639 ();
 sg13g2_fill_2 FILLER_68_2646 ();
 sg13g2_fill_1 FILLER_68_2648 ();
 sg13g2_decap_8 FILLER_68_2673 ();
 sg13g2_decap_4 FILLER_68_2680 ();
 sg13g2_fill_1 FILLER_68_2684 ();
 sg13g2_decap_8 FILLER_68_2744 ();
 sg13g2_decap_8 FILLER_68_2751 ();
 sg13g2_fill_2 FILLER_68_2758 ();
 sg13g2_decap_8 FILLER_68_2782 ();
 sg13g2_decap_8 FILLER_68_2789 ();
 sg13g2_decap_8 FILLER_68_2796 ();
 sg13g2_decap_8 FILLER_68_2803 ();
 sg13g2_decap_8 FILLER_68_2810 ();
 sg13g2_decap_8 FILLER_68_2817 ();
 sg13g2_decap_8 FILLER_68_2824 ();
 sg13g2_decap_8 FILLER_68_2831 ();
 sg13g2_decap_8 FILLER_68_2838 ();
 sg13g2_decap_8 FILLER_68_2845 ();
 sg13g2_decap_8 FILLER_68_2852 ();
 sg13g2_decap_8 FILLER_68_2859 ();
 sg13g2_decap_8 FILLER_68_2866 ();
 sg13g2_decap_8 FILLER_68_2873 ();
 sg13g2_decap_8 FILLER_68_2880 ();
 sg13g2_decap_8 FILLER_68_2887 ();
 sg13g2_decap_8 FILLER_68_2894 ();
 sg13g2_decap_8 FILLER_68_2901 ();
 sg13g2_decap_8 FILLER_68_2908 ();
 sg13g2_decap_8 FILLER_68_2915 ();
 sg13g2_decap_8 FILLER_68_2922 ();
 sg13g2_decap_8 FILLER_68_2929 ();
 sg13g2_fill_1 FILLER_68_2936 ();
 sg13g2_decap_8 FILLER_68_2974 ();
 sg13g2_decap_8 FILLER_68_2981 ();
 sg13g2_decap_8 FILLER_68_2988 ();
 sg13g2_decap_4 FILLER_68_2995 ();
 sg13g2_fill_2 FILLER_68_2999 ();
 sg13g2_decap_8 FILLER_68_3015 ();
 sg13g2_decap_8 FILLER_68_3022 ();
 sg13g2_decap_8 FILLER_68_3029 ();
 sg13g2_fill_2 FILLER_68_3036 ();
 sg13g2_decap_8 FILLER_68_3048 ();
 sg13g2_decap_8 FILLER_68_3055 ();
 sg13g2_decap_8 FILLER_68_3062 ();
 sg13g2_decap_8 FILLER_68_3069 ();
 sg13g2_fill_2 FILLER_68_3076 ();
 sg13g2_decap_8 FILLER_68_3083 ();
 sg13g2_decap_8 FILLER_68_3090 ();
 sg13g2_decap_8 FILLER_68_3097 ();
 sg13g2_decap_8 FILLER_68_3104 ();
 sg13g2_decap_8 FILLER_68_3114 ();
 sg13g2_decap_8 FILLER_68_3121 ();
 sg13g2_decap_4 FILLER_68_3128 ();
 sg13g2_fill_1 FILLER_68_3132 ();
 sg13g2_decap_4 FILLER_68_3142 ();
 sg13g2_fill_2 FILLER_68_3146 ();
 sg13g2_decap_8 FILLER_68_3174 ();
 sg13g2_decap_8 FILLER_68_3181 ();
 sg13g2_fill_2 FILLER_68_3188 ();
 sg13g2_decap_8 FILLER_68_3194 ();
 sg13g2_decap_8 FILLER_68_3201 ();
 sg13g2_decap_8 FILLER_68_3208 ();
 sg13g2_decap_8 FILLER_68_3215 ();
 sg13g2_decap_8 FILLER_68_3222 ();
 sg13g2_decap_8 FILLER_68_3229 ();
 sg13g2_decap_8 FILLER_68_3236 ();
 sg13g2_decap_8 FILLER_68_3243 ();
 sg13g2_decap_8 FILLER_68_3250 ();
 sg13g2_fill_1 FILLER_68_3257 ();
 sg13g2_decap_8 FILLER_68_3268 ();
 sg13g2_decap_8 FILLER_68_3275 ();
 sg13g2_decap_8 FILLER_68_3282 ();
 sg13g2_decap_4 FILLER_68_3289 ();
 sg13g2_decap_8 FILLER_68_3350 ();
 sg13g2_decap_8 FILLER_68_3357 ();
 sg13g2_decap_8 FILLER_68_3364 ();
 sg13g2_decap_8 FILLER_68_3371 ();
 sg13g2_decap_4 FILLER_68_3378 ();
 sg13g2_fill_1 FILLER_68_3382 ();
 sg13g2_decap_4 FILLER_68_3388 ();
 sg13g2_fill_2 FILLER_68_3392 ();
 sg13g2_fill_1 FILLER_68_3404 ();
 sg13g2_decap_8 FILLER_68_3419 ();
 sg13g2_decap_8 FILLER_68_3426 ();
 sg13g2_decap_8 FILLER_68_3433 ();
 sg13g2_decap_8 FILLER_68_3440 ();
 sg13g2_decap_4 FILLER_68_3447 ();
 sg13g2_fill_1 FILLER_68_3451 ();
 sg13g2_decap_8 FILLER_68_3471 ();
 sg13g2_decap_8 FILLER_68_3478 ();
 sg13g2_decap_8 FILLER_68_3485 ();
 sg13g2_decap_8 FILLER_68_3492 ();
 sg13g2_decap_8 FILLER_68_3499 ();
 sg13g2_decap_8 FILLER_68_3506 ();
 sg13g2_decap_4 FILLER_68_3513 ();
 sg13g2_fill_1 FILLER_68_3517 ();
 sg13g2_decap_4 FILLER_68_3521 ();
 sg13g2_decap_8 FILLER_68_3534 ();
 sg13g2_decap_8 FILLER_68_3541 ();
 sg13g2_decap_8 FILLER_68_3548 ();
 sg13g2_decap_8 FILLER_68_3555 ();
 sg13g2_decap_8 FILLER_68_3562 ();
 sg13g2_decap_8 FILLER_68_3569 ();
 sg13g2_decap_4 FILLER_68_3576 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_8 FILLER_69_7 ();
 sg13g2_decap_8 FILLER_69_14 ();
 sg13g2_decap_8 FILLER_69_26 ();
 sg13g2_decap_8 FILLER_69_33 ();
 sg13g2_decap_8 FILLER_69_40 ();
 sg13g2_decap_8 FILLER_69_47 ();
 sg13g2_decap_4 FILLER_69_80 ();
 sg13g2_fill_1 FILLER_69_84 ();
 sg13g2_decap_8 FILLER_69_101 ();
 sg13g2_decap_8 FILLER_69_108 ();
 sg13g2_decap_4 FILLER_69_115 ();
 sg13g2_fill_2 FILLER_69_119 ();
 sg13g2_fill_1 FILLER_69_147 ();
 sg13g2_decap_4 FILLER_69_157 ();
 sg13g2_decap_8 FILLER_69_179 ();
 sg13g2_decap_8 FILLER_69_186 ();
 sg13g2_decap_8 FILLER_69_193 ();
 sg13g2_decap_4 FILLER_69_200 ();
 sg13g2_fill_1 FILLER_69_204 ();
 sg13g2_decap_4 FILLER_69_217 ();
 sg13g2_fill_1 FILLER_69_234 ();
 sg13g2_decap_8 FILLER_69_251 ();
 sg13g2_decap_8 FILLER_69_258 ();
 sg13g2_decap_4 FILLER_69_265 ();
 sg13g2_fill_1 FILLER_69_269 ();
 sg13g2_decap_8 FILLER_69_277 ();
 sg13g2_decap_4 FILLER_69_284 ();
 sg13g2_fill_2 FILLER_69_292 ();
 sg13g2_decap_8 FILLER_69_297 ();
 sg13g2_decap_8 FILLER_69_304 ();
 sg13g2_decap_8 FILLER_69_311 ();
 sg13g2_decap_8 FILLER_69_318 ();
 sg13g2_decap_8 FILLER_69_325 ();
 sg13g2_decap_8 FILLER_69_332 ();
 sg13g2_decap_8 FILLER_69_339 ();
 sg13g2_decap_8 FILLER_69_346 ();
 sg13g2_fill_2 FILLER_69_353 ();
 sg13g2_fill_1 FILLER_69_355 ();
 sg13g2_decap_8 FILLER_69_371 ();
 sg13g2_decap_4 FILLER_69_378 ();
 sg13g2_decap_8 FILLER_69_413 ();
 sg13g2_decap_8 FILLER_69_420 ();
 sg13g2_decap_4 FILLER_69_427 ();
 sg13g2_decap_8 FILLER_69_439 ();
 sg13g2_decap_8 FILLER_69_446 ();
 sg13g2_decap_4 FILLER_69_453 ();
 sg13g2_fill_1 FILLER_69_462 ();
 sg13g2_decap_8 FILLER_69_475 ();
 sg13g2_decap_8 FILLER_69_482 ();
 sg13g2_fill_2 FILLER_69_489 ();
 sg13g2_decap_4 FILLER_69_496 ();
 sg13g2_fill_2 FILLER_69_500 ();
 sg13g2_decap_8 FILLER_69_507 ();
 sg13g2_decap_8 FILLER_69_514 ();
 sg13g2_decap_8 FILLER_69_521 ();
 sg13g2_fill_2 FILLER_69_528 ();
 sg13g2_fill_1 FILLER_69_530 ();
 sg13g2_decap_4 FILLER_69_559 ();
 sg13g2_decap_8 FILLER_69_568 ();
 sg13g2_decap_8 FILLER_69_575 ();
 sg13g2_decap_8 FILLER_69_582 ();
 sg13g2_decap_4 FILLER_69_589 ();
 sg13g2_fill_1 FILLER_69_593 ();
 sg13g2_decap_8 FILLER_69_612 ();
 sg13g2_decap_8 FILLER_69_619 ();
 sg13g2_fill_2 FILLER_69_626 ();
 sg13g2_decap_4 FILLER_69_633 ();
 sg13g2_fill_2 FILLER_69_637 ();
 sg13g2_fill_2 FILLER_69_644 ();
 sg13g2_fill_1 FILLER_69_646 ();
 sg13g2_decap_8 FILLER_69_663 ();
 sg13g2_decap_4 FILLER_69_670 ();
 sg13g2_fill_2 FILLER_69_674 ();
 sg13g2_decap_8 FILLER_69_703 ();
 sg13g2_decap_8 FILLER_69_710 ();
 sg13g2_decap_8 FILLER_69_737 ();
 sg13g2_decap_8 FILLER_69_744 ();
 sg13g2_decap_8 FILLER_69_751 ();
 sg13g2_decap_8 FILLER_69_758 ();
 sg13g2_decap_8 FILLER_69_765 ();
 sg13g2_decap_8 FILLER_69_772 ();
 sg13g2_decap_8 FILLER_69_779 ();
 sg13g2_fill_2 FILLER_69_786 ();
 sg13g2_fill_1 FILLER_69_788 ();
 sg13g2_fill_1 FILLER_69_803 ();
 sg13g2_decap_8 FILLER_69_817 ();
 sg13g2_decap_8 FILLER_69_824 ();
 sg13g2_decap_8 FILLER_69_831 ();
 sg13g2_decap_8 FILLER_69_838 ();
 sg13g2_decap_8 FILLER_69_845 ();
 sg13g2_decap_8 FILLER_69_852 ();
 sg13g2_decap_8 FILLER_69_879 ();
 sg13g2_decap_8 FILLER_69_886 ();
 sg13g2_decap_8 FILLER_69_893 ();
 sg13g2_decap_8 FILLER_69_900 ();
 sg13g2_decap_8 FILLER_69_907 ();
 sg13g2_decap_8 FILLER_69_914 ();
 sg13g2_fill_2 FILLER_69_921 ();
 sg13g2_decap_8 FILLER_69_963 ();
 sg13g2_decap_8 FILLER_69_970 ();
 sg13g2_decap_4 FILLER_69_977 ();
 sg13g2_decap_8 FILLER_69_985 ();
 sg13g2_decap_8 FILLER_69_992 ();
 sg13g2_decap_8 FILLER_69_999 ();
 sg13g2_decap_8 FILLER_69_1006 ();
 sg13g2_decap_8 FILLER_69_1013 ();
 sg13g2_decap_8 FILLER_69_1020 ();
 sg13g2_decap_8 FILLER_69_1027 ();
 sg13g2_decap_4 FILLER_69_1034 ();
 sg13g2_fill_1 FILLER_69_1038 ();
 sg13g2_decap_8 FILLER_69_1051 ();
 sg13g2_decap_8 FILLER_69_1058 ();
 sg13g2_decap_8 FILLER_69_1065 ();
 sg13g2_decap_8 FILLER_69_1072 ();
 sg13g2_decap_8 FILLER_69_1079 ();
 sg13g2_decap_8 FILLER_69_1086 ();
 sg13g2_decap_4 FILLER_69_1093 ();
 sg13g2_fill_2 FILLER_69_1097 ();
 sg13g2_fill_1 FILLER_69_1107 ();
 sg13g2_fill_1 FILLER_69_1123 ();
 sg13g2_decap_8 FILLER_69_1139 ();
 sg13g2_decap_8 FILLER_69_1146 ();
 sg13g2_decap_4 FILLER_69_1153 ();
 sg13g2_fill_2 FILLER_69_1157 ();
 sg13g2_decap_8 FILLER_69_1162 ();
 sg13g2_decap_8 FILLER_69_1169 ();
 sg13g2_decap_8 FILLER_69_1176 ();
 sg13g2_decap_4 FILLER_69_1183 ();
 sg13g2_fill_2 FILLER_69_1187 ();
 sg13g2_decap_8 FILLER_69_1223 ();
 sg13g2_decap_8 FILLER_69_1230 ();
 sg13g2_decap_8 FILLER_69_1240 ();
 sg13g2_decap_8 FILLER_69_1247 ();
 sg13g2_decap_8 FILLER_69_1254 ();
 sg13g2_decap_4 FILLER_69_1261 ();
 sg13g2_fill_1 FILLER_69_1265 ();
 sg13g2_decap_4 FILLER_69_1287 ();
 sg13g2_fill_1 FILLER_69_1291 ();
 sg13g2_decap_8 FILLER_69_1308 ();
 sg13g2_decap_4 FILLER_69_1329 ();
 sg13g2_decap_4 FILLER_69_1342 ();
 sg13g2_fill_1 FILLER_69_1346 ();
 sg13g2_decap_8 FILLER_69_1359 ();
 sg13g2_decap_8 FILLER_69_1366 ();
 sg13g2_decap_8 FILLER_69_1373 ();
 sg13g2_decap_8 FILLER_69_1380 ();
 sg13g2_decap_8 FILLER_69_1387 ();
 sg13g2_decap_8 FILLER_69_1394 ();
 sg13g2_decap_8 FILLER_69_1401 ();
 sg13g2_fill_1 FILLER_69_1408 ();
 sg13g2_decap_8 FILLER_69_1427 ();
 sg13g2_decap_8 FILLER_69_1434 ();
 sg13g2_decap_8 FILLER_69_1441 ();
 sg13g2_decap_8 FILLER_69_1448 ();
 sg13g2_decap_8 FILLER_69_1455 ();
 sg13g2_decap_4 FILLER_69_1462 ();
 sg13g2_decap_8 FILLER_69_1489 ();
 sg13g2_decap_8 FILLER_69_1496 ();
 sg13g2_decap_4 FILLER_69_1503 ();
 sg13g2_decap_8 FILLER_69_1513 ();
 sg13g2_decap_8 FILLER_69_1520 ();
 sg13g2_decap_8 FILLER_69_1527 ();
 sg13g2_decap_8 FILLER_69_1534 ();
 sg13g2_decap_8 FILLER_69_1551 ();
 sg13g2_decap_8 FILLER_69_1558 ();
 sg13g2_decap_8 FILLER_69_1565 ();
 sg13g2_fill_2 FILLER_69_1572 ();
 sg13g2_fill_1 FILLER_69_1574 ();
 sg13g2_decap_8 FILLER_69_1581 ();
 sg13g2_decap_8 FILLER_69_1591 ();
 sg13g2_decap_8 FILLER_69_1598 ();
 sg13g2_decap_8 FILLER_69_1605 ();
 sg13g2_decap_8 FILLER_69_1612 ();
 sg13g2_decap_4 FILLER_69_1624 ();
 sg13g2_decap_8 FILLER_69_1631 ();
 sg13g2_decap_8 FILLER_69_1638 ();
 sg13g2_decap_8 FILLER_69_1645 ();
 sg13g2_decap_8 FILLER_69_1652 ();
 sg13g2_decap_8 FILLER_69_1659 ();
 sg13g2_decap_4 FILLER_69_1666 ();
 sg13g2_fill_2 FILLER_69_1670 ();
 sg13g2_decap_8 FILLER_69_1677 ();
 sg13g2_decap_8 FILLER_69_1697 ();
 sg13g2_decap_8 FILLER_69_1704 ();
 sg13g2_decap_8 FILLER_69_1711 ();
 sg13g2_fill_2 FILLER_69_1718 ();
 sg13g2_decap_8 FILLER_69_1746 ();
 sg13g2_decap_8 FILLER_69_1753 ();
 sg13g2_decap_8 FILLER_69_1760 ();
 sg13g2_fill_2 FILLER_69_1767 ();
 sg13g2_decap_8 FILLER_69_1777 ();
 sg13g2_decap_8 FILLER_69_1784 ();
 sg13g2_decap_8 FILLER_69_1791 ();
 sg13g2_decap_8 FILLER_69_1798 ();
 sg13g2_decap_4 FILLER_69_1805 ();
 sg13g2_fill_2 FILLER_69_1809 ();
 sg13g2_decap_4 FILLER_69_1820 ();
 sg13g2_fill_1 FILLER_69_1824 ();
 sg13g2_fill_1 FILLER_69_1828 ();
 sg13g2_decap_4 FILLER_69_1865 ();
 sg13g2_fill_2 FILLER_69_1869 ();
 sg13g2_decap_8 FILLER_69_1881 ();
 sg13g2_decap_8 FILLER_69_1888 ();
 sg13g2_decap_8 FILLER_69_1895 ();
 sg13g2_decap_8 FILLER_69_1902 ();
 sg13g2_decap_8 FILLER_69_1909 ();
 sg13g2_decap_8 FILLER_69_1916 ();
 sg13g2_fill_2 FILLER_69_1923 ();
 sg13g2_fill_1 FILLER_69_1925 ();
 sg13g2_decap_8 FILLER_69_1952 ();
 sg13g2_decap_8 FILLER_69_1959 ();
 sg13g2_decap_4 FILLER_69_1966 ();
 sg13g2_fill_1 FILLER_69_1970 ();
 sg13g2_decap_8 FILLER_69_2007 ();
 sg13g2_decap_4 FILLER_69_2014 ();
 sg13g2_fill_2 FILLER_69_2018 ();
 sg13g2_fill_2 FILLER_69_2030 ();
 sg13g2_decap_8 FILLER_69_2063 ();
 sg13g2_decap_8 FILLER_69_2070 ();
 sg13g2_decap_4 FILLER_69_2077 ();
 sg13g2_decap_4 FILLER_69_2117 ();
 sg13g2_decap_4 FILLER_69_2147 ();
 sg13g2_fill_2 FILLER_69_2151 ();
 sg13g2_decap_4 FILLER_69_2189 ();
 sg13g2_decap_8 FILLER_69_2196 ();
 sg13g2_decap_8 FILLER_69_2203 ();
 sg13g2_decap_8 FILLER_69_2210 ();
 sg13g2_decap_4 FILLER_69_2217 ();
 sg13g2_decap_8 FILLER_69_2247 ();
 sg13g2_decap_8 FILLER_69_2254 ();
 sg13g2_decap_8 FILLER_69_2261 ();
 sg13g2_fill_2 FILLER_69_2268 ();
 sg13g2_fill_1 FILLER_69_2270 ();
 sg13g2_decap_8 FILLER_69_2297 ();
 sg13g2_decap_8 FILLER_69_2304 ();
 sg13g2_decap_8 FILLER_69_2311 ();
 sg13g2_decap_8 FILLER_69_2318 ();
 sg13g2_fill_1 FILLER_69_2325 ();
 sg13g2_decap_8 FILLER_69_2368 ();
 sg13g2_decap_8 FILLER_69_2375 ();
 sg13g2_decap_8 FILLER_69_2382 ();
 sg13g2_decap_8 FILLER_69_2389 ();
 sg13g2_decap_4 FILLER_69_2396 ();
 sg13g2_fill_2 FILLER_69_2400 ();
 sg13g2_decap_8 FILLER_69_2412 ();
 sg13g2_decap_8 FILLER_69_2419 ();
 sg13g2_decap_8 FILLER_69_2430 ();
 sg13g2_decap_8 FILLER_69_2437 ();
 sg13g2_decap_4 FILLER_69_2444 ();
 sg13g2_fill_2 FILLER_69_2448 ();
 sg13g2_decap_8 FILLER_69_2472 ();
 sg13g2_decap_8 FILLER_69_2479 ();
 sg13g2_fill_1 FILLER_69_2486 ();
 sg13g2_fill_2 FILLER_69_2492 ();
 sg13g2_fill_2 FILLER_69_2499 ();
 sg13g2_decap_8 FILLER_69_2506 ();
 sg13g2_decap_8 FILLER_69_2513 ();
 sg13g2_decap_8 FILLER_69_2520 ();
 sg13g2_decap_8 FILLER_69_2527 ();
 sg13g2_decap_8 FILLER_69_2534 ();
 sg13g2_decap_8 FILLER_69_2541 ();
 sg13g2_decap_8 FILLER_69_2574 ();
 sg13g2_decap_8 FILLER_69_2581 ();
 sg13g2_decap_8 FILLER_69_2588 ();
 sg13g2_decap_8 FILLER_69_2595 ();
 sg13g2_decap_8 FILLER_69_2602 ();
 sg13g2_decap_8 FILLER_69_2609 ();
 sg13g2_decap_8 FILLER_69_2616 ();
 sg13g2_decap_8 FILLER_69_2623 ();
 sg13g2_decap_8 FILLER_69_2630 ();
 sg13g2_decap_8 FILLER_69_2637 ();
 sg13g2_fill_2 FILLER_69_2644 ();
 sg13g2_decap_8 FILLER_69_2676 ();
 sg13g2_decap_8 FILLER_69_2683 ();
 sg13g2_decap_4 FILLER_69_2690 ();
 sg13g2_fill_2 FILLER_69_2694 ();
 sg13g2_decap_8 FILLER_69_2711 ();
 sg13g2_fill_1 FILLER_69_2718 ();
 sg13g2_decap_8 FILLER_69_2738 ();
 sg13g2_decap_8 FILLER_69_2745 ();
 sg13g2_decap_8 FILLER_69_2752 ();
 sg13g2_fill_2 FILLER_69_2759 ();
 sg13g2_fill_1 FILLER_69_2761 ();
 sg13g2_decap_8 FILLER_69_2783 ();
 sg13g2_decap_8 FILLER_69_2790 ();
 sg13g2_decap_8 FILLER_69_2797 ();
 sg13g2_decap_8 FILLER_69_2804 ();
 sg13g2_decap_8 FILLER_69_2811 ();
 sg13g2_decap_8 FILLER_69_2818 ();
 sg13g2_decap_8 FILLER_69_2825 ();
 sg13g2_decap_8 FILLER_69_2832 ();
 sg13g2_decap_8 FILLER_69_2839 ();
 sg13g2_decap_8 FILLER_69_2846 ();
 sg13g2_decap_8 FILLER_69_2853 ();
 sg13g2_fill_1 FILLER_69_2860 ();
 sg13g2_decap_8 FILLER_69_2869 ();
 sg13g2_decap_8 FILLER_69_2876 ();
 sg13g2_decap_8 FILLER_69_2883 ();
 sg13g2_decap_8 FILLER_69_2890 ();
 sg13g2_decap_8 FILLER_69_2897 ();
 sg13g2_decap_8 FILLER_69_2904 ();
 sg13g2_decap_8 FILLER_69_2911 ();
 sg13g2_decap_8 FILLER_69_2918 ();
 sg13g2_decap_8 FILLER_69_2925 ();
 sg13g2_decap_8 FILLER_69_2932 ();
 sg13g2_fill_1 FILLER_69_2939 ();
 sg13g2_decap_8 FILLER_69_2981 ();
 sg13g2_decap_8 FILLER_69_2988 ();
 sg13g2_fill_2 FILLER_69_2995 ();
 sg13g2_fill_1 FILLER_69_3017 ();
 sg13g2_decap_4 FILLER_69_3039 ();
 sg13g2_decap_4 FILLER_69_3058 ();
 sg13g2_fill_1 FILLER_69_3062 ();
 sg13g2_fill_2 FILLER_69_3068 ();
 sg13g2_decap_8 FILLER_69_3096 ();
 sg13g2_decap_8 FILLER_69_3108 ();
 sg13g2_decap_8 FILLER_69_3115 ();
 sg13g2_decap_8 FILLER_69_3122 ();
 sg13g2_decap_8 FILLER_69_3129 ();
 sg13g2_decap_8 FILLER_69_3164 ();
 sg13g2_decap_8 FILLER_69_3171 ();
 sg13g2_decap_4 FILLER_69_3178 ();
 sg13g2_decap_8 FILLER_69_3208 ();
 sg13g2_fill_1 FILLER_69_3215 ();
 sg13g2_decap_8 FILLER_69_3224 ();
 sg13g2_decap_8 FILLER_69_3231 ();
 sg13g2_decap_8 FILLER_69_3238 ();
 sg13g2_decap_8 FILLER_69_3245 ();
 sg13g2_decap_8 FILLER_69_3252 ();
 sg13g2_decap_8 FILLER_69_3259 ();
 sg13g2_decap_8 FILLER_69_3266 ();
 sg13g2_decap_8 FILLER_69_3273 ();
 sg13g2_decap_8 FILLER_69_3280 ();
 sg13g2_decap_8 FILLER_69_3287 ();
 sg13g2_decap_8 FILLER_69_3294 ();
 sg13g2_fill_1 FILLER_69_3301 ();
 sg13g2_decap_8 FILLER_69_3317 ();
 sg13g2_fill_2 FILLER_69_3324 ();
 sg13g2_fill_1 FILLER_69_3326 ();
 sg13g2_decap_8 FILLER_69_3342 ();
 sg13g2_decap_8 FILLER_69_3349 ();
 sg13g2_decap_8 FILLER_69_3356 ();
 sg13g2_fill_2 FILLER_69_3368 ();
 sg13g2_fill_1 FILLER_69_3370 ();
 sg13g2_fill_2 FILLER_69_3381 ();
 sg13g2_decap_8 FILLER_69_3388 ();
 sg13g2_decap_4 FILLER_69_3395 ();
 sg13g2_fill_1 FILLER_69_3399 ();
 sg13g2_decap_8 FILLER_69_3419 ();
 sg13g2_decap_8 FILLER_69_3426 ();
 sg13g2_decap_4 FILLER_69_3433 ();
 sg13g2_fill_2 FILLER_69_3437 ();
 sg13g2_decap_8 FILLER_69_3442 ();
 sg13g2_decap_8 FILLER_69_3449 ();
 sg13g2_decap_8 FILLER_69_3456 ();
 sg13g2_decap_4 FILLER_69_3468 ();
 sg13g2_decap_8 FILLER_69_3498 ();
 sg13g2_decap_8 FILLER_69_3505 ();
 sg13g2_decap_8 FILLER_69_3512 ();
 sg13g2_decap_8 FILLER_69_3519 ();
 sg13g2_decap_8 FILLER_69_3526 ();
 sg13g2_decap_8 FILLER_69_3533 ();
 sg13g2_decap_8 FILLER_69_3540 ();
 sg13g2_decap_8 FILLER_69_3547 ();
 sg13g2_decap_8 FILLER_69_3554 ();
 sg13g2_decap_8 FILLER_69_3561 ();
 sg13g2_decap_8 FILLER_69_3568 ();
 sg13g2_decap_4 FILLER_69_3575 ();
 sg13g2_fill_1 FILLER_69_3579 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_fill_2 FILLER_70_14 ();
 sg13g2_fill_1 FILLER_70_16 ();
 sg13g2_fill_2 FILLER_70_26 ();
 sg13g2_decap_8 FILLER_70_37 ();
 sg13g2_decap_8 FILLER_70_44 ();
 sg13g2_decap_8 FILLER_70_51 ();
 sg13g2_decap_8 FILLER_70_58 ();
 sg13g2_decap_8 FILLER_70_65 ();
 sg13g2_decap_4 FILLER_70_77 ();
 sg13g2_decap_8 FILLER_70_86 ();
 sg13g2_decap_8 FILLER_70_93 ();
 sg13g2_decap_8 FILLER_70_100 ();
 sg13g2_decap_4 FILLER_70_107 ();
 sg13g2_fill_2 FILLER_70_111 ();
 sg13g2_decap_8 FILLER_70_131 ();
 sg13g2_decap_8 FILLER_70_138 ();
 sg13g2_decap_4 FILLER_70_145 ();
 sg13g2_fill_2 FILLER_70_149 ();
 sg13g2_fill_2 FILLER_70_165 ();
 sg13g2_decap_8 FILLER_70_172 ();
 sg13g2_decap_8 FILLER_70_179 ();
 sg13g2_decap_8 FILLER_70_186 ();
 sg13g2_decap_8 FILLER_70_193 ();
 sg13g2_decap_8 FILLER_70_200 ();
 sg13g2_decap_8 FILLER_70_207 ();
 sg13g2_decap_8 FILLER_70_214 ();
 sg13g2_decap_8 FILLER_70_221 ();
 sg13g2_fill_1 FILLER_70_228 ();
 sg13g2_fill_2 FILLER_70_233 ();
 sg13g2_fill_1 FILLER_70_235 ();
 sg13g2_decap_8 FILLER_70_240 ();
 sg13g2_decap_8 FILLER_70_247 ();
 sg13g2_decap_8 FILLER_70_254 ();
 sg13g2_decap_8 FILLER_70_261 ();
 sg13g2_decap_8 FILLER_70_268 ();
 sg13g2_decap_4 FILLER_70_275 ();
 sg13g2_fill_1 FILLER_70_279 ();
 sg13g2_decap_4 FILLER_70_283 ();
 sg13g2_fill_1 FILLER_70_287 ();
 sg13g2_fill_2 FILLER_70_291 ();
 sg13g2_fill_1 FILLER_70_293 ();
 sg13g2_decap_8 FILLER_70_297 ();
 sg13g2_decap_8 FILLER_70_304 ();
 sg13g2_decap_8 FILLER_70_311 ();
 sg13g2_decap_8 FILLER_70_318 ();
 sg13g2_decap_8 FILLER_70_325 ();
 sg13g2_decap_8 FILLER_70_332 ();
 sg13g2_decap_8 FILLER_70_339 ();
 sg13g2_fill_1 FILLER_70_346 ();
 sg13g2_decap_4 FILLER_70_352 ();
 sg13g2_decap_8 FILLER_70_370 ();
 sg13g2_decap_8 FILLER_70_377 ();
 sg13g2_decap_4 FILLER_70_384 ();
 sg13g2_decap_8 FILLER_70_404 ();
 sg13g2_decap_8 FILLER_70_411 ();
 sg13g2_decap_8 FILLER_70_418 ();
 sg13g2_fill_1 FILLER_70_425 ();
 sg13g2_decap_8 FILLER_70_432 ();
 sg13g2_fill_2 FILLER_70_439 ();
 sg13g2_fill_1 FILLER_70_441 ();
 sg13g2_decap_8 FILLER_70_445 ();
 sg13g2_decap_8 FILLER_70_452 ();
 sg13g2_decap_4 FILLER_70_459 ();
 sg13g2_fill_2 FILLER_70_469 ();
 sg13g2_decap_8 FILLER_70_501 ();
 sg13g2_decap_8 FILLER_70_508 ();
 sg13g2_decap_8 FILLER_70_515 ();
 sg13g2_decap_8 FILLER_70_522 ();
 sg13g2_decap_8 FILLER_70_529 ();
 sg13g2_decap_4 FILLER_70_536 ();
 sg13g2_fill_1 FILLER_70_540 ();
 sg13g2_decap_8 FILLER_70_554 ();
 sg13g2_decap_8 FILLER_70_561 ();
 sg13g2_decap_8 FILLER_70_568 ();
 sg13g2_decap_8 FILLER_70_575 ();
 sg13g2_decap_8 FILLER_70_582 ();
 sg13g2_decap_8 FILLER_70_589 ();
 sg13g2_fill_1 FILLER_70_596 ();
 sg13g2_decap_8 FILLER_70_612 ();
 sg13g2_decap_8 FILLER_70_619 ();
 sg13g2_decap_8 FILLER_70_660 ();
 sg13g2_decap_8 FILLER_70_667 ();
 sg13g2_decap_8 FILLER_70_674 ();
 sg13g2_decap_8 FILLER_70_681 ();
 sg13g2_decap_8 FILLER_70_688 ();
 sg13g2_decap_4 FILLER_70_695 ();
 sg13g2_fill_1 FILLER_70_699 ();
 sg13g2_decap_4 FILLER_70_712 ();
 sg13g2_fill_2 FILLER_70_716 ();
 sg13g2_fill_2 FILLER_70_739 ();
 sg13g2_decap_8 FILLER_70_746 ();
 sg13g2_decap_8 FILLER_70_753 ();
 sg13g2_decap_8 FILLER_70_760 ();
 sg13g2_decap_4 FILLER_70_767 ();
 sg13g2_fill_2 FILLER_70_776 ();
 sg13g2_decap_4 FILLER_70_788 ();
 sg13g2_fill_2 FILLER_70_792 ();
 sg13g2_fill_1 FILLER_70_799 ();
 sg13g2_decap_8 FILLER_70_808 ();
 sg13g2_decap_8 FILLER_70_815 ();
 sg13g2_fill_1 FILLER_70_822 ();
 sg13g2_fill_1 FILLER_70_826 ();
 sg13g2_decap_8 FILLER_70_835 ();
 sg13g2_decap_8 FILLER_70_842 ();
 sg13g2_decap_8 FILLER_70_849 ();
 sg13g2_decap_4 FILLER_70_856 ();
 sg13g2_fill_2 FILLER_70_860 ();
 sg13g2_decap_8 FILLER_70_872 ();
 sg13g2_decap_8 FILLER_70_879 ();
 sg13g2_decap_8 FILLER_70_886 ();
 sg13g2_decap_8 FILLER_70_893 ();
 sg13g2_decap_8 FILLER_70_900 ();
 sg13g2_decap_8 FILLER_70_907 ();
 sg13g2_decap_8 FILLER_70_914 ();
 sg13g2_decap_8 FILLER_70_921 ();
 sg13g2_decap_4 FILLER_70_928 ();
 sg13g2_fill_1 FILLER_70_932 ();
 sg13g2_fill_2 FILLER_70_944 ();
 sg13g2_fill_1 FILLER_70_946 ();
 sg13g2_decap_8 FILLER_70_950 ();
 sg13g2_decap_4 FILLER_70_957 ();
 sg13g2_fill_1 FILLER_70_961 ();
 sg13g2_fill_1 FILLER_70_966 ();
 sg13g2_fill_2 FILLER_70_983 ();
 sg13g2_fill_1 FILLER_70_985 ();
 sg13g2_decap_8 FILLER_70_994 ();
 sg13g2_decap_4 FILLER_70_1001 ();
 sg13g2_fill_1 FILLER_70_1005 ();
 sg13g2_decap_8 FILLER_70_1012 ();
 sg13g2_decap_8 FILLER_70_1019 ();
 sg13g2_decap_4 FILLER_70_1026 ();
 sg13g2_fill_2 FILLER_70_1030 ();
 sg13g2_decap_8 FILLER_70_1061 ();
 sg13g2_decap_8 FILLER_70_1068 ();
 sg13g2_decap_8 FILLER_70_1075 ();
 sg13g2_decap_8 FILLER_70_1082 ();
 sg13g2_decap_8 FILLER_70_1089 ();
 sg13g2_decap_8 FILLER_70_1096 ();
 sg13g2_decap_4 FILLER_70_1103 ();
 sg13g2_fill_1 FILLER_70_1107 ();
 sg13g2_decap_8 FILLER_70_1139 ();
 sg13g2_decap_8 FILLER_70_1146 ();
 sg13g2_fill_1 FILLER_70_1153 ();
 sg13g2_decap_8 FILLER_70_1162 ();
 sg13g2_decap_8 FILLER_70_1169 ();
 sg13g2_decap_8 FILLER_70_1176 ();
 sg13g2_decap_8 FILLER_70_1183 ();
 sg13g2_decap_4 FILLER_70_1190 ();
 sg13g2_fill_2 FILLER_70_1194 ();
 sg13g2_decap_4 FILLER_70_1204 ();
 sg13g2_decap_8 FILLER_70_1220 ();
 sg13g2_decap_8 FILLER_70_1227 ();
 sg13g2_fill_2 FILLER_70_1234 ();
 sg13g2_fill_1 FILLER_70_1236 ();
 sg13g2_decap_8 FILLER_70_1240 ();
 sg13g2_decap_8 FILLER_70_1247 ();
 sg13g2_decap_8 FILLER_70_1254 ();
 sg13g2_decap_8 FILLER_70_1261 ();
 sg13g2_decap_8 FILLER_70_1268 ();
 sg13g2_decap_8 FILLER_70_1275 ();
 sg13g2_decap_8 FILLER_70_1282 ();
 sg13g2_decap_4 FILLER_70_1289 ();
 sg13g2_fill_1 FILLER_70_1293 ();
 sg13g2_fill_1 FILLER_70_1339 ();
 sg13g2_decap_8 FILLER_70_1363 ();
 sg13g2_decap_8 FILLER_70_1370 ();
 sg13g2_decap_8 FILLER_70_1377 ();
 sg13g2_decap_8 FILLER_70_1384 ();
 sg13g2_decap_8 FILLER_70_1391 ();
 sg13g2_decap_8 FILLER_70_1398 ();
 sg13g2_decap_8 FILLER_70_1405 ();
 sg13g2_decap_8 FILLER_70_1412 ();
 sg13g2_decap_8 FILLER_70_1419 ();
 sg13g2_decap_8 FILLER_70_1426 ();
 sg13g2_decap_8 FILLER_70_1433 ();
 sg13g2_fill_2 FILLER_70_1440 ();
 sg13g2_fill_1 FILLER_70_1442 ();
 sg13g2_decap_8 FILLER_70_1479 ();
 sg13g2_fill_2 FILLER_70_1486 ();
 sg13g2_fill_1 FILLER_70_1514 ();
 sg13g2_decap_4 FILLER_70_1525 ();
 sg13g2_fill_2 FILLER_70_1529 ();
 sg13g2_decap_4 FILLER_70_1567 ();
 sg13g2_fill_1 FILLER_70_1571 ();
 sg13g2_decap_8 FILLER_70_1598 ();
 sg13g2_decap_8 FILLER_70_1605 ();
 sg13g2_decap_4 FILLER_70_1612 ();
 sg13g2_fill_2 FILLER_70_1616 ();
 sg13g2_decap_8 FILLER_70_1621 ();
 sg13g2_fill_2 FILLER_70_1628 ();
 sg13g2_decap_8 FILLER_70_1638 ();
 sg13g2_decap_8 FILLER_70_1645 ();
 sg13g2_decap_8 FILLER_70_1652 ();
 sg13g2_decap_8 FILLER_70_1659 ();
 sg13g2_fill_1 FILLER_70_1666 ();
 sg13g2_decap_8 FILLER_70_1671 ();
 sg13g2_decap_8 FILLER_70_1678 ();
 sg13g2_decap_8 FILLER_70_1685 ();
 sg13g2_decap_8 FILLER_70_1692 ();
 sg13g2_decap_8 FILLER_70_1699 ();
 sg13g2_decap_8 FILLER_70_1706 ();
 sg13g2_decap_8 FILLER_70_1713 ();
 sg13g2_fill_1 FILLER_70_1720 ();
 sg13g2_fill_2 FILLER_70_1724 ();
 sg13g2_fill_1 FILLER_70_1726 ();
 sg13g2_decap_8 FILLER_70_1736 ();
 sg13g2_decap_8 FILLER_70_1743 ();
 sg13g2_decap_8 FILLER_70_1750 ();
 sg13g2_fill_1 FILLER_70_1757 ();
 sg13g2_fill_2 FILLER_70_1768 ();
 sg13g2_decap_4 FILLER_70_1796 ();
 sg13g2_decap_8 FILLER_70_1826 ();
 sg13g2_decap_8 FILLER_70_1833 ();
 sg13g2_decap_8 FILLER_70_1840 ();
 sg13g2_decap_8 FILLER_70_1847 ();
 sg13g2_decap_8 FILLER_70_1854 ();
 sg13g2_decap_8 FILLER_70_1861 ();
 sg13g2_decap_8 FILLER_70_1894 ();
 sg13g2_decap_8 FILLER_70_1901 ();
 sg13g2_decap_8 FILLER_70_1908 ();
 sg13g2_decap_8 FILLER_70_1915 ();
 sg13g2_decap_8 FILLER_70_1922 ();
 sg13g2_decap_8 FILLER_70_1929 ();
 sg13g2_decap_8 FILLER_70_1936 ();
 sg13g2_decap_8 FILLER_70_1943 ();
 sg13g2_decap_8 FILLER_70_1950 ();
 sg13g2_decap_8 FILLER_70_1957 ();
 sg13g2_decap_8 FILLER_70_1964 ();
 sg13g2_decap_8 FILLER_70_1971 ();
 sg13g2_fill_1 FILLER_70_1978 ();
 sg13g2_decap_8 FILLER_70_1989 ();
 sg13g2_decap_8 FILLER_70_1996 ();
 sg13g2_decap_8 FILLER_70_2003 ();
 sg13g2_decap_8 FILLER_70_2010 ();
 sg13g2_decap_8 FILLER_70_2017 ();
 sg13g2_decap_8 FILLER_70_2024 ();
 sg13g2_decap_8 FILLER_70_2031 ();
 sg13g2_decap_8 FILLER_70_2038 ();
 sg13g2_decap_8 FILLER_70_2045 ();
 sg13g2_decap_8 FILLER_70_2052 ();
 sg13g2_decap_8 FILLER_70_2059 ();
 sg13g2_decap_8 FILLER_70_2066 ();
 sg13g2_fill_2 FILLER_70_2073 ();
 sg13g2_fill_1 FILLER_70_2075 ();
 sg13g2_decap_8 FILLER_70_2086 ();
 sg13g2_decap_8 FILLER_70_2093 ();
 sg13g2_decap_8 FILLER_70_2100 ();
 sg13g2_decap_8 FILLER_70_2107 ();
 sg13g2_decap_8 FILLER_70_2114 ();
 sg13g2_decap_8 FILLER_70_2121 ();
 sg13g2_fill_2 FILLER_70_2128 ();
 sg13g2_decap_8 FILLER_70_2140 ();
 sg13g2_decap_4 FILLER_70_2147 ();
 sg13g2_fill_1 FILLER_70_2151 ();
 sg13g2_decap_8 FILLER_70_2188 ();
 sg13g2_decap_8 FILLER_70_2195 ();
 sg13g2_decap_8 FILLER_70_2202 ();
 sg13g2_decap_8 FILLER_70_2209 ();
 sg13g2_decap_8 FILLER_70_2216 ();
 sg13g2_decap_8 FILLER_70_2223 ();
 sg13g2_decap_8 FILLER_70_2230 ();
 sg13g2_decap_8 FILLER_70_2237 ();
 sg13g2_decap_8 FILLER_70_2244 ();
 sg13g2_decap_8 FILLER_70_2251 ();
 sg13g2_decap_8 FILLER_70_2258 ();
 sg13g2_decap_8 FILLER_70_2265 ();
 sg13g2_decap_8 FILLER_70_2272 ();
 sg13g2_decap_8 FILLER_70_2279 ();
 sg13g2_decap_8 FILLER_70_2286 ();
 sg13g2_decap_8 FILLER_70_2293 ();
 sg13g2_decap_8 FILLER_70_2300 ();
 sg13g2_decap_8 FILLER_70_2307 ();
 sg13g2_decap_8 FILLER_70_2314 ();
 sg13g2_decap_8 FILLER_70_2321 ();
 sg13g2_decap_8 FILLER_70_2328 ();
 sg13g2_fill_1 FILLER_70_2335 ();
 sg13g2_decap_4 FILLER_70_2362 ();
 sg13g2_fill_2 FILLER_70_2366 ();
 sg13g2_decap_8 FILLER_70_2373 ();
 sg13g2_decap_8 FILLER_70_2380 ();
 sg13g2_decap_4 FILLER_70_2387 ();
 sg13g2_fill_1 FILLER_70_2391 ();
 sg13g2_decap_8 FILLER_70_2423 ();
 sg13g2_decap_8 FILLER_70_2430 ();
 sg13g2_decap_8 FILLER_70_2437 ();
 sg13g2_decap_8 FILLER_70_2444 ();
 sg13g2_fill_2 FILLER_70_2472 ();
 sg13g2_fill_2 FILLER_70_2479 ();
 sg13g2_fill_2 FILLER_70_2491 ();
 sg13g2_fill_2 FILLER_70_2514 ();
 sg13g2_fill_1 FILLER_70_2516 ();
 sg13g2_fill_1 FILLER_70_2537 ();
 sg13g2_fill_2 FILLER_70_2542 ();
 sg13g2_decap_8 FILLER_70_2570 ();
 sg13g2_decap_8 FILLER_70_2577 ();
 sg13g2_decap_8 FILLER_70_2584 ();
 sg13g2_decap_8 FILLER_70_2591 ();
 sg13g2_decap_8 FILLER_70_2598 ();
 sg13g2_fill_2 FILLER_70_2605 ();
 sg13g2_fill_1 FILLER_70_2607 ();
 sg13g2_decap_8 FILLER_70_2619 ();
 sg13g2_decap_8 FILLER_70_2626 ();
 sg13g2_decap_8 FILLER_70_2633 ();
 sg13g2_decap_8 FILLER_70_2640 ();
 sg13g2_decap_8 FILLER_70_2647 ();
 sg13g2_fill_2 FILLER_70_2654 ();
 sg13g2_decap_8 FILLER_70_2666 ();
 sg13g2_decap_8 FILLER_70_2673 ();
 sg13g2_decap_8 FILLER_70_2680 ();
 sg13g2_decap_8 FILLER_70_2687 ();
 sg13g2_decap_8 FILLER_70_2699 ();
 sg13g2_decap_8 FILLER_70_2706 ();
 sg13g2_decap_8 FILLER_70_2713 ();
 sg13g2_decap_8 FILLER_70_2720 ();
 sg13g2_fill_1 FILLER_70_2727 ();
 sg13g2_decap_8 FILLER_70_2733 ();
 sg13g2_decap_8 FILLER_70_2740 ();
 sg13g2_decap_8 FILLER_70_2747 ();
 sg13g2_decap_8 FILLER_70_2754 ();
 sg13g2_decap_8 FILLER_70_2761 ();
 sg13g2_decap_8 FILLER_70_2768 ();
 sg13g2_decap_8 FILLER_70_2775 ();
 sg13g2_fill_2 FILLER_70_2782 ();
 sg13g2_decap_8 FILLER_70_2789 ();
 sg13g2_decap_8 FILLER_70_2796 ();
 sg13g2_fill_1 FILLER_70_2803 ();
 sg13g2_decap_4 FILLER_70_2824 ();
 sg13g2_fill_1 FILLER_70_2828 ();
 sg13g2_fill_1 FILLER_70_2855 ();
 sg13g2_decap_4 FILLER_70_2892 ();
 sg13g2_fill_2 FILLER_70_2896 ();
 sg13g2_decap_8 FILLER_70_2924 ();
 sg13g2_fill_2 FILLER_70_2931 ();
 sg13g2_fill_1 FILLER_70_2933 ();
 sg13g2_decap_8 FILLER_70_2939 ();
 sg13g2_decap_4 FILLER_70_2946 ();
 sg13g2_fill_2 FILLER_70_2950 ();
 sg13g2_decap_8 FILLER_70_2976 ();
 sg13g2_decap_8 FILLER_70_2983 ();
 sg13g2_decap_8 FILLER_70_2990 ();
 sg13g2_decap_8 FILLER_70_2997 ();
 sg13g2_decap_8 FILLER_70_3024 ();
 sg13g2_decap_8 FILLER_70_3031 ();
 sg13g2_decap_8 FILLER_70_3048 ();
 sg13g2_decap_8 FILLER_70_3055 ();
 sg13g2_decap_4 FILLER_70_3062 ();
 sg13g2_fill_2 FILLER_70_3066 ();
 sg13g2_decap_4 FILLER_70_3078 ();
 sg13g2_fill_1 FILLER_70_3082 ();
 sg13g2_decap_8 FILLER_70_3088 ();
 sg13g2_decap_8 FILLER_70_3100 ();
 sg13g2_decap_8 FILLER_70_3107 ();
 sg13g2_fill_1 FILLER_70_3114 ();
 sg13g2_decap_8 FILLER_70_3119 ();
 sg13g2_decap_8 FILLER_70_3126 ();
 sg13g2_decap_8 FILLER_70_3133 ();
 sg13g2_fill_2 FILLER_70_3140 ();
 sg13g2_fill_1 FILLER_70_3142 ();
 sg13g2_decap_8 FILLER_70_3147 ();
 sg13g2_fill_2 FILLER_70_3154 ();
 sg13g2_decap_8 FILLER_70_3164 ();
 sg13g2_decap_8 FILLER_70_3171 ();
 sg13g2_decap_8 FILLER_70_3178 ();
 sg13g2_decap_8 FILLER_70_3185 ();
 sg13g2_decap_8 FILLER_70_3200 ();
 sg13g2_decap_8 FILLER_70_3207 ();
 sg13g2_decap_8 FILLER_70_3214 ();
 sg13g2_decap_8 FILLER_70_3221 ();
 sg13g2_decap_8 FILLER_70_3236 ();
 sg13g2_decap_8 FILLER_70_3243 ();
 sg13g2_decap_8 FILLER_70_3250 ();
 sg13g2_decap_8 FILLER_70_3257 ();
 sg13g2_decap_4 FILLER_70_3264 ();
 sg13g2_decap_8 FILLER_70_3293 ();
 sg13g2_decap_8 FILLER_70_3300 ();
 sg13g2_decap_8 FILLER_70_3307 ();
 sg13g2_decap_8 FILLER_70_3314 ();
 sg13g2_decap_8 FILLER_70_3321 ();
 sg13g2_decap_8 FILLER_70_3328 ();
 sg13g2_decap_8 FILLER_70_3335 ();
 sg13g2_decap_8 FILLER_70_3342 ();
 sg13g2_fill_2 FILLER_70_3349 ();
 sg13g2_fill_1 FILLER_70_3351 ();
 sg13g2_decap_8 FILLER_70_3357 ();
 sg13g2_decap_8 FILLER_70_3364 ();
 sg13g2_decap_8 FILLER_70_3371 ();
 sg13g2_decap_8 FILLER_70_3378 ();
 sg13g2_decap_8 FILLER_70_3385 ();
 sg13g2_decap_4 FILLER_70_3392 ();
 sg13g2_fill_1 FILLER_70_3396 ();
 sg13g2_fill_2 FILLER_70_3407 ();
 sg13g2_fill_1 FILLER_70_3409 ();
 sg13g2_fill_2 FILLER_70_3419 ();
 sg13g2_decap_8 FILLER_70_3426 ();
 sg13g2_decap_8 FILLER_70_3433 ();
 sg13g2_decap_8 FILLER_70_3440 ();
 sg13g2_fill_1 FILLER_70_3452 ();
 sg13g2_decap_8 FILLER_70_3462 ();
 sg13g2_decap_8 FILLER_70_3469 ();
 sg13g2_decap_8 FILLER_70_3476 ();
 sg13g2_decap_8 FILLER_70_3483 ();
 sg13g2_decap_8 FILLER_70_3490 ();
 sg13g2_decap_8 FILLER_70_3507 ();
 sg13g2_decap_8 FILLER_70_3514 ();
 sg13g2_decap_8 FILLER_70_3521 ();
 sg13g2_decap_8 FILLER_70_3528 ();
 sg13g2_decap_8 FILLER_70_3535 ();
 sg13g2_decap_8 FILLER_70_3542 ();
 sg13g2_decap_8 FILLER_70_3549 ();
 sg13g2_decap_8 FILLER_70_3556 ();
 sg13g2_decap_8 FILLER_70_3563 ();
 sg13g2_decap_8 FILLER_70_3570 ();
 sg13g2_fill_2 FILLER_70_3577 ();
 sg13g2_fill_1 FILLER_70_3579 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_fill_2 FILLER_71_7 ();
 sg13g2_fill_1 FILLER_71_9 ();
 sg13g2_decap_8 FILLER_71_50 ();
 sg13g2_decap_8 FILLER_71_57 ();
 sg13g2_decap_8 FILLER_71_64 ();
 sg13g2_fill_1 FILLER_71_71 ();
 sg13g2_decap_8 FILLER_71_77 ();
 sg13g2_decap_8 FILLER_71_84 ();
 sg13g2_decap_8 FILLER_71_91 ();
 sg13g2_decap_4 FILLER_71_98 ();
 sg13g2_fill_1 FILLER_71_102 ();
 sg13g2_decap_8 FILLER_71_143 ();
 sg13g2_decap_8 FILLER_71_150 ();
 sg13g2_fill_2 FILLER_71_157 ();
 sg13g2_fill_1 FILLER_71_159 ();
 sg13g2_decap_4 FILLER_71_165 ();
 sg13g2_fill_2 FILLER_71_182 ();
 sg13g2_decap_8 FILLER_71_193 ();
 sg13g2_decap_8 FILLER_71_200 ();
 sg13g2_decap_8 FILLER_71_207 ();
 sg13g2_decap_8 FILLER_71_214 ();
 sg13g2_decap_8 FILLER_71_226 ();
 sg13g2_decap_8 FILLER_71_233 ();
 sg13g2_decap_8 FILLER_71_240 ();
 sg13g2_decap_8 FILLER_71_247 ();
 sg13g2_decap_8 FILLER_71_254 ();
 sg13g2_decap_8 FILLER_71_261 ();
 sg13g2_decap_8 FILLER_71_268 ();
 sg13g2_fill_2 FILLER_71_275 ();
 sg13g2_fill_2 FILLER_71_291 ();
 sg13g2_fill_1 FILLER_71_293 ();
 sg13g2_decap_8 FILLER_71_323 ();
 sg13g2_decap_8 FILLER_71_330 ();
 sg13g2_decap_8 FILLER_71_337 ();
 sg13g2_decap_4 FILLER_71_344 ();
 sg13g2_fill_1 FILLER_71_348 ();
 sg13g2_decap_4 FILLER_71_384 ();
 sg13g2_fill_2 FILLER_71_388 ();
 sg13g2_decap_8 FILLER_71_397 ();
 sg13g2_decap_8 FILLER_71_404 ();
 sg13g2_decap_8 FILLER_71_411 ();
 sg13g2_fill_1 FILLER_71_418 ();
 sg13g2_fill_1 FILLER_71_461 ();
 sg13g2_decap_4 FILLER_71_468 ();
 sg13g2_fill_2 FILLER_71_472 ();
 sg13g2_decap_8 FILLER_71_504 ();
 sg13g2_decap_8 FILLER_71_511 ();
 sg13g2_decap_8 FILLER_71_518 ();
 sg13g2_decap_8 FILLER_71_525 ();
 sg13g2_decap_8 FILLER_71_532 ();
 sg13g2_decap_8 FILLER_71_539 ();
 sg13g2_decap_8 FILLER_71_546 ();
 sg13g2_decap_8 FILLER_71_553 ();
 sg13g2_decap_8 FILLER_71_560 ();
 sg13g2_decap_8 FILLER_71_567 ();
 sg13g2_decap_8 FILLER_71_574 ();
 sg13g2_decap_4 FILLER_71_581 ();
 sg13g2_fill_2 FILLER_71_595 ();
 sg13g2_decap_8 FILLER_71_605 ();
 sg13g2_decap_8 FILLER_71_612 ();
 sg13g2_decap_8 FILLER_71_619 ();
 sg13g2_decap_8 FILLER_71_626 ();
 sg13g2_decap_8 FILLER_71_673 ();
 sg13g2_decap_8 FILLER_71_680 ();
 sg13g2_decap_8 FILLER_71_687 ();
 sg13g2_fill_1 FILLER_71_694 ();
 sg13g2_decap_8 FILLER_71_701 ();
 sg13g2_decap_4 FILLER_71_708 ();
 sg13g2_fill_2 FILLER_71_712 ();
 sg13g2_fill_2 FILLER_71_717 ();
 sg13g2_decap_8 FILLER_71_757 ();
 sg13g2_decap_8 FILLER_71_764 ();
 sg13g2_fill_2 FILLER_71_771 ();
 sg13g2_fill_1 FILLER_71_773 ();
 sg13g2_decap_8 FILLER_71_782 ();
 sg13g2_decap_8 FILLER_71_789 ();
 sg13g2_decap_8 FILLER_71_796 ();
 sg13g2_decap_8 FILLER_71_803 ();
 sg13g2_decap_8 FILLER_71_810 ();
 sg13g2_decap_8 FILLER_71_817 ();
 sg13g2_decap_8 FILLER_71_824 ();
 sg13g2_fill_2 FILLER_71_831 ();
 sg13g2_fill_1 FILLER_71_833 ();
 sg13g2_fill_2 FILLER_71_838 ();
 sg13g2_fill_1 FILLER_71_840 ();
 sg13g2_decap_8 FILLER_71_851 ();
 sg13g2_decap_8 FILLER_71_858 ();
 sg13g2_decap_8 FILLER_71_865 ();
 sg13g2_decap_4 FILLER_71_872 ();
 sg13g2_fill_2 FILLER_71_876 ();
 sg13g2_decap_4 FILLER_71_890 ();
 sg13g2_fill_2 FILLER_71_894 ();
 sg13g2_fill_2 FILLER_71_900 ();
 sg13g2_fill_1 FILLER_71_902 ();
 sg13g2_decap_8 FILLER_71_911 ();
 sg13g2_decap_8 FILLER_71_918 ();
 sg13g2_decap_8 FILLER_71_925 ();
 sg13g2_fill_2 FILLER_71_932 ();
 sg13g2_decap_8 FILLER_71_939 ();
 sg13g2_fill_1 FILLER_71_946 ();
 sg13g2_fill_2 FILLER_71_952 ();
 sg13g2_decap_8 FILLER_71_959 ();
 sg13g2_decap_4 FILLER_71_966 ();
 sg13g2_fill_2 FILLER_71_970 ();
 sg13g2_decap_8 FILLER_71_983 ();
 sg13g2_decap_4 FILLER_71_990 ();
 sg13g2_fill_2 FILLER_71_994 ();
 sg13g2_decap_8 FILLER_71_1002 ();
 sg13g2_fill_2 FILLER_71_1009 ();
 sg13g2_fill_1 FILLER_71_1011 ();
 sg13g2_decap_8 FILLER_71_1017 ();
 sg13g2_decap_8 FILLER_71_1024 ();
 sg13g2_decap_8 FILLER_71_1031 ();
 sg13g2_fill_1 FILLER_71_1038 ();
 sg13g2_fill_1 FILLER_71_1043 ();
 sg13g2_decap_8 FILLER_71_1049 ();
 sg13g2_fill_1 FILLER_71_1056 ();
 sg13g2_decap_8 FILLER_71_1065 ();
 sg13g2_decap_8 FILLER_71_1072 ();
 sg13g2_decap_8 FILLER_71_1079 ();
 sg13g2_decap_8 FILLER_71_1086 ();
 sg13g2_decap_8 FILLER_71_1093 ();
 sg13g2_decap_8 FILLER_71_1100 ();
 sg13g2_decap_4 FILLER_71_1107 ();
 sg13g2_decap_8 FILLER_71_1119 ();
 sg13g2_decap_4 FILLER_71_1126 ();
 sg13g2_decap_8 FILLER_71_1138 ();
 sg13g2_decap_4 FILLER_71_1145 ();
 sg13g2_decap_8 FILLER_71_1155 ();
 sg13g2_decap_8 FILLER_71_1162 ();
 sg13g2_fill_2 FILLER_71_1169 ();
 sg13g2_fill_1 FILLER_71_1171 ();
 sg13g2_decap_8 FILLER_71_1177 ();
 sg13g2_decap_8 FILLER_71_1184 ();
 sg13g2_decap_8 FILLER_71_1191 ();
 sg13g2_decap_4 FILLER_71_1198 ();
 sg13g2_fill_2 FILLER_71_1202 ();
 sg13g2_decap_8 FILLER_71_1208 ();
 sg13g2_decap_8 FILLER_71_1215 ();
 sg13g2_decap_8 FILLER_71_1222 ();
 sg13g2_decap_4 FILLER_71_1229 ();
 sg13g2_decap_8 FILLER_71_1256 ();
 sg13g2_decap_8 FILLER_71_1263 ();
 sg13g2_decap_8 FILLER_71_1270 ();
 sg13g2_decap_8 FILLER_71_1277 ();
 sg13g2_decap_8 FILLER_71_1284 ();
 sg13g2_decap_8 FILLER_71_1291 ();
 sg13g2_decap_8 FILLER_71_1298 ();
 sg13g2_decap_4 FILLER_71_1313 ();
 sg13g2_fill_2 FILLER_71_1345 ();
 sg13g2_fill_1 FILLER_71_1347 ();
 sg13g2_decap_8 FILLER_71_1354 ();
 sg13g2_decap_8 FILLER_71_1361 ();
 sg13g2_decap_4 FILLER_71_1368 ();
 sg13g2_fill_2 FILLER_71_1372 ();
 sg13g2_fill_2 FILLER_71_1380 ();
 sg13g2_fill_2 FILLER_71_1395 ();
 sg13g2_fill_1 FILLER_71_1397 ();
 sg13g2_decap_8 FILLER_71_1424 ();
 sg13g2_decap_8 FILLER_71_1431 ();
 sg13g2_decap_8 FILLER_71_1438 ();
 sg13g2_decap_8 FILLER_71_1481 ();
 sg13g2_decap_8 FILLER_71_1488 ();
 sg13g2_decap_8 FILLER_71_1495 ();
 sg13g2_decap_8 FILLER_71_1502 ();
 sg13g2_fill_1 FILLER_71_1509 ();
 sg13g2_decap_8 FILLER_71_1542 ();
 sg13g2_decap_8 FILLER_71_1549 ();
 sg13g2_decap_8 FILLER_71_1556 ();
 sg13g2_decap_8 FILLER_71_1576 ();
 sg13g2_fill_1 FILLER_71_1583 ();
 sg13g2_decap_8 FILLER_71_1590 ();
 sg13g2_decap_8 FILLER_71_1597 ();
 sg13g2_decap_4 FILLER_71_1604 ();
 sg13g2_fill_1 FILLER_71_1624 ();
 sg13g2_decap_8 FILLER_71_1651 ();
 sg13g2_decap_8 FILLER_71_1658 ();
 sg13g2_fill_2 FILLER_71_1665 ();
 sg13g2_decap_4 FILLER_71_1680 ();
 sg13g2_fill_1 FILLER_71_1684 ();
 sg13g2_decap_8 FILLER_71_1695 ();
 sg13g2_decap_8 FILLER_71_1702 ();
 sg13g2_decap_4 FILLER_71_1709 ();
 sg13g2_fill_1 FILLER_71_1713 ();
 sg13g2_decap_4 FILLER_71_1718 ();
 sg13g2_fill_1 FILLER_71_1722 ();
 sg13g2_decap_8 FILLER_71_1731 ();
 sg13g2_decap_8 FILLER_71_1738 ();
 sg13g2_decap_8 FILLER_71_1745 ();
 sg13g2_decap_4 FILLER_71_1752 ();
 sg13g2_fill_1 FILLER_71_1756 ();
 sg13g2_decap_8 FILLER_71_1783 ();
 sg13g2_decap_8 FILLER_71_1790 ();
 sg13g2_decap_8 FILLER_71_1797 ();
 sg13g2_decap_8 FILLER_71_1804 ();
 sg13g2_decap_8 FILLER_71_1811 ();
 sg13g2_decap_8 FILLER_71_1818 ();
 sg13g2_decap_8 FILLER_71_1825 ();
 sg13g2_decap_8 FILLER_71_1832 ();
 sg13g2_decap_8 FILLER_71_1839 ();
 sg13g2_decap_8 FILLER_71_1846 ();
 sg13g2_decap_8 FILLER_71_1853 ();
 sg13g2_decap_8 FILLER_71_1860 ();
 sg13g2_decap_8 FILLER_71_1867 ();
 sg13g2_decap_8 FILLER_71_1874 ();
 sg13g2_decap_8 FILLER_71_1881 ();
 sg13g2_decap_8 FILLER_71_1888 ();
 sg13g2_decap_8 FILLER_71_1895 ();
 sg13g2_decap_8 FILLER_71_1902 ();
 sg13g2_decap_8 FILLER_71_1909 ();
 sg13g2_decap_4 FILLER_71_1916 ();
 sg13g2_fill_2 FILLER_71_1920 ();
 sg13g2_decap_8 FILLER_71_1926 ();
 sg13g2_decap_8 FILLER_71_1933 ();
 sg13g2_decap_8 FILLER_71_1940 ();
 sg13g2_decap_8 FILLER_71_1947 ();
 sg13g2_decap_8 FILLER_71_1974 ();
 sg13g2_decap_8 FILLER_71_1981 ();
 sg13g2_decap_8 FILLER_71_1988 ();
 sg13g2_decap_8 FILLER_71_1995 ();
 sg13g2_decap_8 FILLER_71_2002 ();
 sg13g2_decap_4 FILLER_71_2009 ();
 sg13g2_fill_1 FILLER_71_2013 ();
 sg13g2_decap_8 FILLER_71_2024 ();
 sg13g2_fill_2 FILLER_71_2031 ();
 sg13g2_fill_1 FILLER_71_2033 ();
 sg13g2_fill_2 FILLER_71_2039 ();
 sg13g2_decap_8 FILLER_71_2056 ();
 sg13g2_decap_8 FILLER_71_2063 ();
 sg13g2_decap_8 FILLER_71_2070 ();
 sg13g2_decap_8 FILLER_71_2077 ();
 sg13g2_decap_8 FILLER_71_2084 ();
 sg13g2_decap_8 FILLER_71_2091 ();
 sg13g2_decap_8 FILLER_71_2098 ();
 sg13g2_decap_8 FILLER_71_2105 ();
 sg13g2_decap_8 FILLER_71_2112 ();
 sg13g2_decap_8 FILLER_71_2119 ();
 sg13g2_fill_2 FILLER_71_2126 ();
 sg13g2_fill_1 FILLER_71_2128 ();
 sg13g2_decap_8 FILLER_71_2139 ();
 sg13g2_decap_8 FILLER_71_2146 ();
 sg13g2_decap_8 FILLER_71_2153 ();
 sg13g2_decap_8 FILLER_71_2160 ();
 sg13g2_decap_8 FILLER_71_2167 ();
 sg13g2_decap_8 FILLER_71_2174 ();
 sg13g2_decap_8 FILLER_71_2181 ();
 sg13g2_decap_8 FILLER_71_2188 ();
 sg13g2_decap_8 FILLER_71_2195 ();
 sg13g2_fill_2 FILLER_71_2202 ();
 sg13g2_fill_1 FILLER_71_2204 ();
 sg13g2_decap_8 FILLER_71_2216 ();
 sg13g2_decap_8 FILLER_71_2223 ();
 sg13g2_decap_8 FILLER_71_2230 ();
 sg13g2_decap_8 FILLER_71_2237 ();
 sg13g2_decap_8 FILLER_71_2244 ();
 sg13g2_decap_8 FILLER_71_2251 ();
 sg13g2_decap_8 FILLER_71_2258 ();
 sg13g2_decap_8 FILLER_71_2265 ();
 sg13g2_decap_8 FILLER_71_2272 ();
 sg13g2_decap_8 FILLER_71_2279 ();
 sg13g2_decap_8 FILLER_71_2286 ();
 sg13g2_decap_8 FILLER_71_2293 ();
 sg13g2_decap_8 FILLER_71_2300 ();
 sg13g2_decap_8 FILLER_71_2307 ();
 sg13g2_decap_8 FILLER_71_2314 ();
 sg13g2_decap_8 FILLER_71_2321 ();
 sg13g2_decap_8 FILLER_71_2328 ();
 sg13g2_fill_1 FILLER_71_2335 ();
 sg13g2_fill_2 FILLER_71_2341 ();
 sg13g2_decap_8 FILLER_71_2358 ();
 sg13g2_decap_8 FILLER_71_2365 ();
 sg13g2_decap_8 FILLER_71_2372 ();
 sg13g2_decap_8 FILLER_71_2379 ();
 sg13g2_decap_8 FILLER_71_2386 ();
 sg13g2_decap_8 FILLER_71_2393 ();
 sg13g2_decap_4 FILLER_71_2400 ();
 sg13g2_fill_1 FILLER_71_2419 ();
 sg13g2_decap_8 FILLER_71_2425 ();
 sg13g2_fill_2 FILLER_71_2432 ();
 sg13g2_decap_8 FILLER_71_2438 ();
 sg13g2_fill_1 FILLER_71_2445 ();
 sg13g2_decap_8 FILLER_71_2455 ();
 sg13g2_decap_8 FILLER_71_2462 ();
 sg13g2_decap_8 FILLER_71_2469 ();
 sg13g2_decap_8 FILLER_71_2476 ();
 sg13g2_decap_8 FILLER_71_2483 ();
 sg13g2_decap_8 FILLER_71_2490 ();
 sg13g2_fill_1 FILLER_71_2497 ();
 sg13g2_decap_8 FILLER_71_2503 ();
 sg13g2_decap_8 FILLER_71_2510 ();
 sg13g2_decap_8 FILLER_71_2517 ();
 sg13g2_decap_4 FILLER_71_2524 ();
 sg13g2_decap_8 FILLER_71_2608 ();
 sg13g2_fill_1 FILLER_71_2615 ();
 sg13g2_fill_2 FILLER_71_2621 ();
 sg13g2_decap_8 FILLER_71_2626 ();
 sg13g2_decap_8 FILLER_71_2633 ();
 sg13g2_decap_8 FILLER_71_2640 ();
 sg13g2_decap_8 FILLER_71_2647 ();
 sg13g2_decap_4 FILLER_71_2654 ();
 sg13g2_fill_1 FILLER_71_2658 ();
 sg13g2_decap_8 FILLER_71_2669 ();
 sg13g2_decap_8 FILLER_71_2676 ();
 sg13g2_fill_1 FILLER_71_2683 ();
 sg13g2_decap_8 FILLER_71_2694 ();
 sg13g2_decap_8 FILLER_71_2701 ();
 sg13g2_decap_8 FILLER_71_2708 ();
 sg13g2_decap_8 FILLER_71_2715 ();
 sg13g2_decap_8 FILLER_71_2722 ();
 sg13g2_decap_8 FILLER_71_2729 ();
 sg13g2_decap_8 FILLER_71_2736 ();
 sg13g2_decap_4 FILLER_71_2743 ();
 sg13g2_fill_2 FILLER_71_2747 ();
 sg13g2_decap_4 FILLER_71_2758 ();
 sg13g2_fill_2 FILLER_71_2762 ();
 sg13g2_decap_4 FILLER_71_2769 ();
 sg13g2_fill_1 FILLER_71_2773 ();
 sg13g2_decap_8 FILLER_71_2784 ();
 sg13g2_decap_8 FILLER_71_2791 ();
 sg13g2_decap_4 FILLER_71_2798 ();
 sg13g2_fill_1 FILLER_71_2802 ();
 sg13g2_decap_4 FILLER_71_2812 ();
 sg13g2_fill_1 FILLER_71_2821 ();
 sg13g2_decap_4 FILLER_71_2837 ();
 sg13g2_fill_2 FILLER_71_2841 ();
 sg13g2_decap_8 FILLER_71_2848 ();
 sg13g2_fill_1 FILLER_71_2855 ();
 sg13g2_fill_1 FILLER_71_2866 ();
 sg13g2_decap_8 FILLER_71_2893 ();
 sg13g2_decap_8 FILLER_71_2900 ();
 sg13g2_decap_8 FILLER_71_2907 ();
 sg13g2_decap_8 FILLER_71_2914 ();
 sg13g2_decap_8 FILLER_71_2921 ();
 sg13g2_decap_8 FILLER_71_2928 ();
 sg13g2_fill_2 FILLER_71_2935 ();
 sg13g2_fill_1 FILLER_71_2937 ();
 sg13g2_decap_8 FILLER_71_2950 ();
 sg13g2_decap_8 FILLER_71_2957 ();
 sg13g2_decap_8 FILLER_71_2969 ();
 sg13g2_decap_8 FILLER_71_2976 ();
 sg13g2_decap_8 FILLER_71_2983 ();
 sg13g2_decap_8 FILLER_71_2990 ();
 sg13g2_decap_8 FILLER_71_2997 ();
 sg13g2_decap_8 FILLER_71_3004 ();
 sg13g2_decap_8 FILLER_71_3011 ();
 sg13g2_decap_4 FILLER_71_3018 ();
 sg13g2_decap_8 FILLER_71_3027 ();
 sg13g2_decap_8 FILLER_71_3034 ();
 sg13g2_decap_8 FILLER_71_3041 ();
 sg13g2_decap_8 FILLER_71_3048 ();
 sg13g2_decap_4 FILLER_71_3055 ();
 sg13g2_decap_8 FILLER_71_3064 ();
 sg13g2_decap_8 FILLER_71_3071 ();
 sg13g2_decap_8 FILLER_71_3078 ();
 sg13g2_decap_8 FILLER_71_3085 ();
 sg13g2_decap_8 FILLER_71_3092 ();
 sg13g2_decap_8 FILLER_71_3099 ();
 sg13g2_decap_8 FILLER_71_3106 ();
 sg13g2_decap_4 FILLER_71_3113 ();
 sg13g2_fill_2 FILLER_71_3117 ();
 sg13g2_decap_8 FILLER_71_3124 ();
 sg13g2_decap_8 FILLER_71_3166 ();
 sg13g2_decap_8 FILLER_71_3173 ();
 sg13g2_decap_4 FILLER_71_3180 ();
 sg13g2_fill_1 FILLER_71_3184 ();
 sg13g2_fill_2 FILLER_71_3189 ();
 sg13g2_decap_8 FILLER_71_3210 ();
 sg13g2_decap_4 FILLER_71_3217 ();
 sg13g2_decap_8 FILLER_71_3252 ();
 sg13g2_decap_4 FILLER_71_3259 ();
 sg13g2_fill_2 FILLER_71_3268 ();
 sg13g2_fill_1 FILLER_71_3270 ();
 sg13g2_decap_4 FILLER_71_3286 ();
 sg13g2_fill_2 FILLER_71_3290 ();
 sg13g2_decap_8 FILLER_71_3302 ();
 sg13g2_decap_4 FILLER_71_3309 ();
 sg13g2_decap_8 FILLER_71_3318 ();
 sg13g2_decap_8 FILLER_71_3325 ();
 sg13g2_decap_8 FILLER_71_3332 ();
 sg13g2_decap_8 FILLER_71_3339 ();
 sg13g2_decap_8 FILLER_71_3346 ();
 sg13g2_decap_8 FILLER_71_3353 ();
 sg13g2_decap_8 FILLER_71_3360 ();
 sg13g2_decap_8 FILLER_71_3367 ();
 sg13g2_decap_8 FILLER_71_3374 ();
 sg13g2_decap_8 FILLER_71_3381 ();
 sg13g2_decap_8 FILLER_71_3388 ();
 sg13g2_decap_8 FILLER_71_3395 ();
 sg13g2_decap_8 FILLER_71_3402 ();
 sg13g2_decap_8 FILLER_71_3409 ();
 sg13g2_decap_8 FILLER_71_3416 ();
 sg13g2_decap_4 FILLER_71_3449 ();
 sg13g2_decap_8 FILLER_71_3487 ();
 sg13g2_fill_2 FILLER_71_3494 ();
 sg13g2_fill_1 FILLER_71_3496 ();
 sg13g2_decap_8 FILLER_71_3523 ();
 sg13g2_decap_8 FILLER_71_3530 ();
 sg13g2_decap_8 FILLER_71_3537 ();
 sg13g2_decap_8 FILLER_71_3544 ();
 sg13g2_decap_8 FILLER_71_3551 ();
 sg13g2_decap_8 FILLER_71_3558 ();
 sg13g2_decap_8 FILLER_71_3565 ();
 sg13g2_decap_8 FILLER_71_3572 ();
 sg13g2_fill_1 FILLER_71_3579 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_fill_1 FILLER_72_14 ();
 sg13g2_decap_8 FILLER_72_41 ();
 sg13g2_decap_8 FILLER_72_48 ();
 sg13g2_decap_8 FILLER_72_55 ();
 sg13g2_decap_8 FILLER_72_62 ();
 sg13g2_fill_1 FILLER_72_69 ();
 sg13g2_decap_4 FILLER_72_78 ();
 sg13g2_decap_8 FILLER_72_90 ();
 sg13g2_decap_8 FILLER_72_97 ();
 sg13g2_decap_8 FILLER_72_104 ();
 sg13g2_decap_8 FILLER_72_111 ();
 sg13g2_decap_4 FILLER_72_118 ();
 sg13g2_fill_1 FILLER_72_122 ();
 sg13g2_decap_8 FILLER_72_144 ();
 sg13g2_decap_8 FILLER_72_151 ();
 sg13g2_fill_2 FILLER_72_158 ();
 sg13g2_decap_8 FILLER_72_200 ();
 sg13g2_decap_8 FILLER_72_207 ();
 sg13g2_decap_8 FILLER_72_214 ();
 sg13g2_fill_1 FILLER_72_221 ();
 sg13g2_decap_8 FILLER_72_230 ();
 sg13g2_fill_2 FILLER_72_237 ();
 sg13g2_decap_8 FILLER_72_265 ();
 sg13g2_fill_1 FILLER_72_272 ();
 sg13g2_decap_4 FILLER_72_291 ();
 sg13g2_decap_8 FILLER_72_321 ();
 sg13g2_decap_8 FILLER_72_328 ();
 sg13g2_decap_8 FILLER_72_335 ();
 sg13g2_decap_8 FILLER_72_342 ();
 sg13g2_decap_8 FILLER_72_349 ();
 sg13g2_fill_2 FILLER_72_356 ();
 sg13g2_fill_1 FILLER_72_358 ();
 sg13g2_decap_8 FILLER_72_364 ();
 sg13g2_decap_8 FILLER_72_371 ();
 sg13g2_fill_2 FILLER_72_389 ();
 sg13g2_decap_8 FILLER_72_404 ();
 sg13g2_decap_8 FILLER_72_411 ();
 sg13g2_decap_8 FILLER_72_418 ();
 sg13g2_decap_4 FILLER_72_425 ();
 sg13g2_fill_2 FILLER_72_429 ();
 sg13g2_fill_1 FILLER_72_438 ();
 sg13g2_decap_8 FILLER_72_447 ();
 sg13g2_decap_8 FILLER_72_454 ();
 sg13g2_decap_8 FILLER_72_461 ();
 sg13g2_decap_8 FILLER_72_468 ();
 sg13g2_decap_4 FILLER_72_475 ();
 sg13g2_decap_8 FILLER_72_503 ();
 sg13g2_decap_8 FILLER_72_510 ();
 sg13g2_decap_8 FILLER_72_517 ();
 sg13g2_decap_8 FILLER_72_524 ();
 sg13g2_decap_8 FILLER_72_531 ();
 sg13g2_decap_8 FILLER_72_538 ();
 sg13g2_decap_8 FILLER_72_545 ();
 sg13g2_fill_1 FILLER_72_552 ();
 sg13g2_decap_8 FILLER_72_566 ();
 sg13g2_decap_8 FILLER_72_573 ();
 sg13g2_fill_2 FILLER_72_580 ();
 sg13g2_decap_8 FILLER_72_626 ();
 sg13g2_fill_1 FILLER_72_633 ();
 sg13g2_decap_4 FILLER_72_659 ();
 sg13g2_fill_1 FILLER_72_663 ();
 sg13g2_decap_8 FILLER_72_687 ();
 sg13g2_fill_2 FILLER_72_694 ();
 sg13g2_fill_1 FILLER_72_700 ();
 sg13g2_fill_1 FILLER_72_706 ();
 sg13g2_decap_8 FILLER_72_721 ();
 sg13g2_decap_8 FILLER_72_728 ();
 sg13g2_decap_4 FILLER_72_735 ();
 sg13g2_fill_2 FILLER_72_739 ();
 sg13g2_decap_8 FILLER_72_746 ();
 sg13g2_decap_8 FILLER_72_753 ();
 sg13g2_decap_8 FILLER_72_760 ();
 sg13g2_decap_8 FILLER_72_767 ();
 sg13g2_decap_8 FILLER_72_774 ();
 sg13g2_decap_8 FILLER_72_803 ();
 sg13g2_decap_4 FILLER_72_810 ();
 sg13g2_fill_2 FILLER_72_814 ();
 sg13g2_fill_2 FILLER_72_825 ();
 sg13g2_fill_1 FILLER_72_831 ();
 sg13g2_decap_4 FILLER_72_837 ();
 sg13g2_fill_1 FILLER_72_841 ();
 sg13g2_fill_1 FILLER_72_852 ();
 sg13g2_decap_8 FILLER_72_863 ();
 sg13g2_decap_8 FILLER_72_870 ();
 sg13g2_decap_8 FILLER_72_877 ();
 sg13g2_fill_2 FILLER_72_884 ();
 sg13g2_fill_1 FILLER_72_897 ();
 sg13g2_decap_8 FILLER_72_923 ();
 sg13g2_fill_2 FILLER_72_930 ();
 sg13g2_fill_1 FILLER_72_932 ();
 sg13g2_decap_8 FILLER_72_967 ();
 sg13g2_fill_1 FILLER_72_974 ();
 sg13g2_decap_8 FILLER_72_988 ();
 sg13g2_decap_8 FILLER_72_995 ();
 sg13g2_decap_8 FILLER_72_1002 ();
 sg13g2_fill_1 FILLER_72_1009 ();
 sg13g2_fill_1 FILLER_72_1015 ();
 sg13g2_fill_2 FILLER_72_1026 ();
 sg13g2_fill_1 FILLER_72_1028 ();
 sg13g2_decap_8 FILLER_72_1034 ();
 sg13g2_fill_2 FILLER_72_1041 ();
 sg13g2_fill_1 FILLER_72_1051 ();
 sg13g2_fill_2 FILLER_72_1062 ();
 sg13g2_fill_2 FILLER_72_1072 ();
 sg13g2_fill_1 FILLER_72_1074 ();
 sg13g2_decap_8 FILLER_72_1080 ();
 sg13g2_decap_8 FILLER_72_1087 ();
 sg13g2_decap_8 FILLER_72_1094 ();
 sg13g2_decap_8 FILLER_72_1101 ();
 sg13g2_decap_8 FILLER_72_1108 ();
 sg13g2_decap_8 FILLER_72_1115 ();
 sg13g2_decap_8 FILLER_72_1122 ();
 sg13g2_decap_8 FILLER_72_1129 ();
 sg13g2_decap_8 FILLER_72_1136 ();
 sg13g2_decap_8 FILLER_72_1143 ();
 sg13g2_decap_8 FILLER_72_1150 ();
 sg13g2_decap_4 FILLER_72_1157 ();
 sg13g2_fill_2 FILLER_72_1161 ();
 sg13g2_fill_1 FILLER_72_1178 ();
 sg13g2_decap_8 FILLER_72_1187 ();
 sg13g2_fill_1 FILLER_72_1194 ();
 sg13g2_decap_8 FILLER_72_1215 ();
 sg13g2_decap_4 FILLER_72_1222 ();
 sg13g2_decap_8 FILLER_72_1258 ();
 sg13g2_decap_8 FILLER_72_1265 ();
 sg13g2_decap_8 FILLER_72_1272 ();
 sg13g2_decap_8 FILLER_72_1279 ();
 sg13g2_decap_8 FILLER_72_1286 ();
 sg13g2_decap_8 FILLER_72_1293 ();
 sg13g2_decap_8 FILLER_72_1300 ();
 sg13g2_decap_8 FILLER_72_1307 ();
 sg13g2_decap_8 FILLER_72_1314 ();
 sg13g2_decap_8 FILLER_72_1321 ();
 sg13g2_decap_8 FILLER_72_1328 ();
 sg13g2_decap_8 FILLER_72_1335 ();
 sg13g2_decap_8 FILLER_72_1342 ();
 sg13g2_decap_8 FILLER_72_1349 ();
 sg13g2_decap_8 FILLER_72_1356 ();
 sg13g2_decap_4 FILLER_72_1363 ();
 sg13g2_fill_1 FILLER_72_1367 ();
 sg13g2_decap_8 FILLER_72_1434 ();
 sg13g2_decap_8 FILLER_72_1441 ();
 sg13g2_decap_8 FILLER_72_1448 ();
 sg13g2_decap_8 FILLER_72_1455 ();
 sg13g2_decap_4 FILLER_72_1462 ();
 sg13g2_decap_8 FILLER_72_1474 ();
 sg13g2_decap_8 FILLER_72_1481 ();
 sg13g2_decap_8 FILLER_72_1488 ();
 sg13g2_decap_8 FILLER_72_1495 ();
 sg13g2_decap_8 FILLER_72_1502 ();
 sg13g2_decap_8 FILLER_72_1509 ();
 sg13g2_decap_8 FILLER_72_1516 ();
 sg13g2_decap_8 FILLER_72_1523 ();
 sg13g2_decap_8 FILLER_72_1530 ();
 sg13g2_decap_8 FILLER_72_1537 ();
 sg13g2_fill_1 FILLER_72_1544 ();
 sg13g2_decap_8 FILLER_72_1576 ();
 sg13g2_decap_8 FILLER_72_1583 ();
 sg13g2_decap_8 FILLER_72_1590 ();
 sg13g2_decap_4 FILLER_72_1597 ();
 sg13g2_fill_1 FILLER_72_1614 ();
 sg13g2_decap_8 FILLER_72_1628 ();
 sg13g2_decap_8 FILLER_72_1635 ();
 sg13g2_decap_8 FILLER_72_1642 ();
 sg13g2_decap_8 FILLER_72_1649 ();
 sg13g2_decap_8 FILLER_72_1656 ();
 sg13g2_decap_8 FILLER_72_1663 ();
 sg13g2_fill_1 FILLER_72_1670 ();
 sg13g2_decap_8 FILLER_72_1697 ();
 sg13g2_decap_8 FILLER_72_1704 ();
 sg13g2_decap_8 FILLER_72_1711 ();
 sg13g2_decap_8 FILLER_72_1718 ();
 sg13g2_decap_8 FILLER_72_1751 ();
 sg13g2_decap_8 FILLER_72_1758 ();
 sg13g2_decap_8 FILLER_72_1765 ();
 sg13g2_decap_8 FILLER_72_1772 ();
 sg13g2_decap_8 FILLER_72_1779 ();
 sg13g2_decap_4 FILLER_72_1786 ();
 sg13g2_fill_1 FILLER_72_1790 ();
 sg13g2_decap_8 FILLER_72_1799 ();
 sg13g2_decap_8 FILLER_72_1806 ();
 sg13g2_decap_8 FILLER_72_1813 ();
 sg13g2_decap_8 FILLER_72_1820 ();
 sg13g2_decap_8 FILLER_72_1827 ();
 sg13g2_fill_2 FILLER_72_1834 ();
 sg13g2_fill_1 FILLER_72_1836 ();
 sg13g2_decap_8 FILLER_72_1873 ();
 sg13g2_fill_2 FILLER_72_1890 ();
 sg13g2_decap_8 FILLER_72_1933 ();
 sg13g2_decap_8 FILLER_72_1940 ();
 sg13g2_decap_8 FILLER_72_1947 ();
 sg13g2_fill_1 FILLER_72_1954 ();
 sg13g2_decap_8 FILLER_72_1981 ();
 sg13g2_decap_8 FILLER_72_1988 ();
 sg13g2_decap_8 FILLER_72_1995 ();
 sg13g2_decap_4 FILLER_72_2002 ();
 sg13g2_fill_1 FILLER_72_2006 ();
 sg13g2_decap_8 FILLER_72_2033 ();
 sg13g2_decap_8 FILLER_72_2040 ();
 sg13g2_decap_4 FILLER_72_2047 ();
 sg13g2_fill_1 FILLER_72_2051 ();
 sg13g2_decap_8 FILLER_72_2078 ();
 sg13g2_decap_8 FILLER_72_2089 ();
 sg13g2_decap_8 FILLER_72_2096 ();
 sg13g2_decap_4 FILLER_72_2103 ();
 sg13g2_fill_1 FILLER_72_2107 ();
 sg13g2_decap_8 FILLER_72_2118 ();
 sg13g2_fill_1 FILLER_72_2125 ();
 sg13g2_decap_8 FILLER_72_2152 ();
 sg13g2_decap_8 FILLER_72_2159 ();
 sg13g2_decap_8 FILLER_72_2166 ();
 sg13g2_decap_8 FILLER_72_2173 ();
 sg13g2_decap_8 FILLER_72_2180 ();
 sg13g2_decap_8 FILLER_72_2187 ();
 sg13g2_decap_4 FILLER_72_2194 ();
 sg13g2_fill_2 FILLER_72_2198 ();
 sg13g2_decap_8 FILLER_72_2211 ();
 sg13g2_decap_8 FILLER_72_2218 ();
 sg13g2_decap_8 FILLER_72_2225 ();
 sg13g2_decap_8 FILLER_72_2232 ();
 sg13g2_fill_1 FILLER_72_2239 ();
 sg13g2_decap_8 FILLER_72_2259 ();
 sg13g2_decap_8 FILLER_72_2266 ();
 sg13g2_decap_8 FILLER_72_2273 ();
 sg13g2_decap_4 FILLER_72_2280 ();
 sg13g2_fill_1 FILLER_72_2284 ();
 sg13g2_decap_8 FILLER_72_2309 ();
 sg13g2_decap_8 FILLER_72_2316 ();
 sg13g2_decap_8 FILLER_72_2323 ();
 sg13g2_fill_2 FILLER_72_2330 ();
 sg13g2_fill_1 FILLER_72_2332 ();
 sg13g2_decap_4 FILLER_72_2337 ();
 sg13g2_fill_1 FILLER_72_2341 ();
 sg13g2_decap_8 FILLER_72_2357 ();
 sg13g2_decap_8 FILLER_72_2364 ();
 sg13g2_decap_8 FILLER_72_2371 ();
 sg13g2_decap_8 FILLER_72_2378 ();
 sg13g2_decap_4 FILLER_72_2385 ();
 sg13g2_fill_2 FILLER_72_2389 ();
 sg13g2_decap_8 FILLER_72_2395 ();
 sg13g2_decap_8 FILLER_72_2402 ();
 sg13g2_decap_8 FILLER_72_2409 ();
 sg13g2_decap_8 FILLER_72_2416 ();
 sg13g2_decap_8 FILLER_72_2423 ();
 sg13g2_decap_8 FILLER_72_2456 ();
 sg13g2_fill_2 FILLER_72_2463 ();
 sg13g2_decap_4 FILLER_72_2475 ();
 sg13g2_fill_2 FILLER_72_2479 ();
 sg13g2_decap_8 FILLER_72_2486 ();
 sg13g2_decap_8 FILLER_72_2493 ();
 sg13g2_decap_8 FILLER_72_2500 ();
 sg13g2_decap_8 FILLER_72_2507 ();
 sg13g2_decap_8 FILLER_72_2514 ();
 sg13g2_decap_8 FILLER_72_2521 ();
 sg13g2_decap_8 FILLER_72_2528 ();
 sg13g2_decap_8 FILLER_72_2535 ();
 sg13g2_fill_1 FILLER_72_2542 ();
 sg13g2_decap_4 FILLER_72_2553 ();
 sg13g2_fill_2 FILLER_72_2557 ();
 sg13g2_fill_2 FILLER_72_2563 ();
 sg13g2_fill_1 FILLER_72_2565 ();
 sg13g2_decap_4 FILLER_72_2575 ();
 sg13g2_fill_1 FILLER_72_2579 ();
 sg13g2_decap_8 FILLER_72_2589 ();
 sg13g2_decap_8 FILLER_72_2596 ();
 sg13g2_decap_4 FILLER_72_2603 ();
 sg13g2_decap_8 FILLER_72_2642 ();
 sg13g2_fill_2 FILLER_72_2649 ();
 sg13g2_decap_4 FILLER_72_2703 ();
 sg13g2_fill_1 FILLER_72_2707 ();
 sg13g2_fill_2 FILLER_72_2712 ();
 sg13g2_fill_1 FILLER_72_2714 ();
 sg13g2_decap_8 FILLER_72_2719 ();
 sg13g2_decap_8 FILLER_72_2726 ();
 sg13g2_decap_8 FILLER_72_2787 ();
 sg13g2_fill_2 FILLER_72_2804 ();
 sg13g2_decap_8 FILLER_72_2837 ();
 sg13g2_decap_8 FILLER_72_2844 ();
 sg13g2_decap_8 FILLER_72_2851 ();
 sg13g2_decap_4 FILLER_72_2861 ();
 sg13g2_fill_1 FILLER_72_2865 ();
 sg13g2_decap_8 FILLER_72_2871 ();
 sg13g2_decap_8 FILLER_72_2878 ();
 sg13g2_decap_8 FILLER_72_2885 ();
 sg13g2_decap_8 FILLER_72_2892 ();
 sg13g2_decap_8 FILLER_72_2899 ();
 sg13g2_decap_4 FILLER_72_2906 ();
 sg13g2_fill_2 FILLER_72_2910 ();
 sg13g2_decap_4 FILLER_72_2938 ();
 sg13g2_fill_2 FILLER_72_2942 ();
 sg13g2_decap_8 FILLER_72_2951 ();
 sg13g2_decap_8 FILLER_72_2972 ();
 sg13g2_decap_8 FILLER_72_2979 ();
 sg13g2_decap_8 FILLER_72_2986 ();
 sg13g2_decap_8 FILLER_72_2993 ();
 sg13g2_decap_8 FILLER_72_3000 ();
 sg13g2_decap_4 FILLER_72_3007 ();
 sg13g2_fill_2 FILLER_72_3011 ();
 sg13g2_decap_8 FILLER_72_3031 ();
 sg13g2_decap_8 FILLER_72_3038 ();
 sg13g2_decap_8 FILLER_72_3045 ();
 sg13g2_decap_8 FILLER_72_3052 ();
 sg13g2_decap_8 FILLER_72_3059 ();
 sg13g2_fill_1 FILLER_72_3066 ();
 sg13g2_fill_1 FILLER_72_3077 ();
 sg13g2_fill_2 FILLER_72_3083 ();
 sg13g2_fill_1 FILLER_72_3085 ();
 sg13g2_decap_8 FILLER_72_3096 ();
 sg13g2_fill_1 FILLER_72_3103 ();
 sg13g2_fill_1 FILLER_72_3114 ();
 sg13g2_decap_4 FILLER_72_3120 ();
 sg13g2_decap_8 FILLER_72_3129 ();
 sg13g2_decap_8 FILLER_72_3136 ();
 sg13g2_fill_2 FILLER_72_3143 ();
 sg13g2_decap_8 FILLER_72_3149 ();
 sg13g2_decap_8 FILLER_72_3156 ();
 sg13g2_decap_8 FILLER_72_3163 ();
 sg13g2_decap_8 FILLER_72_3170 ();
 sg13g2_fill_2 FILLER_72_3177 ();
 sg13g2_fill_1 FILLER_72_3179 ();
 sg13g2_decap_8 FILLER_72_3206 ();
 sg13g2_fill_2 FILLER_72_3213 ();
 sg13g2_decap_8 FILLER_72_3225 ();
 sg13g2_decap_8 FILLER_72_3232 ();
 sg13g2_decap_8 FILLER_72_3239 ();
 sg13g2_decap_8 FILLER_72_3246 ();
 sg13g2_decap_4 FILLER_72_3253 ();
 sg13g2_fill_1 FILLER_72_3257 ();
 sg13g2_fill_2 FILLER_72_3284 ();
 sg13g2_decap_8 FILLER_72_3317 ();
 sg13g2_decap_8 FILLER_72_3324 ();
 sg13g2_decap_8 FILLER_72_3331 ();
 sg13g2_fill_2 FILLER_72_3338 ();
 sg13g2_fill_1 FILLER_72_3340 ();
 sg13g2_fill_1 FILLER_72_3362 ();
 sg13g2_decap_4 FILLER_72_3376 ();
 sg13g2_fill_1 FILLER_72_3380 ();
 sg13g2_decap_8 FILLER_72_3391 ();
 sg13g2_decap_8 FILLER_72_3398 ();
 sg13g2_fill_2 FILLER_72_3405 ();
 sg13g2_decap_8 FILLER_72_3412 ();
 sg13g2_decap_8 FILLER_72_3419 ();
 sg13g2_decap_8 FILLER_72_3426 ();
 sg13g2_decap_8 FILLER_72_3433 ();
 sg13g2_decap_8 FILLER_72_3440 ();
 sg13g2_decap_8 FILLER_72_3447 ();
 sg13g2_decap_8 FILLER_72_3454 ();
 sg13g2_decap_8 FILLER_72_3461 ();
 sg13g2_decap_8 FILLER_72_3468 ();
 sg13g2_decap_8 FILLER_72_3475 ();
 sg13g2_decap_8 FILLER_72_3482 ();
 sg13g2_decap_8 FILLER_72_3489 ();
 sg13g2_decap_8 FILLER_72_3496 ();
 sg13g2_decap_8 FILLER_72_3503 ();
 sg13g2_decap_8 FILLER_72_3510 ();
 sg13g2_decap_8 FILLER_72_3517 ();
 sg13g2_decap_8 FILLER_72_3524 ();
 sg13g2_decap_8 FILLER_72_3531 ();
 sg13g2_decap_8 FILLER_72_3538 ();
 sg13g2_decap_8 FILLER_72_3545 ();
 sg13g2_decap_8 FILLER_72_3552 ();
 sg13g2_decap_8 FILLER_72_3559 ();
 sg13g2_decap_8 FILLER_72_3566 ();
 sg13g2_decap_8 FILLER_72_3573 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_4 FILLER_73_7 ();
 sg13g2_decap_4 FILLER_73_57 ();
 sg13g2_fill_1 FILLER_73_61 ();
 sg13g2_decap_8 FILLER_73_86 ();
 sg13g2_decap_8 FILLER_73_93 ();
 sg13g2_decap_8 FILLER_73_100 ();
 sg13g2_decap_4 FILLER_73_107 ();
 sg13g2_fill_2 FILLER_73_111 ();
 sg13g2_decap_8 FILLER_73_162 ();
 sg13g2_fill_1 FILLER_73_169 ();
 sg13g2_decap_8 FILLER_73_175 ();
 sg13g2_decap_8 FILLER_73_182 ();
 sg13g2_decap_8 FILLER_73_189 ();
 sg13g2_decap_8 FILLER_73_196 ();
 sg13g2_decap_8 FILLER_73_203 ();
 sg13g2_decap_8 FILLER_73_210 ();
 sg13g2_decap_8 FILLER_73_217 ();
 sg13g2_decap_8 FILLER_73_232 ();
 sg13g2_decap_8 FILLER_73_239 ();
 sg13g2_decap_8 FILLER_73_246 ();
 sg13g2_decap_4 FILLER_73_253 ();
 sg13g2_fill_1 FILLER_73_257 ();
 sg13g2_decap_4 FILLER_73_266 ();
 sg13g2_fill_2 FILLER_73_270 ();
 sg13g2_fill_1 FILLER_73_285 ();
 sg13g2_fill_2 FILLER_73_296 ();
 sg13g2_fill_1 FILLER_73_298 ();
 sg13g2_fill_2 FILLER_73_312 ();
 sg13g2_decap_8 FILLER_73_323 ();
 sg13g2_fill_2 FILLER_73_330 ();
 sg13g2_fill_1 FILLER_73_332 ();
 sg13g2_decap_8 FILLER_73_337 ();
 sg13g2_decap_8 FILLER_73_344 ();
 sg13g2_decap_8 FILLER_73_351 ();
 sg13g2_decap_8 FILLER_73_358 ();
 sg13g2_decap_8 FILLER_73_365 ();
 sg13g2_decap_8 FILLER_73_406 ();
 sg13g2_decap_8 FILLER_73_413 ();
 sg13g2_decap_8 FILLER_73_420 ();
 sg13g2_decap_8 FILLER_73_427 ();
 sg13g2_decap_4 FILLER_73_434 ();
 sg13g2_decap_8 FILLER_73_448 ();
 sg13g2_decap_4 FILLER_73_455 ();
 sg13g2_decap_8 FILLER_73_469 ();
 sg13g2_decap_8 FILLER_73_476 ();
 sg13g2_fill_2 FILLER_73_483 ();
 sg13g2_decap_8 FILLER_73_495 ();
 sg13g2_decap_8 FILLER_73_502 ();
 sg13g2_decap_8 FILLER_73_509 ();
 sg13g2_fill_1 FILLER_73_516 ();
 sg13g2_decap_8 FILLER_73_568 ();
 sg13g2_decap_4 FILLER_73_575 ();
 sg13g2_fill_2 FILLER_73_579 ();
 sg13g2_decap_8 FILLER_73_597 ();
 sg13g2_decap_8 FILLER_73_604 ();
 sg13g2_fill_1 FILLER_73_611 ();
 sg13g2_fill_1 FILLER_73_618 ();
 sg13g2_decap_8 FILLER_73_624 ();
 sg13g2_decap_8 FILLER_73_631 ();
 sg13g2_decap_4 FILLER_73_638 ();
 sg13g2_fill_2 FILLER_73_642 ();
 sg13g2_fill_1 FILLER_73_653 ();
 sg13g2_decap_8 FILLER_73_662 ();
 sg13g2_decap_8 FILLER_73_669 ();
 sg13g2_decap_8 FILLER_73_676 ();
 sg13g2_decap_8 FILLER_73_683 ();
 sg13g2_fill_2 FILLER_73_690 ();
 sg13g2_decap_8 FILLER_73_718 ();
 sg13g2_decap_8 FILLER_73_725 ();
 sg13g2_decap_4 FILLER_73_732 ();
 sg13g2_fill_2 FILLER_73_736 ();
 sg13g2_fill_1 FILLER_73_748 ();
 sg13g2_decap_8 FILLER_73_757 ();
 sg13g2_decap_8 FILLER_73_764 ();
 sg13g2_decap_8 FILLER_73_771 ();
 sg13g2_decap_8 FILLER_73_778 ();
 sg13g2_fill_2 FILLER_73_785 ();
 sg13g2_decap_4 FILLER_73_816 ();
 sg13g2_fill_2 FILLER_73_820 ();
 sg13g2_decap_4 FILLER_73_846 ();
 sg13g2_fill_1 FILLER_73_850 ();
 sg13g2_decap_4 FILLER_73_864 ();
 sg13g2_fill_2 FILLER_73_868 ();
 sg13g2_fill_2 FILLER_73_900 ();
 sg13g2_fill_1 FILLER_73_902 ();
 sg13g2_decap_8 FILLER_73_915 ();
 sg13g2_decap_8 FILLER_73_922 ();
 sg13g2_decap_8 FILLER_73_929 ();
 sg13g2_fill_1 FILLER_73_936 ();
 sg13g2_decap_8 FILLER_73_956 ();
 sg13g2_fill_1 FILLER_73_963 ();
 sg13g2_fill_2 FILLER_73_973 ();
 sg13g2_fill_1 FILLER_73_975 ();
 sg13g2_decap_8 FILLER_73_986 ();
 sg13g2_fill_2 FILLER_73_993 ();
 sg13g2_fill_1 FILLER_73_995 ();
 sg13g2_decap_8 FILLER_73_1001 ();
 sg13g2_decap_8 FILLER_73_1008 ();
 sg13g2_fill_2 FILLER_73_1015 ();
 sg13g2_decap_4 FILLER_73_1043 ();
 sg13g2_fill_2 FILLER_73_1047 ();
 sg13g2_fill_2 FILLER_73_1057 ();
 sg13g2_fill_1 FILLER_73_1059 ();
 sg13g2_fill_1 FILLER_73_1068 ();
 sg13g2_decap_8 FILLER_73_1087 ();
 sg13g2_decap_8 FILLER_73_1094 ();
 sg13g2_decap_8 FILLER_73_1114 ();
 sg13g2_fill_1 FILLER_73_1121 ();
 sg13g2_decap_8 FILLER_73_1131 ();
 sg13g2_decap_4 FILLER_73_1138 ();
 sg13g2_fill_2 FILLER_73_1142 ();
 sg13g2_decap_8 FILLER_73_1157 ();
 sg13g2_decap_4 FILLER_73_1164 ();
 sg13g2_fill_1 FILLER_73_1168 ();
 sg13g2_decap_8 FILLER_73_1177 ();
 sg13g2_decap_8 FILLER_73_1184 ();
 sg13g2_decap_8 FILLER_73_1191 ();
 sg13g2_decap_8 FILLER_73_1198 ();
 sg13g2_decap_8 FILLER_73_1205 ();
 sg13g2_decap_4 FILLER_73_1212 ();
 sg13g2_fill_2 FILLER_73_1216 ();
 sg13g2_fill_2 FILLER_73_1236 ();
 sg13g2_decap_8 FILLER_73_1263 ();
 sg13g2_decap_8 FILLER_73_1270 ();
 sg13g2_fill_2 FILLER_73_1277 ();
 sg13g2_decap_8 FILLER_73_1283 ();
 sg13g2_decap_8 FILLER_73_1290 ();
 sg13g2_decap_8 FILLER_73_1297 ();
 sg13g2_decap_8 FILLER_73_1304 ();
 sg13g2_decap_8 FILLER_73_1311 ();
 sg13g2_decap_8 FILLER_73_1318 ();
 sg13g2_decap_8 FILLER_73_1325 ();
 sg13g2_decap_8 FILLER_73_1332 ();
 sg13g2_decap_8 FILLER_73_1339 ();
 sg13g2_decap_8 FILLER_73_1346 ();
 sg13g2_decap_4 FILLER_73_1353 ();
 sg13g2_fill_1 FILLER_73_1357 ();
 sg13g2_decap_8 FILLER_73_1426 ();
 sg13g2_decap_8 FILLER_73_1433 ();
 sg13g2_decap_8 FILLER_73_1440 ();
 sg13g2_decap_8 FILLER_73_1447 ();
 sg13g2_decap_8 FILLER_73_1454 ();
 sg13g2_decap_8 FILLER_73_1461 ();
 sg13g2_decap_8 FILLER_73_1468 ();
 sg13g2_decap_8 FILLER_73_1475 ();
 sg13g2_fill_2 FILLER_73_1482 ();
 sg13g2_fill_1 FILLER_73_1510 ();
 sg13g2_decap_8 FILLER_73_1524 ();
 sg13g2_decap_8 FILLER_73_1531 ();
 sg13g2_decap_8 FILLER_73_1538 ();
 sg13g2_decap_8 FILLER_73_1545 ();
 sg13g2_decap_8 FILLER_73_1552 ();
 sg13g2_decap_8 FILLER_73_1559 ();
 sg13g2_decap_8 FILLER_73_1566 ();
 sg13g2_decap_8 FILLER_73_1573 ();
 sg13g2_decap_8 FILLER_73_1580 ();
 sg13g2_decap_8 FILLER_73_1587 ();
 sg13g2_decap_4 FILLER_73_1594 ();
 sg13g2_fill_1 FILLER_73_1598 ();
 sg13g2_decap_4 FILLER_73_1609 ();
 sg13g2_fill_2 FILLER_73_1613 ();
 sg13g2_decap_8 FILLER_73_1627 ();
 sg13g2_fill_2 FILLER_73_1634 ();
 sg13g2_fill_1 FILLER_73_1636 ();
 sg13g2_decap_8 FILLER_73_1663 ();
 sg13g2_decap_8 FILLER_73_1680 ();
 sg13g2_decap_8 FILLER_73_1687 ();
 sg13g2_decap_8 FILLER_73_1694 ();
 sg13g2_decap_4 FILLER_73_1701 ();
 sg13g2_fill_1 FILLER_73_1705 ();
 sg13g2_decap_8 FILLER_73_1742 ();
 sg13g2_decap_8 FILLER_73_1749 ();
 sg13g2_decap_8 FILLER_73_1756 ();
 sg13g2_decap_8 FILLER_73_1763 ();
 sg13g2_decap_8 FILLER_73_1770 ();
 sg13g2_fill_2 FILLER_73_1777 ();
 sg13g2_decap_8 FILLER_73_1815 ();
 sg13g2_fill_1 FILLER_73_1822 ();
 sg13g2_decap_8 FILLER_73_1859 ();
 sg13g2_decap_8 FILLER_73_1866 ();
 sg13g2_decap_8 FILLER_73_1873 ();
 sg13g2_fill_1 FILLER_73_1916 ();
 sg13g2_decap_8 FILLER_73_1925 ();
 sg13g2_decap_8 FILLER_73_1940 ();
 sg13g2_decap_8 FILLER_73_1947 ();
 sg13g2_decap_4 FILLER_73_1954 ();
 sg13g2_fill_1 FILLER_73_1958 ();
 sg13g2_fill_2 FILLER_73_1995 ();
 sg13g2_fill_1 FILLER_73_1997 ();
 sg13g2_decap_8 FILLER_73_2035 ();
 sg13g2_decap_8 FILLER_73_2042 ();
 sg13g2_decap_8 FILLER_73_2049 ();
 sg13g2_decap_8 FILLER_73_2062 ();
 sg13g2_decap_8 FILLER_73_2069 ();
 sg13g2_fill_2 FILLER_73_2076 ();
 sg13g2_decap_4 FILLER_73_2096 ();
 sg13g2_fill_2 FILLER_73_2100 ();
 sg13g2_decap_8 FILLER_73_2106 ();
 sg13g2_fill_2 FILLER_73_2113 ();
 sg13g2_decap_8 FILLER_73_2141 ();
 sg13g2_decap_8 FILLER_73_2148 ();
 sg13g2_decap_8 FILLER_73_2155 ();
 sg13g2_decap_8 FILLER_73_2176 ();
 sg13g2_decap_8 FILLER_73_2183 ();
 sg13g2_decap_8 FILLER_73_2190 ();
 sg13g2_fill_2 FILLER_73_2197 ();
 sg13g2_fill_1 FILLER_73_2199 ();
 sg13g2_fill_2 FILLER_73_2211 ();
 sg13g2_fill_1 FILLER_73_2213 ();
 sg13g2_fill_2 FILLER_73_2230 ();
 sg13g2_decap_8 FILLER_73_2272 ();
 sg13g2_decap_8 FILLER_73_2279 ();
 sg13g2_fill_2 FILLER_73_2286 ();
 sg13g2_fill_1 FILLER_73_2288 ();
 sg13g2_decap_8 FILLER_73_2324 ();
 sg13g2_decap_4 FILLER_73_2331 ();
 sg13g2_fill_2 FILLER_73_2335 ();
 sg13g2_decap_8 FILLER_73_2372 ();
 sg13g2_decap_4 FILLER_73_2379 ();
 sg13g2_decap_8 FILLER_73_2425 ();
 sg13g2_decap_8 FILLER_73_2432 ();
 sg13g2_decap_8 FILLER_73_2439 ();
 sg13g2_decap_8 FILLER_73_2446 ();
 sg13g2_decap_8 FILLER_73_2453 ();
 sg13g2_decap_8 FILLER_73_2460 ();
 sg13g2_decap_4 FILLER_73_2467 ();
 sg13g2_decap_8 FILLER_73_2507 ();
 sg13g2_decap_8 FILLER_73_2514 ();
 sg13g2_decap_8 FILLER_73_2521 ();
 sg13g2_decap_8 FILLER_73_2528 ();
 sg13g2_decap_8 FILLER_73_2535 ();
 sg13g2_decap_8 FILLER_73_2542 ();
 sg13g2_decap_8 FILLER_73_2549 ();
 sg13g2_decap_8 FILLER_73_2556 ();
 sg13g2_fill_2 FILLER_73_2563 ();
 sg13g2_decap_8 FILLER_73_2576 ();
 sg13g2_decap_8 FILLER_73_2583 ();
 sg13g2_decap_8 FILLER_73_2590 ();
 sg13g2_fill_2 FILLER_73_2597 ();
 sg13g2_fill_1 FILLER_73_2599 ();
 sg13g2_decap_8 FILLER_73_2630 ();
 sg13g2_decap_8 FILLER_73_2637 ();
 sg13g2_decap_8 FILLER_73_2644 ();
 sg13g2_decap_4 FILLER_73_2651 ();
 sg13g2_fill_1 FILLER_73_2655 ();
 sg13g2_fill_1 FILLER_73_2661 ();
 sg13g2_fill_2 FILLER_73_2677 ();
 sg13g2_fill_1 FILLER_73_2684 ();
 sg13g2_decap_8 FILLER_73_2700 ();
 sg13g2_decap_4 FILLER_73_2707 ();
 sg13g2_decap_8 FILLER_73_2742 ();
 sg13g2_decap_8 FILLER_73_2783 ();
 sg13g2_decap_8 FILLER_73_2790 ();
 sg13g2_decap_8 FILLER_73_2802 ();
 sg13g2_decap_8 FILLER_73_2809 ();
 sg13g2_decap_4 FILLER_73_2816 ();
 sg13g2_decap_4 FILLER_73_2835 ();
 sg13g2_fill_2 FILLER_73_2839 ();
 sg13g2_decap_8 FILLER_73_2846 ();
 sg13g2_fill_2 FILLER_73_2853 ();
 sg13g2_decap_8 FILLER_73_2862 ();
 sg13g2_decap_8 FILLER_73_2869 ();
 sg13g2_decap_8 FILLER_73_2887 ();
 sg13g2_decap_8 FILLER_73_2894 ();
 sg13g2_fill_2 FILLER_73_2901 ();
 sg13g2_fill_1 FILLER_73_2903 ();
 sg13g2_decap_8 FILLER_73_2912 ();
 sg13g2_fill_2 FILLER_73_2919 ();
 sg13g2_fill_1 FILLER_73_2921 ();
 sg13g2_decap_8 FILLER_73_2932 ();
 sg13g2_decap_8 FILLER_73_2939 ();
 sg13g2_fill_1 FILLER_73_2946 ();
 sg13g2_fill_2 FILLER_73_2985 ();
 sg13g2_decap_4 FILLER_73_3053 ();
 sg13g2_decap_4 FILLER_73_3085 ();
 sg13g2_decap_8 FILLER_73_3110 ();
 sg13g2_decap_8 FILLER_73_3117 ();
 sg13g2_decap_4 FILLER_73_3124 ();
 sg13g2_fill_2 FILLER_73_3128 ();
 sg13g2_decap_8 FILLER_73_3165 ();
 sg13g2_decap_8 FILLER_73_3172 ();
 sg13g2_fill_2 FILLER_73_3193 ();
 sg13g2_decap_8 FILLER_73_3221 ();
 sg13g2_decap_8 FILLER_73_3228 ();
 sg13g2_decap_8 FILLER_73_3235 ();
 sg13g2_decap_8 FILLER_73_3242 ();
 sg13g2_decap_8 FILLER_73_3249 ();
 sg13g2_fill_2 FILLER_73_3256 ();
 sg13g2_fill_1 FILLER_73_3258 ();
 sg13g2_decap_8 FILLER_73_3295 ();
 sg13g2_decap_4 FILLER_73_3302 ();
 sg13g2_fill_1 FILLER_73_3306 ();
 sg13g2_decap_8 FILLER_73_3312 ();
 sg13g2_fill_2 FILLER_73_3319 ();
 sg13g2_fill_1 FILLER_73_3321 ();
 sg13g2_decap_8 FILLER_73_3326 ();
 sg13g2_decap_4 FILLER_73_3333 ();
 sg13g2_fill_2 FILLER_73_3337 ();
 sg13g2_decap_8 FILLER_73_3385 ();
 sg13g2_fill_2 FILLER_73_3392 ();
 sg13g2_decap_8 FILLER_73_3433 ();
 sg13g2_decap_8 FILLER_73_3440 ();
 sg13g2_fill_2 FILLER_73_3447 ();
 sg13g2_fill_1 FILLER_73_3449 ();
 sg13g2_decap_8 FILLER_73_3458 ();
 sg13g2_decap_8 FILLER_73_3465 ();
 sg13g2_decap_8 FILLER_73_3472 ();
 sg13g2_decap_8 FILLER_73_3479 ();
 sg13g2_decap_8 FILLER_73_3486 ();
 sg13g2_decap_8 FILLER_73_3493 ();
 sg13g2_decap_8 FILLER_73_3500 ();
 sg13g2_decap_8 FILLER_73_3507 ();
 sg13g2_decap_8 FILLER_73_3514 ();
 sg13g2_decap_8 FILLER_73_3521 ();
 sg13g2_decap_8 FILLER_73_3528 ();
 sg13g2_decap_8 FILLER_73_3535 ();
 sg13g2_decap_8 FILLER_73_3542 ();
 sg13g2_decap_8 FILLER_73_3549 ();
 sg13g2_decap_8 FILLER_73_3556 ();
 sg13g2_decap_8 FILLER_73_3563 ();
 sg13g2_decap_8 FILLER_73_3570 ();
 sg13g2_fill_2 FILLER_73_3577 ();
 sg13g2_fill_1 FILLER_73_3579 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_fill_1 FILLER_74_14 ();
 sg13g2_decap_8 FILLER_74_59 ();
 sg13g2_fill_2 FILLER_74_66 ();
 sg13g2_fill_1 FILLER_74_68 ();
 sg13g2_decap_8 FILLER_74_79 ();
 sg13g2_decap_8 FILLER_74_86 ();
 sg13g2_decap_8 FILLER_74_93 ();
 sg13g2_fill_2 FILLER_74_100 ();
 sg13g2_fill_1 FILLER_74_102 ();
 sg13g2_fill_1 FILLER_74_116 ();
 sg13g2_fill_2 FILLER_74_131 ();
 sg13g2_decap_8 FILLER_74_143 ();
 sg13g2_decap_8 FILLER_74_150 ();
 sg13g2_fill_2 FILLER_74_157 ();
 sg13g2_fill_1 FILLER_74_159 ();
 sg13g2_decap_8 FILLER_74_165 ();
 sg13g2_decap_8 FILLER_74_172 ();
 sg13g2_decap_8 FILLER_74_179 ();
 sg13g2_decap_8 FILLER_74_186 ();
 sg13g2_decap_8 FILLER_74_193 ();
 sg13g2_decap_8 FILLER_74_200 ();
 sg13g2_fill_1 FILLER_74_212 ();
 sg13g2_fill_2 FILLER_74_222 ();
 sg13g2_decap_8 FILLER_74_228 ();
 sg13g2_decap_8 FILLER_74_235 ();
 sg13g2_decap_8 FILLER_74_242 ();
 sg13g2_decap_4 FILLER_74_249 ();
 sg13g2_fill_1 FILLER_74_253 ();
 sg13g2_decap_8 FILLER_74_262 ();
 sg13g2_decap_8 FILLER_74_269 ();
 sg13g2_fill_1 FILLER_74_276 ();
 sg13g2_decap_4 FILLER_74_304 ();
 sg13g2_decap_4 FILLER_74_313 ();
 sg13g2_fill_1 FILLER_74_317 ();
 sg13g2_decap_8 FILLER_74_325 ();
 sg13g2_decap_4 FILLER_74_332 ();
 sg13g2_fill_1 FILLER_74_336 ();
 sg13g2_decap_8 FILLER_74_345 ();
 sg13g2_decap_8 FILLER_74_352 ();
 sg13g2_decap_8 FILLER_74_359 ();
 sg13g2_decap_8 FILLER_74_366 ();
 sg13g2_fill_2 FILLER_74_373 ();
 sg13g2_decap_8 FILLER_74_389 ();
 sg13g2_decap_8 FILLER_74_396 ();
 sg13g2_decap_8 FILLER_74_403 ();
 sg13g2_decap_8 FILLER_74_410 ();
 sg13g2_decap_8 FILLER_74_417 ();
 sg13g2_decap_8 FILLER_74_424 ();
 sg13g2_decap_8 FILLER_74_431 ();
 sg13g2_fill_2 FILLER_74_438 ();
 sg13g2_decap_8 FILLER_74_448 ();
 sg13g2_decap_8 FILLER_74_455 ();
 sg13g2_decap_8 FILLER_74_462 ();
 sg13g2_decap_4 FILLER_74_469 ();
 sg13g2_fill_2 FILLER_74_481 ();
 sg13g2_fill_1 FILLER_74_483 ();
 sg13g2_decap_8 FILLER_74_492 ();
 sg13g2_decap_8 FILLER_74_499 ();
 sg13g2_decap_8 FILLER_74_506 ();
 sg13g2_decap_4 FILLER_74_513 ();
 sg13g2_fill_1 FILLER_74_517 ();
 sg13g2_decap_4 FILLER_74_522 ();
 sg13g2_fill_2 FILLER_74_526 ();
 sg13g2_decap_8 FILLER_74_554 ();
 sg13g2_decap_8 FILLER_74_561 ();
 sg13g2_decap_8 FILLER_74_568 ();
 sg13g2_decap_8 FILLER_74_575 ();
 sg13g2_decap_8 FILLER_74_582 ();
 sg13g2_decap_8 FILLER_74_589 ();
 sg13g2_decap_8 FILLER_74_596 ();
 sg13g2_decap_8 FILLER_74_603 ();
 sg13g2_decap_4 FILLER_74_610 ();
 sg13g2_fill_1 FILLER_74_614 ();
 sg13g2_decap_8 FILLER_74_619 ();
 sg13g2_fill_1 FILLER_74_626 ();
 sg13g2_decap_8 FILLER_74_635 ();
 sg13g2_decap_8 FILLER_74_642 ();
 sg13g2_decap_8 FILLER_74_649 ();
 sg13g2_decap_8 FILLER_74_656 ();
 sg13g2_decap_8 FILLER_74_663 ();
 sg13g2_decap_8 FILLER_74_670 ();
 sg13g2_decap_8 FILLER_74_677 ();
 sg13g2_decap_8 FILLER_74_684 ();
 sg13g2_decap_8 FILLER_74_691 ();
 sg13g2_decap_8 FILLER_74_698 ();
 sg13g2_decap_8 FILLER_74_705 ();
 sg13g2_decap_8 FILLER_74_712 ();
 sg13g2_decap_8 FILLER_74_719 ();
 sg13g2_decap_8 FILLER_74_726 ();
 sg13g2_fill_2 FILLER_74_733 ();
 sg13g2_decap_8 FILLER_74_751 ();
 sg13g2_decap_8 FILLER_74_758 ();
 sg13g2_decap_8 FILLER_74_765 ();
 sg13g2_decap_8 FILLER_74_772 ();
 sg13g2_decap_8 FILLER_74_779 ();
 sg13g2_decap_4 FILLER_74_786 ();
 sg13g2_decap_4 FILLER_74_795 ();
 sg13g2_fill_2 FILLER_74_799 ();
 sg13g2_decap_8 FILLER_74_810 ();
 sg13g2_decap_8 FILLER_74_817 ();
 sg13g2_decap_8 FILLER_74_824 ();
 sg13g2_decap_4 FILLER_74_831 ();
 sg13g2_decap_8 FILLER_74_840 ();
 sg13g2_decap_8 FILLER_74_847 ();
 sg13g2_decap_8 FILLER_74_854 ();
 sg13g2_decap_8 FILLER_74_861 ();
 sg13g2_decap_4 FILLER_74_868 ();
 sg13g2_decap_8 FILLER_74_877 ();
 sg13g2_decap_8 FILLER_74_884 ();
 sg13g2_fill_2 FILLER_74_891 ();
 sg13g2_decap_8 FILLER_74_902 ();
 sg13g2_decap_8 FILLER_74_909 ();
 sg13g2_decap_8 FILLER_74_916 ();
 sg13g2_decap_8 FILLER_74_923 ();
 sg13g2_fill_2 FILLER_74_930 ();
 sg13g2_fill_1 FILLER_74_932 ();
 sg13g2_decap_8 FILLER_74_946 ();
 sg13g2_decap_8 FILLER_74_953 ();
 sg13g2_decap_8 FILLER_74_960 ();
 sg13g2_fill_2 FILLER_74_967 ();
 sg13g2_decap_8 FILLER_74_973 ();
 sg13g2_decap_8 FILLER_74_980 ();
 sg13g2_decap_8 FILLER_74_987 ();
 sg13g2_decap_8 FILLER_74_994 ();
 sg13g2_decap_8 FILLER_74_1001 ();
 sg13g2_decap_8 FILLER_74_1008 ();
 sg13g2_decap_8 FILLER_74_1015 ();
 sg13g2_decap_8 FILLER_74_1022 ();
 sg13g2_decap_8 FILLER_74_1029 ();
 sg13g2_decap_8 FILLER_74_1036 ();
 sg13g2_decap_8 FILLER_74_1043 ();
 sg13g2_decap_4 FILLER_74_1050 ();
 sg13g2_fill_1 FILLER_74_1054 ();
 sg13g2_decap_8 FILLER_74_1076 ();
 sg13g2_decap_8 FILLER_74_1083 ();
 sg13g2_decap_8 FILLER_74_1090 ();
 sg13g2_decap_8 FILLER_74_1097 ();
 sg13g2_decap_8 FILLER_74_1104 ();
 sg13g2_decap_8 FILLER_74_1137 ();
 sg13g2_decap_8 FILLER_74_1144 ();
 sg13g2_decap_8 FILLER_74_1151 ();
 sg13g2_decap_8 FILLER_74_1158 ();
 sg13g2_decap_8 FILLER_74_1165 ();
 sg13g2_decap_8 FILLER_74_1172 ();
 sg13g2_fill_2 FILLER_74_1183 ();
 sg13g2_decap_8 FILLER_74_1194 ();
 sg13g2_fill_2 FILLER_74_1201 ();
 sg13g2_fill_1 FILLER_74_1203 ();
 sg13g2_decap_8 FILLER_74_1209 ();
 sg13g2_decap_8 FILLER_74_1216 ();
 sg13g2_decap_4 FILLER_74_1223 ();
 sg13g2_fill_2 FILLER_74_1227 ();
 sg13g2_fill_2 FILLER_74_1234 ();
 sg13g2_decap_8 FILLER_74_1248 ();
 sg13g2_decap_8 FILLER_74_1255 ();
 sg13g2_decap_4 FILLER_74_1262 ();
 sg13g2_decap_8 FILLER_74_1273 ();
 sg13g2_decap_8 FILLER_74_1280 ();
 sg13g2_fill_1 FILLER_74_1287 ();
 sg13g2_decap_8 FILLER_74_1308 ();
 sg13g2_decap_8 FILLER_74_1315 ();
 sg13g2_decap_8 FILLER_74_1322 ();
 sg13g2_decap_8 FILLER_74_1329 ();
 sg13g2_decap_4 FILLER_74_1336 ();
 sg13g2_fill_2 FILLER_74_1340 ();
 sg13g2_decap_8 FILLER_74_1421 ();
 sg13g2_decap_8 FILLER_74_1428 ();
 sg13g2_decap_8 FILLER_74_1435 ();
 sg13g2_decap_8 FILLER_74_1442 ();
 sg13g2_decap_8 FILLER_74_1459 ();
 sg13g2_decap_8 FILLER_74_1466 ();
 sg13g2_decap_8 FILLER_74_1473 ();
 sg13g2_decap_8 FILLER_74_1480 ();
 sg13g2_decap_8 FILLER_74_1487 ();
 sg13g2_decap_8 FILLER_74_1494 ();
 sg13g2_decap_8 FILLER_74_1501 ();
 sg13g2_decap_8 FILLER_74_1508 ();
 sg13g2_decap_8 FILLER_74_1515 ();
 sg13g2_decap_8 FILLER_74_1522 ();
 sg13g2_decap_8 FILLER_74_1529 ();
 sg13g2_decap_8 FILLER_74_1536 ();
 sg13g2_decap_8 FILLER_74_1543 ();
 sg13g2_decap_8 FILLER_74_1550 ();
 sg13g2_decap_8 FILLER_74_1557 ();
 sg13g2_decap_8 FILLER_74_1564 ();
 sg13g2_decap_8 FILLER_74_1571 ();
 sg13g2_decap_8 FILLER_74_1578 ();
 sg13g2_decap_8 FILLER_74_1585 ();
 sg13g2_decap_4 FILLER_74_1592 ();
 sg13g2_fill_2 FILLER_74_1618 ();
 sg13g2_decap_8 FILLER_74_1634 ();
 sg13g2_decap_8 FILLER_74_1641 ();
 sg13g2_decap_8 FILLER_74_1648 ();
 sg13g2_fill_2 FILLER_74_1655 ();
 sg13g2_fill_1 FILLER_74_1657 ();
 sg13g2_decap_8 FILLER_74_1684 ();
 sg13g2_decap_8 FILLER_74_1691 ();
 sg13g2_decap_8 FILLER_74_1698 ();
 sg13g2_decap_8 FILLER_74_1705 ();
 sg13g2_fill_2 FILLER_74_1712 ();
 sg13g2_fill_1 FILLER_74_1743 ();
 sg13g2_decap_8 FILLER_74_1754 ();
 sg13g2_decap_8 FILLER_74_1761 ();
 sg13g2_decap_8 FILLER_74_1774 ();
 sg13g2_fill_2 FILLER_74_1781 ();
 sg13g2_decap_8 FILLER_74_1809 ();
 sg13g2_decap_8 FILLER_74_1816 ();
 sg13g2_decap_8 FILLER_74_1823 ();
 sg13g2_decap_4 FILLER_74_1830 ();
 sg13g2_fill_1 FILLER_74_1834 ();
 sg13g2_decap_4 FILLER_74_1839 ();
 sg13g2_decap_8 FILLER_74_1847 ();
 sg13g2_decap_8 FILLER_74_1854 ();
 sg13g2_decap_8 FILLER_74_1861 ();
 sg13g2_decap_8 FILLER_74_1868 ();
 sg13g2_decap_8 FILLER_74_1875 ();
 sg13g2_decap_8 FILLER_74_1882 ();
 sg13g2_decap_8 FILLER_74_1889 ();
 sg13g2_decap_8 FILLER_74_1896 ();
 sg13g2_fill_2 FILLER_74_1903 ();
 sg13g2_decap_8 FILLER_74_1910 ();
 sg13g2_decap_8 FILLER_74_1917 ();
 sg13g2_fill_2 FILLER_74_1924 ();
 sg13g2_fill_1 FILLER_74_1926 ();
 sg13g2_decap_8 FILLER_74_1932 ();
 sg13g2_decap_8 FILLER_74_1939 ();
 sg13g2_decap_8 FILLER_74_1946 ();
 sg13g2_decap_8 FILLER_74_1953 ();
 sg13g2_decap_8 FILLER_74_1960 ();
 sg13g2_decap_8 FILLER_74_1967 ();
 sg13g2_decap_8 FILLER_74_1974 ();
 sg13g2_decap_8 FILLER_74_1981 ();
 sg13g2_decap_8 FILLER_74_1988 ();
 sg13g2_decap_8 FILLER_74_1995 ();
 sg13g2_decap_8 FILLER_74_2002 ();
 sg13g2_decap_8 FILLER_74_2009 ();
 sg13g2_decap_8 FILLER_74_2016 ();
 sg13g2_decap_8 FILLER_74_2023 ();
 sg13g2_decap_8 FILLER_74_2030 ();
 sg13g2_decap_8 FILLER_74_2037 ();
 sg13g2_decap_8 FILLER_74_2044 ();
 sg13g2_fill_1 FILLER_74_2051 ();
 sg13g2_decap_4 FILLER_74_2067 ();
 sg13g2_fill_1 FILLER_74_2071 ();
 sg13g2_decap_8 FILLER_74_2100 ();
 sg13g2_decap_8 FILLER_74_2107 ();
 sg13g2_decap_8 FILLER_74_2114 ();
 sg13g2_decap_8 FILLER_74_2121 ();
 sg13g2_decap_8 FILLER_74_2128 ();
 sg13g2_decap_8 FILLER_74_2135 ();
 sg13g2_decap_4 FILLER_74_2142 ();
 sg13g2_fill_1 FILLER_74_2146 ();
 sg13g2_decap_8 FILLER_74_2172 ();
 sg13g2_decap_8 FILLER_74_2179 ();
 sg13g2_decap_8 FILLER_74_2186 ();
 sg13g2_fill_2 FILLER_74_2193 ();
 sg13g2_fill_2 FILLER_74_2230 ();
 sg13g2_decap_8 FILLER_74_2258 ();
 sg13g2_decap_8 FILLER_74_2265 ();
 sg13g2_decap_8 FILLER_74_2272 ();
 sg13g2_decap_8 FILLER_74_2279 ();
 sg13g2_fill_2 FILLER_74_2286 ();
 sg13g2_fill_1 FILLER_74_2288 ();
 sg13g2_decap_8 FILLER_74_2300 ();
 sg13g2_decap_8 FILLER_74_2315 ();
 sg13g2_decap_8 FILLER_74_2322 ();
 sg13g2_decap_8 FILLER_74_2329 ();
 sg13g2_decap_4 FILLER_74_2336 ();
 sg13g2_fill_1 FILLER_74_2340 ();
 sg13g2_decap_8 FILLER_74_2356 ();
 sg13g2_decap_8 FILLER_74_2363 ();
 sg13g2_decap_4 FILLER_74_2370 ();
 sg13g2_fill_2 FILLER_74_2374 ();
 sg13g2_decap_8 FILLER_74_2381 ();
 sg13g2_decap_8 FILLER_74_2388 ();
 sg13g2_fill_2 FILLER_74_2395 ();
 sg13g2_fill_2 FILLER_74_2407 ();
 sg13g2_decap_8 FILLER_74_2435 ();
 sg13g2_decap_8 FILLER_74_2442 ();
 sg13g2_decap_8 FILLER_74_2449 ();
 sg13g2_decap_8 FILLER_74_2456 ();
 sg13g2_fill_1 FILLER_74_2463 ();
 sg13g2_decap_4 FILLER_74_2469 ();
 sg13g2_fill_1 FILLER_74_2473 ();
 sg13g2_decap_8 FILLER_74_2484 ();
 sg13g2_decap_8 FILLER_74_2491 ();
 sg13g2_decap_8 FILLER_74_2498 ();
 sg13g2_decap_8 FILLER_74_2505 ();
 sg13g2_decap_8 FILLER_74_2512 ();
 sg13g2_fill_2 FILLER_74_2519 ();
 sg13g2_decap_8 FILLER_74_2531 ();
 sg13g2_decap_8 FILLER_74_2538 ();
 sg13g2_decap_8 FILLER_74_2545 ();
 sg13g2_fill_2 FILLER_74_2552 ();
 sg13g2_fill_1 FILLER_74_2554 ();
 sg13g2_decap_8 FILLER_74_2591 ();
 sg13g2_decap_4 FILLER_74_2598 ();
 sg13g2_fill_2 FILLER_74_2602 ();
 sg13g2_decap_8 FILLER_74_2618 ();
 sg13g2_decap_8 FILLER_74_2625 ();
 sg13g2_decap_8 FILLER_74_2632 ();
 sg13g2_decap_8 FILLER_74_2639 ();
 sg13g2_decap_8 FILLER_74_2646 ();
 sg13g2_decap_4 FILLER_74_2653 ();
 sg13g2_fill_1 FILLER_74_2657 ();
 sg13g2_decap_4 FILLER_74_2663 ();
 sg13g2_decap_8 FILLER_74_2675 ();
 sg13g2_decap_8 FILLER_74_2682 ();
 sg13g2_decap_8 FILLER_74_2689 ();
 sg13g2_decap_8 FILLER_74_2696 ();
 sg13g2_decap_8 FILLER_74_2703 ();
 sg13g2_decap_8 FILLER_74_2710 ();
 sg13g2_decap_8 FILLER_74_2717 ();
 sg13g2_decap_8 FILLER_74_2724 ();
 sg13g2_decap_8 FILLER_74_2731 ();
 sg13g2_decap_8 FILLER_74_2738 ();
 sg13g2_decap_8 FILLER_74_2745 ();
 sg13g2_decap_8 FILLER_74_2752 ();
 sg13g2_decap_8 FILLER_74_2759 ();
 sg13g2_decap_8 FILLER_74_2766 ();
 sg13g2_decap_8 FILLER_74_2773 ();
 sg13g2_decap_8 FILLER_74_2780 ();
 sg13g2_decap_8 FILLER_74_2787 ();
 sg13g2_decap_8 FILLER_74_2794 ();
 sg13g2_decap_8 FILLER_74_2801 ();
 sg13g2_fill_2 FILLER_74_2808 ();
 sg13g2_decap_8 FILLER_74_2815 ();
 sg13g2_decap_8 FILLER_74_2822 ();
 sg13g2_decap_8 FILLER_74_2829 ();
 sg13g2_decap_8 FILLER_74_2836 ();
 sg13g2_decap_8 FILLER_74_2843 ();
 sg13g2_decap_8 FILLER_74_2850 ();
 sg13g2_fill_1 FILLER_74_2857 ();
 sg13g2_decap_8 FILLER_74_2861 ();
 sg13g2_decap_4 FILLER_74_2868 ();
 sg13g2_fill_2 FILLER_74_2872 ();
 sg13g2_decap_8 FILLER_74_2883 ();
 sg13g2_decap_8 FILLER_74_2890 ();
 sg13g2_decap_8 FILLER_74_2897 ();
 sg13g2_fill_2 FILLER_74_2904 ();
 sg13g2_decap_8 FILLER_74_2932 ();
 sg13g2_decap_8 FILLER_74_2939 ();
 sg13g2_decap_4 FILLER_74_2946 ();
 sg13g2_fill_2 FILLER_74_2950 ();
 sg13g2_fill_2 FILLER_74_2957 ();
 sg13g2_decap_8 FILLER_74_2969 ();
 sg13g2_decap_8 FILLER_74_2976 ();
 sg13g2_decap_8 FILLER_74_2983 ();
 sg13g2_decap_8 FILLER_74_2990 ();
 sg13g2_decap_8 FILLER_74_2997 ();
 sg13g2_decap_8 FILLER_74_3004 ();
 sg13g2_decap_4 FILLER_74_3011 ();
 sg13g2_decap_8 FILLER_74_3020 ();
 sg13g2_fill_2 FILLER_74_3027 ();
 sg13g2_fill_1 FILLER_74_3029 ();
 sg13g2_decap_8 FILLER_74_3056 ();
 sg13g2_decap_8 FILLER_74_3063 ();
 sg13g2_decap_4 FILLER_74_3070 ();
 sg13g2_fill_2 FILLER_74_3074 ();
 sg13g2_fill_2 FILLER_74_3102 ();
 sg13g2_decap_8 FILLER_74_3109 ();
 sg13g2_decap_8 FILLER_74_3116 ();
 sg13g2_fill_2 FILLER_74_3123 ();
 sg13g2_fill_1 FILLER_74_3125 ();
 sg13g2_decap_8 FILLER_74_3135 ();
 sg13g2_fill_1 FILLER_74_3142 ();
 sg13g2_decap_4 FILLER_74_3161 ();
 sg13g2_fill_1 FILLER_74_3165 ();
 sg13g2_decap_8 FILLER_74_3174 ();
 sg13g2_decap_8 FILLER_74_3186 ();
 sg13g2_decap_8 FILLER_74_3193 ();
 sg13g2_decap_8 FILLER_74_3200 ();
 sg13g2_fill_2 FILLER_74_3207 ();
 sg13g2_fill_1 FILLER_74_3209 ();
 sg13g2_decap_8 FILLER_74_3219 ();
 sg13g2_decap_8 FILLER_74_3226 ();
 sg13g2_decap_8 FILLER_74_3233 ();
 sg13g2_decap_8 FILLER_74_3240 ();
 sg13g2_decap_8 FILLER_74_3247 ();
 sg13g2_decap_8 FILLER_74_3254 ();
 sg13g2_decap_8 FILLER_74_3261 ();
 sg13g2_fill_2 FILLER_74_3268 ();
 sg13g2_decap_8 FILLER_74_3285 ();
 sg13g2_decap_8 FILLER_74_3292 ();
 sg13g2_decap_8 FILLER_74_3299 ();
 sg13g2_decap_8 FILLER_74_3306 ();
 sg13g2_decap_8 FILLER_74_3313 ();
 sg13g2_fill_2 FILLER_74_3320 ();
 sg13g2_fill_1 FILLER_74_3348 ();
 sg13g2_decap_8 FILLER_74_3380 ();
 sg13g2_decap_8 FILLER_74_3387 ();
 sg13g2_fill_2 FILLER_74_3394 ();
 sg13g2_decap_8 FILLER_74_3422 ();
 sg13g2_decap_8 FILLER_74_3432 ();
 sg13g2_decap_8 FILLER_74_3439 ();
 sg13g2_decap_8 FILLER_74_3446 ();
 sg13g2_decap_8 FILLER_74_3453 ();
 sg13g2_decap_8 FILLER_74_3460 ();
 sg13g2_decap_8 FILLER_74_3467 ();
 sg13g2_decap_8 FILLER_74_3474 ();
 sg13g2_decap_8 FILLER_74_3481 ();
 sg13g2_decap_8 FILLER_74_3488 ();
 sg13g2_decap_8 FILLER_74_3495 ();
 sg13g2_decap_8 FILLER_74_3502 ();
 sg13g2_decap_8 FILLER_74_3509 ();
 sg13g2_decap_8 FILLER_74_3516 ();
 sg13g2_decap_8 FILLER_74_3523 ();
 sg13g2_decap_8 FILLER_74_3530 ();
 sg13g2_decap_8 FILLER_74_3537 ();
 sg13g2_decap_8 FILLER_74_3544 ();
 sg13g2_decap_8 FILLER_74_3551 ();
 sg13g2_decap_8 FILLER_74_3558 ();
 sg13g2_decap_8 FILLER_74_3565 ();
 sg13g2_decap_8 FILLER_74_3572 ();
 sg13g2_fill_1 FILLER_74_3579 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_fill_2 FILLER_75_14 ();
 sg13g2_fill_1 FILLER_75_16 ();
 sg13g2_decap_8 FILLER_75_43 ();
 sg13g2_decap_8 FILLER_75_50 ();
 sg13g2_decap_8 FILLER_75_57 ();
 sg13g2_decap_4 FILLER_75_64 ();
 sg13g2_fill_1 FILLER_75_94 ();
 sg13g2_fill_2 FILLER_75_126 ();
 sg13g2_decap_8 FILLER_75_137 ();
 sg13g2_decap_8 FILLER_75_144 ();
 sg13g2_decap_4 FILLER_75_151 ();
 sg13g2_fill_2 FILLER_75_155 ();
 sg13g2_fill_1 FILLER_75_166 ();
 sg13g2_decap_8 FILLER_75_172 ();
 sg13g2_decap_8 FILLER_75_179 ();
 sg13g2_decap_8 FILLER_75_186 ();
 sg13g2_decap_8 FILLER_75_193 ();
 sg13g2_decap_8 FILLER_75_240 ();
 sg13g2_decap_8 FILLER_75_247 ();
 sg13g2_decap_4 FILLER_75_254 ();
 sg13g2_fill_2 FILLER_75_258 ();
 sg13g2_decap_8 FILLER_75_265 ();
 sg13g2_fill_1 FILLER_75_272 ();
 sg13g2_decap_8 FILLER_75_285 ();
 sg13g2_decap_8 FILLER_75_292 ();
 sg13g2_decap_4 FILLER_75_299 ();
 sg13g2_decap_8 FILLER_75_308 ();
 sg13g2_decap_8 FILLER_75_315 ();
 sg13g2_decap_8 FILLER_75_322 ();
 sg13g2_decap_4 FILLER_75_329 ();
 sg13g2_fill_1 FILLER_75_333 ();
 sg13g2_decap_8 FILLER_75_338 ();
 sg13g2_decap_8 FILLER_75_345 ();
 sg13g2_decap_8 FILLER_75_352 ();
 sg13g2_fill_2 FILLER_75_359 ();
 sg13g2_fill_1 FILLER_75_361 ();
 sg13g2_decap_4 FILLER_75_371 ();
 sg13g2_decap_8 FILLER_75_383 ();
 sg13g2_decap_8 FILLER_75_390 ();
 sg13g2_decap_4 FILLER_75_397 ();
 sg13g2_fill_1 FILLER_75_401 ();
 sg13g2_decap_8 FILLER_75_407 ();
 sg13g2_decap_8 FILLER_75_414 ();
 sg13g2_decap_8 FILLER_75_421 ();
 sg13g2_decap_8 FILLER_75_428 ();
 sg13g2_decap_8 FILLER_75_435 ();
 sg13g2_fill_2 FILLER_75_442 ();
 sg13g2_decap_8 FILLER_75_454 ();
 sg13g2_decap_8 FILLER_75_461 ();
 sg13g2_fill_2 FILLER_75_468 ();
 sg13g2_fill_1 FILLER_75_475 ();
 sg13g2_fill_2 FILLER_75_480 ();
 sg13g2_decap_8 FILLER_75_486 ();
 sg13g2_decap_8 FILLER_75_493 ();
 sg13g2_decap_8 FILLER_75_500 ();
 sg13g2_decap_8 FILLER_75_507 ();
 sg13g2_decap_8 FILLER_75_514 ();
 sg13g2_decap_8 FILLER_75_521 ();
 sg13g2_decap_8 FILLER_75_528 ();
 sg13g2_decap_8 FILLER_75_535 ();
 sg13g2_decap_8 FILLER_75_542 ();
 sg13g2_decap_8 FILLER_75_549 ();
 sg13g2_decap_8 FILLER_75_556 ();
 sg13g2_decap_8 FILLER_75_563 ();
 sg13g2_decap_8 FILLER_75_570 ();
 sg13g2_decap_8 FILLER_75_577 ();
 sg13g2_decap_8 FILLER_75_584 ();
 sg13g2_decap_4 FILLER_75_591 ();
 sg13g2_decap_8 FILLER_75_600 ();
 sg13g2_decap_8 FILLER_75_610 ();
 sg13g2_decap_8 FILLER_75_617 ();
 sg13g2_decap_8 FILLER_75_624 ();
 sg13g2_decap_8 FILLER_75_639 ();
 sg13g2_decap_4 FILLER_75_646 ();
 sg13g2_decap_8 FILLER_75_664 ();
 sg13g2_decap_8 FILLER_75_671 ();
 sg13g2_decap_8 FILLER_75_678 ();
 sg13g2_decap_8 FILLER_75_685 ();
 sg13g2_fill_1 FILLER_75_692 ();
 sg13g2_fill_2 FILLER_75_705 ();
 sg13g2_fill_1 FILLER_75_707 ();
 sg13g2_fill_2 FILLER_75_713 ();
 sg13g2_fill_1 FILLER_75_715 ();
 sg13g2_decap_8 FILLER_75_721 ();
 sg13g2_decap_4 FILLER_75_728 ();
 sg13g2_fill_2 FILLER_75_732 ();
 sg13g2_decap_8 FILLER_75_737 ();
 sg13g2_fill_2 FILLER_75_744 ();
 sg13g2_fill_1 FILLER_75_746 ();
 sg13g2_decap_8 FILLER_75_755 ();
 sg13g2_decap_8 FILLER_75_762 ();
 sg13g2_decap_8 FILLER_75_769 ();
 sg13g2_decap_8 FILLER_75_776 ();
 sg13g2_decap_8 FILLER_75_783 ();
 sg13g2_decap_8 FILLER_75_790 ();
 sg13g2_decap_8 FILLER_75_797 ();
 sg13g2_decap_8 FILLER_75_804 ();
 sg13g2_decap_8 FILLER_75_811 ();
 sg13g2_decap_8 FILLER_75_818 ();
 sg13g2_decap_8 FILLER_75_825 ();
 sg13g2_decap_8 FILLER_75_832 ();
 sg13g2_decap_8 FILLER_75_839 ();
 sg13g2_decap_8 FILLER_75_846 ();
 sg13g2_decap_8 FILLER_75_853 ();
 sg13g2_decap_8 FILLER_75_860 ();
 sg13g2_decap_8 FILLER_75_867 ();
 sg13g2_decap_8 FILLER_75_874 ();
 sg13g2_decap_8 FILLER_75_881 ();
 sg13g2_decap_8 FILLER_75_888 ();
 sg13g2_decap_8 FILLER_75_895 ();
 sg13g2_decap_8 FILLER_75_902 ();
 sg13g2_decap_8 FILLER_75_909 ();
 sg13g2_decap_8 FILLER_75_916 ();
 sg13g2_decap_4 FILLER_75_923 ();
 sg13g2_fill_1 FILLER_75_927 ();
 sg13g2_decap_8 FILLER_75_933 ();
 sg13g2_decap_8 FILLER_75_940 ();
 sg13g2_decap_8 FILLER_75_947 ();
 sg13g2_decap_8 FILLER_75_954 ();
 sg13g2_decap_8 FILLER_75_961 ();
 sg13g2_fill_1 FILLER_75_968 ();
 sg13g2_decap_8 FILLER_75_972 ();
 sg13g2_decap_4 FILLER_75_979 ();
 sg13g2_fill_2 FILLER_75_983 ();
 sg13g2_decap_8 FILLER_75_990 ();
 sg13g2_fill_2 FILLER_75_997 ();
 sg13g2_fill_1 FILLER_75_1004 ();
 sg13g2_decap_4 FILLER_75_1012 ();
 sg13g2_fill_1 FILLER_75_1016 ();
 sg13g2_decap_8 FILLER_75_1024 ();
 sg13g2_decap_8 FILLER_75_1031 ();
 sg13g2_decap_8 FILLER_75_1038 ();
 sg13g2_decap_8 FILLER_75_1045 ();
 sg13g2_decap_8 FILLER_75_1052 ();
 sg13g2_decap_4 FILLER_75_1059 ();
 sg13g2_decap_8 FILLER_75_1067 ();
 sg13g2_decap_8 FILLER_75_1074 ();
 sg13g2_decap_8 FILLER_75_1081 ();
 sg13g2_decap_8 FILLER_75_1088 ();
 sg13g2_decap_8 FILLER_75_1095 ();
 sg13g2_decap_4 FILLER_75_1102 ();
 sg13g2_fill_2 FILLER_75_1124 ();
 sg13g2_decap_8 FILLER_75_1140 ();
 sg13g2_decap_8 FILLER_75_1147 ();
 sg13g2_decap_8 FILLER_75_1154 ();
 sg13g2_decap_8 FILLER_75_1161 ();
 sg13g2_decap_4 FILLER_75_1168 ();
 sg13g2_fill_2 FILLER_75_1172 ();
 sg13g2_decap_8 FILLER_75_1178 ();
 sg13g2_fill_2 FILLER_75_1185 ();
 sg13g2_fill_1 FILLER_75_1187 ();
 sg13g2_decap_8 FILLER_75_1192 ();
 sg13g2_decap_8 FILLER_75_1199 ();
 sg13g2_decap_8 FILLER_75_1206 ();
 sg13g2_decap_8 FILLER_75_1213 ();
 sg13g2_decap_8 FILLER_75_1220 ();
 sg13g2_fill_1 FILLER_75_1227 ();
 sg13g2_decap_8 FILLER_75_1233 ();
 sg13g2_decap_8 FILLER_75_1240 ();
 sg13g2_decap_8 FILLER_75_1247 ();
 sg13g2_decap_8 FILLER_75_1254 ();
 sg13g2_fill_1 FILLER_75_1261 ();
 sg13g2_decap_8 FILLER_75_1270 ();
 sg13g2_fill_1 FILLER_75_1277 ();
 sg13g2_fill_1 FILLER_75_1291 ();
 sg13g2_decap_8 FILLER_75_1300 ();
 sg13g2_decap_8 FILLER_75_1307 ();
 sg13g2_fill_2 FILLER_75_1314 ();
 sg13g2_fill_1 FILLER_75_1316 ();
 sg13g2_decap_8 FILLER_75_1332 ();
 sg13g2_decap_8 FILLER_75_1339 ();
 sg13g2_fill_2 FILLER_75_1346 ();
 sg13g2_fill_1 FILLER_75_1348 ();
 sg13g2_fill_2 FILLER_75_1354 ();
 sg13g2_fill_1 FILLER_75_1356 ();
 sg13g2_fill_1 FILLER_75_1360 ();
 sg13g2_fill_1 FILLER_75_1373 ();
 sg13g2_fill_1 FILLER_75_1405 ();
 sg13g2_decap_8 FILLER_75_1418 ();
 sg13g2_decap_8 FILLER_75_1425 ();
 sg13g2_decap_8 FILLER_75_1432 ();
 sg13g2_decap_4 FILLER_75_1439 ();
 sg13g2_fill_2 FILLER_75_1443 ();
 sg13g2_decap_8 FILLER_75_1481 ();
 sg13g2_decap_8 FILLER_75_1488 ();
 sg13g2_decap_8 FILLER_75_1495 ();
 sg13g2_decap_8 FILLER_75_1502 ();
 sg13g2_decap_4 FILLER_75_1509 ();
 sg13g2_decap_8 FILLER_75_1523 ();
 sg13g2_fill_2 FILLER_75_1530 ();
 sg13g2_fill_1 FILLER_75_1532 ();
 sg13g2_decap_8 FILLER_75_1543 ();
 sg13g2_decap_8 FILLER_75_1550 ();
 sg13g2_decap_8 FILLER_75_1557 ();
 sg13g2_decap_8 FILLER_75_1564 ();
 sg13g2_decap_8 FILLER_75_1571 ();
 sg13g2_decap_8 FILLER_75_1578 ();
 sg13g2_decap_8 FILLER_75_1585 ();
 sg13g2_decap_4 FILLER_75_1592 ();
 sg13g2_decap_8 FILLER_75_1622 ();
 sg13g2_decap_8 FILLER_75_1629 ();
 sg13g2_decap_8 FILLER_75_1636 ();
 sg13g2_decap_8 FILLER_75_1643 ();
 sg13g2_decap_8 FILLER_75_1650 ();
 sg13g2_decap_8 FILLER_75_1657 ();
 sg13g2_decap_8 FILLER_75_1664 ();
 sg13g2_decap_8 FILLER_75_1671 ();
 sg13g2_decap_8 FILLER_75_1678 ();
 sg13g2_decap_8 FILLER_75_1685 ();
 sg13g2_decap_8 FILLER_75_1692 ();
 sg13g2_decap_8 FILLER_75_1699 ();
 sg13g2_decap_8 FILLER_75_1721 ();
 sg13g2_decap_8 FILLER_75_1728 ();
 sg13g2_decap_8 FILLER_75_1735 ();
 sg13g2_decap_8 FILLER_75_1742 ();
 sg13g2_decap_8 FILLER_75_1749 ();
 sg13g2_decap_8 FILLER_75_1756 ();
 sg13g2_decap_8 FILLER_75_1763 ();
 sg13g2_decap_4 FILLER_75_1770 ();
 sg13g2_decap_8 FILLER_75_1780 ();
 sg13g2_decap_8 FILLER_75_1787 ();
 sg13g2_decap_8 FILLER_75_1794 ();
 sg13g2_decap_8 FILLER_75_1801 ();
 sg13g2_decap_8 FILLER_75_1808 ();
 sg13g2_decap_8 FILLER_75_1815 ();
 sg13g2_decap_8 FILLER_75_1822 ();
 sg13g2_fill_2 FILLER_75_1829 ();
 sg13g2_fill_1 FILLER_75_1831 ();
 sg13g2_decap_8 FILLER_75_1849 ();
 sg13g2_decap_8 FILLER_75_1856 ();
 sg13g2_decap_8 FILLER_75_1863 ();
 sg13g2_decap_8 FILLER_75_1870 ();
 sg13g2_decap_8 FILLER_75_1877 ();
 sg13g2_decap_8 FILLER_75_1884 ();
 sg13g2_decap_8 FILLER_75_1891 ();
 sg13g2_decap_8 FILLER_75_1898 ();
 sg13g2_decap_8 FILLER_75_1905 ();
 sg13g2_decap_8 FILLER_75_1912 ();
 sg13g2_decap_8 FILLER_75_1919 ();
 sg13g2_decap_8 FILLER_75_1926 ();
 sg13g2_decap_8 FILLER_75_1933 ();
 sg13g2_decap_8 FILLER_75_1940 ();
 sg13g2_decap_8 FILLER_75_1947 ();
 sg13g2_decap_8 FILLER_75_1954 ();
 sg13g2_decap_8 FILLER_75_1961 ();
 sg13g2_fill_1 FILLER_75_1968 ();
 sg13g2_decap_8 FILLER_75_1979 ();
 sg13g2_decap_8 FILLER_75_1986 ();
 sg13g2_decap_8 FILLER_75_1993 ();
 sg13g2_decap_8 FILLER_75_2000 ();
 sg13g2_decap_8 FILLER_75_2007 ();
 sg13g2_decap_8 FILLER_75_2014 ();
 sg13g2_decap_8 FILLER_75_2021 ();
 sg13g2_decap_8 FILLER_75_2028 ();
 sg13g2_decap_8 FILLER_75_2035 ();
 sg13g2_decap_4 FILLER_75_2042 ();
 sg13g2_fill_1 FILLER_75_2046 ();
 sg13g2_decap_8 FILLER_75_2052 ();
 sg13g2_decap_8 FILLER_75_2067 ();
 sg13g2_decap_8 FILLER_75_2074 ();
 sg13g2_decap_8 FILLER_75_2081 ();
 sg13g2_decap_8 FILLER_75_2088 ();
 sg13g2_decap_8 FILLER_75_2095 ();
 sg13g2_decap_8 FILLER_75_2102 ();
 sg13g2_decap_8 FILLER_75_2109 ();
 sg13g2_decap_8 FILLER_75_2116 ();
 sg13g2_decap_8 FILLER_75_2123 ();
 sg13g2_decap_8 FILLER_75_2130 ();
 sg13g2_decap_8 FILLER_75_2137 ();
 sg13g2_decap_4 FILLER_75_2144 ();
 sg13g2_decap_8 FILLER_75_2165 ();
 sg13g2_decap_8 FILLER_75_2172 ();
 sg13g2_decap_8 FILLER_75_2179 ();
 sg13g2_decap_8 FILLER_75_2186 ();
 sg13g2_decap_8 FILLER_75_2193 ();
 sg13g2_decap_8 FILLER_75_2200 ();
 sg13g2_decap_8 FILLER_75_2207 ();
 sg13g2_decap_8 FILLER_75_2214 ();
 sg13g2_decap_8 FILLER_75_2234 ();
 sg13g2_fill_1 FILLER_75_2241 ();
 sg13g2_decap_8 FILLER_75_2272 ();
 sg13g2_decap_8 FILLER_75_2279 ();
 sg13g2_fill_2 FILLER_75_2286 ();
 sg13g2_fill_1 FILLER_75_2288 ();
 sg13g2_decap_8 FILLER_75_2315 ();
 sg13g2_decap_8 FILLER_75_2322 ();
 sg13g2_decap_8 FILLER_75_2329 ();
 sg13g2_decap_8 FILLER_75_2336 ();
 sg13g2_decap_4 FILLER_75_2343 ();
 sg13g2_decap_8 FILLER_75_2351 ();
 sg13g2_fill_1 FILLER_75_2358 ();
 sg13g2_decap_8 FILLER_75_2368 ();
 sg13g2_decap_8 FILLER_75_2375 ();
 sg13g2_decap_8 FILLER_75_2382 ();
 sg13g2_decap_4 FILLER_75_2389 ();
 sg13g2_fill_2 FILLER_75_2393 ();
 sg13g2_decap_8 FILLER_75_2404 ();
 sg13g2_decap_8 FILLER_75_2411 ();
 sg13g2_decap_8 FILLER_75_2418 ();
 sg13g2_decap_8 FILLER_75_2425 ();
 sg13g2_decap_8 FILLER_75_2432 ();
 sg13g2_fill_2 FILLER_75_2439 ();
 sg13g2_decap_8 FILLER_75_2446 ();
 sg13g2_decap_8 FILLER_75_2453 ();
 sg13g2_decap_4 FILLER_75_2460 ();
 sg13g2_decap_8 FILLER_75_2469 ();
 sg13g2_decap_8 FILLER_75_2476 ();
 sg13g2_decap_8 FILLER_75_2483 ();
 sg13g2_decap_8 FILLER_75_2490 ();
 sg13g2_decap_8 FILLER_75_2497 ();
 sg13g2_decap_8 FILLER_75_2504 ();
 sg13g2_fill_2 FILLER_75_2511 ();
 sg13g2_decap_8 FILLER_75_2549 ();
 sg13g2_fill_1 FILLER_75_2556 ();
 sg13g2_fill_1 FILLER_75_2574 ();
 sg13g2_decap_8 FILLER_75_2584 ();
 sg13g2_decap_8 FILLER_75_2591 ();
 sg13g2_decap_8 FILLER_75_2598 ();
 sg13g2_decap_4 FILLER_75_2605 ();
 sg13g2_decap_8 FILLER_75_2614 ();
 sg13g2_decap_8 FILLER_75_2621 ();
 sg13g2_decap_8 FILLER_75_2628 ();
 sg13g2_decap_8 FILLER_75_2635 ();
 sg13g2_decap_8 FILLER_75_2642 ();
 sg13g2_decap_8 FILLER_75_2649 ();
 sg13g2_decap_8 FILLER_75_2656 ();
 sg13g2_fill_1 FILLER_75_2663 ();
 sg13g2_decap_8 FILLER_75_2671 ();
 sg13g2_decap_4 FILLER_75_2678 ();
 sg13g2_fill_2 FILLER_75_2682 ();
 sg13g2_decap_8 FILLER_75_2701 ();
 sg13g2_decap_8 FILLER_75_2708 ();
 sg13g2_decap_8 FILLER_75_2715 ();
 sg13g2_decap_8 FILLER_75_2722 ();
 sg13g2_decap_8 FILLER_75_2729 ();
 sg13g2_decap_8 FILLER_75_2736 ();
 sg13g2_decap_8 FILLER_75_2743 ();
 sg13g2_decap_8 FILLER_75_2750 ();
 sg13g2_decap_8 FILLER_75_2757 ();
 sg13g2_decap_8 FILLER_75_2764 ();
 sg13g2_decap_8 FILLER_75_2771 ();
 sg13g2_decap_8 FILLER_75_2778 ();
 sg13g2_fill_2 FILLER_75_2795 ();
 sg13g2_fill_1 FILLER_75_2797 ();
 sg13g2_fill_2 FILLER_75_2824 ();
 sg13g2_decap_8 FILLER_75_2829 ();
 sg13g2_decap_8 FILLER_75_2836 ();
 sg13g2_decap_4 FILLER_75_2843 ();
 sg13g2_fill_1 FILLER_75_2847 ();
 sg13g2_decap_8 FILLER_75_2885 ();
 sg13g2_decap_8 FILLER_75_2892 ();
 sg13g2_decap_8 FILLER_75_2899 ();
 sg13g2_decap_8 FILLER_75_2906 ();
 sg13g2_decap_4 FILLER_75_2913 ();
 sg13g2_decap_8 FILLER_75_2926 ();
 sg13g2_decap_4 FILLER_75_2933 ();
 sg13g2_decap_8 FILLER_75_2942 ();
 sg13g2_decap_4 FILLER_75_2949 ();
 sg13g2_fill_2 FILLER_75_2953 ();
 sg13g2_fill_2 FILLER_75_2960 ();
 sg13g2_fill_1 FILLER_75_2962 ();
 sg13g2_decap_8 FILLER_75_2968 ();
 sg13g2_decap_8 FILLER_75_2975 ();
 sg13g2_decap_8 FILLER_75_2982 ();
 sg13g2_decap_8 FILLER_75_2989 ();
 sg13g2_decap_8 FILLER_75_2996 ();
 sg13g2_decap_8 FILLER_75_3003 ();
 sg13g2_fill_1 FILLER_75_3010 ();
 sg13g2_decap_8 FILLER_75_3015 ();
 sg13g2_decap_8 FILLER_75_3022 ();
 sg13g2_decap_8 FILLER_75_3029 ();
 sg13g2_decap_8 FILLER_75_3036 ();
 sg13g2_decap_8 FILLER_75_3043 ();
 sg13g2_decap_8 FILLER_75_3050 ();
 sg13g2_decap_8 FILLER_75_3057 ();
 sg13g2_decap_8 FILLER_75_3064 ();
 sg13g2_decap_8 FILLER_75_3071 ();
 sg13g2_decap_8 FILLER_75_3078 ();
 sg13g2_decap_8 FILLER_75_3085 ();
 sg13g2_decap_8 FILLER_75_3092 ();
 sg13g2_decap_8 FILLER_75_3099 ();
 sg13g2_decap_8 FILLER_75_3106 ();
 sg13g2_fill_2 FILLER_75_3113 ();
 sg13g2_fill_1 FILLER_75_3115 ();
 sg13g2_decap_8 FILLER_75_3121 ();
 sg13g2_decap_8 FILLER_75_3128 ();
 sg13g2_decap_4 FILLER_75_3135 ();
 sg13g2_fill_2 FILLER_75_3139 ();
 sg13g2_decap_8 FILLER_75_3145 ();
 sg13g2_decap_8 FILLER_75_3152 ();
 sg13g2_fill_1 FILLER_75_3159 ();
 sg13g2_decap_8 FILLER_75_3195 ();
 sg13g2_decap_8 FILLER_75_3202 ();
 sg13g2_decap_8 FILLER_75_3209 ();
 sg13g2_decap_4 FILLER_75_3216 ();
 sg13g2_fill_2 FILLER_75_3220 ();
 sg13g2_decap_8 FILLER_75_3232 ();
 sg13g2_decap_8 FILLER_75_3239 ();
 sg13g2_decap_8 FILLER_75_3246 ();
 sg13g2_decap_8 FILLER_75_3253 ();
 sg13g2_decap_4 FILLER_75_3260 ();
 sg13g2_fill_2 FILLER_75_3264 ();
 sg13g2_decap_4 FILLER_75_3271 ();
 sg13g2_decap_8 FILLER_75_3289 ();
 sg13g2_decap_4 FILLER_75_3296 ();
 sg13g2_fill_1 FILLER_75_3300 ();
 sg13g2_decap_8 FILLER_75_3306 ();
 sg13g2_decap_8 FILLER_75_3313 ();
 sg13g2_decap_8 FILLER_75_3320 ();
 sg13g2_decap_8 FILLER_75_3327 ();
 sg13g2_decap_8 FILLER_75_3334 ();
 sg13g2_decap_8 FILLER_75_3341 ();
 sg13g2_decap_8 FILLER_75_3348 ();
 sg13g2_decap_8 FILLER_75_3355 ();
 sg13g2_decap_8 FILLER_75_3362 ();
 sg13g2_decap_8 FILLER_75_3369 ();
 sg13g2_decap_8 FILLER_75_3376 ();
 sg13g2_decap_8 FILLER_75_3383 ();
 sg13g2_decap_8 FILLER_75_3390 ();
 sg13g2_decap_8 FILLER_75_3397 ();
 sg13g2_decap_8 FILLER_75_3404 ();
 sg13g2_decap_8 FILLER_75_3411 ();
 sg13g2_fill_2 FILLER_75_3418 ();
 sg13g2_fill_1 FILLER_75_3420 ();
 sg13g2_decap_8 FILLER_75_3437 ();
 sg13g2_decap_8 FILLER_75_3444 ();
 sg13g2_decap_8 FILLER_75_3451 ();
 sg13g2_decap_8 FILLER_75_3458 ();
 sg13g2_decap_8 FILLER_75_3465 ();
 sg13g2_decap_8 FILLER_75_3472 ();
 sg13g2_decap_8 FILLER_75_3479 ();
 sg13g2_decap_8 FILLER_75_3486 ();
 sg13g2_decap_8 FILLER_75_3493 ();
 sg13g2_decap_8 FILLER_75_3500 ();
 sg13g2_decap_8 FILLER_75_3507 ();
 sg13g2_decap_8 FILLER_75_3514 ();
 sg13g2_decap_8 FILLER_75_3521 ();
 sg13g2_decap_8 FILLER_75_3528 ();
 sg13g2_decap_8 FILLER_75_3535 ();
 sg13g2_decap_8 FILLER_75_3542 ();
 sg13g2_decap_8 FILLER_75_3549 ();
 sg13g2_decap_8 FILLER_75_3556 ();
 sg13g2_decap_8 FILLER_75_3563 ();
 sg13g2_decap_8 FILLER_75_3570 ();
 sg13g2_fill_2 FILLER_75_3577 ();
 sg13g2_fill_1 FILLER_75_3579 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_8 FILLER_76_21 ();
 sg13g2_decap_4 FILLER_76_28 ();
 sg13g2_fill_1 FILLER_76_32 ();
 sg13g2_decap_8 FILLER_76_42 ();
 sg13g2_decap_8 FILLER_76_49 ();
 sg13g2_decap_8 FILLER_76_56 ();
 sg13g2_decap_8 FILLER_76_63 ();
 sg13g2_fill_1 FILLER_76_70 ();
 sg13g2_decap_8 FILLER_76_80 ();
 sg13g2_decap_8 FILLER_76_87 ();
 sg13g2_decap_8 FILLER_76_94 ();
 sg13g2_decap_8 FILLER_76_101 ();
 sg13g2_decap_8 FILLER_76_108 ();
 sg13g2_decap_8 FILLER_76_115 ();
 sg13g2_decap_8 FILLER_76_122 ();
 sg13g2_decap_8 FILLER_76_129 ();
 sg13g2_decap_8 FILLER_76_136 ();
 sg13g2_decap_8 FILLER_76_143 ();
 sg13g2_fill_2 FILLER_76_150 ();
 sg13g2_decap_8 FILLER_76_183 ();
 sg13g2_decap_8 FILLER_76_190 ();
 sg13g2_decap_8 FILLER_76_197 ();
 sg13g2_fill_1 FILLER_76_204 ();
 sg13g2_fill_2 FILLER_76_214 ();
 sg13g2_decap_8 FILLER_76_226 ();
 sg13g2_decap_8 FILLER_76_233 ();
 sg13g2_decap_8 FILLER_76_240 ();
 sg13g2_decap_8 FILLER_76_247 ();
 sg13g2_fill_2 FILLER_76_254 ();
 sg13g2_fill_2 FILLER_76_270 ();
 sg13g2_fill_1 FILLER_76_277 ();
 sg13g2_fill_2 FILLER_76_287 ();
 sg13g2_fill_1 FILLER_76_289 ();
 sg13g2_decap_8 FILLER_76_304 ();
 sg13g2_decap_8 FILLER_76_311 ();
 sg13g2_decap_8 FILLER_76_318 ();
 sg13g2_decap_4 FILLER_76_325 ();
 sg13g2_decap_8 FILLER_76_341 ();
 sg13g2_decap_8 FILLER_76_348 ();
 sg13g2_decap_4 FILLER_76_355 ();
 sg13g2_fill_2 FILLER_76_359 ();
 sg13g2_decap_8 FILLER_76_379 ();
 sg13g2_decap_8 FILLER_76_386 ();
 sg13g2_decap_8 FILLER_76_393 ();
 sg13g2_decap_8 FILLER_76_400 ();
 sg13g2_fill_1 FILLER_76_407 ();
 sg13g2_decap_8 FILLER_76_413 ();
 sg13g2_decap_8 FILLER_76_420 ();
 sg13g2_decap_8 FILLER_76_427 ();
 sg13g2_decap_8 FILLER_76_434 ();
 sg13g2_decap_4 FILLER_76_441 ();
 sg13g2_fill_1 FILLER_76_445 ();
 sg13g2_decap_8 FILLER_76_459 ();
 sg13g2_fill_1 FILLER_76_466 ();
 sg13g2_fill_2 FILLER_76_474 ();
 sg13g2_decap_8 FILLER_76_490 ();
 sg13g2_decap_8 FILLER_76_497 ();
 sg13g2_decap_8 FILLER_76_504 ();
 sg13g2_decap_8 FILLER_76_511 ();
 sg13g2_decap_8 FILLER_76_518 ();
 sg13g2_decap_8 FILLER_76_525 ();
 sg13g2_decap_8 FILLER_76_532 ();
 sg13g2_decap_8 FILLER_76_539 ();
 sg13g2_decap_8 FILLER_76_546 ();
 sg13g2_decap_8 FILLER_76_553 ();
 sg13g2_decap_8 FILLER_76_560 ();
 sg13g2_decap_8 FILLER_76_567 ();
 sg13g2_decap_8 FILLER_76_574 ();
 sg13g2_decap_8 FILLER_76_581 ();
 sg13g2_fill_2 FILLER_76_588 ();
 sg13g2_decap_4 FILLER_76_598 ();
 sg13g2_fill_2 FILLER_76_602 ();
 sg13g2_decap_8 FILLER_76_616 ();
 sg13g2_decap_8 FILLER_76_623 ();
 sg13g2_decap_8 FILLER_76_630 ();
 sg13g2_decap_4 FILLER_76_637 ();
 sg13g2_fill_2 FILLER_76_641 ();
 sg13g2_decap_8 FILLER_76_673 ();
 sg13g2_decap_8 FILLER_76_680 ();
 sg13g2_decap_8 FILLER_76_687 ();
 sg13g2_fill_1 FILLER_76_694 ();
 sg13g2_fill_1 FILLER_76_708 ();
 sg13g2_decap_8 FILLER_76_719 ();
 sg13g2_decap_8 FILLER_76_726 ();
 sg13g2_decap_8 FILLER_76_733 ();
 sg13g2_decap_8 FILLER_76_752 ();
 sg13g2_fill_2 FILLER_76_759 ();
 sg13g2_fill_1 FILLER_76_761 ();
 sg13g2_decap_8 FILLER_76_771 ();
 sg13g2_decap_8 FILLER_76_778 ();
 sg13g2_decap_8 FILLER_76_785 ();
 sg13g2_decap_8 FILLER_76_792 ();
 sg13g2_decap_8 FILLER_76_799 ();
 sg13g2_decap_4 FILLER_76_806 ();
 sg13g2_fill_2 FILLER_76_810 ();
 sg13g2_decap_8 FILLER_76_817 ();
 sg13g2_decap_4 FILLER_76_824 ();
 sg13g2_fill_2 FILLER_76_828 ();
 sg13g2_decap_8 FILLER_76_847 ();
 sg13g2_decap_8 FILLER_76_854 ();
 sg13g2_decap_8 FILLER_76_861 ();
 sg13g2_decap_8 FILLER_76_868 ();
 sg13g2_decap_8 FILLER_76_875 ();
 sg13g2_decap_8 FILLER_76_882 ();
 sg13g2_decap_8 FILLER_76_889 ();
 sg13g2_decap_8 FILLER_76_896 ();
 sg13g2_decap_8 FILLER_76_903 ();
 sg13g2_decap_8 FILLER_76_910 ();
 sg13g2_decap_8 FILLER_76_917 ();
 sg13g2_fill_2 FILLER_76_947 ();
 sg13g2_decap_8 FILLER_76_953 ();
 sg13g2_decap_8 FILLER_76_960 ();
 sg13g2_decap_8 FILLER_76_967 ();
 sg13g2_decap_8 FILLER_76_974 ();
 sg13g2_decap_4 FILLER_76_981 ();
 sg13g2_fill_2 FILLER_76_985 ();
 sg13g2_decap_8 FILLER_76_1022 ();
 sg13g2_decap_8 FILLER_76_1029 ();
 sg13g2_decap_8 FILLER_76_1036 ();
 sg13g2_decap_8 FILLER_76_1043 ();
 sg13g2_decap_8 FILLER_76_1050 ();
 sg13g2_decap_8 FILLER_76_1057 ();
 sg13g2_decap_8 FILLER_76_1064 ();
 sg13g2_decap_8 FILLER_76_1071 ();
 sg13g2_fill_2 FILLER_76_1078 ();
 sg13g2_decap_8 FILLER_76_1093 ();
 sg13g2_decap_8 FILLER_76_1100 ();
 sg13g2_decap_8 FILLER_76_1107 ();
 sg13g2_fill_2 FILLER_76_1114 ();
 sg13g2_fill_1 FILLER_76_1116 ();
 sg13g2_fill_1 FILLER_76_1127 ();
 sg13g2_decap_8 FILLER_76_1141 ();
 sg13g2_decap_8 FILLER_76_1148 ();
 sg13g2_fill_1 FILLER_76_1155 ();
 sg13g2_decap_4 FILLER_76_1159 ();
 sg13g2_fill_1 FILLER_76_1163 ();
 sg13g2_fill_2 FILLER_76_1174 ();
 sg13g2_decap_8 FILLER_76_1191 ();
 sg13g2_decap_4 FILLER_76_1198 ();
 sg13g2_fill_1 FILLER_76_1202 ();
 sg13g2_decap_8 FILLER_76_1206 ();
 sg13g2_fill_2 FILLER_76_1221 ();
 sg13g2_fill_2 FILLER_76_1240 ();
 sg13g2_fill_1 FILLER_76_1242 ();
 sg13g2_decap_8 FILLER_76_1256 ();
 sg13g2_decap_8 FILLER_76_1263 ();
 sg13g2_decap_8 FILLER_76_1270 ();
 sg13g2_decap_8 FILLER_76_1277 ();
 sg13g2_decap_8 FILLER_76_1284 ();
 sg13g2_decap_4 FILLER_76_1291 ();
 sg13g2_fill_2 FILLER_76_1295 ();
 sg13g2_fill_1 FILLER_76_1306 ();
 sg13g2_fill_2 FILLER_76_1312 ();
 sg13g2_fill_1 FILLER_76_1314 ();
 sg13g2_decap_8 FILLER_76_1331 ();
 sg13g2_decap_4 FILLER_76_1344 ();
 sg13g2_decap_8 FILLER_76_1367 ();
 sg13g2_decap_8 FILLER_76_1374 ();
 sg13g2_fill_2 FILLER_76_1381 ();
 sg13g2_fill_1 FILLER_76_1383 ();
 sg13g2_decap_8 FILLER_76_1407 ();
 sg13g2_decap_8 FILLER_76_1414 ();
 sg13g2_decap_8 FILLER_76_1421 ();
 sg13g2_decap_8 FILLER_76_1428 ();
 sg13g2_decap_8 FILLER_76_1435 ();
 sg13g2_decap_8 FILLER_76_1442 ();
 sg13g2_fill_1 FILLER_76_1449 ();
 sg13g2_decap_4 FILLER_76_1456 ();
 sg13g2_decap_8 FILLER_76_1486 ();
 sg13g2_decap_4 FILLER_76_1493 ();
 sg13g2_decap_4 FILLER_76_1502 ();
 sg13g2_fill_2 FILLER_76_1542 ();
 sg13g2_fill_1 FILLER_76_1544 ();
 sg13g2_decap_8 FILLER_76_1584 ();
 sg13g2_decap_8 FILLER_76_1591 ();
 sg13g2_decap_8 FILLER_76_1598 ();
 sg13g2_decap_8 FILLER_76_1605 ();
 sg13g2_decap_8 FILLER_76_1620 ();
 sg13g2_decap_8 FILLER_76_1627 ();
 sg13g2_decap_8 FILLER_76_1634 ();
 sg13g2_decap_8 FILLER_76_1641 ();
 sg13g2_decap_8 FILLER_76_1648 ();
 sg13g2_decap_8 FILLER_76_1655 ();
 sg13g2_decap_8 FILLER_76_1662 ();
 sg13g2_decap_4 FILLER_76_1673 ();
 sg13g2_decap_4 FILLER_76_1681 ();
 sg13g2_decap_8 FILLER_76_1689 ();
 sg13g2_decap_8 FILLER_76_1696 ();
 sg13g2_decap_8 FILLER_76_1703 ();
 sg13g2_fill_2 FILLER_76_1710 ();
 sg13g2_fill_1 FILLER_76_1712 ();
 sg13g2_decap_8 FILLER_76_1719 ();
 sg13g2_decap_8 FILLER_76_1726 ();
 sg13g2_decap_8 FILLER_76_1733 ();
 sg13g2_decap_8 FILLER_76_1740 ();
 sg13g2_decap_8 FILLER_76_1747 ();
 sg13g2_decap_8 FILLER_76_1754 ();
 sg13g2_decap_8 FILLER_76_1761 ();
 sg13g2_decap_8 FILLER_76_1768 ();
 sg13g2_decap_8 FILLER_76_1775 ();
 sg13g2_fill_2 FILLER_76_1782 ();
 sg13g2_fill_1 FILLER_76_1784 ();
 sg13g2_decap_8 FILLER_76_1798 ();
 sg13g2_decap_8 FILLER_76_1805 ();
 sg13g2_decap_8 FILLER_76_1812 ();
 sg13g2_decap_8 FILLER_76_1819 ();
 sg13g2_decap_8 FILLER_76_1826 ();
 sg13g2_decap_8 FILLER_76_1841 ();
 sg13g2_decap_8 FILLER_76_1848 ();
 sg13g2_decap_8 FILLER_76_1855 ();
 sg13g2_decap_8 FILLER_76_1862 ();
 sg13g2_decap_8 FILLER_76_1869 ();
 sg13g2_decap_8 FILLER_76_1876 ();
 sg13g2_decap_8 FILLER_76_1883 ();
 sg13g2_fill_2 FILLER_76_1890 ();
 sg13g2_decap_8 FILLER_76_1906 ();
 sg13g2_decap_8 FILLER_76_1913 ();
 sg13g2_fill_1 FILLER_76_1920 ();
 sg13g2_decap_8 FILLER_76_1931 ();
 sg13g2_decap_8 FILLER_76_1938 ();
 sg13g2_decap_8 FILLER_76_1945 ();
 sg13g2_decap_8 FILLER_76_1952 ();
 sg13g2_decap_8 FILLER_76_1959 ();
 sg13g2_decap_8 FILLER_76_1966 ();
 sg13g2_decap_8 FILLER_76_1993 ();
 sg13g2_decap_8 FILLER_76_2000 ();
 sg13g2_decap_8 FILLER_76_2007 ();
 sg13g2_decap_8 FILLER_76_2014 ();
 sg13g2_decap_8 FILLER_76_2021 ();
 sg13g2_decap_8 FILLER_76_2028 ();
 sg13g2_fill_1 FILLER_76_2035 ();
 sg13g2_fill_2 FILLER_76_2044 ();
 sg13g2_fill_1 FILLER_76_2046 ();
 sg13g2_decap_8 FILLER_76_2064 ();
 sg13g2_decap_8 FILLER_76_2071 ();
 sg13g2_decap_8 FILLER_76_2078 ();
 sg13g2_fill_1 FILLER_76_2085 ();
 sg13g2_decap_8 FILLER_76_2094 ();
 sg13g2_decap_8 FILLER_76_2101 ();
 sg13g2_decap_8 FILLER_76_2108 ();
 sg13g2_decap_8 FILLER_76_2115 ();
 sg13g2_decap_8 FILLER_76_2122 ();
 sg13g2_decap_8 FILLER_76_2129 ();
 sg13g2_fill_2 FILLER_76_2136 ();
 sg13g2_decap_8 FILLER_76_2160 ();
 sg13g2_decap_8 FILLER_76_2167 ();
 sg13g2_decap_8 FILLER_76_2174 ();
 sg13g2_decap_8 FILLER_76_2181 ();
 sg13g2_decap_8 FILLER_76_2188 ();
 sg13g2_decap_8 FILLER_76_2195 ();
 sg13g2_decap_8 FILLER_76_2202 ();
 sg13g2_decap_8 FILLER_76_2209 ();
 sg13g2_fill_2 FILLER_76_2216 ();
 sg13g2_fill_1 FILLER_76_2218 ();
 sg13g2_decap_4 FILLER_76_2228 ();
 sg13g2_fill_2 FILLER_76_2232 ();
 sg13g2_decap_8 FILLER_76_2240 ();
 sg13g2_fill_1 FILLER_76_2247 ();
 sg13g2_fill_2 FILLER_76_2253 ();
 sg13g2_decap_8 FILLER_76_2268 ();
 sg13g2_decap_8 FILLER_76_2275 ();
 sg13g2_decap_8 FILLER_76_2282 ();
 sg13g2_decap_8 FILLER_76_2289 ();
 sg13g2_fill_2 FILLER_76_2296 ();
 sg13g2_fill_1 FILLER_76_2298 ();
 sg13g2_decap_8 FILLER_76_2318 ();
 sg13g2_decap_8 FILLER_76_2325 ();
 sg13g2_decap_8 FILLER_76_2332 ();
 sg13g2_decap_4 FILLER_76_2339 ();
 sg13g2_decap_8 FILLER_76_2369 ();
 sg13g2_decap_8 FILLER_76_2376 ();
 sg13g2_decap_8 FILLER_76_2383 ();
 sg13g2_decap_8 FILLER_76_2390 ();
 sg13g2_decap_8 FILLER_76_2397 ();
 sg13g2_fill_1 FILLER_76_2404 ();
 sg13g2_decap_8 FILLER_76_2431 ();
 sg13g2_decap_8 FILLER_76_2438 ();
 sg13g2_decap_4 FILLER_76_2445 ();
 sg13g2_fill_1 FILLER_76_2457 ();
 sg13g2_decap_8 FILLER_76_2498 ();
 sg13g2_decap_8 FILLER_76_2536 ();
 sg13g2_decap_8 FILLER_76_2543 ();
 sg13g2_decap_8 FILLER_76_2550 ();
 sg13g2_decap_8 FILLER_76_2557 ();
 sg13g2_decap_4 FILLER_76_2564 ();
 sg13g2_decap_8 FILLER_76_2573 ();
 sg13g2_decap_8 FILLER_76_2580 ();
 sg13g2_decap_8 FILLER_76_2587 ();
 sg13g2_decap_8 FILLER_76_2594 ();
 sg13g2_decap_4 FILLER_76_2601 ();
 sg13g2_fill_2 FILLER_76_2605 ();
 sg13g2_fill_2 FILLER_76_2631 ();
 sg13g2_fill_1 FILLER_76_2633 ();
 sg13g2_decap_8 FILLER_76_2647 ();
 sg13g2_decap_8 FILLER_76_2654 ();
 sg13g2_decap_4 FILLER_76_2661 ();
 sg13g2_fill_2 FILLER_76_2665 ();
 sg13g2_decap_8 FILLER_76_2670 ();
 sg13g2_fill_2 FILLER_76_2677 ();
 sg13g2_fill_1 FILLER_76_2679 ();
 sg13g2_decap_4 FILLER_76_2689 ();
 sg13g2_fill_2 FILLER_76_2693 ();
 sg13g2_decap_4 FILLER_76_2702 ();
 sg13g2_fill_1 FILLER_76_2706 ();
 sg13g2_fill_1 FILLER_76_2718 ();
 sg13g2_decap_4 FILLER_76_2727 ();
 sg13g2_fill_1 FILLER_76_2731 ();
 sg13g2_decap_8 FILLER_76_2743 ();
 sg13g2_decap_8 FILLER_76_2750 ();
 sg13g2_fill_2 FILLER_76_2757 ();
 sg13g2_decap_8 FILLER_76_2771 ();
 sg13g2_fill_2 FILLER_76_2778 ();
 sg13g2_fill_1 FILLER_76_2780 ();
 sg13g2_decap_8 FILLER_76_2786 ();
 sg13g2_decap_8 FILLER_76_2793 ();
 sg13g2_decap_8 FILLER_76_2800 ();
 sg13g2_fill_2 FILLER_76_2807 ();
 sg13g2_decap_8 FILLER_76_2830 ();
 sg13g2_decap_8 FILLER_76_2837 ();
 sg13g2_decap_8 FILLER_76_2844 ();
 sg13g2_decap_8 FILLER_76_2851 ();
 sg13g2_decap_8 FILLER_76_2858 ();
 sg13g2_decap_4 FILLER_76_2865 ();
 sg13g2_fill_1 FILLER_76_2869 ();
 sg13g2_decap_8 FILLER_76_2881 ();
 sg13g2_decap_8 FILLER_76_2888 ();
 sg13g2_decap_8 FILLER_76_2895 ();
 sg13g2_decap_8 FILLER_76_2902 ();
 sg13g2_decap_8 FILLER_76_2909 ();
 sg13g2_decap_8 FILLER_76_2916 ();
 sg13g2_decap_8 FILLER_76_2923 ();
 sg13g2_decap_8 FILLER_76_2930 ();
 sg13g2_decap_8 FILLER_76_2937 ();
 sg13g2_fill_1 FILLER_76_2944 ();
 sg13g2_decap_8 FILLER_76_2962 ();
 sg13g2_decap_8 FILLER_76_2969 ();
 sg13g2_decap_8 FILLER_76_2976 ();
 sg13g2_decap_4 FILLER_76_2983 ();
 sg13g2_fill_1 FILLER_76_2987 ();
 sg13g2_fill_1 FILLER_76_2993 ();
 sg13g2_decap_8 FILLER_76_3002 ();
 sg13g2_fill_2 FILLER_76_3009 ();
 sg13g2_decap_8 FILLER_76_3016 ();
 sg13g2_decap_8 FILLER_76_3023 ();
 sg13g2_fill_2 FILLER_76_3030 ();
 sg13g2_fill_1 FILLER_76_3032 ();
 sg13g2_decap_8 FILLER_76_3043 ();
 sg13g2_decap_8 FILLER_76_3050 ();
 sg13g2_decap_8 FILLER_76_3057 ();
 sg13g2_decap_8 FILLER_76_3064 ();
 sg13g2_decap_8 FILLER_76_3071 ();
 sg13g2_decap_8 FILLER_76_3078 ();
 sg13g2_decap_8 FILLER_76_3098 ();
 sg13g2_decap_8 FILLER_76_3105 ();
 sg13g2_decap_8 FILLER_76_3112 ();
 sg13g2_decap_8 FILLER_76_3119 ();
 sg13g2_fill_1 FILLER_76_3126 ();
 sg13g2_fill_1 FILLER_76_3146 ();
 sg13g2_decap_8 FILLER_76_3156 ();
 sg13g2_decap_8 FILLER_76_3163 ();
 sg13g2_decap_8 FILLER_76_3170 ();
 sg13g2_decap_4 FILLER_76_3177 ();
 sg13g2_fill_2 FILLER_76_3181 ();
 sg13g2_decap_8 FILLER_76_3188 ();
 sg13g2_fill_1 FILLER_76_3195 ();
 sg13g2_decap_8 FILLER_76_3199 ();
 sg13g2_decap_8 FILLER_76_3206 ();
 sg13g2_decap_8 FILLER_76_3213 ();
 sg13g2_fill_1 FILLER_76_3220 ();
 sg13g2_decap_8 FILLER_76_3247 ();
 sg13g2_decap_8 FILLER_76_3254 ();
 sg13g2_fill_2 FILLER_76_3261 ();
 sg13g2_decap_8 FILLER_76_3289 ();
 sg13g2_decap_8 FILLER_76_3296 ();
 sg13g2_decap_8 FILLER_76_3303 ();
 sg13g2_decap_8 FILLER_76_3310 ();
 sg13g2_decap_8 FILLER_76_3317 ();
 sg13g2_decap_8 FILLER_76_3324 ();
 sg13g2_decap_8 FILLER_76_3331 ();
 sg13g2_fill_1 FILLER_76_3338 ();
 sg13g2_decap_8 FILLER_76_3348 ();
 sg13g2_decap_8 FILLER_76_3355 ();
 sg13g2_decap_8 FILLER_76_3362 ();
 sg13g2_decap_8 FILLER_76_3369 ();
 sg13g2_decap_8 FILLER_76_3376 ();
 sg13g2_decap_8 FILLER_76_3383 ();
 sg13g2_decap_8 FILLER_76_3390 ();
 sg13g2_fill_2 FILLER_76_3397 ();
 sg13g2_fill_1 FILLER_76_3399 ();
 sg13g2_decap_8 FILLER_76_3408 ();
 sg13g2_decap_8 FILLER_76_3415 ();
 sg13g2_decap_8 FILLER_76_3422 ();
 sg13g2_decap_8 FILLER_76_3432 ();
 sg13g2_decap_8 FILLER_76_3439 ();
 sg13g2_decap_8 FILLER_76_3446 ();
 sg13g2_decap_8 FILLER_76_3453 ();
 sg13g2_decap_8 FILLER_76_3460 ();
 sg13g2_decap_8 FILLER_76_3467 ();
 sg13g2_decap_8 FILLER_76_3474 ();
 sg13g2_decap_8 FILLER_76_3481 ();
 sg13g2_decap_8 FILLER_76_3488 ();
 sg13g2_decap_8 FILLER_76_3495 ();
 sg13g2_decap_8 FILLER_76_3502 ();
 sg13g2_decap_8 FILLER_76_3509 ();
 sg13g2_decap_8 FILLER_76_3516 ();
 sg13g2_decap_8 FILLER_76_3523 ();
 sg13g2_decap_8 FILLER_76_3530 ();
 sg13g2_decap_8 FILLER_76_3537 ();
 sg13g2_decap_8 FILLER_76_3544 ();
 sg13g2_decap_8 FILLER_76_3551 ();
 sg13g2_decap_8 FILLER_76_3558 ();
 sg13g2_decap_8 FILLER_76_3565 ();
 sg13g2_decap_8 FILLER_76_3572 ();
 sg13g2_fill_1 FILLER_76_3579 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_decap_8 FILLER_77_28 ();
 sg13g2_decap_8 FILLER_77_35 ();
 sg13g2_decap_8 FILLER_77_42 ();
 sg13g2_decap_8 FILLER_77_49 ();
 sg13g2_decap_8 FILLER_77_56 ();
 sg13g2_decap_8 FILLER_77_63 ();
 sg13g2_decap_8 FILLER_77_70 ();
 sg13g2_decap_8 FILLER_77_77 ();
 sg13g2_decap_8 FILLER_77_84 ();
 sg13g2_decap_8 FILLER_77_91 ();
 sg13g2_decap_8 FILLER_77_98 ();
 sg13g2_fill_2 FILLER_77_105 ();
 sg13g2_decap_8 FILLER_77_112 ();
 sg13g2_decap_8 FILLER_77_119 ();
 sg13g2_decap_8 FILLER_77_126 ();
 sg13g2_decap_4 FILLER_77_133 ();
 sg13g2_fill_1 FILLER_77_137 ();
 sg13g2_fill_2 FILLER_77_166 ();
 sg13g2_fill_1 FILLER_77_168 ();
 sg13g2_fill_2 FILLER_77_173 ();
 sg13g2_fill_1 FILLER_77_175 ();
 sg13g2_decap_8 FILLER_77_185 ();
 sg13g2_decap_8 FILLER_77_192 ();
 sg13g2_decap_4 FILLER_77_199 ();
 sg13g2_fill_1 FILLER_77_203 ();
 sg13g2_decap_8 FILLER_77_209 ();
 sg13g2_decap_8 FILLER_77_216 ();
 sg13g2_decap_8 FILLER_77_223 ();
 sg13g2_decap_8 FILLER_77_230 ();
 sg13g2_decap_8 FILLER_77_237 ();
 sg13g2_decap_4 FILLER_77_270 ();
 sg13g2_decap_8 FILLER_77_313 ();
 sg13g2_decap_4 FILLER_77_320 ();
 sg13g2_fill_2 FILLER_77_324 ();
 sg13g2_decap_8 FILLER_77_342 ();
 sg13g2_decap_8 FILLER_77_349 ();
 sg13g2_fill_1 FILLER_77_356 ();
 sg13g2_decap_8 FILLER_77_385 ();
 sg13g2_decap_8 FILLER_77_392 ();
 sg13g2_decap_8 FILLER_77_399 ();
 sg13g2_fill_2 FILLER_77_406 ();
 sg13g2_decap_8 FILLER_77_424 ();
 sg13g2_decap_8 FILLER_77_431 ();
 sg13g2_decap_8 FILLER_77_462 ();
 sg13g2_decap_8 FILLER_77_469 ();
 sg13g2_decap_4 FILLER_77_476 ();
 sg13g2_fill_1 FILLER_77_480 ();
 sg13g2_decap_8 FILLER_77_502 ();
 sg13g2_decap_8 FILLER_77_535 ();
 sg13g2_decap_8 FILLER_77_542 ();
 sg13g2_decap_8 FILLER_77_549 ();
 sg13g2_decap_8 FILLER_77_556 ();
 sg13g2_fill_1 FILLER_77_563 ();
 sg13g2_decap_8 FILLER_77_607 ();
 sg13g2_fill_2 FILLER_77_619 ();
 sg13g2_fill_1 FILLER_77_621 ();
 sg13g2_fill_2 FILLER_77_627 ();
 sg13g2_fill_1 FILLER_77_629 ();
 sg13g2_decap_8 FILLER_77_635 ();
 sg13g2_decap_8 FILLER_77_642 ();
 sg13g2_decap_8 FILLER_77_684 ();
 sg13g2_decap_4 FILLER_77_691 ();
 sg13g2_fill_2 FILLER_77_695 ();
 sg13g2_fill_2 FILLER_77_706 ();
 sg13g2_fill_1 FILLER_77_708 ();
 sg13g2_decap_8 FILLER_77_724 ();
 sg13g2_decap_8 FILLER_77_731 ();
 sg13g2_decap_8 FILLER_77_738 ();
 sg13g2_decap_8 FILLER_77_745 ();
 sg13g2_fill_2 FILLER_77_761 ();
 sg13g2_fill_1 FILLER_77_783 ();
 sg13g2_decap_8 FILLER_77_789 ();
 sg13g2_decap_8 FILLER_77_796 ();
 sg13g2_decap_8 FILLER_77_803 ();
 sg13g2_decap_8 FILLER_77_810 ();
 sg13g2_fill_1 FILLER_77_817 ();
 sg13g2_fill_1 FILLER_77_842 ();
 sg13g2_fill_1 FILLER_77_848 ();
 sg13g2_decap_8 FILLER_77_854 ();
 sg13g2_decap_8 FILLER_77_861 ();
 sg13g2_decap_4 FILLER_77_868 ();
 sg13g2_fill_1 FILLER_77_872 ();
 sg13g2_fill_2 FILLER_77_888 ();
 sg13g2_decap_8 FILLER_77_897 ();
 sg13g2_decap_8 FILLER_77_904 ();
 sg13g2_decap_8 FILLER_77_911 ();
 sg13g2_decap_8 FILLER_77_963 ();
 sg13g2_decap_4 FILLER_77_984 ();
 sg13g2_fill_1 FILLER_77_988 ();
 sg13g2_decap_4 FILLER_77_999 ();
 sg13g2_fill_2 FILLER_77_1003 ();
 sg13g2_decap_8 FILLER_77_1043 ();
 sg13g2_decap_8 FILLER_77_1050 ();
 sg13g2_decap_8 FILLER_77_1057 ();
 sg13g2_decap_8 FILLER_77_1064 ();
 sg13g2_decap_8 FILLER_77_1071 ();
 sg13g2_fill_2 FILLER_77_1078 ();
 sg13g2_decap_8 FILLER_77_1083 ();
 sg13g2_decap_8 FILLER_77_1090 ();
 sg13g2_decap_8 FILLER_77_1097 ();
 sg13g2_decap_4 FILLER_77_1104 ();
 sg13g2_decap_8 FILLER_77_1144 ();
 sg13g2_fill_2 FILLER_77_1151 ();
 sg13g2_decap_8 FILLER_77_1201 ();
 sg13g2_decap_8 FILLER_77_1208 ();
 sg13g2_decap_8 FILLER_77_1215 ();
 sg13g2_decap_8 FILLER_77_1222 ();
 sg13g2_fill_2 FILLER_77_1245 ();
 sg13g2_decap_8 FILLER_77_1252 ();
 sg13g2_decap_8 FILLER_77_1259 ();
 sg13g2_decap_8 FILLER_77_1266 ();
 sg13g2_decap_8 FILLER_77_1273 ();
 sg13g2_decap_4 FILLER_77_1280 ();
 sg13g2_fill_2 FILLER_77_1284 ();
 sg13g2_decap_8 FILLER_77_1297 ();
 sg13g2_fill_2 FILLER_77_1312 ();
 sg13g2_fill_1 FILLER_77_1314 ();
 sg13g2_decap_8 FILLER_77_1328 ();
 sg13g2_decap_8 FILLER_77_1335 ();
 sg13g2_fill_2 FILLER_77_1342 ();
 sg13g2_fill_1 FILLER_77_1344 ();
 sg13g2_decap_8 FILLER_77_1353 ();
 sg13g2_decap_8 FILLER_77_1360 ();
 sg13g2_fill_1 FILLER_77_1367 ();
 sg13g2_decap_8 FILLER_77_1376 ();
 sg13g2_fill_2 FILLER_77_1383 ();
 sg13g2_decap_8 FILLER_77_1393 ();
 sg13g2_decap_8 FILLER_77_1400 ();
 sg13g2_decap_4 FILLER_77_1407 ();
 sg13g2_fill_1 FILLER_77_1411 ();
 sg13g2_decap_8 FILLER_77_1425 ();
 sg13g2_fill_2 FILLER_77_1432 ();
 sg13g2_decap_4 FILLER_77_1441 ();
 sg13g2_fill_1 FILLER_77_1459 ();
 sg13g2_decap_8 FILLER_77_1470 ();
 sg13g2_decap_8 FILLER_77_1477 ();
 sg13g2_decap_8 FILLER_77_1484 ();
 sg13g2_decap_8 FILLER_77_1491 ();
 sg13g2_decap_8 FILLER_77_1498 ();
 sg13g2_decap_4 FILLER_77_1505 ();
 sg13g2_fill_2 FILLER_77_1509 ();
 sg13g2_decap_8 FILLER_77_1519 ();
 sg13g2_decap_8 FILLER_77_1526 ();
 sg13g2_decap_8 FILLER_77_1533 ();
 sg13g2_decap_4 FILLER_77_1540 ();
 sg13g2_decap_8 FILLER_77_1575 ();
 sg13g2_decap_8 FILLER_77_1582 ();
 sg13g2_decap_8 FILLER_77_1589 ();
 sg13g2_fill_2 FILLER_77_1596 ();
 sg13g2_fill_1 FILLER_77_1598 ();
 sg13g2_decap_8 FILLER_77_1631 ();
 sg13g2_decap_8 FILLER_77_1638 ();
 sg13g2_decap_4 FILLER_77_1645 ();
 sg13g2_fill_1 FILLER_77_1649 ();
 sg13g2_decap_8 FILLER_77_1653 ();
 sg13g2_fill_2 FILLER_77_1660 ();
 sg13g2_decap_8 FILLER_77_1683 ();
 sg13g2_decap_8 FILLER_77_1690 ();
 sg13g2_decap_8 FILLER_77_1697 ();
 sg13g2_fill_1 FILLER_77_1704 ();
 sg13g2_decap_8 FILLER_77_1729 ();
 sg13g2_decap_8 FILLER_77_1736 ();
 sg13g2_decap_8 FILLER_77_1753 ();
 sg13g2_fill_2 FILLER_77_1760 ();
 sg13g2_decap_8 FILLER_77_1788 ();
 sg13g2_decap_4 FILLER_77_1795 ();
 sg13g2_decap_8 FILLER_77_1802 ();
 sg13g2_decap_8 FILLER_77_1809 ();
 sg13g2_decap_8 FILLER_77_1816 ();
 sg13g2_fill_2 FILLER_77_1823 ();
 sg13g2_fill_1 FILLER_77_1825 ();
 sg13g2_decap_4 FILLER_77_1857 ();
 sg13g2_decap_8 FILLER_77_1867 ();
 sg13g2_decap_8 FILLER_77_1874 ();
 sg13g2_fill_1 FILLER_77_1881 ();
 sg13g2_decap_4 FILLER_77_1906 ();
 sg13g2_fill_1 FILLER_77_1910 ();
 sg13g2_decap_8 FILLER_77_1947 ();
 sg13g2_decap_8 FILLER_77_1954 ();
 sg13g2_fill_1 FILLER_77_1961 ();
 sg13g2_decap_8 FILLER_77_2003 ();
 sg13g2_decap_8 FILLER_77_2010 ();
 sg13g2_decap_8 FILLER_77_2017 ();
 sg13g2_decap_8 FILLER_77_2024 ();
 sg13g2_decap_4 FILLER_77_2031 ();
 sg13g2_fill_2 FILLER_77_2035 ();
 sg13g2_fill_2 FILLER_77_2042 ();
 sg13g2_fill_1 FILLER_77_2044 ();
 sg13g2_fill_2 FILLER_77_2050 ();
 sg13g2_decap_8 FILLER_77_2060 ();
 sg13g2_decap_8 FILLER_77_2067 ();
 sg13g2_decap_8 FILLER_77_2074 ();
 sg13g2_decap_4 FILLER_77_2081 ();
 sg13g2_decap_8 FILLER_77_2106 ();
 sg13g2_decap_4 FILLER_77_2113 ();
 sg13g2_fill_1 FILLER_77_2117 ();
 sg13g2_decap_8 FILLER_77_2167 ();
 sg13g2_decap_8 FILLER_77_2174 ();
 sg13g2_decap_8 FILLER_77_2189 ();
 sg13g2_fill_2 FILLER_77_2196 ();
 sg13g2_decap_8 FILLER_77_2247 ();
 sg13g2_decap_8 FILLER_77_2254 ();
 sg13g2_decap_8 FILLER_77_2261 ();
 sg13g2_decap_8 FILLER_77_2268 ();
 sg13g2_decap_8 FILLER_77_2275 ();
 sg13g2_decap_8 FILLER_77_2311 ();
 sg13g2_decap_8 FILLER_77_2318 ();
 sg13g2_decap_8 FILLER_77_2325 ();
 sg13g2_decap_8 FILLER_77_2332 ();
 sg13g2_decap_8 FILLER_77_2339 ();
 sg13g2_decap_8 FILLER_77_2346 ();
 sg13g2_decap_8 FILLER_77_2353 ();
 sg13g2_decap_8 FILLER_77_2360 ();
 sg13g2_decap_8 FILLER_77_2367 ();
 sg13g2_decap_8 FILLER_77_2374 ();
 sg13g2_fill_1 FILLER_77_2381 ();
 sg13g2_fill_2 FILLER_77_2390 ();
 sg13g2_decap_8 FILLER_77_2402 ();
 sg13g2_decap_8 FILLER_77_2409 ();
 sg13g2_decap_8 FILLER_77_2416 ();
 sg13g2_decap_8 FILLER_77_2423 ();
 sg13g2_decap_8 FILLER_77_2430 ();
 sg13g2_decap_8 FILLER_77_2437 ();
 sg13g2_decap_8 FILLER_77_2444 ();
 sg13g2_decap_8 FILLER_77_2451 ();
 sg13g2_fill_2 FILLER_77_2463 ();
 sg13g2_decap_4 FILLER_77_2470 ();
 sg13g2_fill_2 FILLER_77_2474 ();
 sg13g2_decap_8 FILLER_77_2484 ();
 sg13g2_decap_8 FILLER_77_2491 ();
 sg13g2_decap_8 FILLER_77_2498 ();
 sg13g2_fill_2 FILLER_77_2505 ();
 sg13g2_fill_1 FILLER_77_2507 ();
 sg13g2_decap_4 FILLER_77_2518 ();
 sg13g2_decap_8 FILLER_77_2527 ();
 sg13g2_decap_8 FILLER_77_2534 ();
 sg13g2_fill_1 FILLER_77_2541 ();
 sg13g2_fill_2 FILLER_77_2547 ();
 sg13g2_fill_1 FILLER_77_2549 ();
 sg13g2_decap_8 FILLER_77_2581 ();
 sg13g2_decap_8 FILLER_77_2588 ();
 sg13g2_decap_8 FILLER_77_2595 ();
 sg13g2_fill_1 FILLER_77_2628 ();
 sg13g2_fill_2 FILLER_77_2641 ();
 sg13g2_fill_2 FILLER_77_2680 ();
 sg13g2_decap_4 FILLER_77_2692 ();
 sg13g2_fill_2 FILLER_77_2696 ();
 sg13g2_decap_8 FILLER_77_2701 ();
 sg13g2_decap_4 FILLER_77_2708 ();
 sg13g2_fill_1 FILLER_77_2712 ();
 sg13g2_decap_8 FILLER_77_2724 ();
 sg13g2_decap_4 FILLER_77_2741 ();
 sg13g2_decap_4 FILLER_77_2780 ();
 sg13g2_decap_8 FILLER_77_2792 ();
 sg13g2_decap_8 FILLER_77_2799 ();
 sg13g2_decap_8 FILLER_77_2806 ();
 sg13g2_fill_2 FILLER_77_2813 ();
 sg13g2_fill_1 FILLER_77_2815 ();
 sg13g2_decap_8 FILLER_77_2837 ();
 sg13g2_decap_8 FILLER_77_2844 ();
 sg13g2_decap_4 FILLER_77_2851 ();
 sg13g2_fill_2 FILLER_77_2855 ();
 sg13g2_decap_8 FILLER_77_2897 ();
 sg13g2_decap_8 FILLER_77_2904 ();
 sg13g2_decap_8 FILLER_77_2911 ();
 sg13g2_fill_1 FILLER_77_2918 ();
 sg13g2_decap_8 FILLER_77_2927 ();
 sg13g2_decap_4 FILLER_77_2970 ();
 sg13g2_fill_1 FILLER_77_2974 ();
 sg13g2_decap_4 FILLER_77_2980 ();
 sg13g2_decap_8 FILLER_77_3010 ();
 sg13g2_decap_4 FILLER_77_3017 ();
 sg13g2_fill_1 FILLER_77_3021 ();
 sg13g2_decap_8 FILLER_77_3032 ();
 sg13g2_fill_1 FILLER_77_3073 ();
 sg13g2_decap_4 FILLER_77_3134 ();
 sg13g2_decap_8 FILLER_77_3164 ();
 sg13g2_decap_8 FILLER_77_3171 ();
 sg13g2_decap_4 FILLER_77_3178 ();
 sg13g2_decap_4 FILLER_77_3217 ();
 sg13g2_fill_1 FILLER_77_3221 ();
 sg13g2_decap_8 FILLER_77_3231 ();
 sg13g2_decap_8 FILLER_77_3238 ();
 sg13g2_decap_8 FILLER_77_3245 ();
 sg13g2_decap_8 FILLER_77_3252 ();
 sg13g2_decap_4 FILLER_77_3259 ();
 sg13g2_fill_2 FILLER_77_3263 ();
 sg13g2_fill_2 FILLER_77_3291 ();
 sg13g2_decap_8 FILLER_77_3316 ();
 sg13g2_decap_8 FILLER_77_3323 ();
 sg13g2_fill_1 FILLER_77_3330 ();
 sg13g2_decap_8 FILLER_77_3366 ();
 sg13g2_decap_8 FILLER_77_3373 ();
 sg13g2_decap_8 FILLER_77_3380 ();
 sg13g2_decap_8 FILLER_77_3387 ();
 sg13g2_decap_8 FILLER_77_3394 ();
 sg13g2_decap_8 FILLER_77_3401 ();
 sg13g2_decap_8 FILLER_77_3408 ();
 sg13g2_decap_8 FILLER_77_3415 ();
 sg13g2_decap_8 FILLER_77_3422 ();
 sg13g2_decap_8 FILLER_77_3429 ();
 sg13g2_decap_8 FILLER_77_3436 ();
 sg13g2_decap_8 FILLER_77_3443 ();
 sg13g2_decap_8 FILLER_77_3450 ();
 sg13g2_decap_8 FILLER_77_3457 ();
 sg13g2_decap_8 FILLER_77_3464 ();
 sg13g2_decap_8 FILLER_77_3471 ();
 sg13g2_decap_8 FILLER_77_3478 ();
 sg13g2_decap_8 FILLER_77_3485 ();
 sg13g2_decap_8 FILLER_77_3492 ();
 sg13g2_decap_8 FILLER_77_3499 ();
 sg13g2_decap_8 FILLER_77_3506 ();
 sg13g2_decap_8 FILLER_77_3513 ();
 sg13g2_decap_8 FILLER_77_3520 ();
 sg13g2_decap_8 FILLER_77_3527 ();
 sg13g2_decap_8 FILLER_77_3534 ();
 sg13g2_decap_8 FILLER_77_3541 ();
 sg13g2_decap_8 FILLER_77_3548 ();
 sg13g2_decap_8 FILLER_77_3555 ();
 sg13g2_decap_8 FILLER_77_3562 ();
 sg13g2_decap_8 FILLER_77_3569 ();
 sg13g2_decap_4 FILLER_77_3576 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_decap_8 FILLER_78_28 ();
 sg13g2_decap_8 FILLER_78_35 ();
 sg13g2_decap_8 FILLER_78_42 ();
 sg13g2_decap_8 FILLER_78_49 ();
 sg13g2_decap_8 FILLER_78_56 ();
 sg13g2_decap_8 FILLER_78_63 ();
 sg13g2_decap_8 FILLER_78_70 ();
 sg13g2_decap_8 FILLER_78_77 ();
 sg13g2_decap_8 FILLER_78_84 ();
 sg13g2_decap_8 FILLER_78_91 ();
 sg13g2_decap_8 FILLER_78_98 ();
 sg13g2_decap_8 FILLER_78_105 ();
 sg13g2_decap_4 FILLER_78_112 ();
 sg13g2_fill_2 FILLER_78_116 ();
 sg13g2_fill_2 FILLER_78_144 ();
 sg13g2_fill_1 FILLER_78_146 ();
 sg13g2_decap_8 FILLER_78_175 ();
 sg13g2_decap_8 FILLER_78_182 ();
 sg13g2_decap_8 FILLER_78_189 ();
 sg13g2_fill_2 FILLER_78_196 ();
 sg13g2_fill_1 FILLER_78_198 ();
 sg13g2_decap_8 FILLER_78_224 ();
 sg13g2_decap_8 FILLER_78_231 ();
 sg13g2_decap_8 FILLER_78_238 ();
 sg13g2_decap_8 FILLER_78_245 ();
 sg13g2_decap_8 FILLER_78_252 ();
 sg13g2_fill_2 FILLER_78_259 ();
 sg13g2_fill_2 FILLER_78_275 ();
 sg13g2_fill_1 FILLER_78_277 ();
 sg13g2_decap_8 FILLER_78_313 ();
 sg13g2_decap_8 FILLER_78_320 ();
 sg13g2_decap_8 FILLER_78_327 ();
 sg13g2_decap_8 FILLER_78_334 ();
 sg13g2_decap_8 FILLER_78_341 ();
 sg13g2_fill_2 FILLER_78_348 ();
 sg13g2_fill_2 FILLER_78_395 ();
 sg13g2_fill_1 FILLER_78_397 ();
 sg13g2_decap_4 FILLER_78_419 ();
 sg13g2_fill_1 FILLER_78_423 ();
 sg13g2_fill_1 FILLER_78_444 ();
 sg13g2_fill_2 FILLER_78_450 ();
 sg13g2_decap_8 FILLER_78_464 ();
 sg13g2_decap_8 FILLER_78_471 ();
 sg13g2_decap_8 FILLER_78_478 ();
 sg13g2_fill_2 FILLER_78_485 ();
 sg13g2_fill_1 FILLER_78_487 ();
 sg13g2_decap_8 FILLER_78_491 ();
 sg13g2_decap_4 FILLER_78_498 ();
 sg13g2_fill_2 FILLER_78_502 ();
 sg13g2_decap_4 FILLER_78_520 ();
 sg13g2_fill_1 FILLER_78_563 ();
 sg13g2_fill_1 FILLER_78_610 ();
 sg13g2_fill_1 FILLER_78_637 ();
 sg13g2_fill_1 FILLER_78_642 ();
 sg13g2_decap_8 FILLER_78_653 ();
 sg13g2_decap_8 FILLER_78_660 ();
 sg13g2_decap_8 FILLER_78_667 ();
 sg13g2_decap_8 FILLER_78_674 ();
 sg13g2_decap_8 FILLER_78_681 ();
 sg13g2_decap_8 FILLER_78_688 ();
 sg13g2_decap_8 FILLER_78_695 ();
 sg13g2_fill_1 FILLER_78_702 ();
 sg13g2_decap_8 FILLER_78_731 ();
 sg13g2_decap_8 FILLER_78_738 ();
 sg13g2_decap_4 FILLER_78_745 ();
 sg13g2_fill_1 FILLER_78_791 ();
 sg13g2_decap_8 FILLER_78_816 ();
 sg13g2_fill_2 FILLER_78_823 ();
 sg13g2_fill_1 FILLER_78_825 ();
 sg13g2_fill_2 FILLER_78_848 ();
 sg13g2_fill_2 FILLER_78_858 ();
 sg13g2_fill_1 FILLER_78_860 ();
 sg13g2_decap_8 FILLER_78_905 ();
 sg13g2_decap_8 FILLER_78_912 ();
 sg13g2_decap_4 FILLER_78_919 ();
 sg13g2_fill_2 FILLER_78_923 ();
 sg13g2_fill_2 FILLER_78_960 ();
 sg13g2_fill_1 FILLER_78_962 ();
 sg13g2_fill_2 FILLER_78_972 ();
 sg13g2_decap_4 FILLER_78_992 ();
 sg13g2_decap_8 FILLER_78_1021 ();
 sg13g2_decap_8 FILLER_78_1028 ();
 sg13g2_decap_8 FILLER_78_1035 ();
 sg13g2_decap_8 FILLER_78_1042 ();
 sg13g2_decap_8 FILLER_78_1049 ();
 sg13g2_fill_2 FILLER_78_1056 ();
 sg13g2_fill_1 FILLER_78_1058 ();
 sg13g2_decap_4 FILLER_78_1080 ();
 sg13g2_fill_2 FILLER_78_1084 ();
 sg13g2_decap_8 FILLER_78_1099 ();
 sg13g2_decap_4 FILLER_78_1106 ();
 sg13g2_fill_2 FILLER_78_1154 ();
 sg13g2_decap_8 FILLER_78_1159 ();
 sg13g2_fill_1 FILLER_78_1166 ();
 sg13g2_decap_8 FILLER_78_1198 ();
 sg13g2_decap_8 FILLER_78_1205 ();
 sg13g2_decap_8 FILLER_78_1212 ();
 sg13g2_decap_8 FILLER_78_1219 ();
 sg13g2_fill_2 FILLER_78_1226 ();
 sg13g2_fill_1 FILLER_78_1228 ();
 sg13g2_decap_8 FILLER_78_1245 ();
 sg13g2_decap_8 FILLER_78_1252 ();
 sg13g2_decap_8 FILLER_78_1279 ();
 sg13g2_decap_4 FILLER_78_1286 ();
 sg13g2_fill_1 FILLER_78_1290 ();
 sg13g2_decap_8 FILLER_78_1308 ();
 sg13g2_decap_8 FILLER_78_1315 ();
 sg13g2_decap_8 FILLER_78_1322 ();
 sg13g2_fill_1 FILLER_78_1329 ();
 sg13g2_decap_8 FILLER_78_1338 ();
 sg13g2_decap_8 FILLER_78_1345 ();
 sg13g2_decap_8 FILLER_78_1352 ();
 sg13g2_decap_8 FILLER_78_1359 ();
 sg13g2_decap_4 FILLER_78_1366 ();
 sg13g2_fill_1 FILLER_78_1377 ();
 sg13g2_decap_8 FILLER_78_1394 ();
 sg13g2_decap_8 FILLER_78_1401 ();
 sg13g2_decap_4 FILLER_78_1408 ();
 sg13g2_fill_2 FILLER_78_1412 ();
 sg13g2_decap_8 FILLER_78_1462 ();
 sg13g2_decap_8 FILLER_78_1495 ();
 sg13g2_decap_8 FILLER_78_1502 ();
 sg13g2_decap_8 FILLER_78_1509 ();
 sg13g2_fill_2 FILLER_78_1516 ();
 sg13g2_fill_1 FILLER_78_1518 ();
 sg13g2_decap_4 FILLER_78_1525 ();
 sg13g2_decap_8 FILLER_78_1535 ();
 sg13g2_decap_8 FILLER_78_1542 ();
 sg13g2_decap_8 FILLER_78_1549 ();
 sg13g2_decap_8 FILLER_78_1556 ();
 sg13g2_decap_8 FILLER_78_1563 ();
 sg13g2_decap_8 FILLER_78_1570 ();
 sg13g2_decap_8 FILLER_78_1577 ();
 sg13g2_fill_2 FILLER_78_1584 ();
 sg13g2_fill_1 FILLER_78_1586 ();
 sg13g2_decap_8 FILLER_78_1629 ();
 sg13g2_decap_8 FILLER_78_1636 ();
 sg13g2_fill_1 FILLER_78_1643 ();
 sg13g2_fill_1 FILLER_78_1649 ();
 sg13g2_decap_8 FILLER_78_1671 ();
 sg13g2_decap_8 FILLER_78_1678 ();
 sg13g2_decap_8 FILLER_78_1685 ();
 sg13g2_decap_8 FILLER_78_1692 ();
 sg13g2_fill_1 FILLER_78_1699 ();
 sg13g2_decap_4 FILLER_78_1739 ();
 sg13g2_decap_8 FILLER_78_1769 ();
 sg13g2_decap_8 FILLER_78_1776 ();
 sg13g2_fill_2 FILLER_78_1783 ();
 sg13g2_decap_8 FILLER_78_1824 ();
 sg13g2_fill_2 FILLER_78_1831 ();
 sg13g2_decap_4 FILLER_78_1856 ();
 sg13g2_fill_1 FILLER_78_1874 ();
 sg13g2_decap_8 FILLER_78_1933 ();
 sg13g2_decap_4 FILLER_78_1940 ();
 sg13g2_fill_1 FILLER_78_1944 ();
 sg13g2_decap_8 FILLER_78_1995 ();
 sg13g2_decap_8 FILLER_78_2002 ();
 sg13g2_decap_8 FILLER_78_2009 ();
 sg13g2_decap_8 FILLER_78_2016 ();
 sg13g2_decap_4 FILLER_78_2023 ();
 sg13g2_fill_1 FILLER_78_2027 ();
 sg13g2_decap_8 FILLER_78_2064 ();
 sg13g2_fill_1 FILLER_78_2089 ();
 sg13g2_decap_8 FILLER_78_2110 ();
 sg13g2_decap_8 FILLER_78_2117 ();
 sg13g2_fill_2 FILLER_78_2124 ();
 sg13g2_fill_1 FILLER_78_2126 ();
 sg13g2_decap_8 FILLER_78_2161 ();
 sg13g2_decap_8 FILLER_78_2168 ();
 sg13g2_fill_1 FILLER_78_2175 ();
 sg13g2_decap_4 FILLER_78_2245 ();
 sg13g2_decap_4 FILLER_78_2260 ();
 sg13g2_fill_1 FILLER_78_2264 ();
 sg13g2_fill_2 FILLER_78_2284 ();
 sg13g2_fill_2 FILLER_78_2302 ();
 sg13g2_decap_8 FILLER_78_2320 ();
 sg13g2_fill_1 FILLER_78_2327 ();
 sg13g2_fill_1 FILLER_78_2347 ();
 sg13g2_decap_8 FILLER_78_2367 ();
 sg13g2_fill_1 FILLER_78_2374 ();
 sg13g2_decap_8 FILLER_78_2423 ();
 sg13g2_decap_8 FILLER_78_2430 ();
 sg13g2_decap_4 FILLER_78_2450 ();
 sg13g2_fill_2 FILLER_78_2454 ();
 sg13g2_decap_8 FILLER_78_2486 ();
 sg13g2_decap_4 FILLER_78_2493 ();
 sg13g2_fill_1 FILLER_78_2497 ();
 sg13g2_decap_8 FILLER_78_2524 ();
 sg13g2_decap_8 FILLER_78_2531 ();
 sg13g2_decap_8 FILLER_78_2538 ();
 sg13g2_fill_2 FILLER_78_2545 ();
 sg13g2_decap_8 FILLER_78_2551 ();
 sg13g2_decap_8 FILLER_78_2558 ();
 sg13g2_decap_8 FILLER_78_2565 ();
 sg13g2_fill_1 FILLER_78_2572 ();
 sg13g2_decap_8 FILLER_78_2581 ();
 sg13g2_decap_8 FILLER_78_2588 ();
 sg13g2_fill_1 FILLER_78_2595 ();
 sg13g2_decap_8 FILLER_78_2641 ();
 sg13g2_decap_8 FILLER_78_2648 ();
 sg13g2_decap_8 FILLER_78_2655 ();
 sg13g2_fill_2 FILLER_78_2662 ();
 sg13g2_fill_1 FILLER_78_2664 ();
 sg13g2_decap_8 FILLER_78_2675 ();
 sg13g2_decap_8 FILLER_78_2708 ();
 sg13g2_decap_8 FILLER_78_2715 ();
 sg13g2_decap_4 FILLER_78_2722 ();
 sg13g2_fill_2 FILLER_78_2731 ();
 sg13g2_fill_1 FILLER_78_2733 ();
 sg13g2_decap_8 FILLER_78_2739 ();
 sg13g2_decap_8 FILLER_78_2787 ();
 sg13g2_decap_8 FILLER_78_2794 ();
 sg13g2_fill_2 FILLER_78_2809 ();
 sg13g2_fill_1 FILLER_78_2811 ();
 sg13g2_decap_8 FILLER_78_2838 ();
 sg13g2_decap_8 FILLER_78_2845 ();
 sg13g2_fill_2 FILLER_78_2852 ();
 sg13g2_fill_2 FILLER_78_2906 ();
 sg13g2_fill_2 FILLER_78_2916 ();
 sg13g2_fill_1 FILLER_78_2918 ();
 sg13g2_fill_1 FILLER_78_2935 ();
 sg13g2_decap_8 FILLER_78_2962 ();
 sg13g2_decap_8 FILLER_78_2969 ();
 sg13g2_decap_8 FILLER_78_2976 ();
 sg13g2_fill_1 FILLER_78_2983 ();
 sg13g2_decap_8 FILLER_78_2987 ();
 sg13g2_fill_2 FILLER_78_2994 ();
 sg13g2_fill_1 FILLER_78_2996 ();
 sg13g2_decap_8 FILLER_78_3007 ();
 sg13g2_decap_8 FILLER_78_3014 ();
 sg13g2_decap_8 FILLER_78_3021 ();
 sg13g2_fill_2 FILLER_78_3028 ();
 sg13g2_decap_8 FILLER_78_3056 ();
 sg13g2_decap_4 FILLER_78_3063 ();
 sg13g2_fill_2 FILLER_78_3067 ();
 sg13g2_decap_8 FILLER_78_3105 ();
 sg13g2_decap_8 FILLER_78_3112 ();
 sg13g2_decap_4 FILLER_78_3119 ();
 sg13g2_fill_2 FILLER_78_3123 ();
 sg13g2_decap_8 FILLER_78_3169 ();
 sg13g2_decap_8 FILLER_78_3176 ();
 sg13g2_decap_8 FILLER_78_3183 ();
 sg13g2_decap_8 FILLER_78_3190 ();
 sg13g2_fill_1 FILLER_78_3197 ();
 sg13g2_fill_2 FILLER_78_3216 ();
 sg13g2_decap_8 FILLER_78_3226 ();
 sg13g2_decap_8 FILLER_78_3253 ();
 sg13g2_decap_4 FILLER_78_3286 ();
 sg13g2_fill_2 FILLER_78_3290 ();
 sg13g2_decap_8 FILLER_78_3318 ();
 sg13g2_decap_4 FILLER_78_3325 ();
 sg13g2_fill_1 FILLER_78_3329 ();
 sg13g2_decap_8 FILLER_78_3362 ();
 sg13g2_decap_8 FILLER_78_3369 ();
 sg13g2_decap_8 FILLER_78_3376 ();
 sg13g2_decap_8 FILLER_78_3383 ();
 sg13g2_decap_8 FILLER_78_3390 ();
 sg13g2_decap_8 FILLER_78_3397 ();
 sg13g2_decap_8 FILLER_78_3404 ();
 sg13g2_decap_8 FILLER_78_3411 ();
 sg13g2_decap_8 FILLER_78_3418 ();
 sg13g2_decap_8 FILLER_78_3425 ();
 sg13g2_decap_8 FILLER_78_3432 ();
 sg13g2_decap_8 FILLER_78_3439 ();
 sg13g2_decap_8 FILLER_78_3446 ();
 sg13g2_decap_8 FILLER_78_3453 ();
 sg13g2_decap_8 FILLER_78_3460 ();
 sg13g2_decap_8 FILLER_78_3467 ();
 sg13g2_decap_8 FILLER_78_3474 ();
 sg13g2_decap_8 FILLER_78_3481 ();
 sg13g2_decap_8 FILLER_78_3488 ();
 sg13g2_decap_8 FILLER_78_3495 ();
 sg13g2_decap_8 FILLER_78_3502 ();
 sg13g2_decap_8 FILLER_78_3509 ();
 sg13g2_decap_8 FILLER_78_3516 ();
 sg13g2_decap_8 FILLER_78_3523 ();
 sg13g2_decap_8 FILLER_78_3530 ();
 sg13g2_decap_8 FILLER_78_3537 ();
 sg13g2_decap_8 FILLER_78_3544 ();
 sg13g2_decap_8 FILLER_78_3551 ();
 sg13g2_decap_8 FILLER_78_3558 ();
 sg13g2_decap_8 FILLER_78_3565 ();
 sg13g2_decap_8 FILLER_78_3572 ();
 sg13g2_fill_1 FILLER_78_3579 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_decap_8 FILLER_79_35 ();
 sg13g2_decap_8 FILLER_79_42 ();
 sg13g2_decap_8 FILLER_79_49 ();
 sg13g2_decap_8 FILLER_79_56 ();
 sg13g2_decap_8 FILLER_79_63 ();
 sg13g2_decap_8 FILLER_79_70 ();
 sg13g2_decap_8 FILLER_79_77 ();
 sg13g2_decap_8 FILLER_79_84 ();
 sg13g2_decap_8 FILLER_79_91 ();
 sg13g2_decap_8 FILLER_79_98 ();
 sg13g2_decap_8 FILLER_79_105 ();
 sg13g2_decap_8 FILLER_79_112 ();
 sg13g2_decap_8 FILLER_79_119 ();
 sg13g2_decap_8 FILLER_79_126 ();
 sg13g2_decap_4 FILLER_79_133 ();
 sg13g2_fill_2 FILLER_79_137 ();
 sg13g2_decap_8 FILLER_79_173 ();
 sg13g2_decap_8 FILLER_79_180 ();
 sg13g2_decap_8 FILLER_79_187 ();
 sg13g2_fill_2 FILLER_79_194 ();
 sg13g2_decap_8 FILLER_79_231 ();
 sg13g2_decap_8 FILLER_79_238 ();
 sg13g2_decap_8 FILLER_79_245 ();
 sg13g2_decap_8 FILLER_79_252 ();
 sg13g2_decap_8 FILLER_79_259 ();
 sg13g2_fill_2 FILLER_79_266 ();
 sg13g2_fill_2 FILLER_79_272 ();
 sg13g2_fill_2 FILLER_79_279 ();
 sg13g2_fill_1 FILLER_79_281 ();
 sg13g2_fill_2 FILLER_79_318 ();
 sg13g2_decap_8 FILLER_79_333 ();
 sg13g2_decap_4 FILLER_79_340 ();
 sg13g2_fill_2 FILLER_79_373 ();
 sg13g2_decap_8 FILLER_79_392 ();
 sg13g2_decap_8 FILLER_79_399 ();
 sg13g2_fill_2 FILLER_79_406 ();
 sg13g2_fill_1 FILLER_79_408 ();
 sg13g2_fill_1 FILLER_79_414 ();
 sg13g2_fill_2 FILLER_79_428 ();
 sg13g2_fill_1 FILLER_79_430 ();
 sg13g2_decap_8 FILLER_79_435 ();
 sg13g2_decap_8 FILLER_79_442 ();
 sg13g2_decap_8 FILLER_79_449 ();
 sg13g2_decap_4 FILLER_79_456 ();
 sg13g2_fill_2 FILLER_79_460 ();
 sg13g2_decap_4 FILLER_79_470 ();
 sg13g2_decap_4 FILLER_79_496 ();
 sg13g2_fill_1 FILLER_79_500 ();
 sg13g2_decap_8 FILLER_79_521 ();
 sg13g2_fill_2 FILLER_79_528 ();
 sg13g2_decap_8 FILLER_79_539 ();
 sg13g2_decap_8 FILLER_79_546 ();
 sg13g2_decap_8 FILLER_79_553 ();
 sg13g2_fill_1 FILLER_79_595 ();
 sg13g2_decap_4 FILLER_79_601 ();
 sg13g2_fill_1 FILLER_79_605 ();
 sg13g2_fill_2 FILLER_79_641 ();
 sg13g2_fill_1 FILLER_79_643 ();
 sg13g2_decap_8 FILLER_79_674 ();
 sg13g2_decap_8 FILLER_79_681 ();
 sg13g2_decap_8 FILLER_79_688 ();
 sg13g2_decap_8 FILLER_79_695 ();
 sg13g2_decap_8 FILLER_79_702 ();
 sg13g2_decap_8 FILLER_79_738 ();
 sg13g2_decap_8 FILLER_79_745 ();
 sg13g2_decap_8 FILLER_79_752 ();
 sg13g2_decap_8 FILLER_79_768 ();
 sg13g2_fill_2 FILLER_79_780 ();
 sg13g2_fill_1 FILLER_79_782 ();
 sg13g2_decap_4 FILLER_79_788 ();
 sg13g2_decap_8 FILLER_79_809 ();
 sg13g2_decap_8 FILLER_79_816 ();
 sg13g2_decap_8 FILLER_79_823 ();
 sg13g2_decap_4 FILLER_79_830 ();
 sg13g2_fill_2 FILLER_79_834 ();
 sg13g2_decap_8 FILLER_79_840 ();
 sg13g2_decap_4 FILLER_79_847 ();
 sg13g2_fill_2 FILLER_79_851 ();
 sg13g2_decap_8 FILLER_79_857 ();
 sg13g2_decap_8 FILLER_79_864 ();
 sg13g2_fill_1 FILLER_79_871 ();
 sg13g2_decap_8 FILLER_79_899 ();
 sg13g2_decap_8 FILLER_79_906 ();
 sg13g2_decap_8 FILLER_79_913 ();
 sg13g2_decap_8 FILLER_79_920 ();
 sg13g2_decap_4 FILLER_79_927 ();
 sg13g2_fill_1 FILLER_79_931 ();
 sg13g2_fill_2 FILLER_79_937 ();
 sg13g2_fill_1 FILLER_79_939 ();
 sg13g2_fill_2 FILLER_79_948 ();
 sg13g2_fill_1 FILLER_79_950 ();
 sg13g2_decap_8 FILLER_79_955 ();
 sg13g2_fill_2 FILLER_79_962 ();
 sg13g2_decap_8 FILLER_79_999 ();
 sg13g2_decap_8 FILLER_79_1084 ();
 sg13g2_decap_8 FILLER_79_1091 ();
 sg13g2_decap_8 FILLER_79_1098 ();
 sg13g2_decap_8 FILLER_79_1105 ();
 sg13g2_fill_1 FILLER_79_1112 ();
 sg13g2_decap_8 FILLER_79_1139 ();
 sg13g2_decap_8 FILLER_79_1146 ();
 sg13g2_decap_8 FILLER_79_1153 ();
 sg13g2_decap_8 FILLER_79_1160 ();
 sg13g2_fill_2 FILLER_79_1167 ();
 sg13g2_decap_8 FILLER_79_1208 ();
 sg13g2_decap_8 FILLER_79_1215 ();
 sg13g2_decap_8 FILLER_79_1222 ();
 sg13g2_decap_8 FILLER_79_1229 ();
 sg13g2_decap_8 FILLER_79_1236 ();
 sg13g2_fill_2 FILLER_79_1243 ();
 sg13g2_fill_1 FILLER_79_1245 ();
 sg13g2_decap_8 FILLER_79_1298 ();
 sg13g2_decap_4 FILLER_79_1305 ();
 sg13g2_fill_1 FILLER_79_1309 ();
 sg13g2_decap_4 FILLER_79_1323 ();
 sg13g2_fill_2 FILLER_79_1335 ();
 sg13g2_fill_1 FILLER_79_1342 ();
 sg13g2_decap_8 FILLER_79_1360 ();
 sg13g2_decap_4 FILLER_79_1367 ();
 sg13g2_fill_1 FILLER_79_1371 ();
 sg13g2_decap_8 FILLER_79_1400 ();
 sg13g2_fill_1 FILLER_79_1407 ();
 sg13g2_decap_8 FILLER_79_1428 ();
 sg13g2_decap_8 FILLER_79_1444 ();
 sg13g2_decap_8 FILLER_79_1451 ();
 sg13g2_decap_8 FILLER_79_1458 ();
 sg13g2_decap_8 FILLER_79_1465 ();
 sg13g2_decap_8 FILLER_79_1472 ();
 sg13g2_decap_8 FILLER_79_1479 ();
 sg13g2_decap_8 FILLER_79_1486 ();
 sg13g2_decap_8 FILLER_79_1493 ();
 sg13g2_decap_8 FILLER_79_1500 ();
 sg13g2_fill_1 FILLER_79_1507 ();
 sg13g2_decap_8 FILLER_79_1542 ();
 sg13g2_decap_8 FILLER_79_1549 ();
 sg13g2_decap_8 FILLER_79_1556 ();
 sg13g2_decap_8 FILLER_79_1563 ();
 sg13g2_decap_8 FILLER_79_1570 ();
 sg13g2_decap_8 FILLER_79_1577 ();
 sg13g2_decap_4 FILLER_79_1584 ();
 sg13g2_fill_2 FILLER_79_1588 ();
 sg13g2_decap_8 FILLER_79_1622 ();
 sg13g2_decap_8 FILLER_79_1629 ();
 sg13g2_decap_4 FILLER_79_1636 ();
 sg13g2_fill_1 FILLER_79_1640 ();
 sg13g2_fill_2 FILLER_79_1649 ();
 sg13g2_decap_8 FILLER_79_1668 ();
 sg13g2_decap_8 FILLER_79_1675 ();
 sg13g2_decap_8 FILLER_79_1682 ();
 sg13g2_decap_8 FILLER_79_1689 ();
 sg13g2_decap_4 FILLER_79_1696 ();
 sg13g2_decap_8 FILLER_79_1726 ();
 sg13g2_decap_8 FILLER_79_1733 ();
 sg13g2_decap_8 FILLER_79_1740 ();
 sg13g2_decap_8 FILLER_79_1747 ();
 sg13g2_decap_4 FILLER_79_1754 ();
 sg13g2_decap_8 FILLER_79_1784 ();
 sg13g2_decap_8 FILLER_79_1791 ();
 sg13g2_decap_8 FILLER_79_1798 ();
 sg13g2_decap_8 FILLER_79_1805 ();
 sg13g2_decap_4 FILLER_79_1812 ();
 sg13g2_fill_2 FILLER_79_1816 ();
 sg13g2_decap_8 FILLER_79_1831 ();
 sg13g2_decap_4 FILLER_79_1838 ();
 sg13g2_fill_2 FILLER_79_1842 ();
 sg13g2_decap_8 FILLER_79_1862 ();
 sg13g2_decap_8 FILLER_79_1869 ();
 sg13g2_decap_4 FILLER_79_1876 ();
 sg13g2_fill_1 FILLER_79_1880 ();
 sg13g2_decap_8 FILLER_79_1886 ();
 sg13g2_decap_8 FILLER_79_1893 ();
 sg13g2_decap_8 FILLER_79_1900 ();
 sg13g2_decap_8 FILLER_79_1907 ();
 sg13g2_decap_8 FILLER_79_1914 ();
 sg13g2_decap_8 FILLER_79_1921 ();
 sg13g2_decap_8 FILLER_79_1928 ();
 sg13g2_decap_8 FILLER_79_1935 ();
 sg13g2_decap_8 FILLER_79_1942 ();
 sg13g2_decap_8 FILLER_79_1949 ();
 sg13g2_decap_8 FILLER_79_1956 ();
 sg13g2_decap_8 FILLER_79_2001 ();
 sg13g2_decap_8 FILLER_79_2008 ();
 sg13g2_decap_8 FILLER_79_2015 ();
 sg13g2_decap_8 FILLER_79_2022 ();
 sg13g2_decap_8 FILLER_79_2029 ();
 sg13g2_fill_2 FILLER_79_2036 ();
 sg13g2_fill_1 FILLER_79_2038 ();
 sg13g2_decap_4 FILLER_79_2044 ();
 sg13g2_fill_1 FILLER_79_2048 ();
 sg13g2_decap_8 FILLER_79_2054 ();
 sg13g2_decap_8 FILLER_79_2061 ();
 sg13g2_decap_8 FILLER_79_2068 ();
 sg13g2_decap_4 FILLER_79_2075 ();
 sg13g2_fill_2 FILLER_79_2079 ();
 sg13g2_fill_2 FILLER_79_2086 ();
 sg13g2_fill_1 FILLER_79_2088 ();
 sg13g2_decap_8 FILLER_79_2104 ();
 sg13g2_decap_8 FILLER_79_2111 ();
 sg13g2_decap_8 FILLER_79_2118 ();
 sg13g2_decap_8 FILLER_79_2125 ();
 sg13g2_fill_1 FILLER_79_2132 ();
 sg13g2_decap_8 FILLER_79_2151 ();
 sg13g2_decap_8 FILLER_79_2158 ();
 sg13g2_decap_8 FILLER_79_2165 ();
 sg13g2_decap_8 FILLER_79_2172 ();
 sg13g2_decap_8 FILLER_79_2179 ();
 sg13g2_decap_8 FILLER_79_2186 ();
 sg13g2_decap_8 FILLER_79_2193 ();
 sg13g2_decap_8 FILLER_79_2200 ();
 sg13g2_fill_2 FILLER_79_2207 ();
 sg13g2_fill_1 FILLER_79_2209 ();
 sg13g2_fill_2 FILLER_79_2219 ();
 sg13g2_fill_2 FILLER_79_2234 ();
 sg13g2_decap_8 FILLER_79_2262 ();
 sg13g2_decap_8 FILLER_79_2269 ();
 sg13g2_decap_8 FILLER_79_2276 ();
 sg13g2_fill_1 FILLER_79_2283 ();
 sg13g2_decap_8 FILLER_79_2310 ();
 sg13g2_fill_1 FILLER_79_2317 ();
 sg13g2_fill_2 FILLER_79_2344 ();
 sg13g2_decap_8 FILLER_79_2398 ();
 sg13g2_decap_8 FILLER_79_2405 ();
 sg13g2_decap_8 FILLER_79_2412 ();
 sg13g2_decap_8 FILLER_79_2419 ();
 sg13g2_fill_2 FILLER_79_2439 ();
 sg13g2_decap_8 FILLER_79_2489 ();
 sg13g2_decap_8 FILLER_79_2496 ();
 sg13g2_decap_8 FILLER_79_2503 ();
 sg13g2_decap_4 FILLER_79_2510 ();
 sg13g2_fill_1 FILLER_79_2514 ();
 sg13g2_decap_8 FILLER_79_2541 ();
 sg13g2_decap_4 FILLER_79_2548 ();
 sg13g2_decap_8 FILLER_79_2578 ();
 sg13g2_decap_8 FILLER_79_2585 ();
 sg13g2_decap_8 FILLER_79_2592 ();
 sg13g2_decap_4 FILLER_79_2599 ();
 sg13g2_fill_1 FILLER_79_2603 ();
 sg13g2_decap_8 FILLER_79_2612 ();
 sg13g2_decap_8 FILLER_79_2619 ();
 sg13g2_decap_8 FILLER_79_2626 ();
 sg13g2_decap_8 FILLER_79_2633 ();
 sg13g2_decap_8 FILLER_79_2640 ();
 sg13g2_decap_8 FILLER_79_2647 ();
 sg13g2_decap_4 FILLER_79_2654 ();
 sg13g2_decap_8 FILLER_79_2710 ();
 sg13g2_fill_2 FILLER_79_2717 ();
 sg13g2_fill_1 FILLER_79_2719 ();
 sg13g2_decap_8 FILLER_79_2728 ();
 sg13g2_decap_8 FILLER_79_2735 ();
 sg13g2_decap_8 FILLER_79_2742 ();
 sg13g2_fill_2 FILLER_79_2749 ();
 sg13g2_fill_1 FILLER_79_2751 ();
 sg13g2_decap_8 FILLER_79_2778 ();
 sg13g2_decap_8 FILLER_79_2785 ();
 sg13g2_decap_8 FILLER_79_2792 ();
 sg13g2_fill_1 FILLER_79_2799 ();
 sg13g2_decap_8 FILLER_79_2805 ();
 sg13g2_fill_2 FILLER_79_2812 ();
 sg13g2_decap_8 FILLER_79_2840 ();
 sg13g2_decap_8 FILLER_79_2847 ();
 sg13g2_decap_4 FILLER_79_2854 ();
 sg13g2_decap_8 FILLER_79_2898 ();
 sg13g2_decap_8 FILLER_79_2905 ();
 sg13g2_decap_8 FILLER_79_2912 ();
 sg13g2_fill_2 FILLER_79_2919 ();
 sg13g2_fill_1 FILLER_79_2921 ();
 sg13g2_fill_1 FILLER_79_2926 ();
 sg13g2_decap_8 FILLER_79_2960 ();
 sg13g2_fill_2 FILLER_79_2967 ();
 sg13g2_fill_1 FILLER_79_2969 ();
 sg13g2_decap_8 FILLER_79_2996 ();
 sg13g2_decap_8 FILLER_79_3029 ();
 sg13g2_decap_8 FILLER_79_3036 ();
 sg13g2_decap_8 FILLER_79_3043 ();
 sg13g2_decap_8 FILLER_79_3050 ();
 sg13g2_decap_8 FILLER_79_3057 ();
 sg13g2_decap_8 FILLER_79_3064 ();
 sg13g2_fill_2 FILLER_79_3071 ();
 sg13g2_fill_1 FILLER_79_3073 ();
 sg13g2_decap_8 FILLER_79_3084 ();
 sg13g2_decap_8 FILLER_79_3091 ();
 sg13g2_decap_8 FILLER_79_3098 ();
 sg13g2_decap_8 FILLER_79_3105 ();
 sg13g2_decap_8 FILLER_79_3112 ();
 sg13g2_decap_8 FILLER_79_3119 ();
 sg13g2_decap_8 FILLER_79_3126 ();
 sg13g2_decap_8 FILLER_79_3133 ();
 sg13g2_decap_8 FILLER_79_3140 ();
 sg13g2_fill_1 FILLER_79_3147 ();
 sg13g2_decap_8 FILLER_79_3174 ();
 sg13g2_decap_8 FILLER_79_3181 ();
 sg13g2_decap_4 FILLER_79_3188 ();
 sg13g2_decap_8 FILLER_79_3218 ();
 sg13g2_fill_2 FILLER_79_3225 ();
 sg13g2_decap_8 FILLER_79_3253 ();
 sg13g2_decap_8 FILLER_79_3260 ();
 sg13g2_decap_4 FILLER_79_3267 ();
 sg13g2_fill_1 FILLER_79_3271 ();
 sg13g2_decap_8 FILLER_79_3277 ();
 sg13g2_decap_4 FILLER_79_3284 ();
 sg13g2_decap_8 FILLER_79_3314 ();
 sg13g2_decap_8 FILLER_79_3321 ();
 sg13g2_decap_4 FILLER_79_3328 ();
 sg13g2_fill_1 FILLER_79_3332 ();
 sg13g2_decap_8 FILLER_79_3343 ();
 sg13g2_decap_8 FILLER_79_3350 ();
 sg13g2_decap_8 FILLER_79_3357 ();
 sg13g2_decap_8 FILLER_79_3364 ();
 sg13g2_decap_8 FILLER_79_3371 ();
 sg13g2_decap_8 FILLER_79_3378 ();
 sg13g2_decap_8 FILLER_79_3385 ();
 sg13g2_decap_8 FILLER_79_3392 ();
 sg13g2_decap_8 FILLER_79_3399 ();
 sg13g2_decap_8 FILLER_79_3406 ();
 sg13g2_decap_8 FILLER_79_3413 ();
 sg13g2_decap_8 FILLER_79_3420 ();
 sg13g2_decap_8 FILLER_79_3427 ();
 sg13g2_decap_8 FILLER_79_3434 ();
 sg13g2_decap_8 FILLER_79_3441 ();
 sg13g2_decap_8 FILLER_79_3448 ();
 sg13g2_decap_8 FILLER_79_3455 ();
 sg13g2_decap_8 FILLER_79_3462 ();
 sg13g2_decap_8 FILLER_79_3469 ();
 sg13g2_decap_8 FILLER_79_3476 ();
 sg13g2_decap_8 FILLER_79_3483 ();
 sg13g2_decap_8 FILLER_79_3490 ();
 sg13g2_decap_8 FILLER_79_3497 ();
 sg13g2_decap_8 FILLER_79_3504 ();
 sg13g2_decap_8 FILLER_79_3511 ();
 sg13g2_decap_8 FILLER_79_3518 ();
 sg13g2_decap_8 FILLER_79_3525 ();
 sg13g2_decap_8 FILLER_79_3532 ();
 sg13g2_decap_8 FILLER_79_3539 ();
 sg13g2_decap_8 FILLER_79_3546 ();
 sg13g2_decap_8 FILLER_79_3553 ();
 sg13g2_decap_8 FILLER_79_3560 ();
 sg13g2_decap_8 FILLER_79_3567 ();
 sg13g2_decap_4 FILLER_79_3574 ();
 sg13g2_fill_2 FILLER_79_3578 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_42 ();
 sg13g2_decap_8 FILLER_80_49 ();
 sg13g2_decap_4 FILLER_80_60 ();
 sg13g2_decap_4 FILLER_80_68 ();
 sg13g2_decap_4 FILLER_80_76 ();
 sg13g2_decap_4 FILLER_80_84 ();
 sg13g2_decap_4 FILLER_80_92 ();
 sg13g2_decap_4 FILLER_80_100 ();
 sg13g2_decap_4 FILLER_80_108 ();
 sg13g2_decap_8 FILLER_80_116 ();
 sg13g2_decap_4 FILLER_80_123 ();
 sg13g2_fill_1 FILLER_80_127 ();
 sg13g2_decap_8 FILLER_80_132 ();
 sg13g2_decap_4 FILLER_80_139 ();
 sg13g2_decap_4 FILLER_80_172 ();
 sg13g2_decap_8 FILLER_80_180 ();
 sg13g2_decap_8 FILLER_80_187 ();
 sg13g2_decap_8 FILLER_80_194 ();
 sg13g2_decap_8 FILLER_80_201 ();
 sg13g2_decap_8 FILLER_80_208 ();
 sg13g2_decap_8 FILLER_80_215 ();
 sg13g2_decap_8 FILLER_80_222 ();
 sg13g2_decap_8 FILLER_80_229 ();
 sg13g2_decap_8 FILLER_80_236 ();
 sg13g2_decap_8 FILLER_80_243 ();
 sg13g2_decap_4 FILLER_80_250 ();
 sg13g2_fill_2 FILLER_80_254 ();
 sg13g2_decap_8 FILLER_80_264 ();
 sg13g2_fill_1 FILLER_80_271 ();
 sg13g2_decap_8 FILLER_80_280 ();
 sg13g2_fill_1 FILLER_80_287 ();
 sg13g2_fill_1 FILLER_80_296 ();
 sg13g2_decap_4 FILLER_80_349 ();
 sg13g2_fill_2 FILLER_80_353 ();
 sg13g2_decap_8 FILLER_80_386 ();
 sg13g2_decap_8 FILLER_80_393 ();
 sg13g2_decap_8 FILLER_80_400 ();
 sg13g2_decap_8 FILLER_80_407 ();
 sg13g2_decap_8 FILLER_80_414 ();
 sg13g2_decap_8 FILLER_80_421 ();
 sg13g2_decap_8 FILLER_80_428 ();
 sg13g2_decap_8 FILLER_80_435 ();
 sg13g2_decap_8 FILLER_80_442 ();
 sg13g2_decap_8 FILLER_80_449 ();
 sg13g2_decap_8 FILLER_80_456 ();
 sg13g2_decap_8 FILLER_80_463 ();
 sg13g2_decap_8 FILLER_80_470 ();
 sg13g2_decap_8 FILLER_80_477 ();
 sg13g2_decap_8 FILLER_80_484 ();
 sg13g2_decap_8 FILLER_80_491 ();
 sg13g2_decap_8 FILLER_80_498 ();
 sg13g2_decap_8 FILLER_80_505 ();
 sg13g2_decap_8 FILLER_80_512 ();
 sg13g2_decap_8 FILLER_80_519 ();
 sg13g2_decap_8 FILLER_80_526 ();
 sg13g2_decap_8 FILLER_80_533 ();
 sg13g2_decap_8 FILLER_80_540 ();
 sg13g2_decap_8 FILLER_80_547 ();
 sg13g2_decap_8 FILLER_80_554 ();
 sg13g2_decap_8 FILLER_80_561 ();
 sg13g2_decap_8 FILLER_80_568 ();
 sg13g2_decap_8 FILLER_80_575 ();
 sg13g2_decap_8 FILLER_80_582 ();
 sg13g2_fill_2 FILLER_80_589 ();
 sg13g2_decap_8 FILLER_80_595 ();
 sg13g2_decap_8 FILLER_80_602 ();
 sg13g2_decap_8 FILLER_80_609 ();
 sg13g2_decap_8 FILLER_80_616 ();
 sg13g2_decap_8 FILLER_80_623 ();
 sg13g2_decap_8 FILLER_80_630 ();
 sg13g2_decap_8 FILLER_80_637 ();
 sg13g2_decap_4 FILLER_80_644 ();
 sg13g2_decap_8 FILLER_80_657 ();
 sg13g2_decap_8 FILLER_80_664 ();
 sg13g2_decap_8 FILLER_80_671 ();
 sg13g2_decap_8 FILLER_80_678 ();
 sg13g2_decap_8 FILLER_80_685 ();
 sg13g2_decap_8 FILLER_80_692 ();
 sg13g2_decap_8 FILLER_80_699 ();
 sg13g2_decap_8 FILLER_80_706 ();
 sg13g2_decap_8 FILLER_80_713 ();
 sg13g2_decap_8 FILLER_80_727 ();
 sg13g2_decap_8 FILLER_80_734 ();
 sg13g2_decap_8 FILLER_80_741 ();
 sg13g2_decap_8 FILLER_80_748 ();
 sg13g2_decap_8 FILLER_80_755 ();
 sg13g2_decap_8 FILLER_80_762 ();
 sg13g2_decap_8 FILLER_80_769 ();
 sg13g2_decap_8 FILLER_80_776 ();
 sg13g2_decap_8 FILLER_80_783 ();
 sg13g2_decap_8 FILLER_80_790 ();
 sg13g2_decap_8 FILLER_80_797 ();
 sg13g2_decap_8 FILLER_80_804 ();
 sg13g2_decap_8 FILLER_80_811 ();
 sg13g2_decap_8 FILLER_80_818 ();
 sg13g2_decap_8 FILLER_80_825 ();
 sg13g2_decap_8 FILLER_80_832 ();
 sg13g2_decap_8 FILLER_80_839 ();
 sg13g2_decap_8 FILLER_80_846 ();
 sg13g2_decap_8 FILLER_80_853 ();
 sg13g2_decap_8 FILLER_80_860 ();
 sg13g2_decap_8 FILLER_80_867 ();
 sg13g2_decap_8 FILLER_80_874 ();
 sg13g2_decap_8 FILLER_80_881 ();
 sg13g2_decap_8 FILLER_80_888 ();
 sg13g2_decap_8 FILLER_80_895 ();
 sg13g2_decap_8 FILLER_80_902 ();
 sg13g2_decap_8 FILLER_80_909 ();
 sg13g2_decap_8 FILLER_80_916 ();
 sg13g2_decap_4 FILLER_80_923 ();
 sg13g2_decap_8 FILLER_80_932 ();
 sg13g2_decap_8 FILLER_80_939 ();
 sg13g2_decap_8 FILLER_80_946 ();
 sg13g2_decap_8 FILLER_80_953 ();
 sg13g2_decap_8 FILLER_80_960 ();
 sg13g2_decap_8 FILLER_80_967 ();
 sg13g2_decap_8 FILLER_80_974 ();
 sg13g2_decap_8 FILLER_80_981 ();
 sg13g2_decap_8 FILLER_80_988 ();
 sg13g2_decap_8 FILLER_80_995 ();
 sg13g2_decap_4 FILLER_80_1002 ();
 sg13g2_fill_2 FILLER_80_1006 ();
 sg13g2_decap_8 FILLER_80_1027 ();
 sg13g2_decap_8 FILLER_80_1034 ();
 sg13g2_decap_8 FILLER_80_1041 ();
 sg13g2_decap_8 FILLER_80_1048 ();
 sg13g2_fill_2 FILLER_80_1055 ();
 sg13g2_fill_1 FILLER_80_1057 ();
 sg13g2_decap_8 FILLER_80_1067 ();
 sg13g2_decap_8 FILLER_80_1074 ();
 sg13g2_decap_8 FILLER_80_1081 ();
 sg13g2_decap_8 FILLER_80_1088 ();
 sg13g2_decap_8 FILLER_80_1095 ();
 sg13g2_decap_8 FILLER_80_1102 ();
 sg13g2_decap_8 FILLER_80_1109 ();
 sg13g2_decap_8 FILLER_80_1116 ();
 sg13g2_decap_4 FILLER_80_1123 ();
 sg13g2_fill_1 FILLER_80_1127 ();
 sg13g2_decap_8 FILLER_80_1137 ();
 sg13g2_decap_8 FILLER_80_1144 ();
 sg13g2_decap_8 FILLER_80_1151 ();
 sg13g2_decap_8 FILLER_80_1158 ();
 sg13g2_decap_8 FILLER_80_1165 ();
 sg13g2_decap_8 FILLER_80_1172 ();
 sg13g2_decap_8 FILLER_80_1179 ();
 sg13g2_fill_2 FILLER_80_1186 ();
 sg13g2_decap_8 FILLER_80_1197 ();
 sg13g2_decap_8 FILLER_80_1204 ();
 sg13g2_decap_8 FILLER_80_1211 ();
 sg13g2_decap_8 FILLER_80_1218 ();
 sg13g2_decap_8 FILLER_80_1225 ();
 sg13g2_decap_8 FILLER_80_1232 ();
 sg13g2_decap_8 FILLER_80_1239 ();
 sg13g2_decap_8 FILLER_80_1246 ();
 sg13g2_decap_8 FILLER_80_1253 ();
 sg13g2_decap_8 FILLER_80_1260 ();
 sg13g2_decap_4 FILLER_80_1267 ();
 sg13g2_fill_1 FILLER_80_1271 ();
 sg13g2_decap_8 FILLER_80_1281 ();
 sg13g2_decap_8 FILLER_80_1288 ();
 sg13g2_decap_8 FILLER_80_1295 ();
 sg13g2_decap_8 FILLER_80_1302 ();
 sg13g2_decap_8 FILLER_80_1309 ();
 sg13g2_decap_8 FILLER_80_1316 ();
 sg13g2_decap_8 FILLER_80_1323 ();
 sg13g2_decap_8 FILLER_80_1330 ();
 sg13g2_decap_8 FILLER_80_1337 ();
 sg13g2_decap_8 FILLER_80_1344 ();
 sg13g2_decap_8 FILLER_80_1351 ();
 sg13g2_decap_8 FILLER_80_1358 ();
 sg13g2_decap_8 FILLER_80_1365 ();
 sg13g2_decap_8 FILLER_80_1372 ();
 sg13g2_fill_2 FILLER_80_1379 ();
 sg13g2_decap_8 FILLER_80_1386 ();
 sg13g2_decap_8 FILLER_80_1393 ();
 sg13g2_decap_8 FILLER_80_1400 ();
 sg13g2_decap_8 FILLER_80_1407 ();
 sg13g2_decap_8 FILLER_80_1414 ();
 sg13g2_decap_8 FILLER_80_1421 ();
 sg13g2_decap_8 FILLER_80_1428 ();
 sg13g2_decap_8 FILLER_80_1435 ();
 sg13g2_decap_8 FILLER_80_1442 ();
 sg13g2_decap_8 FILLER_80_1449 ();
 sg13g2_decap_8 FILLER_80_1456 ();
 sg13g2_decap_8 FILLER_80_1463 ();
 sg13g2_decap_8 FILLER_80_1470 ();
 sg13g2_decap_8 FILLER_80_1477 ();
 sg13g2_decap_8 FILLER_80_1484 ();
 sg13g2_decap_8 FILLER_80_1491 ();
 sg13g2_decap_8 FILLER_80_1498 ();
 sg13g2_decap_8 FILLER_80_1505 ();
 sg13g2_decap_8 FILLER_80_1512 ();
 sg13g2_fill_1 FILLER_80_1519 ();
 sg13g2_fill_2 FILLER_80_1525 ();
 sg13g2_decap_8 FILLER_80_1533 ();
 sg13g2_decap_8 FILLER_80_1540 ();
 sg13g2_decap_8 FILLER_80_1547 ();
 sg13g2_decap_8 FILLER_80_1554 ();
 sg13g2_decap_8 FILLER_80_1561 ();
 sg13g2_decap_8 FILLER_80_1568 ();
 sg13g2_decap_8 FILLER_80_1575 ();
 sg13g2_decap_8 FILLER_80_1582 ();
 sg13g2_decap_8 FILLER_80_1589 ();
 sg13g2_decap_8 FILLER_80_1596 ();
 sg13g2_decap_8 FILLER_80_1603 ();
 sg13g2_decap_8 FILLER_80_1610 ();
 sg13g2_decap_8 FILLER_80_1617 ();
 sg13g2_decap_8 FILLER_80_1624 ();
 sg13g2_decap_8 FILLER_80_1631 ();
 sg13g2_decap_8 FILLER_80_1638 ();
 sg13g2_decap_8 FILLER_80_1645 ();
 sg13g2_decap_8 FILLER_80_1652 ();
 sg13g2_decap_8 FILLER_80_1659 ();
 sg13g2_decap_8 FILLER_80_1666 ();
 sg13g2_decap_8 FILLER_80_1673 ();
 sg13g2_decap_8 FILLER_80_1680 ();
 sg13g2_decap_8 FILLER_80_1687 ();
 sg13g2_decap_8 FILLER_80_1694 ();
 sg13g2_decap_8 FILLER_80_1701 ();
 sg13g2_decap_8 FILLER_80_1708 ();
 sg13g2_decap_8 FILLER_80_1715 ();
 sg13g2_decap_8 FILLER_80_1722 ();
 sg13g2_decap_8 FILLER_80_1729 ();
 sg13g2_decap_8 FILLER_80_1736 ();
 sg13g2_decap_8 FILLER_80_1743 ();
 sg13g2_decap_8 FILLER_80_1750 ();
 sg13g2_decap_8 FILLER_80_1757 ();
 sg13g2_decap_8 FILLER_80_1764 ();
 sg13g2_decap_8 FILLER_80_1771 ();
 sg13g2_decap_8 FILLER_80_1778 ();
 sg13g2_decap_8 FILLER_80_1785 ();
 sg13g2_decap_8 FILLER_80_1792 ();
 sg13g2_decap_8 FILLER_80_1799 ();
 sg13g2_decap_8 FILLER_80_1806 ();
 sg13g2_decap_8 FILLER_80_1813 ();
 sg13g2_decap_8 FILLER_80_1820 ();
 sg13g2_decap_8 FILLER_80_1827 ();
 sg13g2_decap_8 FILLER_80_1834 ();
 sg13g2_decap_8 FILLER_80_1841 ();
 sg13g2_decap_8 FILLER_80_1848 ();
 sg13g2_decap_8 FILLER_80_1855 ();
 sg13g2_decap_8 FILLER_80_1862 ();
 sg13g2_decap_8 FILLER_80_1869 ();
 sg13g2_decap_8 FILLER_80_1876 ();
 sg13g2_decap_8 FILLER_80_1883 ();
 sg13g2_decap_8 FILLER_80_1890 ();
 sg13g2_decap_8 FILLER_80_1897 ();
 sg13g2_decap_8 FILLER_80_1904 ();
 sg13g2_decap_8 FILLER_80_1911 ();
 sg13g2_decap_8 FILLER_80_1918 ();
 sg13g2_decap_8 FILLER_80_1925 ();
 sg13g2_decap_8 FILLER_80_1932 ();
 sg13g2_decap_8 FILLER_80_1939 ();
 sg13g2_decap_8 FILLER_80_1946 ();
 sg13g2_decap_8 FILLER_80_1953 ();
 sg13g2_decap_8 FILLER_80_1960 ();
 sg13g2_decap_8 FILLER_80_1967 ();
 sg13g2_decap_8 FILLER_80_1974 ();
 sg13g2_decap_8 FILLER_80_1981 ();
 sg13g2_decap_8 FILLER_80_1988 ();
 sg13g2_decap_8 FILLER_80_1995 ();
 sg13g2_decap_8 FILLER_80_2002 ();
 sg13g2_decap_8 FILLER_80_2009 ();
 sg13g2_decap_8 FILLER_80_2016 ();
 sg13g2_decap_8 FILLER_80_2023 ();
 sg13g2_decap_8 FILLER_80_2030 ();
 sg13g2_decap_8 FILLER_80_2037 ();
 sg13g2_decap_8 FILLER_80_2044 ();
 sg13g2_decap_8 FILLER_80_2051 ();
 sg13g2_decap_8 FILLER_80_2058 ();
 sg13g2_decap_8 FILLER_80_2065 ();
 sg13g2_decap_8 FILLER_80_2072 ();
 sg13g2_decap_8 FILLER_80_2079 ();
 sg13g2_decap_8 FILLER_80_2086 ();
 sg13g2_decap_8 FILLER_80_2093 ();
 sg13g2_decap_8 FILLER_80_2100 ();
 sg13g2_decap_8 FILLER_80_2107 ();
 sg13g2_decap_8 FILLER_80_2114 ();
 sg13g2_decap_8 FILLER_80_2121 ();
 sg13g2_decap_8 FILLER_80_2128 ();
 sg13g2_decap_8 FILLER_80_2135 ();
 sg13g2_decap_8 FILLER_80_2142 ();
 sg13g2_decap_8 FILLER_80_2149 ();
 sg13g2_decap_8 FILLER_80_2156 ();
 sg13g2_decap_8 FILLER_80_2163 ();
 sg13g2_decap_8 FILLER_80_2170 ();
 sg13g2_decap_8 FILLER_80_2177 ();
 sg13g2_decap_8 FILLER_80_2184 ();
 sg13g2_decap_8 FILLER_80_2191 ();
 sg13g2_decap_8 FILLER_80_2198 ();
 sg13g2_decap_8 FILLER_80_2205 ();
 sg13g2_decap_8 FILLER_80_2212 ();
 sg13g2_decap_8 FILLER_80_2219 ();
 sg13g2_decap_8 FILLER_80_2226 ();
 sg13g2_decap_8 FILLER_80_2233 ();
 sg13g2_decap_8 FILLER_80_2240 ();
 sg13g2_decap_4 FILLER_80_2247 ();
 sg13g2_fill_1 FILLER_80_2251 ();
 sg13g2_decap_8 FILLER_80_2261 ();
 sg13g2_decap_8 FILLER_80_2268 ();
 sg13g2_decap_8 FILLER_80_2275 ();
 sg13g2_decap_8 FILLER_80_2282 ();
 sg13g2_decap_8 FILLER_80_2289 ();
 sg13g2_decap_4 FILLER_80_2296 ();
 sg13g2_fill_2 FILLER_80_2300 ();
 sg13g2_decap_8 FILLER_80_2311 ();
 sg13g2_decap_8 FILLER_80_2318 ();
 sg13g2_decap_8 FILLER_80_2325 ();
 sg13g2_decap_8 FILLER_80_2332 ();
 sg13g2_fill_2 FILLER_80_2339 ();
 sg13g2_fill_1 FILLER_80_2341 ();
 sg13g2_decap_8 FILLER_80_2347 ();
 sg13g2_decap_8 FILLER_80_2354 ();
 sg13g2_decap_8 FILLER_80_2361 ();
 sg13g2_decap_8 FILLER_80_2368 ();
 sg13g2_decap_8 FILLER_80_2375 ();
 sg13g2_decap_8 FILLER_80_2382 ();
 sg13g2_decap_8 FILLER_80_2389 ();
 sg13g2_decap_8 FILLER_80_2396 ();
 sg13g2_decap_8 FILLER_80_2403 ();
 sg13g2_decap_8 FILLER_80_2410 ();
 sg13g2_decap_8 FILLER_80_2417 ();
 sg13g2_decap_8 FILLER_80_2424 ();
 sg13g2_decap_8 FILLER_80_2431 ();
 sg13g2_decap_8 FILLER_80_2438 ();
 sg13g2_decap_4 FILLER_80_2445 ();
 sg13g2_decap_8 FILLER_80_2458 ();
 sg13g2_decap_8 FILLER_80_2465 ();
 sg13g2_decap_8 FILLER_80_2472 ();
 sg13g2_decap_8 FILLER_80_2479 ();
 sg13g2_decap_8 FILLER_80_2486 ();
 sg13g2_decap_8 FILLER_80_2493 ();
 sg13g2_decap_8 FILLER_80_2500 ();
 sg13g2_decap_8 FILLER_80_2507 ();
 sg13g2_decap_8 FILLER_80_2514 ();
 sg13g2_decap_8 FILLER_80_2521 ();
 sg13g2_decap_8 FILLER_80_2528 ();
 sg13g2_decap_8 FILLER_80_2535 ();
 sg13g2_decap_8 FILLER_80_2542 ();
 sg13g2_decap_8 FILLER_80_2549 ();
 sg13g2_decap_8 FILLER_80_2556 ();
 sg13g2_decap_8 FILLER_80_2563 ();
 sg13g2_decap_8 FILLER_80_2570 ();
 sg13g2_decap_8 FILLER_80_2577 ();
 sg13g2_decap_8 FILLER_80_2584 ();
 sg13g2_decap_8 FILLER_80_2591 ();
 sg13g2_decap_8 FILLER_80_2598 ();
 sg13g2_decap_8 FILLER_80_2605 ();
 sg13g2_decap_8 FILLER_80_2612 ();
 sg13g2_decap_8 FILLER_80_2619 ();
 sg13g2_decap_8 FILLER_80_2626 ();
 sg13g2_decap_8 FILLER_80_2633 ();
 sg13g2_decap_8 FILLER_80_2640 ();
 sg13g2_decap_8 FILLER_80_2647 ();
 sg13g2_decap_8 FILLER_80_2654 ();
 sg13g2_fill_2 FILLER_80_2661 ();
 sg13g2_fill_1 FILLER_80_2663 ();
 sg13g2_decap_8 FILLER_80_2673 ();
 sg13g2_decap_4 FILLER_80_2680 ();
 sg13g2_fill_2 FILLER_80_2684 ();
 sg13g2_decap_8 FILLER_80_2695 ();
 sg13g2_decap_8 FILLER_80_2702 ();
 sg13g2_decap_8 FILLER_80_2709 ();
 sg13g2_decap_8 FILLER_80_2716 ();
 sg13g2_decap_8 FILLER_80_2723 ();
 sg13g2_decap_8 FILLER_80_2730 ();
 sg13g2_decap_8 FILLER_80_2737 ();
 sg13g2_decap_8 FILLER_80_2744 ();
 sg13g2_decap_8 FILLER_80_2751 ();
 sg13g2_decap_8 FILLER_80_2758 ();
 sg13g2_decap_8 FILLER_80_2765 ();
 sg13g2_decap_8 FILLER_80_2772 ();
 sg13g2_decap_8 FILLER_80_2779 ();
 sg13g2_decap_8 FILLER_80_2786 ();
 sg13g2_decap_8 FILLER_80_2793 ();
 sg13g2_decap_8 FILLER_80_2800 ();
 sg13g2_decap_8 FILLER_80_2807 ();
 sg13g2_decap_4 FILLER_80_2814 ();
 sg13g2_decap_8 FILLER_80_2827 ();
 sg13g2_decap_8 FILLER_80_2834 ();
 sg13g2_decap_8 FILLER_80_2841 ();
 sg13g2_decap_8 FILLER_80_2848 ();
 sg13g2_decap_8 FILLER_80_2855 ();
 sg13g2_decap_8 FILLER_80_2862 ();
 sg13g2_decap_8 FILLER_80_2869 ();
 sg13g2_decap_8 FILLER_80_2876 ();
 sg13g2_decap_8 FILLER_80_2883 ();
 sg13g2_decap_8 FILLER_80_2890 ();
 sg13g2_decap_8 FILLER_80_2897 ();
 sg13g2_decap_8 FILLER_80_2904 ();
 sg13g2_decap_8 FILLER_80_2911 ();
 sg13g2_decap_8 FILLER_80_2918 ();
 sg13g2_decap_8 FILLER_80_2925 ();
 sg13g2_decap_8 FILLER_80_2932 ();
 sg13g2_decap_8 FILLER_80_2939 ();
 sg13g2_decap_8 FILLER_80_2946 ();
 sg13g2_decap_8 FILLER_80_2953 ();
 sg13g2_decap_8 FILLER_80_2960 ();
 sg13g2_decap_8 FILLER_80_2967 ();
 sg13g2_decap_8 FILLER_80_2974 ();
 sg13g2_decap_8 FILLER_80_2981 ();
 sg13g2_fill_2 FILLER_80_2988 ();
 sg13g2_fill_1 FILLER_80_2990 ();
 sg13g2_fill_2 FILLER_80_3000 ();
 sg13g2_fill_1 FILLER_80_3002 ();
 sg13g2_decap_8 FILLER_80_3012 ();
 sg13g2_decap_8 FILLER_80_3019 ();
 sg13g2_decap_8 FILLER_80_3026 ();
 sg13g2_decap_8 FILLER_80_3033 ();
 sg13g2_decap_8 FILLER_80_3040 ();
 sg13g2_decap_8 FILLER_80_3047 ();
 sg13g2_decap_8 FILLER_80_3054 ();
 sg13g2_decap_8 FILLER_80_3061 ();
 sg13g2_decap_8 FILLER_80_3068 ();
 sg13g2_decap_8 FILLER_80_3075 ();
 sg13g2_decap_8 FILLER_80_3082 ();
 sg13g2_decap_8 FILLER_80_3089 ();
 sg13g2_decap_8 FILLER_80_3096 ();
 sg13g2_decap_8 FILLER_80_3103 ();
 sg13g2_decap_8 FILLER_80_3110 ();
 sg13g2_decap_8 FILLER_80_3117 ();
 sg13g2_decap_8 FILLER_80_3124 ();
 sg13g2_decap_8 FILLER_80_3131 ();
 sg13g2_decap_8 FILLER_80_3138 ();
 sg13g2_decap_8 FILLER_80_3145 ();
 sg13g2_decap_8 FILLER_80_3161 ();
 sg13g2_decap_8 FILLER_80_3168 ();
 sg13g2_decap_8 FILLER_80_3175 ();
 sg13g2_decap_8 FILLER_80_3182 ();
 sg13g2_decap_8 FILLER_80_3189 ();
 sg13g2_fill_2 FILLER_80_3196 ();
 sg13g2_decap_8 FILLER_80_3207 ();
 sg13g2_decap_8 FILLER_80_3214 ();
 sg13g2_decap_8 FILLER_80_3221 ();
 sg13g2_decap_8 FILLER_80_3228 ();
 sg13g2_fill_2 FILLER_80_3235 ();
 sg13g2_fill_1 FILLER_80_3237 ();
 sg13g2_decap_8 FILLER_80_3247 ();
 sg13g2_decap_8 FILLER_80_3254 ();
 sg13g2_decap_8 FILLER_80_3261 ();
 sg13g2_decap_8 FILLER_80_3268 ();
 sg13g2_decap_8 FILLER_80_3275 ();
 sg13g2_decap_8 FILLER_80_3282 ();
 sg13g2_decap_4 FILLER_80_3289 ();
 sg13g2_decap_8 FILLER_80_3302 ();
 sg13g2_decap_8 FILLER_80_3309 ();
 sg13g2_decap_8 FILLER_80_3316 ();
 sg13g2_decap_8 FILLER_80_3323 ();
 sg13g2_decap_8 FILLER_80_3330 ();
 sg13g2_decap_8 FILLER_80_3337 ();
 sg13g2_decap_8 FILLER_80_3344 ();
 sg13g2_decap_8 FILLER_80_3351 ();
 sg13g2_decap_8 FILLER_80_3358 ();
 sg13g2_decap_8 FILLER_80_3365 ();
 sg13g2_decap_8 FILLER_80_3372 ();
 sg13g2_decap_8 FILLER_80_3379 ();
 sg13g2_decap_8 FILLER_80_3386 ();
 sg13g2_decap_8 FILLER_80_3393 ();
 sg13g2_decap_8 FILLER_80_3400 ();
 sg13g2_decap_8 FILLER_80_3407 ();
 sg13g2_decap_8 FILLER_80_3414 ();
 sg13g2_decap_8 FILLER_80_3421 ();
 sg13g2_decap_8 FILLER_80_3428 ();
 sg13g2_decap_8 FILLER_80_3435 ();
 sg13g2_decap_8 FILLER_80_3442 ();
 sg13g2_decap_8 FILLER_80_3449 ();
 sg13g2_decap_8 FILLER_80_3456 ();
 sg13g2_decap_8 FILLER_80_3463 ();
 sg13g2_decap_8 FILLER_80_3470 ();
 sg13g2_decap_8 FILLER_80_3477 ();
 sg13g2_decap_8 FILLER_80_3484 ();
 sg13g2_decap_8 FILLER_80_3491 ();
 sg13g2_decap_8 FILLER_80_3498 ();
 sg13g2_decap_8 FILLER_80_3505 ();
 sg13g2_decap_8 FILLER_80_3512 ();
 sg13g2_decap_8 FILLER_80_3519 ();
 sg13g2_decap_8 FILLER_80_3526 ();
 sg13g2_decap_8 FILLER_80_3533 ();
 sg13g2_decap_8 FILLER_80_3540 ();
 sg13g2_decap_8 FILLER_80_3547 ();
 sg13g2_decap_8 FILLER_80_3554 ();
 sg13g2_decap_8 FILLER_80_3561 ();
 sg13g2_decap_8 FILLER_80_3568 ();
 sg13g2_decap_4 FILLER_80_3575 ();
 sg13g2_fill_1 FILLER_80_3579 ();
 assign uio_oe[0] = net16;
 assign uio_oe[1] = net17;
 assign uio_oe[2] = net28;
 assign uio_oe[3] = net18;
 assign uio_oe[4] = net19;
 assign uio_oe[5] = net29;
 assign uio_oe[6] = net20;
 assign uio_oe[7] = net30;
 assign uio_out[0] = net21;
 assign uio_out[1] = net22;
 assign uio_out[3] = net23;
 assign uio_out[4] = net24;
 assign uio_out[6] = net25;
endmodule

module tt_um_bytex64_munch (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire \atick_clock[0] ;
 wire \atick_clock[1] ;
 wire audio;
 wire \audio_mod.audio_gen.ch0_state ;
 wire \audio_mod.audio_gen.ch1_state ;
 wire \audio_mod.audio_gen.ch2_state ;
 wire \audio_mod.audio_gen.ch3_state ;
 wire \audio_mod.audio_gen.chan0.ch_counter[0] ;
 wire \audio_mod.audio_gen.chan0.ch_counter[10] ;
 wire \audio_mod.audio_gen.chan0.ch_counter[11] ;
 wire \audio_mod.audio_gen.chan0.ch_counter[1] ;
 wire \audio_mod.audio_gen.chan0.ch_counter[2] ;
 wire \audio_mod.audio_gen.chan0.ch_counter[3] ;
 wire \audio_mod.audio_gen.chan0.ch_counter[4] ;
 wire \audio_mod.audio_gen.chan0.ch_counter[5] ;
 wire \audio_mod.audio_gen.chan0.ch_counter[6] ;
 wire \audio_mod.audio_gen.chan0.ch_counter[7] ;
 wire \audio_mod.audio_gen.chan0.ch_counter[8] ;
 wire \audio_mod.audio_gen.chan0.ch_counter[9] ;
 wire \audio_mod.audio_gen.chan1.ch_counter[0] ;
 wire \audio_mod.audio_gen.chan1.ch_counter[10] ;
 wire \audio_mod.audio_gen.chan1.ch_counter[11] ;
 wire \audio_mod.audio_gen.chan1.ch_counter[1] ;
 wire \audio_mod.audio_gen.chan1.ch_counter[2] ;
 wire \audio_mod.audio_gen.chan1.ch_counter[3] ;
 wire \audio_mod.audio_gen.chan1.ch_counter[4] ;
 wire \audio_mod.audio_gen.chan1.ch_counter[5] ;
 wire \audio_mod.audio_gen.chan1.ch_counter[6] ;
 wire \audio_mod.audio_gen.chan1.ch_counter[7] ;
 wire \audio_mod.audio_gen.chan1.ch_counter[8] ;
 wire \audio_mod.audio_gen.chan1.ch_counter[9] ;
 wire \audio_mod.audio_gen.chan2.ch_counter[0] ;
 wire \audio_mod.audio_gen.chan2.ch_counter[10] ;
 wire \audio_mod.audio_gen.chan2.ch_counter[11] ;
 wire \audio_mod.audio_gen.chan2.ch_counter[1] ;
 wire \audio_mod.audio_gen.chan2.ch_counter[2] ;
 wire \audio_mod.audio_gen.chan2.ch_counter[3] ;
 wire \audio_mod.audio_gen.chan2.ch_counter[4] ;
 wire \audio_mod.audio_gen.chan2.ch_counter[5] ;
 wire \audio_mod.audio_gen.chan2.ch_counter[6] ;
 wire \audio_mod.audio_gen.chan2.ch_counter[7] ;
 wire \audio_mod.audio_gen.chan2.ch_counter[8] ;
 wire \audio_mod.audio_gen.chan2.ch_counter[9] ;
 wire \audio_mod.audio_gen.chan3.ch_counter[0] ;
 wire \audio_mod.audio_gen.chan3.ch_counter[10] ;
 wire \audio_mod.audio_gen.chan3.ch_counter[11] ;
 wire \audio_mod.audio_gen.chan3.ch_counter[1] ;
 wire \audio_mod.audio_gen.chan3.ch_counter[2] ;
 wire \audio_mod.audio_gen.chan3.ch_counter[3] ;
 wire \audio_mod.audio_gen.chan3.ch_counter[4] ;
 wire \audio_mod.audio_gen.chan3.ch_counter[5] ;
 wire \audio_mod.audio_gen.chan3.ch_counter[6] ;
 wire \audio_mod.audio_gen.chan3.ch_counter[7] ;
 wire \audio_mod.audio_gen.chan3.ch_counter[8] ;
 wire \audio_mod.audio_gen.chan3.ch_counter[9] ;
 wire \audio_mod.audio_gen.chan3.rng ;
 wire \audio_mod.audio_gen.pwm_clock[0] ;
 wire \audio_mod.audio_gen.pwm_clock[1] ;
 wire \audio_mod.audio_gen.pwm_clock[2] ;
 wire \audio_mod.audio_gen.pwm_clock[3] ;
 wire \audio_mod.audio_gen.pwm_clock[4] ;
 wire \audio_mod.audio_gen.pwm_clock[5] ;
 wire \audio_mod.pattern_clock[0] ;
 wire \audio_mod.pattern_clock[1] ;
 wire \audio_mod.pattern_clock[2] ;
 wire \audio_mod.pattern_clock[3] ;
 wire \audio_mod.seq.seq_clock[0] ;
 wire \audio_mod.seq.seq_clock[1] ;
 wire \audio_mod.seq.seq_clock[2] ;
 wire \audio_mod.seq.seq_clock[3] ;
 wire \background_color[0] ;
 wire \background_color[1] ;
 wire \background_color[2] ;
 wire \bright[2][0] ;
 wire \clock_gen.r_atick_clock[0] ;
 wire \clock_gen.vsync ;
 wire \counter[0] ;
 wire \counter[1] ;
 wire \counter[2] ;
 wire \counter[3] ;
 wire \counter[4] ;
 wire \counter[5] ;
 wire \counter[6] ;
 wire \hpos[0] ;
 wire \hpos[1] ;
 wire \hpos[2] ;
 wire \hpos[3] ;
 wire \hpos[4] ;
 wire \hpos[5] ;
 wire \hpos[6] ;
 wire \hpos[7] ;
 wire \hpos[8] ;
 wire \hpos[9] ;
 wire hsync;
 wire \hvsync_gen.vpos[0] ;
 wire \hvsync_gen.vpos[1] ;
 wire \hvsync_gen.vpos[2] ;
 wire \hvsync_gen.vpos[3] ;
 wire \hvsync_gen.vpos[4] ;
 wire \hvsync_gen.vpos[5] ;
 wire \hvsync_gen.vpos[6] ;
 wire \hvsync_gen.vpos[7] ;
 wire \hvsync_gen.vpos[8] ;
 wire \hvsync_gen.vpos[9] ;
 wire \lfsr[1] ;
 wire \lfsr[2] ;
 wire \lfsr[4] ;
 wire \lfsr[5] ;
 wire \lfsr_dev.lfsr[10] ;
 wire \lfsr_dev.lfsr[6] ;
 wire \lfsr_dev.lfsr[7] ;
 wire \lfsr_dev.lfsr[8] ;
 wire \lfsr_dev.lfsr[9] ;
 wire \stage[0] ;
 wire \stage[1] ;
 wire \stage_seq_inst.stage_timer[0] ;
 wire \stage_seq_inst.stage_timer[1] ;
 wire \stage_seq_inst.stage_timer[2] ;
 wire \stage_seq_inst.stage_timer[3] ;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net32;
 wire net33;
 wire net34;
 wire clknet_0_clk;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net1;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;

 sg13g2_inv_2 _1142_ (.Y(_0372_),
    .A(net289));
 sg13g2_inv_1 _1143_ (.Y(_0373_),
    .A(\audio_mod.seq.seq_clock[3] ));
 sg13g2_inv_1 _1144_ (.Y(_0374_),
    .A(\audio_mod.seq.seq_clock[1] ));
 sg13g2_inv_1 _1145_ (.Y(_0051_),
    .A(\audio_mod.seq.seq_clock[0] ));
 sg13g2_inv_1 _1146_ (.Y(_0375_),
    .A(\audio_mod.audio_gen.pwm_clock[1] ));
 sg13g2_inv_1 _1147_ (.Y(_0376_),
    .A(net54));
 sg13g2_inv_1 _1148_ (.Y(_0377_),
    .A(\audio_mod.audio_gen.chan0.ch_counter[7] ));
 sg13g2_inv_1 _1149_ (.Y(_0378_),
    .A(\audio_mod.audio_gen.chan1.ch_counter[7] ));
 sg13g2_inv_1 _1150_ (.Y(_0379_),
    .A(\audio_mod.audio_gen.chan2.ch_counter[7] ));
 sg13g2_inv_1 _1151_ (.Y(_0380_),
    .A(_0074_));
 sg13g2_inv_1 _1152_ (.Y(_0055_),
    .A(net302));
 sg13g2_inv_2 _1153_ (.Y(_0381_),
    .A(\hvsync_gen.vpos[9] ));
 sg13g2_inv_1 _1154_ (.Y(_0382_),
    .A(net324));
 sg13g2_inv_2 _1155_ (.Y(_0383_),
    .A(\hpos[5] ));
 sg13g2_inv_2 _1156_ (.Y(_0384_),
    .A(net80));
 sg13g2_inv_2 _1157_ (.Y(_0385_),
    .A(net318));
 sg13g2_inv_2 _1158_ (.Y(_0386_),
    .A(\hpos[6] ));
 sg13g2_inv_1 _1159_ (.Y(_0387_),
    .A(_0078_));
 sg13g2_inv_2 _1160_ (.Y(_0388_),
    .A(_0080_));
 sg13g2_inv_2 _1161_ (.Y(_0389_),
    .A(_0081_));
 sg13g2_inv_1 _1162_ (.Y(_0390_),
    .A(_0063_));
 sg13g2_and2_2 _1163_ (.A(\stage[1] ),
    .B(\stage[0] ),
    .X(_0391_));
 sg13g2_nand2_2 _1164_ (.Y(_0392_),
    .A(\stage[1] ),
    .B(\stage[0] ));
 sg13g2_or2_1 _1165_ (.X(_0393_),
    .B(\stage_seq_inst.stage_timer[1] ),
    .A(\stage_seq_inst.stage_timer[0] ));
 sg13g2_nor3_1 _1166_ (.A(\stage_seq_inst.stage_timer[2] ),
    .B(_0391_),
    .C(_0393_),
    .Y(_0394_));
 sg13g2_nor2b_1 _1167_ (.A(_0394_),
    .B_N(\stage_seq_inst.stage_timer[3] ),
    .Y(_0182_));
 sg13g2_nor4_2 _1168_ (.A(\stage_seq_inst.stage_timer[3] ),
    .B(\stage_seq_inst.stage_timer[2] ),
    .C(\stage_seq_inst.stage_timer[0] ),
    .Y(_0395_),
    .D(\stage_seq_inst.stage_timer[1] ));
 sg13g2_nand2b_2 _1169_ (.Y(_0396_),
    .B(_0395_),
    .A_N(\stage[1] ));
 sg13g2_nor2b_1 _1170_ (.A(\stage[1] ),
    .B_N(\stage[0] ),
    .Y(_0397_));
 sg13g2_nand2_1 _1171_ (.Y(_0398_),
    .A(_0395_),
    .B(_0397_));
 sg13g2_nand2_1 _1172_ (.Y(_0399_),
    .A(\stage_seq_inst.stage_timer[3] ),
    .B(_0394_));
 sg13g2_o21ai_1 _1173_ (.B1(\stage_seq_inst.stage_timer[2] ),
    .Y(_0400_),
    .A1(_0391_),
    .A2(_0393_));
 sg13g2_nand3_1 _1174_ (.B(_0399_),
    .C(_0400_),
    .A(_0398_),
    .Y(_0181_));
 sg13g2_nand2_1 _1175_ (.Y(_0401_),
    .A(_0103_),
    .B(_0391_));
 sg13g2_nand2_1 _1176_ (.Y(_0402_),
    .A(_0392_),
    .B(_0396_));
 sg13g2_nand2_1 _1177_ (.Y(_0403_),
    .A(\stage_seq_inst.stage_timer[0] ),
    .B(\stage_seq_inst.stage_timer[1] ));
 sg13g2_a21oi_1 _1178_ (.A1(_0393_),
    .A2(_0403_),
    .Y(_0404_),
    .B1(_0395_));
 sg13g2_o21ai_1 _1179_ (.B1(_0401_),
    .Y(_0180_),
    .A1(_0402_),
    .A2(_0404_));
 sg13g2_nand2_1 _1180_ (.Y(_0405_),
    .A(_0102_),
    .B(_0391_));
 sg13g2_nor2_1 _1181_ (.A(\stage_seq_inst.stage_timer[0] ),
    .B(_0395_),
    .Y(_0406_));
 sg13g2_o21ai_1 _1182_ (.B1(_0405_),
    .Y(_0179_),
    .A1(_0402_),
    .A2(_0406_));
 sg13g2_nor3_1 _1183_ (.A(net294),
    .B(_0373_),
    .C(\audio_mod.seq.seq_clock[2] ),
    .Y(_0407_));
 sg13g2_xnor2_1 _1184_ (.Y(_0408_),
    .A(\audio_mod.seq.seq_clock[3] ),
    .B(\audio_mod.seq.seq_clock[2] ));
 sg13g2_xor2_1 _1185_ (.B(\audio_mod.seq.seq_clock[2] ),
    .A(\audio_mod.seq.seq_clock[3] ),
    .X(_0409_));
 sg13g2_nor3_2 _1186_ (.A(net294),
    .B(net293),
    .C(_0408_),
    .Y(_0410_));
 sg13g2_or2_2 _1187_ (.X(_0411_),
    .B(_0410_),
    .A(_0407_));
 sg13g2_inv_1 _1188_ (.Y(_0412_),
    .A(_0411_));
 sg13g2_or3_1 _1189_ (.A(\audio_mod.audio_gen.chan3.ch_counter[5] ),
    .B(\audio_mod.audio_gen.chan3.ch_counter[6] ),
    .C(_0411_),
    .X(_0413_));
 sg13g2_nand3_1 _1190_ (.B(\audio_mod.audio_gen.chan3.ch_counter[6] ),
    .C(_0411_),
    .A(\audio_mod.audio_gen.chan3.ch_counter[5] ),
    .Y(_0414_));
 sg13g2_nand2_1 _1191_ (.Y(_0415_),
    .A(net293),
    .B(_0407_));
 sg13g2_nor2_1 _1192_ (.A(\audio_mod.audio_gen.chan3.ch_counter[0] ),
    .B(\audio_mod.audio_gen.chan3.ch_counter[1] ),
    .Y(_0416_));
 sg13g2_nor4_1 _1193_ (.A(\audio_mod.audio_gen.chan3.ch_counter[7] ),
    .B(\audio_mod.audio_gen.chan3.ch_counter[9] ),
    .C(\audio_mod.audio_gen.chan3.ch_counter[10] ),
    .D(\audio_mod.audio_gen.chan3.ch_counter[11] ),
    .Y(_0417_));
 sg13g2_nor4_1 _1194_ (.A(\audio_mod.audio_gen.chan3.ch_counter[3] ),
    .B(\audio_mod.audio_gen.chan3.ch_counter[4] ),
    .C(\audio_mod.audio_gen.chan3.ch_counter[8] ),
    .D(_0410_),
    .Y(_0418_));
 sg13g2_nand4_1 _1195_ (.B(\audio_mod.audio_gen.chan3.ch_counter[4] ),
    .C(\audio_mod.audio_gen.chan3.ch_counter[8] ),
    .A(\audio_mod.audio_gen.chan3.ch_counter[3] ),
    .Y(_0419_),
    .D(_0410_));
 sg13g2_nand2b_1 _1196_ (.Y(_0420_),
    .B(_0419_),
    .A_N(_0418_));
 sg13g2_xor2_1 _1197_ (.B(_0415_),
    .A(\audio_mod.audio_gen.chan3.ch_counter[2] ),
    .X(_0421_));
 sg13g2_nand4_1 _1198_ (.B(_0417_),
    .C(_0420_),
    .A(_0416_),
    .Y(_0422_),
    .D(_0421_));
 sg13g2_a21oi_2 _1199_ (.B1(_0422_),
    .Y(_0423_),
    .A2(_0414_),
    .A1(_0413_));
 sg13g2_mux2_1 _1200_ (.A0(\audio_mod.audio_gen.ch3_state ),
    .A1(\audio_mod.audio_gen.chan3.rng ),
    .S(_0423_),
    .X(_0168_));
 sg13g2_mux2_1 _1201_ (.A0(\background_color[2] ),
    .A1(\lfsr[2] ),
    .S(_0391_),
    .X(_0167_));
 sg13g2_mux2_1 _1202_ (.A0(\background_color[1] ),
    .A1(\lfsr[1] ),
    .S(_0391_),
    .X(_0166_));
 sg13g2_mux2_1 _1203_ (.A0(\audio_mod.audio_gen.chan3.rng ),
    .A1(\background_color[0] ),
    .S(_0392_),
    .X(_0165_));
 sg13g2_nand2_1 _1204_ (.Y(_0424_),
    .A(\audio_mod.seq.seq_clock[1] ),
    .B(\audio_mod.seq.seq_clock[0] ));
 sg13g2_nand2b_1 _1205_ (.Y(_0425_),
    .B(_0409_),
    .A_N(_0424_));
 sg13g2_nand2_1 _1206_ (.Y(_0426_),
    .A(\audio_mod.pattern_clock[1] ),
    .B(net291));
 sg13g2_and2_1 _1207_ (.A(net294),
    .B(net293),
    .X(_0427_));
 sg13g2_a22oi_1 _1208_ (.Y(_0428_),
    .B1(_0427_),
    .B2(net289),
    .A2(net291),
    .A1(net293));
 sg13g2_nor2b_1 _1209_ (.A(_0425_),
    .B_N(_0428_),
    .Y(_0429_));
 sg13g2_o21ai_1 _1210_ (.B1(net289),
    .Y(_0430_),
    .A1(net291),
    .A2(_0427_));
 sg13g2_and2_1 _1211_ (.A(_0409_),
    .B(_0424_),
    .X(_0431_));
 sg13g2_nor2_1 _1212_ (.A(\audio_mod.seq.seq_clock[1] ),
    .B(_0408_),
    .Y(_0432_));
 sg13g2_nand2_1 _1213_ (.Y(_0433_),
    .A(\audio_mod.seq.seq_clock[0] ),
    .B(_0426_));
 sg13g2_a221oi_1 _1214_ (.B2(_0433_),
    .C1(_0429_),
    .B1(_0432_),
    .A1(_0430_),
    .Y(_0434_),
    .A2(_0431_));
 sg13g2_nand3b_1 _1215_ (.B(net293),
    .C(net291),
    .Y(_0435_),
    .A_N(net294));
 sg13g2_nor2_1 _1216_ (.A(_0372_),
    .B(_0426_),
    .Y(_0436_));
 sg13g2_nand3_1 _1217_ (.B(net289),
    .C(net291),
    .A(net293),
    .Y(_0437_));
 sg13g2_nor2_1 _1218_ (.A(\audio_mod.pattern_clock[0] ),
    .B(_0437_),
    .Y(_0438_));
 sg13g2_nand3_1 _1219_ (.B(_0432_),
    .C(_0438_),
    .A(\audio_mod.seq.seq_clock[0] ),
    .Y(_0439_));
 sg13g2_nor2_1 _1220_ (.A(_0425_),
    .B(_0428_),
    .Y(_0440_));
 sg13g2_nand2b_1 _1221_ (.Y(_0441_),
    .B(\audio_mod.seq.seq_clock[1] ),
    .A_N(\audio_mod.seq.seq_clock[0] ));
 sg13g2_nor2_1 _1222_ (.A(_0430_),
    .B(_0441_),
    .Y(_0442_));
 sg13g2_a22oi_1 _1223_ (.Y(_0443_),
    .B1(_0442_),
    .B2(_0409_),
    .A2(_0440_),
    .A1(_0437_));
 sg13g2_nand2_1 _1224_ (.Y(_0444_),
    .A(_0439_),
    .B(_0443_));
 sg13g2_or2_2 _1225_ (.X(_0445_),
    .B(_0444_),
    .A(_0434_));
 sg13g2_o21ai_1 _1226_ (.B1(_0432_),
    .Y(_0446_),
    .A1(_0051_),
    .A2(_0437_));
 sg13g2_o21ai_1 _1227_ (.B1(_0446_),
    .Y(_0447_),
    .A1(_0425_),
    .A2(_0437_));
 sg13g2_nor2b_1 _1228_ (.A(_0445_),
    .B_N(_0447_),
    .Y(_0448_));
 sg13g2_nand2_1 _1229_ (.Y(_0449_),
    .A(_0443_),
    .B(_0445_));
 sg13g2_nor2b_1 _1230_ (.A(_0444_),
    .B_N(_0445_),
    .Y(_0450_));
 sg13g2_nor2b_2 _1231_ (.A(_0447_),
    .B_N(_0439_),
    .Y(_0451_));
 sg13g2_a21oi_1 _1232_ (.A1(\audio_mod.audio_gen.chan2.ch_counter[4] ),
    .A2(\audio_mod.audio_gen.chan2.ch_counter[7] ),
    .Y(_0452_),
    .B1(_0451_));
 sg13g2_o21ai_1 _1233_ (.B1(_0451_),
    .Y(_0453_),
    .A1(\audio_mod.audio_gen.chan2.ch_counter[4] ),
    .A2(\audio_mod.audio_gen.chan2.ch_counter[7] ));
 sg13g2_nand3_1 _1234_ (.B(_0443_),
    .C(_0451_),
    .A(\audio_mod.audio_gen.chan2.ch_counter[3] ),
    .Y(_0454_));
 sg13g2_a21oi_1 _1235_ (.A1(_0443_),
    .A2(_0451_),
    .Y(_0455_),
    .B1(\audio_mod.audio_gen.chan2.ch_counter[3] ));
 sg13g2_o21ai_1 _1236_ (.B1(_0439_),
    .Y(_0456_),
    .A1(_0445_),
    .A2(_0447_));
 sg13g2_a21oi_1 _1237_ (.A1(_0434_),
    .A2(_0447_),
    .Y(_0457_),
    .B1(_0456_));
 sg13g2_nand2_1 _1238_ (.Y(_0458_),
    .A(\audio_mod.audio_gen.chan2.ch_counter[9] ),
    .B(\audio_mod.audio_gen.chan2.ch_counter[10] ));
 sg13g2_xnor2_1 _1239_ (.Y(_0459_),
    .A(\audio_mod.audio_gen.chan2.ch_counter[5] ),
    .B(_0456_));
 sg13g2_a21oi_1 _1240_ (.A1(\audio_mod.audio_gen.chan2.ch_counter[10] ),
    .A2(_0445_),
    .Y(_0460_),
    .B1(\audio_mod.audio_gen.chan2.ch_counter[9] ));
 sg13g2_o21ai_1 _1241_ (.B1(_0460_),
    .Y(_0461_),
    .A1(\audio_mod.audio_gen.chan2.ch_counter[10] ),
    .A2(_0445_));
 sg13g2_xnor2_1 _1242_ (.Y(_0462_),
    .A(\audio_mod.audio_gen.chan2.ch_counter[0] ),
    .B(_0448_));
 sg13g2_a21oi_1 _1243_ (.A1(\audio_mod.audio_gen.chan2.ch_counter[2] ),
    .A2(_0450_),
    .Y(_0463_),
    .B1(_0452_));
 sg13g2_xor2_1 _1244_ (.B(_0450_),
    .A(\audio_mod.audio_gen.chan2.ch_counter[6] ),
    .X(_0464_));
 sg13g2_nand4_1 _1245_ (.B(_0462_),
    .C(_0463_),
    .A(_0459_),
    .Y(_0465_),
    .D(_0464_));
 sg13g2_mux2_1 _1246_ (.A0(_0458_),
    .A1(_0461_),
    .S(_0457_),
    .X(_0466_));
 sg13g2_o21ai_1 _1247_ (.B1(_0453_),
    .Y(_0467_),
    .A1(\audio_mod.audio_gen.chan2.ch_counter[2] ),
    .A2(_0450_));
 sg13g2_a22oi_1 _1248_ (.Y(_0468_),
    .B1(_0445_),
    .B2(\audio_mod.audio_gen.chan2.ch_counter[8] ),
    .A2(_0443_),
    .A1(_0380_));
 sg13g2_nand3_1 _1249_ (.B(_0443_),
    .C(_0445_),
    .A(\audio_mod.audio_gen.chan2.ch_counter[1] ),
    .Y(_0469_));
 sg13g2_o21ai_1 _1250_ (.B1(\audio_mod.audio_gen.chan2.ch_counter[1] ),
    .Y(_0470_),
    .A1(\audio_mod.audio_gen.chan2.ch_counter[8] ),
    .A2(_0380_));
 sg13g2_a21oi_1 _1251_ (.A1(_0449_),
    .A2(_0470_),
    .Y(_0471_),
    .B1(_0455_));
 sg13g2_nand4_1 _1252_ (.B(_0468_),
    .C(_0469_),
    .A(_0454_),
    .Y(_0472_),
    .D(_0471_));
 sg13g2_nor4_1 _1253_ (.A(_0465_),
    .B(_0466_),
    .C(_0467_),
    .D(_0472_),
    .Y(_0473_));
 sg13g2_mux2_1 _1254_ (.A0(\audio_mod.audio_gen.ch2_state ),
    .A1(_0038_),
    .S(net278),
    .X(_0164_));
 sg13g2_nor2_1 _1255_ (.A(\audio_mod.seq.seq_clock[3] ),
    .B(_0374_),
    .Y(_0474_));
 sg13g2_a21oi_2 _1256_ (.B1(_0374_),
    .Y(_0475_),
    .A2(\audio_mod.seq.seq_clock[2] ),
    .A1(\audio_mod.seq.seq_clock[3] ));
 sg13g2_xor2_1 _1257_ (.B(net293),
    .A(\audio_mod.pattern_clock[0] ),
    .X(_0096_));
 sg13g2_o21ai_1 _1258_ (.B1(_0435_),
    .Y(_0476_),
    .A1(net291),
    .A2(_0096_));
 sg13g2_a22oi_1 _1259_ (.Y(_0477_),
    .B1(_0476_),
    .B2(_0372_),
    .A2(_0436_),
    .A1(net294));
 sg13g2_nor2_1 _1260_ (.A(net293),
    .B(net291),
    .Y(_0478_));
 sg13g2_nor3_1 _1261_ (.A(net294),
    .B(_0372_),
    .C(_0478_),
    .Y(_0479_));
 sg13g2_a221oi_1 _1262_ (.B2(_0372_),
    .C1(_0479_),
    .B1(_0476_),
    .A1(net294),
    .Y(_0480_),
    .A2(_0436_));
 sg13g2_a21oi_1 _1263_ (.A1(\audio_mod.seq.seq_clock[3] ),
    .A2(\audio_mod.seq.seq_clock[2] ),
    .Y(_0481_),
    .B1(_0424_));
 sg13g2_nand3_1 _1264_ (.B(_0476_),
    .C(_0481_),
    .A(net289),
    .Y(_0482_));
 sg13g2_o21ai_1 _1265_ (.B1(_0482_),
    .Y(_0483_),
    .A1(_0475_),
    .A2(_0480_));
 sg13g2_nand3_1 _1266_ (.B(_0475_),
    .C(_0476_),
    .A(_0372_),
    .Y(_0484_));
 sg13g2_a21oi_1 _1267_ (.A1(_0481_),
    .A2(_0484_),
    .Y(_0485_),
    .B1(_0477_));
 sg13g2_nor2_2 _1268_ (.A(net284),
    .B(_0485_),
    .Y(_0486_));
 sg13g2_xnor2_1 _1269_ (.Y(_0487_),
    .A(net284),
    .B(net283));
 sg13g2_nor4_2 _1270_ (.A(\audio_mod.pattern_clock[0] ),
    .B(_0372_),
    .C(_0441_),
    .Y(_0488_),
    .D(_0478_));
 sg13g2_o21ai_1 _1271_ (.B1(_0488_),
    .Y(_0489_),
    .A1(_0409_),
    .A2(_0474_));
 sg13g2_nor2b_1 _1272_ (.A(net284),
    .B_N(_0489_),
    .Y(_0490_));
 sg13g2_xor2_1 _1273_ (.B(_0490_),
    .A(\audio_mod.audio_gen.chan1.ch_counter[2] ),
    .X(_0491_));
 sg13g2_nand2b_1 _1274_ (.Y(_0492_),
    .B(_0489_),
    .A_N(net283));
 sg13g2_and3_1 _1275_ (.X(_0493_),
    .A(\audio_mod.audio_gen.chan1.ch_counter[0] ),
    .B(\audio_mod.audio_gen.chan1.ch_counter[5] ),
    .C(_0492_));
 sg13g2_nor3_1 _1276_ (.A(\audio_mod.audio_gen.chan1.ch_counter[0] ),
    .B(\audio_mod.audio_gen.chan1.ch_counter[5] ),
    .C(_0492_),
    .Y(_0494_));
 sg13g2_nor2_1 _1277_ (.A(_0438_),
    .B(_0488_),
    .Y(_0495_));
 sg13g2_nor2b_1 _1278_ (.A(_0495_),
    .B_N(_0475_),
    .Y(_0496_));
 sg13g2_o21ai_1 _1279_ (.B1(_0475_),
    .Y(_0497_),
    .A1(_0438_),
    .A2(_0488_));
 sg13g2_nand2_2 _1280_ (.Y(_0498_),
    .A(_0483_),
    .B(_0497_));
 sg13g2_nand2b_1 _1281_ (.Y(_0499_),
    .B(_0498_),
    .A_N(_0486_));
 sg13g2_xnor2_1 _1282_ (.Y(_0500_),
    .A(\audio_mod.audio_gen.chan1.ch_counter[3] ),
    .B(net284));
 sg13g2_nor2_1 _1283_ (.A(\audio_mod.audio_gen.chan1.ch_counter[10] ),
    .B(_0489_),
    .Y(_0501_));
 sg13g2_xor2_1 _1284_ (.B(\audio_mod.audio_gen.chan1.ch_counter[1] ),
    .A(\audio_mod.audio_gen.chan1.ch_counter[0] ),
    .X(_0016_));
 sg13g2_nand2_1 _1285_ (.Y(_0502_),
    .A(\audio_mod.audio_gen.chan1.ch_counter[10] ),
    .B(_0489_));
 sg13g2_xor2_1 _1286_ (.B(_0498_),
    .A(\audio_mod.audio_gen.chan1.ch_counter[6] ),
    .X(_0503_));
 sg13g2_xnor2_1 _1287_ (.Y(_0504_),
    .A(\audio_mod.audio_gen.chan1.ch_counter[8] ),
    .B(_0487_));
 sg13g2_nand2_1 _1288_ (.Y(_0505_),
    .A(_0378_),
    .B(net283));
 sg13g2_a21oi_1 _1289_ (.A1(\audio_mod.audio_gen.chan1.ch_counter[9] ),
    .A2(_0505_),
    .Y(_0506_),
    .B1(_0486_));
 sg13g2_a21oi_1 _1290_ (.A1(\audio_mod.audio_gen.chan1.ch_counter[9] ),
    .A2(_0486_),
    .Y(_0507_),
    .B1(_0506_));
 sg13g2_o21ai_1 _1291_ (.B1(_0502_),
    .Y(_0508_),
    .A1(_0378_),
    .A2(net283));
 sg13g2_nor4_1 _1292_ (.A(\audio_mod.audio_gen.chan1.ch_counter[11] ),
    .B(_0501_),
    .C(_0016_),
    .D(_0508_),
    .Y(_0509_));
 sg13g2_nand4_1 _1293_ (.B(_0503_),
    .C(_0507_),
    .A(_0500_),
    .Y(_0510_),
    .D(_0509_));
 sg13g2_o21ai_1 _1294_ (.B1(_0491_),
    .Y(_0511_),
    .A1(_0493_),
    .A2(_0494_));
 sg13g2_xnor2_1 _1295_ (.Y(_0512_),
    .A(\audio_mod.audio_gen.chan1.ch_counter[4] ),
    .B(_0499_));
 sg13g2_nor4_2 _1296_ (.A(_0504_),
    .B(_0510_),
    .C(_0511_),
    .Y(_0513_),
    .D(_0512_));
 sg13g2_mux2_1 _1297_ (.A0(\audio_mod.audio_gen.ch1_state ),
    .A1(_0025_),
    .S(_0513_),
    .X(_0163_));
 sg13g2_xor2_1 _1298_ (.B(_0490_),
    .A(\audio_mod.audio_gen.chan0.ch_counter[3] ),
    .X(_0514_));
 sg13g2_xor2_1 _1299_ (.B(_0499_),
    .A(\audio_mod.audio_gen.chan0.ch_counter[5] ),
    .X(_0515_));
 sg13g2_nand2_1 _1300_ (.Y(_0516_),
    .A(_0514_),
    .B(_0515_));
 sg13g2_nand2_1 _1301_ (.Y(_0517_),
    .A(\audio_mod.audio_gen.chan0.ch_counter[10] ),
    .B(_0486_));
 sg13g2_xor2_1 _1302_ (.B(_0489_),
    .A(\audio_mod.audio_gen.chan0.ch_counter[11] ),
    .X(_0518_));
 sg13g2_xnor2_1 _1303_ (.Y(_0519_),
    .A(\audio_mod.audio_gen.chan0.ch_counter[8] ),
    .B(net283));
 sg13g2_nor2_1 _1304_ (.A(\audio_mod.audio_gen.chan0.ch_counter[10] ),
    .B(_0486_),
    .Y(_0520_));
 sg13g2_nand4_1 _1305_ (.B(\audio_mod.audio_gen.chan0.ch_counter[2] ),
    .C(\audio_mod.audio_gen.chan0.ch_counter[6] ),
    .A(\audio_mod.audio_gen.chan0.ch_counter[1] ),
    .Y(_0521_),
    .D(_0492_));
 sg13g2_or4_1 _1306_ (.A(\audio_mod.audio_gen.chan0.ch_counter[1] ),
    .B(\audio_mod.audio_gen.chan0.ch_counter[2] ),
    .C(\audio_mod.audio_gen.chan0.ch_counter[6] ),
    .D(_0492_),
    .X(_0522_));
 sg13g2_a21oi_1 _1307_ (.A1(_0521_),
    .A2(_0522_),
    .Y(_0523_),
    .B1(_0520_));
 sg13g2_nand4_1 _1308_ (.B(_0518_),
    .C(_0519_),
    .A(_0517_),
    .Y(_0524_),
    .D(_0523_));
 sg13g2_xnor2_1 _1309_ (.Y(_0525_),
    .A(\audio_mod.audio_gen.chan0.ch_counter[9] ),
    .B(_0487_));
 sg13g2_o21ai_1 _1310_ (.B1(net284),
    .Y(_0526_),
    .A1(net283),
    .A2(_0496_));
 sg13g2_xor2_1 _1311_ (.B(_0526_),
    .A(\audio_mod.audio_gen.chan0.ch_counter[0] ),
    .X(_0527_));
 sg13g2_xnor2_1 _1312_ (.Y(_0528_),
    .A(\audio_mod.audio_gen.chan0.ch_counter[4] ),
    .B(net284));
 sg13g2_o21ai_1 _1313_ (.B1(_0528_),
    .Y(_0529_),
    .A1(\audio_mod.audio_gen.chan0.ch_counter[7] ),
    .A2(_0498_));
 sg13g2_a21oi_1 _1314_ (.A1(\audio_mod.audio_gen.chan0.ch_counter[7] ),
    .A2(_0498_),
    .Y(_0530_),
    .B1(_0529_));
 sg13g2_nand2_1 _1315_ (.Y(_0531_),
    .A(_0527_),
    .B(_0530_));
 sg13g2_nor4_1 _1316_ (.A(_0516_),
    .B(_0524_),
    .C(_0525_),
    .D(_0531_),
    .Y(_0532_));
 sg13g2_mux2_1 _1317_ (.A0(\audio_mod.audio_gen.ch0_state ),
    .A1(_0012_),
    .S(net280),
    .X(_0162_));
 sg13g2_nand2b_1 _1318_ (.Y(_0161_),
    .B(_0398_),
    .A_N(\stage[1] ));
 sg13g2_a22oi_1 _1319_ (.Y(_0533_),
    .B1(_0396_),
    .B2(\stage[0] ),
    .A2(_0395_),
    .A1(_0101_));
 sg13g2_inv_1 _1320_ (.Y(_0160_),
    .A(_0533_));
 sg13g2_nand3b_1 _1321_ (.B(net298),
    .C(_0409_),
    .Y(_0534_),
    .A_N(net300));
 sg13g2_nor3_1 _1322_ (.A(net284),
    .B(net283),
    .C(_0496_),
    .Y(_0535_));
 sg13g2_or3_2 _1323_ (.A(net284),
    .B(net283),
    .C(_0496_),
    .X(_0536_));
 sg13g2_nand2_2 _1324_ (.Y(_0537_),
    .A(net300),
    .B(net298));
 sg13g2_and2_1 _1325_ (.A(_0536_),
    .B(_0537_),
    .X(_0538_));
 sg13g2_nand2_1 _1326_ (.Y(_0539_),
    .A(_0536_),
    .B(_0537_));
 sg13g2_nand2_1 _1327_ (.Y(_0540_),
    .A(_0534_),
    .B(_0539_));
 sg13g2_nand3_1 _1328_ (.B(_0536_),
    .C(_0537_),
    .A(\audio_mod.audio_gen.ch1_state ),
    .Y(_0541_));
 sg13g2_nand2_1 _1329_ (.Y(_0542_),
    .A(_0073_),
    .B(_0541_));
 sg13g2_xor2_1 _1330_ (.B(_0541_),
    .A(_0073_),
    .X(_0543_));
 sg13g2_a21oi_1 _1331_ (.A1(_0534_),
    .A2(_0539_),
    .Y(_0544_),
    .B1(_0543_));
 sg13g2_mux2_1 _1332_ (.A0(_0073_),
    .A1(_0543_),
    .S(_0540_),
    .X(_0545_));
 sg13g2_nand2_1 _1333_ (.Y(_0546_),
    .A(_0409_),
    .B(_0537_));
 sg13g2_a21oi_1 _1334_ (.A1(\audio_mod.audio_gen.ch2_state ),
    .A2(net298),
    .Y(_0547_),
    .B1(_0546_));
 sg13g2_a21oi_1 _1335_ (.A1(_0545_),
    .A2(_0547_),
    .Y(_0548_),
    .B1(_0544_));
 sg13g2_nand2b_2 _1336_ (.Y(_0549_),
    .B(_0411_),
    .A_N(net298));
 sg13g2_nor2_2 _1337_ (.A(\audio_mod.audio_gen.ch3_state ),
    .B(_0549_),
    .Y(_0550_));
 sg13g2_nand3_1 _1338_ (.B(_0409_),
    .C(_0537_),
    .A(_0038_),
    .Y(_0551_));
 sg13g2_a221oi_1 _1339_ (.B2(_0497_),
    .C1(\audio_mod.audio_gen.ch1_state ),
    .B1(_0486_),
    .A1(net300),
    .Y(_0552_),
    .A2(net298));
 sg13g2_nor2b_1 _1340_ (.A(_0551_),
    .B_N(_0552_),
    .Y(_0553_));
 sg13g2_xor2_1 _1341_ (.B(_0552_),
    .A(_0551_),
    .X(_0554_));
 sg13g2_nand2_1 _1342_ (.Y(_0555_),
    .A(_0542_),
    .B(_0554_));
 sg13g2_xor2_1 _1343_ (.B(_0554_),
    .A(_0542_),
    .X(_0556_));
 sg13g2_nand2_1 _1344_ (.Y(_0557_),
    .A(_0550_),
    .B(_0556_));
 sg13g2_xnor2_1 _1345_ (.Y(_0558_),
    .A(_0550_),
    .B(_0556_));
 sg13g2_or2_1 _1346_ (.X(_0559_),
    .B(_0558_),
    .A(_0548_));
 sg13g2_nand2_2 _1347_ (.Y(_0560_),
    .A(_0012_),
    .B(_0538_));
 sg13g2_xor2_1 _1348_ (.B(_0558_),
    .A(_0548_),
    .X(_0561_));
 sg13g2_nand2b_1 _1349_ (.Y(_0562_),
    .B(_0561_),
    .A_N(_0560_));
 sg13g2_nand2_1 _1350_ (.Y(_0563_),
    .A(_0559_),
    .B(_0562_));
 sg13g2_nand2_1 _1351_ (.Y(_0564_),
    .A(_0550_),
    .B(_0553_));
 sg13g2_xor2_1 _1352_ (.B(_0553_),
    .A(_0550_),
    .X(_0565_));
 sg13g2_and3_1 _1353_ (.X(_0566_),
    .A(_0555_),
    .B(_0557_),
    .C(_0565_));
 sg13g2_a21oi_1 _1354_ (.A1(_0555_),
    .A2(_0557_),
    .Y(_0567_),
    .B1(_0565_));
 sg13g2_nor2_1 _1355_ (.A(_0566_),
    .B(_0567_),
    .Y(_0568_));
 sg13g2_xor2_1 _1356_ (.B(_0568_),
    .A(_0560_),
    .X(_0569_));
 sg13g2_a21o_1 _1357_ (.A2(_0562_),
    .A1(_0559_),
    .B1(_0569_),
    .X(_0570_));
 sg13g2_nor3_1 _1358_ (.A(net298),
    .B(_0412_),
    .C(_0536_),
    .Y(_0571_));
 sg13g2_xnor2_1 _1359_ (.Y(_0572_),
    .A(_0545_),
    .B(_0547_));
 sg13g2_nor4_1 _1360_ (.A(net298),
    .B(_0412_),
    .C(_0536_),
    .D(_0572_),
    .Y(_0573_));
 sg13g2_xnor2_1 _1361_ (.Y(_0574_),
    .A(\audio_mod.audio_gen.ch3_state ),
    .B(net300));
 sg13g2_nor2_1 _1362_ (.A(_0549_),
    .B(_0574_),
    .Y(_0575_));
 sg13g2_xnor2_1 _1363_ (.Y(_0576_),
    .A(_0571_),
    .B(_0572_));
 sg13g2_a21oi_1 _1364_ (.A1(_0575_),
    .A2(_0576_),
    .Y(_0577_),
    .B1(_0573_));
 sg13g2_xnor2_1 _1365_ (.Y(_0578_),
    .A(_0560_),
    .B(_0561_));
 sg13g2_nor2b_1 _1366_ (.A(_0577_),
    .B_N(_0578_),
    .Y(_0579_));
 sg13g2_xnor2_1 _1367_ (.Y(_0580_),
    .A(_0575_),
    .B(_0576_));
 sg13g2_a221oi_1 _1368_ (.B2(_0549_),
    .C1(_0535_),
    .B1(_0534_),
    .A1(net300),
    .Y(_0581_),
    .A2(net298));
 sg13g2_a21oi_1 _1369_ (.A1(\audio_mod.audio_gen.ch0_state ),
    .A2(_0538_),
    .Y(_0582_),
    .B1(_0581_));
 sg13g2_nand2_1 _1370_ (.Y(_0583_),
    .A(\audio_mod.audio_gen.ch0_state ),
    .B(_0581_));
 sg13g2_o21ai_1 _1371_ (.B1(_0583_),
    .Y(_0584_),
    .A1(_0580_),
    .A2(_0582_));
 sg13g2_xnor2_1 _1372_ (.Y(_0585_),
    .A(_0577_),
    .B(_0578_));
 sg13g2_a21oi_1 _1373_ (.A1(_0584_),
    .A2(_0585_),
    .Y(_0586_),
    .B1(_0579_));
 sg13g2_xor2_1 _1374_ (.B(_0569_),
    .A(_0563_),
    .X(_0587_));
 sg13g2_o21ai_1 _1375_ (.B1(_0570_),
    .Y(_0588_),
    .A1(_0586_),
    .A2(_0587_));
 sg13g2_mux2_1 _1376_ (.A0(_0566_),
    .A1(_0567_),
    .S(_0560_),
    .X(_0589_));
 sg13g2_xnor2_1 _1377_ (.Y(_0590_),
    .A(_0564_),
    .B(_0589_));
 sg13g2_xnor2_1 _1378_ (.Y(_0591_),
    .A(_0588_),
    .B(_0590_));
 sg13g2_or2_1 _1379_ (.X(_0592_),
    .B(_0591_),
    .A(net337));
 sg13g2_and2_1 _1380_ (.A(net336),
    .B(_0591_),
    .X(_0593_));
 sg13g2_xnor2_1 _1381_ (.Y(_0594_),
    .A(_0586_),
    .B(_0587_));
 sg13g2_nor2_1 _1382_ (.A(\audio_mod.audio_gen.pwm_clock[4] ),
    .B(_0594_),
    .Y(_0595_));
 sg13g2_nand2_1 _1383_ (.Y(_0596_),
    .A(\audio_mod.audio_gen.pwm_clock[4] ),
    .B(_0594_));
 sg13g2_xnor2_1 _1384_ (.Y(_0597_),
    .A(_0584_),
    .B(_0585_));
 sg13g2_a21oi_1 _1385_ (.A1(_0534_),
    .A2(_0549_),
    .Y(_0598_),
    .B1(_0375_));
 sg13g2_nand2_1 _1386_ (.Y(_0599_),
    .A(net346),
    .B(_0598_));
 sg13g2_nor2_1 _1387_ (.A(net346),
    .B(_0598_),
    .Y(_0600_));
 sg13g2_nor2b_1 _1388_ (.A(_0582_),
    .B_N(_0583_),
    .Y(_0601_));
 sg13g2_xnor2_1 _1389_ (.Y(_0602_),
    .A(_0580_),
    .B(_0601_));
 sg13g2_o21ai_1 _1390_ (.B1(_0599_),
    .Y(_0603_),
    .A1(_0600_),
    .A2(_0602_));
 sg13g2_a21o_1 _1391_ (.A2(_0597_),
    .A1(\audio_mod.audio_gen.pwm_clock[3] ),
    .B1(_0603_),
    .X(_0604_));
 sg13g2_o21ai_1 _1392_ (.B1(_0604_),
    .Y(_0605_),
    .A1(\audio_mod.audio_gen.pwm_clock[3] ),
    .A2(_0597_));
 sg13g2_a21oi_1 _1393_ (.A1(_0596_),
    .A2(_0605_),
    .Y(_0606_),
    .B1(_0595_));
 sg13g2_a21oi_1 _1394_ (.A1(_0592_),
    .A2(_0606_),
    .Y(audio),
    .B1(_0593_));
 sg13g2_nand2_1 _1395_ (.Y(_0607_),
    .A(_0381_),
    .B(\hvsync_gen.vpos[8] ));
 sg13g2_nor2_1 _1396_ (.A(\hvsync_gen.vpos[2] ),
    .B(_0607_),
    .Y(_0608_));
 sg13g2_nand3_1 _1397_ (.B(\hvsync_gen.vpos[1] ),
    .C(_0608_),
    .A(\hvsync_gen.vpos[3] ),
    .Y(_0609_));
 sg13g2_nand2_1 _1398_ (.Y(_0610_),
    .A(\hvsync_gen.vpos[6] ),
    .B(net325));
 sg13g2_nand3_1 _1399_ (.B(\hvsync_gen.vpos[6] ),
    .C(net324),
    .A(net322),
    .Y(_0611_));
 sg13g2_nor3_1 _1400_ (.A(net49),
    .B(_0609_),
    .C(_0611_),
    .Y(_0059_));
 sg13g2_nand2_1 _1401_ (.Y(_0612_),
    .A(net316),
    .B(\hpos[8] ));
 sg13g2_nand3_1 _1402_ (.B(_0384_),
    .C(_0386_),
    .A(_0383_),
    .Y(_0613_));
 sg13g2_nand3_1 _1403_ (.B(net316),
    .C(_0613_),
    .A(net318),
    .Y(_0614_));
 sg13g2_nand2_2 _1404_ (.Y(_0615_),
    .A(\hpos[5] ),
    .B(\hpos[4] ));
 sg13g2_nand4_1 _1405_ (.B(\hpos[4] ),
    .C(net318),
    .A(\hpos[5] ),
    .Y(_0616_),
    .D(\hpos[6] ));
 sg13g2_nor2b_1 _1406_ (.A(\hpos[8] ),
    .B_N(net316),
    .Y(_0617_));
 sg13g2_a21oi_1 _1407_ (.A1(_0616_),
    .A2(_0617_),
    .Y(_0618_),
    .B1(net60));
 sg13g2_a21oi_1 _1408_ (.A1(_0612_),
    .A2(_0614_),
    .Y(_0058_),
    .B1(net61));
 sg13g2_and2_1 _1409_ (.A(\counter[0] ),
    .B(net306),
    .X(_0619_));
 sg13g2_nand2_1 _1410_ (.Y(_0620_),
    .A(net306),
    .B(net305));
 sg13g2_xor2_1 _1411_ (.B(net297),
    .A(net305),
    .X(_0086_));
 sg13g2_nand4_1 _1412_ (.B(net323),
    .C(\hvsync_gen.vpos[6] ),
    .A(net321),
    .Y(_0621_),
    .D(net325));
 sg13g2_nor2_1 _1413_ (.A(\hpos[7] ),
    .B(\hpos[8] ),
    .Y(_0622_));
 sg13g2_o21ai_1 _1414_ (.B1(_0381_),
    .Y(_0623_),
    .A1(_0075_),
    .A2(_0622_));
 sg13g2_nor2b_1 _1415_ (.A(_0623_),
    .B_N(_0621_),
    .Y(_0624_));
 sg13g2_and2_1 _1416_ (.A(\lfsr[5] ),
    .B(\lfsr[4] ),
    .X(_0625_));
 sg13g2_nand2_1 _1417_ (.Y(_0626_),
    .A(\lfsr[5] ),
    .B(\lfsr[4] ));
 sg13g2_nor3_2 _1418_ (.A(\hpos[3] ),
    .B(net319),
    .C(\hpos[4] ),
    .Y(_0627_));
 sg13g2_or3_1 _1419_ (.A(\hpos[3] ),
    .B(net319),
    .C(\hpos[4] ),
    .X(_0628_));
 sg13g2_nor2_1 _1420_ (.A(_0383_),
    .B(_0627_),
    .Y(_0629_));
 sg13g2_nor3_2 _1421_ (.A(_0383_),
    .B(_0386_),
    .C(_0627_),
    .Y(_0630_));
 sg13g2_nand3_1 _1422_ (.B(\hpos[6] ),
    .C(_0628_),
    .A(\hpos[5] ),
    .Y(_0631_));
 sg13g2_nand3_1 _1423_ (.B(\hpos[8] ),
    .C(_0630_),
    .A(\hpos[7] ),
    .Y(_0632_));
 sg13g2_nand2b_2 _1424_ (.Y(_0633_),
    .B(net290),
    .A_N(net292));
 sg13g2_a21oi_1 _1425_ (.A1(_0397_),
    .A2(_0633_),
    .Y(_0634_),
    .B1(net316));
 sg13g2_nand2_2 _1426_ (.Y(_0635_),
    .A(_0632_),
    .B(_0634_));
 sg13g2_nor2_2 _1427_ (.A(net81),
    .B(net320),
    .Y(_0636_));
 sg13g2_nor2_1 _1428_ (.A(_0383_),
    .B(\hpos[4] ),
    .Y(_0637_));
 sg13g2_nor2b_1 _1429_ (.A(\hpos[3] ),
    .B_N(net319),
    .Y(_0638_));
 sg13g2_nand3_1 _1430_ (.B(_0637_),
    .C(_0638_),
    .A(_0636_),
    .Y(_0639_));
 sg13g2_o21ai_1 _1431_ (.B1(\hpos[2] ),
    .Y(_0640_),
    .A1(\hpos[0] ),
    .A2(net320));
 sg13g2_nor2b_2 _1432_ (.A(\hpos[3] ),
    .B_N(_0640_),
    .Y(_0641_));
 sg13g2_a21o_1 _1433_ (.A2(_0641_),
    .A1(_0637_),
    .B1(_0078_),
    .X(_0642_));
 sg13g2_a21oi_1 _1434_ (.A1(_0639_),
    .A2(_0642_),
    .Y(_0643_),
    .B1(_0386_));
 sg13g2_nor2b_2 _1435_ (.A(_0643_),
    .B_N(_0622_),
    .Y(_0644_));
 sg13g2_nor2_2 _1436_ (.A(net322),
    .B(\hvsync_gen.vpos[6] ),
    .Y(_0645_));
 sg13g2_nor2_2 _1437_ (.A(\hvsync_gen.vpos[0] ),
    .B(\hvsync_gen.vpos[1] ),
    .Y(_0646_));
 sg13g2_nand2b_2 _1438_ (.Y(_0647_),
    .B(_0646_),
    .A_N(\hvsync_gen.vpos[2] ));
 sg13g2_nand3_1 _1439_ (.B(net327),
    .C(_0647_),
    .A(\hvsync_gen.vpos[4] ),
    .Y(_0648_));
 sg13g2_and2_1 _1440_ (.A(_0382_),
    .B(_0648_),
    .X(_0649_));
 sg13g2_and2_1 _1441_ (.A(_0645_),
    .B(_0649_),
    .X(_0650_));
 sg13g2_nand2_1 _1442_ (.Y(_0651_),
    .A(_0645_),
    .B(_0649_));
 sg13g2_a21oi_1 _1443_ (.A1(net321),
    .A2(_0651_),
    .Y(_0652_),
    .B1(\hvsync_gen.vpos[9] ));
 sg13g2_nand3_1 _1444_ (.B(net327),
    .C(_0645_),
    .A(net326),
    .Y(_0653_));
 sg13g2_or4_1 _1445_ (.A(net324),
    .B(_0607_),
    .C(_0647_),
    .D(_0653_),
    .X(_0654_));
 sg13g2_nand2_1 _1446_ (.Y(_0655_),
    .A(_0652_),
    .B(_0654_));
 sg13g2_nor4_2 _1447_ (.A(_0383_),
    .B(net318),
    .C(_0386_),
    .Y(_0656_),
    .D(_0627_));
 sg13g2_nand4_1 _1448_ (.B(_0385_),
    .C(\hpos[6] ),
    .A(\hpos[5] ),
    .Y(_0657_),
    .D(_0628_));
 sg13g2_xnor2_1 _1449_ (.Y(_0658_),
    .A(\hpos[7] ),
    .B(_0630_));
 sg13g2_xnor2_1 _1450_ (.Y(_0659_),
    .A(_0385_),
    .B(_0630_));
 sg13g2_nor3_2 _1451_ (.A(_0388_),
    .B(_0389_),
    .C(_0656_),
    .Y(_0660_));
 sg13g2_a21oi_1 _1452_ (.A1(net317),
    .A2(_0657_),
    .Y(_0661_),
    .B1(_0081_));
 sg13g2_a21oi_2 _1453_ (.B1(_0389_),
    .Y(_0662_),
    .A2(_0657_),
    .A1(net317));
 sg13g2_o21ai_1 _1454_ (.B1(_0081_),
    .Y(_0663_),
    .A1(_0388_),
    .A2(_0656_));
 sg13g2_nor3_2 _1455_ (.A(_0388_),
    .B(_0081_),
    .C(_0656_),
    .Y(_0664_));
 sg13g2_nand3_1 _1456_ (.B(_0389_),
    .C(_0657_),
    .A(net317),
    .Y(_0665_));
 sg13g2_nor2_1 _1457_ (.A(_0662_),
    .B(_0664_),
    .Y(_0666_));
 sg13g2_nand3_1 _1458_ (.B(_0663_),
    .C(_0665_),
    .A(_0658_),
    .Y(_0667_));
 sg13g2_o21ai_1 _1459_ (.B1(_0659_),
    .Y(_0668_),
    .A1(_0662_),
    .A2(_0664_));
 sg13g2_nand2_1 _1460_ (.Y(_0669_),
    .A(_0667_),
    .B(_0668_));
 sg13g2_a21oi_2 _1461_ (.B1(\hpos[6] ),
    .Y(_0670_),
    .A2(_0628_),
    .A1(\hpos[5] ));
 sg13g2_o21ai_1 _1462_ (.B1(_0386_),
    .Y(_0671_),
    .A1(_0383_),
    .A2(_0627_));
 sg13g2_nor2_2 _1463_ (.A(_0630_),
    .B(_0670_),
    .Y(_0672_));
 sg13g2_nand2_1 _1464_ (.Y(_0673_),
    .A(_0631_),
    .B(_0671_));
 sg13g2_nand3_1 _1465_ (.B(_0631_),
    .C(_0671_),
    .A(net318),
    .Y(_0674_));
 sg13g2_a21oi_2 _1466_ (.B1(_0674_),
    .Y(_0675_),
    .A2(_0665_),
    .A1(_0663_));
 sg13g2_a21oi_1 _1467_ (.A1(_0667_),
    .A2(_0668_),
    .Y(_0676_),
    .B1(_0675_));
 sg13g2_a21o_1 _1468_ (.A2(_0668_),
    .A1(_0667_),
    .B1(_0675_),
    .X(_0677_));
 sg13g2_nor2_1 _1469_ (.A(\stage[1] ),
    .B(\stage[0] ),
    .Y(_0678_));
 sg13g2_or2_1 _1470_ (.X(_0679_),
    .B(\stage[0] ),
    .A(\stage[1] ));
 sg13g2_nor2_2 _1471_ (.A(_0392_),
    .B(_0633_),
    .Y(_0680_));
 sg13g2_o21ai_1 _1472_ (.B1(net285),
    .Y(_0681_),
    .A1(_0392_),
    .A2(_0633_));
 sg13g2_nor2_2 _1473_ (.A(\stage[0] ),
    .B(_0396_),
    .Y(_0682_));
 sg13g2_nand2_1 _1474_ (.Y(_0683_),
    .A(net292),
    .B(net285));
 sg13g2_nor2_1 _1475_ (.A(net290),
    .B(_0683_),
    .Y(_0684_));
 sg13g2_inv_1 _1476_ (.Y(_0685_),
    .A(_0684_));
 sg13g2_nor2_1 _1477_ (.A(_0682_),
    .B(_0684_),
    .Y(_0686_));
 sg13g2_nand2_1 _1478_ (.Y(_0687_),
    .A(_0633_),
    .B(net285));
 sg13g2_nor2_1 _1479_ (.A(net318),
    .B(_0673_),
    .Y(_0688_));
 sg13g2_nor4_2 _1480_ (.A(net318),
    .B(_0660_),
    .C(_0661_),
    .Y(_0689_),
    .D(_0673_));
 sg13g2_nand2_1 _1481_ (.Y(_0690_),
    .A(net290),
    .B(net285));
 sg13g2_nand2_1 _1482_ (.Y(_0691_),
    .A(_0683_),
    .B(_0690_));
 sg13g2_o21ai_1 _1483_ (.B1(_0681_),
    .Y(_0692_),
    .A1(_0682_),
    .A2(_0691_));
 sg13g2_and2_1 _1484_ (.A(_0689_),
    .B(_0692_),
    .X(_0693_));
 sg13g2_a221oi_1 _1485_ (.B2(_0686_),
    .C1(_0675_),
    .B1(_0681_),
    .A1(_0667_),
    .Y(_0694_),
    .A2(_0668_));
 sg13g2_o21ai_1 _1486_ (.B1(_0687_),
    .Y(_0695_),
    .A1(_0693_),
    .A2(_0694_));
 sg13g2_nor4_2 _1487_ (.A(_0658_),
    .B(_0662_),
    .C(_0664_),
    .Y(_0696_),
    .D(_0672_));
 sg13g2_nor2_1 _1488_ (.A(\audio_mod.pattern_clock[2] ),
    .B(_0681_),
    .Y(_0697_));
 sg13g2_nor2_1 _1489_ (.A(_0682_),
    .B(_0697_),
    .Y(_0698_));
 sg13g2_nand3_1 _1490_ (.B(_0696_),
    .C(_0698_),
    .A(_0690_),
    .Y(_0699_));
 sg13g2_nand2_1 _1491_ (.Y(_0700_),
    .A(_0658_),
    .B(_0673_));
 sg13g2_nor4_2 _1492_ (.A(_0659_),
    .B(_0660_),
    .C(_0661_),
    .Y(_0701_),
    .D(_0672_));
 sg13g2_nand3_1 _1493_ (.B(net292),
    .C(net285),
    .A(net290),
    .Y(_0702_));
 sg13g2_nand4_1 _1494_ (.B(net292),
    .C(_0679_),
    .A(net290),
    .Y(_0703_),
    .D(_0701_));
 sg13g2_nand2b_1 _1495_ (.Y(_0704_),
    .B(_0675_),
    .A_N(_0686_));
 sg13g2_nand3_1 _1496_ (.B(_0703_),
    .C(_0704_),
    .A(_0699_),
    .Y(_0705_));
 sg13g2_nor2b_2 _1497_ (.A(_0705_),
    .B_N(_0695_),
    .Y(_0706_));
 sg13g2_nand2b_2 _1498_ (.Y(_0707_),
    .B(_0695_),
    .A_N(_0705_));
 sg13g2_nor2_1 _1499_ (.A(_0395_),
    .B(net285),
    .Y(_0708_));
 sg13g2_o21ai_1 _1500_ (.B1(_0708_),
    .Y(_0709_),
    .A1(_0689_),
    .A2(_0696_));
 sg13g2_nor4_1 _1501_ (.A(_0662_),
    .B(_0664_),
    .C(_0674_),
    .D(_0702_),
    .Y(_0710_));
 sg13g2_nor3_1 _1502_ (.A(net290),
    .B(net292),
    .C(_0678_),
    .Y(_0711_));
 sg13g2_or2_1 _1503_ (.X(_0712_),
    .B(_0711_),
    .A(_0680_));
 sg13g2_a21oi_1 _1504_ (.A1(_0701_),
    .A2(_0712_),
    .Y(_0713_),
    .B1(_0710_));
 sg13g2_nand3_1 _1505_ (.B(_0709_),
    .C(_0713_),
    .A(_0677_),
    .Y(_0714_));
 sg13g2_nand2_1 _1506_ (.Y(_0715_),
    .A(_0676_),
    .B(_0697_));
 sg13g2_nand2_2 _1507_ (.Y(_0716_),
    .A(_0714_),
    .B(_0715_));
 sg13g2_nor2_2 _1508_ (.A(_0707_),
    .B(_0716_),
    .Y(_0717_));
 sg13g2_o21ai_1 _1509_ (.B1(_0683_),
    .Y(_0718_),
    .A1(_0395_),
    .A2(net285));
 sg13g2_a22oi_1 _1510_ (.Y(_0719_),
    .B1(_0718_),
    .B2(_0675_),
    .A2(_0701_),
    .A1(net285));
 sg13g2_o21ai_1 _1511_ (.B1(_0684_),
    .Y(_0720_),
    .A1(_0689_),
    .A2(_0696_));
 sg13g2_nand2b_1 _1512_ (.Y(_0721_),
    .B(_0702_),
    .A_N(_0680_));
 sg13g2_a21oi_1 _1513_ (.A1(_0689_),
    .A2(_0721_),
    .Y(_0722_),
    .B1(_0710_));
 sg13g2_nand4_1 _1514_ (.B(_0719_),
    .C(_0720_),
    .A(_0677_),
    .Y(_0723_),
    .D(_0722_));
 sg13g2_or2_1 _1515_ (.X(_0724_),
    .B(_0711_),
    .A(_0682_));
 sg13g2_o21ai_1 _1516_ (.B1(_0723_),
    .Y(_0725_),
    .A1(_0677_),
    .A2(_0724_));
 sg13g2_a22oi_1 _1517_ (.Y(_0726_),
    .B1(_0689_),
    .B2(_0691_),
    .A2(_0685_),
    .A1(_0675_));
 sg13g2_a22oi_1 _1518_ (.Y(_0727_),
    .B1(_0718_),
    .B2(_0696_),
    .A2(_0701_),
    .A1(_0698_));
 sg13g2_nand3_1 _1519_ (.B(_0726_),
    .C(_0727_),
    .A(_0677_),
    .Y(_0728_));
 sg13g2_o21ai_1 _1520_ (.B1(_0676_),
    .Y(_0729_),
    .A1(net289),
    .A2(_0678_));
 sg13g2_and2_2 _1521_ (.A(_0728_),
    .B(_0729_),
    .X(_0730_));
 sg13g2_nand2_2 _1522_ (.Y(_0731_),
    .A(_0728_),
    .B(_0729_));
 sg13g2_nor2_1 _1523_ (.A(net282),
    .B(_0730_),
    .Y(_0732_));
 sg13g2_nor3_2 _1524_ (.A(_0706_),
    .B(_0716_),
    .C(_0730_),
    .Y(_0733_));
 sg13g2_nand4_1 _1525_ (.B(_0714_),
    .C(_0715_),
    .A(_0707_),
    .Y(_0734_),
    .D(_0731_));
 sg13g2_a22oi_1 _1526_ (.Y(_0735_),
    .B1(_0733_),
    .B2(_0725_),
    .A2(_0732_),
    .A1(_0717_));
 sg13g2_nand2_1 _1527_ (.Y(_0736_),
    .A(_0666_),
    .B(_0688_));
 sg13g2_xnor2_1 _1528_ (.Y(_0737_),
    .A(_0666_),
    .B(_0688_));
 sg13g2_xnor2_1 _1529_ (.Y(_0738_),
    .A(_0389_),
    .B(_0737_));
 sg13g2_nand2_1 _1530_ (.Y(_0739_),
    .A(\hpos[9] ),
    .B(_0736_));
 sg13g2_or2_1 _1531_ (.X(_0740_),
    .B(_0736_),
    .A(net316));
 sg13g2_o21ai_1 _1532_ (.B1(_0079_),
    .Y(_0741_),
    .A1(_0630_),
    .A2(_0670_));
 sg13g2_nand3b_1 _1533_ (.B(_0631_),
    .C(_0671_),
    .Y(_0742_),
    .A_N(_0079_));
 sg13g2_and2_1 _1534_ (.A(_0741_),
    .B(_0742_),
    .X(_0743_));
 sg13g2_nand2_1 _1535_ (.Y(_0744_),
    .A(_0741_),
    .B(_0742_));
 sg13g2_and2_1 _1536_ (.A(net327),
    .B(\hvsync_gen.vpos[2] ),
    .X(_0745_));
 sg13g2_nand2_1 _1537_ (.Y(_0746_),
    .A(net327),
    .B(\hvsync_gen.vpos[2] ));
 sg13g2_nand2_2 _1538_ (.Y(_0747_),
    .A(net326),
    .B(_0745_));
 sg13g2_nand2b_1 _1539_ (.Y(_0748_),
    .B(_0646_),
    .A_N(net322));
 sg13g2_nor3_1 _1540_ (.A(_0610_),
    .B(_0646_),
    .C(_0747_),
    .Y(_0749_));
 sg13g2_o21ai_1 _1541_ (.B1(\hvsync_gen.vpos[8] ),
    .Y(_0750_),
    .A1(net323),
    .A2(_0749_));
 sg13g2_and2_1 _1542_ (.A(_0381_),
    .B(_0750_),
    .X(_0751_));
 sg13g2_and3_1 _1543_ (.X(_0752_),
    .A(\hpos[0] ),
    .B(\hpos[3] ),
    .C(net319));
 sg13g2_nor2_1 _1544_ (.A(net320),
    .B(_0615_),
    .Y(_0753_));
 sg13g2_and4_1 _1545_ (.A(_0743_),
    .B(_0751_),
    .C(_0752_),
    .D(_0753_),
    .X(_0754_));
 sg13g2_nand3_1 _1546_ (.B(_0740_),
    .C(_0754_),
    .A(_0739_),
    .Y(_0755_));
 sg13g2_or3_1 _1547_ (.A(_0735_),
    .B(_0738_),
    .C(_0755_),
    .X(_0756_));
 sg13g2_nor2_1 _1548_ (.A(net324),
    .B(net326),
    .Y(_0757_));
 sg13g2_nor3_2 _1549_ (.A(net322),
    .B(net324),
    .C(net326),
    .Y(_0758_));
 sg13g2_and2_1 _1550_ (.A(\hvsync_gen.vpos[0] ),
    .B(\hvsync_gen.vpos[1] ),
    .X(_0759_));
 sg13g2_nand2_2 _1551_ (.Y(_0760_),
    .A(\hvsync_gen.vpos[0] ),
    .B(\hvsync_gen.vpos[1] ));
 sg13g2_o21ai_1 _1552_ (.B1(net327),
    .Y(_0761_),
    .A1(\hvsync_gen.vpos[2] ),
    .A2(_0759_));
 sg13g2_a21oi_2 _1553_ (.B1(_0645_),
    .Y(_0762_),
    .A2(_0761_),
    .A1(_0758_));
 sg13g2_a21o_1 _1554_ (.A2(_0762_),
    .A1(net321),
    .B1(\hvsync_gen.vpos[9] ),
    .X(_0763_));
 sg13g2_xnor2_1 _1555_ (.Y(_0764_),
    .A(_0075_),
    .B(_0667_));
 sg13g2_nor2_1 _1556_ (.A(net317),
    .B(_0700_),
    .Y(_0765_));
 sg13g2_a21oi_1 _1557_ (.A1(_0700_),
    .A2(_0738_),
    .Y(_0766_),
    .B1(_0765_));
 sg13g2_nor3_1 _1558_ (.A(_0385_),
    .B(_0388_),
    .C(_0631_),
    .Y(_0767_));
 sg13g2_xnor2_1 _1559_ (.Y(_0768_),
    .A(net317),
    .B(_0658_));
 sg13g2_and2_1 _1560_ (.A(net320),
    .B(net319),
    .X(_0769_));
 sg13g2_o21ai_1 _1561_ (.B1(\hpos[4] ),
    .Y(_0770_),
    .A1(\hpos[3] ),
    .A2(_0769_));
 sg13g2_or2_1 _1562_ (.X(_0771_),
    .B(_0770_),
    .A(_0387_));
 sg13g2_a21oi_1 _1563_ (.A1(_0741_),
    .A2(_0742_),
    .Y(_0772_),
    .B1(_0771_));
 sg13g2_mux2_1 _1564_ (.A0(_0078_),
    .A1(_0079_),
    .S(_0629_),
    .X(_0773_));
 sg13g2_inv_1 _1565_ (.Y(_0774_),
    .A(_0773_));
 sg13g2_nor2_1 _1566_ (.A(_0772_),
    .B(_0774_),
    .Y(_0775_));
 sg13g2_o21ai_1 _1567_ (.B1(_0768_),
    .Y(_0776_),
    .A1(_0772_),
    .A2(_0774_));
 sg13g2_a21oi_1 _1568_ (.A1(\hpos[8] ),
    .A2(_0669_),
    .Y(_0777_),
    .B1(_0767_));
 sg13g2_nand2_1 _1569_ (.Y(_0778_),
    .A(_0776_),
    .B(_0777_));
 sg13g2_xor2_1 _1570_ (.B(_0778_),
    .A(_0764_),
    .X(_0779_));
 sg13g2_nor2_1 _1571_ (.A(_0069_),
    .B(_0650_),
    .Y(_0780_));
 sg13g2_xor2_1 _1572_ (.B(_0780_),
    .A(_0068_),
    .X(_0781_));
 sg13g2_xnor2_1 _1573_ (.Y(_0782_),
    .A(_0779_),
    .B(_0781_));
 sg13g2_nand3_1 _1574_ (.B(\hpos[4] ),
    .C(_0638_),
    .A(net320),
    .Y(_0783_));
 sg13g2_nor3_1 _1575_ (.A(\hpos[0] ),
    .B(\hpos[5] ),
    .C(_0783_),
    .Y(_0784_));
 sg13g2_and3_1 _1576_ (.X(_0785_),
    .A(_0764_),
    .B(_0766_),
    .C(_0784_));
 sg13g2_nand2_1 _1577_ (.Y(_0786_),
    .A(_0744_),
    .B(_0785_));
 sg13g2_a22oi_1 _1578_ (.Y(_0787_),
    .B1(_0764_),
    .B2(_0778_),
    .A2(_0667_),
    .A1(net316));
 sg13g2_a21oi_1 _1579_ (.A1(_0744_),
    .A2(_0785_),
    .Y(_0788_),
    .B1(_0787_));
 sg13g2_xor2_1 _1580_ (.B(_0736_),
    .A(_0075_),
    .X(_0789_));
 sg13g2_inv_1 _1581_ (.Y(_0790_),
    .A(_0789_));
 sg13g2_xnor2_1 _1582_ (.Y(_0791_),
    .A(_0672_),
    .B(_0768_));
 sg13g2_nand2_1 _1583_ (.Y(_0792_),
    .A(_0629_),
    .B(_0791_));
 sg13g2_nor3_1 _1584_ (.A(_0639_),
    .B(_0789_),
    .C(_0792_),
    .Y(_0793_));
 sg13g2_inv_1 _1585_ (.Y(_0794_),
    .A(_0793_));
 sg13g2_o21ai_1 _1586_ (.B1(_0670_),
    .Y(_0795_),
    .A1(_0385_),
    .A2(net317));
 sg13g2_nand2_1 _1587_ (.Y(_0796_),
    .A(_0387_),
    .B(_0639_));
 sg13g2_nand3_1 _1588_ (.B(_0791_),
    .C(_0796_),
    .A(_0629_),
    .Y(_0797_));
 sg13g2_a21oi_1 _1589_ (.A1(_0795_),
    .A2(_0797_),
    .Y(_0798_),
    .B1(_0738_));
 sg13g2_nor2_1 _1590_ (.A(\hpos[8] ),
    .B(_0737_),
    .Y(_0799_));
 sg13g2_nor2_1 _1591_ (.A(_0798_),
    .B(_0799_),
    .Y(_0800_));
 sg13g2_o21ai_1 _1592_ (.B1(_0790_),
    .Y(_0801_),
    .A1(_0798_),
    .A2(_0799_));
 sg13g2_nand2_1 _1593_ (.Y(_0802_),
    .A(_0740_),
    .B(_0801_));
 sg13g2_a21oi_1 _1594_ (.A1(_0740_),
    .A2(_0801_),
    .Y(_0803_),
    .B1(_0793_));
 sg13g2_or2_1 _1595_ (.X(_0804_),
    .B(_0803_),
    .A(_0788_));
 sg13g2_nor3_1 _1596_ (.A(_0782_),
    .B(_0788_),
    .C(_0803_),
    .Y(_0805_));
 sg13g2_and2_1 _1597_ (.A(_0652_),
    .B(_0787_),
    .X(_0806_));
 sg13g2_nor2_1 _1598_ (.A(_0652_),
    .B(_0787_),
    .Y(_0807_));
 sg13g2_xnor2_1 _1599_ (.Y(_0808_),
    .A(_0768_),
    .B(_0775_));
 sg13g2_nand2_1 _1600_ (.Y(_0809_),
    .A(_0067_),
    .B(_0649_));
 sg13g2_xnor2_1 _1601_ (.Y(_0810_),
    .A(net322),
    .B(_0809_));
 sg13g2_xnor2_1 _1602_ (.Y(_0811_),
    .A(_0808_),
    .B(_0810_));
 sg13g2_xnor2_1 _1603_ (.Y(_0812_),
    .A(_0067_),
    .B(_0649_));
 sg13g2_nand2_1 _1604_ (.Y(_0813_),
    .A(_0078_),
    .B(_0770_));
 sg13g2_xnor2_1 _1605_ (.Y(_0814_),
    .A(_0743_),
    .B(_0813_));
 sg13g2_xor2_1 _1606_ (.B(\hpos[2] ),
    .A(\hpos[1] ),
    .X(_0815_));
 sg13g2_xnor2_1 _1607_ (.Y(_0816_),
    .A(\hvsync_gen.vpos[2] ),
    .B(_0646_));
 sg13g2_xor2_1 _1608_ (.B(net320),
    .A(\hvsync_gen.vpos[1] ),
    .X(_0817_));
 sg13g2_and2_1 _1609_ (.A(\hvsync_gen.vpos[0] ),
    .B(\hpos[0] ),
    .X(_0818_));
 sg13g2_nor2_1 _1610_ (.A(\hvsync_gen.vpos[0] ),
    .B(\hpos[0] ),
    .Y(_0819_));
 sg13g2_mux2_1 _1611_ (.A0(_0818_),
    .A1(_0819_),
    .S(_0817_),
    .X(_0820_));
 sg13g2_xnor2_1 _1612_ (.Y(_0821_),
    .A(_0815_),
    .B(_0816_));
 sg13g2_xnor2_1 _1613_ (.Y(_0822_),
    .A(\hpos[3] ),
    .B(_0769_));
 sg13g2_xor2_1 _1614_ (.B(_0647_),
    .A(_0066_),
    .X(_0823_));
 sg13g2_xnor2_1 _1615_ (.Y(_0824_),
    .A(_0822_),
    .B(_0823_));
 sg13g2_a21o_1 _1616_ (.A2(_0647_),
    .A1(net327),
    .B1(net326),
    .X(_0825_));
 sg13g2_nand2_1 _1617_ (.Y(_0826_),
    .A(_0648_),
    .B(_0825_));
 sg13g2_nand2b_1 _1618_ (.Y(_0827_),
    .B(_0076_),
    .A_N(_0769_));
 sg13g2_xnor2_1 _1619_ (.Y(_0828_),
    .A(_0384_),
    .B(_0827_));
 sg13g2_xnor2_1 _1620_ (.Y(_0829_),
    .A(_0826_),
    .B(_0828_));
 sg13g2_nand4_1 _1621_ (.B(_0821_),
    .C(_0824_),
    .A(_0820_),
    .Y(_0830_),
    .D(_0829_));
 sg13g2_xor2_1 _1622_ (.B(_0078_),
    .A(net325),
    .X(_0831_));
 sg13g2_xnor2_1 _1623_ (.Y(_0832_),
    .A(_0770_),
    .B(_0831_));
 sg13g2_xnor2_1 _1624_ (.Y(_0833_),
    .A(_0648_),
    .B(_0832_));
 sg13g2_xnor2_1 _1625_ (.Y(_0834_),
    .A(_0812_),
    .B(_0814_));
 sg13g2_nor4_1 _1626_ (.A(_0811_),
    .B(_0830_),
    .C(_0833_),
    .D(_0834_),
    .Y(_0835_));
 sg13g2_o21ai_1 _1627_ (.B1(_0776_),
    .Y(_0836_),
    .A1(_0385_),
    .A2(_0631_));
 sg13g2_xnor2_1 _1628_ (.Y(_0837_),
    .A(net321),
    .B(_0650_));
 sg13g2_xnor2_1 _1629_ (.Y(_0838_),
    .A(_0836_),
    .B(_0837_));
 sg13g2_and2_1 _1630_ (.A(net282),
    .B(_0730_),
    .X(_0839_));
 sg13g2_nand2_1 _1631_ (.Y(_0840_),
    .A(_0706_),
    .B(_0716_));
 sg13g2_nand4_1 _1632_ (.B(_0716_),
    .C(net282),
    .A(_0706_),
    .Y(_0841_),
    .D(_0730_));
 sg13g2_and2_1 _1633_ (.A(_0725_),
    .B(_0731_),
    .X(_0842_));
 sg13g2_nand2_1 _1634_ (.Y(_0843_),
    .A(net282),
    .B(_0731_));
 sg13g2_and2_1 _1635_ (.A(_0707_),
    .B(_0716_),
    .X(_0844_));
 sg13g2_nand4_1 _1636_ (.B(_0716_),
    .C(net282),
    .A(_0707_),
    .Y(_0845_),
    .D(_0731_));
 sg13g2_nor2_1 _1637_ (.A(_0725_),
    .B(_0731_),
    .Y(_0846_));
 sg13g2_nand2b_1 _1638_ (.Y(_0847_),
    .B(_0730_),
    .A_N(net282));
 sg13g2_or3_1 _1639_ (.A(_0716_),
    .B(net282),
    .C(_0731_),
    .X(_0848_));
 sg13g2_and4_1 _1640_ (.A(_0734_),
    .B(_0841_),
    .C(_0845_),
    .D(_0848_),
    .X(_0849_));
 sg13g2_a21oi_1 _1641_ (.A1(_0717_),
    .A2(_0842_),
    .Y(_0850_),
    .B1(_0844_));
 sg13g2_a22oi_1 _1642_ (.Y(_0851_),
    .B1(_0844_),
    .B2(_0846_),
    .A2(_0842_),
    .A1(_0717_));
 sg13g2_a21oi_1 _1643_ (.A1(_0849_),
    .A2(_0851_),
    .Y(_0852_),
    .B1(_0786_));
 sg13g2_nor2_1 _1644_ (.A(_0840_),
    .B(_0843_),
    .Y(_0853_));
 sg13g2_nor2_1 _1645_ (.A(_0794_),
    .B(_0853_),
    .Y(_0854_));
 sg13g2_nand3b_1 _1646_ (.B(\hvsync_gen.vpos[6] ),
    .C(_0758_),
    .Y(_0855_),
    .A_N(\hvsync_gen.vpos[0] ));
 sg13g2_nor2_1 _1647_ (.A(_0609_),
    .B(_0855_),
    .Y(_0856_));
 sg13g2_nand3_1 _1648_ (.B(_0716_),
    .C(_0730_),
    .A(_0706_),
    .Y(_0857_));
 sg13g2_nand2_1 _1649_ (.Y(_0858_),
    .A(_0717_),
    .B(_0839_));
 sg13g2_nand4_1 _1650_ (.B(_0851_),
    .C(_0857_),
    .A(_0845_),
    .Y(_0859_),
    .D(_0858_));
 sg13g2_nand2_1 _1651_ (.Y(_0860_),
    .A(_0856_),
    .B(_0859_));
 sg13g2_nor4_1 _1652_ (.A(_0607_),
    .B(_0610_),
    .C(_0747_),
    .D(_0748_),
    .Y(_0861_));
 sg13g2_a221oi_1 _1653_ (.B2(_0717_),
    .C1(_0733_),
    .B1(_0839_),
    .A1(_0675_),
    .Y(_0862_),
    .A2(_0718_));
 sg13g2_o21ai_1 _1654_ (.B1(_0862_),
    .Y(_0863_),
    .A1(net282),
    .A2(_0840_));
 sg13g2_nor2_1 _1655_ (.A(_0654_),
    .B(_0853_),
    .Y(_0864_));
 sg13g2_nand2_1 _1656_ (.Y(_0865_),
    .A(_0707_),
    .B(_0847_));
 sg13g2_a21o_1 _1657_ (.A2(_0865_),
    .A1(_0848_),
    .B1(_0733_),
    .X(_0866_));
 sg13g2_a22oi_1 _1658_ (.Y(_0867_),
    .B1(_0864_),
    .B2(_0866_),
    .A2(_0863_),
    .A1(_0861_));
 sg13g2_a21oi_1 _1659_ (.A1(_0860_),
    .A2(_0867_),
    .Y(_0868_),
    .B1(_0804_));
 sg13g2_or2_1 _1660_ (.X(_0869_),
    .B(_0856_),
    .A(_0763_));
 sg13g2_a21oi_1 _1661_ (.A1(_0849_),
    .A2(_0858_),
    .Y(_0870_),
    .B1(_0786_));
 sg13g2_nand2b_1 _1662_ (.Y(_0871_),
    .B(_0843_),
    .A_N(_0717_));
 sg13g2_a21oi_1 _1663_ (.A1(_0850_),
    .A2(_0871_),
    .Y(_0872_),
    .B1(_0794_));
 sg13g2_o21ai_1 _1664_ (.B1(_0869_),
    .Y(_0873_),
    .A1(_0870_),
    .A2(_0872_));
 sg13g2_xnor2_1 _1665_ (.Y(_0874_),
    .A(_0789_),
    .B(_0800_));
 sg13g2_nand2b_1 _1666_ (.Y(_0875_),
    .B(_0762_),
    .A_N(_0069_));
 sg13g2_xnor2_1 _1667_ (.Y(_0876_),
    .A(_0068_),
    .B(_0875_));
 sg13g2_xnor2_1 _1668_ (.Y(_0877_),
    .A(_0874_),
    .B(_0876_));
 sg13g2_nand3_1 _1669_ (.B(_0795_),
    .C(_0797_),
    .A(_0738_),
    .Y(_0878_));
 sg13g2_nand2b_1 _1670_ (.Y(_0879_),
    .B(_0878_),
    .A_N(_0798_));
 sg13g2_xor2_1 _1671_ (.B(_0762_),
    .A(net321),
    .X(_0880_));
 sg13g2_a21oi_1 _1672_ (.A1(_0757_),
    .A2(_0761_),
    .Y(_0881_),
    .B1(_0067_));
 sg13g2_nand2_1 _1673_ (.Y(_0882_),
    .A(_0639_),
    .B(_0671_));
 sg13g2_xor2_1 _1674_ (.B(_0882_),
    .A(net323),
    .X(_0883_));
 sg13g2_xnor2_1 _1675_ (.Y(_0884_),
    .A(_0881_),
    .B(_0883_));
 sg13g2_nand2_1 _1676_ (.Y(_0885_),
    .A(_0077_),
    .B(_0641_));
 sg13g2_nand2_1 _1677_ (.Y(_0886_),
    .A(_0071_),
    .B(_0761_));
 sg13g2_xor2_1 _1678_ (.B(_0886_),
    .A(_0831_),
    .X(_0887_));
 sg13g2_nand3_1 _1679_ (.B(_0757_),
    .C(_0761_),
    .A(_0067_),
    .Y(_0888_));
 sg13g2_nor2b_1 _1680_ (.A(_0881_),
    .B_N(_0888_),
    .Y(_0889_));
 sg13g2_xnor2_1 _1681_ (.Y(_0890_),
    .A(_0077_),
    .B(_0641_));
 sg13g2_xor2_1 _1682_ (.B(_0761_),
    .A(_0071_),
    .X(_0891_));
 sg13g2_xnor2_1 _1683_ (.Y(_0892_),
    .A(_0890_),
    .B(_0891_));
 sg13g2_nand2_1 _1684_ (.Y(_0893_),
    .A(_0070_),
    .B(_0760_));
 sg13g2_xnor2_1 _1685_ (.Y(_0894_),
    .A(_0070_),
    .B(_0760_));
 sg13g2_xnor2_1 _1686_ (.Y(_0895_),
    .A(net319),
    .B(_0636_));
 sg13g2_nor2_1 _1687_ (.A(_0818_),
    .B(_0819_),
    .Y(_0896_));
 sg13g2_xnor2_1 _1688_ (.Y(_0897_),
    .A(_0076_),
    .B(_0640_));
 sg13g2_xor2_1 _1689_ (.B(_0893_),
    .A(_0066_),
    .X(_0898_));
 sg13g2_xnor2_1 _1690_ (.Y(_0899_),
    .A(_0894_),
    .B(_0895_));
 sg13g2_o21ai_1 _1691_ (.B1(_0899_),
    .Y(_0900_),
    .A1(_0897_),
    .A2(_0898_));
 sg13g2_a21oi_1 _1692_ (.A1(_0897_),
    .A2(_0898_),
    .Y(_0901_),
    .B1(_0896_));
 sg13g2_nand2_1 _1693_ (.Y(_0902_),
    .A(_0817_),
    .B(_0901_));
 sg13g2_mux2_1 _1694_ (.A0(_0717_),
    .A1(_0844_),
    .S(_0839_),
    .X(_0903_));
 sg13g2_nor2_2 _1695_ (.A(\lfsr[2] ),
    .B(\lfsr[1] ),
    .Y(_0904_));
 sg13g2_xor2_1 _1696_ (.B(_0802_),
    .A(_0763_),
    .X(_0905_));
 sg13g2_nand2_1 _1697_ (.Y(_0906_),
    .A(_0791_),
    .B(_0884_));
 sg13g2_nor2_1 _1698_ (.A(_0791_),
    .B(_0884_),
    .Y(_0907_));
 sg13g2_xnor2_1 _1699_ (.Y(_0908_),
    .A(_0885_),
    .B(_0887_));
 sg13g2_xnor2_1 _1700_ (.Y(_0909_),
    .A(_0639_),
    .B(_0889_));
 sg13g2_xnor2_1 _1701_ (.Y(_0910_),
    .A(_0879_),
    .B(_0880_));
 sg13g2_xnor2_1 _1702_ (.Y(_0911_),
    .A(_0766_),
    .B(_0838_));
 sg13g2_nand4_1 _1703_ (.B(_0835_),
    .C(_0839_),
    .A(_0707_),
    .Y(_0912_),
    .D(_0911_));
 sg13g2_nor3_1 _1704_ (.A(_0806_),
    .B(_0807_),
    .C(_0912_),
    .Y(_0913_));
 sg13g2_a221oi_1 _1705_ (.B2(_0805_),
    .C1(_0852_),
    .B1(_0913_),
    .A1(_0735_),
    .Y(_0914_),
    .A2(_0854_));
 sg13g2_o21ai_1 _1706_ (.B1(_0756_),
    .Y(_0915_),
    .A1(_0763_),
    .A2(_0914_));
 sg13g2_nor4_1 _1707_ (.A(_0892_),
    .B(_0900_),
    .C(_0902_),
    .D(_0909_),
    .Y(_0916_));
 sg13g2_nand4_1 _1708_ (.B(_0906_),
    .C(_0908_),
    .A(_0869_),
    .Y(_0917_),
    .D(_0916_));
 sg13g2_nor3_1 _1709_ (.A(_0732_),
    .B(_0907_),
    .C(_0917_),
    .Y(_0918_));
 sg13g2_nand4_1 _1710_ (.B(_0905_),
    .C(_0910_),
    .A(_0877_),
    .Y(_0919_),
    .D(_0918_));
 sg13g2_nand2b_1 _1711_ (.Y(_0920_),
    .B(_0903_),
    .A_N(_0804_));
 sg13g2_o21ai_1 _1712_ (.B1(_0873_),
    .Y(_0921_),
    .A1(_0919_),
    .A2(_0920_));
 sg13g2_a221oi_1 _1713_ (.B2(_0751_),
    .C1(_0868_),
    .B1(_0921_),
    .A1(_0655_),
    .Y(_0922_),
    .A2(_0915_));
 sg13g2_nor3_1 _1714_ (.A(_0635_),
    .B(_0644_),
    .C(_0922_),
    .Y(_0923_));
 sg13g2_nor4_1 _1715_ (.A(_0626_),
    .B(_0635_),
    .C(_0644_),
    .D(_0922_),
    .Y(_0924_));
 sg13g2_nor4_2 _1716_ (.A(_0635_),
    .B(_0644_),
    .C(_0904_),
    .Y(_0925_),
    .D(_0922_));
 sg13g2_nor4_2 _1717_ (.A(_0635_),
    .B(_0644_),
    .C(_0680_),
    .Y(_0926_),
    .D(_0922_));
 sg13g2_nand4_1 _1718_ (.B(_0680_),
    .C(_0904_),
    .A(_0625_),
    .Y(_0927_),
    .D(_0923_));
 sg13g2_nand2_1 _1719_ (.Y(_0928_),
    .A(_0624_),
    .B(_0927_));
 sg13g2_xor2_1 _1720_ (.B(net317),
    .A(\counter[5] ),
    .X(_0929_));
 sg13g2_xnor2_1 _1721_ (.Y(_0930_),
    .A(\hvsync_gen.vpos[7] ),
    .B(_0929_));
 sg13g2_xor2_1 _1722_ (.B(_0081_),
    .A(net321),
    .X(_0931_));
 sg13g2_xor2_1 _1723_ (.B(_0931_),
    .A(\counter[6] ),
    .X(_0932_));
 sg13g2_xor2_1 _1724_ (.B(_0831_),
    .A(net303),
    .X(_0933_));
 sg13g2_xnor2_1 _1725_ (.Y(_0934_),
    .A(net319),
    .B(\counter[0] ));
 sg13g2_xnor2_1 _1726_ (.Y(_0935_),
    .A(\hvsync_gen.vpos[2] ),
    .B(_0934_));
 sg13g2_xor2_1 _1727_ (.B(_0076_),
    .A(net327),
    .X(_0936_));
 sg13g2_xnor2_1 _1728_ (.Y(_0937_),
    .A(net306),
    .B(_0936_));
 sg13g2_xnor2_1 _1729_ (.Y(_0938_),
    .A(net326),
    .B(net304));
 sg13g2_xnor2_1 _1730_ (.Y(_0939_),
    .A(_0077_),
    .B(_0938_));
 sg13g2_xnor2_1 _1731_ (.Y(_0940_),
    .A(\hvsync_gen.vpos[6] ),
    .B(_0079_));
 sg13g2_xnor2_1 _1732_ (.Y(_0941_),
    .A(\counter[4] ),
    .B(_0940_));
 sg13g2_nand4_1 _1733_ (.B(_0933_),
    .C(_0939_),
    .A(_0932_),
    .Y(_0942_),
    .D(_0941_));
 sg13g2_nor4_1 _1734_ (.A(_0930_),
    .B(_0935_),
    .C(_0937_),
    .D(_0942_),
    .Y(_0943_));
 sg13g2_nor2_1 _1735_ (.A(net306),
    .B(net305),
    .Y(_0944_));
 sg13g2_xnor2_1 _1736_ (.Y(_0945_),
    .A(net325),
    .B(_0082_));
 sg13g2_xnor2_1 _1737_ (.Y(_0946_),
    .A(_0082_),
    .B(_0831_));
 sg13g2_xor2_1 _1738_ (.B(_0940_),
    .A(_0083_),
    .X(_0947_));
 sg13g2_nor2b_1 _1739_ (.A(\counter[3] ),
    .B_N(_0947_),
    .Y(_0948_));
 sg13g2_nor2_1 _1740_ (.A(net303),
    .B(\counter[4] ),
    .Y(_0949_));
 sg13g2_nand2b_1 _1741_ (.Y(_0950_),
    .B(_0949_),
    .A_N(\counter[5] ));
 sg13g2_xor2_1 _1742_ (.B(_0931_),
    .A(_0061_),
    .X(_0951_));
 sg13g2_a21oi_1 _1743_ (.A1(\counter[6] ),
    .A2(_0951_),
    .Y(_0952_),
    .B1(_0950_));
 sg13g2_xor2_1 _1744_ (.B(_0084_),
    .A(net317),
    .X(_0953_));
 sg13g2_xnor2_1 _1745_ (.Y(_0954_),
    .A(\hvsync_gen.vpos[7] ),
    .B(_0953_));
 sg13g2_and2_1 _1746_ (.A(_0949_),
    .B(_0954_),
    .X(_0955_));
 sg13g2_or3_1 _1747_ (.A(_0948_),
    .B(_0952_),
    .C(_0955_),
    .X(_0956_));
 sg13g2_nor4_1 _1748_ (.A(_0946_),
    .B(_0948_),
    .C(_0952_),
    .D(_0955_),
    .Y(_0957_));
 sg13g2_nor2b_1 _1749_ (.A(_0957_),
    .B_N(_0944_),
    .Y(_0958_));
 sg13g2_nor2b_1 _1750_ (.A(_0951_),
    .B_N(_0954_),
    .Y(_0959_));
 sg13g2_a21oi_1 _1751_ (.A1(_0946_),
    .A2(_0959_),
    .Y(_0960_),
    .B1(_0944_));
 sg13g2_nand2_1 _1752_ (.Y(_0961_),
    .A(_0950_),
    .B(_0951_));
 sg13g2_nor2_1 _1753_ (.A(net304),
    .B(net303),
    .Y(_0962_));
 sg13g2_nor2_1 _1754_ (.A(net296),
    .B(_0962_),
    .Y(_0963_));
 sg13g2_nor3_1 _1755_ (.A(net306),
    .B(net305),
    .C(net303),
    .Y(_0964_));
 sg13g2_o21ai_1 _1756_ (.B1(_0961_),
    .Y(_0965_),
    .A1(net296),
    .A2(_0964_));
 sg13g2_o21ai_1 _1757_ (.B1(_0937_),
    .Y(_0966_),
    .A1(_0949_),
    .A2(net295));
 sg13g2_nor2_1 _1758_ (.A(_0935_),
    .B(_0966_),
    .Y(_0967_));
 sg13g2_xnor2_1 _1759_ (.Y(_0968_),
    .A(\counter[1] ),
    .B(_0939_));
 sg13g2_nand2_1 _1760_ (.Y(_0969_),
    .A(_0967_),
    .B(_0968_));
 sg13g2_nor4_2 _1761_ (.A(_0958_),
    .B(_0960_),
    .C(_0965_),
    .Y(_0970_),
    .D(_0969_));
 sg13g2_nor2_1 _1762_ (.A(_0943_),
    .B(_0970_),
    .Y(_0971_));
 sg13g2_nor3_2 _1763_ (.A(net304),
    .B(net303),
    .C(\counter[4] ),
    .Y(_0972_));
 sg13g2_nor2_1 _1764_ (.A(\counter[5] ),
    .B(\counter[6] ),
    .Y(_0973_));
 sg13g2_a22oi_1 _1765_ (.Y(_0974_),
    .B1(_0972_),
    .B2(_0973_),
    .A2(_0962_),
    .A1(net296));
 sg13g2_a21oi_1 _1766_ (.A1(net295),
    .A2(_0972_),
    .Y(_0975_),
    .B1(net297));
 sg13g2_a21oi_1 _1767_ (.A1(_0974_),
    .A2(_0975_),
    .Y(_0976_),
    .B1(_0939_));
 sg13g2_nand2b_1 _1768_ (.Y(_0977_),
    .B(_0062_),
    .A_N(_0619_));
 sg13g2_xnor2_1 _1769_ (.Y(_0978_),
    .A(_0946_),
    .B(_0977_));
 sg13g2_nor2_1 _1770_ (.A(net295),
    .B(_0972_),
    .Y(_0979_));
 sg13g2_nor2_1 _1771_ (.A(_0963_),
    .B(_0979_),
    .Y(_0980_));
 sg13g2_nor3_1 _1772_ (.A(net304),
    .B(net297),
    .C(_0950_),
    .Y(_0981_));
 sg13g2_xnor2_1 _1773_ (.Y(_0982_),
    .A(_0951_),
    .B(_0981_));
 sg13g2_nand3_1 _1774_ (.B(net296),
    .C(net295),
    .A(net297),
    .Y(_0983_));
 sg13g2_xnor2_1 _1775_ (.Y(_0984_),
    .A(\counter[0] ),
    .B(_0937_));
 sg13g2_nand2_1 _1776_ (.Y(_0985_),
    .A(_0935_),
    .B(_0984_));
 sg13g2_a21oi_1 _1777_ (.A1(_0939_),
    .A2(_0983_),
    .Y(_0986_),
    .B1(_0985_));
 sg13g2_nand4_1 _1778_ (.B(_0980_),
    .C(_0982_),
    .A(_0978_),
    .Y(_0987_),
    .D(_0986_));
 sg13g2_nor2_2 _1779_ (.A(\counter[0] ),
    .B(net306),
    .Y(_0988_));
 sg13g2_nor3_2 _1780_ (.A(\counter[0] ),
    .B(net306),
    .C(net304),
    .Y(_0989_));
 sg13g2_nor2b_1 _1781_ (.A(_0984_),
    .B_N(_0935_),
    .Y(_0990_));
 sg13g2_nor2_1 _1782_ (.A(net296),
    .B(_0988_),
    .Y(_0991_));
 sg13g2_a21oi_1 _1783_ (.A1(_0972_),
    .A2(_0988_),
    .Y(_0992_),
    .B1(net295));
 sg13g2_xor2_1 _1784_ (.B(_0988_),
    .A(_0077_),
    .X(_0993_));
 sg13g2_xnor2_1 _1785_ (.Y(_0994_),
    .A(net326),
    .B(_0062_));
 sg13g2_xnor2_1 _1786_ (.Y(_0995_),
    .A(_0993_),
    .B(_0994_));
 sg13g2_nor3_1 _1787_ (.A(_0991_),
    .B(_0992_),
    .C(_0995_),
    .Y(_0996_));
 sg13g2_nand2b_1 _1788_ (.Y(_0997_),
    .B(_0989_),
    .A_N(_0950_));
 sg13g2_a21oi_1 _1789_ (.A1(_0951_),
    .A2(_0997_),
    .Y(_0998_),
    .B1(_0963_));
 sg13g2_xnor2_1 _1790_ (.Y(_0999_),
    .A(_0945_),
    .B(_0989_));
 sg13g2_xnor2_1 _1791_ (.Y(_1000_),
    .A(_0078_),
    .B(_0999_));
 sg13g2_nand4_1 _1792_ (.B(_0996_),
    .C(_0998_),
    .A(_0990_),
    .Y(_1001_),
    .D(_1000_));
 sg13g2_a21oi_1 _1793_ (.A1(_0956_),
    .A2(_0989_),
    .Y(_1002_),
    .B1(_1001_));
 sg13g2_o21ai_1 _1794_ (.B1(_0971_),
    .Y(_1003_),
    .A1(_0976_),
    .A2(_0987_));
 sg13g2_nor2_1 _1795_ (.A(_1002_),
    .B(_1003_),
    .Y(_1004_));
 sg13g2_nor3_1 _1796_ (.A(_0935_),
    .B(_0937_),
    .C(_0939_),
    .Y(_1005_));
 sg13g2_nor2_1 _1797_ (.A(_0933_),
    .B(_0955_),
    .Y(_1006_));
 sg13g2_nor2_1 _1798_ (.A(\counter[5] ),
    .B(net295),
    .Y(_1007_));
 sg13g2_xnor2_1 _1799_ (.Y(_1008_),
    .A(_0951_),
    .B(_1007_));
 sg13g2_mux2_1 _1800_ (.A0(_1006_),
    .A1(_0933_),
    .S(net304),
    .X(_1009_));
 sg13g2_and3_1 _1801_ (.X(_1010_),
    .A(_0974_),
    .B(_0980_),
    .C(_1005_));
 sg13g2_nand3_1 _1802_ (.B(_1009_),
    .C(_1010_),
    .A(_1008_),
    .Y(_1011_));
 sg13g2_nor2b_1 _1803_ (.A(_0943_),
    .B_N(_1011_),
    .Y(_1012_));
 sg13g2_nor2b_1 _1804_ (.A(_1002_),
    .B_N(_1012_),
    .Y(_1013_));
 sg13g2_o21ai_1 _1805_ (.B1(net304),
    .Y(_1014_),
    .A1(\counter[0] ),
    .A2(net306));
 sg13g2_o21ai_1 _1806_ (.B1(_0082_),
    .Y(_1015_),
    .A1(net303),
    .A2(_1014_));
 sg13g2_nor2_1 _1807_ (.A(\counter[4] ),
    .B(_1015_),
    .Y(_1016_));
 sg13g2_o21ai_1 _1808_ (.B1(_1016_),
    .Y(_1017_),
    .A1(net295),
    .A2(_0973_));
 sg13g2_nor2_1 _1809_ (.A(net295),
    .B(_1016_),
    .Y(_1018_));
 sg13g2_xor2_1 _1810_ (.B(_1015_),
    .A(net296),
    .X(_1019_));
 sg13g2_xnor2_1 _1811_ (.Y(_1020_),
    .A(_0933_),
    .B(_1014_));
 sg13g2_xnor2_1 _1812_ (.Y(_1021_),
    .A(_0939_),
    .B(_0988_));
 sg13g2_nand4_1 _1813_ (.B(_1008_),
    .C(_1017_),
    .A(_0990_),
    .Y(_1022_),
    .D(_1021_));
 sg13g2_nor4_1 _1814_ (.A(_1018_),
    .B(_1019_),
    .C(_1020_),
    .D(_1022_),
    .Y(_1023_));
 sg13g2_nor2b_1 _1815_ (.A(_1023_),
    .B_N(_1013_),
    .Y(_1024_));
 sg13g2_nand2_1 _1816_ (.Y(_1025_),
    .A(_0082_),
    .B(net296));
 sg13g2_nand3_1 _1817_ (.B(_1006_),
    .C(_1025_),
    .A(_0961_),
    .Y(_1026_));
 sg13g2_o21ai_1 _1818_ (.B1(_0620_),
    .Y(_1027_),
    .A1(_0952_),
    .A2(_1026_));
 sg13g2_a21o_1 _1819_ (.A2(_0959_),
    .A1(_0933_),
    .B1(_0620_),
    .X(_1028_));
 sg13g2_a21oi_1 _1820_ (.A1(_0082_),
    .A2(_0620_),
    .Y(_1029_),
    .B1(net296));
 sg13g2_nor2_1 _1821_ (.A(_0968_),
    .B(_1029_),
    .Y(_1030_));
 sg13g2_nand4_1 _1822_ (.B(_1027_),
    .C(_1028_),
    .A(_0967_),
    .Y(_1031_),
    .D(_1030_));
 sg13g2_and2_1 _1823_ (.A(_0971_),
    .B(_1031_),
    .X(_1032_));
 sg13g2_nand2b_1 _1824_ (.Y(_1033_),
    .B(_0625_),
    .A_N(_1032_));
 sg13g2_nand3_1 _1825_ (.B(_1011_),
    .C(_1032_),
    .A(\bright[2][0] ),
    .Y(_1034_));
 sg13g2_mux2_1 _1826_ (.A0(_1034_),
    .A1(_1033_),
    .S(_1024_),
    .X(_1035_));
 sg13g2_nor2b_1 _1827_ (.A(_1035_),
    .B_N(_1004_),
    .Y(_0193_));
 sg13g2_a21oi_1 _1828_ (.A1(_0971_),
    .A2(_1012_),
    .Y(_0194_),
    .B1(_0904_));
 sg13g2_a21oi_1 _1829_ (.A1(_0985_),
    .A2(_1012_),
    .Y(_0195_),
    .B1(_1004_));
 sg13g2_nor3_2 _1830_ (.A(_0193_),
    .B(_0194_),
    .C(_0195_),
    .Y(_0196_));
 sg13g2_and3_1 _1831_ (.X(_0197_),
    .A(_0063_),
    .B(_0065_),
    .C(_0391_));
 sg13g2_nor2_1 _1832_ (.A(_0065_),
    .B(_0392_),
    .Y(_0198_));
 sg13g2_a21o_1 _1833_ (.A2(_0198_),
    .A1(_0064_),
    .B1(_0197_),
    .X(_0199_));
 sg13g2_nand2b_1 _1834_ (.Y(_0200_),
    .B(_0199_),
    .A_N(_0196_));
 sg13g2_nand2b_1 _1835_ (.Y(_0201_),
    .B(\background_color[0] ),
    .A_N(\background_color[1] ));
 sg13g2_nand2_1 _1836_ (.Y(_0202_),
    .A(\background_color[2] ),
    .B(\background_color[1] ));
 sg13g2_nand2_1 _1837_ (.Y(_0203_),
    .A(_0201_),
    .B(_0202_));
 sg13g2_a21oi_2 _1838_ (.B1(_1004_),
    .Y(_0204_),
    .A2(_1033_),
    .A1(_1013_));
 sg13g2_o21ai_1 _1839_ (.B1(_0679_),
    .Y(_0205_),
    .A1(_0065_),
    .A2(_0392_));
 sg13g2_o21ai_1 _1840_ (.B1(_0205_),
    .Y(_0206_),
    .A1(_0390_),
    .A2(_0392_));
 sg13g2_nand2_1 _1841_ (.Y(_0207_),
    .A(_0064_),
    .B(_0391_));
 sg13g2_inv_1 _1842_ (.Y(_0208_),
    .A(_0207_));
 sg13g2_o21ai_1 _1843_ (.B1(_0206_),
    .Y(_0209_),
    .A1(_0197_),
    .A2(_0207_));
 sg13g2_nor2b_1 _1844_ (.A(_0209_),
    .B_N(_0204_),
    .Y(_0210_));
 sg13g2_nand2_1 _1845_ (.Y(_0211_),
    .A(_0199_),
    .B(_0204_));
 sg13g2_o21ai_1 _1846_ (.B1(_0206_),
    .Y(_0212_),
    .A1(_0205_),
    .A2(_0208_));
 sg13g2_inv_1 _1847_ (.Y(_0213_),
    .A(_0212_));
 sg13g2_o21ai_1 _1848_ (.B1(_0204_),
    .Y(_0214_),
    .A1(_0199_),
    .A2(_0213_));
 sg13g2_nor2b_1 _1849_ (.A(_0210_),
    .B_N(_0214_),
    .Y(_0215_));
 sg13g2_or2_1 _1850_ (.X(_0216_),
    .B(_0209_),
    .A(_0196_));
 sg13g2_nand2b_1 _1851_ (.Y(_0217_),
    .B(_0213_),
    .A_N(_0196_));
 sg13g2_and4_1 _1852_ (.A(_0200_),
    .B(_0215_),
    .C(_0216_),
    .D(_0217_),
    .X(_0218_));
 sg13g2_nand2_1 _1853_ (.Y(_0219_),
    .A(_0203_),
    .B(_0218_));
 sg13g2_nor3_2 _1854_ (.A(_0924_),
    .B(_0925_),
    .C(_0926_),
    .Y(_0220_));
 sg13g2_and2_1 _1855_ (.A(_0219_),
    .B(_0220_),
    .X(_0221_));
 sg13g2_a21oi_2 _1856_ (.B1(_0928_),
    .Y(uo_out[4]),
    .A2(_0221_),
    .A1(_0200_));
 sg13g2_nand3_1 _1857_ (.B(_0680_),
    .C(_0925_),
    .A(_0626_),
    .Y(_0222_));
 sg13g2_nand2_1 _1858_ (.Y(_0223_),
    .A(_0624_),
    .B(_0222_));
 sg13g2_a21oi_2 _1859_ (.B1(_0223_),
    .Y(uo_out[0]),
    .A2(_0221_),
    .A1(_0211_));
 sg13g2_o21ai_1 _1860_ (.B1(_0624_),
    .Y(_0224_),
    .A1(_0926_),
    .A2(_0220_));
 sg13g2_nor2_1 _1861_ (.A(\background_color[0] ),
    .B(_0390_),
    .Y(_0225_));
 sg13g2_a22oi_1 _1862_ (.Y(_0226_),
    .B1(_0225_),
    .B2(\background_color[1] ),
    .A2(_0201_),
    .A1(\background_color[2] ));
 sg13g2_nand2b_1 _1863_ (.Y(_0227_),
    .B(_0218_),
    .A_N(_0226_));
 sg13g2_nand3_1 _1864_ (.B(_0220_),
    .C(_0227_),
    .A(_0216_),
    .Y(_0228_));
 sg13g2_nor2b_2 _1865_ (.A(_0224_),
    .B_N(_0228_),
    .Y(uo_out[5]));
 sg13g2_nor2b_1 _1866_ (.A(_0210_),
    .B_N(_0227_),
    .Y(_0229_));
 sg13g2_a21oi_2 _1867_ (.B1(_0224_),
    .Y(uo_out[1]),
    .A2(_0229_),
    .A1(_0220_));
 sg13g2_nand2b_1 _1868_ (.Y(_0230_),
    .B(\background_color[1] ),
    .A_N(_0064_));
 sg13g2_o21ai_1 _1869_ (.B1(_0230_),
    .Y(_0231_),
    .A1(\background_color[1] ),
    .A2(_0063_));
 sg13g2_nand2_1 _1870_ (.Y(_0232_),
    .A(_0218_),
    .B(_0231_));
 sg13g2_nand3_1 _1871_ (.B(_0220_),
    .C(_0232_),
    .A(_0217_),
    .Y(_0233_));
 sg13g2_nor2b_2 _1872_ (.A(_0928_),
    .B_N(_0233_),
    .Y(uo_out[6]));
 sg13g2_a22oi_1 _1873_ (.Y(_0234_),
    .B1(_0218_),
    .B2(_0231_),
    .A2(_0213_),
    .A1(_0204_));
 sg13g2_a21oi_2 _1874_ (.B1(_0223_),
    .Y(uo_out[2]),
    .A2(_0234_),
    .A1(_0220_));
 sg13g2_nor2_1 _1875_ (.A(net301),
    .B(net302),
    .Y(_0235_));
 sg13g2_nand2b_1 _1876_ (.Y(_0236_),
    .B(_0072_),
    .A_N(net301));
 sg13g2_a21oi_1 _1877_ (.A1(net302),
    .A2(_0236_),
    .Y(_0056_),
    .B1(_0235_));
 sg13g2_a21oi_1 _1878_ (.A1(net301),
    .A2(net302),
    .Y(_0237_),
    .B1(net299));
 sg13g2_nand3_1 _1879_ (.B(net302),
    .C(_0236_),
    .A(net299),
    .Y(_0238_));
 sg13g2_nor2b_1 _1880_ (.A(_0237_),
    .B_N(_0238_),
    .Y(_0057_));
 sg13g2_nor2_1 _1881_ (.A(\audio_mod.audio_gen.chan0.ch_counter[0] ),
    .B(net279),
    .Y(_0000_));
 sg13g2_xnor2_1 _1882_ (.Y(_0239_),
    .A(\audio_mod.audio_gen.chan0.ch_counter[0] ),
    .B(\audio_mod.audio_gen.chan0.ch_counter[1] ));
 sg13g2_nor2_1 _1883_ (.A(net279),
    .B(_0239_),
    .Y(_0003_));
 sg13g2_and3_1 _1884_ (.X(_0240_),
    .A(\audio_mod.audio_gen.chan0.ch_counter[0] ),
    .B(\audio_mod.audio_gen.chan0.ch_counter[1] ),
    .C(\audio_mod.audio_gen.chan0.ch_counter[2] ));
 sg13g2_a21oi_1 _1885_ (.A1(\audio_mod.audio_gen.chan0.ch_counter[0] ),
    .A2(\audio_mod.audio_gen.chan0.ch_counter[1] ),
    .Y(_0241_),
    .B1(\audio_mod.audio_gen.chan0.ch_counter[2] ));
 sg13g2_nor3_1 _1886_ (.A(net279),
    .B(_0240_),
    .C(_0241_),
    .Y(_0004_));
 sg13g2_nor2_1 _1887_ (.A(\audio_mod.audio_gen.chan0.ch_counter[3] ),
    .B(_0240_),
    .Y(_0242_));
 sg13g2_and2_1 _1888_ (.A(\audio_mod.audio_gen.chan0.ch_counter[3] ),
    .B(_0240_),
    .X(_0243_));
 sg13g2_nor3_1 _1889_ (.A(net279),
    .B(_0242_),
    .C(_0243_),
    .Y(_0005_));
 sg13g2_and2_1 _1890_ (.A(\audio_mod.audio_gen.chan0.ch_counter[4] ),
    .B(_0243_),
    .X(_0244_));
 sg13g2_nor2_1 _1891_ (.A(\audio_mod.audio_gen.chan0.ch_counter[4] ),
    .B(_0243_),
    .Y(_0245_));
 sg13g2_nor3_1 _1892_ (.A(net279),
    .B(_0244_),
    .C(_0245_),
    .Y(_0006_));
 sg13g2_xnor2_1 _1893_ (.Y(_0246_),
    .A(\audio_mod.audio_gen.chan0.ch_counter[5] ),
    .B(_0244_));
 sg13g2_nor2_1 _1894_ (.A(net279),
    .B(_0246_),
    .Y(_0007_));
 sg13g2_nand3_1 _1895_ (.B(\audio_mod.audio_gen.chan0.ch_counter[6] ),
    .C(_0244_),
    .A(\audio_mod.audio_gen.chan0.ch_counter[5] ),
    .Y(_0247_));
 sg13g2_a21o_1 _1896_ (.A2(_0244_),
    .A1(\audio_mod.audio_gen.chan0.ch_counter[5] ),
    .B1(\audio_mod.audio_gen.chan0.ch_counter[6] ),
    .X(_0248_));
 sg13g2_nand2_1 _1897_ (.Y(_0249_),
    .A(_0247_),
    .B(_0248_));
 sg13g2_nor2_1 _1898_ (.A(net279),
    .B(_0249_),
    .Y(_0008_));
 sg13g2_nor2_1 _1899_ (.A(_0377_),
    .B(_0247_),
    .Y(_0250_));
 sg13g2_and2_1 _1900_ (.A(_0377_),
    .B(_0247_),
    .X(_0251_));
 sg13g2_nor3_1 _1901_ (.A(net280),
    .B(_0250_),
    .C(_0251_),
    .Y(_0009_));
 sg13g2_nor2_1 _1902_ (.A(\audio_mod.audio_gen.chan0.ch_counter[8] ),
    .B(_0250_),
    .Y(_0252_));
 sg13g2_and2_1 _1903_ (.A(\audio_mod.audio_gen.chan0.ch_counter[8] ),
    .B(_0250_),
    .X(_0253_));
 sg13g2_nor3_1 _1904_ (.A(net280),
    .B(_0252_),
    .C(_0253_),
    .Y(_0010_));
 sg13g2_xnor2_1 _1905_ (.Y(_0254_),
    .A(\audio_mod.audio_gen.chan0.ch_counter[9] ),
    .B(_0253_));
 sg13g2_nor2_1 _1906_ (.A(net280),
    .B(_0254_),
    .Y(_0011_));
 sg13g2_a21oi_1 _1907_ (.A1(\audio_mod.audio_gen.chan0.ch_counter[9] ),
    .A2(_0253_),
    .Y(_0255_),
    .B1(\audio_mod.audio_gen.chan0.ch_counter[10] ));
 sg13g2_nand3_1 _1908_ (.B(\audio_mod.audio_gen.chan0.ch_counter[10] ),
    .C(_0253_),
    .A(\audio_mod.audio_gen.chan0.ch_counter[9] ),
    .Y(_0256_));
 sg13g2_nand2b_1 _1909_ (.Y(_0257_),
    .B(_0256_),
    .A_N(_0255_));
 sg13g2_nor2_1 _1910_ (.A(net279),
    .B(_0257_),
    .Y(_0001_));
 sg13g2_xor2_1 _1911_ (.B(_0256_),
    .A(\audio_mod.audio_gen.chan0.ch_counter[11] ),
    .X(_0258_));
 sg13g2_nor2_1 _1912_ (.A(net280),
    .B(_0258_),
    .Y(_0002_));
 sg13g2_nor2_1 _1913_ (.A(\audio_mod.audio_gen.chan1.ch_counter[0] ),
    .B(net281),
    .Y(_0013_));
 sg13g2_and3_1 _1914_ (.X(_0259_),
    .A(\audio_mod.audio_gen.chan1.ch_counter[0] ),
    .B(\audio_mod.audio_gen.chan1.ch_counter[1] ),
    .C(\audio_mod.audio_gen.chan1.ch_counter[2] ));
 sg13g2_a21oi_1 _1915_ (.A1(\audio_mod.audio_gen.chan1.ch_counter[0] ),
    .A2(\audio_mod.audio_gen.chan1.ch_counter[1] ),
    .Y(_0260_),
    .B1(\audio_mod.audio_gen.chan1.ch_counter[2] ));
 sg13g2_nor3_1 _1916_ (.A(net281),
    .B(_0259_),
    .C(_0260_),
    .Y(_0017_));
 sg13g2_nor2_1 _1917_ (.A(\audio_mod.audio_gen.chan1.ch_counter[3] ),
    .B(_0259_),
    .Y(_0261_));
 sg13g2_and2_1 _1918_ (.A(\audio_mod.audio_gen.chan1.ch_counter[3] ),
    .B(_0259_),
    .X(_0262_));
 sg13g2_nor3_1 _1919_ (.A(net281),
    .B(_0261_),
    .C(_0262_),
    .Y(_0018_));
 sg13g2_and2_1 _1920_ (.A(\audio_mod.audio_gen.chan1.ch_counter[4] ),
    .B(_0262_),
    .X(_0263_));
 sg13g2_nor2_1 _1921_ (.A(\audio_mod.audio_gen.chan1.ch_counter[4] ),
    .B(_0262_),
    .Y(_0264_));
 sg13g2_nor3_1 _1922_ (.A(net281),
    .B(_0263_),
    .C(_0264_),
    .Y(_0019_));
 sg13g2_xnor2_1 _1923_ (.Y(_0265_),
    .A(\audio_mod.audio_gen.chan1.ch_counter[5] ),
    .B(_0263_));
 sg13g2_nor2_1 _1924_ (.A(net281),
    .B(_0265_),
    .Y(_0020_));
 sg13g2_nand3_1 _1925_ (.B(\audio_mod.audio_gen.chan1.ch_counter[6] ),
    .C(_0263_),
    .A(\audio_mod.audio_gen.chan1.ch_counter[5] ),
    .Y(_0266_));
 sg13g2_a21o_1 _1926_ (.A2(_0263_),
    .A1(\audio_mod.audio_gen.chan1.ch_counter[5] ),
    .B1(\audio_mod.audio_gen.chan1.ch_counter[6] ),
    .X(_0267_));
 sg13g2_nand2_1 _1927_ (.Y(_0268_),
    .A(_0266_),
    .B(_0267_));
 sg13g2_nor2_1 _1928_ (.A(net281),
    .B(_0268_),
    .Y(_0021_));
 sg13g2_nor2_1 _1929_ (.A(_0378_),
    .B(_0266_),
    .Y(_0269_));
 sg13g2_and2_1 _1930_ (.A(_0378_),
    .B(_0266_),
    .X(_0270_));
 sg13g2_nor3_1 _1931_ (.A(net281),
    .B(_0269_),
    .C(_0270_),
    .Y(_0022_));
 sg13g2_nor2_1 _1932_ (.A(\audio_mod.audio_gen.chan1.ch_counter[8] ),
    .B(_0269_),
    .Y(_0271_));
 sg13g2_and2_1 _1933_ (.A(\audio_mod.audio_gen.chan1.ch_counter[8] ),
    .B(_0269_),
    .X(_0272_));
 sg13g2_nor3_1 _1934_ (.A(_0513_),
    .B(_0271_),
    .C(_0272_),
    .Y(_0023_));
 sg13g2_xnor2_1 _1935_ (.Y(_0273_),
    .A(\audio_mod.audio_gen.chan1.ch_counter[9] ),
    .B(_0272_));
 sg13g2_nor2_1 _1936_ (.A(_0513_),
    .B(_0273_),
    .Y(_0024_));
 sg13g2_a21oi_1 _1937_ (.A1(\audio_mod.audio_gen.chan1.ch_counter[9] ),
    .A2(_0272_),
    .Y(_0274_),
    .B1(\audio_mod.audio_gen.chan1.ch_counter[10] ));
 sg13g2_nand3_1 _1938_ (.B(\audio_mod.audio_gen.chan1.ch_counter[10] ),
    .C(_0272_),
    .A(\audio_mod.audio_gen.chan1.ch_counter[9] ),
    .Y(_0275_));
 sg13g2_nand2b_1 _1939_ (.Y(_0276_),
    .B(_0275_),
    .A_N(_0274_));
 sg13g2_nor2_1 _1940_ (.A(net281),
    .B(_0276_),
    .Y(_0014_));
 sg13g2_xnor2_1 _1941_ (.Y(_0015_),
    .A(\audio_mod.audio_gen.chan1.ch_counter[11] ),
    .B(_0275_));
 sg13g2_nor2_1 _1942_ (.A(\audio_mod.audio_gen.chan2.ch_counter[0] ),
    .B(net277),
    .Y(_0026_));
 sg13g2_xnor2_1 _1943_ (.Y(_0277_),
    .A(\audio_mod.audio_gen.chan2.ch_counter[0] ),
    .B(\audio_mod.audio_gen.chan2.ch_counter[1] ));
 sg13g2_nor2_1 _1944_ (.A(net277),
    .B(_0277_),
    .Y(_0029_));
 sg13g2_and3_1 _1945_ (.X(_0278_),
    .A(\audio_mod.audio_gen.chan2.ch_counter[0] ),
    .B(\audio_mod.audio_gen.chan2.ch_counter[1] ),
    .C(\audio_mod.audio_gen.chan2.ch_counter[2] ));
 sg13g2_a21oi_1 _1946_ (.A1(\audio_mod.audio_gen.chan2.ch_counter[0] ),
    .A2(\audio_mod.audio_gen.chan2.ch_counter[1] ),
    .Y(_0279_),
    .B1(\audio_mod.audio_gen.chan2.ch_counter[2] ));
 sg13g2_nor3_1 _1947_ (.A(net277),
    .B(_0278_),
    .C(_0279_),
    .Y(_0030_));
 sg13g2_nor2_1 _1948_ (.A(\audio_mod.audio_gen.chan2.ch_counter[3] ),
    .B(_0278_),
    .Y(_0280_));
 sg13g2_and2_1 _1949_ (.A(\audio_mod.audio_gen.chan2.ch_counter[3] ),
    .B(_0278_),
    .X(_0281_));
 sg13g2_nor3_1 _1950_ (.A(net278),
    .B(_0280_),
    .C(_0281_),
    .Y(_0031_));
 sg13g2_and2_1 _1951_ (.A(\audio_mod.audio_gen.chan2.ch_counter[4] ),
    .B(_0281_),
    .X(_0282_));
 sg13g2_nor2_1 _1952_ (.A(\audio_mod.audio_gen.chan2.ch_counter[4] ),
    .B(_0281_),
    .Y(_0283_));
 sg13g2_nor3_1 _1953_ (.A(net277),
    .B(_0282_),
    .C(_0283_),
    .Y(_0032_));
 sg13g2_xnor2_1 _1954_ (.Y(_0284_),
    .A(\audio_mod.audio_gen.chan2.ch_counter[5] ),
    .B(_0282_));
 sg13g2_nor2_1 _1955_ (.A(net277),
    .B(_0284_),
    .Y(_0033_));
 sg13g2_nand3_1 _1956_ (.B(\audio_mod.audio_gen.chan2.ch_counter[6] ),
    .C(_0282_),
    .A(\audio_mod.audio_gen.chan2.ch_counter[5] ),
    .Y(_0285_));
 sg13g2_a21o_1 _1957_ (.A2(_0282_),
    .A1(\audio_mod.audio_gen.chan2.ch_counter[5] ),
    .B1(\audio_mod.audio_gen.chan2.ch_counter[6] ),
    .X(_0286_));
 sg13g2_nand2_1 _1958_ (.Y(_0287_),
    .A(_0285_),
    .B(_0286_));
 sg13g2_nor2_1 _1959_ (.A(net277),
    .B(_0287_),
    .Y(_0034_));
 sg13g2_and2_1 _1960_ (.A(_0379_),
    .B(_0285_),
    .X(_0288_));
 sg13g2_nor2_1 _1961_ (.A(_0379_),
    .B(_0285_),
    .Y(_0289_));
 sg13g2_nor3_1 _1962_ (.A(net278),
    .B(_0288_),
    .C(_0289_),
    .Y(_0035_));
 sg13g2_nor2_1 _1963_ (.A(\audio_mod.audio_gen.chan2.ch_counter[8] ),
    .B(_0289_),
    .Y(_0290_));
 sg13g2_and2_1 _1964_ (.A(\audio_mod.audio_gen.chan2.ch_counter[8] ),
    .B(_0289_),
    .X(_0291_));
 sg13g2_nor3_1 _1965_ (.A(net277),
    .B(_0290_),
    .C(_0291_),
    .Y(_0036_));
 sg13g2_xnor2_1 _1966_ (.Y(_0292_),
    .A(\audio_mod.audio_gen.chan2.ch_counter[9] ),
    .B(_0291_));
 sg13g2_nor2_1 _1967_ (.A(net278),
    .B(_0292_),
    .Y(_0037_));
 sg13g2_a21oi_1 _1968_ (.A1(\audio_mod.audio_gen.chan2.ch_counter[9] ),
    .A2(_0291_),
    .Y(_0293_),
    .B1(\audio_mod.audio_gen.chan2.ch_counter[10] ));
 sg13g2_nand2b_1 _1969_ (.Y(_0294_),
    .B(_0291_),
    .A_N(_0458_));
 sg13g2_nand2b_1 _1970_ (.Y(_0295_),
    .B(_0294_),
    .A_N(_0293_));
 sg13g2_nor2_1 _1971_ (.A(net278),
    .B(_0295_),
    .Y(_0027_));
 sg13g2_xnor2_1 _1972_ (.Y(_0296_),
    .A(_0074_),
    .B(_0294_));
 sg13g2_nor2_1 _1973_ (.A(net277),
    .B(_0296_),
    .Y(_0028_));
 sg13g2_nor2_1 _1974_ (.A(\audio_mod.audio_gen.chan3.ch_counter[0] ),
    .B(_0423_),
    .Y(_0039_));
 sg13g2_xor2_1 _1975_ (.B(\audio_mod.audio_gen.chan3.ch_counter[1] ),
    .A(\audio_mod.audio_gen.chan3.ch_counter[0] ),
    .X(_0042_));
 sg13g2_and3_1 _1976_ (.X(_0297_),
    .A(\audio_mod.audio_gen.chan3.ch_counter[0] ),
    .B(\audio_mod.audio_gen.chan3.ch_counter[1] ),
    .C(\audio_mod.audio_gen.chan3.ch_counter[2] ));
 sg13g2_a21oi_1 _1977_ (.A1(\audio_mod.audio_gen.chan3.ch_counter[0] ),
    .A2(\audio_mod.audio_gen.chan3.ch_counter[1] ),
    .Y(_0298_),
    .B1(\audio_mod.audio_gen.chan3.ch_counter[2] ));
 sg13g2_nor3_1 _1978_ (.A(_0423_),
    .B(_0297_),
    .C(_0298_),
    .Y(_0043_));
 sg13g2_nor2_1 _1979_ (.A(\audio_mod.audio_gen.chan3.ch_counter[3] ),
    .B(_0297_),
    .Y(_0299_));
 sg13g2_and2_1 _1980_ (.A(\audio_mod.audio_gen.chan3.ch_counter[3] ),
    .B(_0297_),
    .X(_0300_));
 sg13g2_nor3_1 _1981_ (.A(_0423_),
    .B(_0299_),
    .C(_0300_),
    .Y(_0044_));
 sg13g2_and2_1 _1982_ (.A(\audio_mod.audio_gen.chan3.ch_counter[4] ),
    .B(_0300_),
    .X(_0301_));
 sg13g2_nor2_1 _1983_ (.A(\audio_mod.audio_gen.chan3.ch_counter[4] ),
    .B(_0300_),
    .Y(_0302_));
 sg13g2_nor3_1 _1984_ (.A(_0423_),
    .B(_0301_),
    .C(_0302_),
    .Y(_0045_));
 sg13g2_nor2_1 _1985_ (.A(\audio_mod.audio_gen.chan3.ch_counter[5] ),
    .B(_0301_),
    .Y(_0303_));
 sg13g2_and2_1 _1986_ (.A(\audio_mod.audio_gen.chan3.ch_counter[5] ),
    .B(_0301_),
    .X(_0304_));
 sg13g2_nor3_1 _1987_ (.A(_0423_),
    .B(_0303_),
    .C(_0304_),
    .Y(_0046_));
 sg13g2_and2_1 _1988_ (.A(\audio_mod.audio_gen.chan3.ch_counter[6] ),
    .B(_0304_),
    .X(_0305_));
 sg13g2_nor2_1 _1989_ (.A(\audio_mod.audio_gen.chan3.ch_counter[6] ),
    .B(_0304_),
    .Y(_0306_));
 sg13g2_nor3_1 _1990_ (.A(_0423_),
    .B(_0305_),
    .C(_0306_),
    .Y(_0047_));
 sg13g2_xor2_1 _1991_ (.B(_0305_),
    .A(\audio_mod.audio_gen.chan3.ch_counter[7] ),
    .X(_0048_));
 sg13g2_a21oi_1 _1992_ (.A1(\audio_mod.audio_gen.chan3.ch_counter[7] ),
    .A2(_0305_),
    .Y(_0307_),
    .B1(\audio_mod.audio_gen.chan3.ch_counter[8] ));
 sg13g2_and3_1 _1993_ (.X(_0308_),
    .A(\audio_mod.audio_gen.chan3.ch_counter[7] ),
    .B(\audio_mod.audio_gen.chan3.ch_counter[8] ),
    .C(_0305_));
 sg13g2_nor3_1 _1994_ (.A(_0423_),
    .B(_0307_),
    .C(_0308_),
    .Y(_0049_));
 sg13g2_xor2_1 _1995_ (.B(_0308_),
    .A(\audio_mod.audio_gen.chan3.ch_counter[9] ),
    .X(_0050_));
 sg13g2_nand3_1 _1996_ (.B(\audio_mod.audio_gen.chan3.ch_counter[10] ),
    .C(_0308_),
    .A(\audio_mod.audio_gen.chan3.ch_counter[9] ),
    .Y(_0309_));
 sg13g2_a21o_1 _1997_ (.A2(_0308_),
    .A1(\audio_mod.audio_gen.chan3.ch_counter[9] ),
    .B1(\audio_mod.audio_gen.chan3.ch_counter[10] ),
    .X(_0310_));
 sg13g2_and2_1 _1998_ (.A(_0309_),
    .B(_0310_),
    .X(_0040_));
 sg13g2_xnor2_1 _1999_ (.Y(_0041_),
    .A(\audio_mod.audio_gen.chan3.ch_counter[11] ),
    .B(_0309_));
 sg13g2_xor2_1 _2000_ (.B(\audio_mod.seq.seq_clock[0] ),
    .A(\audio_mod.seq.seq_clock[1] ),
    .X(_0052_));
 sg13g2_nand3_1 _2001_ (.B(\audio_mod.seq.seq_clock[1] ),
    .C(\audio_mod.seq.seq_clock[0] ),
    .A(\audio_mod.seq.seq_clock[2] ),
    .Y(_0311_));
 sg13g2_a21o_1 _2002_ (.A2(_0474_),
    .A1(\audio_mod.seq.seq_clock[0] ),
    .B1(\audio_mod.seq.seq_clock[2] ),
    .X(_0312_));
 sg13g2_and2_1 _2003_ (.A(_0311_),
    .B(_0312_),
    .X(_0053_));
 sg13g2_xnor2_1 _2004_ (.Y(_0054_),
    .A(\audio_mod.seq.seq_clock[3] ),
    .B(_0311_));
 sg13g2_xnor2_1 _2005_ (.Y(_0060_),
    .A(net51),
    .B(net48));
 sg13g2_nor2_1 _2006_ (.A(net297),
    .B(_0988_),
    .Y(_0085_));
 sg13g2_xor2_1 _2007_ (.B(net52),
    .A(\audio_mod.audio_gen.pwm_clock[1] ),
    .X(_0091_));
 sg13g2_nand3_1 _2008_ (.B(net52),
    .C(net344),
    .A(net74),
    .Y(_0313_));
 sg13g2_a21o_1 _2009_ (.A2(net52),
    .A1(net74),
    .B1(net344),
    .X(_0314_));
 sg13g2_and2_1 _2010_ (.A(_0313_),
    .B(_0314_),
    .X(_0092_));
 sg13g2_nand4_1 _2011_ (.B(net52),
    .C(net56),
    .A(net74),
    .Y(_0315_),
    .D(net344));
 sg13g2_xnor2_1 _2012_ (.Y(_0093_),
    .A(net56),
    .B(_0313_));
 sg13g2_nor2_1 _2013_ (.A(_0376_),
    .B(_0315_),
    .Y(_0316_));
 sg13g2_xnor2_1 _2014_ (.Y(_0094_),
    .A(net54),
    .B(_0315_));
 sg13g2_xor2_1 _2015_ (.B(_0316_),
    .A(net336),
    .X(_0095_));
 sg13g2_nand2b_1 _2016_ (.Y(_0317_),
    .B(net297),
    .A_N(_0062_));
 sg13g2_xnor2_1 _2017_ (.Y(_0087_),
    .A(net303),
    .B(_0317_));
 sg13g2_and2_1 _2018_ (.A(net304),
    .B(net303),
    .X(_0318_));
 sg13g2_nand2_1 _2019_ (.Y(_0319_),
    .A(net297),
    .B(_0318_));
 sg13g2_xnor2_1 _2020_ (.Y(_0088_),
    .A(\counter[4] ),
    .B(_0319_));
 sg13g2_nor2_1 _2021_ (.A(_0083_),
    .B(_0319_),
    .Y(_0320_));
 sg13g2_xor2_1 _2022_ (.B(_0320_),
    .A(\counter[5] ),
    .X(_0089_));
 sg13g2_nand4_1 _2023_ (.B(\counter[5] ),
    .C(net297),
    .A(\counter[4] ),
    .Y(_0321_),
    .D(_0318_));
 sg13g2_xnor2_1 _2024_ (.Y(_0090_),
    .A(\counter[6] ),
    .B(_0321_));
 sg13g2_xor2_1 _2025_ (.B(_0427_),
    .A(net292),
    .X(_0097_));
 sg13g2_a21oi_1 _2026_ (.A1(net291),
    .A2(_0427_),
    .Y(_0322_),
    .B1(net289));
 sg13g2_a21oi_1 _2027_ (.A1(net294),
    .A2(_0436_),
    .Y(_0098_),
    .B1(_0322_));
 sg13g2_nor3_1 _2028_ (.A(net300),
    .B(net299),
    .C(net302),
    .Y(_0104_));
 sg13g2_or4_1 _2029_ (.A(\audio_mod.audio_gen.pwm_clock[1] ),
    .B(\audio_mod.audio_gen.pwm_clock[0] ),
    .C(\audio_mod.audio_gen.pwm_clock[3] ),
    .D(\audio_mod.audio_gen.pwm_clock[4] ),
    .X(_0323_));
 sg13g2_nor3_1 _2030_ (.A(net338),
    .B(net329),
    .C(net307),
    .Y(_0108_));
 sg13g2_and2_1 _2031_ (.A(net81),
    .B(net320),
    .X(_0324_));
 sg13g2_and2_1 _2032_ (.A(net81),
    .B(_0769_),
    .X(_0325_));
 sg13g2_nand2_2 _2033_ (.Y(_0326_),
    .A(net320),
    .B(_0752_));
 sg13g2_nand3_1 _2034_ (.B(_0385_),
    .C(_0386_),
    .A(_0383_),
    .Y(_0327_));
 sg13g2_nor4_2 _2035_ (.A(_0384_),
    .B(_0612_),
    .C(_0326_),
    .Y(_0328_),
    .D(_0327_));
 sg13g2_nor2b_1 _2036_ (.A(_0328_),
    .B_N(net365),
    .Y(_0329_));
 sg13g2_nand2b_2 _2037_ (.Y(_0330_),
    .B(net365),
    .A_N(_0328_));
 sg13g2_nor3_1 _2038_ (.A(_0381_),
    .B(net321),
    .C(\hvsync_gen.vpos[6] ),
    .Y(_0331_));
 sg13g2_nand4_1 _2039_ (.B(_0745_),
    .C(_0758_),
    .A(_0646_),
    .Y(_0332_),
    .D(_0331_));
 sg13g2_nand2_1 _2040_ (.Y(_0333_),
    .A(net365),
    .B(_0332_));
 sg13g2_inv_1 _2041_ (.Y(_0334_),
    .A(_0333_));
 sg13g2_nand2_2 _2042_ (.Y(_0335_),
    .A(_0328_),
    .B(_0334_));
 sg13g2_inv_1 _2043_ (.Y(_0336_),
    .A(_0335_));
 sg13g2_a22oi_1 _2044_ (.Y(_0337_),
    .B1(_0336_),
    .B2(net45),
    .A2(net287),
    .A1(\hvsync_gen.vpos[0] ));
 sg13g2_inv_1 _2045_ (.Y(_0169_),
    .A(net46));
 sg13g2_nor3_1 _2046_ (.A(_0646_),
    .B(_0759_),
    .C(_0335_),
    .Y(_0338_));
 sg13g2_a21o_1 _2047_ (.A2(net286),
    .A1(net65),
    .B1(_0338_),
    .X(_0170_));
 sg13g2_nor2_2 _2048_ (.A(net286),
    .B(_0334_),
    .Y(_0339_));
 sg13g2_nor2_1 _2049_ (.A(_0760_),
    .B(net286),
    .Y(_0340_));
 sg13g2_xnor2_1 _2050_ (.Y(_0341_),
    .A(net75),
    .B(_0340_));
 sg13g2_nor2_1 _2051_ (.A(_0339_),
    .B(_0341_),
    .Y(_0171_));
 sg13g2_nor3_1 _2052_ (.A(net63),
    .B(_0760_),
    .C(net286),
    .Y(_0342_));
 sg13g2_xnor2_1 _2053_ (.Y(_0343_),
    .A(net327),
    .B(_0342_));
 sg13g2_nor2_1 _2054_ (.A(_0339_),
    .B(net64),
    .Y(_0172_));
 sg13g2_a21oi_1 _2055_ (.A1(_0745_),
    .A2(_0340_),
    .Y(_0344_),
    .B1(net326));
 sg13g2_nor3_2 _2056_ (.A(_0747_),
    .B(_0760_),
    .C(net286),
    .Y(_0345_));
 sg13g2_nor3_1 _2057_ (.A(_0339_),
    .B(_0344_),
    .C(_0345_),
    .Y(_0173_));
 sg13g2_nand2_1 _2058_ (.Y(_0346_),
    .A(net324),
    .B(net286));
 sg13g2_nor3_1 _2059_ (.A(net71),
    .B(_0746_),
    .C(_0760_),
    .Y(_0347_));
 sg13g2_xnor2_1 _2060_ (.Y(_0348_),
    .A(net324),
    .B(_0347_));
 sg13g2_o21ai_1 _2061_ (.B1(_0346_),
    .Y(_0174_),
    .A1(_0335_),
    .A2(_0348_));
 sg13g2_a21oi_1 _2062_ (.A1(net324),
    .A2(_0345_),
    .Y(_0349_),
    .B1(net67));
 sg13g2_nor2b_1 _2063_ (.A(_0610_),
    .B_N(_0345_),
    .Y(_0350_));
 sg13g2_nor3_1 _2064_ (.A(_0339_),
    .B(_0349_),
    .C(_0350_),
    .Y(_0175_));
 sg13g2_nand2_1 _2065_ (.Y(_0351_),
    .A(net322),
    .B(net286));
 sg13g2_or4_1 _2066_ (.A(_0382_),
    .B(_0067_),
    .C(_0747_),
    .D(_0760_),
    .X(_0352_));
 sg13g2_xor2_1 _2067_ (.B(_0352_),
    .A(net322),
    .X(_0353_));
 sg13g2_o21ai_1 _2068_ (.B1(_0351_),
    .Y(_0176_),
    .A1(_0335_),
    .A2(_0353_));
 sg13g2_nand2_1 _2069_ (.Y(_0354_),
    .A(net322),
    .B(_0350_));
 sg13g2_xor2_1 _2070_ (.B(_0354_),
    .A(net321),
    .X(_0355_));
 sg13g2_nor2_1 _2071_ (.A(_0339_),
    .B(_0355_),
    .Y(_0177_));
 sg13g2_nand2_1 _2072_ (.Y(_0356_),
    .A(net58),
    .B(net287));
 sg13g2_nor4_1 _2073_ (.A(_0069_),
    .B(_0611_),
    .C(_0747_),
    .D(_0760_),
    .Y(_0357_));
 sg13g2_xnor2_1 _2074_ (.Y(_0358_),
    .A(net58),
    .B(_0357_));
 sg13g2_o21ai_1 _2075_ (.B1(_0356_),
    .Y(_0178_),
    .A1(_0335_),
    .A2(_0358_));
 sg13g2_and2_1 _2076_ (.A(net43),
    .B(net286),
    .X(_0183_));
 sg13g2_nor3_1 _2077_ (.A(_0636_),
    .B(_0324_),
    .C(_0330_),
    .Y(_0184_));
 sg13g2_nor2_1 _2078_ (.A(net319),
    .B(_0324_),
    .Y(_0359_));
 sg13g2_nor3_1 _2079_ (.A(_0325_),
    .B(_0330_),
    .C(_0359_),
    .Y(_0185_));
 sg13g2_o21ai_1 _2080_ (.B1(net365),
    .Y(_0360_),
    .A1(net76),
    .A2(_0325_));
 sg13g2_nor2b_1 _2081_ (.A(_0360_),
    .B_N(_0326_),
    .Y(_0186_));
 sg13g2_o21ai_1 _2082_ (.B1(net365),
    .Y(_0361_),
    .A1(_0384_),
    .A2(_0326_));
 sg13g2_a21oi_1 _2083_ (.A1(_0384_),
    .A2(_0326_),
    .Y(_0187_),
    .B1(_0361_));
 sg13g2_nor2_1 _2084_ (.A(_0077_),
    .B(_0326_),
    .Y(_0362_));
 sg13g2_xnor2_1 _2085_ (.Y(_0363_),
    .A(net72),
    .B(_0362_));
 sg13g2_nor2_1 _2086_ (.A(_0330_),
    .B(net73),
    .Y(_0188_));
 sg13g2_nor2_1 _2087_ (.A(_0615_),
    .B(_0326_),
    .Y(_0364_));
 sg13g2_xnor2_1 _2088_ (.Y(_0365_),
    .A(net66),
    .B(_0364_));
 sg13g2_nor2_1 _2089_ (.A(_0330_),
    .B(_0365_),
    .Y(_0189_));
 sg13g2_nor3_1 _2090_ (.A(net69),
    .B(_0615_),
    .C(_0326_),
    .Y(_0366_));
 sg13g2_xnor2_1 _2091_ (.Y(_0367_),
    .A(net318),
    .B(_0366_));
 sg13g2_nor2_1 _2092_ (.A(_0330_),
    .B(net70),
    .Y(_0190_));
 sg13g2_or2_1 _2093_ (.X(_0368_),
    .B(_0326_),
    .A(_0616_));
 sg13g2_xor2_1 _2094_ (.B(_0368_),
    .A(net68),
    .X(_0369_));
 sg13g2_nor2_1 _2095_ (.A(_0330_),
    .B(_0369_),
    .Y(_0191_));
 sg13g2_nor2_1 _2096_ (.A(_0081_),
    .B(_0368_),
    .Y(_0370_));
 sg13g2_o21ai_1 _2097_ (.B1(net287),
    .Y(_0371_),
    .A1(net316),
    .A2(_0370_));
 sg13g2_a21oi_1 _2098_ (.A1(net316),
    .A2(_0370_),
    .Y(_0192_),
    .B1(_0371_));
 sg13g2_nor3_1 _2099_ (.A(net301),
    .B(net299),
    .C(net302),
    .Y(_0105_));
 sg13g2_nor3_1 _2100_ (.A(net300),
    .B(net299),
    .C(net302),
    .Y(_0106_));
 sg13g2_nor3_1 _2101_ (.A(net300),
    .B(net299),
    .C(\clock_gen.r_atick_clock[0] ),
    .Y(_0107_));
 sg13g2_nor3_1 _2102_ (.A(net338),
    .B(net329),
    .C(net307),
    .Y(_0109_));
 sg13g2_nor3_1 _2103_ (.A(net338),
    .B(net329),
    .C(net307),
    .Y(_0110_));
 sg13g2_nor3_1 _2104_ (.A(net338),
    .B(net329),
    .C(net307),
    .Y(_0111_));
 sg13g2_nor3_1 _2105_ (.A(net338),
    .B(net329),
    .C(net307),
    .Y(_0112_));
 sg13g2_nor3_1 _2106_ (.A(net338),
    .B(net329),
    .C(net307),
    .Y(_0113_));
 sg13g2_nor3_1 _2107_ (.A(net338),
    .B(net329),
    .C(net312),
    .Y(_0114_));
 sg13g2_nor3_1 _2108_ (.A(net340),
    .B(net331),
    .C(net309),
    .Y(_0115_));
 sg13g2_nor3_1 _2109_ (.A(net343),
    .B(net334),
    .C(net312),
    .Y(_0116_));
 sg13g2_nor3_1 _2110_ (.A(net343),
    .B(net334),
    .C(net309),
    .Y(_0117_));
 sg13g2_nor3_1 _2111_ (.A(net340),
    .B(net331),
    .C(net309),
    .Y(_0118_));
 sg13g2_nor3_1 _2112_ (.A(net340),
    .B(net331),
    .C(net313),
    .Y(_0119_));
 sg13g2_nor3_1 _2113_ (.A(net339),
    .B(net330),
    .C(net308),
    .Y(_0120_));
 sg13g2_nor3_1 _2114_ (.A(net341),
    .B(net332),
    .C(net310),
    .Y(_0121_));
 sg13g2_nor3_1 _2115_ (.A(net341),
    .B(net332),
    .C(net310),
    .Y(_0122_));
 sg13g2_nor3_1 _2116_ (.A(net339),
    .B(net330),
    .C(net308),
    .Y(_0123_));
 sg13g2_nor3_1 _2117_ (.A(net339),
    .B(net330),
    .C(net308),
    .Y(_0124_));
 sg13g2_nor3_1 _2118_ (.A(net339),
    .B(net330),
    .C(net307),
    .Y(_0125_));
 sg13g2_nor3_1 _2119_ (.A(net338),
    .B(net329),
    .C(net307),
    .Y(_0126_));
 sg13g2_nor3_1 _2120_ (.A(net339),
    .B(net330),
    .C(net308),
    .Y(_0127_));
 sg13g2_nor3_1 _2121_ (.A(net340),
    .B(net331),
    .C(net309),
    .Y(_0128_));
 sg13g2_nor3_1 _2122_ (.A(net340),
    .B(net331),
    .C(net309),
    .Y(_0129_));
 sg13g2_nor3_1 _2123_ (.A(net342),
    .B(net333),
    .C(net312),
    .Y(_0130_));
 sg13g2_nor3_1 _2124_ (.A(net341),
    .B(net332),
    .C(net310),
    .Y(_0131_));
 sg13g2_nor3_1 _2125_ (.A(net344),
    .B(net336),
    .C(net314),
    .Y(_0132_));
 sg13g2_nor3_1 _2126_ (.A(net342),
    .B(net333),
    .C(net310),
    .Y(_0133_));
 sg13g2_nor3_1 _2127_ (.A(net342),
    .B(net333),
    .C(net311),
    .Y(_0134_));
 sg13g2_nor3_1 _2128_ (.A(net341),
    .B(net332),
    .C(net310),
    .Y(_0135_));
 sg13g2_nor3_1 _2129_ (.A(net341),
    .B(net332),
    .C(net311),
    .Y(_0136_));
 sg13g2_nor3_1 _2130_ (.A(net341),
    .B(net332),
    .C(net310),
    .Y(_0137_));
 sg13g2_nor3_1 _2131_ (.A(net341),
    .B(net332),
    .C(net310),
    .Y(_0138_));
 sg13g2_nor3_1 _2132_ (.A(net341),
    .B(net333),
    .C(net310),
    .Y(_0139_));
 sg13g2_nor3_1 _2133_ (.A(net342),
    .B(net332),
    .C(net311),
    .Y(_0140_));
 sg13g2_nor3_1 _2134_ (.A(net342),
    .B(net333),
    .C(net311),
    .Y(_0141_));
 sg13g2_nor3_1 _2135_ (.A(net342),
    .B(net333),
    .C(net311),
    .Y(_0142_));
 sg13g2_nor3_1 _2136_ (.A(net342),
    .B(net333),
    .C(net311),
    .Y(_0143_));
 sg13g2_nor3_1 _2137_ (.A(net343),
    .B(net334),
    .C(net311),
    .Y(_0144_));
 sg13g2_nor3_1 _2138_ (.A(net340),
    .B(net331),
    .C(net309),
    .Y(_0145_));
 sg13g2_nor3_1 _2139_ (.A(net345),
    .B(net335),
    .C(net314),
    .Y(_0146_));
 sg13g2_nor3_1 _2140_ (.A(net345),
    .B(net335),
    .C(net313),
    .Y(_0147_));
 sg13g2_nor3_1 _2141_ (.A(net344),
    .B(net336),
    .C(net314),
    .Y(_0148_));
 sg13g2_nor3_1 _2142_ (.A(net344),
    .B(net336),
    .C(net314),
    .Y(_0149_));
 sg13g2_nor3_1 _2143_ (.A(net344),
    .B(net336),
    .C(net314),
    .Y(_0150_));
 sg13g2_nor3_1 _2144_ (.A(net344),
    .B(net336),
    .C(net314),
    .Y(_0151_));
 sg13g2_nor3_1 _2145_ (.A(net345),
    .B(net335),
    .C(net313),
    .Y(_0152_));
 sg13g2_nor3_1 _2146_ (.A(net345),
    .B(net335),
    .C(net313),
    .Y(_0153_));
 sg13g2_nor3_1 _2147_ (.A(net345),
    .B(net335),
    .C(net313),
    .Y(_0154_));
 sg13g2_nor3_1 _2148_ (.A(net345),
    .B(net335),
    .C(net313),
    .Y(_0155_));
 sg13g2_nor3_1 _2149_ (.A(net345),
    .B(net335),
    .C(net313),
    .Y(_0156_));
 sg13g2_nor3_1 _2150_ (.A(net345),
    .B(net335),
    .C(net313),
    .Y(_0157_));
 sg13g2_nor3_1 _2151_ (.A(net347),
    .B(net337),
    .C(net315),
    .Y(_0158_));
 sg13g2_nor3_1 _2152_ (.A(net346),
    .B(net336),
    .C(net314),
    .Y(_0159_));
 sg13g2_dfrbp_1 _2153_ (.CLK(\clock_gen.vsync ),
    .RESET_B(net364),
    .D(_1037_),
    .Q_N(_1037_),
    .Q(\counter[0] ));
 sg13g2_dfrbp_1 _2154_ (.CLK(\clock_gen.vsync ),
    .RESET_B(net364),
    .D(_0085_),
    .Q_N(_1100_),
    .Q(\counter[1] ));
 sg13g2_dfrbp_1 _2155_ (.CLK(net328),
    .RESET_B(net364),
    .D(_0086_),
    .Q_N(_0062_),
    .Q(\counter[2] ));
 sg13g2_dfrbp_1 _2156_ (.CLK(net328),
    .RESET_B(net364),
    .D(_0087_),
    .Q_N(_0082_),
    .Q(\counter[3] ));
 sg13g2_dfrbp_1 _2157_ (.CLK(net328),
    .RESET_B(net363),
    .D(_0088_),
    .Q_N(_0083_),
    .Q(\counter[4] ));
 sg13g2_dfrbp_1 _2158_ (.CLK(net328),
    .RESET_B(net363),
    .D(_0089_),
    .Q_N(_0084_),
    .Q(\counter[5] ));
 sg13g2_dfrbp_1 _2159_ (.CLK(net328),
    .RESET_B(net363),
    .D(_0090_),
    .Q_N(_0061_),
    .Q(\counter[6] ));
 sg13g2_dfrbp_1 _2160_ (.CLK(_1104_),
    .RESET_B(net359),
    .D(_0160_),
    .Q_N(_0101_),
    .Q(\stage[0] ));
 sg13g2_dfrbp_1 _2161_ (.CLK(_1104_),
    .RESET_B(net359),
    .D(_0161_),
    .Q_N(_1101_),
    .Q(\stage[1] ));
 sg13g2_dfrbp_1 _2162_ (.CLK(net328),
    .RESET_B(net361),
    .D(_0055_),
    .Q_N(_1102_),
    .Q(\clock_gen.r_atick_clock[0] ));
 sg13g2_dfrbp_1 _2163_ (.CLK(net328),
    .RESET_B(net361),
    .D(_0056_),
    .Q_N(_1103_),
    .Q(\atick_clock[0] ));
 sg13g2_dfrbp_1 _2164_ (.CLK(net328),
    .RESET_B(net361),
    .D(_0057_),
    .Q_N(_0072_),
    .Q(\atick_clock[1] ));
 sg13g2_dfrbp_1 _2165_ (.CLK(_0104_),
    .RESET_B(net361),
    .D(_1038_),
    .Q_N(_1038_),
    .Q(\audio_mod.pattern_clock[0] ));
 sg13g2_dfrbp_1 _2166_ (.CLK(_0105_),
    .RESET_B(net361),
    .D(_0096_),
    .Q_N(_1099_),
    .Q(\audio_mod.pattern_clock[1] ));
 sg13g2_dfrbp_1 _2167_ (.CLK(_0106_),
    .RESET_B(net363),
    .D(_0097_),
    .Q_N(_1098_),
    .Q(\audio_mod.pattern_clock[2] ));
 sg13g2_dfrbp_1 _2168_ (.CLK(_0107_),
    .RESET_B(net361),
    .D(_0098_),
    .Q_N(_1104_),
    .Q(\audio_mod.pattern_clock[3] ));
 sg13g2_dfrbp_1 _2169_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net356),
    .D(net35),
    .Q_N(_1036_),
    .Q(\audio_mod.audio_gen.pwm_clock[0] ));
 sg13g2_dfrbp_1 _2170_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net356),
    .D(net53),
    .Q_N(_1105_),
    .Q(\audio_mod.audio_gen.pwm_clock[1] ));
 sg13g2_dfrbp_1 _2171_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net356),
    .D(_0092_),
    .Q_N(_1106_),
    .Q(\audio_mod.audio_gen.pwm_clock[2] ));
 sg13g2_dfrbp_1 _2172_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net356),
    .D(net57),
    .Q_N(_1107_),
    .Q(\audio_mod.audio_gen.pwm_clock[3] ));
 sg13g2_dfrbp_1 _2173_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net356),
    .D(net55),
    .Q_N(_1108_),
    .Q(\audio_mod.audio_gen.pwm_clock[4] ));
 sg13g2_dfrbp_1 _2174_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net356),
    .D(_0095_),
    .Q_N(_1109_),
    .Q(\audio_mod.audio_gen.pwm_clock[5] ));
 sg13g2_dfrbp_1 _2175_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net359),
    .D(net44),
    .Q_N(_0073_),
    .Q(\audio_mod.audio_gen.chan3.rng ));
 sg13g2_dfrbp_1 _2176_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net357),
    .D(net48),
    .Q_N(_1110_),
    .Q(\lfsr[1] ));
 sg13g2_dfrbp_1 _2177_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net360),
    .D(net47),
    .Q_N(_1111_),
    .Q(\lfsr[2] ));
 sg13g2_dfrbp_1 _2178_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net360),
    .D(net41),
    .Q_N(_1112_),
    .Q(\bright[2][0] ));
 sg13g2_dfrbp_1 _2179_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net360),
    .D(net42),
    .Q_N(_1113_),
    .Q(\lfsr[4] ));
 sg13g2_dfrbp_1 _2180_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net359),
    .D(net36),
    .Q_N(_1114_),
    .Q(\lfsr[5] ));
 sg13g2_dfrbp_1 _2181_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net357),
    .D(net40),
    .Q_N(_1115_),
    .Q(\lfsr_dev.lfsr[6] ));
 sg13g2_dfrbp_1 _2182_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net357),
    .D(net39),
    .Q_N(_1116_),
    .Q(\lfsr_dev.lfsr[7] ));
 sg13g2_dfrbp_1 _2183_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net357),
    .D(net38),
    .Q_N(_1117_),
    .Q(\lfsr_dev.lfsr[8] ));
 sg13g2_dfrbp_1 _2184_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net356),
    .D(net37),
    .Q_N(_1118_),
    .Q(\lfsr_dev.lfsr[9] ));
 sg13g2_dfrbp_1 _2185_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net356),
    .D(_0060_),
    .Q_N(_1097_),
    .Q(\lfsr_dev.lfsr[10] ));
 sg13g2_dfrbp_1 _2186_ (.CLK(_0108_),
    .RESET_B(net348),
    .D(_0000_),
    .Q_N(_1096_),
    .Q(\audio_mod.audio_gen.chan0.ch_counter[0] ));
 sg13g2_dfrbp_1 _2187_ (.CLK(_0109_),
    .RESET_B(net348),
    .D(_0003_),
    .Q_N(_1095_),
    .Q(\audio_mod.audio_gen.chan0.ch_counter[1] ));
 sg13g2_dfrbp_1 _2188_ (.CLK(_0110_),
    .RESET_B(net348),
    .D(_0004_),
    .Q_N(_1094_),
    .Q(\audio_mod.audio_gen.chan0.ch_counter[2] ));
 sg13g2_dfrbp_1 _2189_ (.CLK(_0111_),
    .RESET_B(net348),
    .D(_0005_),
    .Q_N(_1093_),
    .Q(\audio_mod.audio_gen.chan0.ch_counter[3] ));
 sg13g2_dfrbp_1 _2190_ (.CLK(_0112_),
    .RESET_B(net348),
    .D(_0006_),
    .Q_N(_1092_),
    .Q(\audio_mod.audio_gen.chan0.ch_counter[4] ));
 sg13g2_dfrbp_1 _2191_ (.CLK(_0113_),
    .RESET_B(net348),
    .D(_0007_),
    .Q_N(_1091_),
    .Q(\audio_mod.audio_gen.chan0.ch_counter[5] ));
 sg13g2_dfrbp_1 _2192_ (.CLK(_0114_),
    .RESET_B(net348),
    .D(_0008_),
    .Q_N(_1090_),
    .Q(\audio_mod.audio_gen.chan0.ch_counter[6] ));
 sg13g2_dfrbp_1 _2193_ (.CLK(_0115_),
    .RESET_B(net350),
    .D(_0009_),
    .Q_N(_1089_),
    .Q(\audio_mod.audio_gen.chan0.ch_counter[7] ));
 sg13g2_dfrbp_1 _2194_ (.CLK(_0116_),
    .RESET_B(net350),
    .D(_0010_),
    .Q_N(_1088_),
    .Q(\audio_mod.audio_gen.chan0.ch_counter[8] ));
 sg13g2_dfrbp_1 _2195_ (.CLK(_0117_),
    .RESET_B(net350),
    .D(_0011_),
    .Q_N(_1087_),
    .Q(\audio_mod.audio_gen.chan0.ch_counter[9] ));
 sg13g2_dfrbp_1 _2196_ (.CLK(_0118_),
    .RESET_B(net350),
    .D(_0001_),
    .Q_N(_1086_),
    .Q(\audio_mod.audio_gen.chan0.ch_counter[10] ));
 sg13g2_dfrbp_1 _2197_ (.CLK(_0119_),
    .RESET_B(net350),
    .D(_0002_),
    .Q_N(_1085_),
    .Q(\audio_mod.audio_gen.chan0.ch_counter[11] ));
 sg13g2_dfrbp_1 _2198_ (.CLK(_0120_),
    .RESET_B(net349),
    .D(_0013_),
    .Q_N(_1084_),
    .Q(\audio_mod.audio_gen.chan1.ch_counter[0] ));
 sg13g2_dfrbp_1 _2199_ (.CLK(_0121_),
    .RESET_B(net353),
    .D(_0016_),
    .Q_N(_1083_),
    .Q(\audio_mod.audio_gen.chan1.ch_counter[1] ));
 sg13g2_dfrbp_1 _2200_ (.CLK(_0122_),
    .RESET_B(net353),
    .D(_0017_),
    .Q_N(_1082_),
    .Q(\audio_mod.audio_gen.chan1.ch_counter[2] ));
 sg13g2_dfrbp_1 _2201_ (.CLK(_0123_),
    .RESET_B(net349),
    .D(_0018_),
    .Q_N(_1081_),
    .Q(\audio_mod.audio_gen.chan1.ch_counter[3] ));
 sg13g2_dfrbp_1 _2202_ (.CLK(_0124_),
    .RESET_B(net349),
    .D(_0019_),
    .Q_N(_1080_),
    .Q(\audio_mod.audio_gen.chan1.ch_counter[4] ));
 sg13g2_dfrbp_1 _2203_ (.CLK(_0125_),
    .RESET_B(net349),
    .D(_0020_),
    .Q_N(_1079_),
    .Q(\audio_mod.audio_gen.chan1.ch_counter[5] ));
 sg13g2_dfrbp_1 _2204_ (.CLK(_0126_),
    .RESET_B(net349),
    .D(_0021_),
    .Q_N(_1078_),
    .Q(\audio_mod.audio_gen.chan1.ch_counter[6] ));
 sg13g2_dfrbp_1 _2205_ (.CLK(_0127_),
    .RESET_B(net348),
    .D(_0022_),
    .Q_N(_1077_),
    .Q(\audio_mod.audio_gen.chan1.ch_counter[7] ));
 sg13g2_dfrbp_1 _2206_ (.CLK(_0128_),
    .RESET_B(net351),
    .D(_0023_),
    .Q_N(_1076_),
    .Q(\audio_mod.audio_gen.chan1.ch_counter[8] ));
 sg13g2_dfrbp_1 _2207_ (.CLK(_0129_),
    .RESET_B(net351),
    .D(_0024_),
    .Q_N(_1075_),
    .Q(\audio_mod.audio_gen.chan1.ch_counter[9] ));
 sg13g2_dfrbp_1 _2208_ (.CLK(_0130_),
    .RESET_B(net353),
    .D(_0014_),
    .Q_N(_1074_),
    .Q(\audio_mod.audio_gen.chan1.ch_counter[10] ));
 sg13g2_dfrbp_1 _2209_ (.CLK(_0131_),
    .RESET_B(net353),
    .D(_0015_),
    .Q_N(_1073_),
    .Q(\audio_mod.audio_gen.chan1.ch_counter[11] ));
 sg13g2_dfrbp_1 _2210_ (.CLK(_0132_),
    .RESET_B(net358),
    .D(_0162_),
    .Q_N(_0012_),
    .Q(\audio_mod.audio_gen.ch0_state ));
 sg13g2_dfrbp_1 _2211_ (.CLK(_0133_),
    .RESET_B(net354),
    .D(_0026_),
    .Q_N(_1072_),
    .Q(\audio_mod.audio_gen.chan2.ch_counter[0] ));
 sg13g2_dfrbp_1 _2212_ (.CLK(_0134_),
    .RESET_B(net354),
    .D(_0029_),
    .Q_N(_1071_),
    .Q(\audio_mod.audio_gen.chan2.ch_counter[1] ));
 sg13g2_dfrbp_1 _2213_ (.CLK(_0135_),
    .RESET_B(net353),
    .D(_0030_),
    .Q_N(_1070_),
    .Q(\audio_mod.audio_gen.chan2.ch_counter[2] ));
 sg13g2_dfrbp_1 _2214_ (.CLK(_0136_),
    .RESET_B(net353),
    .D(_0031_),
    .Q_N(_1069_),
    .Q(\audio_mod.audio_gen.chan2.ch_counter[3] ));
 sg13g2_dfrbp_1 _2215_ (.CLK(_0137_),
    .RESET_B(net353),
    .D(_0032_),
    .Q_N(_1068_),
    .Q(\audio_mod.audio_gen.chan2.ch_counter[4] ));
 sg13g2_dfrbp_1 _2216_ (.CLK(_0138_),
    .RESET_B(net353),
    .D(_0033_),
    .Q_N(_1067_),
    .Q(\audio_mod.audio_gen.chan2.ch_counter[5] ));
 sg13g2_dfrbp_1 _2217_ (.CLK(_0139_),
    .RESET_B(net363),
    .D(_0034_),
    .Q_N(_1066_),
    .Q(\audio_mod.audio_gen.chan2.ch_counter[6] ));
 sg13g2_dfrbp_1 _2218_ (.CLK(_0140_),
    .RESET_B(net363),
    .D(_0035_),
    .Q_N(_1065_),
    .Q(\audio_mod.audio_gen.chan2.ch_counter[7] ));
 sg13g2_dfrbp_1 _2219_ (.CLK(_0141_),
    .RESET_B(net363),
    .D(_0036_),
    .Q_N(_1064_),
    .Q(\audio_mod.audio_gen.chan2.ch_counter[8] ));
 sg13g2_dfrbp_1 _2220_ (.CLK(_0142_),
    .RESET_B(net363),
    .D(_0037_),
    .Q_N(_1063_),
    .Q(\audio_mod.audio_gen.chan2.ch_counter[9] ));
 sg13g2_dfrbp_1 _2221_ (.CLK(_0143_),
    .RESET_B(net354),
    .D(_0027_),
    .Q_N(_1062_),
    .Q(\audio_mod.audio_gen.chan2.ch_counter[10] ));
 sg13g2_dfrbp_1 _2222_ (.CLK(_0144_),
    .RESET_B(net354),
    .D(_0028_),
    .Q_N(_0074_),
    .Q(\audio_mod.audio_gen.chan2.ch_counter[11] ));
 sg13g2_dfrbp_1 _2223_ (.CLK(_0145_),
    .RESET_B(net351),
    .D(_0163_),
    .Q_N(_0025_),
    .Q(\audio_mod.audio_gen.ch1_state ));
 sg13g2_dfrbp_1 _2224_ (.CLK(_0146_),
    .RESET_B(net355),
    .D(_0039_),
    .Q_N(_1061_),
    .Q(\audio_mod.audio_gen.chan3.ch_counter[0] ));
 sg13g2_dfrbp_1 _2225_ (.CLK(_0147_),
    .RESET_B(net355),
    .D(_0042_),
    .Q_N(_1060_),
    .Q(\audio_mod.audio_gen.chan3.ch_counter[1] ));
 sg13g2_dfrbp_1 _2226_ (.CLK(_0148_),
    .RESET_B(net355),
    .D(_0043_),
    .Q_N(_1059_),
    .Q(\audio_mod.audio_gen.chan3.ch_counter[2] ));
 sg13g2_dfrbp_1 _2227_ (.CLK(_0149_),
    .RESET_B(net355),
    .D(_0044_),
    .Q_N(_1058_),
    .Q(\audio_mod.audio_gen.chan3.ch_counter[3] ));
 sg13g2_dfrbp_1 _2228_ (.CLK(_0150_),
    .RESET_B(net355),
    .D(_0045_),
    .Q_N(_1057_),
    .Q(\audio_mod.audio_gen.chan3.ch_counter[4] ));
 sg13g2_dfrbp_1 _2229_ (.CLK(_0151_),
    .RESET_B(net355),
    .D(_0046_),
    .Q_N(_1056_),
    .Q(\audio_mod.audio_gen.chan3.ch_counter[5] ));
 sg13g2_dfrbp_1 _2230_ (.CLK(_0152_),
    .RESET_B(net358),
    .D(_0047_),
    .Q_N(_1055_),
    .Q(\audio_mod.audio_gen.chan3.ch_counter[6] ));
 sg13g2_dfrbp_1 _2231_ (.CLK(_0153_),
    .RESET_B(net351),
    .D(_0048_),
    .Q_N(_1054_),
    .Q(\audio_mod.audio_gen.chan3.ch_counter[7] ));
 sg13g2_dfrbp_1 _2232_ (.CLK(_0154_),
    .RESET_B(net355),
    .D(_0049_),
    .Q_N(_1053_),
    .Q(\audio_mod.audio_gen.chan3.ch_counter[8] ));
 sg13g2_dfrbp_1 _2233_ (.CLK(_0155_),
    .RESET_B(net350),
    .D(_0050_),
    .Q_N(_1052_),
    .Q(\audio_mod.audio_gen.chan3.ch_counter[9] ));
 sg13g2_dfrbp_1 _2234_ (.CLK(_0156_),
    .RESET_B(net350),
    .D(_0040_),
    .Q_N(_1051_),
    .Q(\audio_mod.audio_gen.chan3.ch_counter[10] ));
 sg13g2_dfrbp_1 _2235_ (.CLK(_0157_),
    .RESET_B(net350),
    .D(_0041_),
    .Q_N(_1050_),
    .Q(\audio_mod.audio_gen.chan3.ch_counter[11] ));
 sg13g2_dfrbp_1 _2236_ (.CLK(_0158_),
    .RESET_B(net361),
    .D(_0164_),
    .Q_N(_0038_),
    .Q(\audio_mod.audio_gen.ch2_state ));
 sg13g2_dfrbp_1 _2237_ (.CLK(net288),
    .RESET_B(net354),
    .D(_0051_),
    .Q_N(_1049_),
    .Q(\audio_mod.seq.seq_clock[0] ));
 sg13g2_dfrbp_1 _2238_ (.CLK(net288),
    .RESET_B(net354),
    .D(_0052_),
    .Q_N(_1048_),
    .Q(\audio_mod.seq.seq_clock[1] ));
 sg13g2_dfrbp_1 _2239_ (.CLK(net288),
    .RESET_B(net354),
    .D(_0053_),
    .Q_N(_1047_),
    .Q(\audio_mod.seq.seq_clock[2] ));
 sg13g2_dfrbp_1 _2240_ (.CLK(net288),
    .RESET_B(net351),
    .D(_0054_),
    .Q_N(_1046_),
    .Q(\audio_mod.seq.seq_clock[3] ));
 sg13g2_dfrbp_1 _2241_ (.CLK(_1099_),
    .RESET_B(net360),
    .D(_0165_),
    .Q_N(_0064_),
    .Q(\background_color[0] ));
 sg13g2_dfrbp_1 _2242_ (.CLK(_1099_),
    .RESET_B(net360),
    .D(_0166_),
    .Q_N(_0065_),
    .Q(\background_color[1] ));
 sg13g2_dfrbp_1 _2243_ (.CLK(_1099_),
    .RESET_B(net359),
    .D(_0167_),
    .Q_N(_0063_),
    .Q(\background_color[2] ));
 sg13g2_dfrbp_1 _2244_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net27),
    .D(net62),
    .Q_N(uo_out[7]),
    .Q(hsync));
 sg13g2_dfrbp_1 _2245_ (.CLK(_0159_),
    .RESET_B(net355),
    .D(_0168_),
    .Q_N(_1119_),
    .Q(\audio_mod.audio_gen.ch3_state ));
 sg13g2_dfrbp_1 _2246_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net25),
    .D(net50),
    .Q_N(uo_out[3]),
    .Q(\clock_gen.vsync ));
 sg13g2_dfrbp_1 _2247_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net24),
    .D(_0169_),
    .Q_N(_0100_),
    .Q(\hvsync_gen.vpos[0] ));
 sg13g2_dfrbp_1 _2248_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net22),
    .D(_0170_),
    .Q_N(_1045_),
    .Q(\hvsync_gen.vpos[1] ));
 sg13g2_dfrbp_1 _2249_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net20),
    .D(_0171_),
    .Q_N(_0070_),
    .Q(\hvsync_gen.vpos[2] ));
 sg13g2_dfrbp_1 _2250_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net18),
    .D(_0172_),
    .Q_N(_0066_),
    .Q(\hvsync_gen.vpos[3] ));
 sg13g2_dfrbp_1 _2251_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net17),
    .D(_0173_),
    .Q_N(_0071_),
    .Q(\hvsync_gen.vpos[4] ));
 sg13g2_dfrbp_1 _2252_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net15),
    .D(_0174_),
    .Q_N(_1044_),
    .Q(\hvsync_gen.vpos[5] ));
 sg13g2_dfrbp_1 _2253_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net14),
    .D(_0175_),
    .Q_N(_0067_),
    .Q(\hvsync_gen.vpos[6] ));
 sg13g2_dfrbp_1 _2254_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net13),
    .D(_0176_),
    .Q_N(_1043_),
    .Q(\hvsync_gen.vpos[7] ));
 sg13g2_dfrbp_1 _2255_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net11),
    .D(_0177_),
    .Q_N(_0069_),
    .Q(\hvsync_gen.vpos[8] ));
 sg13g2_dfrbp_1 _2256_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net9),
    .D(net59),
    .Q_N(_0068_),
    .Q(\hvsync_gen.vpos[9] ));
 sg13g2_dfrbp_1 _2257_ (.CLK(net288),
    .RESET_B(net359),
    .D(_0179_),
    .Q_N(\stage_seq_inst.stage_timer[0] ),
    .Q(_0102_));
 sg13g2_dfrbp_1 _2258_ (.CLK(net288),
    .RESET_B(net359),
    .D(_0180_),
    .Q_N(\stage_seq_inst.stage_timer[1] ),
    .Q(_0103_));
 sg13g2_dfrbp_1 _2259_ (.CLK(net288),
    .RESET_B(net359),
    .D(_0181_),
    .Q_N(_1042_),
    .Q(\stage_seq_inst.stage_timer[2] ));
 sg13g2_dfrbp_1 _2260_ (.CLK(net288),
    .RESET_B(net357),
    .D(_0182_),
    .Q_N(_1041_),
    .Q(\stage_seq_inst.stage_timer[3] ));
 sg13g2_dfrbp_1 _2261_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net12),
    .D(_0183_),
    .Q_N(_0099_),
    .Q(\hpos[0] ));
 sg13g2_dfrbp_1 _2262_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net10),
    .D(_0184_),
    .Q_N(_1040_),
    .Q(\hpos[1] ));
 sg13g2_dfrbp_1 _2263_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net30),
    .D(_0185_),
    .Q_N(_1039_),
    .Q(\hpos[2] ));
 sg13g2_dfrbp_1 _2264_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net29),
    .D(_0186_),
    .Q_N(_0076_),
    .Q(\hpos[3] ));
 sg13g2_dfrbp_1 _2265_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net28),
    .D(_0187_),
    .Q_N(_0077_),
    .Q(\hpos[4] ));
 sg13g2_dfrbp_1 _2266_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net26),
    .D(_0188_),
    .Q_N(_0078_),
    .Q(\hpos[5] ));
 sg13g2_dfrbp_1 _2267_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net23),
    .D(_0189_),
    .Q_N(_0079_),
    .Q(\hpos[6] ));
 sg13g2_dfrbp_1 _2268_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net21),
    .D(_0190_),
    .Q_N(_0080_),
    .Q(\hpos[7] ));
 sg13g2_dfrbp_1 _2269_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net19),
    .D(_0191_),
    .Q_N(_0081_),
    .Q(\hpos[8] ));
 sg13g2_dfrbp_1 _2270_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net16),
    .D(net78),
    .Q_N(_0075_),
    .Q(\hpos[9] ));
 sg13g2_tiehi _2262__10 (.L_HI(net10));
 sg13g2_tiehi _2255__11 (.L_HI(net11));
 sg13g2_tiehi _2261__12 (.L_HI(net12));
 sg13g2_tiehi _2254__13 (.L_HI(net13));
 sg13g2_tiehi _2253__14 (.L_HI(net14));
 sg13g2_tiehi _2252__15 (.L_HI(net15));
 sg13g2_tiehi _2270__16 (.L_HI(net16));
 sg13g2_tiehi _2251__17 (.L_HI(net17));
 sg13g2_tiehi _2250__18 (.L_HI(net18));
 sg13g2_tiehi _2269__19 (.L_HI(net19));
 sg13g2_tiehi _2249__20 (.L_HI(net20));
 sg13g2_tiehi _2268__21 (.L_HI(net21));
 sg13g2_tiehi _2248__22 (.L_HI(net22));
 sg13g2_tiehi _2267__23 (.L_HI(net23));
 sg13g2_tiehi _2247__24 (.L_HI(net24));
 sg13g2_tiehi _2246__25 (.L_HI(net25));
 sg13g2_tiehi _2266__26 (.L_HI(net26));
 sg13g2_tiehi _2244__27 (.L_HI(net27));
 sg13g2_tiehi _2265__28 (.L_HI(net28));
 sg13g2_tiehi _2264__29 (.L_HI(net29));
 sg13g2_tiehi _2263__30 (.L_HI(net30));
 sg13g2_tiehi tt_um_bytex64_munch_31 (.L_HI(net31));
 sg13g2_tiehi tt_um_bytex64_munch_32 (.L_HI(net32));
 sg13g2_tiehi tt_um_bytex64_munch_33 (.L_HI(net33));
 sg13g2_tiehi tt_um_bytex64_munch_34 (.L_HI(net34));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_bytex64_munch_2 (.L_LO(net2));
 sg13g2_tielo tt_um_bytex64_munch_3 (.L_LO(net3));
 sg13g2_tielo tt_um_bytex64_munch_4 (.L_LO(net4));
 sg13g2_tielo tt_um_bytex64_munch_5 (.L_LO(net5));
 sg13g2_tielo tt_um_bytex64_munch_6 (.L_LO(net6));
 sg13g2_tielo tt_um_bytex64_munch_7 (.L_LO(net7));
 sg13g2_tielo tt_um_bytex64_munch_8 (.L_LO(net8));
 sg13g2_tiehi _2256__9 (.L_HI(net9));
 sg13g2_buf_2 _2305_ (.A(\audio_mod.pattern_clock[1] ),
    .X(uio_out[4]));
 sg13g2_buf_2 _2306_ (.A(net292),
    .X(uio_out[5]));
 sg13g2_buf_2 _2307_ (.A(net289),
    .X(uio_out[6]));
 sg13g2_buf_1 _2308_ (.A(audio),
    .X(uio_out[7]));
 sg13g2_buf_2 fanout277 (.A(net278),
    .X(net277));
 sg13g2_buf_2 fanout278 (.A(_0473_),
    .X(net278));
 sg13g2_buf_2 fanout279 (.A(net280),
    .X(net279));
 sg13g2_buf_2 fanout280 (.A(_0532_),
    .X(net280));
 sg13g2_buf_2 fanout281 (.A(_0513_),
    .X(net281));
 sg13g2_buf_2 fanout282 (.A(_0725_),
    .X(net282));
 sg13g2_buf_4 fanout283 (.X(net283),
    .A(_0485_));
 sg13g2_buf_4 fanout284 (.X(net284),
    .A(_0483_));
 sg13g2_buf_2 fanout285 (.A(_0679_),
    .X(net285));
 sg13g2_buf_2 fanout286 (.A(net287),
    .X(net286));
 sg13g2_buf_2 fanout287 (.A(_0329_),
    .X(net287));
 sg13g2_buf_4 fanout288 (.X(net288),
    .A(_1104_));
 sg13g2_buf_4 fanout289 (.X(net289),
    .A(\audio_mod.pattern_clock[3] ));
 sg13g2_buf_2 fanout290 (.A(\audio_mod.pattern_clock[3] ),
    .X(net290));
 sg13g2_buf_2 fanout291 (.A(net292),
    .X(net291));
 sg13g2_buf_4 fanout292 (.X(net292),
    .A(\audio_mod.pattern_clock[2] ));
 sg13g2_buf_2 fanout293 (.A(\audio_mod.pattern_clock[1] ),
    .X(net293));
 sg13g2_buf_2 fanout294 (.A(\audio_mod.pattern_clock[0] ),
    .X(net294));
 sg13g2_buf_2 fanout295 (.A(_0954_),
    .X(net295));
 sg13g2_buf_2 fanout296 (.A(_0947_),
    .X(net296));
 sg13g2_buf_2 fanout297 (.A(_0619_),
    .X(net297));
 sg13g2_buf_2 fanout298 (.A(\atick_clock[1] ),
    .X(net298));
 sg13g2_buf_2 fanout299 (.A(\atick_clock[1] ),
    .X(net299));
 sg13g2_buf_2 fanout300 (.A(\atick_clock[0] ),
    .X(net300));
 sg13g2_buf_1 fanout301 (.A(\atick_clock[0] ),
    .X(net301));
 sg13g2_buf_2 fanout302 (.A(\clock_gen.r_atick_clock[0] ),
    .X(net302));
 sg13g2_buf_4 fanout303 (.X(net303),
    .A(\counter[3] ));
 sg13g2_buf_4 fanout304 (.X(net304),
    .A(\counter[2] ));
 sg13g2_buf_1 fanout305 (.A(\counter[2] ),
    .X(net305));
 sg13g2_buf_2 fanout306 (.A(\counter[1] ),
    .X(net306));
 sg13g2_buf_2 fanout307 (.A(net309),
    .X(net307));
 sg13g2_buf_1 fanout308 (.A(net309),
    .X(net308));
 sg13g2_buf_2 fanout309 (.A(net312),
    .X(net309));
 sg13g2_buf_2 fanout310 (.A(net311),
    .X(net310));
 sg13g2_buf_2 fanout311 (.A(net312),
    .X(net311));
 sg13g2_buf_2 fanout312 (.A(net315),
    .X(net312));
 sg13g2_buf_2 fanout313 (.A(net315),
    .X(net313));
 sg13g2_buf_2 fanout314 (.A(net315),
    .X(net314));
 sg13g2_buf_2 fanout315 (.A(_0323_),
    .X(net315));
 sg13g2_buf_2 fanout316 (.A(net77),
    .X(net316));
 sg13g2_buf_4 fanout317 (.X(net317),
    .A(_0080_));
 sg13g2_buf_4 fanout318 (.X(net318),
    .A(\hpos[7] ));
 sg13g2_buf_2 fanout319 (.A(net82),
    .X(net319));
 sg13g2_buf_2 fanout320 (.A(\hpos[1] ),
    .X(net320));
 sg13g2_buf_4 fanout321 (.X(net321),
    .A(net79));
 sg13g2_buf_4 fanout322 (.X(net322),
    .A(net323));
 sg13g2_buf_2 fanout323 (.A(\hvsync_gen.vpos[7] ),
    .X(net323));
 sg13g2_buf_2 fanout324 (.A(net325),
    .X(net324));
 sg13g2_buf_2 fanout325 (.A(\hvsync_gen.vpos[5] ),
    .X(net325));
 sg13g2_buf_4 fanout326 (.X(net326),
    .A(net49));
 sg13g2_buf_2 fanout327 (.A(\hvsync_gen.vpos[3] ),
    .X(net327));
 sg13g2_buf_4 fanout328 (.X(net328),
    .A(\clock_gen.vsync ));
 sg13g2_buf_2 fanout329 (.A(net331),
    .X(net329));
 sg13g2_buf_1 fanout330 (.A(net331),
    .X(net330));
 sg13g2_buf_2 fanout331 (.A(net334),
    .X(net331));
 sg13g2_buf_2 fanout332 (.A(net333),
    .X(net332));
 sg13g2_buf_2 fanout333 (.A(net334),
    .X(net333));
 sg13g2_buf_2 fanout334 (.A(\audio_mod.audio_gen.pwm_clock[5] ),
    .X(net334));
 sg13g2_buf_2 fanout335 (.A(net337),
    .X(net335));
 sg13g2_buf_2 fanout336 (.A(net337),
    .X(net336));
 sg13g2_buf_2 fanout337 (.A(\audio_mod.audio_gen.pwm_clock[5] ),
    .X(net337));
 sg13g2_buf_2 fanout338 (.A(net340),
    .X(net338));
 sg13g2_buf_1 fanout339 (.A(net340),
    .X(net339));
 sg13g2_buf_2 fanout340 (.A(net343),
    .X(net340));
 sg13g2_buf_2 fanout341 (.A(net342),
    .X(net341));
 sg13g2_buf_2 fanout342 (.A(net343),
    .X(net342));
 sg13g2_buf_2 fanout343 (.A(net347),
    .X(net343));
 sg13g2_buf_2 fanout344 (.A(net346),
    .X(net344));
 sg13g2_buf_2 fanout345 (.A(net347),
    .X(net345));
 sg13g2_buf_1 fanout346 (.A(net347),
    .X(net346));
 sg13g2_buf_2 fanout347 (.A(\audio_mod.audio_gen.pwm_clock[2] ),
    .X(net347));
 sg13g2_buf_4 fanout348 (.X(net348),
    .A(net352));
 sg13g2_buf_2 fanout349 (.A(net352),
    .X(net349));
 sg13g2_buf_4 fanout350 (.X(net350),
    .A(net352));
 sg13g2_buf_2 fanout351 (.A(net352),
    .X(net351));
 sg13g2_buf_2 fanout352 (.A(net362),
    .X(net352));
 sg13g2_buf_4 fanout353 (.X(net353),
    .A(net354));
 sg13g2_buf_4 fanout354 (.X(net354),
    .A(net362));
 sg13g2_buf_4 fanout355 (.X(net355),
    .A(net358));
 sg13g2_buf_4 fanout356 (.X(net356),
    .A(net357));
 sg13g2_buf_4 fanout357 (.X(net357),
    .A(net358));
 sg13g2_buf_2 fanout358 (.A(net362),
    .X(net358));
 sg13g2_buf_4 fanout359 (.X(net359),
    .A(net362));
 sg13g2_buf_4 fanout360 (.X(net360),
    .A(net361));
 sg13g2_buf_4 fanout361 (.X(net361),
    .A(net362));
 sg13g2_buf_2 fanout362 (.A(rst_n),
    .X(net362));
 sg13g2_buf_4 fanout363 (.X(net363),
    .A(net365));
 sg13g2_buf_2 fanout364 (.A(net365),
    .X(net364));
 sg13g2_buf_4 fanout365 (.X(net365),
    .A(rst_n));
 sg13g2_tielo tt_um_bytex64_munch_1 (.L_LO(net1));
 sg13g2_buf_2 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sg13g2_buf_2 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sg13g2_buf_2 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sg13g2_buf_2 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sg13g2_buf_2 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sg13g2_buf_2 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sg13g2_buf_2 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sg13g2_buf_2 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_3_7__leaf_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(_1036_),
    .X(net35));
 sg13g2_dlygate4sd3_1 hold2 (.A(\lfsr_dev.lfsr[6] ),
    .X(net36));
 sg13g2_dlygate4sd3_1 hold3 (.A(\lfsr_dev.lfsr[10] ),
    .X(net37));
 sg13g2_dlygate4sd3_1 hold4 (.A(\lfsr_dev.lfsr[9] ),
    .X(net38));
 sg13g2_dlygate4sd3_1 hold5 (.A(\lfsr_dev.lfsr[8] ),
    .X(net39));
 sg13g2_dlygate4sd3_1 hold6 (.A(\lfsr_dev.lfsr[7] ),
    .X(net40));
 sg13g2_dlygate4sd3_1 hold7 (.A(\lfsr[4] ),
    .X(net41));
 sg13g2_dlygate4sd3_1 hold8 (.A(\lfsr[5] ),
    .X(net42));
 sg13g2_dlygate4sd3_1 hold9 (.A(_0099_),
    .X(net43));
 sg13g2_dlygate4sd3_1 hold10 (.A(\lfsr[1] ),
    .X(net44));
 sg13g2_dlygate4sd3_1 hold11 (.A(_0100_),
    .X(net45));
 sg13g2_dlygate4sd3_1 hold12 (.A(_0337_),
    .X(net46));
 sg13g2_dlygate4sd3_1 hold13 (.A(\bright[2][0] ),
    .X(net47));
 sg13g2_dlygate4sd3_1 hold14 (.A(\lfsr[2] ),
    .X(net48));
 sg13g2_dlygate4sd3_1 hold15 (.A(\hvsync_gen.vpos[4] ),
    .X(net49));
 sg13g2_dlygate4sd3_1 hold16 (.A(_0059_),
    .X(net50));
 sg13g2_dlygate4sd3_1 hold17 (.A(\audio_mod.audio_gen.chan3.rng ),
    .X(net51));
 sg13g2_dlygate4sd3_1 hold18 (.A(\audio_mod.audio_gen.pwm_clock[0] ),
    .X(net52));
 sg13g2_dlygate4sd3_1 hold19 (.A(_0091_),
    .X(net53));
 sg13g2_dlygate4sd3_1 hold20 (.A(\audio_mod.audio_gen.pwm_clock[4] ),
    .X(net54));
 sg13g2_dlygate4sd3_1 hold21 (.A(_0094_),
    .X(net55));
 sg13g2_dlygate4sd3_1 hold22 (.A(\audio_mod.audio_gen.pwm_clock[3] ),
    .X(net56));
 sg13g2_dlygate4sd3_1 hold23 (.A(_0093_),
    .X(net57));
 sg13g2_dlygate4sd3_1 hold24 (.A(\hvsync_gen.vpos[9] ),
    .X(net58));
 sg13g2_dlygate4sd3_1 hold25 (.A(_0178_),
    .X(net59));
 sg13g2_dlygate4sd3_1 hold26 (.A(_0075_),
    .X(net60));
 sg13g2_dlygate4sd3_1 hold27 (.A(_0618_),
    .X(net61));
 sg13g2_dlygate4sd3_1 hold28 (.A(_0058_),
    .X(net62));
 sg13g2_dlygate4sd3_1 hold29 (.A(_0070_),
    .X(net63));
 sg13g2_dlygate4sd3_1 hold30 (.A(_0343_),
    .X(net64));
 sg13g2_dlygate4sd3_1 hold31 (.A(\hvsync_gen.vpos[1] ),
    .X(net65));
 sg13g2_dlygate4sd3_1 hold32 (.A(\hpos[6] ),
    .X(net66));
 sg13g2_dlygate4sd3_1 hold33 (.A(\hvsync_gen.vpos[6] ),
    .X(net67));
 sg13g2_dlygate4sd3_1 hold34 (.A(\hpos[8] ),
    .X(net68));
 sg13g2_dlygate4sd3_1 hold35 (.A(_0079_),
    .X(net69));
 sg13g2_dlygate4sd3_1 hold36 (.A(_0367_),
    .X(net70));
 sg13g2_dlygate4sd3_1 hold37 (.A(_0071_),
    .X(net71));
 sg13g2_dlygate4sd3_1 hold38 (.A(\hpos[5] ),
    .X(net72));
 sg13g2_dlygate4sd3_1 hold39 (.A(_0363_),
    .X(net73));
 sg13g2_dlygate4sd3_1 hold40 (.A(\audio_mod.audio_gen.pwm_clock[1] ),
    .X(net74));
 sg13g2_dlygate4sd3_1 hold41 (.A(\hvsync_gen.vpos[2] ),
    .X(net75));
 sg13g2_dlygate4sd3_1 hold42 (.A(\hpos[3] ),
    .X(net76));
 sg13g2_dlygate4sd3_1 hold43 (.A(\hpos[9] ),
    .X(net77));
 sg13g2_dlygate4sd3_1 hold44 (.A(_0192_),
    .X(net78));
 sg13g2_dlygate4sd3_1 hold45 (.A(\hvsync_gen.vpos[8] ),
    .X(net79));
 sg13g2_dlygate4sd3_1 hold46 (.A(\hpos[4] ),
    .X(net80));
 sg13g2_dlygate4sd3_1 hold47 (.A(\hpos[0] ),
    .X(net81));
 sg13g2_dlygate4sd3_1 hold48 (.A(\hpos[2] ),
    .X(net82));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_fill_1 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_17 ();
 sg13g2_decap_4 FILLER_2_24 ();
 sg13g2_fill_1 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_37 ();
 sg13g2_decap_8 FILLER_2_44 ();
 sg13g2_fill_2 FILLER_2_56 ();
 sg13g2_fill_2 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_134 ();
 sg13g2_fill_1 FILLER_2_141 ();
 sg13g2_decap_8 FILLER_2_151 ();
 sg13g2_decap_8 FILLER_2_158 ();
 sg13g2_decap_8 FILLER_2_165 ();
 sg13g2_decap_8 FILLER_2_172 ();
 sg13g2_decap_8 FILLER_2_179 ();
 sg13g2_decap_8 FILLER_2_186 ();
 sg13g2_decap_8 FILLER_2_193 ();
 sg13g2_decap_8 FILLER_2_200 ();
 sg13g2_decap_8 FILLER_2_207 ();
 sg13g2_decap_8 FILLER_2_214 ();
 sg13g2_decap_8 FILLER_2_221 ();
 sg13g2_decap_8 FILLER_2_228 ();
 sg13g2_decap_8 FILLER_2_235 ();
 sg13g2_decap_8 FILLER_2_242 ();
 sg13g2_decap_8 FILLER_2_249 ();
 sg13g2_decap_8 FILLER_2_256 ();
 sg13g2_decap_8 FILLER_2_263 ();
 sg13g2_decap_8 FILLER_2_270 ();
 sg13g2_decap_8 FILLER_2_277 ();
 sg13g2_decap_8 FILLER_2_284 ();
 sg13g2_decap_8 FILLER_2_291 ();
 sg13g2_decap_8 FILLER_2_298 ();
 sg13g2_decap_8 FILLER_2_305 ();
 sg13g2_decap_8 FILLER_2_312 ();
 sg13g2_decap_8 FILLER_2_319 ();
 sg13g2_decap_8 FILLER_2_326 ();
 sg13g2_decap_8 FILLER_2_333 ();
 sg13g2_decap_8 FILLER_2_340 ();
 sg13g2_decap_8 FILLER_2_347 ();
 sg13g2_decap_8 FILLER_2_354 ();
 sg13g2_decap_8 FILLER_2_361 ();
 sg13g2_decap_8 FILLER_2_368 ();
 sg13g2_decap_8 FILLER_2_375 ();
 sg13g2_decap_8 FILLER_2_382 ();
 sg13g2_decap_8 FILLER_2_389 ();
 sg13g2_decap_8 FILLER_2_396 ();
 sg13g2_decap_4 FILLER_2_403 ();
 sg13g2_fill_2 FILLER_2_407 ();
 sg13g2_fill_2 FILLER_3_0 ();
 sg13g2_fill_1 FILLER_3_28 ();
 sg13g2_fill_2 FILLER_3_60 ();
 sg13g2_decap_8 FILLER_3_79 ();
 sg13g2_decap_8 FILLER_3_86 ();
 sg13g2_decap_4 FILLER_3_93 ();
 sg13g2_fill_2 FILLER_3_97 ();
 sg13g2_decap_8 FILLER_3_178 ();
 sg13g2_decap_8 FILLER_3_185 ();
 sg13g2_decap_8 FILLER_3_192 ();
 sg13g2_decap_8 FILLER_3_199 ();
 sg13g2_decap_8 FILLER_3_206 ();
 sg13g2_decap_8 FILLER_3_213 ();
 sg13g2_decap_8 FILLER_3_220 ();
 sg13g2_decap_8 FILLER_3_227 ();
 sg13g2_decap_8 FILLER_3_234 ();
 sg13g2_decap_8 FILLER_3_241 ();
 sg13g2_decap_8 FILLER_3_248 ();
 sg13g2_decap_8 FILLER_3_255 ();
 sg13g2_decap_8 FILLER_3_262 ();
 sg13g2_decap_8 FILLER_3_269 ();
 sg13g2_decap_8 FILLER_3_276 ();
 sg13g2_decap_8 FILLER_3_283 ();
 sg13g2_decap_8 FILLER_3_290 ();
 sg13g2_decap_8 FILLER_3_297 ();
 sg13g2_decap_8 FILLER_3_304 ();
 sg13g2_decap_8 FILLER_3_311 ();
 sg13g2_decap_8 FILLER_3_318 ();
 sg13g2_decap_8 FILLER_3_325 ();
 sg13g2_decap_8 FILLER_3_332 ();
 sg13g2_decap_8 FILLER_3_339 ();
 sg13g2_decap_8 FILLER_3_346 ();
 sg13g2_decap_8 FILLER_3_353 ();
 sg13g2_decap_8 FILLER_3_360 ();
 sg13g2_decap_8 FILLER_3_367 ();
 sg13g2_decap_8 FILLER_3_374 ();
 sg13g2_decap_8 FILLER_3_381 ();
 sg13g2_decap_8 FILLER_3_388 ();
 sg13g2_decap_8 FILLER_3_395 ();
 sg13g2_decap_8 FILLER_3_402 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_fill_2 FILLER_4_28 ();
 sg13g2_decap_4 FILLER_4_39 ();
 sg13g2_fill_2 FILLER_4_43 ();
 sg13g2_fill_1 FILLER_4_55 ();
 sg13g2_fill_2 FILLER_4_92 ();
 sg13g2_fill_1 FILLER_4_94 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_4 FILLER_4_112 ();
 sg13g2_fill_2 FILLER_4_125 ();
 sg13g2_decap_4 FILLER_4_136 ();
 sg13g2_fill_1 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_187 ();
 sg13g2_decap_8 FILLER_4_194 ();
 sg13g2_decap_8 FILLER_4_201 ();
 sg13g2_decap_8 FILLER_4_208 ();
 sg13g2_decap_8 FILLER_4_215 ();
 sg13g2_decap_8 FILLER_4_222 ();
 sg13g2_decap_8 FILLER_4_229 ();
 sg13g2_decap_8 FILLER_4_236 ();
 sg13g2_decap_8 FILLER_4_243 ();
 sg13g2_decap_8 FILLER_4_250 ();
 sg13g2_decap_8 FILLER_4_257 ();
 sg13g2_decap_8 FILLER_4_264 ();
 sg13g2_decap_8 FILLER_4_271 ();
 sg13g2_decap_8 FILLER_4_278 ();
 sg13g2_decap_8 FILLER_4_285 ();
 sg13g2_decap_8 FILLER_4_292 ();
 sg13g2_decap_8 FILLER_4_299 ();
 sg13g2_decap_8 FILLER_4_306 ();
 sg13g2_decap_8 FILLER_4_313 ();
 sg13g2_decap_8 FILLER_4_320 ();
 sg13g2_decap_8 FILLER_4_327 ();
 sg13g2_decap_8 FILLER_4_334 ();
 sg13g2_decap_8 FILLER_4_341 ();
 sg13g2_decap_8 FILLER_4_348 ();
 sg13g2_decap_8 FILLER_4_355 ();
 sg13g2_decap_8 FILLER_4_362 ();
 sg13g2_decap_8 FILLER_4_369 ();
 sg13g2_decap_8 FILLER_4_376 ();
 sg13g2_decap_8 FILLER_4_383 ();
 sg13g2_decap_8 FILLER_4_390 ();
 sg13g2_decap_8 FILLER_4_397 ();
 sg13g2_decap_4 FILLER_4_404 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_fill_2 FILLER_5_0 ();
 sg13g2_fill_1 FILLER_5_2 ();
 sg13g2_fill_1 FILLER_5_47 ();
 sg13g2_decap_8 FILLER_5_82 ();
 sg13g2_fill_1 FILLER_5_89 ();
 sg13g2_fill_2 FILLER_5_103 ();
 sg13g2_fill_1 FILLER_5_105 ();
 sg13g2_fill_2 FILLER_5_114 ();
 sg13g2_decap_8 FILLER_5_176 ();
 sg13g2_decap_8 FILLER_5_183 ();
 sg13g2_decap_8 FILLER_5_190 ();
 sg13g2_decap_8 FILLER_5_197 ();
 sg13g2_decap_8 FILLER_5_204 ();
 sg13g2_decap_8 FILLER_5_211 ();
 sg13g2_decap_8 FILLER_5_218 ();
 sg13g2_decap_8 FILLER_5_225 ();
 sg13g2_decap_8 FILLER_5_232 ();
 sg13g2_decap_8 FILLER_5_239 ();
 sg13g2_decap_8 FILLER_5_246 ();
 sg13g2_decap_8 FILLER_5_253 ();
 sg13g2_decap_8 FILLER_5_260 ();
 sg13g2_decap_8 FILLER_5_267 ();
 sg13g2_decap_8 FILLER_5_274 ();
 sg13g2_decap_8 FILLER_5_281 ();
 sg13g2_decap_8 FILLER_5_288 ();
 sg13g2_decap_8 FILLER_5_295 ();
 sg13g2_decap_8 FILLER_5_302 ();
 sg13g2_decap_8 FILLER_5_309 ();
 sg13g2_decap_8 FILLER_5_316 ();
 sg13g2_decap_8 FILLER_5_323 ();
 sg13g2_decap_8 FILLER_5_330 ();
 sg13g2_decap_8 FILLER_5_337 ();
 sg13g2_decap_8 FILLER_5_344 ();
 sg13g2_decap_8 FILLER_5_351 ();
 sg13g2_decap_8 FILLER_5_358 ();
 sg13g2_decap_8 FILLER_5_365 ();
 sg13g2_decap_8 FILLER_5_372 ();
 sg13g2_decap_8 FILLER_5_379 ();
 sg13g2_decap_8 FILLER_5_386 ();
 sg13g2_decap_8 FILLER_5_393 ();
 sg13g2_decap_8 FILLER_5_400 ();
 sg13g2_fill_2 FILLER_5_407 ();
 sg13g2_fill_1 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_52 ();
 sg13g2_fill_2 FILLER_6_64 ();
 sg13g2_fill_1 FILLER_6_80 ();
 sg13g2_decap_4 FILLER_6_86 ();
 sg13g2_fill_2 FILLER_6_98 ();
 sg13g2_decap_4 FILLER_6_104 ();
 sg13g2_decap_4 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_143 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_fill_2 FILLER_6_168 ();
 sg13g2_fill_1 FILLER_6_170 ();
 sg13g2_decap_4 FILLER_6_191 ();
 sg13g2_fill_1 FILLER_6_195 ();
 sg13g2_decap_8 FILLER_6_222 ();
 sg13g2_decap_8 FILLER_6_229 ();
 sg13g2_decap_8 FILLER_6_236 ();
 sg13g2_decap_8 FILLER_6_243 ();
 sg13g2_decap_8 FILLER_6_250 ();
 sg13g2_decap_8 FILLER_6_257 ();
 sg13g2_decap_8 FILLER_6_264 ();
 sg13g2_decap_8 FILLER_6_271 ();
 sg13g2_decap_8 FILLER_6_278 ();
 sg13g2_decap_8 FILLER_6_285 ();
 sg13g2_decap_8 FILLER_6_292 ();
 sg13g2_decap_8 FILLER_6_299 ();
 sg13g2_decap_8 FILLER_6_306 ();
 sg13g2_decap_8 FILLER_6_313 ();
 sg13g2_decap_8 FILLER_6_320 ();
 sg13g2_decap_8 FILLER_6_327 ();
 sg13g2_decap_8 FILLER_6_334 ();
 sg13g2_decap_8 FILLER_6_341 ();
 sg13g2_decap_8 FILLER_6_348 ();
 sg13g2_decap_8 FILLER_6_355 ();
 sg13g2_decap_8 FILLER_6_362 ();
 sg13g2_decap_8 FILLER_6_369 ();
 sg13g2_decap_8 FILLER_6_376 ();
 sg13g2_decap_8 FILLER_6_383 ();
 sg13g2_decap_8 FILLER_6_390 ();
 sg13g2_decap_8 FILLER_6_397 ();
 sg13g2_decap_4 FILLER_6_404 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_17 ();
 sg13g2_decap_4 FILLER_7_24 ();
 sg13g2_fill_2 FILLER_7_28 ();
 sg13g2_decap_4 FILLER_7_35 ();
 sg13g2_fill_2 FILLER_7_48 ();
 sg13g2_decap_8 FILLER_7_53 ();
 sg13g2_decap_8 FILLER_7_60 ();
 sg13g2_fill_2 FILLER_7_67 ();
 sg13g2_fill_1 FILLER_7_69 ();
 sg13g2_fill_2 FILLER_7_75 ();
 sg13g2_fill_1 FILLER_7_85 ();
 sg13g2_fill_2 FILLER_7_98 ();
 sg13g2_decap_4 FILLER_7_110 ();
 sg13g2_fill_1 FILLER_7_114 ();
 sg13g2_decap_4 FILLER_7_123 ();
 sg13g2_fill_1 FILLER_7_127 ();
 sg13g2_fill_2 FILLER_7_136 ();
 sg13g2_fill_1 FILLER_7_138 ();
 sg13g2_decap_8 FILLER_7_158 ();
 sg13g2_decap_8 FILLER_7_165 ();
 sg13g2_fill_2 FILLER_7_172 ();
 sg13g2_fill_1 FILLER_7_174 ();
 sg13g2_decap_8 FILLER_7_180 ();
 sg13g2_fill_2 FILLER_7_187 ();
 sg13g2_fill_2 FILLER_7_215 ();
 sg13g2_decap_8 FILLER_7_222 ();
 sg13g2_fill_2 FILLER_7_229 ();
 sg13g2_decap_8 FILLER_7_257 ();
 sg13g2_fill_1 FILLER_7_264 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_fill_1 FILLER_8_0 ();
 sg13g2_fill_2 FILLER_8_72 ();
 sg13g2_decap_8 FILLER_8_97 ();
 sg13g2_decap_8 FILLER_8_109 ();
 sg13g2_fill_2 FILLER_8_116 ();
 sg13g2_fill_1 FILLER_8_118 ();
 sg13g2_fill_2 FILLER_8_131 ();
 sg13g2_fill_1 FILLER_8_133 ();
 sg13g2_fill_2 FILLER_8_148 ();
 sg13g2_fill_1 FILLER_8_192 ();
 sg13g2_decap_4 FILLER_8_208 ();
 sg13g2_decap_4 FILLER_8_243 ();
 sg13g2_fill_2 FILLER_8_247 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_11 ();
 sg13g2_fill_2 FILLER_9_18 ();
 sg13g2_fill_1 FILLER_9_20 ();
 sg13g2_fill_2 FILLER_9_36 ();
 sg13g2_fill_1 FILLER_9_38 ();
 sg13g2_decap_8 FILLER_9_48 ();
 sg13g2_decap_8 FILLER_9_55 ();
 sg13g2_decap_4 FILLER_9_62 ();
 sg13g2_decap_8 FILLER_9_92 ();
 sg13g2_decap_4 FILLER_9_120 ();
 sg13g2_decap_4 FILLER_9_138 ();
 sg13g2_fill_2 FILLER_9_142 ();
 sg13g2_fill_2 FILLER_9_159 ();
 sg13g2_fill_1 FILLER_9_161 ();
 sg13g2_fill_2 FILLER_9_188 ();
 sg13g2_fill_1 FILLER_9_190 ();
 sg13g2_fill_1 FILLER_9_211 ();
 sg13g2_decap_8 FILLER_9_227 ();
 sg13g2_decap_8 FILLER_9_234 ();
 sg13g2_fill_1 FILLER_9_241 ();
 sg13g2_fill_1 FILLER_9_269 ();
 sg13g2_decap_8 FILLER_9_279 ();
 sg13g2_decap_8 FILLER_9_286 ();
 sg13g2_decap_8 FILLER_9_293 ();
 sg13g2_decap_8 FILLER_9_300 ();
 sg13g2_decap_8 FILLER_9_307 ();
 sg13g2_decap_8 FILLER_9_314 ();
 sg13g2_decap_8 FILLER_9_321 ();
 sg13g2_decap_8 FILLER_9_328 ();
 sg13g2_decap_8 FILLER_9_335 ();
 sg13g2_decap_8 FILLER_9_342 ();
 sg13g2_decap_8 FILLER_9_349 ();
 sg13g2_decap_8 FILLER_9_356 ();
 sg13g2_decap_8 FILLER_9_363 ();
 sg13g2_decap_8 FILLER_9_370 ();
 sg13g2_decap_8 FILLER_9_377 ();
 sg13g2_decap_8 FILLER_9_384 ();
 sg13g2_decap_8 FILLER_9_391 ();
 sg13g2_decap_8 FILLER_9_398 ();
 sg13g2_decap_4 FILLER_9_405 ();
 sg13g2_fill_1 FILLER_10_34 ();
 sg13g2_fill_2 FILLER_10_69 ();
 sg13g2_decap_8 FILLER_10_79 ();
 sg13g2_decap_4 FILLER_10_86 ();
 sg13g2_decap_4 FILLER_10_95 ();
 sg13g2_fill_1 FILLER_10_134 ();
 sg13g2_decap_8 FILLER_10_143 ();
 sg13g2_decap_8 FILLER_10_150 ();
 sg13g2_decap_8 FILLER_10_171 ();
 sg13g2_fill_1 FILLER_10_178 ();
 sg13g2_decap_8 FILLER_10_187 ();
 sg13g2_fill_1 FILLER_10_202 ();
 sg13g2_decap_4 FILLER_10_208 ();
 sg13g2_decap_4 FILLER_10_217 ();
 sg13g2_fill_2 FILLER_10_221 ();
 sg13g2_fill_2 FILLER_10_254 ();
 sg13g2_fill_2 FILLER_10_261 ();
 sg13g2_decap_8 FILLER_10_300 ();
 sg13g2_decap_8 FILLER_10_307 ();
 sg13g2_decap_8 FILLER_10_314 ();
 sg13g2_decap_8 FILLER_10_321 ();
 sg13g2_decap_8 FILLER_10_328 ();
 sg13g2_decap_8 FILLER_10_335 ();
 sg13g2_decap_8 FILLER_10_342 ();
 sg13g2_decap_8 FILLER_10_349 ();
 sg13g2_decap_8 FILLER_10_356 ();
 sg13g2_decap_8 FILLER_10_363 ();
 sg13g2_decap_8 FILLER_10_370 ();
 sg13g2_decap_8 FILLER_10_377 ();
 sg13g2_decap_8 FILLER_10_384 ();
 sg13g2_decap_8 FILLER_10_391 ();
 sg13g2_decap_8 FILLER_10_398 ();
 sg13g2_decap_4 FILLER_10_405 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_fill_1 FILLER_11_12 ();
 sg13g2_fill_2 FILLER_11_23 ();
 sg13g2_decap_8 FILLER_11_29 ();
 sg13g2_fill_1 FILLER_11_45 ();
 sg13g2_fill_2 FILLER_11_51 ();
 sg13g2_fill_1 FILLER_11_53 ();
 sg13g2_fill_2 FILLER_11_85 ();
 sg13g2_fill_1 FILLER_11_97 ();
 sg13g2_decap_8 FILLER_11_108 ();
 sg13g2_fill_2 FILLER_11_115 ();
 sg13g2_fill_1 FILLER_11_153 ();
 sg13g2_fill_2 FILLER_11_195 ();
 sg13g2_decap_8 FILLER_11_227 ();
 sg13g2_decap_8 FILLER_11_234 ();
 sg13g2_fill_1 FILLER_11_241 ();
 sg13g2_fill_2 FILLER_11_254 ();
 sg13g2_fill_1 FILLER_11_256 ();
 sg13g2_decap_8 FILLER_11_306 ();
 sg13g2_decap_8 FILLER_11_313 ();
 sg13g2_decap_8 FILLER_11_320 ();
 sg13g2_decap_8 FILLER_11_327 ();
 sg13g2_decap_8 FILLER_11_334 ();
 sg13g2_decap_8 FILLER_11_341 ();
 sg13g2_decap_8 FILLER_11_348 ();
 sg13g2_decap_8 FILLER_11_355 ();
 sg13g2_decap_8 FILLER_11_362 ();
 sg13g2_decap_8 FILLER_11_369 ();
 sg13g2_decap_8 FILLER_11_376 ();
 sg13g2_decap_8 FILLER_11_383 ();
 sg13g2_decap_8 FILLER_11_390 ();
 sg13g2_decap_8 FILLER_11_397 ();
 sg13g2_decap_4 FILLER_11_404 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_4 FILLER_12_31 ();
 sg13g2_fill_1 FILLER_12_35 ();
 sg13g2_fill_1 FILLER_12_41 ();
 sg13g2_fill_2 FILLER_12_59 ();
 sg13g2_decap_8 FILLER_12_66 ();
 sg13g2_decap_8 FILLER_12_73 ();
 sg13g2_decap_4 FILLER_12_80 ();
 sg13g2_fill_1 FILLER_12_84 ();
 sg13g2_decap_4 FILLER_12_93 ();
 sg13g2_decap_8 FILLER_12_149 ();
 sg13g2_decap_8 FILLER_12_156 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_4 FILLER_12_182 ();
 sg13g2_decap_4 FILLER_12_194 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_fill_2 FILLER_12_231 ();
 sg13g2_fill_1 FILLER_12_233 ();
 sg13g2_decap_4 FILLER_12_249 ();
 sg13g2_fill_1 FILLER_12_253 ();
 sg13g2_decap_8 FILLER_12_267 ();
 sg13g2_fill_1 FILLER_12_274 ();
 sg13g2_decap_8 FILLER_12_288 ();
 sg13g2_decap_8 FILLER_12_295 ();
 sg13g2_decap_8 FILLER_12_302 ();
 sg13g2_decap_8 FILLER_12_309 ();
 sg13g2_decap_8 FILLER_12_316 ();
 sg13g2_decap_8 FILLER_12_323 ();
 sg13g2_decap_8 FILLER_12_330 ();
 sg13g2_decap_8 FILLER_12_337 ();
 sg13g2_decap_8 FILLER_12_344 ();
 sg13g2_decap_8 FILLER_12_351 ();
 sg13g2_decap_8 FILLER_12_358 ();
 sg13g2_decap_8 FILLER_12_365 ();
 sg13g2_decap_8 FILLER_12_372 ();
 sg13g2_decap_8 FILLER_12_379 ();
 sg13g2_decap_8 FILLER_12_386 ();
 sg13g2_decap_8 FILLER_12_393 ();
 sg13g2_decap_8 FILLER_12_400 ();
 sg13g2_fill_2 FILLER_12_407 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_fill_1 FILLER_13_12 ();
 sg13g2_decap_8 FILLER_13_86 ();
 sg13g2_fill_1 FILLER_13_93 ();
 sg13g2_decap_4 FILLER_13_99 ();
 sg13g2_fill_1 FILLER_13_103 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_fill_2 FILLER_13_119 ();
 sg13g2_decap_4 FILLER_13_126 ();
 sg13g2_fill_1 FILLER_13_130 ();
 sg13g2_decap_8 FILLER_13_165 ();
 sg13g2_fill_2 FILLER_13_198 ();
 sg13g2_decap_8 FILLER_13_212 ();
 sg13g2_fill_2 FILLER_13_219 ();
 sg13g2_fill_2 FILLER_13_224 ();
 sg13g2_decap_4 FILLER_13_247 ();
 sg13g2_fill_2 FILLER_13_276 ();
 sg13g2_decap_8 FILLER_13_304 ();
 sg13g2_decap_8 FILLER_13_311 ();
 sg13g2_decap_8 FILLER_13_318 ();
 sg13g2_decap_8 FILLER_13_325 ();
 sg13g2_decap_8 FILLER_13_332 ();
 sg13g2_decap_8 FILLER_13_339 ();
 sg13g2_decap_8 FILLER_13_346 ();
 sg13g2_decap_8 FILLER_13_353 ();
 sg13g2_decap_8 FILLER_13_360 ();
 sg13g2_decap_8 FILLER_13_367 ();
 sg13g2_decap_8 FILLER_13_374 ();
 sg13g2_decap_8 FILLER_13_381 ();
 sg13g2_decap_8 FILLER_13_388 ();
 sg13g2_decap_8 FILLER_13_395 ();
 sg13g2_decap_8 FILLER_13_402 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_fill_2 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_4 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_30 ();
 sg13g2_decap_4 FILLER_14_42 ();
 sg13g2_fill_1 FILLER_14_52 ();
 sg13g2_fill_1 FILLER_14_58 ();
 sg13g2_fill_1 FILLER_14_69 ();
 sg13g2_decap_4 FILLER_14_122 ();
 sg13g2_fill_1 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_144 ();
 sg13g2_decap_4 FILLER_14_180 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_fill_1 FILLER_14_196 ();
 sg13g2_fill_2 FILLER_14_228 ();
 sg13g2_fill_1 FILLER_14_230 ();
 sg13g2_fill_1 FILLER_14_236 ();
 sg13g2_fill_2 FILLER_14_247 ();
 sg13g2_fill_1 FILLER_14_249 ();
 sg13g2_decap_8 FILLER_14_255 ();
 sg13g2_fill_1 FILLER_14_262 ();
 sg13g2_decap_4 FILLER_14_271 ();
 sg13g2_fill_2 FILLER_14_275 ();
 sg13g2_decap_8 FILLER_14_282 ();
 sg13g2_decap_8 FILLER_14_289 ();
 sg13g2_decap_8 FILLER_14_296 ();
 sg13g2_decap_8 FILLER_14_303 ();
 sg13g2_decap_8 FILLER_14_310 ();
 sg13g2_decap_8 FILLER_14_317 ();
 sg13g2_decap_8 FILLER_14_324 ();
 sg13g2_decap_8 FILLER_14_331 ();
 sg13g2_decap_8 FILLER_14_338 ();
 sg13g2_decap_8 FILLER_14_345 ();
 sg13g2_decap_8 FILLER_14_352 ();
 sg13g2_decap_8 FILLER_14_359 ();
 sg13g2_decap_8 FILLER_14_366 ();
 sg13g2_decap_8 FILLER_14_373 ();
 sg13g2_decap_8 FILLER_14_380 ();
 sg13g2_decap_8 FILLER_14_387 ();
 sg13g2_decap_8 FILLER_14_394 ();
 sg13g2_decap_8 FILLER_14_401 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_fill_2 FILLER_15_34 ();
 sg13g2_fill_2 FILLER_15_69 ();
 sg13g2_decap_8 FILLER_15_79 ();
 sg13g2_fill_1 FILLER_15_86 ();
 sg13g2_decap_8 FILLER_15_92 ();
 sg13g2_fill_2 FILLER_15_99 ();
 sg13g2_fill_1 FILLER_15_101 ();
 sg13g2_decap_8 FILLER_15_118 ();
 sg13g2_fill_2 FILLER_15_125 ();
 sg13g2_fill_2 FILLER_15_136 ();
 sg13g2_fill_2 FILLER_15_157 ();
 sg13g2_fill_2 FILLER_15_168 ();
 sg13g2_fill_1 FILLER_15_180 ();
 sg13g2_decap_4 FILLER_15_197 ();
 sg13g2_fill_2 FILLER_15_205 ();
 sg13g2_fill_1 FILLER_15_207 ();
 sg13g2_fill_2 FILLER_15_213 ();
 sg13g2_decap_8 FILLER_15_265 ();
 sg13g2_fill_2 FILLER_15_272 ();
 sg13g2_decap_8 FILLER_15_308 ();
 sg13g2_decap_8 FILLER_15_315 ();
 sg13g2_decap_8 FILLER_15_322 ();
 sg13g2_decap_8 FILLER_15_329 ();
 sg13g2_decap_8 FILLER_15_336 ();
 sg13g2_decap_8 FILLER_15_343 ();
 sg13g2_decap_8 FILLER_15_350 ();
 sg13g2_decap_8 FILLER_15_357 ();
 sg13g2_decap_8 FILLER_15_364 ();
 sg13g2_decap_8 FILLER_15_371 ();
 sg13g2_decap_8 FILLER_15_378 ();
 sg13g2_decap_8 FILLER_15_385 ();
 sg13g2_decap_8 FILLER_15_392 ();
 sg13g2_decap_8 FILLER_15_399 ();
 sg13g2_fill_2 FILLER_15_406 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_fill_2 FILLER_16_0 ();
 sg13g2_decap_4 FILLER_16_33 ();
 sg13g2_fill_1 FILLER_16_37 ();
 sg13g2_fill_2 FILLER_16_43 ();
 sg13g2_fill_1 FILLER_16_45 ();
 sg13g2_decap_8 FILLER_16_51 ();
 sg13g2_decap_4 FILLER_16_58 ();
 sg13g2_fill_1 FILLER_16_62 ();
 sg13g2_fill_2 FILLER_16_94 ();
 sg13g2_fill_2 FILLER_16_102 ();
 sg13g2_fill_1 FILLER_16_104 ();
 sg13g2_decap_8 FILLER_16_113 ();
 sg13g2_fill_2 FILLER_16_131 ();
 sg13g2_fill_1 FILLER_16_133 ();
 sg13g2_decap_4 FILLER_16_154 ();
 sg13g2_fill_1 FILLER_16_158 ();
 sg13g2_fill_1 FILLER_16_175 ();
 sg13g2_decap_4 FILLER_16_201 ();
 sg13g2_decap_8 FILLER_16_231 ();
 sg13g2_decap_4 FILLER_16_238 ();
 sg13g2_fill_2 FILLER_16_242 ();
 sg13g2_fill_1 FILLER_16_291 ();
 sg13g2_fill_2 FILLER_16_300 ();
 sg13g2_decap_4 FILLER_16_310 ();
 sg13g2_decap_8 FILLER_16_324 ();
 sg13g2_fill_2 FILLER_16_331 ();
 sg13g2_fill_1 FILLER_16_333 ();
 sg13g2_decap_8 FILLER_16_348 ();
 sg13g2_decap_4 FILLER_16_355 ();
 sg13g2_fill_1 FILLER_16_359 ();
 sg13g2_decap_8 FILLER_16_368 ();
 sg13g2_decap_8 FILLER_16_375 ();
 sg13g2_decap_8 FILLER_16_382 ();
 sg13g2_decap_8 FILLER_16_389 ();
 sg13g2_decap_8 FILLER_16_396 ();
 sg13g2_decap_4 FILLER_16_403 ();
 sg13g2_fill_2 FILLER_16_407 ();
 sg13g2_decap_4 FILLER_17_0 ();
 sg13g2_fill_1 FILLER_17_4 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_fill_2 FILLER_17_28 ();
 sg13g2_fill_1 FILLER_17_30 ();
 sg13g2_decap_4 FILLER_17_35 ();
 sg13g2_fill_2 FILLER_17_53 ();
 sg13g2_fill_1 FILLER_17_55 ();
 sg13g2_decap_4 FILLER_17_64 ();
 sg13g2_fill_2 FILLER_17_68 ();
 sg13g2_fill_2 FILLER_17_84 ();
 sg13g2_fill_1 FILLER_17_86 ();
 sg13g2_fill_2 FILLER_17_92 ();
 sg13g2_fill_2 FILLER_17_102 ();
 sg13g2_fill_1 FILLER_17_104 ();
 sg13g2_decap_4 FILLER_17_114 ();
 sg13g2_fill_2 FILLER_17_163 ();
 sg13g2_fill_2 FILLER_17_179 ();
 sg13g2_decap_8 FILLER_17_197 ();
 sg13g2_decap_4 FILLER_17_204 ();
 sg13g2_fill_2 FILLER_17_208 ();
 sg13g2_decap_4 FILLER_17_214 ();
 sg13g2_fill_2 FILLER_17_218 ();
 sg13g2_decap_4 FILLER_17_228 ();
 sg13g2_fill_2 FILLER_17_232 ();
 sg13g2_decap_8 FILLER_17_250 ();
 sg13g2_fill_2 FILLER_17_257 ();
 sg13g2_fill_2 FILLER_17_263 ();
 sg13g2_fill_1 FILLER_17_265 ();
 sg13g2_fill_2 FILLER_17_270 ();
 sg13g2_decap_4 FILLER_17_282 ();
 sg13g2_decap_8 FILLER_17_291 ();
 sg13g2_fill_2 FILLER_17_298 ();
 sg13g2_decap_4 FILLER_17_319 ();
 sg13g2_decap_4 FILLER_17_329 ();
 sg13g2_fill_2 FILLER_17_355 ();
 sg13g2_fill_1 FILLER_17_357 ();
 sg13g2_decap_8 FILLER_17_392 ();
 sg13g2_decap_8 FILLER_17_399 ();
 sg13g2_fill_2 FILLER_17_406 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_fill_2 FILLER_18_0 ();
 sg13g2_decap_4 FILLER_18_33 ();
 sg13g2_decap_8 FILLER_18_54 ();
 sg13g2_decap_4 FILLER_18_61 ();
 sg13g2_fill_1 FILLER_18_65 ();
 sg13g2_fill_2 FILLER_18_86 ();
 sg13g2_fill_1 FILLER_18_88 ();
 sg13g2_decap_8 FILLER_18_94 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_4 FILLER_18_140 ();
 sg13g2_decap_8 FILLER_18_158 ();
 sg13g2_fill_1 FILLER_18_165 ();
 sg13g2_decap_4 FILLER_18_200 ();
 sg13g2_fill_1 FILLER_18_230 ();
 sg13g2_decap_4 FILLER_18_247 ();
 sg13g2_fill_2 FILLER_18_251 ();
 sg13g2_fill_1 FILLER_18_289 ();
 sg13g2_fill_2 FILLER_18_313 ();
 sg13g2_decap_4 FILLER_18_333 ();
 sg13g2_fill_1 FILLER_18_337 ();
 sg13g2_fill_2 FILLER_18_350 ();
 sg13g2_fill_1 FILLER_18_352 ();
 sg13g2_fill_1 FILLER_18_370 ();
 sg13g2_decap_8 FILLER_18_397 ();
 sg13g2_decap_4 FILLER_18_404 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_fill_2 FILLER_19_0 ();
 sg13g2_fill_1 FILLER_19_2 ();
 sg13g2_fill_2 FILLER_19_17 ();
 sg13g2_fill_1 FILLER_19_19 ();
 sg13g2_decap_4 FILLER_19_34 ();
 sg13g2_fill_2 FILLER_19_38 ();
 sg13g2_decap_8 FILLER_19_80 ();
 sg13g2_decap_4 FILLER_19_87 ();
 sg13g2_fill_1 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_136 ();
 sg13g2_fill_1 FILLER_19_143 ();
 sg13g2_decap_8 FILLER_19_152 ();
 sg13g2_decap_8 FILLER_19_159 ();
 sg13g2_decap_4 FILLER_19_166 ();
 sg13g2_decap_4 FILLER_19_175 ();
 sg13g2_fill_2 FILLER_19_179 ();
 sg13g2_fill_1 FILLER_19_189 ();
 sg13g2_decap_4 FILLER_19_195 ();
 sg13g2_fill_1 FILLER_19_199 ();
 sg13g2_decap_8 FILLER_19_213 ();
 sg13g2_decap_8 FILLER_19_220 ();
 sg13g2_decap_8 FILLER_19_227 ();
 sg13g2_fill_2 FILLER_19_234 ();
 sg13g2_decap_4 FILLER_19_241 ();
 sg13g2_fill_1 FILLER_19_245 ();
 sg13g2_fill_2 FILLER_19_256 ();
 sg13g2_fill_1 FILLER_19_258 ();
 sg13g2_fill_1 FILLER_19_273 ();
 sg13g2_fill_1 FILLER_19_278 ();
 sg13g2_decap_8 FILLER_19_292 ();
 sg13g2_decap_8 FILLER_19_320 ();
 sg13g2_fill_1 FILLER_19_327 ();
 sg13g2_fill_2 FILLER_19_350 ();
 sg13g2_fill_1 FILLER_19_352 ();
 sg13g2_fill_2 FILLER_19_361 ();
 sg13g2_decap_8 FILLER_19_371 ();
 sg13g2_fill_2 FILLER_19_378 ();
 sg13g2_fill_1 FILLER_19_380 ();
 sg13g2_fill_2 FILLER_19_407 ();
 sg13g2_decap_4 FILLER_20_0 ();
 sg13g2_decap_4 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_4 FILLER_20_63 ();
 sg13g2_fill_1 FILLER_20_67 ();
 sg13g2_decap_4 FILLER_20_78 ();
 sg13g2_fill_2 FILLER_20_82 ();
 sg13g2_fill_2 FILLER_20_109 ();
 sg13g2_fill_2 FILLER_20_123 ();
 sg13g2_fill_1 FILLER_20_125 ();
 sg13g2_fill_2 FILLER_20_139 ();
 sg13g2_fill_1 FILLER_20_141 ();
 sg13g2_fill_2 FILLER_20_168 ();
 sg13g2_fill_1 FILLER_20_170 ();
 sg13g2_decap_8 FILLER_20_197 ();
 sg13g2_fill_2 FILLER_20_204 ();
 sg13g2_decap_4 FILLER_20_214 ();
 sg13g2_decap_4 FILLER_20_231 ();
 sg13g2_fill_2 FILLER_20_235 ();
 sg13g2_decap_8 FILLER_20_246 ();
 sg13g2_fill_1 FILLER_20_253 ();
 sg13g2_fill_2 FILLER_20_266 ();
 sg13g2_fill_2 FILLER_20_301 ();
 sg13g2_fill_1 FILLER_20_303 ();
 sg13g2_decap_8 FILLER_20_322 ();
 sg13g2_fill_1 FILLER_20_329 ();
 sg13g2_decap_8 FILLER_20_346 ();
 sg13g2_decap_4 FILLER_20_353 ();
 sg13g2_fill_1 FILLER_20_372 ();
 sg13g2_fill_1 FILLER_20_378 ();
 sg13g2_decap_4 FILLER_20_405 ();
 sg13g2_fill_2 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_4 FILLER_21_35 ();
 sg13g2_fill_1 FILLER_21_39 ();
 sg13g2_decap_8 FILLER_21_45 ();
 sg13g2_fill_2 FILLER_21_88 ();
 sg13g2_decap_8 FILLER_21_106 ();
 sg13g2_decap_4 FILLER_21_167 ();
 sg13g2_fill_1 FILLER_21_212 ();
 sg13g2_fill_1 FILLER_21_253 ();
 sg13g2_fill_2 FILLER_21_275 ();
 sg13g2_fill_1 FILLER_21_277 ();
 sg13g2_decap_4 FILLER_21_316 ();
 sg13g2_decap_4 FILLER_21_328 ();
 sg13g2_decap_8 FILLER_21_345 ();
 sg13g2_fill_2 FILLER_21_352 ();
 sg13g2_fill_2 FILLER_21_377 ();
 sg13g2_decap_8 FILLER_21_387 ();
 sg13g2_decap_8 FILLER_21_394 ();
 sg13g2_decap_8 FILLER_21_401 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_decap_4 FILLER_22_0 ();
 sg13g2_fill_1 FILLER_22_4 ();
 sg13g2_decap_8 FILLER_22_23 ();
 sg13g2_decap_4 FILLER_22_66 ();
 sg13g2_fill_2 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_82 ();
 sg13g2_fill_1 FILLER_22_89 ();
 sg13g2_decap_4 FILLER_22_102 ();
 sg13g2_fill_1 FILLER_22_106 ();
 sg13g2_decap_8 FILLER_22_137 ();
 sg13g2_fill_2 FILLER_22_149 ();
 sg13g2_fill_1 FILLER_22_151 ();
 sg13g2_decap_8 FILLER_22_157 ();
 sg13g2_decap_8 FILLER_22_187 ();
 sg13g2_fill_1 FILLER_22_194 ();
 sg13g2_decap_8 FILLER_22_208 ();
 sg13g2_decap_8 FILLER_22_215 ();
 sg13g2_decap_8 FILLER_22_222 ();
 sg13g2_fill_1 FILLER_22_229 ();
 sg13g2_decap_8 FILLER_22_248 ();
 sg13g2_decap_4 FILLER_22_255 ();
 sg13g2_fill_1 FILLER_22_259 ();
 sg13g2_decap_8 FILLER_22_264 ();
 sg13g2_decap_8 FILLER_22_271 ();
 sg13g2_decap_4 FILLER_22_278 ();
 sg13g2_fill_2 FILLER_22_282 ();
 sg13g2_decap_4 FILLER_22_289 ();
 sg13g2_fill_2 FILLER_22_293 ();
 sg13g2_decap_4 FILLER_22_309 ();
 sg13g2_fill_1 FILLER_22_313 ();
 sg13g2_decap_4 FILLER_22_322 ();
 sg13g2_fill_2 FILLER_22_335 ();
 sg13g2_fill_2 FILLER_22_345 ();
 sg13g2_fill_1 FILLER_22_347 ();
 sg13g2_fill_2 FILLER_22_380 ();
 sg13g2_fill_1 FILLER_22_382 ();
 sg13g2_decap_4 FILLER_23_0 ();
 sg13g2_fill_1 FILLER_23_4 ();
 sg13g2_fill_2 FILLER_23_31 ();
 sg13g2_fill_1 FILLER_23_33 ();
 sg13g2_fill_2 FILLER_23_53 ();
 sg13g2_fill_2 FILLER_23_82 ();
 sg13g2_fill_2 FILLER_23_111 ();
 sg13g2_fill_1 FILLER_23_113 ();
 sg13g2_fill_2 FILLER_23_123 ();
 sg13g2_fill_2 FILLER_23_167 ();
 sg13g2_decap_8 FILLER_23_205 ();
 sg13g2_decap_4 FILLER_23_212 ();
 sg13g2_fill_1 FILLER_23_216 ();
 sg13g2_decap_4 FILLER_23_299 ();
 sg13g2_decap_8 FILLER_23_327 ();
 sg13g2_fill_1 FILLER_23_350 ();
 sg13g2_fill_2 FILLER_23_386 ();
 sg13g2_decap_8 FILLER_23_397 ();
 sg13g2_decap_4 FILLER_23_404 ();
 sg13g2_fill_1 FILLER_23_408 ();
 sg13g2_fill_1 FILLER_24_0 ();
 sg13g2_fill_1 FILLER_24_13 ();
 sg13g2_fill_2 FILLER_24_33 ();
 sg13g2_fill_1 FILLER_24_40 ();
 sg13g2_fill_1 FILLER_24_62 ();
 sg13g2_decap_8 FILLER_24_67 ();
 sg13g2_decap_4 FILLER_24_74 ();
 sg13g2_fill_1 FILLER_24_78 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_fill_2 FILLER_24_91 ();
 sg13g2_fill_1 FILLER_24_93 ();
 sg13g2_decap_4 FILLER_24_115 ();
 sg13g2_decap_8 FILLER_24_139 ();
 sg13g2_decap_4 FILLER_24_151 ();
 sg13g2_fill_2 FILLER_24_155 ();
 sg13g2_decap_8 FILLER_24_165 ();
 sg13g2_fill_1 FILLER_24_172 ();
 sg13g2_fill_1 FILLER_24_178 ();
 sg13g2_fill_2 FILLER_24_196 ();
 sg13g2_fill_1 FILLER_24_198 ();
 sg13g2_decap_4 FILLER_24_204 ();
 sg13g2_decap_4 FILLER_24_212 ();
 sg13g2_fill_1 FILLER_24_216 ();
 sg13g2_fill_2 FILLER_24_243 ();
 sg13g2_fill_1 FILLER_24_245 ();
 sg13g2_decap_4 FILLER_24_270 ();
 sg13g2_fill_2 FILLER_24_283 ();
 sg13g2_fill_1 FILLER_24_285 ();
 sg13g2_fill_1 FILLER_24_330 ();
 sg13g2_fill_2 FILLER_24_355 ();
 sg13g2_fill_1 FILLER_24_357 ();
 sg13g2_decap_4 FILLER_24_366 ();
 sg13g2_decap_4 FILLER_24_374 ();
 sg13g2_fill_2 FILLER_24_378 ();
 sg13g2_fill_2 FILLER_24_406 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_fill_1 FILLER_25_0 ();
 sg13g2_decap_4 FILLER_25_13 ();
 sg13g2_fill_2 FILLER_25_41 ();
 sg13g2_fill_2 FILLER_25_85 ();
 sg13g2_fill_1 FILLER_25_87 ();
 sg13g2_fill_1 FILLER_25_96 ();
 sg13g2_decap_8 FILLER_25_109 ();
 sg13g2_fill_1 FILLER_25_116 ();
 sg13g2_fill_1 FILLER_25_137 ();
 sg13g2_fill_2 FILLER_25_190 ();
 sg13g2_fill_2 FILLER_25_223 ();
 sg13g2_fill_1 FILLER_25_225 ();
 sg13g2_fill_1 FILLER_25_240 ();
 sg13g2_fill_2 FILLER_25_250 ();
 sg13g2_fill_1 FILLER_25_252 ();
 sg13g2_fill_2 FILLER_25_263 ();
 sg13g2_fill_1 FILLER_25_291 ();
 sg13g2_decap_4 FILLER_25_299 ();
 sg13g2_decap_8 FILLER_25_311 ();
 sg13g2_fill_1 FILLER_25_318 ();
 sg13g2_decap_8 FILLER_25_342 ();
 sg13g2_decap_8 FILLER_25_349 ();
 sg13g2_fill_2 FILLER_25_376 ();
 sg13g2_decap_4 FILLER_26_26 ();
 sg13g2_fill_1 FILLER_26_66 ();
 sg13g2_decap_4 FILLER_26_88 ();
 sg13g2_fill_2 FILLER_26_92 ();
 sg13g2_decap_4 FILLER_26_110 ();
 sg13g2_fill_2 FILLER_26_114 ();
 sg13g2_decap_8 FILLER_26_138 ();
 sg13g2_decap_8 FILLER_26_145 ();
 sg13g2_decap_8 FILLER_26_152 ();
 sg13g2_decap_8 FILLER_26_159 ();
 sg13g2_fill_1 FILLER_26_166 ();
 sg13g2_fill_1 FILLER_26_171 ();
 sg13g2_fill_1 FILLER_26_180 ();
 sg13g2_fill_2 FILLER_26_199 ();
 sg13g2_decap_4 FILLER_26_213 ();
 sg13g2_decap_4 FILLER_26_223 ();
 sg13g2_fill_1 FILLER_26_263 ();
 sg13g2_fill_2 FILLER_26_271 ();
 sg13g2_fill_1 FILLER_26_273 ();
 sg13g2_fill_2 FILLER_26_283 ();
 sg13g2_fill_1 FILLER_26_285 ();
 sg13g2_fill_2 FILLER_26_321 ();
 sg13g2_fill_2 FILLER_26_366 ();
 sg13g2_fill_2 FILLER_26_392 ();
 sg13g2_decap_4 FILLER_26_403 ();
 sg13g2_fill_2 FILLER_26_407 ();
 sg13g2_fill_2 FILLER_27_0 ();
 sg13g2_fill_1 FILLER_27_2 ();
 sg13g2_fill_1 FILLER_27_20 ();
 sg13g2_fill_1 FILLER_27_39 ();
 sg13g2_fill_2 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_83 ();
 sg13g2_decap_8 FILLER_27_90 ();
 sg13g2_fill_2 FILLER_27_97 ();
 sg13g2_fill_1 FILLER_27_99 ();
 sg13g2_decap_4 FILLER_27_104 ();
 sg13g2_decap_8 FILLER_27_125 ();
 sg13g2_decap_4 FILLER_27_132 ();
 sg13g2_fill_1 FILLER_27_136 ();
 sg13g2_fill_2 FILLER_27_163 ();
 sg13g2_fill_2 FILLER_27_173 ();
 sg13g2_fill_1 FILLER_27_233 ();
 sg13g2_decap_4 FILLER_27_254 ();
 sg13g2_fill_2 FILLER_27_263 ();
 sg13g2_decap_4 FILLER_27_284 ();
 sg13g2_decap_8 FILLER_27_296 ();
 sg13g2_fill_1 FILLER_27_303 ();
 sg13g2_fill_2 FILLER_27_308 ();
 sg13g2_fill_1 FILLER_27_310 ();
 sg13g2_decap_8 FILLER_27_319 ();
 sg13g2_fill_1 FILLER_27_326 ();
 sg13g2_fill_1 FILLER_27_333 ();
 sg13g2_decap_8 FILLER_27_342 ();
 sg13g2_fill_2 FILLER_27_349 ();
 sg13g2_fill_2 FILLER_27_357 ();
 sg13g2_fill_1 FILLER_27_359 ();
 sg13g2_fill_2 FILLER_27_366 ();
 sg13g2_fill_2 FILLER_27_379 ();
 sg13g2_decap_8 FILLER_27_400 ();
 sg13g2_fill_2 FILLER_27_407 ();
 sg13g2_fill_2 FILLER_28_26 ();
 sg13g2_fill_1 FILLER_28_28 ();
 sg13g2_decap_4 FILLER_28_107 ();
 sg13g2_fill_2 FILLER_28_137 ();
 sg13g2_fill_1 FILLER_28_144 ();
 sg13g2_fill_2 FILLER_28_190 ();
 sg13g2_fill_2 FILLER_28_211 ();
 sg13g2_fill_1 FILLER_28_222 ();
 sg13g2_decap_8 FILLER_28_233 ();
 sg13g2_decap_8 FILLER_28_248 ();
 sg13g2_fill_1 FILLER_28_255 ();
 sg13g2_fill_2 FILLER_28_264 ();
 sg13g2_fill_2 FILLER_28_318 ();
 sg13g2_fill_1 FILLER_28_320 ();
 sg13g2_fill_2 FILLER_28_337 ();
 sg13g2_fill_1 FILLER_28_366 ();
 sg13g2_fill_2 FILLER_29_0 ();
 sg13g2_fill_1 FILLER_29_2 ();
 sg13g2_fill_1 FILLER_29_43 ();
 sg13g2_fill_2 FILLER_29_134 ();
 sg13g2_fill_2 FILLER_29_171 ();
 sg13g2_fill_1 FILLER_29_173 ();
 sg13g2_fill_1 FILLER_29_195 ();
 sg13g2_fill_1 FILLER_29_210 ();
 sg13g2_decap_4 FILLER_29_223 ();
 sg13g2_decap_8 FILLER_29_234 ();
 sg13g2_fill_1 FILLER_29_241 ();
 sg13g2_decap_8 FILLER_29_273 ();
 sg13g2_fill_2 FILLER_29_280 ();
 sg13g2_decap_4 FILLER_29_296 ();
 sg13g2_fill_2 FILLER_29_300 ();
 sg13g2_fill_1 FILLER_29_308 ();
 sg13g2_decap_8 FILLER_29_313 ();
 sg13g2_fill_2 FILLER_29_320 ();
 sg13g2_decap_8 FILLER_29_334 ();
 sg13g2_fill_2 FILLER_29_345 ();
 sg13g2_fill_2 FILLER_29_356 ();
 sg13g2_fill_1 FILLER_29_358 ();
 sg13g2_fill_2 FILLER_29_367 ();
 sg13g2_fill_1 FILLER_29_369 ();
 sg13g2_fill_2 FILLER_29_375 ();
 sg13g2_fill_1 FILLER_29_377 ();
 sg13g2_fill_1 FILLER_29_408 ();
 sg13g2_decap_4 FILLER_30_26 ();
 sg13g2_fill_2 FILLER_30_47 ();
 sg13g2_fill_1 FILLER_30_110 ();
 sg13g2_fill_2 FILLER_30_129 ();
 sg13g2_fill_1 FILLER_30_131 ();
 sg13g2_fill_1 FILLER_30_136 ();
 sg13g2_fill_2 FILLER_30_153 ();
 sg13g2_fill_2 FILLER_30_194 ();
 sg13g2_fill_2 FILLER_30_212 ();
 sg13g2_fill_1 FILLER_30_214 ();
 sg13g2_decap_4 FILLER_30_226 ();
 sg13g2_fill_2 FILLER_30_263 ();
 sg13g2_fill_1 FILLER_30_265 ();
 sg13g2_decap_4 FILLER_30_275 ();
 sg13g2_fill_1 FILLER_30_279 ();
 sg13g2_fill_2 FILLER_30_288 ();
 sg13g2_fill_1 FILLER_30_290 ();
 sg13g2_fill_2 FILLER_30_315 ();
 sg13g2_fill_2 FILLER_30_335 ();
 sg13g2_decap_4 FILLER_30_355 ();
 sg13g2_fill_1 FILLER_30_359 ();
 sg13g2_fill_2 FILLER_30_380 ();
 sg13g2_fill_1 FILLER_30_382 ();
 sg13g2_fill_2 FILLER_31_0 ();
 sg13g2_decap_4 FILLER_31_28 ();
 sg13g2_fill_1 FILLER_31_32 ();
 sg13g2_fill_2 FILLER_31_64 ();
 sg13g2_decap_8 FILLER_31_92 ();
 sg13g2_fill_1 FILLER_31_122 ();
 sg13g2_fill_1 FILLER_31_128 ();
 sg13g2_fill_2 FILLER_31_136 ();
 sg13g2_fill_1 FILLER_31_138 ();
 sg13g2_fill_2 FILLER_31_152 ();
 sg13g2_fill_2 FILLER_31_169 ();
 sg13g2_fill_2 FILLER_31_183 ();
 sg13g2_fill_1 FILLER_31_185 ();
 sg13g2_decap_4 FILLER_31_195 ();
 sg13g2_decap_4 FILLER_31_207 ();
 sg13g2_fill_2 FILLER_31_211 ();
 sg13g2_decap_4 FILLER_31_245 ();
 sg13g2_fill_1 FILLER_31_249 ();
 sg13g2_decap_8 FILLER_31_254 ();
 sg13g2_decap_4 FILLER_31_261 ();
 sg13g2_fill_1 FILLER_31_265 ();
 sg13g2_decap_8 FILLER_31_286 ();
 sg13g2_fill_2 FILLER_31_293 ();
 sg13g2_decap_8 FILLER_31_303 ();
 sg13g2_decap_8 FILLER_31_310 ();
 sg13g2_fill_2 FILLER_31_334 ();
 sg13g2_fill_1 FILLER_31_336 ();
 sg13g2_fill_1 FILLER_31_342 ();
 sg13g2_fill_1 FILLER_31_352 ();
 sg13g2_fill_2 FILLER_31_359 ();
 sg13g2_fill_2 FILLER_31_406 ();
 sg13g2_fill_1 FILLER_31_408 ();
 sg13g2_fill_2 FILLER_32_0 ();
 sg13g2_fill_2 FILLER_32_11 ();
 sg13g2_fill_1 FILLER_32_13 ();
 sg13g2_fill_2 FILLER_32_48 ();
 sg13g2_fill_1 FILLER_32_50 ();
 sg13g2_decap_4 FILLER_32_70 ();
 sg13g2_fill_1 FILLER_32_74 ();
 sg13g2_fill_1 FILLER_32_126 ();
 sg13g2_fill_2 FILLER_32_169 ();
 sg13g2_fill_1 FILLER_32_180 ();
 sg13g2_fill_2 FILLER_32_193 ();
 sg13g2_fill_1 FILLER_32_195 ();
 sg13g2_fill_1 FILLER_32_224 ();
 sg13g2_fill_1 FILLER_32_229 ();
 sg13g2_fill_2 FILLER_32_246 ();
 sg13g2_fill_1 FILLER_32_248 ();
 sg13g2_decap_4 FILLER_32_287 ();
 sg13g2_decap_4 FILLER_32_310 ();
 sg13g2_fill_2 FILLER_32_314 ();
 sg13g2_decap_4 FILLER_32_329 ();
 sg13g2_fill_1 FILLER_32_333 ();
 sg13g2_decap_8 FILLER_32_356 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_4 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_34 ();
 sg13g2_decap_4 FILLER_33_50 ();
 sg13g2_decap_4 FILLER_33_59 ();
 sg13g2_fill_2 FILLER_33_103 ();
 sg13g2_fill_2 FILLER_33_127 ();
 sg13g2_fill_2 FILLER_33_137 ();
 sg13g2_fill_1 FILLER_33_162 ();
 sg13g2_decap_8 FILLER_33_167 ();
 sg13g2_decap_4 FILLER_33_174 ();
 sg13g2_fill_1 FILLER_33_178 ();
 sg13g2_fill_2 FILLER_33_235 ();
 sg13g2_fill_1 FILLER_33_237 ();
 sg13g2_decap_8 FILLER_33_255 ();
 sg13g2_fill_2 FILLER_33_262 ();
 sg13g2_fill_2 FILLER_33_273 ();
 sg13g2_fill_1 FILLER_33_275 ();
 sg13g2_decap_4 FILLER_33_286 ();
 sg13g2_fill_1 FILLER_33_290 ();
 sg13g2_decap_4 FILLER_33_313 ();
 sg13g2_fill_2 FILLER_33_330 ();
 sg13g2_fill_1 FILLER_33_348 ();
 sg13g2_fill_2 FILLER_33_369 ();
 sg13g2_fill_2 FILLER_33_395 ();
 sg13g2_fill_1 FILLER_33_397 ();
 sg13g2_fill_2 FILLER_33_407 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_fill_1 FILLER_34_97 ();
 sg13g2_fill_2 FILLER_34_105 ();
 sg13g2_decap_8 FILLER_34_127 ();
 sg13g2_decap_8 FILLER_34_134 ();
 sg13g2_decap_4 FILLER_34_141 ();
 sg13g2_fill_1 FILLER_34_156 ();
 sg13g2_decap_4 FILLER_34_162 ();
 sg13g2_fill_1 FILLER_34_166 ();
 sg13g2_decap_4 FILLER_34_172 ();
 sg13g2_fill_1 FILLER_34_176 ();
 sg13g2_decap_8 FILLER_34_182 ();
 sg13g2_decap_4 FILLER_34_189 ();
 sg13g2_fill_2 FILLER_34_208 ();
 sg13g2_fill_1 FILLER_34_240 ();
 sg13g2_decap_4 FILLER_34_248 ();
 sg13g2_fill_1 FILLER_34_252 ();
 sg13g2_fill_2 FILLER_34_276 ();
 sg13g2_fill_1 FILLER_34_291 ();
 sg13g2_decap_4 FILLER_34_300 ();
 sg13g2_fill_1 FILLER_34_304 ();
 sg13g2_fill_2 FILLER_34_314 ();
 sg13g2_fill_1 FILLER_34_316 ();
 sg13g2_fill_2 FILLER_34_329 ();
 sg13g2_fill_1 FILLER_34_364 ();
 sg13g2_fill_1 FILLER_34_377 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_fill_1 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_71 ();
 sg13g2_decap_4 FILLER_35_78 ();
 sg13g2_fill_2 FILLER_35_82 ();
 sg13g2_decap_8 FILLER_35_94 ();
 sg13g2_decap_8 FILLER_35_101 ();
 sg13g2_fill_2 FILLER_35_108 ();
 sg13g2_fill_1 FILLER_35_110 ();
 sg13g2_decap_4 FILLER_35_120 ();
 sg13g2_fill_1 FILLER_35_124 ();
 sg13g2_fill_2 FILLER_35_134 ();
 sg13g2_decap_8 FILLER_35_155 ();
 sg13g2_fill_1 FILLER_35_172 ();
 sg13g2_decap_8 FILLER_35_188 ();
 sg13g2_fill_2 FILLER_35_195 ();
 sg13g2_fill_2 FILLER_35_204 ();
 sg13g2_decap_8 FILLER_35_211 ();
 sg13g2_decap_8 FILLER_35_218 ();
 sg13g2_decap_4 FILLER_35_225 ();
 sg13g2_fill_1 FILLER_35_229 ();
 sg13g2_fill_2 FILLER_35_267 ();
 sg13g2_decap_8 FILLER_35_285 ();
 sg13g2_fill_1 FILLER_35_292 ();
 sg13g2_decap_4 FILLER_35_317 ();
 sg13g2_fill_2 FILLER_35_392 ();
 sg13g2_decap_8 FILLER_35_398 ();
 sg13g2_decap_4 FILLER_35_405 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_4 FILLER_36_28 ();
 sg13g2_fill_1 FILLER_36_32 ();
 sg13g2_fill_2 FILLER_36_59 ();
 sg13g2_fill_2 FILLER_36_77 ();
 sg13g2_fill_1 FILLER_36_79 ();
 sg13g2_fill_2 FILLER_36_85 ();
 sg13g2_fill_2 FILLER_36_91 ();
 sg13g2_decap_4 FILLER_36_139 ();
 sg13g2_fill_2 FILLER_36_143 ();
 sg13g2_fill_1 FILLER_36_180 ();
 sg13g2_fill_2 FILLER_36_192 ();
 sg13g2_decap_8 FILLER_36_215 ();
 sg13g2_fill_2 FILLER_36_222 ();
 sg13g2_decap_8 FILLER_36_236 ();
 sg13g2_decap_4 FILLER_36_243 ();
 sg13g2_decap_8 FILLER_36_258 ();
 sg13g2_fill_2 FILLER_36_265 ();
 sg13g2_fill_2 FILLER_36_299 ();
 sg13g2_fill_1 FILLER_36_301 ();
 sg13g2_decap_8 FILLER_36_317 ();
 sg13g2_decap_8 FILLER_36_324 ();
 sg13g2_fill_2 FILLER_36_331 ();
 sg13g2_fill_1 FILLER_36_333 ();
 sg13g2_fill_2 FILLER_36_338 ();
 sg13g2_fill_2 FILLER_36_357 ();
 sg13g2_fill_2 FILLER_36_381 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_fill_1 FILLER_37_35 ();
 sg13g2_fill_1 FILLER_37_67 ();
 sg13g2_fill_1 FILLER_37_94 ();
 sg13g2_fill_2 FILLER_37_116 ();
 sg13g2_decap_4 FILLER_37_124 ();
 sg13g2_fill_1 FILLER_37_128 ();
 sg13g2_fill_2 FILLER_37_135 ();
 sg13g2_fill_1 FILLER_37_159 ();
 sg13g2_fill_2 FILLER_37_187 ();
 sg13g2_fill_1 FILLER_37_197 ();
 sg13g2_fill_2 FILLER_37_203 ();
 sg13g2_decap_8 FILLER_37_209 ();
 sg13g2_fill_2 FILLER_37_216 ();
 sg13g2_fill_1 FILLER_37_218 ();
 sg13g2_fill_2 FILLER_37_231 ();
 sg13g2_fill_1 FILLER_37_233 ();
 sg13g2_fill_2 FILLER_37_268 ();
 sg13g2_fill_2 FILLER_37_284 ();
 sg13g2_fill_1 FILLER_37_286 ();
 sg13g2_fill_2 FILLER_37_313 ();
 sg13g2_fill_2 FILLER_37_353 ();
 sg13g2_fill_2 FILLER_37_391 ();
 sg13g2_fill_1 FILLER_37_393 ();
 sg13g2_decap_8 FILLER_37_398 ();
 sg13g2_decap_4 FILLER_37_405 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_fill_2 FILLER_38_42 ();
 sg13g2_fill_1 FILLER_38_44 ();
 sg13g2_fill_1 FILLER_38_84 ();
 sg13g2_fill_2 FILLER_38_93 ();
 sg13g2_fill_1 FILLER_38_95 ();
 sg13g2_decap_4 FILLER_38_130 ();
 sg13g2_fill_2 FILLER_38_134 ();
 sg13g2_fill_2 FILLER_38_152 ();
 sg13g2_fill_2 FILLER_38_158 ();
 sg13g2_fill_2 FILLER_38_177 ();
 sg13g2_decap_4 FILLER_38_188 ();
 sg13g2_fill_2 FILLER_38_192 ();
 sg13g2_fill_2 FILLER_38_220 ();
 sg13g2_fill_1 FILLER_38_222 ();
 sg13g2_decap_8 FILLER_38_238 ();
 sg13g2_decap_8 FILLER_38_257 ();
 sg13g2_fill_2 FILLER_38_264 ();
 sg13g2_fill_1 FILLER_38_266 ();
 sg13g2_decap_4 FILLER_38_287 ();
 sg13g2_fill_2 FILLER_38_291 ();
 sg13g2_fill_2 FILLER_38_297 ();
 sg13g2_fill_1 FILLER_38_299 ();
 sg13g2_decap_8 FILLER_38_314 ();
 sg13g2_decap_4 FILLER_38_321 ();
 sg13g2_fill_1 FILLER_38_325 ();
 sg13g2_decap_8 FILLER_38_391 ();
 sg13g2_decap_8 FILLER_38_398 ();
 sg13g2_decap_4 FILLER_38_405 ();
 assign uio_oe[0] = net1;
 assign uio_oe[1] = net2;
 assign uio_oe[2] = net3;
 assign uio_oe[3] = net4;
 assign uio_oe[4] = net31;
 assign uio_oe[5] = net32;
 assign uio_oe[6] = net33;
 assign uio_oe[7] = net34;
 assign uio_out[0] = net5;
 assign uio_out[1] = net6;
 assign uio_out[2] = net7;
 assign uio_out[3] = net8;
endmodule

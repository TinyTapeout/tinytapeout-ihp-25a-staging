module tt_um_emilian_muxpga (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire clknet_0_clk;
 wire \cell_cfg[0][0] ;
 wire \cell_cfg[0][1] ;
 wire \cell_cfg[0][2] ;
 wire \cell_cfg[0][3] ;
 wire \cell_cfg[10][0] ;
 wire \cell_cfg[10][1] ;
 wire \cell_cfg[10][2] ;
 wire \cell_cfg[10][3] ;
 wire \cell_cfg[11][0] ;
 wire \cell_cfg[11][1] ;
 wire \cell_cfg[11][2] ;
 wire \cell_cfg[11][3] ;
 wire \cell_cfg[12][0] ;
 wire \cell_cfg[12][1] ;
 wire \cell_cfg[12][2] ;
 wire \cell_cfg[12][3] ;
 wire \cell_cfg[13][0] ;
 wire \cell_cfg[13][1] ;
 wire \cell_cfg[13][2] ;
 wire \cell_cfg[13][3] ;
 wire \cell_cfg[14][0] ;
 wire \cell_cfg[14][1] ;
 wire \cell_cfg[14][2] ;
 wire \cell_cfg[14][3] ;
 wire \cell_cfg[15][0] ;
 wire \cell_cfg[15][1] ;
 wire \cell_cfg[15][2] ;
 wire \cell_cfg[15][3] ;
 wire \cell_cfg[16][0] ;
 wire \cell_cfg[16][1] ;
 wire \cell_cfg[16][2] ;
 wire \cell_cfg[16][3] ;
 wire \cell_cfg[17][0] ;
 wire \cell_cfg[17][1] ;
 wire \cell_cfg[17][2] ;
 wire \cell_cfg[17][3] ;
 wire \cell_cfg[18][0] ;
 wire \cell_cfg[18][1] ;
 wire \cell_cfg[18][2] ;
 wire \cell_cfg[18][3] ;
 wire \cell_cfg[19][0] ;
 wire \cell_cfg[19][1] ;
 wire \cell_cfg[19][2] ;
 wire \cell_cfg[19][3] ;
 wire \cell_cfg[1][0] ;
 wire \cell_cfg[1][1] ;
 wire \cell_cfg[1][2] ;
 wire \cell_cfg[1][3] ;
 wire \cell_cfg[20][0] ;
 wire \cell_cfg[20][1] ;
 wire \cell_cfg[20][2] ;
 wire \cell_cfg[20][3] ;
 wire \cell_cfg[21][0] ;
 wire \cell_cfg[21][1] ;
 wire \cell_cfg[21][2] ;
 wire \cell_cfg[21][3] ;
 wire \cell_cfg[22][0] ;
 wire \cell_cfg[22][1] ;
 wire \cell_cfg[22][2] ;
 wire \cell_cfg[22][3] ;
 wire \cell_cfg[23][0] ;
 wire \cell_cfg[23][1] ;
 wire \cell_cfg[23][2] ;
 wire \cell_cfg[23][3] ;
 wire \cell_cfg[24][0] ;
 wire \cell_cfg[24][1] ;
 wire \cell_cfg[24][2] ;
 wire \cell_cfg[24][3] ;
 wire \cell_cfg[25][0] ;
 wire \cell_cfg[25][1] ;
 wire \cell_cfg[25][2] ;
 wire \cell_cfg[25][3] ;
 wire \cell_cfg[26][0] ;
 wire \cell_cfg[26][1] ;
 wire \cell_cfg[26][2] ;
 wire \cell_cfg[26][3] ;
 wire \cell_cfg[27][0] ;
 wire \cell_cfg[27][1] ;
 wire \cell_cfg[27][2] ;
 wire \cell_cfg[27][3] ;
 wire \cell_cfg[28][0] ;
 wire \cell_cfg[28][1] ;
 wire \cell_cfg[28][2] ;
 wire \cell_cfg[28][3] ;
 wire \cell_cfg[29][0] ;
 wire \cell_cfg[29][1] ;
 wire \cell_cfg[29][2] ;
 wire \cell_cfg[29][3] ;
 wire \cell_cfg[2][0] ;
 wire \cell_cfg[2][1] ;
 wire \cell_cfg[2][2] ;
 wire \cell_cfg[2][3] ;
 wire \cell_cfg[30][0] ;
 wire \cell_cfg[30][1] ;
 wire \cell_cfg[30][2] ;
 wire \cell_cfg[30][3] ;
 wire \cell_cfg[31][0] ;
 wire \cell_cfg[31][1] ;
 wire \cell_cfg[31][2] ;
 wire \cell_cfg[31][3] ;
 wire \cell_cfg[32][0] ;
 wire \cell_cfg[32][1] ;
 wire \cell_cfg[32][2] ;
 wire \cell_cfg[32][3] ;
 wire \cell_cfg[33][0] ;
 wire \cell_cfg[33][1] ;
 wire \cell_cfg[33][2] ;
 wire \cell_cfg[33][3] ;
 wire \cell_cfg[34][0] ;
 wire \cell_cfg[34][1] ;
 wire \cell_cfg[34][2] ;
 wire \cell_cfg[34][3] ;
 wire \cell_cfg[35][0] ;
 wire \cell_cfg[35][1] ;
 wire \cell_cfg[35][2] ;
 wire \cell_cfg[35][3] ;
 wire \cell_cfg[3][0] ;
 wire \cell_cfg[3][1] ;
 wire \cell_cfg[3][2] ;
 wire \cell_cfg[3][3] ;
 wire \cell_cfg[4][0] ;
 wire \cell_cfg[4][1] ;
 wire \cell_cfg[4][2] ;
 wire \cell_cfg[4][3] ;
 wire \cell_cfg[5][0] ;
 wire \cell_cfg[5][1] ;
 wire \cell_cfg[5][2] ;
 wire \cell_cfg[5][3] ;
 wire \cell_cfg[6][0] ;
 wire \cell_cfg[6][1] ;
 wire \cell_cfg[6][2] ;
 wire \cell_cfg[6][3] ;
 wire \cell_cfg[7][0] ;
 wire \cell_cfg[7][1] ;
 wire \cell_cfg[7][2] ;
 wire \cell_cfg[7][3] ;
 wire \cell_cfg[8][0] ;
 wire \cell_cfg[8][1] ;
 wire \cell_cfg[8][2] ;
 wire \cell_cfg[8][3] ;
 wire \cell_cfg[9][0] ;
 wire \cell_cfg[9][1] ;
 wire \cell_cfg[9][2] ;
 wire \cell_cfg[9][3] ;
 wire en_cells;
 wire \genrow[1].gencol[0].genblk1.c.bufs[0].A ;
 wire \genrow[1].gencol[1].genblk1.c.bufs[0].A ;
 wire \genrow[1].gencol[2].genblk1.c.bufs[0].A ;
 wire \genrow[1].gencol[3].genblk1.c.bufs[0].A ;
 wire \genrow[1].gencol[4].genblk1.c.bufs[0].A ;
 wire \genrow[2].gencol[0].genblk1.c.bufs[0].A ;
 wire \genrow[2].gencol[1].genblk1.c.bufs[0].A ;
 wire \genrow[2].gencol[2].genblk1.c.bufs[0].A ;
 wire \genrow[2].gencol[3].genblk1.c.bufs[0].A ;
 wire \genrow[2].gencol[4].genblk1.c.bufs[0].A ;
 wire \genrow[2].gencol[5].genblk1.c.bufs[0].A ;
 wire \genrow[3].gencol[0].genblk1.c.bufs[0].A ;
 wire \genrow[3].gencol[1].genblk1.c.bufs[0].A ;
 wire \genrow[3].gencol[2].genblk1.c.bufs[0].A ;
 wire \genrow[3].gencol[3].genblk1.c.bufs[0].A ;
 wire \genrow[3].gencol[4].genblk1.c.bufs[0].A ;
 wire \genrow[3].gencol[5].genblk1.c.bufs[0].A ;
 wire \genrow[4].gencol[0].genblk1.c.bufs[0].A ;
 wire \genrow[4].gencol[1].genblk1.c.bufs[0].A ;
 wire \genrow[4].gencol[2].genblk1.c.bufs[0].A ;
 wire \genrow[4].gencol[3].genblk1.c.bufs[0].A ;
 wire \genrow[4].gencol[4].genblk1.c.bufs[0].A ;
 wire \genrow[4].gencol[5].genblk1.c.bufs[0].A ;
 wire \genrow[5].gencol[0].genblk1.c.bufs[0].A ;
 wire \genrow[5].gencol[1].genblk1.c.bufs[0].A ;
 wire \genrow[5].gencol[2].genblk1.c.bufs[0].A ;
 wire \genrow[5].gencol[3].genblk1.c.bufs[0].A ;
 wire \genrow[5].gencol[4].genblk1.c.bufs[0].A ;
 wire \genrow[6].gencol[0].genblk1.c.bufs[0].A ;
 wire \genrow[6].gencol[1].genblk1.c.bufs[0].A ;
 wire \genrow[6].gencol[2].genblk1.c.bufs[0].A ;
 wire \genrow[6].gencol[3].genblk1.c.bufs[0].A ;
 wire \genrow[6].gencol[5].genblk1.c.bufs[0].A ;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_5_0__leaf_clk;
 wire clknet_5_1__leaf_clk;
 wire clknet_5_2__leaf_clk;
 wire clknet_5_3__leaf_clk;
 wire clknet_5_4__leaf_clk;
 wire clknet_5_5__leaf_clk;
 wire clknet_5_6__leaf_clk;
 wire clknet_5_7__leaf_clk;
 wire clknet_5_8__leaf_clk;
 wire clknet_5_9__leaf_clk;
 wire clknet_5_10__leaf_clk;
 wire clknet_5_11__leaf_clk;
 wire clknet_5_12__leaf_clk;
 wire clknet_5_13__leaf_clk;
 wire clknet_5_14__leaf_clk;
 wire clknet_5_15__leaf_clk;
 wire clknet_5_16__leaf_clk;
 wire clknet_5_17__leaf_clk;
 wire clknet_5_18__leaf_clk;
 wire clknet_5_19__leaf_clk;
 wire clknet_5_20__leaf_clk;
 wire clknet_5_21__leaf_clk;
 wire clknet_5_22__leaf_clk;
 wire clknet_5_23__leaf_clk;
 wire clknet_5_24__leaf_clk;
 wire clknet_5_25__leaf_clk;
 wire clknet_5_26__leaf_clk;
 wire clknet_5_27__leaf_clk;
 wire clknet_5_28__leaf_clk;
 wire clknet_5_29__leaf_clk;
 wire clknet_5_30__leaf_clk;
 wire clknet_5_31__leaf_clk;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net180;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;

 sg13g2_inv_1 _1169_ (.Y(_0334_),
    .A(\cell_cfg[20][3] ));
 sg13g2_inv_1 _1170_ (.Y(_0335_),
    .A(\cell_cfg[12][3] ));
 sg13g2_inv_1 _1171_ (.Y(_0336_),
    .A(\cell_cfg[21][3] ));
 sg13g2_inv_1 _1172_ (.Y(_0337_),
    .A(\cell_cfg[22][3] ));
 sg13g2_inv_1 _1173_ (.Y(_0338_),
    .A(\cell_cfg[23][2] ));
 sg13g2_inv_1 _1174_ (.Y(_0339_),
    .A(net468));
 sg13g2_inv_1 _1175_ (.Y(_0340_),
    .A(net438));
 sg13g2_inv_1 _1176_ (.Y(_0341_),
    .A(\cell_cfg[25][3] ));
 sg13g2_inv_1 _1177_ (.Y(_0342_),
    .A(net392));
 sg13g2_inv_1 _1178_ (.Y(_0343_),
    .A(net245));
 sg13g2_inv_1 _1179_ (.Y(_0344_),
    .A(\cell_cfg[26][3] ));
 sg13g2_inv_1 _1180_ (.Y(_0345_),
    .A(net249));
 sg13g2_inv_1 _1181_ (.Y(_0346_),
    .A(net334));
 sg13g2_inv_1 _1182_ (.Y(_0347_),
    .A(\cell_cfg[27][3] ));
 sg13g2_inv_1 _1183_ (.Y(_0348_),
    .A(\cell_cfg[28][2] ));
 sg13g2_inv_1 _1184_ (.Y(_0349_),
    .A(\cell_cfg[30][3] ));
 sg13g2_inv_1 _1185_ (.Y(_0350_),
    .A(\cell_cfg[31][3] ));
 sg13g2_inv_1 _1186_ (.Y(_0351_),
    .A(\cell_cfg[35][3] ));
 sg13g2_inv_1 _1187_ (.Y(_0352_),
    .A(\cell_cfg[35][2] ));
 sg13g2_inv_1 _1188_ (.Y(_0353_),
    .A(\cell_cfg[2][2] ));
 sg13g2_inv_1 _1189_ (.Y(_0354_),
    .A(\cell_cfg[10][3] ));
 sg13g2_inv_1 _1190_ (.Y(_0355_),
    .A(\cell_cfg[14][3] ));
 sg13g2_inv_1 _1191_ (.Y(_0356_),
    .A(\cell_cfg[1][2] ));
 sg13g2_inv_1 _1192_ (.Y(_0357_),
    .A(\cell_cfg[9][3] ));
 sg13g2_inv_1 _1193_ (.Y(_0358_),
    .A(net223));
 sg13g2_inv_1 _1194_ (.Y(_0359_),
    .A(net439));
 sg13g2_inv_1 _1195_ (.Y(_0360_),
    .A(\cell_cfg[0][3] ));
 sg13g2_inv_1 _1196_ (.Y(_0361_),
    .A(\cell_cfg[8][3] ));
 sg13g2_inv_2 _1197_ (.Y(_0362_),
    .A(net318));
 sg13g2_inv_1 _1198_ (.Y(_0363_),
    .A(\cell_cfg[3][1] ));
 sg13g2_inv_1 _1199_ (.Y(_0364_),
    .A(\cell_cfg[4][0] ));
 sg13g2_inv_1 _1200_ (.Y(_0365_),
    .A(\cell_cfg[6][1] ));
 sg13g2_inv_1 _1201_ (.Y(_0366_),
    .A(\cell_cfg[8][0] ));
 sg13g2_inv_1 _1202_ (.Y(_0367_),
    .A(\cell_cfg[10][0] ));
 sg13g2_inv_1 _1203_ (.Y(_0368_),
    .A(\cell_cfg[11][0] ));
 sg13g2_inv_1 _1204_ (.Y(_0369_),
    .A(\cell_cfg[12][0] ));
 sg13g2_inv_1 _1205_ (.Y(_0370_),
    .A(\cell_cfg[14][0] ));
 sg13g2_inv_1 _1206_ (.Y(_0371_),
    .A(\cell_cfg[20][0] ));
 sg13g2_inv_1 _1207_ (.Y(_0372_),
    .A(net398));
 sg13g2_inv_1 _1208_ (.Y(_0373_),
    .A(\cell_cfg[26][0] ));
 sg13g2_inv_1 _1209_ (.Y(_0374_),
    .A(\cell_cfg[28][1] ));
 sg13g2_inv_1 _1210_ (.Y(_0375_),
    .A(\cell_cfg[29][1] ));
 sg13g2_inv_1 _1211_ (.Y(_0376_),
    .A(\cell_cfg[32][1] ));
 sg13g2_inv_1 _1212_ (.Y(_0377_),
    .A(\cell_cfg[32][0] ));
 sg13g2_inv_1 _1213_ (.Y(_0378_),
    .A(net459));
 sg13g2_inv_1 _1214_ (.Y(_0379_),
    .A(\cell_cfg[35][0] ));
 sg13g2_inv_1 _1215_ (.Y(_0380_),
    .A(\cell_cfg[19][3] ));
 sg13g2_inv_1 _1216_ (.Y(_0381_),
    .A(net382));
 sg13g2_inv_1 _1217_ (.Y(_0382_),
    .A(net388));
 sg13g2_inv_1 _1218_ (.Y(_0383_),
    .A(net346));
 sg13g2_inv_1 _1219_ (.Y(_0384_),
    .A(net374));
 sg13g2_inv_1 _1220_ (.Y(_0385_),
    .A(\cell_cfg[7][3] ));
 sg13g2_inv_1 _1221_ (.Y(_0386_),
    .A(net376));
 sg13g2_inv_1 _1222_ (.Y(_0387_),
    .A(net401));
 sg13g2_inv_1 _1223_ (.Y(_0388_),
    .A(\cell_cfg[18][3] ));
 sg13g2_inv_1 _1224_ (.Y(_0389_),
    .A(net349));
 sg13g2_inv_1 _1225_ (.Y(_0390_),
    .A(net355));
 sg13g2_inv_1 _1226_ (.Y(_0391_),
    .A(net405));
 sg13g2_inv_1 _1227_ (.Y(_0392_),
    .A(net380));
 sg13g2_inv_1 _1228_ (.Y(_0393_),
    .A(net486));
 sg13g2_inv_2 _1229_ (.Y(_0394_),
    .A(net253));
 sg13g2_inv_1 _1230_ (.Y(_0395_),
    .A(net3));
 sg13g2_inv_1 _1231_ (.Y(_0396_),
    .A(net328));
 sg13g2_inv_4 _1232_ (.A(\genrow[6].gencol[0].genblk1.c.bufs[0].A ),
    .Y(_0397_));
 sg13g2_inv_2 _1233_ (.Y(_0398_),
    .A(net172));
 sg13g2_inv_2 _1234_ (.Y(_0399_),
    .A(\genrow[2].gencol[0].genblk1.c.bufs[0].A ));
 sg13g2_inv_1 _1235_ (.Y(_0400_),
    .A(\genrow[2].gencol[1].genblk1.c.bufs[0].A ));
 sg13g2_inv_2 _1236_ (.Y(_0401_),
    .A(\genrow[2].gencol[2].genblk1.c.bufs[0].A ));
 sg13g2_inv_2 _1237_ (.Y(_0402_),
    .A(\genrow[2].gencol[3].genblk1.c.bufs[0].A ));
 sg13g2_inv_1 _1238_ (.Y(_0403_),
    .A(\genrow[3].gencol[0].genblk1.c.bufs[0].A ));
 sg13g2_inv_1 _1239_ (.Y(_0404_),
    .A(\genrow[3].gencol[1].genblk1.c.bufs[0].A ));
 sg13g2_inv_1 _1240_ (.Y(_0405_),
    .A(\genrow[3].gencol[2].genblk1.c.bufs[0].A ));
 sg13g2_inv_1 _1241_ (.Y(_0406_),
    .A(\genrow[3].gencol[3].genblk1.c.bufs[0].A ));
 sg13g2_inv_1 _1242_ (.Y(_0407_),
    .A(\genrow[3].gencol[4].genblk1.c.bufs[0].A ));
 sg13g2_inv_1 _1243_ (.Y(_0408_),
    .A(\genrow[3].gencol[5].genblk1.c.bufs[0].A ));
 sg13g2_inv_2 _1244_ (.Y(_0409_),
    .A(\genrow[4].gencol[0].genblk1.c.bufs[0].A ));
 sg13g2_inv_1 _1245_ (.Y(_0410_),
    .A(\genrow[4].gencol[1].genblk1.c.bufs[0].A ));
 sg13g2_inv_1 _1246_ (.Y(_0411_),
    .A(\genrow[4].gencol[2].genblk1.c.bufs[0].A ));
 sg13g2_inv_1 _1247_ (.Y(_0412_),
    .A(\genrow[4].gencol[3].genblk1.c.bufs[0].A ));
 sg13g2_inv_1 _1248_ (.Y(_0413_),
    .A(\genrow[4].gencol[4].genblk1.c.bufs[0].A ));
 sg13g2_inv_1 _1249_ (.Y(_0414_),
    .A(net199));
 sg13g2_inv_2 _1250_ (.Y(_0415_),
    .A(\genrow[5].gencol[0].genblk1.c.bufs[0].A ));
 sg13g2_inv_2 _1251_ (.Y(_0416_),
    .A(\genrow[5].gencol[1].genblk1.c.bufs[0].A ));
 sg13g2_inv_1 _1252_ (.Y(_0417_),
    .A(\genrow[5].gencol[2].genblk1.c.bufs[0].A ));
 sg13g2_inv_1 _1253_ (.Y(_0418_),
    .A(\genrow[5].gencol[3].genblk1.c.bufs[0].A ));
 sg13g2_inv_1 _1254_ (.Y(_0419_),
    .A(net174));
 sg13g2_inv_1 _1255_ (.Y(_0420_),
    .A(\genrow[6].gencol[1].genblk1.c.bufs[0].A ));
 sg13g2_inv_4 _1256_ (.A(\genrow[1].gencol[0].genblk1.c.bufs[0].A ),
    .Y(_0421_));
 sg13g2_inv_1 _1257_ (.Y(_0422_),
    .A(\genrow[1].gencol[1].genblk1.c.bufs[0].A ));
 sg13g2_inv_1 _1258_ (.Y(_0423_),
    .A(\genrow[1].gencol[2].genblk1.c.bufs[0].A ));
 sg13g2_inv_1 _1259_ (.Y(_0424_),
    .A(\genrow[1].gencol[3].genblk1.c.bufs[0].A ));
 sg13g2_inv_1 _1260_ (.Y(_0425_),
    .A(\genrow[1].gencol[4].genblk1.c.bufs[0].A ));
 sg13g2_mux4_1 _1261_ (.S0(\cell_cfg[34][1] ),
    .A0(net208),
    .A1(net172),
    .A2(net318),
    .A3(\genrow[6].gencol[0].genblk1.c.bufs[0].A ),
    .S1(\cell_cfg[34][0] ),
    .X(_0426_));
 sg13g2_and2_1 _1262_ (.A(\cell_cfg[34][1] ),
    .B(\genrow[6].gencol[3].genblk1.c.bufs[0].A ),
    .X(_0427_));
 sg13g2_mux4_1 _1263_ (.S0(\cell_cfg[34][2] ),
    .A0(\cell_cfg[34][0] ),
    .A1(_0426_),
    .A2(_0427_),
    .A3(net208),
    .S1(\cell_cfg[34][3] ),
    .X(_0428_));
 sg13g2_and2_2 _1264_ (.A(_0394_),
    .B(_0428_),
    .X(_0429_));
 sg13g2_nand4_1 _1265_ (.B(\cell_cfg[29][0] ),
    .C(_0394_),
    .A(\cell_cfg[29][1] ),
    .Y(_0430_),
    .D(_0428_));
 sg13g2_o21ai_1 _1266_ (.B1(\cell_cfg[29][0] ),
    .Y(_0431_),
    .A1(\cell_cfg[29][1] ),
    .A2(_0398_));
 sg13g2_o21ai_1 _1267_ (.B1(_0431_),
    .Y(_0432_),
    .A1(_0375_),
    .A2(net216));
 sg13g2_nor2_1 _1268_ (.A(\cell_cfg[29][1] ),
    .B(\cell_cfg[29][0] ),
    .Y(_0433_));
 sg13g2_a221oi_1 _1269_ (.B2(_0414_),
    .C1(\cell_cfg[29][3] ),
    .B1(_0433_),
    .A1(_0430_),
    .Y(_0434_),
    .A2(_0432_));
 sg13g2_nand2_1 _1270_ (.Y(_0435_),
    .A(\cell_cfg[29][3] ),
    .B(\genrow[4].gencol[5].genblk1.c.bufs[0].A ));
 sg13g2_nand2_1 _1271_ (.Y(_0436_),
    .A(\cell_cfg[29][1] ),
    .B(net175));
 sg13g2_nor2b_1 _1272_ (.A(\cell_cfg[29][2] ),
    .B_N(\cell_cfg[29][3] ),
    .Y(_0437_));
 sg13g2_a22oi_1 _1273_ (.Y(_0438_),
    .B1(_0436_),
    .B2(_0437_),
    .A2(_0435_),
    .A1(\cell_cfg[29][2] ));
 sg13g2_nor3_1 _1274_ (.A(\cell_cfg[29][3] ),
    .B(\cell_cfg[29][2] ),
    .C(\cell_cfg[29][0] ),
    .Y(_0439_));
 sg13g2_nor2_1 _1275_ (.A(net255),
    .B(_0439_),
    .Y(_0440_));
 sg13g2_o21ai_1 _1276_ (.B1(_0440_),
    .Y(_0441_),
    .A1(_0434_),
    .A2(_0438_));
 sg13g2_nand2b_1 _1277_ (.Y(_0442_),
    .B(\cell_cfg[28][1] ),
    .A_N(\cell_cfg[28][0] ));
 sg13g2_nand3_1 _1278_ (.B(\cell_cfg[28][0] ),
    .C(net216),
    .A(\cell_cfg[28][1] ),
    .Y(_0443_));
 sg13g2_o21ai_1 _1279_ (.B1(_0443_),
    .Y(_0444_),
    .A1(\cell_cfg[28][1] ),
    .A2(\cell_cfg[28][0] ));
 sg13g2_a21oi_1 _1280_ (.A1(_0374_),
    .A2(_0429_),
    .Y(_0445_),
    .B1(_0444_));
 sg13g2_o21ai_1 _1281_ (.B1(_0445_),
    .Y(_0446_),
    .A1(_0441_),
    .A2(_0442_));
 sg13g2_nor3_1 _1282_ (.A(\cell_cfg[28][1] ),
    .B(\cell_cfg[28][0] ),
    .C(net222),
    .Y(_0447_));
 sg13g2_nor3_1 _1283_ (.A(\cell_cfg[28][3] ),
    .B(_0348_),
    .C(_0447_),
    .Y(_0448_));
 sg13g2_nand2_1 _1284_ (.Y(_0449_),
    .A(\cell_cfg[28][3] ),
    .B(net222));
 sg13g2_nand2_1 _1285_ (.Y(_0450_),
    .A(\cell_cfg[28][1] ),
    .B(\genrow[5].gencol[3].genblk1.c.bufs[0].A ));
 sg13g2_nor2b_1 _1286_ (.A(\cell_cfg[28][2] ),
    .B_N(\cell_cfg[28][3] ),
    .Y(_0451_));
 sg13g2_a22oi_1 _1287_ (.Y(_0452_),
    .B1(_0450_),
    .B2(_0451_),
    .A2(_0449_),
    .A1(\cell_cfg[28][2] ));
 sg13g2_a21oi_1 _1288_ (.A1(_0446_),
    .A2(_0448_),
    .Y(_0453_),
    .B1(_0452_));
 sg13g2_nor3_1 _1289_ (.A(\cell_cfg[28][3] ),
    .B(\cell_cfg[28][2] ),
    .C(\cell_cfg[28][0] ),
    .Y(_0454_));
 sg13g2_nor3_2 _1290_ (.A(_0453_),
    .B(net255),
    .C(_0454_),
    .Y(\genrow[5].gencol[4].genblk1.c.bufs[0].A ));
 sg13g2_and2_1 _1291_ (.A(\cell_cfg[33][1] ),
    .B(\genrow[6].gencol[2].genblk1.c.bufs[0].A ),
    .X(_0455_));
 sg13g2_mux4_1 _1292_ (.S0(\cell_cfg[33][1] ),
    .A0(\genrow[5].gencol[3].genblk1.c.bufs[0].A ),
    .A1(_0429_),
    .A2(net318),
    .A3(\genrow[6].gencol[0].genblk1.c.bufs[0].A ),
    .S1(\cell_cfg[33][0] ),
    .X(_0456_));
 sg13g2_nor2_1 _1293_ (.A(net336),
    .B(net330),
    .Y(_0457_));
 sg13g2_mux4_1 _1294_ (.S0(\cell_cfg[33][3] ),
    .A0(\cell_cfg[33][0] ),
    .A1(_0455_),
    .A2(_0456_),
    .A3(\genrow[5].gencol[3].genblk1.c.bufs[0].A ),
    .S1(\cell_cfg[33][2] ),
    .X(_0458_));
 sg13g2_and2_2 _1295_ (.A(_0394_),
    .B(_0458_),
    .X(\genrow[6].gencol[3].genblk1.c.bufs[0].A ));
 sg13g2_o21ai_1 _1296_ (.B1(_0349_),
    .Y(_0459_),
    .A1(\cell_cfg[30][1] ),
    .A2(\cell_cfg[30][0] ));
 sg13g2_a21oi_1 _1297_ (.A1(\cell_cfg[30][1] ),
    .A2(\genrow[6].gencol[5].genblk1.c.bufs[0].A ),
    .Y(_0460_),
    .B1(\cell_cfg[30][2] ));
 sg13g2_a21oi_1 _1298_ (.A1(\cell_cfg[30][2] ),
    .A2(_0415_),
    .Y(_0461_),
    .B1(_0460_));
 sg13g2_nand3_1 _1299_ (.B(\cell_cfg[30][0] ),
    .C(_0397_),
    .A(\cell_cfg[30][1] ),
    .Y(_0462_));
 sg13g2_o21ai_1 _1300_ (.B1(_0462_),
    .Y(_0463_),
    .A1(net318),
    .A2(\cell_cfg[30][1] ));
 sg13g2_a21o_1 _1301_ (.A2(net180),
    .A1(\cell_cfg[30][2] ),
    .B1(\cell_cfg[30][0] ),
    .X(_0464_));
 sg13g2_a21oi_1 _1302_ (.A1(\cell_cfg[30][2] ),
    .A2(_0463_),
    .Y(_0465_),
    .B1(_0459_));
 sg13g2_a22oi_1 _1303_ (.Y(_0466_),
    .B1(_0464_),
    .B2(_0465_),
    .A2(_0461_),
    .A1(_0459_));
 sg13g2_nor2_2 _1304_ (.A(net252),
    .B(_0466_),
    .Y(\genrow[6].gencol[0].genblk1.c.bufs[0].A ));
 sg13g2_mux4_1 _1305_ (.S0(\cell_cfg[35][1] ),
    .A0(_0362_),
    .A1(_0398_),
    .A2(net201),
    .A3(_0397_),
    .S1(_0379_),
    .X(_0467_));
 sg13g2_nand2b_1 _1306_ (.Y(_0468_),
    .B(_0351_),
    .A_N(_0467_));
 sg13g2_nor3_1 _1307_ (.A(_0351_),
    .B(_0352_),
    .C(net201),
    .Y(_0469_));
 sg13g2_nor2_1 _1308_ (.A(\cell_cfg[35][3] ),
    .B(\cell_cfg[35][2] ),
    .Y(_0470_));
 sg13g2_nor2_1 _1309_ (.A(\cell_cfg[35][2] ),
    .B(_0378_),
    .Y(_0471_));
 sg13g2_a221oi_1 _1310_ (.B2(_0471_),
    .C1(_0469_),
    .B1(_0429_),
    .A1(_0351_),
    .Y(_0472_),
    .A2(_0352_));
 sg13g2_a221oi_1 _1311_ (.B2(_0472_),
    .C1(net252),
    .B1(_0468_),
    .A1(_0379_),
    .Y(\genrow[6].gencol[5].genblk1.c.bufs[0].A ),
    .A2(_0470_));
 sg13g2_o21ai_1 _1312_ (.B1(_0347_),
    .Y(_0473_),
    .A1(\cell_cfg[27][1] ),
    .A2(\cell_cfg[27][0] ));
 sg13g2_a21oi_1 _1313_ (.A1(\cell_cfg[27][1] ),
    .A2(\genrow[5].gencol[2].genblk1.c.bufs[0].A ),
    .Y(_0474_),
    .B1(\cell_cfg[27][2] ));
 sg13g2_a21oi_1 _1314_ (.A1(\cell_cfg[27][2] ),
    .A2(_0412_),
    .Y(_0475_),
    .B1(_0474_));
 sg13g2_nand3_1 _1315_ (.B(\cell_cfg[27][0] ),
    .C(_0415_),
    .A(\cell_cfg[27][1] ),
    .Y(_0476_));
 sg13g2_o21ai_1 _1316_ (.B1(_0476_),
    .Y(_0477_),
    .A1(\cell_cfg[27][1] ),
    .A2(\genrow[6].gencol[3].genblk1.c.bufs[0].A ));
 sg13g2_a21o_1 _1317_ (.A2(\genrow[5].gencol[4].genblk1.c.bufs[0].A ),
    .A1(\cell_cfg[27][2] ),
    .B1(\cell_cfg[27][0] ),
    .X(_0478_));
 sg13g2_a21oi_1 _1318_ (.A1(\cell_cfg[27][2] ),
    .A2(_0477_),
    .Y(_0479_),
    .B1(_0473_));
 sg13g2_a22oi_1 _1319_ (.Y(_0480_),
    .B1(_0478_),
    .B2(_0479_),
    .A2(_0475_),
    .A1(_0473_));
 sg13g2_nor2_2 _1320_ (.A(net255),
    .B(_0480_),
    .Y(\genrow[5].gencol[3].genblk1.c.bufs[0].A ));
 sg13g2_a21oi_1 _1321_ (.A1(\cell_cfg[32][1] ),
    .A2(\genrow[6].gencol[1].genblk1.c.bufs[0].A ),
    .Y(_0481_),
    .B1(\cell_cfg[32][2] ));
 sg13g2_a21o_1 _1322_ (.A2(_0377_),
    .A1(_0376_),
    .B1(\cell_cfg[32][3] ),
    .X(_0482_));
 sg13g2_a21oi_1 _1323_ (.A1(\cell_cfg[32][2] ),
    .A2(_0417_),
    .Y(_0483_),
    .B1(_0481_));
 sg13g2_nand3_1 _1324_ (.B(\cell_cfg[32][0] ),
    .C(_0397_),
    .A(\cell_cfg[32][1] ),
    .Y(_0484_));
 sg13g2_o21ai_1 _1325_ (.B1(_0484_),
    .Y(_0485_),
    .A1(net318),
    .A2(\cell_cfg[32][1] ));
 sg13g2_nand2_1 _1326_ (.Y(_0486_),
    .A(\cell_cfg[32][2] ),
    .B(\genrow[6].gencol[3].genblk1.c.bufs[0].A ));
 sg13g2_a221oi_1 _1327_ (.B2(_0377_),
    .C1(_0482_),
    .B1(_0486_),
    .A1(\cell_cfg[32][2] ),
    .Y(_0487_),
    .A2(_0485_));
 sg13g2_a21oi_1 _1328_ (.A1(_0482_),
    .A2(_0483_),
    .Y(_0488_),
    .B1(_0487_));
 sg13g2_nor2_2 _1329_ (.A(net252),
    .B(_0488_),
    .Y(\genrow[6].gencol[2].genblk1.c.bufs[0].A ));
 sg13g2_a21oi_1 _1330_ (.A1(\cell_cfg[26][1] ),
    .A2(\genrow[5].gencol[1].genblk1.c.bufs[0].A ),
    .Y(_0489_),
    .B1(\cell_cfg[26][2] ));
 sg13g2_o21ai_1 _1331_ (.B1(_0344_),
    .Y(_0490_),
    .A1(\cell_cfg[26][1] ),
    .A2(\cell_cfg[26][0] ));
 sg13g2_a21oi_1 _1332_ (.A1(\cell_cfg[26][2] ),
    .A2(_0411_),
    .Y(_0491_),
    .B1(_0489_));
 sg13g2_nand3_1 _1333_ (.B(\cell_cfg[26][0] ),
    .C(_0415_),
    .A(\cell_cfg[26][1] ),
    .Y(_0492_));
 sg13g2_o21ai_1 _1334_ (.B1(_0492_),
    .Y(_0493_),
    .A1(\cell_cfg[26][1] ),
    .A2(net214));
 sg13g2_nand3_1 _1335_ (.B(\cell_cfg[26][1] ),
    .C(\genrow[5].gencol[3].genblk1.c.bufs[0].A ),
    .A(\cell_cfg[26][2] ),
    .Y(_0494_));
 sg13g2_a22oi_1 _1336_ (.Y(_0495_),
    .B1(_0494_),
    .B2(_0373_),
    .A2(_0493_),
    .A1(\cell_cfg[26][2] ));
 sg13g2_a22oi_1 _1337_ (.Y(_0496_),
    .B1(_0495_),
    .B2(_0344_),
    .A2(_0491_),
    .A1(_0490_));
 sg13g2_nor2_2 _1338_ (.A(net251),
    .B(_0496_),
    .Y(\genrow[5].gencol[2].genblk1.c.bufs[0].A ));
 sg13g2_nand3_1 _1339_ (.B(\cell_cfg[31][0] ),
    .C(_0420_),
    .A(\cell_cfg[31][1] ),
    .Y(_0497_));
 sg13g2_o21ai_1 _1340_ (.B1(_0497_),
    .Y(_0498_),
    .A1(net318),
    .A2(\cell_cfg[31][1] ));
 sg13g2_a21o_1 _1341_ (.A2(\genrow[6].gencol[2].genblk1.c.bufs[0].A ),
    .A1(\cell_cfg[31][2] ),
    .B1(\cell_cfg[31][0] ),
    .X(_0499_));
 sg13g2_o21ai_1 _1342_ (.B1(_0350_),
    .Y(_0500_),
    .A1(\cell_cfg[31][1] ),
    .A2(\cell_cfg[31][0] ));
 sg13g2_a21oi_1 _1343_ (.A1(\cell_cfg[31][2] ),
    .A2(_0498_),
    .Y(_0501_),
    .B1(_0500_));
 sg13g2_a21oi_1 _1344_ (.A1(\cell_cfg[31][1] ),
    .A2(\genrow[6].gencol[0].genblk1.c.bufs[0].A ),
    .Y(_0502_),
    .B1(\cell_cfg[31][2] ));
 sg13g2_a21oi_1 _1345_ (.A1(\cell_cfg[31][2] ),
    .A2(_0416_),
    .Y(_0503_),
    .B1(_0502_));
 sg13g2_a22oi_1 _1346_ (.Y(_0504_),
    .B1(_0503_),
    .B2(_0500_),
    .A2(_0501_),
    .A1(_0499_));
 sg13g2_nor2_2 _1347_ (.A(net252),
    .B(_0504_),
    .Y(\genrow[6].gencol[1].genblk1.c.bufs[0].A ));
 sg13g2_nand3_1 _1348_ (.B(\cell_cfg[25][0] ),
    .C(_0397_),
    .A(\cell_cfg[25][1] ),
    .Y(_0505_));
 sg13g2_o21ai_1 _1349_ (.B1(_0505_),
    .Y(_0506_),
    .A1(\cell_cfg[25][1] ),
    .A2(net180));
 sg13g2_a21o_1 _1350_ (.A2(\genrow[5].gencol[2].genblk1.c.bufs[0].A ),
    .A1(\cell_cfg[25][2] ),
    .B1(\cell_cfg[25][0] ),
    .X(_0507_));
 sg13g2_o21ai_1 _1351_ (.B1(_0341_),
    .Y(_0508_),
    .A1(\cell_cfg[25][1] ),
    .A2(\cell_cfg[25][0] ));
 sg13g2_a21oi_1 _1352_ (.A1(\cell_cfg[25][2] ),
    .A2(_0506_),
    .Y(_0509_),
    .B1(_0508_));
 sg13g2_a21oi_1 _1353_ (.A1(\cell_cfg[25][1] ),
    .A2(\genrow[5].gencol[0].genblk1.c.bufs[0].A ),
    .Y(_0510_),
    .B1(\cell_cfg[25][2] ));
 sg13g2_a21oi_1 _1354_ (.A1(\cell_cfg[25][2] ),
    .A2(_0410_),
    .Y(_0511_),
    .B1(_0510_));
 sg13g2_a22oi_1 _1355_ (.Y(_0512_),
    .B1(_0511_),
    .B2(_0508_),
    .A2(_0509_),
    .A1(_0507_));
 sg13g2_nor2_1 _1356_ (.A(net251),
    .B(_0512_),
    .Y(\genrow[5].gencol[1].genblk1.c.bufs[0].A ));
 sg13g2_nor3_1 _1357_ (.A(\cell_cfg[24][2] ),
    .B(_0372_),
    .C(net212),
    .Y(_0513_));
 sg13g2_nor2_1 _1358_ (.A(\cell_cfg[24][0] ),
    .B(\genrow[5].gencol[1].genblk1.c.bufs[0].A ),
    .Y(_0514_));
 sg13g2_a21oi_1 _1359_ (.A1(\cell_cfg[24][0] ),
    .A2(_0398_),
    .Y(_0515_),
    .B1(_0514_));
 sg13g2_nor2_1 _1360_ (.A(\cell_cfg[24][1] ),
    .B(_0397_),
    .Y(_0516_));
 sg13g2_a22oi_1 _1361_ (.Y(_0517_),
    .B1(_0516_),
    .B2(\cell_cfg[24][0] ),
    .A2(_0515_),
    .A1(\cell_cfg[24][1] ));
 sg13g2_o21ai_1 _1362_ (.B1(_0339_),
    .Y(_0518_),
    .A1(\cell_cfg[24][1] ),
    .A2(\cell_cfg[24][0] ));
 sg13g2_and3_1 _1363_ (.X(_0519_),
    .A(\cell_cfg[24][2] ),
    .B(net210),
    .C(_0518_));
 sg13g2_a21oi_1 _1364_ (.A1(\cell_cfg[24][2] ),
    .A2(_0517_),
    .Y(_0520_),
    .B1(\cell_cfg[24][3] ));
 sg13g2_nor3_1 _1365_ (.A(_0513_),
    .B(_0519_),
    .C(_0520_),
    .Y(_0521_));
 sg13g2_nor3_1 _1366_ (.A(\cell_cfg[24][3] ),
    .B(\cell_cfg[24][2] ),
    .C(\cell_cfg[24][0] ),
    .Y(_0522_));
 sg13g2_nor3_2 _1367_ (.A(net251),
    .B(_0521_),
    .C(_0522_),
    .Y(\genrow[5].gencol[0].genblk1.c.bufs[0].A ));
 sg13g2_nand3_1 _1368_ (.B(\cell_cfg[23][0] ),
    .C(\genrow[6].gencol[3].genblk1.c.bufs[0].A ),
    .A(\cell_cfg[23][1] ),
    .Y(_0523_));
 sg13g2_a21oi_1 _1369_ (.A1(\cell_cfg[23][1] ),
    .A2(_0409_),
    .Y(_0524_),
    .B1(\cell_cfg[23][0] ));
 sg13g2_nor2b_1 _1370_ (.A(_0524_),
    .B_N(_0523_),
    .Y(_0525_));
 sg13g2_o21ai_1 _1371_ (.B1(_0525_),
    .Y(_0526_),
    .A1(\cell_cfg[23][1] ),
    .A2(net200));
 sg13g2_nor3_1 _1372_ (.A(\cell_cfg[23][1] ),
    .B(\cell_cfg[23][0] ),
    .C(net211),
    .Y(_0527_));
 sg13g2_nor3_1 _1373_ (.A(\cell_cfg[23][3] ),
    .B(_0338_),
    .C(_0527_),
    .Y(_0528_));
 sg13g2_nand2_1 _1374_ (.Y(_0529_),
    .A(\cell_cfg[23][3] ),
    .B(net211));
 sg13g2_nand2_1 _1375_ (.Y(_0530_),
    .A(\cell_cfg[23][1] ),
    .B(\genrow[4].gencol[4].genblk1.c.bufs[0].A ));
 sg13g2_nor2b_1 _1376_ (.A(\cell_cfg[23][2] ),
    .B_N(\cell_cfg[23][3] ),
    .Y(_0531_));
 sg13g2_a22oi_1 _1377_ (.Y(_0532_),
    .B1(_0530_),
    .B2(_0531_),
    .A2(_0529_),
    .A1(\cell_cfg[23][2] ));
 sg13g2_a21oi_1 _1378_ (.A1(_0526_),
    .A2(_0528_),
    .Y(_0533_),
    .B1(_0532_));
 sg13g2_nor3_1 _1379_ (.A(\cell_cfg[23][3] ),
    .B(\cell_cfg[23][2] ),
    .C(\cell_cfg[23][0] ),
    .Y(_0534_));
 sg13g2_nor3_2 _1380_ (.A(net251),
    .B(_0533_),
    .C(_0534_),
    .Y(\genrow[4].gencol[5].genblk1.c.bufs[0].A ));
 sg13g2_o21ai_1 _1381_ (.B1(_0337_),
    .Y(_0535_),
    .A1(\cell_cfg[22][1] ),
    .A2(\cell_cfg[22][0] ));
 sg13g2_a21oi_1 _1382_ (.A1(\cell_cfg[22][1] ),
    .A2(\genrow[4].gencol[3].genblk1.c.bufs[0].A ),
    .Y(_0536_),
    .B1(\cell_cfg[22][2] ));
 sg13g2_a21oi_1 _1383_ (.A1(\cell_cfg[22][2] ),
    .A2(_0407_),
    .Y(_0537_),
    .B1(_0536_));
 sg13g2_nand3_1 _1384_ (.B(\cell_cfg[22][0] ),
    .C(_0409_),
    .A(\cell_cfg[22][1] ),
    .Y(_0538_));
 sg13g2_o21ai_1 _1385_ (.B1(_0538_),
    .Y(_0539_),
    .A1(\cell_cfg[22][1] ),
    .A2(\genrow[5].gencol[4].genblk1.c.bufs[0].A ));
 sg13g2_a21o_1 _1386_ (.A2(\genrow[4].gencol[5].genblk1.c.bufs[0].A ),
    .A1(\cell_cfg[22][2] ),
    .B1(\cell_cfg[22][0] ),
    .X(_0540_));
 sg13g2_a21oi_1 _1387_ (.A1(\cell_cfg[22][2] ),
    .A2(_0539_),
    .Y(_0541_),
    .B1(_0535_));
 sg13g2_a22oi_1 _1388_ (.Y(_0542_),
    .B1(_0540_),
    .B2(_0541_),
    .A2(_0537_),
    .A1(_0535_));
 sg13g2_nor2_2 _1389_ (.A(net251),
    .B(_0542_),
    .Y(\genrow[4].gencol[4].genblk1.c.bufs[0].A ));
 sg13g2_o21ai_1 _1390_ (.B1(_0336_),
    .Y(_0543_),
    .A1(\cell_cfg[21][1] ),
    .A2(\cell_cfg[21][0] ));
 sg13g2_a21oi_1 _1391_ (.A1(\cell_cfg[21][1] ),
    .A2(\genrow[4].gencol[2].genblk1.c.bufs[0].A ),
    .Y(_0544_),
    .B1(\cell_cfg[21][2] ));
 sg13g2_a21oi_1 _1392_ (.A1(\cell_cfg[21][2] ),
    .A2(_0406_),
    .Y(_0545_),
    .B1(_0544_));
 sg13g2_nand3_1 _1393_ (.B(\cell_cfg[21][0] ),
    .C(_0409_),
    .A(\cell_cfg[21][1] ),
    .Y(_0546_));
 sg13g2_o21ai_1 _1394_ (.B1(_0546_),
    .Y(_0547_),
    .A1(\cell_cfg[21][1] ),
    .A2(net209));
 sg13g2_a21o_1 _1395_ (.A2(\genrow[4].gencol[4].genblk1.c.bufs[0].A ),
    .A1(\cell_cfg[21][2] ),
    .B1(\cell_cfg[21][0] ),
    .X(_0548_));
 sg13g2_a21oi_1 _1396_ (.A1(\cell_cfg[21][2] ),
    .A2(_0547_),
    .Y(_0549_),
    .B1(_0543_));
 sg13g2_a22oi_1 _1397_ (.Y(_0550_),
    .B1(_0548_),
    .B2(_0549_),
    .A2(_0545_),
    .A1(_0543_));
 sg13g2_nor2_2 _1398_ (.A(net251),
    .B(_0550_),
    .Y(\genrow[4].gencol[3].genblk1.c.bufs[0].A ));
 sg13g2_a21oi_1 _1399_ (.A1(\cell_cfg[20][1] ),
    .A2(\genrow[4].gencol[1].genblk1.c.bufs[0].A ),
    .Y(_0551_),
    .B1(\cell_cfg[20][2] ));
 sg13g2_o21ai_1 _1400_ (.B1(_0334_),
    .Y(_0552_),
    .A1(\cell_cfg[20][1] ),
    .A2(\cell_cfg[20][0] ));
 sg13g2_a21oi_1 _1401_ (.A1(\cell_cfg[20][2] ),
    .A2(_0405_),
    .Y(_0553_),
    .B1(_0551_));
 sg13g2_nand3_1 _1402_ (.B(\cell_cfg[20][0] ),
    .C(_0409_),
    .A(\cell_cfg[20][1] ),
    .Y(_0554_));
 sg13g2_o21ai_1 _1403_ (.B1(_0554_),
    .Y(_0555_),
    .A1(\cell_cfg[20][1] ),
    .A2(\genrow[5].gencol[2].genblk1.c.bufs[0].A ));
 sg13g2_nand3_1 _1404_ (.B(\cell_cfg[20][1] ),
    .C(\genrow[4].gencol[3].genblk1.c.bufs[0].A ),
    .A(\cell_cfg[20][2] ),
    .Y(_0556_));
 sg13g2_a22oi_1 _1405_ (.Y(_0557_),
    .B1(_0556_),
    .B2(_0371_),
    .A2(_0555_),
    .A1(\cell_cfg[20][2] ));
 sg13g2_a22oi_1 _1406_ (.Y(_0558_),
    .B1(_0557_),
    .B2(_0334_),
    .A2(_0553_),
    .A1(_0552_));
 sg13g2_nor2_2 _1407_ (.A(net251),
    .B(_0558_),
    .Y(\genrow[4].gencol[2].genblk1.c.bufs[0].A ));
 sg13g2_or2_1 _1408_ (.X(_0559_),
    .B(\cell_cfg[19][2] ),
    .A(\cell_cfg[19][3] ));
 sg13g2_nor2b_1 _1409_ (.A(\genrow[4].gencol[2].genblk1.c.bufs[0].A ),
    .B_N(\cell_cfg[19][1] ),
    .Y(_0560_));
 sg13g2_nor3_1 _1410_ (.A(\cell_cfg[19][0] ),
    .B(\cell_cfg[19][3] ),
    .C(_0560_),
    .Y(_0561_));
 sg13g2_o21ai_1 _1411_ (.B1(_0561_),
    .Y(_0562_),
    .A1(\cell_cfg[19][1] ),
    .A2(\genrow[3].gencol[1].genblk1.c.bufs[0].A ));
 sg13g2_a21oi_1 _1412_ (.A1(\cell_cfg[19][1] ),
    .A2(\genrow[4].gencol[0].genblk1.c.bufs[0].A ),
    .Y(_0563_),
    .B1(\cell_cfg[19][2] ));
 sg13g2_a21o_1 _1413_ (.A2(_0404_),
    .A1(\cell_cfg[19][2] ),
    .B1(_0380_),
    .X(_0564_));
 sg13g2_o21ai_1 _1414_ (.B1(_0562_),
    .Y(_0565_),
    .A1(_0563_),
    .A2(_0564_));
 sg13g2_o21ai_1 _1415_ (.B1(\cell_cfg[19][2] ),
    .Y(_0566_),
    .A1(\cell_cfg[19][1] ),
    .A2(_0416_));
 sg13g2_a21oi_1 _1416_ (.A1(\cell_cfg[19][1] ),
    .A2(net173),
    .Y(_0567_),
    .B1(_0566_));
 sg13g2_nor2b_1 _1417_ (.A(_0567_),
    .B_N(\cell_cfg[19][0] ),
    .Y(_0568_));
 sg13g2_a22oi_1 _1418_ (.Y(_0569_),
    .B1(_0568_),
    .B2(_0380_),
    .A2(_0565_),
    .A1(_0559_));
 sg13g2_nor2_2 _1419_ (.A(net252),
    .B(_0569_),
    .Y(\genrow[4].gencol[1].genblk1.c.bufs[0].A ));
 sg13g2_nand2_1 _1420_ (.Y(_0570_),
    .A(\cell_cfg[18][3] ),
    .B(\genrow[3].gencol[0].genblk1.c.bufs[0].A ));
 sg13g2_nand2_1 _1421_ (.Y(_0571_),
    .A(\cell_cfg[18][1] ),
    .B(net198));
 sg13g2_nor2_1 _1422_ (.A(_0388_),
    .B(\cell_cfg[18][2] ),
    .Y(_0572_));
 sg13g2_a22oi_1 _1423_ (.Y(_0573_),
    .B1(_0571_),
    .B2(_0572_),
    .A2(_0570_),
    .A1(\cell_cfg[18][2] ));
 sg13g2_mux4_1 _1424_ (.S0(\cell_cfg[18][1] ),
    .A0(\genrow[3].gencol[0].genblk1.c.bufs[0].A ),
    .A1(\genrow[4].gencol[1].genblk1.c.bufs[0].A ),
    .A2(\genrow[5].gencol[0].genblk1.c.bufs[0].A ),
    .A3(_0429_),
    .S1(\cell_cfg[18][0] ),
    .X(_0574_));
 sg13g2_a21oi_1 _1425_ (.A1(_0388_),
    .A2(_0574_),
    .Y(_0575_),
    .B1(_0573_));
 sg13g2_nor2_1 _1426_ (.A(\cell_cfg[18][3] ),
    .B(\cell_cfg[18][2] ),
    .Y(_0576_));
 sg13g2_nor3_1 _1427_ (.A(\cell_cfg[18][0] ),
    .B(\cell_cfg[18][3] ),
    .C(\cell_cfg[18][2] ),
    .Y(_0577_));
 sg13g2_nor3_2 _1428_ (.A(net252),
    .B(_0575_),
    .C(_0577_),
    .Y(\genrow[4].gencol[0].genblk1.c.bufs[0].A ));
 sg13g2_nor2_1 _1429_ (.A(net346),
    .B(net374),
    .Y(_0578_));
 sg13g2_nor2b_1 _1430_ (.A(net211),
    .B_N(\cell_cfg[16][1] ),
    .Y(_0579_));
 sg13g2_nor3_1 _1431_ (.A(\cell_cfg[16][0] ),
    .B(\cell_cfg[16][3] ),
    .C(_0579_),
    .Y(_0580_));
 sg13g2_o21ai_1 _1432_ (.B1(_0580_),
    .Y(_0581_),
    .A1(\cell_cfg[16][1] ),
    .A2(\genrow[2].gencol[4].genblk1.c.bufs[0].A ));
 sg13g2_a21oi_1 _1433_ (.A1(\cell_cfg[16][1] ),
    .A2(\genrow[3].gencol[3].genblk1.c.bufs[0].A ),
    .Y(_0582_),
    .B1(\cell_cfg[16][2] ));
 sg13g2_o21ai_1 _1434_ (.B1(\cell_cfg[16][3] ),
    .Y(_0583_),
    .A1(_0384_),
    .A2(\genrow[2].gencol[4].genblk1.c.bufs[0].A ));
 sg13g2_o21ai_1 _1435_ (.B1(_0581_),
    .Y(_0584_),
    .A1(_0582_),
    .A2(_0583_));
 sg13g2_nand2b_1 _1436_ (.Y(_0585_),
    .B(_0584_),
    .A_N(_0578_));
 sg13g2_o21ai_1 _1437_ (.B1(\cell_cfg[16][2] ),
    .Y(_0586_),
    .A1(\cell_cfg[16][1] ),
    .A2(_0413_));
 sg13g2_a21oi_1 _1438_ (.A1(\cell_cfg[16][1] ),
    .A2(\genrow[3].gencol[0].genblk1.c.bufs[0].A ),
    .Y(_0587_),
    .B1(_0586_));
 sg13g2_nand3b_1 _1439_ (.B(\cell_cfg[16][0] ),
    .C(_0383_),
    .Y(_0588_),
    .A_N(_0587_));
 sg13g2_a21oi_2 _1440_ (.B1(net252),
    .Y(\genrow[3].gencol[4].genblk1.c.bufs[0].A ),
    .A2(_0588_),
    .A1(_0585_));
 sg13g2_a21oi_1 _1441_ (.A1(\cell_cfg[15][1] ),
    .A2(\genrow[3].gencol[2].genblk1.c.bufs[0].A ),
    .Y(_0589_),
    .B1(\cell_cfg[15][2] ));
 sg13g2_o21ai_1 _1442_ (.B1(_0358_),
    .Y(_0590_),
    .A1(\cell_cfg[15][1] ),
    .A2(\cell_cfg[15][0] ));
 sg13g2_a21oi_1 _1443_ (.A1(\cell_cfg[15][2] ),
    .A2(_0402_),
    .Y(_0591_),
    .B1(_0589_));
 sg13g2_nand3_1 _1444_ (.B(\cell_cfg[15][0] ),
    .C(_0403_),
    .A(\cell_cfg[15][1] ),
    .Y(_0592_));
 sg13g2_o21ai_1 _1445_ (.B1(_0592_),
    .Y(_0593_),
    .A1(\cell_cfg[15][1] ),
    .A2(\genrow[4].gencol[3].genblk1.c.bufs[0].A ));
 sg13g2_a21o_1 _1446_ (.A2(\genrow[3].gencol[4].genblk1.c.bufs[0].A ),
    .A1(\cell_cfg[15][2] ),
    .B1(\cell_cfg[15][0] ),
    .X(_0594_));
 sg13g2_a21oi_1 _1447_ (.A1(\cell_cfg[15][2] ),
    .A2(_0593_),
    .Y(_0595_),
    .B1(_0590_));
 sg13g2_a22oi_1 _1448_ (.Y(_0596_),
    .B1(_0594_),
    .B2(_0595_),
    .A2(_0591_),
    .A1(_0590_));
 sg13g2_nor2_2 _1449_ (.A(net253),
    .B(_0596_),
    .Y(\genrow[3].gencol[3].genblk1.c.bufs[0].A ));
 sg13g2_a21oi_1 _1450_ (.A1(\cell_cfg[14][1] ),
    .A2(\genrow[3].gencol[1].genblk1.c.bufs[0].A ),
    .Y(_0597_),
    .B1(\cell_cfg[14][2] ));
 sg13g2_o21ai_1 _1451_ (.B1(_0355_),
    .Y(_0598_),
    .A1(\cell_cfg[14][1] ),
    .A2(\cell_cfg[14][0] ));
 sg13g2_a21oi_1 _1452_ (.A1(\cell_cfg[14][2] ),
    .A2(_0401_),
    .Y(_0599_),
    .B1(_0597_));
 sg13g2_nand3_1 _1453_ (.B(\cell_cfg[14][0] ),
    .C(_0403_),
    .A(\cell_cfg[14][1] ),
    .Y(_0600_));
 sg13g2_o21ai_1 _1454_ (.B1(_0600_),
    .Y(_0601_),
    .A1(\cell_cfg[14][1] ),
    .A2(\genrow[4].gencol[2].genblk1.c.bufs[0].A ));
 sg13g2_nand3_1 _1455_ (.B(\cell_cfg[14][1] ),
    .C(\genrow[3].gencol[3].genblk1.c.bufs[0].A ),
    .A(\cell_cfg[14][2] ),
    .Y(_0602_));
 sg13g2_a22oi_1 _1456_ (.Y(_0603_),
    .B1(_0602_),
    .B2(_0370_),
    .A2(_0601_),
    .A1(\cell_cfg[14][2] ));
 sg13g2_a22oi_1 _1457_ (.Y(_0604_),
    .B1(_0603_),
    .B2(_0355_),
    .A2(_0599_),
    .A1(_0598_));
 sg13g2_nor2_2 _1458_ (.A(net253),
    .B(_0604_),
    .Y(\genrow[3].gencol[2].genblk1.c.bufs[0].A ));
 sg13g2_and2_1 _1459_ (.A(\cell_cfg[13][1] ),
    .B(\genrow[3].gencol[0].genblk1.c.bufs[0].A ),
    .X(_0605_));
 sg13g2_mux4_1 _1460_ (.S0(\cell_cfg[13][1] ),
    .A0(\genrow[2].gencol[1].genblk1.c.bufs[0].A ),
    .A1(\genrow[3].gencol[2].genblk1.c.bufs[0].A ),
    .A2(\genrow[4].gencol[1].genblk1.c.bufs[0].A ),
    .A3(_0429_),
    .S1(\cell_cfg[13][0] ),
    .X(_0606_));
 sg13g2_nor2_1 _1461_ (.A(\cell_cfg[13][3] ),
    .B(net396),
    .Y(_0607_));
 sg13g2_or2_1 _1462_ (.X(_0608_),
    .B(\cell_cfg[13][2] ),
    .A(\cell_cfg[13][3] ));
 sg13g2_mux4_1 _1463_ (.S0(\cell_cfg[13][3] ),
    .A0(\cell_cfg[13][0] ),
    .A1(_0605_),
    .A2(_0606_),
    .A3(\genrow[2].gencol[1].genblk1.c.bufs[0].A ),
    .S1(\cell_cfg[13][2] ),
    .X(_0609_));
 sg13g2_and2_2 _1464_ (.A(_0394_),
    .B(_0609_),
    .X(\genrow[3].gencol[1].genblk1.c.bufs[0].A ));
 sg13g2_nand3b_1 _1465_ (.B(\cell_cfg[12][0] ),
    .C(\cell_cfg[12][1] ),
    .Y(_0610_),
    .A_N(\genrow[6].gencol[3].genblk1.c.bufs[0].A ));
 sg13g2_o21ai_1 _1466_ (.B1(_0610_),
    .Y(_0611_),
    .A1(\cell_cfg[12][1] ),
    .A2(\genrow[4].gencol[0].genblk1.c.bufs[0].A ));
 sg13g2_o21ai_1 _1467_ (.B1(_0335_),
    .Y(_0612_),
    .A1(\cell_cfg[12][1] ),
    .A2(\cell_cfg[12][0] ));
 sg13g2_nand3_1 _1468_ (.B(\cell_cfg[12][1] ),
    .C(\genrow[3].gencol[1].genblk1.c.bufs[0].A ),
    .A(\cell_cfg[12][2] ),
    .Y(_0613_));
 sg13g2_a22oi_1 _1469_ (.Y(_0614_),
    .B1(_0613_),
    .B2(_0369_),
    .A2(_0611_),
    .A1(\cell_cfg[12][2] ));
 sg13g2_a21oi_1 _1470_ (.A1(\cell_cfg[12][1] ),
    .A2(\genrow[3].gencol[5].genblk1.c.bufs[0].A ),
    .Y(_0615_),
    .B1(\cell_cfg[12][2] ));
 sg13g2_a21oi_1 _1471_ (.A1(\cell_cfg[12][2] ),
    .A2(_0399_),
    .Y(_0616_),
    .B1(_0615_));
 sg13g2_a22oi_1 _1472_ (.Y(_0617_),
    .B1(_0616_),
    .B2(_0612_),
    .A2(_0614_),
    .A1(_0335_));
 sg13g2_nor2_2 _1473_ (.A(net253),
    .B(_0617_),
    .Y(\genrow[3].gencol[0].genblk1.c.bufs[0].A ));
 sg13g2_nor2_1 _1474_ (.A(net380),
    .B(net486),
    .Y(_0618_));
 sg13g2_nor2b_1 _1475_ (.A(\genrow[3].gencol[0].genblk1.c.bufs[0].A ),
    .B_N(\cell_cfg[17][1] ),
    .Y(_0619_));
 sg13g2_nor3_1 _1476_ (.A(\cell_cfg[17][0] ),
    .B(\cell_cfg[17][3] ),
    .C(_0619_),
    .Y(_0620_));
 sg13g2_o21ai_1 _1477_ (.B1(_0620_),
    .Y(_0621_),
    .A1(\cell_cfg[17][1] ),
    .A2(net171));
 sg13g2_a21oi_1 _1478_ (.A1(\cell_cfg[17][1] ),
    .A2(net221),
    .Y(_0622_),
    .B1(\cell_cfg[17][2] ));
 sg13g2_o21ai_1 _1479_ (.B1(\cell_cfg[17][3] ),
    .Y(_0623_),
    .A1(_0393_),
    .A2(net171));
 sg13g2_o21ai_1 _1480_ (.B1(_0621_),
    .Y(_0624_),
    .A1(_0622_),
    .A2(_0623_));
 sg13g2_nand2b_1 _1481_ (.Y(_0625_),
    .B(_0624_),
    .A_N(_0618_));
 sg13g2_a21oi_1 _1482_ (.A1(\cell_cfg[17][1] ),
    .A2(net213),
    .Y(_0626_),
    .B1(_0393_));
 sg13g2_o21ai_1 _1483_ (.B1(_0626_),
    .Y(_0627_),
    .A1(\cell_cfg[17][1] ),
    .A2(_0414_));
 sg13g2_nand3_1 _1484_ (.B(_0392_),
    .C(_0627_),
    .A(\cell_cfg[17][0] ),
    .Y(_0628_));
 sg13g2_a21oi_2 _1485_ (.B1(net251),
    .Y(\genrow[3].gencol[5].genblk1.c.bufs[0].A ),
    .A2(_0628_),
    .A1(_0625_));
 sg13g2_nand3_1 _1486_ (.B(\cell_cfg[10][0] ),
    .C(_0399_),
    .A(\cell_cfg[10][1] ),
    .Y(_0629_));
 sg13g2_o21ai_1 _1487_ (.B1(_0629_),
    .Y(_0630_),
    .A1(\cell_cfg[10][1] ),
    .A2(net221));
 sg13g2_o21ai_1 _1488_ (.B1(_0354_),
    .Y(_0631_),
    .A1(\cell_cfg[10][1] ),
    .A2(\cell_cfg[10][0] ));
 sg13g2_nand3_1 _1489_ (.B(\cell_cfg[10][1] ),
    .C(\genrow[2].gencol[5].genblk1.c.bufs[0].A ),
    .A(\cell_cfg[10][2] ),
    .Y(_0632_));
 sg13g2_a22oi_1 _1490_ (.Y(_0633_),
    .B1(_0632_),
    .B2(_0367_),
    .A2(_0630_),
    .A1(\cell_cfg[10][2] ));
 sg13g2_a21oi_1 _1491_ (.A1(\cell_cfg[10][1] ),
    .A2(\genrow[2].gencol[3].genblk1.c.bufs[0].A ),
    .Y(_0634_),
    .B1(\cell_cfg[10][2] ));
 sg13g2_a21oi_1 _1492_ (.A1(\cell_cfg[10][2] ),
    .A2(_0425_),
    .Y(_0635_),
    .B1(_0634_));
 sg13g2_a22oi_1 _1493_ (.Y(_0636_),
    .B1(_0635_),
    .B2(_0631_),
    .A2(_0633_),
    .A1(_0354_));
 sg13g2_nor2_2 _1494_ (.A(net254),
    .B(_0636_),
    .Y(\genrow[2].gencol[4].genblk1.c.bufs[0].A ));
 sg13g2_a21oi_1 _1495_ (.A1(\cell_cfg[9][1] ),
    .A2(\genrow[2].gencol[2].genblk1.c.bufs[0].A ),
    .Y(_0637_),
    .B1(\cell_cfg[9][2] ));
 sg13g2_o21ai_1 _1496_ (.B1(_0357_),
    .Y(_0638_),
    .A1(\cell_cfg[9][1] ),
    .A2(\cell_cfg[9][0] ));
 sg13g2_a21oi_1 _1497_ (.A1(\cell_cfg[9][2] ),
    .A2(_0424_),
    .Y(_0639_),
    .B1(_0637_));
 sg13g2_nand3_1 _1498_ (.B(\cell_cfg[9][0] ),
    .C(_0399_),
    .A(\cell_cfg[9][1] ),
    .Y(_0640_));
 sg13g2_o21ai_1 _1499_ (.B1(_0640_),
    .Y(_0641_),
    .A1(\cell_cfg[9][1] ),
    .A2(\genrow[3].gencol[3].genblk1.c.bufs[0].A ));
 sg13g2_a21o_1 _1500_ (.A2(\genrow[2].gencol[4].genblk1.c.bufs[0].A ),
    .A1(\cell_cfg[9][2] ),
    .B1(\cell_cfg[9][0] ),
    .X(_0642_));
 sg13g2_a21oi_1 _1501_ (.A1(\cell_cfg[9][2] ),
    .A2(_0641_),
    .Y(_0643_),
    .B1(_0638_));
 sg13g2_a22oi_1 _1502_ (.Y(_0644_),
    .B1(_0642_),
    .B2(_0643_),
    .A2(_0639_),
    .A1(_0638_));
 sg13g2_nor2_1 _1503_ (.A(net253),
    .B(_0644_),
    .Y(\genrow[2].gencol[3].genblk1.c.bufs[0].A ));
 sg13g2_nand3_1 _1504_ (.B(\cell_cfg[8][0] ),
    .C(_0399_),
    .A(\cell_cfg[8][1] ),
    .Y(_0645_));
 sg13g2_o21ai_1 _1505_ (.B1(_0645_),
    .Y(_0646_),
    .A1(\cell_cfg[8][1] ),
    .A2(\genrow[3].gencol[2].genblk1.c.bufs[0].A ));
 sg13g2_o21ai_1 _1506_ (.B1(_0361_),
    .Y(_0647_),
    .A1(\cell_cfg[8][1] ),
    .A2(\cell_cfg[8][0] ));
 sg13g2_nand3_1 _1507_ (.B(\cell_cfg[8][1] ),
    .C(\genrow[2].gencol[3].genblk1.c.bufs[0].A ),
    .A(\cell_cfg[8][2] ),
    .Y(_0648_));
 sg13g2_a22oi_1 _1508_ (.Y(_0649_),
    .B1(_0648_),
    .B2(_0366_),
    .A2(_0646_),
    .A1(\cell_cfg[8][2] ));
 sg13g2_a21oi_1 _1509_ (.A1(\cell_cfg[8][1] ),
    .A2(\genrow[2].gencol[1].genblk1.c.bufs[0].A ),
    .Y(_0650_),
    .B1(\cell_cfg[8][2] ));
 sg13g2_a21oi_1 _1510_ (.A1(\cell_cfg[8][2] ),
    .A2(_0423_),
    .Y(_0651_),
    .B1(_0650_));
 sg13g2_a22oi_1 _1511_ (.Y(_0652_),
    .B1(_0651_),
    .B2(_0647_),
    .A2(_0649_),
    .A1(_0361_));
 sg13g2_nor2_2 _1512_ (.A(net253),
    .B(_0652_),
    .Y(\genrow[2].gencol[2].genblk1.c.bufs[0].A ));
 sg13g2_or2_1 _1513_ (.X(_0653_),
    .B(\cell_cfg[7][2] ),
    .A(\cell_cfg[7][3] ));
 sg13g2_nor2b_1 _1514_ (.A(\genrow[2].gencol[2].genblk1.c.bufs[0].A ),
    .B_N(\cell_cfg[7][1] ),
    .Y(_0654_));
 sg13g2_nor3_1 _1515_ (.A(\cell_cfg[7][0] ),
    .B(\cell_cfg[7][3] ),
    .C(_0654_),
    .Y(_0655_));
 sg13g2_o21ai_1 _1516_ (.B1(_0655_),
    .Y(_0656_),
    .A1(\cell_cfg[7][1] ),
    .A2(\genrow[1].gencol[1].genblk1.c.bufs[0].A ));
 sg13g2_a21oi_1 _1517_ (.A1(\cell_cfg[7][1] ),
    .A2(\genrow[2].gencol[0].genblk1.c.bufs[0].A ),
    .Y(_0657_),
    .B1(\cell_cfg[7][2] ));
 sg13g2_a21o_1 _1518_ (.A2(_0422_),
    .A1(\cell_cfg[7][2] ),
    .B1(_0385_),
    .X(_0658_));
 sg13g2_o21ai_1 _1519_ (.B1(_0656_),
    .Y(_0659_),
    .A1(_0657_),
    .A2(_0658_));
 sg13g2_o21ai_1 _1520_ (.B1(\cell_cfg[7][2] ),
    .Y(_0660_),
    .A1(\cell_cfg[7][1] ),
    .A2(_0404_));
 sg13g2_a21oi_1 _1521_ (.A1(\cell_cfg[7][1] ),
    .A2(\genrow[6].gencol[3].genblk1.c.bufs[0].A ),
    .Y(_0661_),
    .B1(_0660_));
 sg13g2_nor2b_1 _1522_ (.A(_0661_),
    .B_N(\cell_cfg[7][0] ),
    .Y(_0662_));
 sg13g2_a22oi_1 _1523_ (.Y(_0663_),
    .B1(_0662_),
    .B2(_0385_),
    .A2(_0659_),
    .A1(_0653_));
 sg13g2_nor2_2 _1524_ (.A(net253),
    .B(_0663_),
    .Y(\genrow[2].gencol[1].genblk1.c.bufs[0].A ));
 sg13g2_nor2_1 _1525_ (.A(net376),
    .B(net401),
    .Y(_0664_));
 sg13g2_a21oi_1 _1526_ (.A1(_0365_),
    .A2(_0421_),
    .Y(_0665_),
    .B1(\cell_cfg[6][0] ));
 sg13g2_a21oi_1 _1527_ (.A1(\cell_cfg[6][1] ),
    .A2(_0400_),
    .Y(_0666_),
    .B1(\cell_cfg[6][3] ));
 sg13g2_a21oi_1 _1528_ (.A1(\cell_cfg[6][1] ),
    .A2(net171),
    .Y(_0667_),
    .B1(\cell_cfg[6][2] ));
 sg13g2_a21oi_1 _1529_ (.A1(\cell_cfg[6][2] ),
    .A2(_0421_),
    .Y(_0668_),
    .B1(_0667_));
 sg13g2_a22oi_1 _1530_ (.Y(_0669_),
    .B1(_0668_),
    .B2(\cell_cfg[6][3] ),
    .A2(_0666_),
    .A1(_0665_));
 sg13g2_a21oi_1 _1531_ (.A1(\cell_cfg[6][1] ),
    .A2(net213),
    .Y(_0670_),
    .B1(_0387_));
 sg13g2_o21ai_1 _1532_ (.B1(_0670_),
    .Y(_0671_),
    .A1(\cell_cfg[6][1] ),
    .A2(_0403_));
 sg13g2_nand3_1 _1533_ (.B(_0386_),
    .C(_0671_),
    .A(\cell_cfg[6][0] ),
    .Y(_0672_));
 sg13g2_o21ai_1 _1534_ (.B1(_0672_),
    .Y(_0673_),
    .A1(_0664_),
    .A2(_0669_));
 sg13g2_and2_2 _1535_ (.A(_0394_),
    .B(_0673_),
    .X(\genrow[2].gencol[0].genblk1.c.bufs[0].A ));
 sg13g2_o21ai_1 _1536_ (.B1(\cell_cfg[5][1] ),
    .Y(_0674_),
    .A1(\cell_cfg[5][0] ),
    .A2(\genrow[1].gencol[0].genblk1.c.bufs[0].A ));
 sg13g2_a21oi_1 _1537_ (.A1(\cell_cfg[5][0] ),
    .A2(_0397_),
    .Y(_0675_),
    .B1(_0674_));
 sg13g2_nor2b_1 _1538_ (.A(net171),
    .B_N(\cell_cfg[5][0] ),
    .Y(_0676_));
 sg13g2_nor2_1 _1539_ (.A(net317),
    .B(\cell_cfg[5][0] ),
    .Y(_0677_));
 sg13g2_nor3_1 _1540_ (.A(\cell_cfg[5][1] ),
    .B(_0676_),
    .C(_0677_),
    .Y(_0678_));
 sg13g2_nor4_1 _1541_ (.A(\cell_cfg[5][3] ),
    .B(_0391_),
    .C(_0675_),
    .D(_0678_),
    .Y(_0679_));
 sg13g2_o21ai_1 _1542_ (.B1(\cell_cfg[5][1] ),
    .Y(_0680_),
    .A1(_0391_),
    .A2(net1));
 sg13g2_a21oi_1 _1543_ (.A1(_0391_),
    .A2(_0425_),
    .Y(_0681_),
    .B1(_0680_));
 sg13g2_nand2b_1 _1544_ (.Y(_0682_),
    .B(net317),
    .A_N(\cell_cfg[5][1] ));
 sg13g2_o21ai_1 _1545_ (.B1(\cell_cfg[5][3] ),
    .Y(_0683_),
    .A1(_0391_),
    .A2(_0682_));
 sg13g2_nor2_1 _1546_ (.A(net355),
    .B(net405),
    .Y(_0684_));
 sg13g2_a21oi_1 _1547_ (.A1(_0000_),
    .A2(_0684_),
    .Y(_0685_),
    .B1(net254));
 sg13g2_o21ai_1 _1548_ (.B1(_0685_),
    .Y(_0686_),
    .A1(_0681_),
    .A2(_0683_));
 sg13g2_nor2_2 _1549_ (.A(_0679_),
    .B(_0686_),
    .Y(_0687_));
 sg13g2_mux4_1 _1550_ (.S0(_0368_),
    .A0(\genrow[3].gencol[5].genblk1.c.bufs[0].A ),
    .A1(_0687_),
    .A2(\genrow[6].gencol[1].genblk1.c.bufs[0].A ),
    .A3(\genrow[2].gencol[0].genblk1.c.bufs[0].A ),
    .S1(\cell_cfg[11][1] ),
    .X(_0688_));
 sg13g2_nand3_1 _1551_ (.B(\cell_cfg[11][2] ),
    .C(_0687_),
    .A(\cell_cfg[11][3] ),
    .Y(_0689_));
 sg13g2_a21o_1 _1552_ (.A2(\genrow[2].gencol[4].genblk1.c.bufs[0].A ),
    .A1(\cell_cfg[11][1] ),
    .B1(_0345_),
    .X(_0690_));
 sg13g2_a22oi_1 _1553_ (.Y(_0691_),
    .B1(_0690_),
    .B2(_0346_),
    .A2(_0688_),
    .A1(_0345_));
 sg13g2_nor2_1 _1554_ (.A(\cell_cfg[11][3] ),
    .B(\cell_cfg[11][2] ),
    .Y(_0692_));
 sg13g2_a221oi_1 _1555_ (.B2(_0368_),
    .C1(net253),
    .B1(_0692_),
    .A1(_0691_),
    .Y(\genrow[2].gencol[5].genblk1.c.bufs[0].A ),
    .A2(_0689_));
 sg13g2_mux2_1 _1556_ (.A0(net318),
    .A1(_0687_),
    .S(\cell_cfg[4][1] ),
    .X(_0693_));
 sg13g2_nand2_1 _1557_ (.Y(_0694_),
    .A(\cell_cfg[4][1] ),
    .B(_0421_));
 sg13g2_o21ai_1 _1558_ (.B1(_0694_),
    .Y(_0695_),
    .A1(\cell_cfg[4][1] ),
    .A2(\genrow[2].gencol[4].genblk1.c.bufs[0].A ));
 sg13g2_a21oi_1 _1559_ (.A1(\cell_cfg[4][0] ),
    .A2(_0695_),
    .Y(_0696_),
    .B1(net482));
 sg13g2_o21ai_1 _1560_ (.B1(_0696_),
    .Y(_0697_),
    .A1(\cell_cfg[4][0] ),
    .A2(_0693_));
 sg13g2_nor2_1 _1561_ (.A(net382),
    .B(net388),
    .Y(_0698_));
 sg13g2_nand3b_1 _1562_ (.B(\cell_cfg[4][2] ),
    .C(\cell_cfg[4][1] ),
    .Y(_0699_),
    .A_N(net1));
 sg13g2_a21oi_1 _1563_ (.A1(net317),
    .A2(\cell_cfg[4][2] ),
    .Y(_0700_),
    .B1(\cell_cfg[4][1] ));
 sg13g2_nor2_1 _1564_ (.A(\cell_cfg[4][2] ),
    .B(\genrow[1].gencol[3].genblk1.c.bufs[0].A ),
    .Y(_0701_));
 sg13g2_nor3_1 _1565_ (.A(_0381_),
    .B(_0700_),
    .C(_0701_),
    .Y(_0702_));
 sg13g2_a21oi_1 _1566_ (.A1(_0699_),
    .A2(_0702_),
    .Y(_0703_),
    .B1(_0698_));
 sg13g2_a221oi_1 _1567_ (.B2(_0697_),
    .C1(net254),
    .B1(_0703_),
    .A1(_0364_),
    .Y(\genrow[1].gencol[4].genblk1.c.bufs[0].A ),
    .A2(_0698_));
 sg13g2_nand2_1 _1568_ (.Y(_0704_),
    .A(_0342_),
    .B(\cell_cfg[3][0] ));
 sg13g2_o21ai_1 _1569_ (.B1(\cell_cfg[3][1] ),
    .Y(_0705_),
    .A1(\cell_cfg[3][3] ),
    .A2(_0425_));
 sg13g2_a21oi_1 _1570_ (.A1(\cell_cfg[3][3] ),
    .A2(net1),
    .Y(_0706_),
    .B1(_0705_));
 sg13g2_o21ai_1 _1571_ (.B1(_0704_),
    .Y(_0707_),
    .A1(net317),
    .A2(\cell_cfg[3][1] ));
 sg13g2_or3_1 _1572_ (.A(_0343_),
    .B(_0706_),
    .C(_0707_),
    .X(_0708_));
 sg13g2_nand4_1 _1573_ (.B(_0343_),
    .C(\cell_cfg[3][1] ),
    .A(\cell_cfg[3][3] ),
    .Y(_0709_),
    .D(\genrow[1].gencol[2].genblk1.c.bufs[0].A ));
 sg13g2_mux2_1 _1574_ (.A0(_0402_),
    .A1(_0421_),
    .S(\cell_cfg[3][1] ),
    .X(_0710_));
 sg13g2_a22oi_1 _1575_ (.Y(_0711_),
    .B1(_0710_),
    .B2(\cell_cfg[3][2] ),
    .A2(_0709_),
    .A1(_0704_));
 sg13g2_inv_1 _1576_ (.Y(_0712_),
    .A(_0711_));
 sg13g2_a21oi_1 _1577_ (.A1(_0708_),
    .A2(_0712_),
    .Y(\genrow[1].gencol[3].genblk1.c.bufs[0].A ),
    .B1(net254));
 sg13g2_nand2b_1 _1578_ (.Y(_0713_),
    .B(\cell_cfg[2][0] ),
    .A_N(\cell_cfg[2][3] ));
 sg13g2_o21ai_1 _1579_ (.B1(\cell_cfg[2][1] ),
    .Y(_0714_),
    .A1(\cell_cfg[2][3] ),
    .A2(_0424_));
 sg13g2_a21oi_1 _1580_ (.A1(\cell_cfg[2][3] ),
    .A2(net1),
    .Y(_0715_),
    .B1(_0714_));
 sg13g2_nor2_1 _1581_ (.A(net317),
    .B(\cell_cfg[2][1] ),
    .Y(_0716_));
 sg13g2_nand2_1 _1582_ (.Y(_0717_),
    .A(\cell_cfg[2][2] ),
    .B(_0713_));
 sg13g2_nor3_1 _1583_ (.A(_0715_),
    .B(_0716_),
    .C(_0717_),
    .Y(_0718_));
 sg13g2_nand4_1 _1584_ (.B(_0353_),
    .C(\cell_cfg[2][1] ),
    .A(\cell_cfg[2][3] ),
    .Y(_0719_),
    .D(\genrow[1].gencol[1].genblk1.c.bufs[0].A ));
 sg13g2_mux2_1 _1585_ (.A0(_0401_),
    .A1(_0421_),
    .S(\cell_cfg[2][1] ),
    .X(_0720_));
 sg13g2_a22oi_1 _1586_ (.Y(_0721_),
    .B1(_0720_),
    .B2(\cell_cfg[2][2] ),
    .A2(_0719_),
    .A1(_0713_));
 sg13g2_nor2_1 _1587_ (.A(_0718_),
    .B(_0721_),
    .Y(_0722_));
 sg13g2_nor2_1 _1588_ (.A(net254),
    .B(_0722_),
    .Y(\genrow[1].gencol[2].genblk1.c.bufs[0].A ));
 sg13g2_nand2b_1 _1589_ (.Y(_0723_),
    .B(\cell_cfg[1][0] ),
    .A_N(\cell_cfg[1][3] ));
 sg13g2_o21ai_1 _1590_ (.B1(\cell_cfg[1][1] ),
    .Y(_0724_),
    .A1(\cell_cfg[1][3] ),
    .A2(_0423_));
 sg13g2_a21oi_1 _1591_ (.A1(\cell_cfg[1][3] ),
    .A2(net1),
    .Y(_0725_),
    .B1(_0724_));
 sg13g2_nor2_1 _1592_ (.A(net317),
    .B(\cell_cfg[1][1] ),
    .Y(_0726_));
 sg13g2_nand2_1 _1593_ (.Y(_0727_),
    .A(\cell_cfg[1][2] ),
    .B(_0723_));
 sg13g2_nor3_1 _1594_ (.A(_0725_),
    .B(_0726_),
    .C(_0727_),
    .Y(_0728_));
 sg13g2_nand4_1 _1595_ (.B(_0356_),
    .C(\cell_cfg[1][1] ),
    .A(\cell_cfg[1][3] ),
    .Y(_0729_),
    .D(\genrow[1].gencol[0].genblk1.c.bufs[0].A ));
 sg13g2_o21ai_1 _1596_ (.B1(\cell_cfg[1][2] ),
    .Y(_0730_),
    .A1(\cell_cfg[1][1] ),
    .A2(_0400_));
 sg13g2_a21oi_1 _1597_ (.A1(\cell_cfg[1][1] ),
    .A2(net215),
    .Y(_0731_),
    .B1(_0730_));
 sg13g2_a21oi_1 _1598_ (.A1(_0723_),
    .A2(_0729_),
    .Y(_0732_),
    .B1(_0731_));
 sg13g2_nor2_1 _1599_ (.A(_0728_),
    .B(_0732_),
    .Y(_0733_));
 sg13g2_nor2_2 _1600_ (.A(net254),
    .B(_0733_),
    .Y(\genrow[1].gencol[1].genblk1.c.bufs[0].A ));
 sg13g2_nor2_1 _1601_ (.A(\cell_cfg[0][3] ),
    .B(net429),
    .Y(_0734_));
 sg13g2_nor3_1 _1602_ (.A(\cell_cfg[0][3] ),
    .B(\cell_cfg[0][2] ),
    .C(\cell_cfg[0][0] ),
    .Y(_0735_));
 sg13g2_mux4_1 _1603_ (.S0(\cell_cfg[0][0] ),
    .A0(net317),
    .A1(\genrow[2].gencol[0].genblk1.c.bufs[0].A ),
    .A2(\genrow[1].gencol[1].genblk1.c.bufs[0].A ),
    .A3(\genrow[6].gencol[1].genblk1.c.bufs[0].A ),
    .S1(\cell_cfg[0][1] ),
    .X(_0736_));
 sg13g2_nand2b_1 _1604_ (.Y(_0737_),
    .B(\cell_cfg[0][3] ),
    .A_N(\cell_cfg[0][2] ));
 sg13g2_a21oi_1 _1605_ (.A1(\cell_cfg[0][1] ),
    .A2(_0687_),
    .Y(_0738_),
    .B1(_0737_));
 sg13g2_a21oi_1 _1606_ (.A1(\cell_cfg[0][1] ),
    .A2(net1),
    .Y(_0739_),
    .B1(_0360_));
 sg13g2_o21ai_1 _1607_ (.B1(_0739_),
    .Y(_0740_),
    .A1(_0362_),
    .A2(\cell_cfg[0][1] ));
 sg13g2_o21ai_1 _1608_ (.B1(_0740_),
    .Y(_0741_),
    .A1(\cell_cfg[0][3] ),
    .A2(_0736_));
 sg13g2_and2_1 _1609_ (.A(\cell_cfg[0][2] ),
    .B(_0741_),
    .X(_0742_));
 sg13g2_nor4_2 _1610_ (.A(net254),
    .B(_0735_),
    .C(_0742_),
    .Y(\genrow[1].gencol[0].genblk1.c.bufs[0].A ),
    .D(_0738_));
 sg13g2_nor2b_2 _1611_ (.A(net5),
    .B_N(net4),
    .Y(_0743_));
 sg13g2_nand2_1 _1612_ (.Y(_0744_),
    .A(\genrow[6].gencol[0].genblk1.c.bufs[0].A ),
    .B(_0743_));
 sg13g2_o21ai_1 _1613_ (.B1(_0744_),
    .Y(uo_out[4]),
    .A1(_0379_),
    .A2(_0743_));
 sg13g2_o21ai_1 _1614_ (.B1(_0744_),
    .Y(uo_out[5]),
    .A1(_0378_),
    .A2(_0743_));
 sg13g2_nand2_1 _1615_ (.Y(_0745_),
    .A(net172),
    .B(_0743_));
 sg13g2_o21ai_1 _1616_ (.B1(_0745_),
    .Y(uo_out[6]),
    .A1(_0352_),
    .A2(_0743_));
 sg13g2_o21ai_1 _1617_ (.B1(_0745_),
    .Y(uo_out[7]),
    .A1(_0351_),
    .A2(_0743_));
 sg13g2_nor2_2 _1618_ (.A(net4),
    .B(net5),
    .Y(_0746_));
 sg13g2_or2_1 _1619_ (.X(_0747_),
    .B(net5),
    .A(net4));
 sg13g2_o21ai_1 _1620_ (.B1(net320),
    .Y(_0748_),
    .A1(\cell_cfg[17][2] ),
    .A2(net278));
 sg13g2_a21oi_1 _1621_ (.A1(_0384_),
    .A2(net278),
    .Y(_0002_),
    .B1(_0748_));
 sg13g2_o21ai_1 _1622_ (.B1(net320),
    .Y(_0749_),
    .A1(net380),
    .A2(net278));
 sg13g2_a21oi_1 _1623_ (.A1(_0383_),
    .A2(net277),
    .Y(_0003_),
    .B1(_0749_));
 sg13g2_o21ai_1 _1624_ (.B1(net327),
    .Y(_0750_),
    .A1(net405),
    .A2(net301));
 sg13g2_a21oi_1 _1625_ (.A1(_0382_),
    .A2(net300),
    .Y(_0004_),
    .B1(_0750_));
 sg13g2_o21ai_1 _1626_ (.B1(net327),
    .Y(_0751_),
    .A1(net355),
    .A2(net300));
 sg13g2_a21oi_1 _1627_ (.A1(_0381_),
    .A2(net300),
    .Y(_0005_),
    .B1(_0751_));
 sg13g2_o21ai_1 _1628_ (.B1(net320),
    .Y(_0752_),
    .A1(net349),
    .A2(net281));
 sg13g2_a21oi_1 _1629_ (.A1(_0393_),
    .A2(net279),
    .Y(_0006_),
    .B1(_0752_));
 sg13g2_o21ai_1 _1630_ (.B1(net326),
    .Y(_0753_),
    .A1(\cell_cfg[18][3] ),
    .A2(net292));
 sg13g2_a21oi_1 _1631_ (.A1(_0392_),
    .A2(net292),
    .Y(_0007_),
    .B1(_0753_));
 sg13g2_o21ai_1 _1632_ (.B1(net328),
    .Y(_0754_),
    .A1(net401),
    .A2(net299));
 sg13g2_a21oi_1 _1633_ (.A1(_0391_),
    .A2(net299),
    .Y(_0008_),
    .B1(_0754_));
 sg13g2_o21ai_1 _1634_ (.B1(net328),
    .Y(_0755_),
    .A1(\cell_cfg[6][3] ),
    .A2(net299));
 sg13g2_a21oi_1 _1635_ (.A1(_0390_),
    .A2(net299),
    .Y(_0009_),
    .B1(_0755_));
 sg13g2_o21ai_1 _1636_ (.B1(net326),
    .Y(_0756_),
    .A1(net391),
    .A2(net291));
 sg13g2_a21oi_1 _1637_ (.A1(_0387_),
    .A2(net299),
    .Y(_0010_),
    .B1(_0756_));
 sg13g2_o21ai_1 _1638_ (.B1(net329),
    .Y(_0757_),
    .A1(\cell_cfg[7][3] ),
    .A2(net301));
 sg13g2_a21oi_1 _1639_ (.A1(_0386_),
    .A2(net301),
    .Y(_0011_),
    .B1(_0757_));
 sg13g2_o21ai_1 _1640_ (.B1(net320),
    .Y(_0758_),
    .A1(net374),
    .A2(net277));
 sg13g2_a21oi_1 _1641_ (.A1(_0359_),
    .A2(net277),
    .Y(_0012_),
    .B1(_0758_));
 sg13g2_o21ai_1 _1642_ (.B1(net320),
    .Y(_0759_),
    .A1(net346),
    .A2(net277));
 sg13g2_a21oi_1 _1643_ (.A1(_0358_),
    .A2(net277),
    .Y(_0013_),
    .B1(_0759_));
 sg13g2_o21ai_1 _1644_ (.B1(net327),
    .Y(_0760_),
    .A1(net388),
    .A2(net301));
 sg13g2_a21oi_1 _1645_ (.A1(_0343_),
    .A2(net300),
    .Y(_0014_),
    .B1(_0760_));
 sg13g2_o21ai_1 _1646_ (.B1(net327),
    .Y(_0761_),
    .A1(net382),
    .A2(net300));
 sg13g2_a21oi_1 _1647_ (.A1(_0342_),
    .A2(net300),
    .Y(_0015_),
    .B1(_0761_));
 sg13g2_o21ai_1 _1648_ (.B1(net320),
    .Y(_0762_),
    .A1(\cell_cfg[19][2] ),
    .A2(net281));
 sg13g2_a21oi_1 _1649_ (.A1(_0389_),
    .A2(net288),
    .Y(_0016_),
    .B1(_0762_));
 sg13g2_o21ai_1 _1650_ (.B1(net321),
    .Y(_0763_),
    .A1(net466),
    .A2(net279));
 sg13g2_a21oi_1 _1651_ (.A1(_0388_),
    .A2(net279),
    .Y(_0017_),
    .B1(_0763_));
 sg13g2_nand2_1 _1652_ (.Y(_0764_),
    .A(_0429_),
    .B(net263));
 sg13g2_nor3_1 _1653_ (.A(net353),
    .B(net344),
    .C(_0764_),
    .Y(_0765_));
 sg13g2_nand2_1 _1654_ (.Y(_0766_),
    .A(net344),
    .B(net261));
 sg13g2_nand2_1 _1655_ (.Y(_0767_),
    .A(net353),
    .B(net263));
 sg13g2_nor2_1 _1656_ (.A(_0470_),
    .B(net286),
    .Y(_0768_));
 sg13g2_a221oi_1 _1657_ (.B2(net369),
    .C1(_0765_),
    .B1(_0768_),
    .A1(\cell_cfg[34][0] ),
    .Y(_0769_),
    .A2(net286));
 sg13g2_nor2_1 _1658_ (.A(net310),
    .B(net370),
    .Y(_0018_));
 sg13g2_a21oi_1 _1659_ (.A1(\cell_cfg[34][1] ),
    .A2(net286),
    .Y(_0770_),
    .B1(_0768_));
 sg13g2_a221oi_1 _1660_ (.B2(_0764_),
    .C1(net309),
    .B1(_0770_),
    .A1(_0378_),
    .Y(_0019_),
    .A2(_0768_));
 sg13g2_nand2_1 _1661_ (.Y(_0771_),
    .A(net373),
    .B(net263));
 sg13g2_nand2_1 _1662_ (.Y(_0772_),
    .A(net357),
    .B(net261));
 sg13g2_o21ai_1 _1663_ (.B1(net263),
    .Y(_0773_),
    .A1(\cell_cfg[34][3] ),
    .A2(\cell_cfg[34][2] ));
 sg13g2_and2_1 _1664_ (.A(\genrow[6].gencol[3].genblk1.c.bufs[0].A ),
    .B(net262),
    .X(_0774_));
 sg13g2_a21oi_1 _1665_ (.A1(net443),
    .A2(net285),
    .Y(_0775_),
    .B1(_0774_));
 sg13g2_o21ai_1 _1666_ (.B1(net322),
    .Y(_0776_),
    .A1(net478),
    .A2(_0773_));
 sg13g2_a21oi_1 _1667_ (.A1(_0773_),
    .A2(_0775_),
    .Y(_0020_),
    .B1(_0776_));
 sg13g2_a21oi_1 _1668_ (.A1(net359),
    .A2(net285),
    .Y(_0777_),
    .B1(_0774_));
 sg13g2_o21ai_1 _1669_ (.B1(net322),
    .Y(_0778_),
    .A1(net490),
    .A2(_0773_));
 sg13g2_a21oi_1 _1670_ (.A1(_0773_),
    .A2(_0777_),
    .Y(_0021_),
    .B1(_0778_));
 sg13g2_nand2_1 _1671_ (.Y(_0779_),
    .A(net330),
    .B(net262));
 sg13g2_nand2_1 _1672_ (.Y(_0780_),
    .A(net336),
    .B(net272));
 sg13g2_nor2_1 _1673_ (.A(_0457_),
    .B(net285),
    .Y(_0781_));
 sg13g2_nand3_1 _1674_ (.B(_0457_),
    .C(net262),
    .A(\genrow[6].gencol[2].genblk1.c.bufs[0].A ),
    .Y(_0782_));
 sg13g2_a22oi_1 _1675_ (.Y(_0783_),
    .B1(_0781_),
    .B2(net443),
    .A2(net285),
    .A1(\cell_cfg[32][0] ));
 sg13g2_a21oi_1 _1676_ (.A1(_0782_),
    .A2(net444),
    .Y(_0022_),
    .B1(net309));
 sg13g2_o21ai_1 _1677_ (.B1(_0782_),
    .Y(_0784_),
    .A1(_0376_),
    .A2(net262));
 sg13g2_a21oi_1 _1678_ (.A1(net359),
    .A2(_0781_),
    .Y(_0785_),
    .B1(_0784_));
 sg13g2_nor2_1 _1679_ (.A(net309),
    .B(net360),
    .Y(_0023_));
 sg13g2_nand2_1 _1680_ (.Y(_0786_),
    .A(net233),
    .B(net272));
 sg13g2_nand2_1 _1681_ (.Y(_0787_),
    .A(net480),
    .B(net262));
 sg13g2_o21ai_1 _1682_ (.B1(net272),
    .Y(_0788_),
    .A1(\cell_cfg[32][3] ),
    .A2(\cell_cfg[32][2] ));
 sg13g2_o21ai_1 _1683_ (.B1(_0788_),
    .Y(_0789_),
    .A1(_0420_),
    .A2(net286));
 sg13g2_a21oi_1 _1684_ (.A1(net409),
    .A2(net285),
    .Y(_0790_),
    .B1(_0789_));
 sg13g2_o21ai_1 _1685_ (.B1(net328),
    .Y(_0791_),
    .A1(\cell_cfg[32][0] ),
    .A2(_0788_));
 sg13g2_nor2_1 _1686_ (.A(_0790_),
    .B(_0791_),
    .Y(_0024_));
 sg13g2_a21oi_1 _1687_ (.A1(net453),
    .A2(net298),
    .Y(_0792_),
    .B1(_0789_));
 sg13g2_o21ai_1 _1688_ (.B1(net328),
    .Y(_0793_),
    .A1(\cell_cfg[32][1] ),
    .A2(_0788_));
 sg13g2_nor2_1 _1689_ (.A(_0792_),
    .B(_0793_),
    .Y(_0025_));
 sg13g2_nand2_1 _1690_ (.Y(_0794_),
    .A(net332),
    .B(net262));
 sg13g2_nand2_1 _1691_ (.Y(_0795_),
    .A(net431),
    .B(net262));
 sg13g2_o21ai_1 _1692_ (.B1(net262),
    .Y(_0796_),
    .A1(net332),
    .A2(\cell_cfg[31][2] ));
 sg13g2_o21ai_1 _1693_ (.B1(_0796_),
    .Y(_0797_),
    .A1(_0397_),
    .A2(net287));
 sg13g2_a21oi_1 _1694_ (.A1(net386),
    .A2(net286),
    .Y(_0798_),
    .B1(_0797_));
 sg13g2_o21ai_1 _1695_ (.B1(net324),
    .Y(_0799_),
    .A1(\cell_cfg[31][0] ),
    .A2(_0796_));
 sg13g2_nor2_1 _1696_ (.A(_0798_),
    .B(_0799_),
    .Y(_0026_));
 sg13g2_a21oi_1 _1697_ (.A1(net498),
    .A2(net287),
    .Y(_0800_),
    .B1(_0797_));
 sg13g2_o21ai_1 _1698_ (.B1(net324),
    .Y(_0801_),
    .A1(net453),
    .A2(_0796_));
 sg13g2_nor2_1 _1699_ (.A(_0800_),
    .B(_0801_),
    .Y(_0027_));
 sg13g2_nand2_1 _1700_ (.Y(_0802_),
    .A(net351),
    .B(net261));
 sg13g2_nand2_1 _1701_ (.Y(_0803_),
    .A(net422),
    .B(net261));
 sg13g2_o21ai_1 _1702_ (.B1(net260),
    .Y(_0804_),
    .A1(\cell_cfg[30][3] ),
    .A2(\cell_cfg[30][2] ));
 sg13g2_o21ai_1 _1703_ (.B1(_0804_),
    .Y(_0805_),
    .A1(_0398_),
    .A2(net284));
 sg13g2_a21oi_1 _1704_ (.A1(net472),
    .A2(net284),
    .Y(_0806_),
    .B1(_0805_));
 sg13g2_o21ai_1 _1705_ (.B1(net323),
    .Y(_0807_),
    .A1(net386),
    .A2(_0804_));
 sg13g2_nor2_1 _1706_ (.A(_0806_),
    .B(_0807_),
    .Y(_0028_));
 sg13g2_a21oi_1 _1707_ (.A1(net510),
    .A2(net283),
    .Y(_0808_),
    .B1(_0805_));
 sg13g2_o21ai_1 _1708_ (.B1(net323),
    .Y(_0809_),
    .A1(net498),
    .A2(_0804_));
 sg13g2_nor2_1 _1709_ (.A(_0808_),
    .B(_0809_),
    .Y(_0029_));
 sg13g2_nand2_1 _1710_ (.Y(_0810_),
    .A(net464),
    .B(net261));
 sg13g2_nand2_1 _1711_ (.Y(_0811_),
    .A(net363),
    .B(net261));
 sg13g2_o21ai_1 _1712_ (.B1(net261),
    .Y(_0812_),
    .A1(\cell_cfg[29][3] ),
    .A2(\cell_cfg[29][2] ));
 sg13g2_o21ai_1 _1713_ (.B1(_0812_),
    .Y(_0813_),
    .A1(_0419_),
    .A2(net283));
 sg13g2_a21oi_1 _1714_ (.A1(net505),
    .A2(net283),
    .Y(_0814_),
    .B1(_0813_));
 sg13g2_o21ai_1 _1715_ (.B1(net323),
    .Y(_0815_),
    .A1(net472),
    .A2(_0812_));
 sg13g2_nor2_1 _1716_ (.A(_0814_),
    .B(_0815_),
    .Y(_0030_));
 sg13g2_a21oi_1 _1717_ (.A1(net508),
    .A2(net283),
    .Y(_0816_),
    .B1(_0813_));
 sg13g2_o21ai_1 _1718_ (.B1(net323),
    .Y(_0817_),
    .A1(\cell_cfg[29][1] ),
    .A2(_0812_));
 sg13g2_nor2_1 _1719_ (.A(_0816_),
    .B(_0817_),
    .Y(_0031_));
 sg13g2_nand2_1 _1720_ (.Y(_0818_),
    .A(net242),
    .B(net260));
 sg13g2_nand2_1 _1721_ (.Y(_0819_),
    .A(net427),
    .B(net260));
 sg13g2_o21ai_1 _1722_ (.B1(net260),
    .Y(_0820_),
    .A1(\cell_cfg[28][3] ),
    .A2(\cell_cfg[28][2] ));
 sg13g2_o21ai_1 _1723_ (.B1(_0820_),
    .Y(_0821_),
    .A1(_0418_),
    .A2(net282));
 sg13g2_a21oi_1 _1724_ (.A1(net347),
    .A2(net282),
    .Y(_0822_),
    .B1(_0821_));
 sg13g2_o21ai_1 _1725_ (.B1(net322),
    .Y(_0823_),
    .A1(\cell_cfg[28][0] ),
    .A2(_0820_));
 sg13g2_nor2_1 _1726_ (.A(_0822_),
    .B(_0823_),
    .Y(_0032_));
 sg13g2_a21oi_1 _1727_ (.A1(net473),
    .A2(net282),
    .Y(_0824_),
    .B1(_0821_));
 sg13g2_o21ai_1 _1728_ (.B1(net322),
    .Y(_0825_),
    .A1(\cell_cfg[28][1] ),
    .A2(_0820_));
 sg13g2_nor2_1 _1729_ (.A(_0824_),
    .B(_0825_),
    .Y(_0033_));
 sg13g2_nand2_1 _1730_ (.Y(_0826_),
    .A(net228),
    .B(net260));
 sg13g2_nand2_1 _1731_ (.Y(_0827_),
    .A(net423),
    .B(net260));
 sg13g2_o21ai_1 _1732_ (.B1(net260),
    .Y(_0828_),
    .A1(net516),
    .A2(\cell_cfg[27][2] ));
 sg13g2_o21ai_1 _1733_ (.B1(_0828_),
    .Y(_0829_),
    .A1(_0417_),
    .A2(net284));
 sg13g2_a21oi_1 _1734_ (.A1(net417),
    .A2(net282),
    .Y(_0830_),
    .B1(_0829_));
 sg13g2_o21ai_1 _1735_ (.B1(net322),
    .Y(_0831_),
    .A1(net347),
    .A2(_0828_));
 sg13g2_nor2_1 _1736_ (.A(_0830_),
    .B(_0831_),
    .Y(_0034_));
 sg13g2_a21oi_1 _1737_ (.A1(net497),
    .A2(net284),
    .Y(_0832_),
    .B1(_0829_));
 sg13g2_o21ai_1 _1738_ (.B1(net322),
    .Y(_0833_),
    .A1(net473),
    .A2(_0828_));
 sg13g2_nor2_1 _1739_ (.A(_0832_),
    .B(_0833_),
    .Y(_0035_));
 sg13g2_nand2_1 _1740_ (.Y(_0834_),
    .A(net337),
    .B(net257));
 sg13g2_nand2_1 _1741_ (.Y(_0835_),
    .A(net432),
    .B(net256));
 sg13g2_o21ai_1 _1742_ (.B1(net260),
    .Y(_0836_),
    .A1(\cell_cfg[26][3] ),
    .A2(\cell_cfg[26][2] ));
 sg13g2_o21ai_1 _1743_ (.B1(_0836_),
    .Y(_0837_),
    .A1(_0416_),
    .A2(net285));
 sg13g2_a21oi_1 _1744_ (.A1(net406),
    .A2(net285),
    .Y(_0838_),
    .B1(_0837_));
 sg13g2_o21ai_1 _1745_ (.B1(net322),
    .Y(_0839_),
    .A1(\cell_cfg[26][0] ),
    .A2(_0836_));
 sg13g2_nor2_1 _1746_ (.A(_0838_),
    .B(_0839_),
    .Y(_0036_));
 sg13g2_a21oi_1 _1747_ (.A1(net457),
    .A2(net285),
    .Y(_0840_),
    .B1(_0837_));
 sg13g2_o21ai_1 _1748_ (.B1(net322),
    .Y(_0841_),
    .A1(\cell_cfg[26][1] ),
    .A2(_0836_));
 sg13g2_nor2_1 _1749_ (.A(_0840_),
    .B(_0841_),
    .Y(_0037_));
 sg13g2_nand2_1 _1750_ (.Y(_0842_),
    .A(net341),
    .B(net256));
 sg13g2_nand2_1 _1751_ (.Y(_0843_),
    .A(net442),
    .B(net257));
 sg13g2_o21ai_1 _1752_ (.B1(net257),
    .Y(_0844_),
    .A1(\cell_cfg[25][3] ),
    .A2(\cell_cfg[25][2] ));
 sg13g2_o21ai_1 _1753_ (.B1(_0844_),
    .Y(_0845_),
    .A1(_0415_),
    .A2(net275));
 sg13g2_a21oi_1 _1754_ (.A1(net491),
    .A2(net275),
    .Y(_0846_),
    .B1(_0845_));
 sg13g2_o21ai_1 _1755_ (.B1(net321),
    .Y(_0847_),
    .A1(net406),
    .A2(_0844_));
 sg13g2_nor2_1 _1756_ (.A(_0846_),
    .B(_0847_),
    .Y(_0038_));
 sg13g2_a21oi_1 _1757_ (.A1(net398),
    .A2(net276),
    .Y(_0848_),
    .B1(_0845_));
 sg13g2_o21ai_1 _1758_ (.B1(net321),
    .Y(_0849_),
    .A1(\cell_cfg[25][1] ),
    .A2(_0844_));
 sg13g2_nor2_1 _1759_ (.A(_0848_),
    .B(_0849_),
    .Y(_0039_));
 sg13g2_nand2b_1 _1760_ (.Y(_0850_),
    .B(net256),
    .A_N(net200));
 sg13g2_o21ai_1 _1761_ (.B1(net256),
    .Y(_0851_),
    .A1(net468),
    .A2(\cell_cfg[24][2] ));
 sg13g2_inv_1 _1762_ (.Y(_0852_),
    .A(_0851_));
 sg13g2_a21oi_1 _1763_ (.A1(net511),
    .A2(net275),
    .Y(_0853_),
    .B1(_0852_));
 sg13g2_o21ai_1 _1764_ (.B1(net321),
    .Y(_0854_),
    .A1(net491),
    .A2(_0851_));
 sg13g2_a21oi_1 _1765_ (.A1(_0850_),
    .A2(_0853_),
    .Y(_0040_),
    .B1(_0854_));
 sg13g2_a21oi_1 _1766_ (.A1(net449),
    .A2(net275),
    .Y(_0855_),
    .B1(_0852_));
 sg13g2_a221oi_1 _1767_ (.B2(_0850_),
    .C1(net307),
    .B1(_0855_),
    .A1(_0372_),
    .Y(_0041_),
    .A2(_0852_));
 sg13g2_nand2_1 _1768_ (.Y(_0856_),
    .A(net241),
    .B(net258));
 sg13g2_nand2_1 _1769_ (.Y(_0857_),
    .A(net428),
    .B(net258));
 sg13g2_o21ai_1 _1770_ (.B1(net258),
    .Y(_0858_),
    .A1(\cell_cfg[23][3] ),
    .A2(\cell_cfg[23][2] ));
 sg13g2_o21ai_1 _1771_ (.B1(_0858_),
    .Y(_0859_),
    .A1(_0413_),
    .A2(net273));
 sg13g2_a21oi_1 _1772_ (.A1(net418),
    .A2(net273),
    .Y(_0860_),
    .B1(_0859_));
 sg13g2_o21ai_1 _1773_ (.B1(net319),
    .Y(_0861_),
    .A1(\cell_cfg[23][0] ),
    .A2(_0858_));
 sg13g2_nor2_1 _1774_ (.A(_0860_),
    .B(_0861_),
    .Y(_0042_));
 sg13g2_a21oi_1 _1775_ (.A1(net463),
    .A2(net273),
    .Y(_0862_),
    .B1(_0859_));
 sg13g2_o21ai_1 _1776_ (.B1(net319),
    .Y(_0863_),
    .A1(net449),
    .A2(_0858_));
 sg13g2_nor2_1 _1777_ (.A(_0862_),
    .B(_0863_),
    .Y(_0043_));
 sg13g2_nand2_1 _1778_ (.Y(_0864_),
    .A(net230),
    .B(net258));
 sg13g2_nand2_1 _1779_ (.Y(_0865_),
    .A(net414),
    .B(net258));
 sg13g2_o21ai_1 _1780_ (.B1(net258),
    .Y(_0866_),
    .A1(net230),
    .A2(\cell_cfg[22][2] ));
 sg13g2_o21ai_1 _1781_ (.B1(_0866_),
    .Y(_0867_),
    .A1(_0412_),
    .A2(net274));
 sg13g2_a21oi_1 _1782_ (.A1(net365),
    .A2(net274),
    .Y(_0868_),
    .B1(_0867_));
 sg13g2_o21ai_1 _1783_ (.B1(net319),
    .Y(_0869_),
    .A1(\cell_cfg[22][0] ),
    .A2(_0866_));
 sg13g2_nor2_1 _1784_ (.A(_0868_),
    .B(_0869_),
    .Y(_0044_));
 sg13g2_a21oi_1 _1785_ (.A1(net455),
    .A2(net274),
    .Y(_0870_),
    .B1(_0867_));
 sg13g2_o21ai_1 _1786_ (.B1(net319),
    .Y(_0871_),
    .A1(\cell_cfg[22][1] ),
    .A2(_0866_));
 sg13g2_nor2_1 _1787_ (.A(_0870_),
    .B(_0871_),
    .Y(_0045_));
 sg13g2_nand2_1 _1788_ (.Y(_0872_),
    .A(net237),
    .B(net258));
 sg13g2_nand2_1 _1789_ (.Y(_0873_),
    .A(net437),
    .B(net265));
 sg13g2_o21ai_1 _1790_ (.B1(net258),
    .Y(_0874_),
    .A1(net237),
    .A2(\cell_cfg[21][2] ));
 sg13g2_o21ai_1 _1791_ (.B1(_0874_),
    .Y(_0875_),
    .A1(_0411_),
    .A2(net273));
 sg13g2_a21oi_1 _1792_ (.A1(net436),
    .A2(net273),
    .Y(_0876_),
    .B1(_0875_));
 sg13g2_o21ai_1 _1793_ (.B1(net319),
    .Y(_0877_),
    .A1(net365),
    .A2(_0874_));
 sg13g2_nor2_1 _1794_ (.A(_0876_),
    .B(_0877_),
    .Y(_0046_));
 sg13g2_a21oi_1 _1795_ (.A1(net501),
    .A2(net273),
    .Y(_0878_),
    .B1(_0875_));
 sg13g2_o21ai_1 _1796_ (.B1(net319),
    .Y(_0879_),
    .A1(net455),
    .A2(_0874_));
 sg13g2_nor2_1 _1797_ (.A(_0878_),
    .B(_0879_),
    .Y(_0047_));
 sg13g2_nand2_1 _1798_ (.Y(_0880_),
    .A(net226),
    .B(net265));
 sg13g2_nand2_1 _1799_ (.Y(_0147_),
    .A(net378),
    .B(net259));
 sg13g2_o21ai_1 _1800_ (.B1(net259),
    .Y(_0148_),
    .A1(net226),
    .A2(\cell_cfg[20][2] ));
 sg13g2_o21ai_1 _1801_ (.B1(_0148_),
    .Y(_0149_),
    .A1(_0410_),
    .A2(net280));
 sg13g2_a21oi_1 _1802_ (.A1(net339),
    .A2(net280),
    .Y(_0150_),
    .B1(_0149_));
 sg13g2_o21ai_1 _1803_ (.B1(net320),
    .Y(_0151_),
    .A1(\cell_cfg[20][0] ),
    .A2(_0148_));
 sg13g2_nor2_1 _1804_ (.A(_0150_),
    .B(_0151_),
    .Y(_0048_));
 sg13g2_a21oi_1 _1805_ (.A1(net507),
    .A2(net280),
    .Y(_0152_),
    .B1(_0149_));
 sg13g2_o21ai_1 _1806_ (.B1(net320),
    .Y(_0153_),
    .A1(net501),
    .A2(_0148_));
 sg13g2_nor2_1 _1807_ (.A(_0152_),
    .B(_0153_),
    .Y(_0049_));
 sg13g2_and2_1 _1808_ (.A(_0559_),
    .B(net259),
    .X(_0154_));
 sg13g2_or3_1 _1809_ (.A(_0409_),
    .B(_0559_),
    .C(net280),
    .X(_0155_));
 sg13g2_a22oi_1 _1810_ (.Y(_0156_),
    .B1(_0154_),
    .B2(net339),
    .A2(net280),
    .A1(net371));
 sg13g2_a21oi_1 _1811_ (.A1(_0155_),
    .A2(_0156_),
    .Y(_0050_),
    .B1(net307));
 sg13g2_a22oi_1 _1812_ (.Y(_0157_),
    .B1(_0154_),
    .B2(\cell_cfg[19][1] ),
    .A2(net280),
    .A1(net484));
 sg13g2_a21oi_1 _1813_ (.A1(_0155_),
    .A2(net485),
    .Y(_0051_),
    .B1(net306));
 sg13g2_nor2_1 _1814_ (.A(_0576_),
    .B(net281),
    .Y(_0158_));
 sg13g2_and3_1 _1815_ (.X(_0159_),
    .A(net199),
    .B(_0576_),
    .C(net259));
 sg13g2_a221oi_1 _1816_ (.B2(net371),
    .C1(_0159_),
    .B1(_0158_),
    .A1(net411),
    .Y(_0160_),
    .A2(net279));
 sg13g2_nor2_1 _1817_ (.A(net306),
    .B(_0160_),
    .Y(_0052_));
 sg13g2_a221oi_1 _1818_ (.B2(net484),
    .C1(_0159_),
    .B1(_0158_),
    .A1(net499),
    .Y(_0161_),
    .A2(net279));
 sg13g2_nor2_1 _1819_ (.A(net306),
    .B(_0161_),
    .Y(_0053_));
 sg13g2_nor2_1 _1820_ (.A(_0618_),
    .B(net279),
    .Y(_0162_));
 sg13g2_nand3_1 _1821_ (.B(_0618_),
    .C(net259),
    .A(\genrow[3].gencol[4].genblk1.c.bufs[0].A ),
    .Y(_0163_));
 sg13g2_a22oi_1 _1822_ (.Y(_0164_),
    .B1(_0162_),
    .B2(net411),
    .A2(net279),
    .A1(\cell_cfg[16][0] ));
 sg13g2_a21oi_1 _1823_ (.A1(_0163_),
    .A2(net412),
    .Y(_0054_),
    .B1(net307));
 sg13g2_a22oi_1 _1824_ (.Y(_0165_),
    .B1(_0162_),
    .B2(net499),
    .A2(net279),
    .A1(\cell_cfg[16][1] ));
 sg13g2_a21oi_1 _1825_ (.A1(_0163_),
    .A2(net500),
    .Y(_0055_),
    .B1(net307));
 sg13g2_nor2_1 _1826_ (.A(_0578_),
    .B(net277),
    .Y(_0166_));
 sg13g2_nand3_1 _1827_ (.B(_0578_),
    .C(net259),
    .A(\genrow[3].gencol[3].genblk1.c.bufs[0].A ),
    .Y(_0167_));
 sg13g2_a22oi_1 _1828_ (.Y(_0168_),
    .B1(_0166_),
    .B2(net461),
    .A2(net277),
    .A1(\cell_cfg[15][0] ));
 sg13g2_a21oi_1 _1829_ (.A1(_0167_),
    .A2(net462),
    .Y(_0056_),
    .B1(net306));
 sg13g2_a22oi_1 _1830_ (.Y(_0169_),
    .B1(_0166_),
    .B2(net503),
    .A2(net277),
    .A1(\cell_cfg[15][1] ));
 sg13g2_a21oi_1 _1831_ (.A1(_0167_),
    .A2(net504),
    .Y(_0057_),
    .B1(net306));
 sg13g2_nand2_1 _1832_ (.Y(_0170_),
    .A(net223),
    .B(net266));
 sg13g2_nand2_1 _1833_ (.Y(_0171_),
    .A(net439),
    .B(net266));
 sg13g2_o21ai_1 _1834_ (.B1(net266),
    .Y(_0172_),
    .A1(net223),
    .A2(\cell_cfg[15][2] ));
 sg13g2_o21ai_1 _1835_ (.B1(_0172_),
    .Y(_0173_),
    .A1(_0405_),
    .A2(net290));
 sg13g2_a21oi_1 _1836_ (.A1(net404),
    .A2(net290),
    .Y(_0174_),
    .B1(_0173_));
 sg13g2_o21ai_1 _1837_ (.B1(net326),
    .Y(_0175_),
    .A1(net513),
    .A2(_0172_));
 sg13g2_nor2_1 _1838_ (.A(_0174_),
    .B(_0175_),
    .Y(_0058_));
 sg13g2_a21oi_1 _1839_ (.A1(net483),
    .A2(net290),
    .Y(_0176_),
    .B1(_0173_));
 sg13g2_o21ai_1 _1840_ (.B1(net326),
    .Y(_0177_),
    .A1(net514),
    .A2(_0172_));
 sg13g2_nor2_1 _1841_ (.A(_0176_),
    .B(_0177_),
    .Y(_0059_));
 sg13g2_nand2_1 _1842_ (.Y(_0178_),
    .A(net247),
    .B(net266));
 sg13g2_nand2_1 _1843_ (.Y(_0179_),
    .A(net421),
    .B(net266));
 sg13g2_o21ai_1 _1844_ (.B1(net266),
    .Y(_0180_),
    .A1(net517),
    .A2(\cell_cfg[14][2] ));
 sg13g2_o21ai_1 _1845_ (.B1(_0180_),
    .Y(_0181_),
    .A1(_0404_),
    .A2(net291));
 sg13g2_a21oi_1 _1846_ (.A1(net416),
    .A2(net291),
    .Y(_0182_),
    .B1(_0181_));
 sg13g2_o21ai_1 _1847_ (.B1(net326),
    .Y(_0183_),
    .A1(net404),
    .A2(_0180_));
 sg13g2_nor2_1 _1848_ (.A(_0182_),
    .B(_0183_),
    .Y(_0060_));
 sg13g2_a21oi_1 _1849_ (.A1(net408),
    .A2(net291),
    .Y(_0184_),
    .B1(_0181_));
 sg13g2_o21ai_1 _1850_ (.B1(net326),
    .Y(_0185_),
    .A1(net483),
    .A2(_0180_));
 sg13g2_nor2_1 _1851_ (.A(_0184_),
    .B(_0185_),
    .Y(_0061_));
 sg13g2_nand2_1 _1852_ (.Y(_0186_),
    .A(net396),
    .B(net266));
 sg13g2_nand2_1 _1853_ (.Y(_0187_),
    .A(\cell_cfg[13][3] ),
    .B(net266));
 sg13g2_nor2_1 _1854_ (.A(_0607_),
    .B(net291),
    .Y(_0188_));
 sg13g2_nand3_1 _1855_ (.B(_0607_),
    .C(net269),
    .A(\genrow[3].gencol[0].genblk1.c.bufs[0].A ),
    .Y(_0189_));
 sg13g2_a22oi_1 _1856_ (.Y(_0190_),
    .B1(_0188_),
    .B2(net416),
    .A2(net291),
    .A1(net425));
 sg13g2_a21oi_1 _1857_ (.A1(_0189_),
    .A2(_0190_),
    .Y(_0062_),
    .B1(net313));
 sg13g2_nand3_1 _1858_ (.B(_0608_),
    .C(net269),
    .A(net408),
    .Y(_0191_));
 sg13g2_nand2_1 _1859_ (.Y(_0192_),
    .A(_0189_),
    .B(_0191_));
 sg13g2_a21oi_1 _1860_ (.A1(net465),
    .A2(net291),
    .Y(_0193_),
    .B1(_0192_));
 sg13g2_nor2_1 _1861_ (.A(net311),
    .B(_0193_),
    .Y(_0063_));
 sg13g2_nand2_1 _1862_ (.Y(_0194_),
    .A(net243),
    .B(net267));
 sg13g2_nand2_1 _1863_ (.Y(_0195_),
    .A(\cell_cfg[12][2] ),
    .B(net267));
 sg13g2_o21ai_1 _1864_ (.B1(net267),
    .Y(_0196_),
    .A1(\cell_cfg[12][3] ),
    .A2(\cell_cfg[12][2] ));
 sg13g2_o21ai_1 _1865_ (.B1(_0196_),
    .Y(_0197_),
    .A1(_0408_),
    .A2(net293));
 sg13g2_a21oi_1 _1866_ (.A1(net239),
    .A2(net293),
    .Y(_0198_),
    .B1(_0197_));
 sg13g2_o21ai_1 _1867_ (.B1(net325),
    .Y(_0199_),
    .A1(\cell_cfg[12][0] ),
    .A2(_0196_));
 sg13g2_nor2_1 _1868_ (.A(_0198_),
    .B(_0199_),
    .Y(_0064_));
 sg13g2_a21oi_1 _1869_ (.A1(net394),
    .A2(net293),
    .Y(_0200_),
    .B1(_0197_));
 sg13g2_o21ai_1 _1870_ (.B1(net325),
    .Y(_0201_),
    .A1(\cell_cfg[12][1] ),
    .A2(_0196_));
 sg13g2_nor2_1 _1871_ (.A(_0200_),
    .B(_0201_),
    .Y(_0065_));
 sg13g2_a21oi_1 _1872_ (.A1(_0345_),
    .A2(_0346_),
    .Y(_0202_),
    .B1(net294));
 sg13g2_nand4_1 _1873_ (.B(_0346_),
    .C(_0345_),
    .A(\genrow[2].gencol[4].genblk1.c.bufs[0].A ),
    .Y(_0203_),
    .D(net268));
 sg13g2_a22oi_1 _1874_ (.Y(_0204_),
    .B1(_0202_),
    .B2(net239),
    .A2(net294),
    .A1(net358));
 sg13g2_a21oi_1 _1875_ (.A1(_0203_),
    .A2(_0204_),
    .Y(_0066_),
    .B1(net312));
 sg13g2_a22oi_1 _1876_ (.Y(_0205_),
    .B1(_0202_),
    .B2(net394),
    .A2(net293),
    .A1(net469));
 sg13g2_a21oi_1 _1877_ (.A1(_0203_),
    .A2(_0205_),
    .Y(_0067_),
    .B1(net312));
 sg13g2_nand2_1 _1878_ (.Y(_0206_),
    .A(net250),
    .B(net267));
 sg13g2_nand2_1 _1879_ (.Y(_0207_),
    .A(net445),
    .B(net269));
 sg13g2_o21ai_1 _1880_ (.B1(net267),
    .Y(_0208_),
    .A1(net448),
    .A2(\cell_cfg[10][2] ));
 sg13g2_o21ai_1 _1881_ (.B1(_0208_),
    .Y(_0209_),
    .A1(_0402_),
    .A2(net293));
 sg13g2_a21oi_1 _1882_ (.A1(net402),
    .A2(net294),
    .Y(_0210_),
    .B1(_0209_));
 sg13g2_o21ai_1 _1883_ (.B1(net325),
    .Y(_0211_),
    .A1(net358),
    .A2(_0208_));
 sg13g2_nor2_1 _1884_ (.A(_0210_),
    .B(_0211_),
    .Y(_0068_));
 sg13g2_a21oi_1 _1885_ (.A1(net481),
    .A2(net294),
    .Y(_0212_),
    .B1(_0209_));
 sg13g2_o21ai_1 _1886_ (.B1(net325),
    .Y(_0213_),
    .A1(net469),
    .A2(_0208_));
 sg13g2_nor2_1 _1887_ (.A(_0212_),
    .B(_0213_),
    .Y(_0069_));
 sg13g2_nand2_1 _1888_ (.Y(_0214_),
    .A(net238),
    .B(net268));
 sg13g2_nand2_1 _1889_ (.Y(_0215_),
    .A(net447),
    .B(net268));
 sg13g2_o21ai_1 _1890_ (.B1(net269),
    .Y(_0216_),
    .A1(net238),
    .A2(\cell_cfg[9][2] ));
 sg13g2_o21ai_1 _1891_ (.B1(_0216_),
    .Y(_0217_),
    .A1(_0401_),
    .A2(net296));
 sg13g2_a21oi_1 _1892_ (.A1(net400),
    .A2(net296),
    .Y(_0218_),
    .B1(_0217_));
 sg13g2_o21ai_1 _1893_ (.B1(net326),
    .Y(_0219_),
    .A1(net402),
    .A2(_0216_));
 sg13g2_nor2_1 _1894_ (.A(_0218_),
    .B(_0219_),
    .Y(_0070_));
 sg13g2_a21oi_1 _1895_ (.A1(net479),
    .A2(net295),
    .Y(_0220_),
    .B1(_0217_));
 sg13g2_o21ai_1 _1896_ (.B1(net329),
    .Y(_0221_),
    .A1(net481),
    .A2(_0216_));
 sg13g2_nor2_1 _1897_ (.A(_0220_),
    .B(_0221_),
    .Y(_0071_));
 sg13g2_nand2_1 _1898_ (.Y(_0222_),
    .A(net235),
    .B(net268));
 sg13g2_nand2_1 _1899_ (.Y(_0223_),
    .A(net420),
    .B(net268));
 sg13g2_o21ai_1 _1900_ (.B1(net268),
    .Y(_0224_),
    .A1(\cell_cfg[8][3] ),
    .A2(\cell_cfg[8][2] ));
 sg13g2_o21ai_1 _1901_ (.B1(_0224_),
    .Y(_0225_),
    .A1(_0400_),
    .A2(net295));
 sg13g2_a21oi_1 _1902_ (.A1(net361),
    .A2(net295),
    .Y(_0226_),
    .B1(_0225_));
 sg13g2_o21ai_1 _1903_ (.B1(net325),
    .Y(_0227_),
    .A1(\cell_cfg[8][0] ),
    .A2(_0224_));
 sg13g2_nor2_1 _1904_ (.A(_0226_),
    .B(_0227_),
    .Y(_0072_));
 sg13g2_a21oi_1 _1905_ (.A1(net492),
    .A2(net295),
    .Y(_0228_),
    .B1(_0225_));
 sg13g2_o21ai_1 _1906_ (.B1(net325),
    .Y(_0229_),
    .A1(net479),
    .A2(_0224_));
 sg13g2_nor2_1 _1907_ (.A(_0228_),
    .B(_0229_),
    .Y(_0073_));
 sg13g2_and2_1 _1908_ (.A(_0653_),
    .B(net269),
    .X(_0230_));
 sg13g2_or3_1 _1909_ (.A(_0399_),
    .B(_0653_),
    .C(net292),
    .X(_0231_));
 sg13g2_a22oi_1 _1910_ (.Y(_0232_),
    .B1(_0230_),
    .B2(net361),
    .A2(net291),
    .A1(net383));
 sg13g2_a21oi_1 _1911_ (.A1(_0231_),
    .A2(_0232_),
    .Y(_0074_),
    .B1(net311));
 sg13g2_a22oi_1 _1912_ (.Y(_0233_),
    .B1(_0230_),
    .B2(net492),
    .A2(net292),
    .A1(net502));
 sg13g2_a21oi_1 _1913_ (.A1(_0231_),
    .A2(_0233_),
    .Y(_0075_),
    .B1(net313));
 sg13g2_nor2_1 _1914_ (.A(_0664_),
    .B(net299),
    .Y(_0234_));
 sg13g2_nand3_1 _1915_ (.B(_0664_),
    .C(net272),
    .A(net171),
    .Y(_0235_));
 sg13g2_a22oi_1 _1916_ (.Y(_0236_),
    .B1(_0234_),
    .B2(net383),
    .A2(net299),
    .A1(\cell_cfg[5][0] ));
 sg13g2_a21oi_1 _1917_ (.A1(_0235_),
    .A2(net384),
    .Y(_0076_),
    .B1(net315));
 sg13g2_a22oi_1 _1918_ (.Y(_0237_),
    .B1(_0234_),
    .B2(net502),
    .A2(net299),
    .A1(net487));
 sg13g2_a21oi_1 _1919_ (.A1(_0235_),
    .A2(_0237_),
    .Y(_0077_),
    .B1(net315));
 sg13g2_nor2_1 _1920_ (.A(_0684_),
    .B(net301),
    .Y(_0238_));
 sg13g2_nand3_1 _1921_ (.B(_0684_),
    .C(net271),
    .A(\genrow[1].gencol[4].genblk1.c.bufs[0].A ),
    .Y(_0239_));
 sg13g2_a22oi_1 _1922_ (.Y(_0240_),
    .B1(_0238_),
    .B2(net450),
    .A2(net301),
    .A1(\cell_cfg[4][0] ));
 sg13g2_a21oi_1 _1923_ (.A1(_0239_),
    .A2(net451),
    .Y(_0078_),
    .B1(net314));
 sg13g2_a22oi_1 _1924_ (.Y(_0241_),
    .B1(_0238_),
    .B2(net487),
    .A2(net301),
    .A1(\cell_cfg[4][1] ));
 sg13g2_a21oi_1 _1925_ (.A1(_0239_),
    .A2(net488),
    .Y(_0079_),
    .B1(net314));
 sg13g2_nor2_1 _1926_ (.A(_0698_),
    .B(net300),
    .Y(_0242_));
 sg13g2_nand3_1 _1927_ (.B(_0698_),
    .C(net271),
    .A(\genrow[1].gencol[3].genblk1.c.bufs[0].A ),
    .Y(_0243_));
 sg13g2_a22oi_1 _1928_ (.Y(_0244_),
    .B1(_0242_),
    .B2(\cell_cfg[4][0] ),
    .A2(net300),
    .A1(net434));
 sg13g2_a21oi_1 _1929_ (.A1(_0243_),
    .A2(net435),
    .Y(_0080_),
    .B1(net314));
 sg13g2_o21ai_1 _1930_ (.B1(_0243_),
    .Y(_0245_),
    .A1(_0363_),
    .A2(net271));
 sg13g2_a21oi_1 _1931_ (.A1(net495),
    .A2(_0242_),
    .Y(_0246_),
    .B1(_0245_));
 sg13g2_nor2_1 _1932_ (.A(net314),
    .B(net496),
    .Y(_0081_));
 sg13g2_nand2_1 _1933_ (.Y(_0247_),
    .A(net392),
    .B(net271));
 sg13g2_nand2_1 _1934_ (.Y(_0248_),
    .A(net245),
    .B(net270));
 sg13g2_o21ai_1 _1935_ (.B1(net271),
    .Y(_0249_),
    .A1(\cell_cfg[3][3] ),
    .A2(net245));
 sg13g2_o21ai_1 _1936_ (.B1(_0249_),
    .Y(_0250_),
    .A1(_0423_),
    .A2(net302));
 sg13g2_a21oi_1 _1937_ (.A1(net232),
    .A2(net302),
    .Y(_0251_),
    .B1(_0250_));
 sg13g2_o21ai_1 _1938_ (.B1(net327),
    .Y(_0252_),
    .A1(net434),
    .A2(_0249_));
 sg13g2_nor2_1 _1939_ (.A(_0251_),
    .B(_0252_),
    .Y(_0082_));
 sg13g2_a21oi_1 _1940_ (.A1(net475),
    .A2(net302),
    .Y(_0253_),
    .B1(_0250_));
 sg13g2_o21ai_1 _1941_ (.B1(net327),
    .Y(_0254_),
    .A1(net515),
    .A2(_0249_));
 sg13g2_nor2_1 _1942_ (.A(_0253_),
    .B(_0254_),
    .Y(_0083_));
 sg13g2_nand2_1 _1943_ (.Y(_0255_),
    .A(net476),
    .B(net270));
 sg13g2_nand2_1 _1944_ (.Y(_0256_),
    .A(net372),
    .B(net270));
 sg13g2_o21ai_1 _1945_ (.B1(net270),
    .Y(_0257_),
    .A1(\cell_cfg[2][3] ),
    .A2(\cell_cfg[2][2] ));
 sg13g2_o21ai_1 _1946_ (.B1(_0257_),
    .Y(_0258_),
    .A1(_0422_),
    .A2(net303));
 sg13g2_a21oi_1 _1947_ (.A1(net343),
    .A2(net303),
    .Y(_0259_),
    .B1(_0258_));
 sg13g2_o21ai_1 _1948_ (.B1(net329),
    .Y(_0260_),
    .A1(net232),
    .A2(_0257_));
 sg13g2_nor2_1 _1949_ (.A(_0259_),
    .B(_0260_),
    .Y(_0084_));
 sg13g2_a21oi_1 _1950_ (.A1(net477),
    .A2(net303),
    .Y(_0261_),
    .B1(_0258_));
 sg13g2_o21ai_1 _1951_ (.B1(net329),
    .Y(_0262_),
    .A1(net475),
    .A2(_0257_));
 sg13g2_nor2_1 _1952_ (.A(_0261_),
    .B(_0262_),
    .Y(_0085_));
 sg13g2_nand2_1 _1953_ (.Y(_0263_),
    .A(net440),
    .B(net270));
 sg13g2_nand2_1 _1954_ (.Y(_0264_),
    .A(net367),
    .B(net270));
 sg13g2_o21ai_1 _1955_ (.B1(net270),
    .Y(_0265_),
    .A1(\cell_cfg[1][3] ),
    .A2(\cell_cfg[1][2] ));
 sg13g2_o21ai_1 _1956_ (.B1(_0265_),
    .Y(_0266_),
    .A1(_0421_),
    .A2(net304));
 sg13g2_a21oi_1 _1957_ (.A1(net389),
    .A2(net298),
    .Y(_0267_),
    .B1(_0266_));
 sg13g2_o21ai_1 _1958_ (.B1(net328),
    .Y(_0268_),
    .A1(net343),
    .A2(_0265_));
 sg13g2_nor2_1 _1959_ (.A(_0267_),
    .B(_0268_),
    .Y(_0086_));
 sg13g2_a21oi_1 _1960_ (.A1(net470),
    .A2(net298),
    .Y(_0269_),
    .B1(_0266_));
 sg13g2_o21ai_1 _1961_ (.B1(net328),
    .Y(_0270_),
    .A1(\cell_cfg[1][1] ),
    .A2(_0265_));
 sg13g2_nor2_1 _1962_ (.A(_0269_),
    .B(_0270_),
    .Y(_0087_));
 sg13g2_nor2_1 _1963_ (.A(net429),
    .B(net303),
    .Y(_0271_));
 sg13g2_nand3b_1 _1964_ (.B(_0687_),
    .C(_0271_),
    .Y(_0272_),
    .A_N(\cell_cfg[0][3] ));
 sg13g2_nor2_1 _1965_ (.A(_0734_),
    .B(net298),
    .Y(_0273_));
 sg13g2_a22oi_1 _1966_ (.Y(_0274_),
    .B1(_0273_),
    .B2(net389),
    .A2(net298),
    .A1(net317));
 sg13g2_a21oi_1 _1967_ (.A1(net430),
    .A2(_0274_),
    .Y(_0088_),
    .B1(net315));
 sg13g2_a22oi_1 _1968_ (.Y(_0275_),
    .B1(_0273_),
    .B2(net470),
    .A2(net298),
    .A1(net1));
 sg13g2_a21oi_1 _1969_ (.A1(net430),
    .A2(_0275_),
    .Y(_0089_),
    .B1(net315));
 sg13g2_nor2b_1 _1970_ (.A(net4),
    .B_N(net5),
    .Y(_0276_));
 sg13g2_o21ai_1 _1971_ (.B1(net328),
    .Y(_0277_),
    .A1(net225),
    .A2(_0276_));
 sg13g2_a21oi_1 _1972_ (.A1(_0362_),
    .A2(_0276_),
    .Y(_0090_),
    .B1(_0277_));
 sg13g2_nand2_1 _1973_ (.Y(_0278_),
    .A(net391),
    .B(net295));
 sg13g2_a21oi_1 _1974_ (.A1(_0223_),
    .A2(_0278_),
    .Y(_0091_),
    .B1(net312));
 sg13g2_nand2_1 _1975_ (.Y(_0279_),
    .A(\cell_cfg[7][3] ),
    .B(net295));
 sg13g2_a21oi_1 _1976_ (.A1(_0222_),
    .A2(_0279_),
    .Y(_0092_),
    .B1(net312));
 sg13g2_o21ai_1 _1977_ (.B1(net327),
    .Y(_0280_),
    .A1(net2),
    .A2(net270));
 sg13g2_nor2_1 _1978_ (.A(_0271_),
    .B(_0280_),
    .Y(_0093_));
 sg13g2_o21ai_1 _1979_ (.B1(net327),
    .Y(_0281_),
    .A1(net494),
    .A2(net302));
 sg13g2_a21oi_1 _1980_ (.A1(_0395_),
    .A2(net302),
    .Y(_0094_),
    .B1(_0281_));
 sg13g2_nand2_1 _1981_ (.Y(_0282_),
    .A(net421),
    .B(net290));
 sg13g2_a21oi_1 _1982_ (.A1(_0171_),
    .A2(_0282_),
    .Y(_0095_),
    .B1(net311));
 sg13g2_nand2_1 _1983_ (.Y(_0283_),
    .A(\cell_cfg[14][3] ),
    .B(net290));
 sg13g2_a21oi_1 _1984_ (.A1(_0170_),
    .A2(_0283_),
    .Y(_0096_),
    .B1(net311));
 sg13g2_nand2_1 _1985_ (.Y(_0284_),
    .A(net420),
    .B(net295));
 sg13g2_a21oi_1 _1986_ (.A1(_0215_),
    .A2(_0284_),
    .Y(_0097_),
    .B1(net312));
 sg13g2_nand2_1 _1987_ (.Y(_0285_),
    .A(net235),
    .B(net296));
 sg13g2_a21oi_1 _1988_ (.A1(_0214_),
    .A2(_0285_),
    .Y(_0098_),
    .B1(net313));
 sg13g2_nand2_1 _1989_ (.Y(_0286_),
    .A(\cell_cfg[0][2] ),
    .B(net303));
 sg13g2_a21oi_1 _1990_ (.A1(_0264_),
    .A2(_0286_),
    .Y(_0099_),
    .B1(net314));
 sg13g2_nand2_1 _1991_ (.Y(_0287_),
    .A(\cell_cfg[0][3] ),
    .B(net302));
 sg13g2_a21oi_1 _1992_ (.A1(_0263_),
    .A2(_0287_),
    .Y(_0100_),
    .B1(net314));
 sg13g2_nand2_1 _1993_ (.Y(_0288_),
    .A(net396),
    .B(net290));
 sg13g2_a21oi_1 _1994_ (.A1(_0179_),
    .A2(_0288_),
    .Y(_0101_),
    .B1(net311));
 sg13g2_nand2_1 _1995_ (.Y(_0289_),
    .A(\cell_cfg[13][3] ),
    .B(net297));
 sg13g2_a21oi_1 _1996_ (.A1(_0178_),
    .A2(_0289_),
    .Y(_0102_),
    .B1(net311));
 sg13g2_nand2_1 _1997_ (.Y(_0290_),
    .A(\cell_cfg[9][2] ),
    .B(net295));
 sg13g2_a21oi_1 _1998_ (.A1(_0207_),
    .A2(_0290_),
    .Y(_0103_),
    .B1(net313));
 sg13g2_nand2_1 _1999_ (.Y(_0291_),
    .A(net238),
    .B(net293));
 sg13g2_a21oi_1 _2000_ (.A1(_0206_),
    .A2(_0291_),
    .Y(_0104_),
    .B1(net312));
 sg13g2_nand2_1 _2001_ (.Y(_0292_),
    .A(net367),
    .B(net303));
 sg13g2_a21oi_1 _2002_ (.A1(_0256_),
    .A2(_0292_),
    .Y(_0105_),
    .B1(net314));
 sg13g2_nand2_1 _2003_ (.Y(_0293_),
    .A(net440),
    .B(net302));
 sg13g2_a21oi_1 _2004_ (.A1(_0255_),
    .A2(_0293_),
    .Y(_0106_),
    .B1(net314));
 sg13g2_nand2_1 _2005_ (.Y(_0294_),
    .A(\cell_cfg[34][2] ),
    .B(net284));
 sg13g2_a21oi_1 _2006_ (.A1(_0766_),
    .A2(_0294_),
    .Y(_0107_),
    .B1(net310));
 sg13g2_nand2_1 _2007_ (.Y(_0295_),
    .A(\cell_cfg[34][3] ),
    .B(net286));
 sg13g2_a21oi_1 _2008_ (.A1(_0767_),
    .A2(_0295_),
    .Y(_0108_),
    .B1(net309));
 sg13g2_nand2_1 _2009_ (.Y(_0296_),
    .A(\cell_cfg[12][2] ),
    .B(net290));
 sg13g2_a21oi_1 _2010_ (.A1(_0186_),
    .A2(_0296_),
    .Y(_0109_),
    .B1(net311));
 sg13g2_nand2_1 _2011_ (.Y(_0297_),
    .A(net243),
    .B(net290));
 sg13g2_a21oi_1 _2012_ (.A1(_0187_),
    .A2(_0297_),
    .Y(_0110_),
    .B1(net311));
 sg13g2_nand2_1 _2013_ (.Y(_0298_),
    .A(net330),
    .B(net286));
 sg13g2_a21oi_1 _2014_ (.A1(_0772_),
    .A2(_0298_),
    .Y(_0111_),
    .B1(net308));
 sg13g2_nand2_1 _2015_ (.Y(_0299_),
    .A(net336),
    .B(net286));
 sg13g2_a21oi_1 _2016_ (.A1(_0771_),
    .A2(_0299_),
    .Y(_0112_),
    .B1(net309));
 sg13g2_nand2_1 _2017_ (.Y(_0300_),
    .A(\cell_cfg[32][2] ),
    .B(net288));
 sg13g2_a21oi_1 _2018_ (.A1(_0779_),
    .A2(_0300_),
    .Y(_0113_),
    .B1(net309));
 sg13g2_nand2_1 _2019_ (.Y(_0301_),
    .A(net233),
    .B(net298));
 sg13g2_a21oi_1 _2020_ (.A1(_0780_),
    .A2(_0301_),
    .Y(_0114_),
    .B1(net315));
 sg13g2_nand2_1 _2021_ (.Y(_0302_),
    .A(net431),
    .B(net287));
 sg13g2_a21oi_1 _2022_ (.A1(_0787_),
    .A2(_0302_),
    .Y(_0115_),
    .B1(net315));
 sg13g2_nand2_1 _2023_ (.Y(_0303_),
    .A(\cell_cfg[31][3] ),
    .B(net298));
 sg13g2_a21oi_1 _2024_ (.A1(_0786_),
    .A2(_0303_),
    .Y(_0116_),
    .B1(net315));
 sg13g2_nand2_1 _2025_ (.Y(_0304_),
    .A(net422),
    .B(net287));
 sg13g2_a21oi_1 _2026_ (.A1(_0795_),
    .A2(_0304_),
    .Y(_0117_),
    .B1(net309));
 sg13g2_nand2_1 _2027_ (.Y(_0305_),
    .A(\cell_cfg[30][3] ),
    .B(net287));
 sg13g2_a21oi_1 _2028_ (.A1(_0794_),
    .A2(_0305_),
    .Y(_0118_),
    .B1(net309));
 sg13g2_nand2_1 _2029_ (.Y(_0306_),
    .A(net363),
    .B(net283));
 sg13g2_a21oi_1 _2030_ (.A1(_0803_),
    .A2(_0306_),
    .Y(_0119_),
    .B1(net308));
 sg13g2_nand2_1 _2031_ (.Y(_0307_),
    .A(\cell_cfg[29][3] ),
    .B(net283));
 sg13g2_a21oi_1 _2032_ (.A1(_0802_),
    .A2(_0307_),
    .Y(_0120_),
    .B1(net308));
 sg13g2_nand2_1 _2033_ (.Y(_0308_),
    .A(\cell_cfg[28][2] ),
    .B(net283));
 sg13g2_a21oi_1 _2034_ (.A1(_0811_),
    .A2(_0308_),
    .Y(_0121_),
    .B1(net310));
 sg13g2_nand2_1 _2035_ (.Y(_0309_),
    .A(net242),
    .B(net283));
 sg13g2_a21oi_1 _2036_ (.A1(_0810_),
    .A2(_0309_),
    .Y(_0122_),
    .B1(net310));
 sg13g2_nand2_1 _2037_ (.Y(_0310_),
    .A(net423),
    .B(net282));
 sg13g2_a21oi_1 _2038_ (.A1(_0819_),
    .A2(_0310_),
    .Y(_0123_),
    .B1(net308));
 sg13g2_nand2_1 _2039_ (.Y(_0311_),
    .A(net228),
    .B(net282));
 sg13g2_a21oi_1 _2040_ (.A1(_0818_),
    .A2(_0311_),
    .Y(_0124_),
    .B1(net308));
 sg13g2_nand2_1 _2041_ (.Y(_0312_),
    .A(\cell_cfg[26][2] ),
    .B(net282));
 sg13g2_a21oi_1 _2042_ (.A1(_0827_),
    .A2(_0312_),
    .Y(_0125_),
    .B1(net308));
 sg13g2_nand2_1 _2043_ (.Y(_0313_),
    .A(\cell_cfg[26][3] ),
    .B(net282));
 sg13g2_a21oi_1 _2044_ (.A1(_0826_),
    .A2(_0313_),
    .Y(_0126_),
    .B1(net308));
 sg13g2_o21ai_1 _2045_ (.B1(net325),
    .Y(_0314_),
    .A1(net445),
    .A2(net267));
 sg13g2_a21oi_1 _2046_ (.A1(_0346_),
    .A2(net267),
    .Y(_0127_),
    .B1(_0314_));
 sg13g2_o21ai_1 _2047_ (.B1(net325),
    .Y(_0315_),
    .A1(net250),
    .A2(net268));
 sg13g2_a21oi_1 _2048_ (.A1(_0345_),
    .A2(net267),
    .Y(_0128_),
    .B1(_0315_));
 sg13g2_nand2_1 _2049_ (.Y(_0316_),
    .A(\cell_cfg[25][2] ),
    .B(net275));
 sg13g2_a21oi_1 _2050_ (.A1(_0835_),
    .A2(_0316_),
    .Y(_0129_),
    .B1(net305));
 sg13g2_nand2_1 _2051_ (.Y(_0317_),
    .A(\cell_cfg[25][3] ),
    .B(net275));
 sg13g2_a21oi_1 _2052_ (.A1(_0834_),
    .A2(_0317_),
    .Y(_0130_),
    .B1(net308));
 sg13g2_nand2_1 _2053_ (.Y(_0318_),
    .A(\cell_cfg[2][2] ),
    .B(net303));
 sg13g2_a21oi_1 _2054_ (.A1(_0248_),
    .A2(_0318_),
    .Y(_0131_),
    .B1(net316));
 sg13g2_nand2_1 _2055_ (.Y(_0319_),
    .A(\cell_cfg[2][3] ),
    .B(net302));
 sg13g2_a21oi_1 _2056_ (.A1(_0247_),
    .A2(_0319_),
    .Y(_0132_),
    .B1(net316));
 sg13g2_nand2_1 _2057_ (.Y(_0320_),
    .A(net438),
    .B(net275));
 sg13g2_a21oi_1 _2058_ (.A1(_0843_),
    .A2(_0320_),
    .Y(_0133_),
    .B1(net305));
 sg13g2_nand2_1 _2059_ (.Y(_0321_),
    .A(\cell_cfg[24][3] ),
    .B(net275));
 sg13g2_a21oi_1 _2060_ (.A1(_0842_),
    .A2(_0321_),
    .Y(_0134_),
    .B1(net305));
 sg13g2_o21ai_1 _2061_ (.B1(net319),
    .Y(_0322_),
    .A1(net428),
    .A2(net256));
 sg13g2_a21oi_1 _2062_ (.A1(_0340_),
    .A2(net256),
    .Y(_0135_),
    .B1(_0322_));
 sg13g2_o21ai_1 _2063_ (.B1(net319),
    .Y(_0323_),
    .A1(net241),
    .A2(net256));
 sg13g2_a21oi_1 _2064_ (.A1(_0339_),
    .A2(net256),
    .Y(_0136_),
    .B1(_0323_));
 sg13g2_nand2_1 _2065_ (.Y(_0324_),
    .A(net414),
    .B(net273));
 sg13g2_a21oi_1 _2066_ (.A1(_0857_),
    .A2(_0324_),
    .Y(_0137_),
    .B1(net305));
 sg13g2_nand2_1 _2067_ (.Y(_0325_),
    .A(net230),
    .B(net273));
 sg13g2_a21oi_1 _2068_ (.A1(_0856_),
    .A2(_0325_),
    .Y(_0138_),
    .B1(net305));
 sg13g2_nand2_1 _2069_ (.Y(_0326_),
    .A(\cell_cfg[21][2] ),
    .B(net274));
 sg13g2_a21oi_1 _2070_ (.A1(_0865_),
    .A2(_0326_),
    .Y(_0139_),
    .B1(net305));
 sg13g2_nand2_1 _2071_ (.Y(_0327_),
    .A(\cell_cfg[21][3] ),
    .B(net274));
 sg13g2_a21oi_1 _2072_ (.A1(_0864_),
    .A2(_0327_),
    .Y(_0140_),
    .B1(net305));
 sg13g2_nand2_1 _2073_ (.Y(_0328_),
    .A(net378),
    .B(net278));
 sg13g2_a21oi_1 _2074_ (.A1(_0873_),
    .A2(_0328_),
    .Y(_0141_),
    .B1(net306));
 sg13g2_nand2_1 _2075_ (.Y(_0329_),
    .A(net226),
    .B(net278));
 sg13g2_a21oi_1 _2076_ (.A1(_0872_),
    .A2(_0329_),
    .Y(_0142_),
    .B1(net305));
 sg13g2_nand2_1 _2077_ (.Y(_0330_),
    .A(net334),
    .B(net293));
 sg13g2_a21oi_1 _2078_ (.A1(_0195_),
    .A2(_0330_),
    .Y(_0143_),
    .B1(net312));
 sg13g2_nand2_1 _2079_ (.Y(_0331_),
    .A(net249),
    .B(net293));
 sg13g2_a21oi_1 _2080_ (.A1(_0194_),
    .A2(_0331_),
    .Y(_0144_),
    .B1(net312));
 sg13g2_nand2_1 _2081_ (.Y(_0332_),
    .A(\cell_cfg[19][2] ),
    .B(net280));
 sg13g2_a21oi_1 _2082_ (.A1(_0147_),
    .A2(_0332_),
    .Y(_0145_),
    .B1(net306));
 sg13g2_nand2_1 _2083_ (.Y(_0333_),
    .A(\cell_cfg[19][3] ),
    .B(net278));
 sg13g2_a21oi_1 _2084_ (.A1(_0880_),
    .A2(_0333_),
    .Y(_0146_),
    .B1(net306));
 sg13g2_dfrbp_1 _2085_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net92),
    .D(net375),
    .Q_N(_1023_),
    .Q(\cell_cfg[17][2] ));
 sg13g2_dfrbp_1 _2086_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net125),
    .D(_0003_),
    .Q_N(_1022_),
    .Q(\cell_cfg[17][3] ));
 sg13g2_dfrbp_1 _2087_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net123),
    .D(_0004_),
    .Q_N(_1021_),
    .Q(\cell_cfg[5][2] ));
 sg13g2_dfrbp_1 _2088_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net121),
    .D(_0005_),
    .Q_N(_1020_),
    .Q(\cell_cfg[5][3] ));
 sg13g2_dfrbp_1 _2089_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net119),
    .D(_0006_),
    .Q_N(_1019_),
    .Q(\cell_cfg[18][2] ));
 sg13g2_dfrbp_1 _2090_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net117),
    .D(net381),
    .Q_N(_1018_),
    .Q(\cell_cfg[18][3] ));
 sg13g2_dfrbp_1 _2091_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net115),
    .D(_0008_),
    .Q_N(_1017_),
    .Q(\cell_cfg[6][2] ));
 sg13g2_dfrbp_1 _2092_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net113),
    .D(net356),
    .Q_N(_1016_),
    .Q(\cell_cfg[6][3] ));
 sg13g2_dfrbp_1 _2093_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net111),
    .D(_0010_),
    .Q_N(_1015_),
    .Q(\cell_cfg[7][2] ));
 sg13g2_dfrbp_1 _2094_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net109),
    .D(net377),
    .Q_N(_1014_),
    .Q(\cell_cfg[7][3] ));
 sg13g2_dfrbp_1 _2095_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net107),
    .D(_0012_),
    .Q_N(_1013_),
    .Q(\cell_cfg[16][2] ));
 sg13g2_dfrbp_1 _2096_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net105),
    .D(_0013_),
    .Q_N(_1012_),
    .Q(\cell_cfg[16][3] ));
 sg13g2_dfrbp_1 _2097_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net103),
    .D(_0014_),
    .Q_N(_1011_),
    .Q(\cell_cfg[4][2] ));
 sg13g2_dfrbp_1 _2098_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net101),
    .D(_0015_),
    .Q_N(_1010_),
    .Q(\cell_cfg[4][3] ));
 sg13g2_dfrbp_1 _2099_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net99),
    .D(net350),
    .Q_N(_1009_),
    .Q(\cell_cfg[19][2] ));
 sg13g2_dfrbp_1 _2100_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net97),
    .D(net467),
    .Q_N(_1008_),
    .Q(\cell_cfg[19][3] ));
 sg13g2_dfrbp_1 _2101_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net95),
    .D(_0018_),
    .Q_N(_1007_),
    .Q(\cell_cfg[35][0] ));
 sg13g2_dfrbp_1 _2102_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net93),
    .D(net460),
    .Q_N(_1006_),
    .Q(\cell_cfg[35][1] ));
 sg13g2_dfrbp_1 _2103_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net91),
    .D(_0020_),
    .Q_N(_1005_),
    .Q(\cell_cfg[34][0] ));
 sg13g2_dfrbp_1 _2104_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net89),
    .D(_0021_),
    .Q_N(_1004_),
    .Q(\cell_cfg[34][1] ));
 sg13g2_dfrbp_1 _2105_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net87),
    .D(_0022_),
    .Q_N(_1003_),
    .Q(\cell_cfg[33][0] ));
 sg13g2_dfrbp_1 _2106_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net85),
    .D(_0023_),
    .Q_N(_1002_),
    .Q(\cell_cfg[33][1] ));
 sg13g2_dfrbp_1 _2107_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net83),
    .D(net410),
    .Q_N(_1001_),
    .Q(\cell_cfg[32][0] ));
 sg13g2_dfrbp_1 _2108_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net81),
    .D(net454),
    .Q_N(_1000_),
    .Q(\cell_cfg[32][1] ));
 sg13g2_dfrbp_1 _2109_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net79),
    .D(net387),
    .Q_N(_0999_),
    .Q(\cell_cfg[31][0] ));
 sg13g2_dfrbp_1 _2110_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net77),
    .D(_0027_),
    .Q_N(_0998_),
    .Q(\cell_cfg[31][1] ));
 sg13g2_dfrbp_1 _2111_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net75),
    .D(_0028_),
    .Q_N(_0997_),
    .Q(\cell_cfg[30][0] ));
 sg13g2_dfrbp_1 _2112_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net73),
    .D(_0029_),
    .Q_N(_0996_),
    .Q(\cell_cfg[30][1] ));
 sg13g2_dfrbp_1 _2113_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net71),
    .D(net506),
    .Q_N(_0995_),
    .Q(\cell_cfg[29][0] ));
 sg13g2_dfrbp_1 _2114_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net69),
    .D(net509),
    .Q_N(_0994_),
    .Q(\cell_cfg[29][1] ));
 sg13g2_dfrbp_1 _2115_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net67),
    .D(net348),
    .Q_N(_0993_),
    .Q(\cell_cfg[28][0] ));
 sg13g2_dfrbp_1 _2116_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net65),
    .D(net474),
    .Q_N(_0992_),
    .Q(\cell_cfg[28][1] ));
 sg13g2_dfrbp_1 _2117_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net63),
    .D(_0034_),
    .Q_N(_0991_),
    .Q(\cell_cfg[27][0] ));
 sg13g2_dfrbp_1 _2118_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net61),
    .D(_0035_),
    .Q_N(_0990_),
    .Q(\cell_cfg[27][1] ));
 sg13g2_dfrbp_1 _2119_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net59),
    .D(net407),
    .Q_N(_0989_),
    .Q(\cell_cfg[26][0] ));
 sg13g2_dfrbp_1 _2120_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net57),
    .D(net458),
    .Q_N(_0988_),
    .Q(\cell_cfg[26][1] ));
 sg13g2_dfrbp_1 _2121_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net55),
    .D(_0038_),
    .Q_N(_0987_),
    .Q(\cell_cfg[25][0] ));
 sg13g2_dfrbp_1 _2122_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net53),
    .D(net399),
    .Q_N(_0986_),
    .Q(\cell_cfg[25][1] ));
 sg13g2_dfrbp_1 _2123_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net51),
    .D(net512),
    .Q_N(_0985_),
    .Q(\cell_cfg[24][0] ));
 sg13g2_dfrbp_1 _2124_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net49),
    .D(_0041_),
    .Q_N(_0984_),
    .Q(\cell_cfg[24][1] ));
 sg13g2_dfrbp_1 _2125_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net47),
    .D(net419),
    .Q_N(_0983_),
    .Q(\cell_cfg[23][0] ));
 sg13g2_dfrbp_1 _2126_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net45),
    .D(_0043_),
    .Q_N(_0982_),
    .Q(\cell_cfg[23][1] ));
 sg13g2_dfrbp_1 _2127_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net43),
    .D(net366),
    .Q_N(_0981_),
    .Q(\cell_cfg[22][0] ));
 sg13g2_dfrbp_1 _2128_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net41),
    .D(net456),
    .Q_N(_0980_),
    .Q(\cell_cfg[22][1] ));
 sg13g2_dfrbp_1 _2129_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net39),
    .D(_0046_),
    .Q_N(_0979_),
    .Q(\cell_cfg[21][0] ));
 sg13g2_dfrbp_1 _2130_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net37),
    .D(_0047_),
    .Q_N(_0978_),
    .Q(\cell_cfg[21][1] ));
 sg13g2_dfrbp_1 _2131_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net35),
    .D(net340),
    .Q_N(_0977_),
    .Q(\cell_cfg[20][0] ));
 sg13g2_dfrbp_1 _2132_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net33),
    .D(_0049_),
    .Q_N(_0976_),
    .Q(\cell_cfg[20][1] ));
 sg13g2_dfrbp_1 _2133_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net31),
    .D(_0050_),
    .Q_N(_0975_),
    .Q(\cell_cfg[19][0] ));
 sg13g2_dfrbp_1 _2134_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net29),
    .D(_0051_),
    .Q_N(_0974_),
    .Q(\cell_cfg[19][1] ));
 sg13g2_dfrbp_1 _2135_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net27),
    .D(_0052_),
    .Q_N(_0973_),
    .Q(\cell_cfg[18][0] ));
 sg13g2_dfrbp_1 _2136_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net170),
    .D(_0053_),
    .Q_N(_0972_),
    .Q(\cell_cfg[18][1] ));
 sg13g2_dfrbp_1 _2137_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net168),
    .D(net413),
    .Q_N(_0971_),
    .Q(\cell_cfg[17][0] ));
 sg13g2_dfrbp_1 _2138_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net166),
    .D(_0055_),
    .Q_N(_0970_),
    .Q(\cell_cfg[17][1] ));
 sg13g2_dfrbp_1 _2139_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net164),
    .D(_0056_),
    .Q_N(_0969_),
    .Q(\cell_cfg[16][0] ));
 sg13g2_dfrbp_1 _2140_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net162),
    .D(_0057_),
    .Q_N(_0968_),
    .Q(\cell_cfg[16][1] ));
 sg13g2_dfrbp_1 _2141_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net160),
    .D(_0058_),
    .Q_N(_0967_),
    .Q(\cell_cfg[15][0] ));
 sg13g2_dfrbp_1 _2142_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net158),
    .D(_0059_),
    .Q_N(_0966_),
    .Q(\cell_cfg[15][1] ));
 sg13g2_dfrbp_1 _2143_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net156),
    .D(_0060_),
    .Q_N(_0965_),
    .Q(\cell_cfg[14][0] ));
 sg13g2_dfrbp_1 _2144_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net154),
    .D(_0061_),
    .Q_N(_0964_),
    .Q(\cell_cfg[14][1] ));
 sg13g2_dfrbp_1 _2145_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net152),
    .D(net426),
    .Q_N(_0963_),
    .Q(\cell_cfg[13][0] ));
 sg13g2_dfrbp_1 _2146_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net150),
    .D(_0063_),
    .Q_N(_0962_),
    .Q(\cell_cfg[13][1] ));
 sg13g2_dfrbp_1 _2147_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net148),
    .D(net240),
    .Q_N(_0961_),
    .Q(\cell_cfg[12][0] ));
 sg13g2_dfrbp_1 _2148_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net146),
    .D(net395),
    .Q_N(_0960_),
    .Q(\cell_cfg[12][1] ));
 sg13g2_dfrbp_1 _2149_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net144),
    .D(_0066_),
    .Q_N(_0959_),
    .Q(\cell_cfg[11][0] ));
 sg13g2_dfrbp_1 _2150_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net142),
    .D(_0067_),
    .Q_N(_0958_),
    .Q(\cell_cfg[11][1] ));
 sg13g2_dfrbp_1 _2151_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net140),
    .D(net403),
    .Q_N(_0957_),
    .Q(\cell_cfg[10][0] ));
 sg13g2_dfrbp_1 _2152_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net138),
    .D(_0069_),
    .Q_N(_0956_),
    .Q(\cell_cfg[10][1] ));
 sg13g2_dfrbp_1 _2153_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net136),
    .D(_0070_),
    .Q_N(_0955_),
    .Q(\cell_cfg[9][0] ));
 sg13g2_dfrbp_1 _2154_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net134),
    .D(_0071_),
    .Q_N(_0954_),
    .Q(\cell_cfg[9][1] ));
 sg13g2_dfrbp_1 _2155_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net132),
    .D(net362),
    .Q_N(_0953_),
    .Q(\cell_cfg[8][0] ));
 sg13g2_dfrbp_1 _2156_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net130),
    .D(net493),
    .Q_N(_0952_),
    .Q(\cell_cfg[8][1] ));
 sg13g2_dfrbp_1 _2157_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net128),
    .D(_0074_),
    .Q_N(_0951_),
    .Q(\cell_cfg[7][0] ));
 sg13g2_dfrbp_1 _2158_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net126),
    .D(_0075_),
    .Q_N(_0950_),
    .Q(\cell_cfg[7][1] ));
 sg13g2_dfrbp_1 _2159_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net122),
    .D(net385),
    .Q_N(_0949_),
    .Q(\cell_cfg[6][0] ));
 sg13g2_dfrbp_1 _2160_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net118),
    .D(_0077_),
    .Q_N(_0948_),
    .Q(\cell_cfg[6][1] ));
 sg13g2_dfrbp_1 _2161_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net114),
    .D(net452),
    .Q_N(_0000_),
    .Q(\cell_cfg[5][0] ));
 sg13g2_dfrbp_1 _2162_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net110),
    .D(net489),
    .Q_N(_0947_),
    .Q(\cell_cfg[5][1] ));
 sg13g2_dfrbp_1 _2163_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net106),
    .D(_0080_),
    .Q_N(_0946_),
    .Q(\cell_cfg[4][0] ));
 sg13g2_dfrbp_1 _2164_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net102),
    .D(_0081_),
    .Q_N(_0945_),
    .Q(\cell_cfg[4][1] ));
 sg13g2_dfrbp_1 _2165_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net98),
    .D(_0082_),
    .Q_N(_0944_),
    .Q(\cell_cfg[3][0] ));
 sg13g2_dfrbp_1 _2166_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net94),
    .D(_0083_),
    .Q_N(_0943_),
    .Q(\cell_cfg[3][1] ));
 sg13g2_dfrbp_1 _2167_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net90),
    .D(_0084_),
    .Q_N(_0942_),
    .Q(\cell_cfg[2][0] ));
 sg13g2_dfrbp_1 _2168_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net86),
    .D(_0085_),
    .Q_N(_0941_),
    .Q(\cell_cfg[2][1] ));
 sg13g2_dfrbp_1 _2169_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net82),
    .D(net390),
    .Q_N(_0940_),
    .Q(\cell_cfg[1][0] ));
 sg13g2_dfrbp_1 _2170_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net78),
    .D(net471),
    .Q_N(_0939_),
    .Q(\cell_cfg[1][1] ));
 sg13g2_dfrbp_1 _2171_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net74),
    .D(_0088_),
    .Q_N(_0938_),
    .Q(\cell_cfg[0][0] ));
 sg13g2_dfrbp_1 _2172_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net70),
    .D(_0089_),
    .Q_N(_0937_),
    .Q(\cell_cfg[0][1] ));
 sg13g2_dfrbp_1 _2173_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net66),
    .D(_0090_),
    .Q_N(_0001_),
    .Q(en_cells));
 sg13g2_dfrbp_1 _2174_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net62),
    .D(_0091_),
    .Q_N(_0936_),
    .Q(\cell_cfg[8][2] ));
 sg13g2_dfrbp_1 _2175_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net58),
    .D(net236),
    .Q_N(_0935_),
    .Q(\cell_cfg[8][3] ));
 sg13g2_dfrbp_1 _2176_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net54),
    .D(_0093_),
    .Q_N(_0934_),
    .Q(\cell_cfg[0][2] ));
 sg13g2_dfrbp_1 _2177_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net50),
    .D(_0094_),
    .Q_N(_0933_),
    .Q(\cell_cfg[0][3] ));
 sg13g2_dfrbp_1 _2178_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net46),
    .D(_0095_),
    .Q_N(_0932_),
    .Q(\cell_cfg[15][2] ));
 sg13g2_dfrbp_1 _2179_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net42),
    .D(net224),
    .Q_N(_0931_),
    .Q(\cell_cfg[15][3] ));
 sg13g2_dfrbp_1 _2180_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net38),
    .D(_0097_),
    .Q_N(_0930_),
    .Q(\cell_cfg[9][2] ));
 sg13g2_dfrbp_1 _2181_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net34),
    .D(_0098_),
    .Q_N(_0929_),
    .Q(\cell_cfg[9][3] ));
 sg13g2_dfrbp_1 _2182_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net30),
    .D(net368),
    .Q_N(_0928_),
    .Q(\cell_cfg[1][2] ));
 sg13g2_dfrbp_1 _2183_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net26),
    .D(net441),
    .Q_N(_0927_),
    .Q(\cell_cfg[1][3] ));
 sg13g2_dfrbp_1 _2184_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net167),
    .D(_0101_),
    .Q_N(_0926_),
    .Q(\cell_cfg[14][2] ));
 sg13g2_dfrbp_1 _2185_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net163),
    .D(net248),
    .Q_N(_0925_),
    .Q(\cell_cfg[14][3] ));
 sg13g2_dfrbp_1 _2186_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net159),
    .D(net446),
    .Q_N(_0924_),
    .Q(\cell_cfg[10][2] ));
 sg13g2_dfrbp_1 _2187_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net155),
    .D(_0104_),
    .Q_N(_0923_),
    .Q(\cell_cfg[10][3] ));
 sg13g2_dfrbp_1 _2188_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net151),
    .D(_0105_),
    .Q_N(_0922_),
    .Q(\cell_cfg[2][2] ));
 sg13g2_dfrbp_1 _2189_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net147),
    .D(_0106_),
    .Q_N(_0921_),
    .Q(\cell_cfg[2][3] ));
 sg13g2_dfrbp_1 _2190_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net143),
    .D(net345),
    .Q_N(_0920_),
    .Q(\cell_cfg[35][2] ));
 sg13g2_dfrbp_1 _2191_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net139),
    .D(net354),
    .Q_N(_0919_),
    .Q(\cell_cfg[35][3] ));
 sg13g2_dfrbp_1 _2192_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net135),
    .D(net397),
    .Q_N(_0918_),
    .Q(\cell_cfg[13][2] ));
 sg13g2_dfrbp_1 _2193_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net131),
    .D(net244),
    .Q_N(_0917_),
    .Q(\cell_cfg[13][3] ));
 sg13g2_dfrbp_1 _2194_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net127),
    .D(_0111_),
    .Q_N(_0916_),
    .Q(\cell_cfg[34][2] ));
 sg13g2_dfrbp_1 _2195_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net120),
    .D(_0112_),
    .Q_N(_0915_),
    .Q(\cell_cfg[34][3] ));
 sg13g2_dfrbp_1 _2196_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net112),
    .D(net331),
    .Q_N(_0914_),
    .Q(\cell_cfg[33][2] ));
 sg13g2_dfrbp_1 _2197_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net104),
    .D(_0114_),
    .Q_N(_0913_),
    .Q(\cell_cfg[33][3] ));
 sg13g2_dfrbp_1 _2198_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net96),
    .D(_0115_),
    .Q_N(_0912_),
    .Q(\cell_cfg[32][2] ));
 sg13g2_dfrbp_1 _2199_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net88),
    .D(net234),
    .Q_N(_0911_),
    .Q(\cell_cfg[32][3] ));
 sg13g2_dfrbp_1 _2200_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net80),
    .D(_0117_),
    .Q_N(_0910_),
    .Q(\cell_cfg[31][2] ));
 sg13g2_dfrbp_1 _2201_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net72),
    .D(net333),
    .Q_N(_0909_),
    .Q(\cell_cfg[31][3] ));
 sg13g2_dfrbp_1 _2202_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net64),
    .D(_0119_),
    .Q_N(_0908_),
    .Q(\cell_cfg[30][2] ));
 sg13g2_dfrbp_1 _2203_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net56),
    .D(net352),
    .Q_N(_0907_),
    .Q(\cell_cfg[30][3] ));
 sg13g2_dfrbp_1 _2204_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net48),
    .D(net364),
    .Q_N(_0906_),
    .Q(\cell_cfg[29][2] ));
 sg13g2_dfrbp_1 _2205_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net40),
    .D(_0122_),
    .Q_N(_0905_),
    .Q(\cell_cfg[29][3] ));
 sg13g2_dfrbp_1 _2206_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net32),
    .D(_0123_),
    .Q_N(_0904_),
    .Q(\cell_cfg[28][2] ));
 sg13g2_dfrbp_1 _2207_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net169),
    .D(_0124_),
    .Q_N(_0903_),
    .Q(\cell_cfg[28][3] ));
 sg13g2_dfrbp_1 _2208_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net161),
    .D(net424),
    .Q_N(_0902_),
    .Q(\cell_cfg[27][2] ));
 sg13g2_dfrbp_1 _2209_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net153),
    .D(net229),
    .Q_N(_0901_),
    .Q(\cell_cfg[27][3] ));
 sg13g2_dfrbp_1 _2210_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net145),
    .D(_0127_),
    .Q_N(_0900_),
    .Q(\cell_cfg[11][2] ));
 sg13g2_dfrbp_1 _2211_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net137),
    .D(_0128_),
    .Q_N(_0899_),
    .Q(\cell_cfg[11][3] ));
 sg13g2_dfrbp_1 _2212_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net129),
    .D(net433),
    .Q_N(_0898_),
    .Q(\cell_cfg[26][2] ));
 sg13g2_dfrbp_1 _2213_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net116),
    .D(net338),
    .Q_N(_0897_),
    .Q(\cell_cfg[26][3] ));
 sg13g2_dfrbp_1 _2214_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net100),
    .D(net246),
    .Q_N(_0896_),
    .Q(\cell_cfg[3][2] ));
 sg13g2_dfrbp_1 _2215_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net84),
    .D(net393),
    .Q_N(_0895_),
    .Q(\cell_cfg[3][3] ));
 sg13g2_dfrbp_1 _2216_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net68),
    .D(_0133_),
    .Q_N(_0894_),
    .Q(\cell_cfg[25][2] ));
 sg13g2_dfrbp_1 _2217_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net52),
    .D(net342),
    .Q_N(_0893_),
    .Q(\cell_cfg[25][3] ));
 sg13g2_dfrbp_1 _2218_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net36),
    .D(_0135_),
    .Q_N(_0892_),
    .Q(\cell_cfg[24][2] ));
 sg13g2_dfrbp_1 _2219_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net165),
    .D(_0136_),
    .Q_N(_0891_),
    .Q(\cell_cfg[24][3] ));
 sg13g2_dfrbp_1 _2220_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net149),
    .D(_0137_),
    .Q_N(_0890_),
    .Q(\cell_cfg[23][2] ));
 sg13g2_dfrbp_1 _2221_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net133),
    .D(_0138_),
    .Q_N(_0889_),
    .Q(\cell_cfg[23][3] ));
 sg13g2_dfrbp_1 _2222_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net108),
    .D(net415),
    .Q_N(_0888_),
    .Q(\cell_cfg[22][2] ));
 sg13g2_dfrbp_1 _2223_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net76),
    .D(net231),
    .Q_N(_0887_),
    .Q(\cell_cfg[22][3] ));
 sg13g2_dfrbp_1 _2224_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net44),
    .D(_0141_),
    .Q_N(_0886_),
    .Q(\cell_cfg[21][2] ));
 sg13g2_dfrbp_1 _2225_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net157),
    .D(_0142_),
    .Q_N(_0885_),
    .Q(\cell_cfg[21][3] ));
 sg13g2_dfrbp_1 _2226_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net124),
    .D(net335),
    .Q_N(_0884_),
    .Q(\cell_cfg[12][2] ));
 sg13g2_dfrbp_1 _2227_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net60),
    .D(_0144_),
    .Q_N(_0883_),
    .Q(\cell_cfg[12][3] ));
 sg13g2_dfrbp_1 _2228_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net141),
    .D(net379),
    .Q_N(_0882_),
    .Q(\cell_cfg[20][2] ));
 sg13g2_dfrbp_1 _2229_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net28),
    .D(net227),
    .Q_N(_0881_),
    .Q(\cell_cfg[20][3] ));
 sg13g2_tiehi _2135__27 (.L_HI(net27));
 sg13g2_tiehi _2229__28 (.L_HI(net28));
 sg13g2_tiehi _2134__29 (.L_HI(net29));
 sg13g2_tiehi _2182__30 (.L_HI(net30));
 sg13g2_tiehi _2133__31 (.L_HI(net31));
 sg13g2_tiehi _2206__32 (.L_HI(net32));
 sg13g2_tiehi _2132__33 (.L_HI(net33));
 sg13g2_tiehi _2181__34 (.L_HI(net34));
 sg13g2_tiehi _2131__35 (.L_HI(net35));
 sg13g2_tiehi _2218__36 (.L_HI(net36));
 sg13g2_tiehi _2130__37 (.L_HI(net37));
 sg13g2_tiehi _2180__38 (.L_HI(net38));
 sg13g2_tiehi _2129__39 (.L_HI(net39));
 sg13g2_tiehi _2205__40 (.L_HI(net40));
 sg13g2_tiehi _2128__41 (.L_HI(net41));
 sg13g2_tiehi _2179__42 (.L_HI(net42));
 sg13g2_tiehi _2127__43 (.L_HI(net43));
 sg13g2_tiehi _2224__44 (.L_HI(net44));
 sg13g2_tiehi _2126__45 (.L_HI(net45));
 sg13g2_tiehi _2178__46 (.L_HI(net46));
 sg13g2_tiehi _2125__47 (.L_HI(net47));
 sg13g2_tiehi _2204__48 (.L_HI(net48));
 sg13g2_tiehi _2124__49 (.L_HI(net49));
 sg13g2_tiehi _2177__50 (.L_HI(net50));
 sg13g2_tiehi _2123__51 (.L_HI(net51));
 sg13g2_tiehi _2217__52 (.L_HI(net52));
 sg13g2_tiehi _2122__53 (.L_HI(net53));
 sg13g2_tiehi _2176__54 (.L_HI(net54));
 sg13g2_tiehi _2121__55 (.L_HI(net55));
 sg13g2_tiehi _2203__56 (.L_HI(net56));
 sg13g2_tiehi _2120__57 (.L_HI(net57));
 sg13g2_tiehi _2175__58 (.L_HI(net58));
 sg13g2_tiehi _2119__59 (.L_HI(net59));
 sg13g2_tiehi _2227__60 (.L_HI(net60));
 sg13g2_tiehi _2118__61 (.L_HI(net61));
 sg13g2_tiehi _2174__62 (.L_HI(net62));
 sg13g2_tiehi _2117__63 (.L_HI(net63));
 sg13g2_tiehi _2202__64 (.L_HI(net64));
 sg13g2_tiehi _2116__65 (.L_HI(net65));
 sg13g2_tiehi _2173__66 (.L_HI(net66));
 sg13g2_tiehi _2115__67 (.L_HI(net67));
 sg13g2_tiehi _2216__68 (.L_HI(net68));
 sg13g2_tiehi _2114__69 (.L_HI(net69));
 sg13g2_tiehi _2172__70 (.L_HI(net70));
 sg13g2_tiehi _2113__71 (.L_HI(net71));
 sg13g2_tiehi _2201__72 (.L_HI(net72));
 sg13g2_tiehi _2112__73 (.L_HI(net73));
 sg13g2_tiehi _2171__74 (.L_HI(net74));
 sg13g2_tiehi _2111__75 (.L_HI(net75));
 sg13g2_tiehi _2223__76 (.L_HI(net76));
 sg13g2_tiehi _2110__77 (.L_HI(net77));
 sg13g2_tiehi _2170__78 (.L_HI(net78));
 sg13g2_tiehi _2109__79 (.L_HI(net79));
 sg13g2_tiehi _2200__80 (.L_HI(net80));
 sg13g2_tiehi _2108__81 (.L_HI(net81));
 sg13g2_tiehi _2169__82 (.L_HI(net82));
 sg13g2_tiehi _2107__83 (.L_HI(net83));
 sg13g2_tiehi _2215__84 (.L_HI(net84));
 sg13g2_tiehi _2106__85 (.L_HI(net85));
 sg13g2_tiehi _2168__86 (.L_HI(net86));
 sg13g2_tiehi _2105__87 (.L_HI(net87));
 sg13g2_tiehi _2199__88 (.L_HI(net88));
 sg13g2_tiehi _2104__89 (.L_HI(net89));
 sg13g2_tiehi _2167__90 (.L_HI(net90));
 sg13g2_tiehi _2103__91 (.L_HI(net91));
 sg13g2_tiehi _2085__92 (.L_HI(net92));
 sg13g2_tiehi _2102__93 (.L_HI(net93));
 sg13g2_tiehi _2166__94 (.L_HI(net94));
 sg13g2_tiehi _2101__95 (.L_HI(net95));
 sg13g2_tiehi _2198__96 (.L_HI(net96));
 sg13g2_tiehi _2100__97 (.L_HI(net97));
 sg13g2_tiehi _2165__98 (.L_HI(net98));
 sg13g2_tiehi _2099__99 (.L_HI(net99));
 sg13g2_tiehi _2214__100 (.L_HI(net100));
 sg13g2_tiehi _2098__101 (.L_HI(net101));
 sg13g2_tiehi _2164__102 (.L_HI(net102));
 sg13g2_tiehi _2097__103 (.L_HI(net103));
 sg13g2_tiehi _2197__104 (.L_HI(net104));
 sg13g2_tiehi _2096__105 (.L_HI(net105));
 sg13g2_tiehi _2163__106 (.L_HI(net106));
 sg13g2_tiehi _2095__107 (.L_HI(net107));
 sg13g2_tiehi _2222__108 (.L_HI(net108));
 sg13g2_tiehi _2094__109 (.L_HI(net109));
 sg13g2_tiehi _2162__110 (.L_HI(net110));
 sg13g2_tiehi _2093__111 (.L_HI(net111));
 sg13g2_tiehi _2196__112 (.L_HI(net112));
 sg13g2_tiehi _2092__113 (.L_HI(net113));
 sg13g2_tiehi _2161__114 (.L_HI(net114));
 sg13g2_tiehi _2091__115 (.L_HI(net115));
 sg13g2_tiehi _2213__116 (.L_HI(net116));
 sg13g2_tiehi _2090__117 (.L_HI(net117));
 sg13g2_tiehi _2160__118 (.L_HI(net118));
 sg13g2_tiehi _2089__119 (.L_HI(net119));
 sg13g2_tiehi _2195__120 (.L_HI(net120));
 sg13g2_tiehi _2088__121 (.L_HI(net121));
 sg13g2_tiehi _2159__122 (.L_HI(net122));
 sg13g2_tiehi _2087__123 (.L_HI(net123));
 sg13g2_tiehi _2226__124 (.L_HI(net124));
 sg13g2_tiehi _2086__125 (.L_HI(net125));
 sg13g2_tiehi _2158__126 (.L_HI(net126));
 sg13g2_tiehi _2194__127 (.L_HI(net127));
 sg13g2_tiehi _2157__128 (.L_HI(net128));
 sg13g2_tiehi _2212__129 (.L_HI(net129));
 sg13g2_tiehi _2156__130 (.L_HI(net130));
 sg13g2_tiehi _2193__131 (.L_HI(net131));
 sg13g2_tiehi _2155__132 (.L_HI(net132));
 sg13g2_tiehi _2221__133 (.L_HI(net133));
 sg13g2_tiehi _2154__134 (.L_HI(net134));
 sg13g2_tiehi _2192__135 (.L_HI(net135));
 sg13g2_tiehi _2153__136 (.L_HI(net136));
 sg13g2_tiehi _2211__137 (.L_HI(net137));
 sg13g2_tiehi _2152__138 (.L_HI(net138));
 sg13g2_tiehi _2191__139 (.L_HI(net139));
 sg13g2_tiehi _2151__140 (.L_HI(net140));
 sg13g2_tiehi _2228__141 (.L_HI(net141));
 sg13g2_tiehi _2150__142 (.L_HI(net142));
 sg13g2_tiehi _2190__143 (.L_HI(net143));
 sg13g2_tiehi _2149__144 (.L_HI(net144));
 sg13g2_tiehi _2210__145 (.L_HI(net145));
 sg13g2_tiehi _2148__146 (.L_HI(net146));
 sg13g2_tiehi _2189__147 (.L_HI(net147));
 sg13g2_tiehi _2147__148 (.L_HI(net148));
 sg13g2_tiehi _2220__149 (.L_HI(net149));
 sg13g2_tiehi _2146__150 (.L_HI(net150));
 sg13g2_tiehi _2188__151 (.L_HI(net151));
 sg13g2_tiehi _2145__152 (.L_HI(net152));
 sg13g2_tiehi _2209__153 (.L_HI(net153));
 sg13g2_tiehi _2144__154 (.L_HI(net154));
 sg13g2_tiehi _2187__155 (.L_HI(net155));
 sg13g2_tiehi _2143__156 (.L_HI(net156));
 sg13g2_tiehi _2225__157 (.L_HI(net157));
 sg13g2_tiehi _2142__158 (.L_HI(net158));
 sg13g2_tiehi _2186__159 (.L_HI(net159));
 sg13g2_tiehi _2141__160 (.L_HI(net160));
 sg13g2_tiehi _2208__161 (.L_HI(net161));
 sg13g2_tiehi _2140__162 (.L_HI(net162));
 sg13g2_tiehi _2185__163 (.L_HI(net163));
 sg13g2_tiehi _2139__164 (.L_HI(net164));
 sg13g2_tiehi _2219__165 (.L_HI(net165));
 sg13g2_tiehi _2138__166 (.L_HI(net166));
 sg13g2_tiehi _2184__167 (.L_HI(net167));
 sg13g2_tiehi _2137__168 (.L_HI(net168));
 sg13g2_tiehi _2207__169 (.L_HI(net169));
 sg13g2_tiehi _2136__170 (.L_HI(net170));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_emilian_muxpga_7 (.L_LO(net7));
 sg13g2_tielo tt_um_emilian_muxpga_8 (.L_LO(net8));
 sg13g2_tielo tt_um_emilian_muxpga_9 (.L_LO(net9));
 sg13g2_tielo tt_um_emilian_muxpga_10 (.L_LO(net10));
 sg13g2_tielo tt_um_emilian_muxpga_11 (.L_LO(net11));
 sg13g2_tielo tt_um_emilian_muxpga_12 (.L_LO(net12));
 sg13g2_tielo tt_um_emilian_muxpga_13 (.L_LO(net13));
 sg13g2_tielo tt_um_emilian_muxpga_14 (.L_LO(net14));
 sg13g2_tielo tt_um_emilian_muxpga_15 (.L_LO(net15));
 sg13g2_tielo tt_um_emilian_muxpga_16 (.L_LO(net16));
 sg13g2_tielo tt_um_emilian_muxpga_17 (.L_LO(net17));
 sg13g2_tielo tt_um_emilian_muxpga_18 (.L_LO(net18));
 sg13g2_tielo tt_um_emilian_muxpga_19 (.L_LO(net19));
 sg13g2_tielo tt_um_emilian_muxpga_20 (.L_LO(net20));
 sg13g2_tielo tt_um_emilian_muxpga_21 (.L_LO(net21));
 sg13g2_tielo tt_um_emilian_muxpga_22 (.L_LO(net22));
 sg13g2_tielo tt_um_emilian_muxpga_23 (.L_LO(net23));
 sg13g2_tielo tt_um_emilian_muxpga_24 (.L_LO(net24));
 sg13g2_tielo tt_um_emilian_muxpga_25 (.L_LO(net25));
 sg13g2_tiehi _2183__26 (.L_HI(net26));
 sg13g2_buf_4 fanout251 (.X(net251),
    .A(net252));
 sg13g2_buf_4 fanout252 (.X(net252),
    .A(net255));
 sg13g2_buf_4 fanout253 (.X(net253),
    .A(net254));
 sg13g2_buf_4 fanout254 (.X(net254),
    .A(net255));
 sg13g2_buf_2 fanout255 (.A(_0001_),
    .X(net255));
 sg13g2_buf_2 fanout256 (.A(net257),
    .X(net256));
 sg13g2_buf_1 fanout257 (.A(net259),
    .X(net257));
 sg13g2_buf_2 fanout258 (.A(net259),
    .X(net258));
 sg13g2_buf_4 fanout259 (.X(net259),
    .A(net265));
 sg13g2_buf_4 fanout260 (.X(net260),
    .A(net264));
 sg13g2_buf_2 fanout261 (.A(net264),
    .X(net261));
 sg13g2_buf_2 fanout262 (.A(net264),
    .X(net262));
 sg13g2_buf_1 fanout263 (.A(net264),
    .X(net263));
 sg13g2_buf_2 fanout264 (.A(net265),
    .X(net264));
 sg13g2_buf_2 fanout265 (.A(_0747_),
    .X(net265));
 sg13g2_buf_2 fanout266 (.A(net269),
    .X(net266));
 sg13g2_buf_2 fanout267 (.A(net268),
    .X(net267));
 sg13g2_buf_2 fanout268 (.A(net269),
    .X(net268));
 sg13g2_buf_2 fanout269 (.A(_0747_),
    .X(net269));
 sg13g2_buf_2 fanout270 (.A(net271),
    .X(net270));
 sg13g2_buf_2 fanout271 (.A(net272),
    .X(net271));
 sg13g2_buf_2 fanout272 (.A(_0747_),
    .X(net272));
 sg13g2_buf_2 fanout273 (.A(net276),
    .X(net273));
 sg13g2_buf_1 fanout274 (.A(net276),
    .X(net274));
 sg13g2_buf_2 fanout275 (.A(net276),
    .X(net275));
 sg13g2_buf_1 fanout276 (.A(net289),
    .X(net276));
 sg13g2_buf_2 fanout277 (.A(net278),
    .X(net277));
 sg13g2_buf_2 fanout278 (.A(net281),
    .X(net278));
 sg13g2_buf_2 fanout279 (.A(net280),
    .X(net279));
 sg13g2_buf_2 fanout280 (.A(net281),
    .X(net280));
 sg13g2_buf_2 fanout281 (.A(net289),
    .X(net281));
 sg13g2_buf_2 fanout282 (.A(net284),
    .X(net282));
 sg13g2_buf_2 fanout283 (.A(net284),
    .X(net283));
 sg13g2_buf_2 fanout284 (.A(net289),
    .X(net284));
 sg13g2_buf_2 fanout285 (.A(net288),
    .X(net285));
 sg13g2_buf_2 fanout286 (.A(net288),
    .X(net286));
 sg13g2_buf_1 fanout287 (.A(net288),
    .X(net287));
 sg13g2_buf_2 fanout288 (.A(net289),
    .X(net288));
 sg13g2_buf_2 fanout289 (.A(_0746_),
    .X(net289));
 sg13g2_buf_2 fanout290 (.A(net297),
    .X(net290));
 sg13g2_buf_2 fanout291 (.A(net292),
    .X(net291));
 sg13g2_buf_2 fanout292 (.A(net297),
    .X(net292));
 sg13g2_buf_2 fanout293 (.A(net296),
    .X(net293));
 sg13g2_buf_1 fanout294 (.A(net296),
    .X(net294));
 sg13g2_buf_2 fanout295 (.A(net296),
    .X(net295));
 sg13g2_buf_2 fanout296 (.A(net297),
    .X(net296));
 sg13g2_buf_2 fanout297 (.A(_0746_),
    .X(net297));
 sg13g2_buf_2 fanout298 (.A(net304),
    .X(net298));
 sg13g2_buf_2 fanout299 (.A(net304),
    .X(net299));
 sg13g2_buf_2 fanout300 (.A(net301),
    .X(net300));
 sg13g2_buf_2 fanout301 (.A(net304),
    .X(net301));
 sg13g2_buf_2 fanout302 (.A(net303),
    .X(net302));
 sg13g2_buf_2 fanout303 (.A(net304),
    .X(net303));
 sg13g2_buf_2 fanout304 (.A(_0746_),
    .X(net304));
 sg13g2_buf_2 fanout305 (.A(net307),
    .X(net305));
 sg13g2_buf_2 fanout306 (.A(net307),
    .X(net306));
 sg13g2_buf_2 fanout307 (.A(_0396_),
    .X(net307));
 sg13g2_buf_2 fanout308 (.A(net310),
    .X(net308));
 sg13g2_buf_2 fanout309 (.A(net310),
    .X(net309));
 sg13g2_buf_2 fanout310 (.A(_0396_),
    .X(net310));
 sg13g2_buf_2 fanout311 (.A(net313),
    .X(net311));
 sg13g2_buf_2 fanout312 (.A(net313),
    .X(net312));
 sg13g2_buf_2 fanout313 (.A(net316),
    .X(net313));
 sg13g2_buf_4 fanout314 (.X(net314),
    .A(net315));
 sg13g2_buf_2 fanout315 (.A(net316),
    .X(net315));
 sg13g2_buf_2 fanout316 (.A(_0396_),
    .X(net316));
 sg13g2_buf_2 fanout317 (.A(net318),
    .X(net317));
 sg13g2_buf_4 fanout318 (.X(net318),
    .A(ui_in[0]));
 sg13g2_buf_2 fanout319 (.A(net321),
    .X(net319));
 sg13g2_buf_4 fanout320 (.X(net320),
    .A(net321));
 sg13g2_buf_2 fanout321 (.A(rst_n),
    .X(net321));
 sg13g2_buf_2 fanout322 (.A(net324),
    .X(net322));
 sg13g2_buf_1 fanout323 (.A(net324),
    .X(net323));
 sg13g2_buf_2 fanout324 (.A(rst_n),
    .X(net324));
 sg13g2_buf_2 fanout325 (.A(net326),
    .X(net325));
 sg13g2_buf_4 fanout326 (.X(net326),
    .A(net329));
 sg13g2_buf_2 fanout327 (.A(net329),
    .X(net327));
 sg13g2_buf_2 fanout328 (.A(net329),
    .X(net328));
 sg13g2_buf_4 fanout329 (.X(net329),
    .A(rst_n));
 sg13g2_buf_2 input1 (.A(ui_in[1]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[2]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[3]),
    .X(net3));
 sg13g2_buf_2 input4 (.A(ui_in[6]),
    .X(net4));
 sg13g2_buf_2 input5 (.A(ui_in[7]),
    .X(net5));
 sg13g2_tielo tt_um_emilian_muxpga_6 (.L_LO(net6));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_buf_2 clkbuf_5_0__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_0__leaf_clk));
 sg13g2_buf_2 clkbuf_5_1__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_1__leaf_clk));
 sg13g2_buf_2 clkbuf_5_2__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_2__leaf_clk));
 sg13g2_buf_2 clkbuf_5_3__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_3__leaf_clk));
 sg13g2_buf_2 clkbuf_5_4__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_4__leaf_clk));
 sg13g2_buf_2 clkbuf_5_5__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_5__leaf_clk));
 sg13g2_buf_2 clkbuf_5_6__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_6__leaf_clk));
 sg13g2_buf_2 clkbuf_5_7__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_7__leaf_clk));
 sg13g2_buf_2 clkbuf_5_8__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_8__leaf_clk));
 sg13g2_buf_2 clkbuf_5_9__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_9__leaf_clk));
 sg13g2_buf_2 clkbuf_5_10__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_10__leaf_clk));
 sg13g2_buf_2 clkbuf_5_11__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_11__leaf_clk));
 sg13g2_buf_2 clkbuf_5_12__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_12__leaf_clk));
 sg13g2_buf_2 clkbuf_5_13__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_13__leaf_clk));
 sg13g2_buf_2 clkbuf_5_14__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_14__leaf_clk));
 sg13g2_buf_2 clkbuf_5_15__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_15__leaf_clk));
 sg13g2_buf_2 clkbuf_5_16__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_16__leaf_clk));
 sg13g2_buf_2 clkbuf_5_17__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_17__leaf_clk));
 sg13g2_buf_2 clkbuf_5_18__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_18__leaf_clk));
 sg13g2_buf_2 clkbuf_5_19__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_19__leaf_clk));
 sg13g2_buf_2 clkbuf_5_20__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_20__leaf_clk));
 sg13g2_buf_2 clkbuf_5_21__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_21__leaf_clk));
 sg13g2_buf_2 clkbuf_5_22__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_22__leaf_clk));
 sg13g2_buf_2 clkbuf_5_23__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_23__leaf_clk));
 sg13g2_buf_2 clkbuf_5_24__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_24__leaf_clk));
 sg13g2_buf_2 clkbuf_5_25__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_25__leaf_clk));
 sg13g2_buf_2 clkbuf_5_26__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_26__leaf_clk));
 sg13g2_buf_2 clkbuf_5_27__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_27__leaf_clk));
 sg13g2_buf_2 clkbuf_5_28__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_28__leaf_clk));
 sg13g2_buf_2 clkbuf_5_29__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_29__leaf_clk));
 sg13g2_buf_2 clkbuf_5_30__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_30__leaf_clk));
 sg13g2_buf_2 clkbuf_5_31__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_31__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_5_3__leaf_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_5_5__leaf_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_5_7__leaf_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_5_9__leaf_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_5_11__leaf_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_5_13__leaf_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_5_15__leaf_clk));
 sg13g2_inv_1 clkload7 (.A(clknet_5_17__leaf_clk));
 sg13g2_inv_1 clkload8 (.A(clknet_5_19__leaf_clk));
 sg13g2_inv_1 clkload9 (.A(clknet_5_21__leaf_clk));
 sg13g2_inv_1 clkload10 (.A(clknet_5_23__leaf_clk));
 sg13g2_inv_1 clkload11 (.A(clknet_5_25__leaf_clk));
 sg13g2_inv_1 clkload12 (.A(clknet_5_27__leaf_clk));
 sg13g2_inv_1 clkload13 (.A(clknet_5_29__leaf_clk));
 sg13g2_inv_1 clkload14 (.A(clknet_5_31__leaf_clk));
 sg13g2_buf_2 rebuffer1 (.A(\genrow[2].gencol[5].genblk1.c.bufs[0].A ),
    .X(net171));
 sg13g2_buf_2 rebuffer2 (.A(\genrow[6].gencol[5].genblk1.c.bufs[0].A ),
    .X(net172));
 sg13g2_dlygate4sd1_1 rebuffer3 (.A(net172),
    .X(net173));
 sg13g2_dlygate4sd1_1 rebuffer4 (.A(\genrow[5].gencol[4].genblk1.c.bufs[0].A ),
    .X(net174));
 sg13g2_dlygate4sd1_1 rebuffer5 (.A(\genrow[5].gencol[4].genblk1.c.bufs[0].A ),
    .X(net175));
 sg13g2_dlygate4sd1_1 rebuffer10 (.A(\genrow[6].gencol[1].genblk1.c.bufs[0].A ),
    .X(net180));
 sg13g2_dlygate4sd1_1 rebuffer28 (.A(\genrow[4].gencol[5].genblk1.c.bufs[0].A ),
    .X(net198));
 sg13g2_dlygate4sd1_1 rebuffer29 (.A(net198),
    .X(net199));
 sg13g2_dlygate4sd1_1 rebuffer30 (.A(net212),
    .X(net200));
 sg13g2_dlygate4sd1_1 rebuffer31 (.A(_0441_),
    .X(net201));
 sg13g2_dlygate4sd1_1 rebuffer38 (.A(\genrow[5].gencol[4].genblk1.c.bufs[0].A ),
    .X(net208));
 sg13g2_dlygate4sd1_1 rebuffer39 (.A(\genrow[5].gencol[3].genblk1.c.bufs[0].A ),
    .X(net209));
 sg13g2_dlygate4sd1_1 rebuffer40 (.A(\genrow[4].gencol[0].genblk1.c.bufs[0].A ),
    .X(net210));
 sg13g2_dlygate4sd1_1 rebuffer41 (.A(\genrow[3].gencol[5].genblk1.c.bufs[0].A ),
    .X(net211));
 sg13g2_dlygate4sd1_1 rebuffer42 (.A(_0441_),
    .X(net212));
 sg13g2_dlygate4sd1_1 rebuffer43 (.A(\genrow[6].gencol[2].genblk1.c.bufs[0].A ),
    .X(net213));
 sg13g2_dlygate4sd1_1 rebuffer44 (.A(\genrow[6].gencol[2].genblk1.c.bufs[0].A ),
    .X(net214));
 sg13g2_dlygate4sd1_1 rebuffer45 (.A(\genrow[6].gencol[2].genblk1.c.bufs[0].A ),
    .X(net215));
 sg13g2_dlygate4sd1_1 rebuffer46 (.A(\genrow[5].gencol[0].genblk1.c.bufs[0].A ),
    .X(net216));
 sg13g2_buf_1 rebuffer51 (.A(\genrow[3].gencol[4].genblk1.c.bufs[0].A ),
    .X(net221));
 sg13g2_dlygate4sd1_1 rebuffer52 (.A(\genrow[4].gencol[4].genblk1.c.bufs[0].A ),
    .X(net222));
 sg13g2_dlygate4sd3_1 hold53 (.A(\cell_cfg[15][3] ),
    .X(net223));
 sg13g2_dlygate4sd3_1 hold54 (.A(_0096_),
    .X(net224));
 sg13g2_dlygate4sd3_1 hold55 (.A(en_cells),
    .X(net225));
 sg13g2_dlygate4sd3_1 hold56 (.A(\cell_cfg[20][3] ),
    .X(net226));
 sg13g2_dlygate4sd3_1 hold57 (.A(_0146_),
    .X(net227));
 sg13g2_dlygate4sd3_1 hold58 (.A(\cell_cfg[27][3] ),
    .X(net228));
 sg13g2_dlygate4sd3_1 hold59 (.A(_0126_),
    .X(net229));
 sg13g2_dlygate4sd3_1 hold60 (.A(\cell_cfg[22][3] ),
    .X(net230));
 sg13g2_dlygate4sd3_1 hold61 (.A(_0140_),
    .X(net231));
 sg13g2_dlygate4sd3_1 hold62 (.A(\cell_cfg[2][0] ),
    .X(net232));
 sg13g2_dlygate4sd3_1 hold63 (.A(\cell_cfg[32][3] ),
    .X(net233));
 sg13g2_dlygate4sd3_1 hold64 (.A(_0116_),
    .X(net234));
 sg13g2_dlygate4sd3_1 hold65 (.A(\cell_cfg[8][3] ),
    .X(net235));
 sg13g2_dlygate4sd3_1 hold66 (.A(_0092_),
    .X(net236));
 sg13g2_dlygate4sd3_1 hold67 (.A(\cell_cfg[21][3] ),
    .X(net237));
 sg13g2_dlygate4sd3_1 hold68 (.A(\cell_cfg[9][3] ),
    .X(net238));
 sg13g2_dlygate4sd3_1 hold69 (.A(\cell_cfg[11][0] ),
    .X(net239));
 sg13g2_dlygate4sd3_1 hold70 (.A(_0064_),
    .X(net240));
 sg13g2_dlygate4sd3_1 hold71 (.A(\cell_cfg[23][3] ),
    .X(net241));
 sg13g2_dlygate4sd3_1 hold72 (.A(\cell_cfg[28][3] ),
    .X(net242));
 sg13g2_dlygate4sd3_1 hold73 (.A(\cell_cfg[12][3] ),
    .X(net243));
 sg13g2_dlygate4sd3_1 hold74 (.A(_0110_),
    .X(net244));
 sg13g2_dlygate4sd3_1 hold75 (.A(\cell_cfg[3][2] ),
    .X(net245));
 sg13g2_dlygate4sd3_1 hold76 (.A(_0131_),
    .X(net246));
 sg13g2_dlygate4sd3_1 hold77 (.A(\cell_cfg[14][3] ),
    .X(net247));
 sg13g2_dlygate4sd3_1 hold78 (.A(_0102_),
    .X(net248));
 sg13g2_dlygate4sd3_1 hold79 (.A(\cell_cfg[11][3] ),
    .X(net249));
 sg13g2_dlygate4sd3_1 hold80 (.A(\cell_cfg[10][3] ),
    .X(net250));
 sg13g2_dlygate4sd3_1 hold81 (.A(\cell_cfg[33][2] ),
    .X(net330));
 sg13g2_dlygate4sd3_1 hold82 (.A(_0113_),
    .X(net331));
 sg13g2_dlygate4sd3_1 hold83 (.A(\cell_cfg[31][3] ),
    .X(net332));
 sg13g2_dlygate4sd3_1 hold84 (.A(_0118_),
    .X(net333));
 sg13g2_dlygate4sd3_1 hold85 (.A(\cell_cfg[11][2] ),
    .X(net334));
 sg13g2_dlygate4sd3_1 hold86 (.A(_0143_),
    .X(net335));
 sg13g2_dlygate4sd3_1 hold87 (.A(\cell_cfg[33][3] ),
    .X(net336));
 sg13g2_dlygate4sd3_1 hold88 (.A(\cell_cfg[26][3] ),
    .X(net337));
 sg13g2_dlygate4sd3_1 hold89 (.A(_0130_),
    .X(net338));
 sg13g2_dlygate4sd3_1 hold90 (.A(\cell_cfg[19][0] ),
    .X(net339));
 sg13g2_dlygate4sd3_1 hold91 (.A(_0048_),
    .X(net340));
 sg13g2_dlygate4sd3_1 hold92 (.A(\cell_cfg[25][3] ),
    .X(net341));
 sg13g2_dlygate4sd3_1 hold93 (.A(_0134_),
    .X(net342));
 sg13g2_dlygate4sd3_1 hold94 (.A(\cell_cfg[1][0] ),
    .X(net343));
 sg13g2_dlygate4sd3_1 hold95 (.A(\cell_cfg[35][2] ),
    .X(net344));
 sg13g2_dlygate4sd3_1 hold96 (.A(_0107_),
    .X(net345));
 sg13g2_dlygate4sd3_1 hold97 (.A(\cell_cfg[16][3] ),
    .X(net346));
 sg13g2_dlygate4sd3_1 hold98 (.A(\cell_cfg[27][0] ),
    .X(net347));
 sg13g2_dlygate4sd3_1 hold99 (.A(_0032_),
    .X(net348));
 sg13g2_dlygate4sd3_1 hold100 (.A(\cell_cfg[18][2] ),
    .X(net349));
 sg13g2_dlygate4sd3_1 hold101 (.A(_0016_),
    .X(net350));
 sg13g2_dlygate4sd3_1 hold102 (.A(\cell_cfg[30][3] ),
    .X(net351));
 sg13g2_dlygate4sd3_1 hold103 (.A(_0120_),
    .X(net352));
 sg13g2_dlygate4sd3_1 hold104 (.A(\cell_cfg[35][3] ),
    .X(net353));
 sg13g2_dlygate4sd3_1 hold105 (.A(_0108_),
    .X(net354));
 sg13g2_dlygate4sd3_1 hold106 (.A(\cell_cfg[5][3] ),
    .X(net355));
 sg13g2_dlygate4sd3_1 hold107 (.A(_0009_),
    .X(net356));
 sg13g2_dlygate4sd3_1 hold108 (.A(\cell_cfg[34][2] ),
    .X(net357));
 sg13g2_dlygate4sd3_1 hold109 (.A(\cell_cfg[10][0] ),
    .X(net358));
 sg13g2_dlygate4sd3_1 hold110 (.A(\cell_cfg[33][1] ),
    .X(net359));
 sg13g2_dlygate4sd3_1 hold111 (.A(_0785_),
    .X(net360));
 sg13g2_dlygate4sd3_1 hold112 (.A(\cell_cfg[7][0] ),
    .X(net361));
 sg13g2_dlygate4sd3_1 hold113 (.A(_0072_),
    .X(net362));
 sg13g2_dlygate4sd3_1 hold114 (.A(\cell_cfg[29][2] ),
    .X(net363));
 sg13g2_dlygate4sd3_1 hold115 (.A(_0121_),
    .X(net364));
 sg13g2_dlygate4sd3_1 hold116 (.A(\cell_cfg[21][0] ),
    .X(net365));
 sg13g2_dlygate4sd3_1 hold117 (.A(_0044_),
    .X(net366));
 sg13g2_dlygate4sd3_1 hold118 (.A(\cell_cfg[1][2] ),
    .X(net367));
 sg13g2_dlygate4sd3_1 hold119 (.A(_0099_),
    .X(net368));
 sg13g2_dlygate4sd3_1 hold120 (.A(\cell_cfg[35][0] ),
    .X(net369));
 sg13g2_dlygate4sd3_1 hold121 (.A(_0769_),
    .X(net370));
 sg13g2_dlygate4sd3_1 hold122 (.A(\cell_cfg[18][0] ),
    .X(net371));
 sg13g2_dlygate4sd3_1 hold123 (.A(\cell_cfg[2][2] ),
    .X(net372));
 sg13g2_dlygate4sd3_1 hold124 (.A(\cell_cfg[34][3] ),
    .X(net373));
 sg13g2_dlygate4sd3_1 hold125 (.A(\cell_cfg[16][2] ),
    .X(net374));
 sg13g2_dlygate4sd3_1 hold126 (.A(_0002_),
    .X(net375));
 sg13g2_dlygate4sd3_1 hold127 (.A(\cell_cfg[6][3] ),
    .X(net376));
 sg13g2_dlygate4sd3_1 hold128 (.A(_0011_),
    .X(net377));
 sg13g2_dlygate4sd3_1 hold129 (.A(\cell_cfg[20][2] ),
    .X(net378));
 sg13g2_dlygate4sd3_1 hold130 (.A(_0145_),
    .X(net379));
 sg13g2_dlygate4sd3_1 hold131 (.A(\cell_cfg[17][3] ),
    .X(net380));
 sg13g2_dlygate4sd3_1 hold132 (.A(_0007_),
    .X(net381));
 sg13g2_dlygate4sd3_1 hold133 (.A(\cell_cfg[4][3] ),
    .X(net382));
 sg13g2_dlygate4sd3_1 hold134 (.A(\cell_cfg[6][0] ),
    .X(net383));
 sg13g2_dlygate4sd3_1 hold135 (.A(_0236_),
    .X(net384));
 sg13g2_dlygate4sd3_1 hold136 (.A(_0076_),
    .X(net385));
 sg13g2_dlygate4sd3_1 hold137 (.A(\cell_cfg[30][0] ),
    .X(net386));
 sg13g2_dlygate4sd3_1 hold138 (.A(_0026_),
    .X(net387));
 sg13g2_dlygate4sd3_1 hold139 (.A(\cell_cfg[4][2] ),
    .X(net388));
 sg13g2_dlygate4sd3_1 hold140 (.A(\cell_cfg[0][0] ),
    .X(net389));
 sg13g2_dlygate4sd3_1 hold141 (.A(_0086_),
    .X(net390));
 sg13g2_dlygate4sd3_1 hold142 (.A(\cell_cfg[7][2] ),
    .X(net391));
 sg13g2_dlygate4sd3_1 hold143 (.A(\cell_cfg[3][3] ),
    .X(net392));
 sg13g2_dlygate4sd3_1 hold144 (.A(_0132_),
    .X(net393));
 sg13g2_dlygate4sd3_1 hold145 (.A(\cell_cfg[11][1] ),
    .X(net394));
 sg13g2_dlygate4sd3_1 hold146 (.A(_0065_),
    .X(net395));
 sg13g2_dlygate4sd3_1 hold147 (.A(\cell_cfg[13][2] ),
    .X(net396));
 sg13g2_dlygate4sd3_1 hold148 (.A(_0109_),
    .X(net397));
 sg13g2_dlygate4sd3_1 hold149 (.A(\cell_cfg[24][1] ),
    .X(net398));
 sg13g2_dlygate4sd3_1 hold150 (.A(_0039_),
    .X(net399));
 sg13g2_dlygate4sd3_1 hold151 (.A(\cell_cfg[8][0] ),
    .X(net400));
 sg13g2_dlygate4sd3_1 hold152 (.A(\cell_cfg[6][2] ),
    .X(net401));
 sg13g2_dlygate4sd3_1 hold153 (.A(\cell_cfg[9][0] ),
    .X(net402));
 sg13g2_dlygate4sd3_1 hold154 (.A(_0068_),
    .X(net403));
 sg13g2_dlygate4sd3_1 hold155 (.A(\cell_cfg[14][0] ),
    .X(net404));
 sg13g2_dlygate4sd3_1 hold156 (.A(\cell_cfg[5][2] ),
    .X(net405));
 sg13g2_dlygate4sd3_1 hold157 (.A(\cell_cfg[25][0] ),
    .X(net406));
 sg13g2_dlygate4sd3_1 hold158 (.A(_0036_),
    .X(net407));
 sg13g2_dlygate4sd3_1 hold159 (.A(\cell_cfg[13][1] ),
    .X(net408));
 sg13g2_dlygate4sd3_1 hold160 (.A(\cell_cfg[31][0] ),
    .X(net409));
 sg13g2_dlygate4sd3_1 hold161 (.A(_0024_),
    .X(net410));
 sg13g2_dlygate4sd3_1 hold162 (.A(\cell_cfg[17][0] ),
    .X(net411));
 sg13g2_dlygate4sd3_1 hold163 (.A(_0164_),
    .X(net412));
 sg13g2_dlygate4sd3_1 hold164 (.A(_0054_),
    .X(net413));
 sg13g2_dlygate4sd3_1 hold165 (.A(\cell_cfg[22][2] ),
    .X(net414));
 sg13g2_dlygate4sd3_1 hold166 (.A(_0139_),
    .X(net415));
 sg13g2_dlygate4sd3_1 hold167 (.A(\cell_cfg[13][0] ),
    .X(net416));
 sg13g2_dlygate4sd3_1 hold168 (.A(\cell_cfg[26][0] ),
    .X(net417));
 sg13g2_dlygate4sd3_1 hold169 (.A(\cell_cfg[22][0] ),
    .X(net418));
 sg13g2_dlygate4sd3_1 hold170 (.A(_0042_),
    .X(net419));
 sg13g2_dlygate4sd3_1 hold171 (.A(\cell_cfg[8][2] ),
    .X(net420));
 sg13g2_dlygate4sd3_1 hold172 (.A(\cell_cfg[14][2] ),
    .X(net421));
 sg13g2_dlygate4sd3_1 hold173 (.A(\cell_cfg[30][2] ),
    .X(net422));
 sg13g2_dlygate4sd3_1 hold174 (.A(\cell_cfg[27][2] ),
    .X(net423));
 sg13g2_dlygate4sd3_1 hold175 (.A(_0125_),
    .X(net424));
 sg13g2_dlygate4sd3_1 hold176 (.A(\cell_cfg[12][0] ),
    .X(net425));
 sg13g2_dlygate4sd3_1 hold177 (.A(_0062_),
    .X(net426));
 sg13g2_dlygate4sd3_1 hold178 (.A(\cell_cfg[28][2] ),
    .X(net427));
 sg13g2_dlygate4sd3_1 hold179 (.A(\cell_cfg[23][2] ),
    .X(net428));
 sg13g2_dlygate4sd3_1 hold180 (.A(\cell_cfg[0][2] ),
    .X(net429));
 sg13g2_dlygate4sd3_1 hold181 (.A(_0272_),
    .X(net430));
 sg13g2_dlygate4sd3_1 hold182 (.A(\cell_cfg[31][2] ),
    .X(net431));
 sg13g2_dlygate4sd3_1 hold183 (.A(\cell_cfg[26][2] ),
    .X(net432));
 sg13g2_dlygate4sd3_1 hold184 (.A(_0129_),
    .X(net433));
 sg13g2_dlygate4sd3_1 hold185 (.A(\cell_cfg[3][0] ),
    .X(net434));
 sg13g2_dlygate4sd3_1 hold186 (.A(_0244_),
    .X(net435));
 sg13g2_dlygate4sd3_1 hold187 (.A(\cell_cfg[20][0] ),
    .X(net436));
 sg13g2_dlygate4sd3_1 hold188 (.A(\cell_cfg[21][2] ),
    .X(net437));
 sg13g2_dlygate4sd3_1 hold189 (.A(\cell_cfg[24][2] ),
    .X(net438));
 sg13g2_dlygate4sd3_1 hold190 (.A(\cell_cfg[15][2] ),
    .X(net439));
 sg13g2_dlygate4sd3_1 hold191 (.A(\cell_cfg[1][3] ),
    .X(net440));
 sg13g2_dlygate4sd3_1 hold192 (.A(_0100_),
    .X(net441));
 sg13g2_dlygate4sd3_1 hold193 (.A(\cell_cfg[25][2] ),
    .X(net442));
 sg13g2_dlygate4sd3_1 hold194 (.A(\cell_cfg[33][0] ),
    .X(net443));
 sg13g2_dlygate4sd3_1 hold195 (.A(_0783_),
    .X(net444));
 sg13g2_dlygate4sd3_1 hold196 (.A(\cell_cfg[10][2] ),
    .X(net445));
 sg13g2_dlygate4sd3_1 hold197 (.A(_0103_),
    .X(net446));
 sg13g2_dlygate4sd3_1 hold198 (.A(\cell_cfg[9][2] ),
    .X(net447));
 sg13g2_dlygate4sd3_1 hold199 (.A(\cell_cfg[10][3] ),
    .X(net448));
 sg13g2_dlygate4sd3_1 hold200 (.A(\cell_cfg[23][1] ),
    .X(net449));
 sg13g2_dlygate4sd3_1 hold201 (.A(\cell_cfg[5][0] ),
    .X(net450));
 sg13g2_dlygate4sd3_1 hold202 (.A(_0240_),
    .X(net451));
 sg13g2_dlygate4sd3_1 hold203 (.A(_0078_),
    .X(net452));
 sg13g2_dlygate4sd3_1 hold204 (.A(\cell_cfg[31][1] ),
    .X(net453));
 sg13g2_dlygate4sd3_1 hold205 (.A(_0025_),
    .X(net454));
 sg13g2_dlygate4sd3_1 hold206 (.A(\cell_cfg[21][1] ),
    .X(net455));
 sg13g2_dlygate4sd3_1 hold207 (.A(_0045_),
    .X(net456));
 sg13g2_dlygate4sd3_1 hold208 (.A(\cell_cfg[25][1] ),
    .X(net457));
 sg13g2_dlygate4sd3_1 hold209 (.A(_0037_),
    .X(net458));
 sg13g2_dlygate4sd3_1 hold210 (.A(\cell_cfg[35][1] ),
    .X(net459));
 sg13g2_dlygate4sd3_1 hold211 (.A(_0019_),
    .X(net460));
 sg13g2_dlygate4sd3_1 hold212 (.A(\cell_cfg[16][0] ),
    .X(net461));
 sg13g2_dlygate4sd3_1 hold213 (.A(_0168_),
    .X(net462));
 sg13g2_dlygate4sd3_1 hold214 (.A(\cell_cfg[22][1] ),
    .X(net463));
 sg13g2_dlygate4sd3_1 hold215 (.A(\cell_cfg[29][3] ),
    .X(net464));
 sg13g2_dlygate4sd3_1 hold216 (.A(\cell_cfg[12][1] ),
    .X(net465));
 sg13g2_dlygate4sd3_1 hold217 (.A(\cell_cfg[19][3] ),
    .X(net466));
 sg13g2_dlygate4sd3_1 hold218 (.A(_0017_),
    .X(net467));
 sg13g2_dlygate4sd3_1 hold219 (.A(\cell_cfg[24][3] ),
    .X(net468));
 sg13g2_dlygate4sd3_1 hold220 (.A(\cell_cfg[10][1] ),
    .X(net469));
 sg13g2_dlygate4sd3_1 hold221 (.A(\cell_cfg[0][1] ),
    .X(net470));
 sg13g2_dlygate4sd3_1 hold222 (.A(_0087_),
    .X(net471));
 sg13g2_dlygate4sd3_1 hold223 (.A(\cell_cfg[29][0] ),
    .X(net472));
 sg13g2_dlygate4sd3_1 hold224 (.A(\cell_cfg[27][1] ),
    .X(net473));
 sg13g2_dlygate4sd3_1 hold225 (.A(_0033_),
    .X(net474));
 sg13g2_dlygate4sd3_1 hold226 (.A(\cell_cfg[2][1] ),
    .X(net475));
 sg13g2_dlygate4sd3_1 hold227 (.A(\cell_cfg[2][3] ),
    .X(net476));
 sg13g2_dlygate4sd3_1 hold228 (.A(\cell_cfg[1][1] ),
    .X(net477));
 sg13g2_dlygate4sd3_1 hold229 (.A(\cell_cfg[34][0] ),
    .X(net478));
 sg13g2_dlygate4sd3_1 hold230 (.A(\cell_cfg[8][1] ),
    .X(net479));
 sg13g2_dlygate4sd3_1 hold231 (.A(\cell_cfg[32][2] ),
    .X(net480));
 sg13g2_dlygate4sd3_1 hold232 (.A(\cell_cfg[9][1] ),
    .X(net481));
 sg13g2_dlygate4sd3_1 hold233 (.A(\cell_cfg[4][3] ),
    .X(net482));
 sg13g2_dlygate4sd3_1 hold234 (.A(\cell_cfg[14][1] ),
    .X(net483));
 sg13g2_dlygate4sd3_1 hold235 (.A(\cell_cfg[18][1] ),
    .X(net484));
 sg13g2_dlygate4sd3_1 hold236 (.A(_0157_),
    .X(net485));
 sg13g2_dlygate4sd3_1 hold237 (.A(\cell_cfg[17][2] ),
    .X(net486));
 sg13g2_dlygate4sd3_1 hold238 (.A(\cell_cfg[5][1] ),
    .X(net487));
 sg13g2_dlygate4sd3_1 hold239 (.A(_0241_),
    .X(net488));
 sg13g2_dlygate4sd3_1 hold240 (.A(_0079_),
    .X(net489));
 sg13g2_dlygate4sd3_1 hold241 (.A(\cell_cfg[34][1] ),
    .X(net490));
 sg13g2_dlygate4sd3_1 hold242 (.A(\cell_cfg[24][0] ),
    .X(net491));
 sg13g2_dlygate4sd3_1 hold243 (.A(\cell_cfg[7][1] ),
    .X(net492));
 sg13g2_dlygate4sd3_1 hold244 (.A(_0073_),
    .X(net493));
 sg13g2_dlygate4sd3_1 hold245 (.A(\cell_cfg[0][3] ),
    .X(net494));
 sg13g2_dlygate4sd3_1 hold246 (.A(\cell_cfg[4][1] ),
    .X(net495));
 sg13g2_dlygate4sd3_1 hold247 (.A(_0246_),
    .X(net496));
 sg13g2_dlygate4sd3_1 hold248 (.A(\cell_cfg[26][1] ),
    .X(net497));
 sg13g2_dlygate4sd3_1 hold249 (.A(\cell_cfg[30][1] ),
    .X(net498));
 sg13g2_dlygate4sd3_1 hold250 (.A(\cell_cfg[17][1] ),
    .X(net499));
 sg13g2_dlygate4sd3_1 hold251 (.A(_0165_),
    .X(net500));
 sg13g2_dlygate4sd3_1 hold252 (.A(\cell_cfg[20][1] ),
    .X(net501));
 sg13g2_dlygate4sd3_1 hold253 (.A(\cell_cfg[6][1] ),
    .X(net502));
 sg13g2_dlygate4sd3_1 hold254 (.A(\cell_cfg[16][1] ),
    .X(net503));
 sg13g2_dlygate4sd3_1 hold255 (.A(_0169_),
    .X(net504));
 sg13g2_dlygate4sd3_1 hold256 (.A(\cell_cfg[28][0] ),
    .X(net505));
 sg13g2_dlygate4sd3_1 hold257 (.A(_0030_),
    .X(net506));
 sg13g2_dlygate4sd3_1 hold258 (.A(\cell_cfg[19][1] ),
    .X(net507));
 sg13g2_dlygate4sd3_1 hold259 (.A(\cell_cfg[28][1] ),
    .X(net508));
 sg13g2_dlygate4sd3_1 hold260 (.A(_0031_),
    .X(net509));
 sg13g2_dlygate4sd3_1 hold261 (.A(\cell_cfg[29][1] ),
    .X(net510));
 sg13g2_dlygate4sd3_1 hold262 (.A(\cell_cfg[23][0] ),
    .X(net511));
 sg13g2_dlygate4sd3_1 hold263 (.A(_0040_),
    .X(net512));
 sg13g2_dlygate4sd3_1 hold264 (.A(\cell_cfg[15][0] ),
    .X(net513));
 sg13g2_dlygate4sd3_1 hold265 (.A(\cell_cfg[15][1] ),
    .X(net514));
 sg13g2_dlygate4sd3_1 hold266 (.A(\cell_cfg[3][1] ),
    .X(net515));
 sg13g2_dlygate4sd3_1 hold267 (.A(\cell_cfg[27][3] ),
    .X(net516));
 sg13g2_dlygate4sd3_1 hold268 (.A(\cell_cfg[14][3] ),
    .X(net517));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_4 FILLER_5_42 ();
 sg13g2_decap_4 FILLER_5_50 ();
 sg13g2_fill_1 FILLER_5_54 ();
 sg13g2_fill_2 FILLER_5_59 ();
 sg13g2_decap_8 FILLER_5_65 ();
 sg13g2_decap_8 FILLER_5_72 ();
 sg13g2_decap_8 FILLER_5_79 ();
 sg13g2_decap_8 FILLER_5_86 ();
 sg13g2_decap_8 FILLER_5_93 ();
 sg13g2_decap_8 FILLER_5_100 ();
 sg13g2_decap_8 FILLER_5_107 ();
 sg13g2_decap_8 FILLER_5_114 ();
 sg13g2_decap_8 FILLER_5_121 ();
 sg13g2_decap_8 FILLER_5_128 ();
 sg13g2_decap_8 FILLER_5_135 ();
 sg13g2_decap_8 FILLER_5_142 ();
 sg13g2_decap_8 FILLER_5_149 ();
 sg13g2_decap_8 FILLER_5_156 ();
 sg13g2_decap_8 FILLER_5_163 ();
 sg13g2_decap_8 FILLER_5_170 ();
 sg13g2_decap_8 FILLER_5_177 ();
 sg13g2_decap_8 FILLER_5_184 ();
 sg13g2_decap_8 FILLER_5_191 ();
 sg13g2_decap_8 FILLER_5_198 ();
 sg13g2_decap_8 FILLER_5_205 ();
 sg13g2_decap_8 FILLER_5_212 ();
 sg13g2_decap_8 FILLER_5_219 ();
 sg13g2_decap_8 FILLER_5_226 ();
 sg13g2_decap_8 FILLER_5_233 ();
 sg13g2_decap_8 FILLER_5_240 ();
 sg13g2_decap_8 FILLER_5_247 ();
 sg13g2_decap_8 FILLER_5_254 ();
 sg13g2_decap_8 FILLER_5_261 ();
 sg13g2_fill_1 FILLER_5_268 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_fill_2 FILLER_6_35 ();
 sg13g2_fill_2 FILLER_6_55 ();
 sg13g2_fill_1 FILLER_6_57 ();
 sg13g2_fill_2 FILLER_6_110 ();
 sg13g2_decap_8 FILLER_6_116 ();
 sg13g2_decap_8 FILLER_6_123 ();
 sg13g2_decap_8 FILLER_6_130 ();
 sg13g2_decap_8 FILLER_6_137 ();
 sg13g2_decap_4 FILLER_6_144 ();
 sg13g2_fill_2 FILLER_6_148 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_4 FILLER_6_206 ();
 sg13g2_decap_8 FILLER_6_214 ();
 sg13g2_decap_8 FILLER_6_221 ();
 sg13g2_fill_1 FILLER_6_235 ();
 sg13g2_decap_8 FILLER_6_249 ();
 sg13g2_decap_4 FILLER_6_256 ();
 sg13g2_decap_8 FILLER_6_298 ();
 sg13g2_fill_2 FILLER_6_305 ();
 sg13g2_fill_1 FILLER_6_307 ();
 sg13g2_decap_8 FILLER_6_312 ();
 sg13g2_decap_8 FILLER_6_319 ();
 sg13g2_decap_8 FILLER_6_326 ();
 sg13g2_decap_8 FILLER_6_333 ();
 sg13g2_decap_8 FILLER_6_340 ();
 sg13g2_decap_8 FILLER_6_347 ();
 sg13g2_decap_8 FILLER_6_354 ();
 sg13g2_decap_8 FILLER_6_361 ();
 sg13g2_decap_8 FILLER_6_368 ();
 sg13g2_decap_8 FILLER_6_375 ();
 sg13g2_decap_8 FILLER_6_382 ();
 sg13g2_decap_8 FILLER_6_389 ();
 sg13g2_decap_8 FILLER_6_396 ();
 sg13g2_decap_4 FILLER_6_403 ();
 sg13g2_fill_2 FILLER_6_407 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_4 FILLER_7_14 ();
 sg13g2_fill_1 FILLER_7_70 ();
 sg13g2_fill_2 FILLER_7_88 ();
 sg13g2_fill_1 FILLER_7_94 ();
 sg13g2_fill_2 FILLER_7_99 ();
 sg13g2_decap_8 FILLER_7_127 ();
 sg13g2_fill_2 FILLER_7_134 ();
 sg13g2_fill_1 FILLER_7_188 ();
 sg13g2_fill_2 FILLER_7_270 ();
 sg13g2_fill_2 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_4 FILLER_8_14 ();
 sg13g2_fill_2 FILLER_8_57 ();
 sg13g2_fill_2 FILLER_8_113 ();
 sg13g2_fill_2 FILLER_8_123 ();
 sg13g2_fill_1 FILLER_8_125 ();
 sg13g2_fill_2 FILLER_8_146 ();
 sg13g2_fill_2 FILLER_8_218 ();
 sg13g2_decap_4 FILLER_8_224 ();
 sg13g2_fill_2 FILLER_8_228 ();
 sg13g2_decap_4 FILLER_8_233 ();
 sg13g2_fill_2 FILLER_8_246 ();
 sg13g2_fill_2 FILLER_8_274 ();
 sg13g2_fill_1 FILLER_8_276 ();
 sg13g2_decap_8 FILLER_8_334 ();
 sg13g2_decap_8 FILLER_8_341 ();
 sg13g2_decap_8 FILLER_8_348 ();
 sg13g2_decap_8 FILLER_8_355 ();
 sg13g2_decap_8 FILLER_8_362 ();
 sg13g2_decap_8 FILLER_8_369 ();
 sg13g2_decap_8 FILLER_8_376 ();
 sg13g2_decap_8 FILLER_8_383 ();
 sg13g2_decap_8 FILLER_8_390 ();
 sg13g2_decap_8 FILLER_8_397 ();
 sg13g2_decap_4 FILLER_8_404 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_4 FILLER_9_7 ();
 sg13g2_fill_2 FILLER_9_15 ();
 sg13g2_fill_2 FILLER_9_70 ();
 sg13g2_fill_1 FILLER_9_77 ();
 sg13g2_fill_2 FILLER_9_245 ();
 sg13g2_fill_2 FILLER_9_266 ();
 sg13g2_fill_1 FILLER_9_268 ();
 sg13g2_fill_1 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_347 ();
 sg13g2_decap_8 FILLER_9_354 ();
 sg13g2_decap_8 FILLER_9_361 ();
 sg13g2_decap_8 FILLER_9_368 ();
 sg13g2_decap_8 FILLER_9_375 ();
 sg13g2_decap_8 FILLER_9_382 ();
 sg13g2_decap_8 FILLER_9_389 ();
 sg13g2_decap_8 FILLER_9_396 ();
 sg13g2_decap_4 FILLER_9_403 ();
 sg13g2_fill_2 FILLER_9_407 ();
 sg13g2_fill_1 FILLER_10_0 ();
 sg13g2_fill_1 FILLER_10_36 ();
 sg13g2_fill_2 FILLER_10_60 ();
 sg13g2_fill_2 FILLER_10_72 ();
 sg13g2_fill_1 FILLER_10_79 ();
 sg13g2_fill_2 FILLER_10_102 ();
 sg13g2_fill_1 FILLER_10_104 ();
 sg13g2_fill_2 FILLER_10_149 ();
 sg13g2_fill_1 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_fill_1 FILLER_10_224 ();
 sg13g2_decap_4 FILLER_10_239 ();
 sg13g2_fill_2 FILLER_10_288 ();
 sg13g2_fill_1 FILLER_10_299 ();
 sg13g2_decap_4 FILLER_10_335 ();
 sg13g2_fill_2 FILLER_10_343 ();
 sg13g2_fill_1 FILLER_10_345 ();
 sg13g2_decap_8 FILLER_10_349 ();
 sg13g2_decap_8 FILLER_10_360 ();
 sg13g2_decap_8 FILLER_10_367 ();
 sg13g2_decap_8 FILLER_10_374 ();
 sg13g2_decap_8 FILLER_10_381 ();
 sg13g2_decap_8 FILLER_10_388 ();
 sg13g2_decap_8 FILLER_10_395 ();
 sg13g2_decap_8 FILLER_10_402 ();
 sg13g2_decap_4 FILLER_11_0 ();
 sg13g2_fill_1 FILLER_11_4 ();
 sg13g2_fill_2 FILLER_11_60 ();
 sg13g2_fill_2 FILLER_11_77 ();
 sg13g2_fill_1 FILLER_11_90 ();
 sg13g2_fill_2 FILLER_11_102 ();
 sg13g2_fill_1 FILLER_11_114 ();
 sg13g2_fill_2 FILLER_11_146 ();
 sg13g2_fill_2 FILLER_11_179 ();
 sg13g2_fill_2 FILLER_11_227 ();
 sg13g2_fill_2 FILLER_11_249 ();
 sg13g2_fill_1 FILLER_11_251 ();
 sg13g2_fill_2 FILLER_11_301 ();
 sg13g2_fill_1 FILLER_11_334 ();
 sg13g2_fill_1 FILLER_11_344 ();
 sg13g2_decap_4 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_387 ();
 sg13g2_decap_8 FILLER_11_394 ();
 sg13g2_decap_8 FILLER_11_401 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_fill_2 FILLER_12_35 ();
 sg13g2_fill_2 FILLER_12_83 ();
 sg13g2_fill_1 FILLER_12_85 ();
 sg13g2_fill_2 FILLER_12_97 ();
 sg13g2_decap_4 FILLER_12_122 ();
 sg13g2_fill_1 FILLER_12_126 ();
 sg13g2_fill_1 FILLER_12_141 ();
 sg13g2_fill_1 FILLER_12_164 ();
 sg13g2_fill_2 FILLER_12_178 ();
 sg13g2_fill_1 FILLER_12_195 ();
 sg13g2_decap_8 FILLER_12_216 ();
 sg13g2_decap_8 FILLER_12_223 ();
 sg13g2_decap_4 FILLER_12_230 ();
 sg13g2_fill_1 FILLER_12_234 ();
 sg13g2_fill_2 FILLER_12_252 ();
 sg13g2_fill_1 FILLER_12_254 ();
 sg13g2_fill_2 FILLER_12_264 ();
 sg13g2_fill_1 FILLER_12_266 ();
 sg13g2_fill_2 FILLER_12_285 ();
 sg13g2_fill_1 FILLER_12_287 ();
 sg13g2_fill_1 FILLER_12_307 ();
 sg13g2_fill_2 FILLER_12_317 ();
 sg13g2_decap_4 FILLER_12_396 ();
 sg13g2_decap_4 FILLER_13_0 ();
 sg13g2_fill_2 FILLER_13_39 ();
 sg13g2_fill_1 FILLER_13_41 ();
 sg13g2_fill_2 FILLER_13_76 ();
 sg13g2_fill_1 FILLER_13_78 ();
 sg13g2_decap_4 FILLER_13_112 ();
 sg13g2_fill_2 FILLER_13_121 ();
 sg13g2_fill_2 FILLER_13_159 ();
 sg13g2_decap_4 FILLER_13_226 ();
 sg13g2_fill_1 FILLER_13_230 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_fill_1 FILLER_13_245 ();
 sg13g2_fill_2 FILLER_13_260 ();
 sg13g2_fill_1 FILLER_13_262 ();
 sg13g2_fill_2 FILLER_13_294 ();
 sg13g2_fill_1 FILLER_13_335 ();
 sg13g2_fill_1 FILLER_13_393 ();
 sg13g2_decap_4 FILLER_13_403 ();
 sg13g2_fill_2 FILLER_13_407 ();
 sg13g2_decap_4 FILLER_14_0 ();
 sg13g2_fill_2 FILLER_14_4 ();
 sg13g2_fill_2 FILLER_14_39 ();
 sg13g2_fill_1 FILLER_14_50 ();
 sg13g2_decap_8 FILLER_14_81 ();
 sg13g2_fill_2 FILLER_14_88 ();
 sg13g2_fill_1 FILLER_14_153 ();
 sg13g2_fill_2 FILLER_14_164 ();
 sg13g2_fill_1 FILLER_14_166 ();
 sg13g2_fill_1 FILLER_14_175 ();
 sg13g2_fill_1 FILLER_14_193 ();
 sg13g2_fill_2 FILLER_14_199 ();
 sg13g2_fill_1 FILLER_14_206 ();
 sg13g2_fill_1 FILLER_14_219 ();
 sg13g2_fill_2 FILLER_14_265 ();
 sg13g2_fill_1 FILLER_14_286 ();
 sg13g2_fill_1 FILLER_14_344 ();
 sg13g2_fill_1 FILLER_14_380 ();
 sg13g2_fill_2 FILLER_14_407 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_fill_1 FILLER_15_91 ();
 sg13g2_fill_2 FILLER_15_109 ();
 sg13g2_fill_1 FILLER_15_111 ();
 sg13g2_decap_4 FILLER_15_134 ();
 sg13g2_fill_1 FILLER_15_155 ();
 sg13g2_fill_2 FILLER_15_163 ();
 sg13g2_fill_1 FILLER_15_254 ();
 sg13g2_fill_1 FILLER_15_284 ();
 sg13g2_fill_2 FILLER_15_348 ();
 sg13g2_fill_1 FILLER_15_381 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_4 FILLER_16_0 ();
 sg13g2_fill_1 FILLER_16_4 ();
 sg13g2_fill_1 FILLER_16_70 ();
 sg13g2_fill_1 FILLER_16_76 ();
 sg13g2_fill_1 FILLER_16_103 ();
 sg13g2_fill_2 FILLER_16_143 ();
 sg13g2_fill_1 FILLER_16_192 ();
 sg13g2_fill_1 FILLER_16_271 ();
 sg13g2_fill_2 FILLER_16_278 ();
 sg13g2_decap_4 FILLER_16_290 ();
 sg13g2_decap_4 FILLER_16_300 ();
 sg13g2_fill_1 FILLER_16_304 ();
 sg13g2_fill_2 FILLER_16_321 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_fill_1 FILLER_17_0 ();
 sg13g2_fill_1 FILLER_17_31 ();
 sg13g2_decap_8 FILLER_17_104 ();
 sg13g2_decap_4 FILLER_17_111 ();
 sg13g2_decap_4 FILLER_17_119 ();
 sg13g2_fill_1 FILLER_17_123 ();
 sg13g2_fill_1 FILLER_17_145 ();
 sg13g2_fill_2 FILLER_17_235 ();
 sg13g2_fill_1 FILLER_17_237 ();
 sg13g2_decap_4 FILLER_17_306 ();
 sg13g2_fill_2 FILLER_17_341 ();
 sg13g2_fill_2 FILLER_17_363 ();
 sg13g2_fill_2 FILLER_17_370 ();
 sg13g2_fill_1 FILLER_17_372 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_fill_1 FILLER_18_26 ();
 sg13g2_fill_1 FILLER_18_46 ();
 sg13g2_fill_1 FILLER_18_69 ();
 sg13g2_decap_4 FILLER_18_100 ();
 sg13g2_fill_1 FILLER_18_130 ();
 sg13g2_fill_2 FILLER_18_220 ();
 sg13g2_fill_1 FILLER_18_222 ();
 sg13g2_decap_8 FILLER_18_240 ();
 sg13g2_fill_1 FILLER_18_247 ();
 sg13g2_fill_1 FILLER_18_252 ();
 sg13g2_decap_8 FILLER_18_276 ();
 sg13g2_fill_2 FILLER_18_283 ();
 sg13g2_decap_8 FILLER_18_289 ();
 sg13g2_decap_8 FILLER_18_296 ();
 sg13g2_fill_1 FILLER_18_303 ();
 sg13g2_decap_8 FILLER_18_314 ();
 sg13g2_fill_1 FILLER_18_321 ();
 sg13g2_fill_1 FILLER_18_327 ();
 sg13g2_fill_2 FILLER_18_355 ();
 sg13g2_fill_1 FILLER_18_357 ();
 sg13g2_decap_4 FILLER_18_404 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_decap_4 FILLER_19_0 ();
 sg13g2_fill_1 FILLER_19_4 ();
 sg13g2_fill_2 FILLER_19_22 ();
 sg13g2_fill_1 FILLER_19_24 ();
 sg13g2_fill_1 FILLER_19_30 ();
 sg13g2_fill_2 FILLER_19_67 ();
 sg13g2_fill_1 FILLER_19_69 ();
 sg13g2_fill_1 FILLER_19_75 ();
 sg13g2_fill_2 FILLER_19_81 ();
 sg13g2_fill_2 FILLER_19_97 ();
 sg13g2_decap_4 FILLER_19_107 ();
 sg13g2_fill_1 FILLER_19_111 ();
 sg13g2_fill_2 FILLER_19_116 ();
 sg13g2_fill_1 FILLER_19_118 ();
 sg13g2_fill_2 FILLER_19_159 ();
 sg13g2_fill_1 FILLER_19_216 ();
 sg13g2_fill_2 FILLER_19_260 ();
 sg13g2_fill_1 FILLER_19_314 ();
 sg13g2_fill_1 FILLER_19_334 ();
 sg13g2_fill_1 FILLER_19_343 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_fill_1 FILLER_20_0 ();
 sg13g2_fill_1 FILLER_20_44 ();
 sg13g2_fill_2 FILLER_20_58 ();
 sg13g2_fill_1 FILLER_20_65 ();
 sg13g2_fill_2 FILLER_20_92 ();
 sg13g2_fill_2 FILLER_20_109 ();
 sg13g2_fill_1 FILLER_20_129 ();
 sg13g2_fill_1 FILLER_20_134 ();
 sg13g2_decap_4 FILLER_20_139 ();
 sg13g2_fill_2 FILLER_20_176 ();
 sg13g2_fill_2 FILLER_20_183 ();
 sg13g2_fill_2 FILLER_20_190 ();
 sg13g2_decap_8 FILLER_20_206 ();
 sg13g2_decap_8 FILLER_20_213 ();
 sg13g2_decap_4 FILLER_20_220 ();
 sg13g2_fill_1 FILLER_20_224 ();
 sg13g2_decap_8 FILLER_20_234 ();
 sg13g2_decap_8 FILLER_20_241 ();
 sg13g2_fill_1 FILLER_20_248 ();
 sg13g2_decap_4 FILLER_20_269 ();
 sg13g2_decap_4 FILLER_20_277 ();
 sg13g2_fill_2 FILLER_20_281 ();
 sg13g2_fill_2 FILLER_20_315 ();
 sg13g2_fill_1 FILLER_20_326 ();
 sg13g2_fill_2 FILLER_20_354 ();
 sg13g2_fill_2 FILLER_20_365 ();
 sg13g2_fill_1 FILLER_20_367 ();
 sg13g2_fill_2 FILLER_20_373 ();
 sg13g2_fill_1 FILLER_20_375 ();
 sg13g2_fill_2 FILLER_20_385 ();
 sg13g2_fill_1 FILLER_20_387 ();
 sg13g2_decap_4 FILLER_20_405 ();
 sg13g2_decap_4 FILLER_21_0 ();
 sg13g2_fill_1 FILLER_21_4 ();
 sg13g2_fill_2 FILLER_21_45 ();
 sg13g2_fill_1 FILLER_21_47 ();
 sg13g2_fill_1 FILLER_21_80 ();
 sg13g2_fill_2 FILLER_21_113 ();
 sg13g2_fill_1 FILLER_21_124 ();
 sg13g2_decap_8 FILLER_21_135 ();
 sg13g2_decap_4 FILLER_21_142 ();
 sg13g2_fill_1 FILLER_21_156 ();
 sg13g2_fill_2 FILLER_21_165 ();
 sg13g2_decap_8 FILLER_21_211 ();
 sg13g2_fill_1 FILLER_21_218 ();
 sg13g2_fill_2 FILLER_21_249 ();
 sg13g2_fill_1 FILLER_21_251 ();
 sg13g2_fill_2 FILLER_21_258 ();
 sg13g2_fill_1 FILLER_21_279 ();
 sg13g2_fill_1 FILLER_21_318 ();
 sg13g2_fill_2 FILLER_21_333 ();
 sg13g2_fill_1 FILLER_21_335 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_4 FILLER_22_7 ();
 sg13g2_fill_1 FILLER_22_24 ();
 sg13g2_fill_2 FILLER_22_65 ();
 sg13g2_fill_1 FILLER_22_107 ();
 sg13g2_fill_2 FILLER_22_160 ();
 sg13g2_fill_1 FILLER_22_202 ();
 sg13g2_fill_1 FILLER_22_238 ();
 sg13g2_fill_2 FILLER_22_274 ();
 sg13g2_decap_4 FILLER_22_291 ();
 sg13g2_fill_1 FILLER_22_339 ();
 sg13g2_fill_1 FILLER_22_345 ();
 sg13g2_fill_1 FILLER_22_363 ();
 sg13g2_fill_1 FILLER_23_35 ();
 sg13g2_fill_1 FILLER_23_40 ();
 sg13g2_fill_1 FILLER_23_57 ();
 sg13g2_fill_1 FILLER_23_65 ();
 sg13g2_decap_4 FILLER_23_81 ();
 sg13g2_fill_1 FILLER_23_90 ();
 sg13g2_decap_4 FILLER_23_159 ();
 sg13g2_fill_2 FILLER_23_163 ();
 sg13g2_fill_1 FILLER_23_170 ();
 sg13g2_fill_1 FILLER_23_176 ();
 sg13g2_decap_8 FILLER_23_198 ();
 sg13g2_fill_1 FILLER_23_205 ();
 sg13g2_decap_8 FILLER_23_211 ();
 sg13g2_decap_4 FILLER_23_218 ();
 sg13g2_fill_2 FILLER_23_222 ();
 sg13g2_decap_8 FILLER_23_236 ();
 sg13g2_fill_1 FILLER_23_248 ();
 sg13g2_decap_4 FILLER_23_254 ();
 sg13g2_fill_1 FILLER_23_266 ();
 sg13g2_decap_4 FILLER_23_316 ();
 sg13g2_fill_1 FILLER_23_320 ();
 sg13g2_fill_2 FILLER_23_344 ();
 sg13g2_fill_1 FILLER_23_382 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_fill_1 FILLER_24_7 ();
 sg13g2_fill_1 FILLER_24_106 ();
 sg13g2_decap_8 FILLER_24_182 ();
 sg13g2_decap_8 FILLER_24_189 ();
 sg13g2_fill_2 FILLER_24_196 ();
 sg13g2_fill_2 FILLER_24_211 ();
 sg13g2_fill_2 FILLER_24_239 ();
 sg13g2_fill_2 FILLER_24_255 ();
 sg13g2_decap_4 FILLER_24_271 ();
 sg13g2_fill_2 FILLER_24_275 ();
 sg13g2_fill_1 FILLER_24_295 ();
 sg13g2_decap_8 FILLER_24_351 ();
 sg13g2_fill_2 FILLER_24_366 ();
 sg13g2_fill_2 FILLER_24_372 ();
 sg13g2_fill_2 FILLER_25_26 ();
 sg13g2_fill_1 FILLER_25_42 ();
 sg13g2_fill_2 FILLER_25_79 ();
 sg13g2_fill_2 FILLER_25_92 ();
 sg13g2_fill_1 FILLER_25_141 ();
 sg13g2_decap_8 FILLER_25_151 ();
 sg13g2_fill_2 FILLER_25_158 ();
 sg13g2_fill_2 FILLER_25_168 ();
 sg13g2_fill_1 FILLER_25_170 ();
 sg13g2_fill_2 FILLER_25_180 ();
 sg13g2_fill_1 FILLER_25_182 ();
 sg13g2_decap_8 FILLER_25_214 ();
 sg13g2_fill_1 FILLER_25_221 ();
 sg13g2_fill_1 FILLER_25_248 ();
 sg13g2_fill_2 FILLER_25_270 ();
 sg13g2_fill_1 FILLER_25_297 ();
 sg13g2_fill_2 FILLER_26_0 ();
 sg13g2_fill_1 FILLER_26_2 ();
 sg13g2_fill_2 FILLER_26_46 ();
 sg13g2_fill_1 FILLER_26_57 ();
 sg13g2_fill_2 FILLER_26_68 ();
 sg13g2_fill_1 FILLER_26_75 ();
 sg13g2_fill_2 FILLER_26_103 ();
 sg13g2_fill_1 FILLER_26_114 ();
 sg13g2_fill_2 FILLER_26_130 ();
 sg13g2_decap_8 FILLER_26_220 ();
 sg13g2_fill_1 FILLER_26_312 ();
 sg13g2_fill_2 FILLER_26_319 ();
 sg13g2_fill_1 FILLER_26_382 ();
 sg13g2_fill_2 FILLER_27_63 ();
 sg13g2_fill_2 FILLER_27_122 ();
 sg13g2_fill_2 FILLER_27_138 ();
 sg13g2_fill_1 FILLER_27_155 ();
 sg13g2_fill_2 FILLER_27_222 ();
 sg13g2_fill_1 FILLER_27_224 ();
 sg13g2_fill_1 FILLER_27_255 ();
 sg13g2_fill_2 FILLER_27_310 ();
 sg13g2_fill_1 FILLER_27_350 ();
 sg13g2_fill_2 FILLER_27_373 ();
 sg13g2_fill_1 FILLER_27_408 ();
 sg13g2_fill_1 FILLER_28_0 ();
 sg13g2_fill_2 FILLER_28_27 ();
 sg13g2_fill_1 FILLER_28_58 ();
 sg13g2_fill_1 FILLER_28_102 ();
 sg13g2_fill_2 FILLER_28_117 ();
 sg13g2_fill_2 FILLER_28_129 ();
 sg13g2_fill_1 FILLER_28_131 ();
 sg13g2_fill_2 FILLER_28_158 ();
 sg13g2_fill_1 FILLER_28_160 ();
 sg13g2_fill_2 FILLER_28_169 ();
 sg13g2_fill_1 FILLER_28_171 ();
 sg13g2_fill_2 FILLER_28_212 ();
 sg13g2_decap_4 FILLER_28_223 ();
 sg13g2_fill_1 FILLER_28_253 ();
 sg13g2_fill_1 FILLER_28_269 ();
 sg13g2_fill_2 FILLER_28_294 ();
 sg13g2_fill_2 FILLER_28_320 ();
 sg13g2_fill_2 FILLER_29_77 ();
 sg13g2_fill_1 FILLER_29_79 ();
 sg13g2_fill_1 FILLER_29_88 ();
 sg13g2_fill_2 FILLER_29_137 ();
 sg13g2_fill_1 FILLER_29_139 ();
 sg13g2_fill_2 FILLER_29_145 ();
 sg13g2_fill_1 FILLER_29_147 ();
 sg13g2_fill_2 FILLER_29_175 ();
 sg13g2_fill_1 FILLER_29_177 ();
 sg13g2_fill_2 FILLER_29_218 ();
 sg13g2_fill_2 FILLER_29_232 ();
 sg13g2_fill_1 FILLER_29_234 ();
 sg13g2_fill_1 FILLER_29_323 ();
 sg13g2_fill_2 FILLER_29_333 ();
 sg13g2_fill_1 FILLER_29_373 ();
 sg13g2_fill_2 FILLER_30_0 ();
 sg13g2_fill_2 FILLER_30_26 ();
 sg13g2_fill_2 FILLER_30_73 ();
 sg13g2_fill_1 FILLER_30_112 ();
 sg13g2_decap_4 FILLER_30_128 ();
 sg13g2_fill_2 FILLER_30_137 ();
 sg13g2_fill_1 FILLER_30_144 ();
 sg13g2_decap_4 FILLER_30_150 ();
 sg13g2_fill_1 FILLER_30_176 ();
 sg13g2_fill_1 FILLER_30_204 ();
 sg13g2_decap_4 FILLER_30_226 ();
 sg13g2_fill_1 FILLER_30_230 ();
 sg13g2_decap_8 FILLER_30_235 ();
 sg13g2_fill_1 FILLER_30_242 ();
 sg13g2_fill_1 FILLER_30_261 ();
 sg13g2_fill_2 FILLER_30_286 ();
 sg13g2_fill_1 FILLER_30_288 ();
 sg13g2_decap_4 FILLER_30_300 ();
 sg13g2_fill_2 FILLER_30_319 ();
 sg13g2_fill_1 FILLER_31_26 ();
 sg13g2_fill_2 FILLER_31_63 ();
 sg13g2_fill_1 FILLER_31_74 ();
 sg13g2_fill_1 FILLER_31_132 ();
 sg13g2_fill_2 FILLER_31_189 ();
 sg13g2_fill_1 FILLER_31_191 ();
 sg13g2_fill_1 FILLER_31_197 ();
 sg13g2_decap_8 FILLER_31_219 ();
 sg13g2_decap_4 FILLER_31_226 ();
 sg13g2_fill_1 FILLER_31_230 ();
 sg13g2_fill_2 FILLER_31_251 ();
 sg13g2_fill_1 FILLER_31_253 ();
 sg13g2_fill_2 FILLER_31_282 ();
 sg13g2_fill_1 FILLER_31_284 ();
 sg13g2_decap_8 FILLER_31_290 ();
 sg13g2_fill_2 FILLER_31_311 ();
 sg13g2_fill_1 FILLER_31_337 ();
 sg13g2_fill_1 FILLER_31_343 ();
 sg13g2_fill_1 FILLER_31_350 ();
 sg13g2_fill_2 FILLER_31_365 ();
 sg13g2_fill_2 FILLER_31_372 ();
 sg13g2_fill_1 FILLER_32_0 ();
 sg13g2_fill_1 FILLER_32_41 ();
 sg13g2_fill_2 FILLER_32_149 ();
 sg13g2_fill_1 FILLER_32_151 ();
 sg13g2_decap_4 FILLER_32_160 ();
 sg13g2_fill_1 FILLER_32_164 ();
 sg13g2_fill_2 FILLER_32_174 ();
 sg13g2_fill_2 FILLER_32_224 ();
 sg13g2_fill_1 FILLER_32_226 ();
 sg13g2_fill_2 FILLER_32_253 ();
 sg13g2_fill_1 FILLER_32_255 ();
 sg13g2_fill_1 FILLER_32_271 ();
 sg13g2_fill_2 FILLER_32_313 ();
 sg13g2_fill_2 FILLER_32_331 ();
 sg13g2_fill_1 FILLER_33_97 ();
 sg13g2_fill_1 FILLER_33_131 ();
 sg13g2_fill_2 FILLER_33_155 ();
 sg13g2_fill_2 FILLER_33_176 ();
 sg13g2_decap_4 FILLER_33_228 ();
 sg13g2_fill_1 FILLER_33_232 ();
 sg13g2_fill_2 FILLER_33_247 ();
 sg13g2_fill_1 FILLER_33_249 ();
 sg13g2_fill_2 FILLER_33_260 ();
 sg13g2_fill_2 FILLER_33_276 ();
 sg13g2_fill_1 FILLER_33_278 ();
 sg13g2_fill_1 FILLER_33_397 ();
 sg13g2_fill_2 FILLER_33_406 ();
 sg13g2_fill_1 FILLER_33_408 ();
 sg13g2_fill_1 FILLER_34_0 ();
 sg13g2_fill_2 FILLER_34_18 ();
 sg13g2_fill_1 FILLER_34_20 ();
 sg13g2_fill_1 FILLER_34_66 ();
 sg13g2_fill_1 FILLER_34_81 ();
 sg13g2_fill_1 FILLER_34_92 ();
 sg13g2_fill_1 FILLER_34_146 ();
 sg13g2_fill_2 FILLER_34_169 ();
 sg13g2_fill_2 FILLER_34_190 ();
 sg13g2_fill_1 FILLER_34_202 ();
 sg13g2_decap_4 FILLER_34_221 ();
 sg13g2_fill_1 FILLER_34_225 ();
 sg13g2_fill_2 FILLER_34_319 ();
 sg13g2_fill_1 FILLER_34_321 ();
 sg13g2_fill_2 FILLER_34_327 ();
 sg13g2_fill_1 FILLER_34_329 ();
 sg13g2_fill_1 FILLER_34_339 ();
 sg13g2_fill_2 FILLER_34_349 ();
 sg13g2_fill_2 FILLER_34_365 ();
 sg13g2_fill_2 FILLER_34_381 ();
 sg13g2_fill_1 FILLER_35_35 ();
 sg13g2_fill_1 FILLER_35_45 ();
 sg13g2_fill_1 FILLER_35_76 ();
 sg13g2_fill_2 FILLER_35_217 ();
 sg13g2_fill_1 FILLER_35_249 ();
 sg13g2_fill_1 FILLER_35_258 ();
 sg13g2_fill_1 FILLER_35_322 ();
 sg13g2_fill_1 FILLER_35_354 ();
 sg13g2_fill_2 FILLER_35_406 ();
 sg13g2_fill_1 FILLER_35_408 ();
 sg13g2_decap_4 FILLER_36_0 ();
 sg13g2_fill_2 FILLER_36_47 ();
 sg13g2_fill_1 FILLER_36_49 ();
 sg13g2_fill_2 FILLER_36_160 ();
 sg13g2_fill_2 FILLER_36_180 ();
 sg13g2_fill_1 FILLER_36_182 ();
 sg13g2_decap_8 FILLER_36_235 ();
 sg13g2_fill_1 FILLER_36_242 ();
 sg13g2_fill_1 FILLER_36_339 ();
 sg13g2_fill_2 FILLER_36_348 ();
 sg13g2_fill_1 FILLER_36_350 ();
 sg13g2_fill_1 FILLER_36_382 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_fill_1 FILLER_37_14 ();
 sg13g2_fill_2 FILLER_37_203 ();
 sg13g2_decap_4 FILLER_37_218 ();
 sg13g2_fill_2 FILLER_37_313 ();
 sg13g2_fill_1 FILLER_37_315 ();
 sg13g2_fill_1 FILLER_37_338 ();
 sg13g2_fill_2 FILLER_37_406 ();
 sg13g2_fill_1 FILLER_37_408 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_4 FILLER_38_21 ();
 sg13g2_fill_1 FILLER_38_46 ();
 sg13g2_fill_2 FILLER_38_101 ();
 sg13g2_fill_2 FILLER_38_138 ();
 sg13g2_fill_1 FILLER_38_153 ();
 sg13g2_fill_2 FILLER_38_166 ();
 sg13g2_fill_2 FILLER_38_176 ();
 sg13g2_fill_1 FILLER_38_178 ();
 sg13g2_fill_2 FILLER_38_192 ();
 sg13g2_decap_4 FILLER_38_228 ();
 sg13g2_fill_1 FILLER_38_232 ();
 sg13g2_fill_2 FILLER_38_241 ();
 sg13g2_fill_2 FILLER_38_256 ();
 sg13g2_fill_1 FILLER_38_258 ();
 sg13g2_fill_1 FILLER_38_271 ();
 sg13g2_fill_2 FILLER_38_317 ();
 assign uio_oe[0] = net6;
 assign uio_oe[1] = net7;
 assign uio_oe[2] = net8;
 assign uio_oe[3] = net9;
 assign uio_oe[4] = net10;
 assign uio_oe[5] = net11;
 assign uio_oe[6] = net12;
 assign uio_oe[7] = net13;
 assign uio_out[0] = net14;
 assign uio_out[1] = net15;
 assign uio_out[2] = net16;
 assign uio_out[3] = net17;
 assign uio_out[4] = net18;
 assign uio_out[5] = net19;
 assign uio_out[6] = net20;
 assign uio_out[7] = net21;
 assign uo_out[0] = net22;
 assign uo_out[1] = net23;
 assign uo_out[2] = net24;
 assign uo_out[3] = net25;
endmodule

module tt_um_kch_cd101 (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire clknet_0_clk;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire data;
 wire \stop.adsr_ai[0] ;
 wire \stop.adsr_ai[1] ;
 wire \stop.adsr_ai[2] ;
 wire \stop.adsr_ai[3] ;
 wire \stop.adsr_ai[4] ;
 wire \stop.adsr_ai[5] ;
 wire \stop.adsr_ai[6] ;
 wire \stop.adsr_ai[7] ;
 wire \stop.adsr_di[0] ;
 wire \stop.adsr_di[1] ;
 wire \stop.adsr_di[2] ;
 wire \stop.adsr_di[3] ;
 wire \stop.adsr_di[4] ;
 wire \stop.adsr_di[5] ;
 wire \stop.adsr_di[6] ;
 wire \stop.adsr_di[7] ;
 wire \stop.adsr_ri[0] ;
 wire \stop.adsr_ri[1] ;
 wire \stop.adsr_ri[2] ;
 wire \stop.adsr_ri[3] ;
 wire \stop.adsr_ri[4] ;
 wire \stop.adsr_ri[5] ;
 wire \stop.adsr_ri[6] ;
 wire \stop.adsr_ri[7] ;
 wire \stop.adsr_s[0] ;
 wire \stop.adsr_s[1] ;
 wire \stop.adsr_s[2] ;
 wire \stop.adsr_s[3] ;
 wire \stop.adsr_s[4] ;
 wire \stop.adsr_s[5] ;
 wire \stop.adsr_s[6] ;
 wire \stop.adsr_s[7] ;
 wire \stop.ctrl.cfg[32] ;
 wire \stop.ctrl.cfg[33] ;
 wire \stop.ctrl.cfg[34] ;
 wire \stop.ctrl.cfg[35] ;
 wire \stop.ctrl.cfg[36] ;
 wire \stop.ctrl.cfg[37] ;
 wire \stop.ctrl.cfg[38] ;
 wire \stop.ctrl.cfg[39] ;
 wire \stop.ctrl.cfg[40] ;
 wire \stop.ctrl.cfg[41] ;
 wire \stop.ctrl.cfg[42] ;
 wire \stop.ctrl.cfg[43] ;
 wire \stop.ctrl.cfg[44] ;
 wire \stop.ctrl.cfg[45] ;
 wire \stop.ctrl.cfg[46] ;
 wire \stop.ctrl.cfg[47] ;
 wire \stop.ctrl.cfg[48] ;
 wire \stop.ctrl.cfg[49] ;
 wire \stop.ctrl.cfg[50] ;
 wire \stop.ctrl.cfg[51] ;
 wire \stop.ctrl.cfg[52] ;
 wire \stop.ctrl.cfg[53] ;
 wire \stop.ctrl.cfg[54] ;
 wire \stop.ctrl.cfg[55] ;
 wire \stop.ctrl.cfg[56] ;
 wire \stop.ctrl.cfg[57] ;
 wire \stop.ctrl.cfg[58] ;
 wire \stop.ctrl.cfg[59] ;
 wire \stop.ctrl.first_bit ;
 wire \stop.ctrl.first_bit_reg ;
 wire \stop.ctrl.trig ;
 wire \stop.merge_rstn ;
 wire \stop.merge_trig ;
 wire \stop.syn.adsr_data[0] ;
 wire \stop.syn.adsr_data[10] ;
 wire \stop.syn.adsr_data[11] ;
 wire \stop.syn.adsr_data[12] ;
 wire \stop.syn.adsr_data[13] ;
 wire \stop.syn.adsr_data[14] ;
 wire \stop.syn.adsr_data[15] ;
 wire \stop.syn.adsr_data[1] ;
 wire \stop.syn.adsr_data[2] ;
 wire \stop.syn.adsr_data[3] ;
 wire \stop.syn.adsr_data[4] ;
 wire \stop.syn.adsr_data[5] ;
 wire \stop.syn.adsr_data[6] ;
 wire \stop.syn.adsr_data[7] ;
 wire \stop.syn.adsr_data[8] ;
 wire \stop.syn.adsr_data[9] ;
 wire \stop.syn.adsr_data_reg[0] ;
 wire \stop.syn.adsr_data_reg[10] ;
 wire \stop.syn.adsr_data_reg[11] ;
 wire \stop.syn.adsr_data_reg[12] ;
 wire \stop.syn.adsr_data_reg[13] ;
 wire \stop.syn.adsr_data_reg[14] ;
 wire \stop.syn.adsr_data_reg[15] ;
 wire \stop.syn.adsr_data_reg[1] ;
 wire \stop.syn.adsr_data_reg[2] ;
 wire \stop.syn.adsr_data_reg[3] ;
 wire \stop.syn.adsr_data_reg[4] ;
 wire \stop.syn.adsr_data_reg[5] ;
 wire \stop.syn.adsr_data_reg[6] ;
 wire \stop.syn.adsr_data_reg[7] ;
 wire \stop.syn.adsr_data_reg[8] ;
 wire \stop.syn.adsr_data_reg[9] ;
 wire \stop.syn.adsri.clk ;
 wire \stop.syn.adsri.envelope[0] ;
 wire \stop.syn.adsri.envelope[1] ;
 wire \stop.syn.adsri.envelope[2] ;
 wire \stop.syn.adsri.envelope[3] ;
 wire \stop.syn.adsri.envelope[4] ;
 wire \stop.syn.adsri.envelope[5] ;
 wire \stop.syn.adsri.envelope[6] ;
 wire \stop.syn.adsri.envelope[7] ;
 wire \stop.syn.adsri.rstn ;
 wire \stop.syn.adsri.state[0] ;
 wire \stop.syn.adsri.state[1] ;
 wire \stop.syn.adsri.state[2] ;
 wire \stop.syn.adsri.state[3] ;
 wire \stop.syn.adsri.state[4] ;
 wire \stop.syn.adsri.trig ;
 wire \stop.syn.clk_mult ;
 wire \stop.syn.clk_sample ;
 wire \stop.syn.clk_sample_x2 ;
 wire \stop.syn.clki.arstn ;
 wire \stop.syn.clki.gen[0].inst.q ;
 wire \stop.syn.clki.gen[10].inst.clk ;
 wire \stop.syn.clki.gen[10].inst.q ;
 wire \stop.syn.clki.gen[11].inst.q ;
 wire \stop.syn.clki.gen[12].inst.q ;
 wire \stop.syn.clki.gen[13].inst.q ;
 wire \stop.syn.clki.gen[14].inst.q ;
 wire \stop.syn.clki.gen[1].inst.q ;
 wire \stop.syn.clki.gen[2].inst.q ;
 wire \stop.syn.clki.gen[3].inst.q ;
 wire \stop.syn.clki.gen[5].inst.q ;
 wire \stop.syn.clki.gen[6].inst.q ;
 wire \stop.syn.daci.accumulator[0] ;
 wire \stop.syn.daci.accumulator[10] ;
 wire \stop.syn.daci.accumulator[11] ;
 wire \stop.syn.daci.accumulator[12] ;
 wire \stop.syn.daci.accumulator[13] ;
 wire \stop.syn.daci.accumulator[14] ;
 wire \stop.syn.daci.accumulator[15] ;
 wire \stop.syn.daci.accumulator[1] ;
 wire \stop.syn.daci.accumulator[2] ;
 wire \stop.syn.daci.accumulator[3] ;
 wire \stop.syn.daci.accumulator[4] ;
 wire \stop.syn.daci.accumulator[5] ;
 wire \stop.syn.daci.accumulator[6] ;
 wire \stop.syn.daci.accumulator[7] ;
 wire \stop.syn.daci.accumulator[8] ;
 wire \stop.syn.daci.accumulator[9] ;
 wire \stop.syn.daci.din[0] ;
 wire \stop.syn.daci.din[10] ;
 wire \stop.syn.daci.din[11] ;
 wire \stop.syn.daci.din[12] ;
 wire \stop.syn.daci.din[13] ;
 wire \stop.syn.daci.din[14] ;
 wire \stop.syn.daci.din[15] ;
 wire \stop.syn.daci.din[1] ;
 wire \stop.syn.daci.din[2] ;
 wire \stop.syn.daci.din[3] ;
 wire \stop.syn.daci.din[4] ;
 wire \stop.syn.daci.din[5] ;
 wire \stop.syn.daci.din[6] ;
 wire \stop.syn.daci.din[7] ;
 wire \stop.syn.daci.din[8] ;
 wire \stop.syn.daci.din[9] ;
 wire \stop.syn.filt.m1.b_bit ;
 wire \stop.syn.filt.m1.b_latched[1] ;
 wire \stop.syn.filt.m1.b_latched[2] ;
 wire \stop.syn.filt.m1.b_latched[3] ;
 wire \stop.syn.filt.m1.b_latched[4] ;
 wire \stop.syn.filt.m1.b_latched[5] ;
 wire \stop.syn.filt.m1.b_latched[6] ;
 wire \stop.syn.filt.m1.b_latched[7] ;
 wire \stop.syn.filt.m1.sum[10] ;
 wire \stop.syn.filt.m1.sum[11] ;
 wire \stop.syn.filt.m1.sum[12] ;
 wire \stop.syn.filt.m1.sum[13] ;
 wire \stop.syn.filt.m1.sum[14] ;
 wire \stop.syn.filt.m1.sum[15] ;
 wire \stop.syn.filt.m1.sum[16] ;
 wire \stop.syn.filt.m1.sum[1] ;
 wire \stop.syn.filt.m1.sum[2] ;
 wire \stop.syn.filt.m1.sum[3] ;
 wire \stop.syn.filt.m1.sum[4] ;
 wire \stop.syn.filt.m1.sum[5] ;
 wire \stop.syn.filt.m1.sum[6] ;
 wire \stop.syn.filt.m1.sum[7] ;
 wire \stop.syn.filt.m1.sum[8] ;
 wire \stop.syn.filt.m1.sum[9] ;
 wire \stop.syn.filt.m1.sum_in2[0] ;
 wire \stop.syn.filt.m1.sum_in2[10] ;
 wire \stop.syn.filt.m1.sum_in2[11] ;
 wire \stop.syn.filt.m1.sum_in2[12] ;
 wire \stop.syn.filt.m1.sum_in2[13] ;
 wire \stop.syn.filt.m1.sum_in2[14] ;
 wire \stop.syn.filt.m1.sum_in2[15] ;
 wire \stop.syn.filt.m1.sum_in2[1] ;
 wire \stop.syn.filt.m1.sum_in2[2] ;
 wire \stop.syn.filt.m1.sum_in2[3] ;
 wire \stop.syn.filt.m1.sum_in2[4] ;
 wire \stop.syn.filt.m1.sum_in2[5] ;
 wire \stop.syn.filt.m1.sum_in2[6] ;
 wire \stop.syn.filt.m1.sum_in2[7] ;
 wire \stop.syn.filt.m1.sum_in2[8] ;
 wire \stop.syn.filt.m1.sum_in2[9] ;
 wire \stop.syn.filt.m2.b_bit ;
 wire \stop.syn.filt.m2.b_latched[1] ;
 wire \stop.syn.filt.m2.b_latched[2] ;
 wire \stop.syn.filt.m2.b_latched[3] ;
 wire \stop.syn.filt.m2.b_latched[4] ;
 wire \stop.syn.filt.m2.b_latched[5] ;
 wire \stop.syn.filt.m2.b_latched[6] ;
 wire \stop.syn.filt.m2.b_latched[7] ;
 wire \stop.syn.filt.m2.sum[10] ;
 wire \stop.syn.filt.m2.sum[11] ;
 wire \stop.syn.filt.m2.sum[12] ;
 wire \stop.syn.filt.m2.sum[13] ;
 wire \stop.syn.filt.m2.sum[14] ;
 wire \stop.syn.filt.m2.sum[15] ;
 wire \stop.syn.filt.m2.sum[16] ;
 wire \stop.syn.filt.m2.sum[1] ;
 wire \stop.syn.filt.m2.sum[2] ;
 wire \stop.syn.filt.m2.sum[3] ;
 wire \stop.syn.filt.m2.sum[4] ;
 wire \stop.syn.filt.m2.sum[5] ;
 wire \stop.syn.filt.m2.sum[6] ;
 wire \stop.syn.filt.m2.sum[7] ;
 wire \stop.syn.filt.m2.sum[8] ;
 wire \stop.syn.filt.m2.sum[9] ;
 wire \stop.syn.filt.m2.sum_in2[0] ;
 wire \stop.syn.filt.m2.sum_in2[10] ;
 wire \stop.syn.filt.m2.sum_in2[11] ;
 wire \stop.syn.filt.m2.sum_in2[12] ;
 wire \stop.syn.filt.m2.sum_in2[13] ;
 wire \stop.syn.filt.m2.sum_in2[14] ;
 wire \stop.syn.filt.m2.sum_in2[15] ;
 wire \stop.syn.filt.m2.sum_in2[1] ;
 wire \stop.syn.filt.m2.sum_in2[2] ;
 wire \stop.syn.filt.m2.sum_in2[3] ;
 wire \stop.syn.filt.m2.sum_in2[4] ;
 wire \stop.syn.filt.m2.sum_in2[5] ;
 wire \stop.syn.filt.m2.sum_in2[6] ;
 wire \stop.syn.filt.m2.sum_in2[7] ;
 wire \stop.syn.filt.m2.sum_in2[8] ;
 wire \stop.syn.filt.m2.sum_in2[9] ;
 wire \stop.syn.osci.counter[0] ;
 wire \stop.syn.osci.counter[10] ;
 wire \stop.syn.osci.counter[11] ;
 wire \stop.syn.osci.counter[1] ;
 wire \stop.syn.osci.counter[2] ;
 wire \stop.syn.osci.counter[3] ;
 wire \stop.syn.osci.counter[4] ;
 wire \stop.syn.osci.counter[5] ;
 wire \stop.syn.osci.counter[6] ;
 wire \stop.syn.osci.counter[7] ;
 wire \stop.syn.osci.counter[8] ;
 wire \stop.syn.osci.counter[9] ;
 wire \stop.syn.osci.data_buf ;
 wire \stop.syn.rstn_fst_reg1 ;
 wire \stop.syn.rstn_fst_reg2 ;
 wire \stop.syn.rstn_reg1 ;
 wire \stop.syn.smul8.b_bit ;
 wire \stop.syn.smul8.b_latched[1] ;
 wire \stop.syn.smul8.b_latched[2] ;
 wire \stop.syn.smul8.b_latched[3] ;
 wire \stop.syn.smul8.b_latched[4] ;
 wire \stop.syn.smul8.b_latched[5] ;
 wire \stop.syn.smul8.b_latched[6] ;
 wire \stop.syn.smul8.b_latched[7] ;
 wire \stop.syn.trig_reg1 ;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;

 sg13g2_inv_1 _0986_ (.Y(_0299_),
    .A(\stop.syn.adsri.envelope[1] ));
 sg13g2_inv_1 _0987_ (.Y(_0300_),
    .A(\stop.syn.adsri.envelope[0] ));
 sg13g2_inv_1 _0988_ (.Y(_0082_),
    .A(\stop.ctrl.first_bit ));
 sg13g2_inv_1 _0989_ (.Y(_0301_),
    .A(\stop.syn.adsri.state[0] ));
 sg13g2_inv_1 _0990_ (.Y(_0302_),
    .A(\stop.syn.adsri.trig ));
 sg13g2_inv_2 _0991_ (.Y(_0303_),
    .A(\stop.syn.adsri.state[3] ));
 sg13g2_inv_1 _0992_ (.Y(_0304_),
    .A(\stop.adsr_ai[2] ));
 sg13g2_inv_1 _0993_ (.Y(_0305_),
    .A(\stop.adsr_ai[3] ));
 sg13g2_inv_1 _0994_ (.Y(_0306_),
    .A(\stop.adsr_ai[4] ));
 sg13g2_inv_1 _0995_ (.Y(_0307_),
    .A(\stop.adsr_ai[5] ));
 sg13g2_inv_1 _0996_ (.Y(_0308_),
    .A(\stop.adsr_ai[6] ));
 sg13g2_inv_1 _0997_ (.Y(_0309_),
    .A(\stop.adsr_ai[7] ));
 sg13g2_inv_1 _0998_ (.Y(_0083_),
    .A(net2));
 sg13g2_inv_1 _0999_ (.Y(_0310_),
    .A(\stop.syn.filt.m1.sum_in2[6] ));
 sg13g2_inv_1 _1000_ (.Y(_0311_),
    .A(_0052_));
 sg13g2_inv_1 _1001_ (.Y(_0312_),
    .A(_0053_));
 sg13g2_nor2b_1 _1002_ (.A(\stop.syn.clk_sample_x2 ),
    .B_N(net298),
    .Y(_0313_));
 sg13g2_inv_4 _1003_ (.A(net296),
    .Y(_0133_));
 sg13g2_and2_1 _1004_ (.A(\stop.ctrl.cfg[51] ),
    .B(net288),
    .X(_0158_));
 sg13g2_and2_1 _1005_ (.A(\stop.ctrl.cfg[59] ),
    .B(net295),
    .X(_0156_));
 sg13g2_and2_1 _1006_ (.A(\stop.syn.adsri.envelope[7] ),
    .B(net294),
    .X(_0134_));
 sg13g2_a22oi_1 _1007_ (.Y(_0314_),
    .B1(\stop.adsr_di[6] ),
    .B2(net282),
    .A2(\stop.adsr_ri[6] ),
    .A1(net283));
 sg13g2_o21ai_1 _1008_ (.B1(_0314_),
    .Y(_0315_),
    .A1(_0303_),
    .A2(_0308_));
 sg13g2_and2_1 _1009_ (.A(\stop.syn.adsri.envelope[6] ),
    .B(_0315_),
    .X(_0316_));
 sg13g2_xor2_1 _1010_ (.B(_0315_),
    .A(\stop.syn.adsri.envelope[6] ),
    .X(_0317_));
 sg13g2_a22oi_1 _1011_ (.Y(_0318_),
    .B1(\stop.adsr_di[5] ),
    .B2(net282),
    .A2(\stop.adsr_ri[5] ),
    .A1(net283));
 sg13g2_o21ai_1 _1012_ (.B1(_0318_),
    .Y(_0319_),
    .A1(_0303_),
    .A2(_0307_));
 sg13g2_and2_1 _1013_ (.A(\stop.syn.adsri.envelope[5] ),
    .B(_0319_),
    .X(_0320_));
 sg13g2_a22oi_1 _1014_ (.Y(_0321_),
    .B1(\stop.adsr_di[4] ),
    .B2(net282),
    .A2(\stop.adsr_ri[4] ),
    .A1(net283));
 sg13g2_o21ai_1 _1015_ (.B1(_0321_),
    .Y(_0322_),
    .A1(_0303_),
    .A2(_0306_));
 sg13g2_and2_1 _1016_ (.A(\stop.syn.adsri.envelope[4] ),
    .B(_0322_),
    .X(_0323_));
 sg13g2_a22oi_1 _1017_ (.Y(_0324_),
    .B1(\stop.adsr_di[3] ),
    .B2(\stop.syn.adsri.state[2] ),
    .A2(\stop.adsr_ri[3] ),
    .A1(net284));
 sg13g2_o21ai_1 _1018_ (.B1(_0324_),
    .Y(_0325_),
    .A1(_0303_),
    .A2(_0305_));
 sg13g2_nand2_1 _1019_ (.Y(_0326_),
    .A(\stop.syn.adsri.envelope[3] ),
    .B(_0325_));
 sg13g2_nor2_1 _1020_ (.A(\stop.syn.adsri.envelope[3] ),
    .B(_0325_),
    .Y(_0327_));
 sg13g2_a22oi_1 _1021_ (.Y(_0328_),
    .B1(\stop.adsr_di[2] ),
    .B2(\stop.syn.adsri.state[2] ),
    .A2(\stop.adsr_ri[2] ),
    .A1(net284));
 sg13g2_o21ai_1 _1022_ (.B1(_0328_),
    .Y(_0329_),
    .A1(_0303_),
    .A2(_0304_));
 sg13g2_and2_1 _1023_ (.A(\stop.syn.adsri.envelope[2] ),
    .B(_0329_),
    .X(_0330_));
 sg13g2_nand2_1 _1024_ (.Y(_0331_),
    .A(\stop.syn.adsri.state[3] ),
    .B(\stop.adsr_ai[1] ));
 sg13g2_a22oi_1 _1025_ (.Y(_0332_),
    .B1(\stop.adsr_di[1] ),
    .B2(\stop.syn.adsri.state[2] ),
    .A2(\stop.adsr_ri[1] ),
    .A1(net284));
 sg13g2_a21oi_1 _1026_ (.A1(_0331_),
    .A2(_0332_),
    .Y(_0333_),
    .B1(_0299_));
 sg13g2_a21o_1 _1027_ (.A2(_0332_),
    .A1(_0331_),
    .B1(_0299_),
    .X(_0334_));
 sg13g2_nand2_1 _1028_ (.Y(_0335_),
    .A(\stop.adsr_ri[0] ),
    .B(net284));
 sg13g2_a22oi_1 _1029_ (.Y(_0336_),
    .B1(\stop.adsr_ai[0] ),
    .B2(\stop.syn.adsri.state[3] ),
    .A2(\stop.adsr_di[0] ),
    .A1(net282));
 sg13g2_a21o_1 _1030_ (.A2(_0336_),
    .A1(_0335_),
    .B1(_0300_),
    .X(_0337_));
 sg13g2_and3_1 _1031_ (.X(_0338_),
    .A(_0299_),
    .B(_0331_),
    .C(_0332_));
 sg13g2_nor2_1 _1032_ (.A(_0333_),
    .B(_0338_),
    .Y(_0339_));
 sg13g2_o21ai_1 _1033_ (.B1(_0334_),
    .Y(_0340_),
    .A1(_0337_),
    .A2(_0338_));
 sg13g2_xor2_1 _1034_ (.B(_0329_),
    .A(\stop.syn.adsri.envelope[2] ),
    .X(_0341_));
 sg13g2_a21oi_2 _1035_ (.B1(_0330_),
    .Y(_0342_),
    .A2(_0341_),
    .A1(_0340_));
 sg13g2_a21oi_2 _1036_ (.B1(_0327_),
    .Y(_0343_),
    .A2(_0342_),
    .A1(_0326_));
 sg13g2_xor2_1 _1037_ (.B(_0322_),
    .A(\stop.syn.adsri.envelope[4] ),
    .X(_0344_));
 sg13g2_a21oi_1 _1038_ (.A1(_0343_),
    .A2(_0344_),
    .Y(_0345_),
    .B1(_0323_));
 sg13g2_xor2_1 _1039_ (.B(_0319_),
    .A(\stop.syn.adsri.envelope[5] ),
    .X(_0346_));
 sg13g2_and2_1 _1040_ (.A(_0344_),
    .B(_0346_),
    .X(_0347_));
 sg13g2_a21o_1 _1041_ (.A2(_0346_),
    .A1(_0323_),
    .B1(_0320_),
    .X(_0348_));
 sg13g2_a21o_1 _1042_ (.A2(_0347_),
    .A1(_0343_),
    .B1(_0348_),
    .X(_0349_));
 sg13g2_a21oi_1 _1043_ (.A1(_0317_),
    .A2(_0349_),
    .Y(_0350_),
    .B1(_0316_));
 sg13g2_a22oi_1 _1044_ (.Y(_0351_),
    .B1(\stop.adsr_di[7] ),
    .B2(net282),
    .A2(\stop.adsr_ri[7] ),
    .A1(net283));
 sg13g2_o21ai_1 _1045_ (.B1(_0351_),
    .Y(_0352_),
    .A1(_0303_),
    .A2(_0309_));
 sg13g2_xor2_1 _1046_ (.B(_0352_),
    .A(\stop.syn.adsri.envelope[7] ),
    .X(_0353_));
 sg13g2_nor2b_1 _1047_ (.A(_0350_),
    .B_N(_0353_),
    .Y(_0354_));
 sg13g2_xnor2_1 _1048_ (.Y(_0355_),
    .A(_0350_),
    .B(_0353_));
 sg13g2_inv_1 _1049_ (.Y(_0356_),
    .A(_0355_));
 sg13g2_xnor2_1 _1050_ (.Y(_0357_),
    .A(\stop.adsr_s[7] ),
    .B(_0355_));
 sg13g2_xnor2_1 _1051_ (.Y(_0358_),
    .A(_0317_),
    .B(_0349_));
 sg13g2_xor2_1 _1052_ (.B(_0346_),
    .A(_0345_),
    .X(_0359_));
 sg13g2_xnor2_1 _1053_ (.Y(_0360_),
    .A(_0343_),
    .B(_0344_));
 sg13g2_xnor2_1 _1054_ (.Y(_0361_),
    .A(\stop.syn.adsri.envelope[3] ),
    .B(_0325_));
 sg13g2_xnor2_1 _1055_ (.Y(_0362_),
    .A(_0342_),
    .B(_0361_));
 sg13g2_xnor2_1 _1056_ (.Y(_0363_),
    .A(_0340_),
    .B(_0341_));
 sg13g2_xor2_1 _1057_ (.B(_0339_),
    .A(_0337_),
    .X(_0364_));
 sg13g2_nand3_1 _1058_ (.B(_0335_),
    .C(_0336_),
    .A(_0300_),
    .Y(_0365_));
 sg13g2_nand2_2 _1059_ (.Y(_0366_),
    .A(_0337_),
    .B(_0365_));
 sg13g2_xnor2_1 _1060_ (.Y(_0367_),
    .A(\stop.adsr_s[0] ),
    .B(_0366_));
 sg13g2_xnor2_1 _1061_ (.Y(_0368_),
    .A(\stop.adsr_s[1] ),
    .B(_0364_));
 sg13g2_xnor2_1 _1062_ (.Y(_0369_),
    .A(\stop.adsr_s[2] ),
    .B(_0363_));
 sg13g2_xnor2_1 _1063_ (.Y(_0370_),
    .A(\stop.adsr_s[3] ),
    .B(_0362_));
 sg13g2_nor4_1 _1064_ (.A(_0367_),
    .B(_0368_),
    .C(_0369_),
    .D(_0370_),
    .Y(_0371_));
 sg13g2_xor2_1 _1065_ (.B(_0360_),
    .A(\stop.adsr_s[4] ),
    .X(_0372_));
 sg13g2_xor2_1 _1066_ (.B(_0359_),
    .A(\stop.adsr_s[5] ),
    .X(_0373_));
 sg13g2_xor2_1 _1067_ (.B(_0358_),
    .A(\stop.adsr_s[6] ),
    .X(_0374_));
 sg13g2_nand4_1 _1068_ (.B(_0372_),
    .C(_0373_),
    .A(_0371_),
    .Y(_0375_),
    .D(_0374_));
 sg13g2_nand2b_1 _1069_ (.Y(_0376_),
    .B(_0357_),
    .A_N(_0375_));
 sg13g2_nor2b_1 _1070_ (.A(\stop.syn.adsri.state[4] ),
    .B_N(_0376_),
    .Y(_0377_));
 sg13g2_nand2_1 _1071_ (.Y(_0378_),
    .A(net281),
    .B(\stop.syn.adsri.trig ));
 sg13g2_nor2_1 _1072_ (.A(net282),
    .B(\stop.syn.adsri.state[4] ),
    .Y(_0379_));
 sg13g2_nor3_1 _1073_ (.A(_0377_),
    .B(_0378_),
    .C(_0379_),
    .Y(_0004_));
 sg13g2_a21oi_2 _1074_ (.B1(_0354_),
    .Y(_0380_),
    .A2(_0352_),
    .A1(\stop.syn.adsri.envelope[7] ));
 sg13g2_nor2_1 _1075_ (.A(net282),
    .B(net283),
    .Y(_0381_));
 sg13g2_xor2_1 _1076_ (.B(_0381_),
    .A(_0380_),
    .X(_0382_));
 sg13g2_o21ai_1 _1077_ (.B1(_0301_),
    .Y(_0383_),
    .A1(_0303_),
    .A2(_0382_));
 sg13g2_nor2b_1 _1078_ (.A(_0378_),
    .B_N(_0383_),
    .Y(_0003_));
 sg13g2_a22oi_1 _1079_ (.Y(_0384_),
    .B1(_0382_),
    .B2(\stop.syn.adsri.state[3] ),
    .A2(_0376_),
    .A1(net282));
 sg13g2_nor2_1 _1080_ (.A(_0378_),
    .B(_0384_),
    .Y(_0002_));
 sg13g2_nor2b_1 _1081_ (.A(\stop.syn.adsri.trig ),
    .B_N(net281),
    .Y(_0385_));
 sg13g2_nand2_1 _1082_ (.Y(_0386_),
    .A(_0303_),
    .B(_0379_));
 sg13g2_nand2_1 _1083_ (.Y(_0387_),
    .A(_0385_),
    .B(_0386_));
 sg13g2_nand2_1 _1084_ (.Y(_0388_),
    .A(net281),
    .B(net283));
 sg13g2_o21ai_1 _1085_ (.B1(_0387_),
    .Y(_0001_),
    .A1(_0380_),
    .A2(_0388_));
 sg13g2_nand2_1 _1086_ (.Y(_0389_),
    .A(net283),
    .B(_0380_));
 sg13g2_a21oi_1 _1087_ (.A1(\stop.syn.adsri.state[0] ),
    .A2(_0385_),
    .Y(_0390_),
    .B1(_0047_));
 sg13g2_nand2_1 _1088_ (.Y(_0000_),
    .A(_0389_),
    .B(_0390_));
 sg13g2_nor2_1 _1089_ (.A(\stop.syn.smul8.b_latched[1] ),
    .B(net292),
    .Y(_0391_));
 sg13g2_a21oi_2 _1090_ (.B1(_0391_),
    .Y(_0019_),
    .A2(net292),
    .A1(_0300_));
 sg13g2_nand2_1 _1091_ (.Y(_0392_),
    .A(\stop.syn.smul8.b_latched[2] ),
    .B(_0133_));
 sg13g2_o21ai_1 _1092_ (.B1(_0392_),
    .Y(_0020_),
    .A1(_0299_),
    .A2(_0133_));
 sg13g2_mux2_1 _1093_ (.A0(\stop.syn.adsri.envelope[2] ),
    .A1(\stop.syn.smul8.b_latched[3] ),
    .S(_0133_),
    .X(_0021_));
 sg13g2_mux2_1 _1094_ (.A0(\stop.syn.adsri.envelope[3] ),
    .A1(\stop.syn.smul8.b_latched[4] ),
    .S(_0133_),
    .X(_0022_));
 sg13g2_mux2_1 _1095_ (.A0(\stop.syn.adsri.envelope[4] ),
    .A1(\stop.syn.smul8.b_latched[5] ),
    .S(_0133_),
    .X(_0023_));
 sg13g2_mux2_1 _1096_ (.A0(\stop.syn.adsri.envelope[5] ),
    .A1(\stop.syn.smul8.b_latched[6] ),
    .S(_0133_),
    .X(_0024_));
 sg13g2_mux2_1 _1097_ (.A0(\stop.syn.adsri.envelope[6] ),
    .A1(\stop.syn.smul8.b_latched[7] ),
    .S(_0133_),
    .X(_0025_));
 sg13g2_mux2_1 _1098_ (.A0(\stop.syn.filt.m2.b_latched[1] ),
    .A1(\stop.ctrl.cfg[52] ),
    .S(net295),
    .X(_0012_));
 sg13g2_mux2_1 _1099_ (.A0(\stop.syn.filt.m2.b_latched[2] ),
    .A1(\stop.ctrl.cfg[53] ),
    .S(net295),
    .X(_0013_));
 sg13g2_mux2_1 _1100_ (.A0(\stop.syn.filt.m2.b_latched[3] ),
    .A1(\stop.ctrl.cfg[54] ),
    .S(net295),
    .X(_0014_));
 sg13g2_mux2_1 _1101_ (.A0(\stop.syn.filt.m2.b_latched[4] ),
    .A1(\stop.ctrl.cfg[55] ),
    .S(net295),
    .X(_0015_));
 sg13g2_mux2_1 _1102_ (.A0(\stop.syn.filt.m2.b_latched[5] ),
    .A1(\stop.ctrl.cfg[56] ),
    .S(net295),
    .X(_0016_));
 sg13g2_mux2_1 _1103_ (.A0(\stop.syn.filt.m2.b_latched[6] ),
    .A1(\stop.ctrl.cfg[57] ),
    .S(net295),
    .X(_0017_));
 sg13g2_mux2_1 _1104_ (.A0(\stop.syn.filt.m2.b_latched[7] ),
    .A1(\stop.ctrl.cfg[58] ),
    .S(net295),
    .X(_0018_));
 sg13g2_mux2_1 _1105_ (.A0(\stop.syn.filt.m1.b_latched[1] ),
    .A1(\stop.ctrl.cfg[44] ),
    .S(net287),
    .X(_0005_));
 sg13g2_mux2_1 _1106_ (.A0(\stop.syn.filt.m1.b_latched[2] ),
    .A1(\stop.ctrl.cfg[45] ),
    .S(net287),
    .X(_0006_));
 sg13g2_mux2_1 _1107_ (.A0(\stop.syn.filt.m1.b_latched[3] ),
    .A1(\stop.ctrl.cfg[46] ),
    .S(net287),
    .X(_0007_));
 sg13g2_mux2_1 _1108_ (.A0(\stop.syn.filt.m1.b_latched[4] ),
    .A1(\stop.ctrl.cfg[47] ),
    .S(net287),
    .X(_0008_));
 sg13g2_mux2_1 _1109_ (.A0(\stop.syn.filt.m1.b_latched[5] ),
    .A1(\stop.ctrl.cfg[48] ),
    .S(net287),
    .X(_0009_));
 sg13g2_mux2_1 _1110_ (.A0(\stop.syn.filt.m1.b_latched[6] ),
    .A1(\stop.ctrl.cfg[49] ),
    .S(net288),
    .X(_0010_));
 sg13g2_mux2_1 _1111_ (.A0(\stop.syn.filt.m1.b_latched[7] ),
    .A1(\stop.ctrl.cfg[50] ),
    .S(net287),
    .X(_0011_));
 sg13g2_nand3_1 _1112_ (.B(\stop.syn.daci.din[0] ),
    .C(\stop.syn.filt.m1.sum_in2[0] ),
    .A(net313),
    .Y(_0393_));
 sg13g2_and3_1 _1113_ (.X(_0394_),
    .A(net313),
    .B(\stop.syn.daci.din[1] ),
    .C(\stop.syn.filt.m1.sum_in2[1] ));
 sg13g2_nand3_1 _1114_ (.B(\stop.syn.daci.din[1] ),
    .C(\stop.syn.filt.m1.sum_in2[1] ),
    .A(net313),
    .Y(_0395_));
 sg13g2_a21oi_1 _1115_ (.A1(net312),
    .A2(\stop.syn.daci.din[1] ),
    .Y(_0396_),
    .B1(\stop.syn.filt.m1.sum_in2[1] ));
 sg13g2_nor2_1 _1116_ (.A(_0394_),
    .B(_0396_),
    .Y(_0397_));
 sg13g2_xnor2_1 _1117_ (.Y(\stop.syn.filt.m1.sum[1] ),
    .A(_0393_),
    .B(_0397_));
 sg13g2_o21ai_1 _1118_ (.B1(_0395_),
    .Y(_0398_),
    .A1(_0393_),
    .A2(_0396_));
 sg13g2_and3_1 _1119_ (.X(_0399_),
    .A(net312),
    .B(\stop.syn.daci.din[2] ),
    .C(\stop.syn.filt.m1.sum_in2[2] ));
 sg13g2_a21o_1 _1120_ (.A2(\stop.syn.daci.din[2] ),
    .A1(net312),
    .B1(\stop.syn.filt.m1.sum_in2[2] ),
    .X(_0400_));
 sg13g2_nand2b_1 _1121_ (.Y(_0401_),
    .B(_0400_),
    .A_N(_0399_));
 sg13g2_xnor2_1 _1122_ (.Y(\stop.syn.filt.m1.sum[2] ),
    .A(_0398_),
    .B(_0401_));
 sg13g2_a21o_1 _1123_ (.A2(_0400_),
    .A1(_0398_),
    .B1(_0399_),
    .X(_0402_));
 sg13g2_nand2_1 _1124_ (.Y(_0403_),
    .A(net312),
    .B(\stop.syn.daci.din[3] ));
 sg13g2_nor2_1 _1125_ (.A(_0048_),
    .B(_0403_),
    .Y(_0404_));
 sg13g2_xor2_1 _1126_ (.B(_0403_),
    .A(_0048_),
    .X(_0405_));
 sg13g2_xor2_1 _1127_ (.B(_0405_),
    .A(_0402_),
    .X(\stop.syn.filt.m1.sum[3] ));
 sg13g2_a21oi_2 _1128_ (.B1(_0404_),
    .Y(_0406_),
    .A2(_0405_),
    .A1(_0402_));
 sg13g2_nand3_1 _1129_ (.B(\stop.syn.daci.din[4] ),
    .C(\stop.syn.filt.m1.sum_in2[4] ),
    .A(net312),
    .Y(_0407_));
 sg13g2_a21o_1 _1130_ (.A2(\stop.syn.daci.din[4] ),
    .A1(net312),
    .B1(\stop.syn.filt.m1.sum_in2[4] ),
    .X(_0408_));
 sg13g2_nand2_1 _1131_ (.Y(_0409_),
    .A(_0407_),
    .B(_0408_));
 sg13g2_xor2_1 _1132_ (.B(_0409_),
    .A(_0406_),
    .X(\stop.syn.filt.m1.sum[4] ));
 sg13g2_nand2_1 _1133_ (.Y(_0410_),
    .A(net312),
    .B(\stop.syn.daci.din[5] ));
 sg13g2_nor2_1 _1134_ (.A(_0049_),
    .B(_0410_),
    .Y(_0411_));
 sg13g2_xor2_1 _1135_ (.B(_0410_),
    .A(_0049_),
    .X(_0412_));
 sg13g2_o21ai_1 _1136_ (.B1(_0407_),
    .Y(_0413_),
    .A1(_0406_),
    .A2(_0409_));
 sg13g2_xor2_1 _1137_ (.B(_0413_),
    .A(_0412_),
    .X(\stop.syn.filt.m1.sum[5] ));
 sg13g2_nand2b_1 _1138_ (.Y(_0414_),
    .B(_0412_),
    .A_N(_0409_));
 sg13g2_a21oi_1 _1139_ (.A1(_0049_),
    .A2(_0410_),
    .Y(_0415_),
    .B1(_0407_));
 sg13g2_nor2_1 _1140_ (.A(_0411_),
    .B(_0415_),
    .Y(_0416_));
 sg13g2_o21ai_1 _1141_ (.B1(_0416_),
    .Y(_0417_),
    .A1(_0406_),
    .A2(_0414_));
 sg13g2_nand2_1 _1142_ (.Y(_0418_),
    .A(net312),
    .B(\stop.syn.daci.din[6] ));
 sg13g2_xnor2_1 _1143_ (.Y(_0419_),
    .A(_0310_),
    .B(_0418_));
 sg13g2_nand2b_1 _1144_ (.Y(_0420_),
    .B(_0417_),
    .A_N(_0419_));
 sg13g2_xnor2_1 _1145_ (.Y(\stop.syn.filt.m1.sum[6] ),
    .A(_0417_),
    .B(_0419_));
 sg13g2_o21ai_1 _1146_ (.B1(_0420_),
    .Y(_0421_),
    .A1(_0310_),
    .A2(_0418_));
 sg13g2_and3_1 _1147_ (.X(_0422_),
    .A(net311),
    .B(\stop.syn.daci.din[7] ),
    .C(\stop.syn.filt.m1.sum_in2[7] ));
 sg13g2_a21o_1 _1148_ (.A2(\stop.syn.daci.din[7] ),
    .A1(net311),
    .B1(\stop.syn.filt.m1.sum_in2[7] ),
    .X(_0423_));
 sg13g2_nand2b_1 _1149_ (.Y(_0424_),
    .B(_0423_),
    .A_N(_0422_));
 sg13g2_xnor2_1 _1150_ (.Y(\stop.syn.filt.m1.sum[7] ),
    .A(_0421_),
    .B(_0424_));
 sg13g2_a21o_2 _1151_ (.A2(_0423_),
    .A1(_0421_),
    .B1(_0422_),
    .X(_0425_));
 sg13g2_inv_1 _1152_ (.Y(_0426_),
    .A(_0425_));
 sg13g2_nand3_1 _1153_ (.B(\stop.syn.daci.din[8] ),
    .C(\stop.syn.filt.m1.sum_in2[8] ),
    .A(net311),
    .Y(_0427_));
 sg13g2_a21o_1 _1154_ (.A2(\stop.syn.daci.din[8] ),
    .A1(net311),
    .B1(\stop.syn.filt.m1.sum_in2[8] ),
    .X(_0428_));
 sg13g2_nand2_1 _1155_ (.Y(_0429_),
    .A(_0427_),
    .B(_0428_));
 sg13g2_xnor2_1 _1156_ (.Y(\stop.syn.filt.m1.sum[8] ),
    .A(_0425_),
    .B(_0429_));
 sg13g2_nand2_1 _1157_ (.Y(_0430_),
    .A(net309),
    .B(\stop.syn.daci.din[9] ));
 sg13g2_nand2_1 _1158_ (.Y(_0431_),
    .A(_0050_),
    .B(_0430_));
 sg13g2_xor2_1 _1159_ (.B(_0430_),
    .A(_0050_),
    .X(_0432_));
 sg13g2_o21ai_1 _1160_ (.B1(_0427_),
    .Y(_0433_),
    .A1(_0426_),
    .A2(_0429_));
 sg13g2_xor2_1 _1161_ (.B(_0433_),
    .A(_0432_),
    .X(\stop.syn.filt.m1.sum[9] ));
 sg13g2_nand3_1 _1162_ (.B(\stop.syn.daci.din[10] ),
    .C(\stop.syn.filt.m1.sum_in2[10] ),
    .A(net309),
    .Y(_0434_));
 sg13g2_a21o_1 _1163_ (.A2(\stop.syn.daci.din[10] ),
    .A1(net309),
    .B1(\stop.syn.filt.m1.sum_in2[10] ),
    .X(_0435_));
 sg13g2_nand2_1 _1164_ (.Y(_0436_),
    .A(_0434_),
    .B(_0435_));
 sg13g2_nand2b_1 _1165_ (.Y(_0437_),
    .B(_0432_),
    .A_N(_0429_));
 sg13g2_nand2b_1 _1166_ (.Y(_0438_),
    .B(_0425_),
    .A_N(_0437_));
 sg13g2_o21ai_1 _1167_ (.B1(_0427_),
    .Y(_0439_),
    .A1(_0050_),
    .A2(_0430_));
 sg13g2_nand2_1 _1168_ (.Y(_0440_),
    .A(_0431_),
    .B(_0439_));
 sg13g2_and2_1 _1169_ (.A(_0438_),
    .B(_0440_),
    .X(_0441_));
 sg13g2_xor2_1 _1170_ (.B(_0441_),
    .A(_0436_),
    .X(\stop.syn.filt.m1.sum[10] ));
 sg13g2_a21o_1 _1171_ (.A2(\stop.syn.daci.din[11] ),
    .A1(net309),
    .B1(\stop.syn.filt.m1.sum_in2[11] ),
    .X(_0442_));
 sg13g2_nand3_1 _1172_ (.B(\stop.syn.daci.din[11] ),
    .C(\stop.syn.filt.m1.sum_in2[11] ),
    .A(net309),
    .Y(_0443_));
 sg13g2_nand2_1 _1173_ (.Y(_0444_),
    .A(_0442_),
    .B(_0443_));
 sg13g2_o21ai_1 _1174_ (.B1(_0434_),
    .Y(_0445_),
    .A1(_0436_),
    .A2(_0441_));
 sg13g2_xnor2_1 _1175_ (.Y(\stop.syn.filt.m1.sum[11] ),
    .A(_0444_),
    .B(_0445_));
 sg13g2_nand3_1 _1176_ (.B(\stop.syn.daci.din[12] ),
    .C(\stop.syn.filt.m1.sum_in2[12] ),
    .A(net310),
    .Y(_0446_));
 sg13g2_a21o_1 _1177_ (.A2(\stop.syn.daci.din[12] ),
    .A1(net310),
    .B1(\stop.syn.filt.m1.sum_in2[12] ),
    .X(_0447_));
 sg13g2_nand2_1 _1178_ (.Y(_0448_),
    .A(_0446_),
    .B(_0447_));
 sg13g2_nand2_1 _1179_ (.Y(_0449_),
    .A(_0434_),
    .B(_0443_));
 sg13g2_or2_1 _1180_ (.X(_0450_),
    .B(_0444_),
    .A(_0436_));
 sg13g2_nor2_1 _1181_ (.A(_0440_),
    .B(_0450_),
    .Y(_0451_));
 sg13g2_nor2_1 _1182_ (.A(_0437_),
    .B(_0450_),
    .Y(_0452_));
 sg13g2_a221oi_1 _1183_ (.B2(_0425_),
    .C1(_0451_),
    .B1(_0452_),
    .A1(_0442_),
    .Y(_0453_),
    .A2(_0449_));
 sg13g2_xor2_1 _1184_ (.B(_0453_),
    .A(_0448_),
    .X(\stop.syn.filt.m1.sum[12] ));
 sg13g2_o21ai_1 _1185_ (.B1(_0446_),
    .Y(_0454_),
    .A1(_0448_),
    .A2(_0453_));
 sg13g2_nand2_1 _1186_ (.Y(_0455_),
    .A(net310),
    .B(\stop.syn.daci.din[13] ));
 sg13g2_nor2_1 _1187_ (.A(_0051_),
    .B(_0455_),
    .Y(_0456_));
 sg13g2_xor2_1 _1188_ (.B(_0455_),
    .A(_0051_),
    .X(_0457_));
 sg13g2_xor2_1 _1189_ (.B(_0457_),
    .A(_0454_),
    .X(\stop.syn.filt.m1.sum[13] ));
 sg13g2_nand2b_1 _1190_ (.Y(_0458_),
    .B(_0457_),
    .A_N(_0448_));
 sg13g2_a21oi_1 _1191_ (.A1(_0051_),
    .A2(_0455_),
    .Y(_0459_),
    .B1(_0446_));
 sg13g2_nor2_1 _1192_ (.A(_0456_),
    .B(_0459_),
    .Y(_0460_));
 sg13g2_o21ai_1 _1193_ (.B1(_0460_),
    .Y(_0461_),
    .A1(_0453_),
    .A2(_0458_));
 sg13g2_and3_1 _1194_ (.X(_0462_),
    .A(net310),
    .B(\stop.syn.daci.din[14] ),
    .C(\stop.syn.filt.m1.sum_in2[14] ));
 sg13g2_a21o_1 _1195_ (.A2(\stop.syn.daci.din[14] ),
    .A1(net310),
    .B1(\stop.syn.filt.m1.sum_in2[14] ),
    .X(_0463_));
 sg13g2_nand2b_1 _1196_ (.Y(_0464_),
    .B(_0463_),
    .A_N(_0462_));
 sg13g2_xnor2_1 _1197_ (.Y(\stop.syn.filt.m1.sum[14] ),
    .A(_0461_),
    .B(_0464_));
 sg13g2_and3_1 _1198_ (.X(_0465_),
    .A(net309),
    .B(\stop.syn.daci.din[15] ),
    .C(\stop.syn.filt.m1.sum_in2[15] ));
 sg13g2_nand3_1 _1199_ (.B(\stop.syn.daci.din[15] ),
    .C(\stop.syn.filt.m1.sum_in2[15] ),
    .A(net309),
    .Y(_0466_));
 sg13g2_a21oi_1 _1200_ (.A1(net309),
    .A2(\stop.syn.daci.din[15] ),
    .Y(_0467_),
    .B1(\stop.syn.filt.m1.sum_in2[15] ));
 sg13g2_nor2_1 _1201_ (.A(_0465_),
    .B(_0467_),
    .Y(_0468_));
 sg13g2_a21oi_1 _1202_ (.A1(_0461_),
    .A2(_0463_),
    .Y(_0469_),
    .B1(_0462_));
 sg13g2_xnor2_1 _1203_ (.Y(\stop.syn.filt.m1.sum[15] ),
    .A(_0468_),
    .B(_0469_));
 sg13g2_nand2_1 _1204_ (.Y(_0470_),
    .A(\stop.syn.filt.m1.sum_in2[0] ),
    .B(\stop.syn.filt.m2.sum_in2[0] ));
 sg13g2_xor2_1 _1205_ (.B(\stop.syn.filt.m2.sum_in2[0] ),
    .A(\stop.syn.filt.m1.sum_in2[0] ),
    .X(_0054_));
 sg13g2_nand2_1 _1206_ (.Y(_0471_),
    .A(\stop.syn.filt.m1.sum_in2[1] ),
    .B(\stop.syn.filt.m2.sum_in2[1] ));
 sg13g2_nor2_1 _1207_ (.A(\stop.syn.filt.m1.sum_in2[1] ),
    .B(\stop.syn.filt.m2.sum_in2[1] ),
    .Y(_0472_));
 sg13g2_xor2_1 _1208_ (.B(\stop.syn.filt.m2.sum_in2[1] ),
    .A(\stop.syn.filt.m1.sum_in2[1] ),
    .X(_0473_));
 sg13g2_xnor2_1 _1209_ (.Y(_0061_),
    .A(_0470_),
    .B(_0473_));
 sg13g2_o21ai_1 _1210_ (.B1(_0471_),
    .Y(_0474_),
    .A1(_0470_),
    .A2(_0472_));
 sg13g2_and2_1 _1211_ (.A(\stop.syn.filt.m1.sum_in2[2] ),
    .B(\stop.syn.filt.m2.sum_in2[2] ),
    .X(_0475_));
 sg13g2_or2_1 _1212_ (.X(_0476_),
    .B(\stop.syn.filt.m2.sum_in2[2] ),
    .A(\stop.syn.filt.m1.sum_in2[2] ));
 sg13g2_nand2b_1 _1213_ (.Y(_0477_),
    .B(_0476_),
    .A_N(_0475_));
 sg13g2_xnor2_1 _1214_ (.Y(_0062_),
    .A(_0474_),
    .B(_0477_));
 sg13g2_a21o_1 _1215_ (.A2(_0476_),
    .A1(_0474_),
    .B1(_0475_),
    .X(_0478_));
 sg13g2_and2_1 _1216_ (.A(\stop.syn.filt.m1.sum_in2[3] ),
    .B(\stop.syn.filt.m2.sum_in2[3] ),
    .X(_0479_));
 sg13g2_or2_1 _1217_ (.X(_0480_),
    .B(\stop.syn.filt.m2.sum_in2[3] ),
    .A(\stop.syn.filt.m1.sum_in2[3] ));
 sg13g2_nand2b_1 _1218_ (.Y(_0481_),
    .B(_0480_),
    .A_N(_0479_));
 sg13g2_xnor2_1 _1219_ (.Y(_0063_),
    .A(_0478_),
    .B(_0481_));
 sg13g2_nand2_1 _1220_ (.Y(_0482_),
    .A(\stop.syn.filt.m1.sum_in2[4] ),
    .B(\stop.syn.filt.m2.sum_in2[4] ));
 sg13g2_xnor2_1 _1221_ (.Y(_0483_),
    .A(\stop.syn.filt.m1.sum_in2[4] ),
    .B(\stop.syn.filt.m2.sum_in2[4] ));
 sg13g2_a21oi_2 _1222_ (.B1(_0479_),
    .Y(_0484_),
    .A2(_0480_),
    .A1(_0478_));
 sg13g2_xor2_1 _1223_ (.B(_0484_),
    .A(_0483_),
    .X(_0064_));
 sg13g2_or2_1 _1224_ (.X(_0485_),
    .B(\stop.syn.filt.m2.sum_in2[5] ),
    .A(\stop.syn.filt.m1.sum_in2[5] ));
 sg13g2_xnor2_1 _1225_ (.Y(_0486_),
    .A(\stop.syn.filt.m1.sum_in2[5] ),
    .B(\stop.syn.filt.m2.sum_in2[5] ));
 sg13g2_o21ai_1 _1226_ (.B1(_0482_),
    .Y(_0487_),
    .A1(_0483_),
    .A2(_0484_));
 sg13g2_xnor2_1 _1227_ (.Y(_0065_),
    .A(_0486_),
    .B(_0487_));
 sg13g2_nand2_1 _1228_ (.Y(_0488_),
    .A(\stop.syn.filt.m1.sum_in2[6] ),
    .B(\stop.syn.filt.m2.sum_in2[6] ));
 sg13g2_xnor2_1 _1229_ (.Y(_0489_),
    .A(\stop.syn.filt.m1.sum_in2[6] ),
    .B(\stop.syn.filt.m2.sum_in2[6] ));
 sg13g2_inv_1 _1230_ (.Y(_0490_),
    .A(_0489_));
 sg13g2_a22oi_1 _1231_ (.Y(_0491_),
    .B1(\stop.syn.filt.m2.sum_in2[5] ),
    .B2(\stop.syn.filt.m1.sum_in2[5] ),
    .A2(\stop.syn.filt.m2.sum_in2[4] ),
    .A1(\stop.syn.filt.m1.sum_in2[4] ));
 sg13g2_o21ai_1 _1232_ (.B1(_0491_),
    .Y(_0492_),
    .A1(_0483_),
    .A2(_0484_));
 sg13g2_nand2_1 _1233_ (.Y(_0493_),
    .A(_0485_),
    .B(_0492_));
 sg13g2_nand3_1 _1234_ (.B(_0490_),
    .C(_0492_),
    .A(_0485_),
    .Y(_0494_));
 sg13g2_xnor2_1 _1235_ (.Y(_0066_),
    .A(_0490_),
    .B(_0493_));
 sg13g2_and2_1 _1236_ (.A(\stop.syn.filt.m1.sum_in2[7] ),
    .B(\stop.syn.filt.m2.sum_in2[7] ),
    .X(_0495_));
 sg13g2_xnor2_1 _1237_ (.Y(_0496_),
    .A(\stop.syn.filt.m1.sum_in2[7] ),
    .B(\stop.syn.filt.m2.sum_in2[7] ));
 sg13g2_a21oi_2 _1238_ (.B1(_0496_),
    .Y(_0497_),
    .A2(_0494_),
    .A1(_0488_));
 sg13g2_nand3_1 _1239_ (.B(_0494_),
    .C(_0496_),
    .A(_0488_),
    .Y(_0498_));
 sg13g2_nor2b_1 _1240_ (.A(_0497_),
    .B_N(_0498_),
    .Y(_0067_));
 sg13g2_nor2_1 _1241_ (.A(_0495_),
    .B(_0497_),
    .Y(_0499_));
 sg13g2_nand2_1 _1242_ (.Y(_0500_),
    .A(\stop.syn.filt.m1.sum_in2[8] ),
    .B(\stop.syn.filt.m2.sum_in2[8] ));
 sg13g2_xnor2_1 _1243_ (.Y(_0501_),
    .A(\stop.syn.filt.m1.sum_in2[8] ),
    .B(\stop.syn.filt.m2.sum_in2[8] ));
 sg13g2_xor2_1 _1244_ (.B(_0501_),
    .A(_0499_),
    .X(_0068_));
 sg13g2_xnor2_1 _1245_ (.Y(_0502_),
    .A(\stop.syn.filt.m1.sum_in2[9] ),
    .B(\stop.syn.filt.m2.sum_in2[9] ));
 sg13g2_o21ai_1 _1246_ (.B1(_0500_),
    .Y(_0503_),
    .A1(_0499_),
    .A2(_0501_));
 sg13g2_xnor2_1 _1247_ (.Y(_0069_),
    .A(_0502_),
    .B(_0503_));
 sg13g2_nand2_1 _1248_ (.Y(_0504_),
    .A(\stop.syn.filt.m1.sum_in2[10] ),
    .B(\stop.syn.filt.m2.sum_in2[10] ));
 sg13g2_nor2_1 _1249_ (.A(\stop.syn.filt.m1.sum_in2[10] ),
    .B(\stop.syn.filt.m2.sum_in2[10] ),
    .Y(_0505_));
 sg13g2_xor2_1 _1250_ (.B(\stop.syn.filt.m2.sum_in2[10] ),
    .A(\stop.syn.filt.m1.sum_in2[10] ),
    .X(_0506_));
 sg13g2_nor2_1 _1251_ (.A(_0501_),
    .B(_0502_),
    .Y(_0507_));
 sg13g2_o21ai_1 _1252_ (.B1(_0507_),
    .Y(_0508_),
    .A1(_0495_),
    .A2(_0497_));
 sg13g2_a22oi_1 _1253_ (.Y(_0509_),
    .B1(\stop.syn.filt.m2.sum_in2[9] ),
    .B2(\stop.syn.filt.m1.sum_in2[9] ),
    .A2(\stop.syn.filt.m2.sum_in2[8] ),
    .A1(\stop.syn.filt.m1.sum_in2[8] ));
 sg13g2_inv_1 _1254_ (.Y(_0510_),
    .A(_0509_));
 sg13g2_o21ai_1 _1255_ (.B1(_0510_),
    .Y(_0511_),
    .A1(\stop.syn.filt.m1.sum_in2[9] ),
    .A2(\stop.syn.filt.m2.sum_in2[9] ));
 sg13g2_and2_1 _1256_ (.A(_0508_),
    .B(_0511_),
    .X(_0512_));
 sg13g2_xnor2_1 _1257_ (.Y(_0055_),
    .A(_0506_),
    .B(_0512_));
 sg13g2_nor2_1 _1258_ (.A(\stop.syn.filt.m1.sum_in2[11] ),
    .B(\stop.syn.filt.m2.sum_in2[11] ),
    .Y(_0513_));
 sg13g2_nand2_1 _1259_ (.Y(_0514_),
    .A(\stop.syn.filt.m1.sum_in2[11] ),
    .B(\stop.syn.filt.m2.sum_in2[11] ));
 sg13g2_nand2b_1 _1260_ (.Y(_0515_),
    .B(_0514_),
    .A_N(_0513_));
 sg13g2_o21ai_1 _1261_ (.B1(_0504_),
    .Y(_0516_),
    .A1(_0505_),
    .A2(_0512_));
 sg13g2_xnor2_1 _1262_ (.Y(_0056_),
    .A(_0515_),
    .B(_0516_));
 sg13g2_and2_1 _1263_ (.A(\stop.syn.filt.m1.sum_in2[12] ),
    .B(\stop.syn.filt.m2.sum_in2[12] ),
    .X(_0517_));
 sg13g2_xor2_1 _1264_ (.B(\stop.syn.filt.m2.sum_in2[12] ),
    .A(\stop.syn.filt.m1.sum_in2[12] ),
    .X(_0518_));
 sg13g2_nand2_1 _1265_ (.Y(_0519_),
    .A(_0504_),
    .B(_0514_));
 sg13g2_nand2b_1 _1266_ (.Y(_0520_),
    .B(_0519_),
    .A_N(_0513_));
 sg13g2_and2_1 _1267_ (.A(_0511_),
    .B(_0520_),
    .X(_0521_));
 sg13g2_a221oi_1 _1268_ (.B2(_0508_),
    .C1(_0513_),
    .B1(_0521_),
    .A1(_0505_),
    .Y(_0522_),
    .A2(_0514_));
 sg13g2_xor2_1 _1269_ (.B(_0522_),
    .A(_0518_),
    .X(_0057_));
 sg13g2_nand2_1 _1270_ (.Y(_0523_),
    .A(\stop.syn.filt.m1.sum_in2[13] ),
    .B(\stop.syn.filt.m2.sum_in2[13] ));
 sg13g2_xor2_1 _1271_ (.B(\stop.syn.filt.m2.sum_in2[13] ),
    .A(\stop.syn.filt.m1.sum_in2[13] ),
    .X(_0524_));
 sg13g2_a21oi_1 _1272_ (.A1(_0518_),
    .A2(_0522_),
    .Y(_0525_),
    .B1(_0517_));
 sg13g2_xnor2_1 _1273_ (.Y(_0058_),
    .A(_0524_),
    .B(_0525_));
 sg13g2_and2_1 _1274_ (.A(_0518_),
    .B(_0524_),
    .X(_0526_));
 sg13g2_o21ai_1 _1275_ (.B1(_0517_),
    .Y(_0527_),
    .A1(\stop.syn.filt.m1.sum_in2[13] ),
    .A2(\stop.syn.filt.m2.sum_in2[13] ));
 sg13g2_nand2_1 _1276_ (.Y(_0528_),
    .A(_0523_),
    .B(_0527_));
 sg13g2_a21o_1 _1277_ (.A2(_0526_),
    .A1(_0522_),
    .B1(_0528_),
    .X(_0529_));
 sg13g2_and2_1 _1278_ (.A(\stop.syn.filt.m1.sum_in2[14] ),
    .B(\stop.syn.filt.m2.sum_in2[14] ),
    .X(_0530_));
 sg13g2_xor2_1 _1279_ (.B(\stop.syn.filt.m2.sum_in2[14] ),
    .A(\stop.syn.filt.m1.sum_in2[14] ),
    .X(_0531_));
 sg13g2_xor2_1 _1280_ (.B(_0531_),
    .A(_0529_),
    .X(_0059_));
 sg13g2_a21oi_1 _1281_ (.A1(_0529_),
    .A2(_0531_),
    .Y(_0532_),
    .B1(_0530_));
 sg13g2_xor2_1 _1282_ (.B(\stop.syn.filt.m2.sum_in2[15] ),
    .A(\stop.syn.filt.m1.sum_in2[15] ),
    .X(_0533_));
 sg13g2_xnor2_1 _1283_ (.Y(_0060_),
    .A(_0532_),
    .B(_0533_));
 sg13g2_nand2_2 _1284_ (.Y(_0534_),
    .A(\stop.syn.osci.data_buf ),
    .B(\stop.syn.smul8.b_bit ));
 sg13g2_xnor2_1 _1285_ (.Y(_0071_),
    .A(\stop.syn.adsr_data[8] ),
    .B(_0534_));
 sg13g2_nor3_2 _1286_ (.A(\stop.syn.adsr_data[8] ),
    .B(\stop.syn.adsr_data[9] ),
    .C(_0534_),
    .Y(_0535_));
 sg13g2_o21ai_1 _1287_ (.B1(\stop.syn.adsr_data[9] ),
    .Y(_0536_),
    .A1(\stop.syn.adsr_data[8] ),
    .A2(_0534_));
 sg13g2_nand2b_1 _1288_ (.Y(_0072_),
    .B(_0536_),
    .A_N(_0535_));
 sg13g2_nor2b_1 _1289_ (.A(\stop.syn.adsr_data[10] ),
    .B_N(_0535_),
    .Y(_0537_));
 sg13g2_xor2_1 _1290_ (.B(_0535_),
    .A(\stop.syn.adsr_data[10] ),
    .X(_0073_));
 sg13g2_nand2_1 _1291_ (.Y(_0538_),
    .A(_0052_),
    .B(_0537_));
 sg13g2_xnor2_1 _1292_ (.Y(_0074_),
    .A(_0052_),
    .B(_0537_));
 sg13g2_xnor2_1 _1293_ (.Y(_0075_),
    .A(\stop.syn.adsr_data[12] ),
    .B(_0538_));
 sg13g2_o21ai_1 _1294_ (.B1(_0312_),
    .Y(_0539_),
    .A1(\stop.syn.adsr_data[12] ),
    .A2(_0538_));
 sg13g2_or3_1 _1295_ (.A(\stop.syn.adsr_data[12] ),
    .B(_0312_),
    .C(_0538_),
    .X(_0540_));
 sg13g2_nand2_1 _1296_ (.Y(_0076_),
    .A(_0539_),
    .B(_0540_));
 sg13g2_nor2_1 _1297_ (.A(\stop.syn.adsr_data[14] ),
    .B(_0540_),
    .Y(_0541_));
 sg13g2_xnor2_1 _1298_ (.Y(_0077_),
    .A(\stop.syn.adsr_data[14] ),
    .B(_0540_));
 sg13g2_xor2_1 _1299_ (.B(_0541_),
    .A(\stop.syn.adsr_data[15] ),
    .X(_0078_));
 sg13g2_nand3_1 _1300_ (.B(net308),
    .C(\stop.syn.adsr_data_reg[0] ),
    .A(\stop.syn.filt.m2.sum_in2[0] ),
    .Y(_0542_));
 sg13g2_and3_1 _1301_ (.X(_0543_),
    .A(\stop.syn.filt.m2.sum_in2[1] ),
    .B(\stop.syn.adsr_data_reg[1] ),
    .C(net307));
 sg13g2_nand3_1 _1302_ (.B(\stop.syn.adsr_data_reg[1] ),
    .C(net307),
    .A(\stop.syn.filt.m2.sum_in2[1] ),
    .Y(_0544_));
 sg13g2_a21oi_1 _1303_ (.A1(\stop.syn.adsr_data_reg[1] ),
    .A2(net307),
    .Y(_0545_),
    .B1(\stop.syn.filt.m2.sum_in2[1] ));
 sg13g2_nor2_1 _1304_ (.A(_0543_),
    .B(_0545_),
    .Y(_0546_));
 sg13g2_xnor2_1 _1305_ (.Y(\stop.syn.filt.m2.sum[1] ),
    .A(_0542_),
    .B(_0546_));
 sg13g2_o21ai_1 _1306_ (.B1(_0544_),
    .Y(_0547_),
    .A1(_0542_),
    .A2(_0545_));
 sg13g2_and3_1 _1307_ (.X(_0548_),
    .A(\stop.syn.filt.m2.sum_in2[2] ),
    .B(net307),
    .C(\stop.syn.adsr_data_reg[2] ));
 sg13g2_a21o_1 _1308_ (.A2(\stop.syn.adsr_data_reg[2] ),
    .A1(net307),
    .B1(\stop.syn.filt.m2.sum_in2[2] ),
    .X(_0549_));
 sg13g2_nand2b_1 _1309_ (.Y(_0550_),
    .B(_0549_),
    .A_N(_0548_));
 sg13g2_xnor2_1 _1310_ (.Y(\stop.syn.filt.m2.sum[2] ),
    .A(_0547_),
    .B(_0550_));
 sg13g2_nand2_1 _1311_ (.Y(_0551_),
    .A(net308),
    .B(\stop.syn.adsr_data_reg[3] ));
 sg13g2_nor2_1 _1312_ (.A(_0043_),
    .B(_0551_),
    .Y(_0552_));
 sg13g2_xor2_1 _1313_ (.B(_0551_),
    .A(_0043_),
    .X(_0553_));
 sg13g2_a21o_1 _1314_ (.A2(_0549_),
    .A1(_0547_),
    .B1(_0548_),
    .X(_0554_));
 sg13g2_xor2_1 _1315_ (.B(_0554_),
    .A(_0553_),
    .X(\stop.syn.filt.m2.sum[3] ));
 sg13g2_a21oi_2 _1316_ (.B1(_0552_),
    .Y(_0555_),
    .A2(_0554_),
    .A1(_0553_));
 sg13g2_nand3_1 _1317_ (.B(net307),
    .C(\stop.syn.adsr_data_reg[4] ),
    .A(\stop.syn.filt.m2.sum_in2[4] ),
    .Y(_0556_));
 sg13g2_a21o_1 _1318_ (.A2(\stop.syn.adsr_data_reg[4] ),
    .A1(net307),
    .B1(\stop.syn.filt.m2.sum_in2[4] ),
    .X(_0557_));
 sg13g2_nand2_1 _1319_ (.Y(_0558_),
    .A(_0556_),
    .B(_0557_));
 sg13g2_xor2_1 _1320_ (.B(_0558_),
    .A(_0555_),
    .X(\stop.syn.filt.m2.sum[4] ));
 sg13g2_nand2_1 _1321_ (.Y(_0559_),
    .A(net307),
    .B(\stop.syn.adsr_data_reg[5] ));
 sg13g2_nor2_1 _1322_ (.A(_0044_),
    .B(_0559_),
    .Y(_0560_));
 sg13g2_xor2_1 _1323_ (.B(_0559_),
    .A(_0044_),
    .X(_0561_));
 sg13g2_o21ai_1 _1324_ (.B1(_0556_),
    .Y(_0562_),
    .A1(_0555_),
    .A2(_0558_));
 sg13g2_xor2_1 _1325_ (.B(_0562_),
    .A(_0561_),
    .X(\stop.syn.filt.m2.sum[5] ));
 sg13g2_and3_1 _1326_ (.X(_0563_),
    .A(\stop.syn.filt.m2.sum_in2[6] ),
    .B(net306),
    .C(\stop.syn.adsr_data_reg[6] ));
 sg13g2_a21o_1 _1327_ (.A2(\stop.syn.adsr_data_reg[6] ),
    .A1(net306),
    .B1(\stop.syn.filt.m2.sum_in2[6] ),
    .X(_0564_));
 sg13g2_nand2b_1 _1328_ (.Y(_0565_),
    .B(_0564_),
    .A_N(_0563_));
 sg13g2_nand2b_1 _1329_ (.Y(_0566_),
    .B(_0561_),
    .A_N(_0558_));
 sg13g2_a21oi_1 _1330_ (.A1(_0044_),
    .A2(_0559_),
    .Y(_0567_),
    .B1(_0556_));
 sg13g2_nor2_1 _1331_ (.A(_0560_),
    .B(_0567_),
    .Y(_0568_));
 sg13g2_o21ai_1 _1332_ (.B1(_0568_),
    .Y(_0569_),
    .A1(_0555_),
    .A2(_0566_));
 sg13g2_xnor2_1 _1333_ (.Y(\stop.syn.filt.m2.sum[6] ),
    .A(_0565_),
    .B(_0569_));
 sg13g2_a21oi_2 _1334_ (.B1(_0563_),
    .Y(_0570_),
    .A2(_0569_),
    .A1(_0564_));
 sg13g2_nand3_1 _1335_ (.B(net306),
    .C(\stop.syn.adsr_data_reg[7] ),
    .A(\stop.syn.filt.m2.sum_in2[7] ),
    .Y(_0571_));
 sg13g2_a21o_1 _1336_ (.A2(\stop.syn.adsr_data_reg[7] ),
    .A1(net306),
    .B1(\stop.syn.filt.m2.sum_in2[7] ),
    .X(_0572_));
 sg13g2_nand2_1 _1337_ (.Y(_0573_),
    .A(_0571_),
    .B(_0572_));
 sg13g2_xor2_1 _1338_ (.B(_0573_),
    .A(_0570_),
    .X(\stop.syn.filt.m2.sum[7] ));
 sg13g2_o21ai_1 _1339_ (.B1(_0571_),
    .Y(_0574_),
    .A1(_0570_),
    .A2(_0573_));
 sg13g2_inv_1 _1340_ (.Y(_0575_),
    .A(_0574_));
 sg13g2_nand3_1 _1341_ (.B(net306),
    .C(\stop.syn.adsr_data_reg[8] ),
    .A(\stop.syn.filt.m2.sum_in2[8] ),
    .Y(_0576_));
 sg13g2_a21o_1 _1342_ (.A2(\stop.syn.adsr_data_reg[8] ),
    .A1(net306),
    .B1(\stop.syn.filt.m2.sum_in2[8] ),
    .X(_0577_));
 sg13g2_nand2_1 _1343_ (.Y(_0578_),
    .A(_0576_),
    .B(_0577_));
 sg13g2_xnor2_1 _1344_ (.Y(\stop.syn.filt.m2.sum[8] ),
    .A(_0574_),
    .B(_0578_));
 sg13g2_nand2_1 _1345_ (.Y(_0579_),
    .A(net306),
    .B(\stop.syn.adsr_data_reg[9] ));
 sg13g2_nand2_1 _1346_ (.Y(_0580_),
    .A(_0045_),
    .B(_0579_));
 sg13g2_xor2_1 _1347_ (.B(_0579_),
    .A(_0045_),
    .X(_0581_));
 sg13g2_o21ai_1 _1348_ (.B1(_0576_),
    .Y(_0582_),
    .A1(_0575_),
    .A2(_0578_));
 sg13g2_xor2_1 _1349_ (.B(_0582_),
    .A(_0581_),
    .X(\stop.syn.filt.m2.sum[9] ));
 sg13g2_nand3_1 _1350_ (.B(net304),
    .C(\stop.syn.adsr_data_reg[10] ),
    .A(\stop.syn.filt.m2.sum_in2[10] ),
    .Y(_0583_));
 sg13g2_a21o_1 _1351_ (.A2(\stop.syn.adsr_data_reg[10] ),
    .A1(net304),
    .B1(\stop.syn.filt.m2.sum_in2[10] ),
    .X(_0584_));
 sg13g2_nand2_1 _1352_ (.Y(_0585_),
    .A(_0583_),
    .B(_0584_));
 sg13g2_nand2b_1 _1353_ (.Y(_0586_),
    .B(_0581_),
    .A_N(_0578_));
 sg13g2_nand2b_1 _1354_ (.Y(_0587_),
    .B(_0574_),
    .A_N(_0586_));
 sg13g2_o21ai_1 _1355_ (.B1(_0576_),
    .Y(_0588_),
    .A1(_0045_),
    .A2(_0579_));
 sg13g2_nand2_1 _1356_ (.Y(_0589_),
    .A(_0580_),
    .B(_0588_));
 sg13g2_and2_1 _1357_ (.A(_0587_),
    .B(_0589_),
    .X(_0590_));
 sg13g2_xor2_1 _1358_ (.B(_0590_),
    .A(_0585_),
    .X(\stop.syn.filt.m2.sum[10] ));
 sg13g2_a21o_1 _1359_ (.A2(\stop.syn.adsr_data_reg[11] ),
    .A1(net304),
    .B1(\stop.syn.filt.m2.sum_in2[11] ),
    .X(_0591_));
 sg13g2_nand3_1 _1360_ (.B(net304),
    .C(\stop.syn.adsr_data_reg[11] ),
    .A(\stop.syn.filt.m2.sum_in2[11] ),
    .Y(_0592_));
 sg13g2_nand2_1 _1361_ (.Y(_0593_),
    .A(_0591_),
    .B(_0592_));
 sg13g2_o21ai_1 _1362_ (.B1(_0583_),
    .Y(_0594_),
    .A1(_0585_),
    .A2(_0590_));
 sg13g2_xnor2_1 _1363_ (.Y(\stop.syn.filt.m2.sum[11] ),
    .A(_0593_),
    .B(_0594_));
 sg13g2_nand3_1 _1364_ (.B(net304),
    .C(\stop.syn.adsr_data_reg[12] ),
    .A(\stop.syn.filt.m2.sum_in2[12] ),
    .Y(_0595_));
 sg13g2_a21o_1 _1365_ (.A2(\stop.syn.adsr_data_reg[12] ),
    .A1(net304),
    .B1(\stop.syn.filt.m2.sum_in2[12] ),
    .X(_0596_));
 sg13g2_nand2_1 _1366_ (.Y(_0597_),
    .A(_0595_),
    .B(_0596_));
 sg13g2_nand2_1 _1367_ (.Y(_0598_),
    .A(_0583_),
    .B(_0592_));
 sg13g2_or2_1 _1368_ (.X(_0599_),
    .B(_0593_),
    .A(_0585_));
 sg13g2_nor2_1 _1369_ (.A(_0589_),
    .B(_0599_),
    .Y(_0600_));
 sg13g2_nor2_1 _1370_ (.A(_0586_),
    .B(_0599_),
    .Y(_0601_));
 sg13g2_a221oi_1 _1371_ (.B2(_0574_),
    .C1(_0600_),
    .B1(_0601_),
    .A1(_0591_),
    .Y(_0602_),
    .A2(_0598_));
 sg13g2_xor2_1 _1372_ (.B(_0602_),
    .A(_0597_),
    .X(\stop.syn.filt.m2.sum[12] ));
 sg13g2_nand2_1 _1373_ (.Y(_0603_),
    .A(net304),
    .B(\stop.syn.adsr_data_reg[13] ));
 sg13g2_nor2_1 _1374_ (.A(_0046_),
    .B(_0603_),
    .Y(_0604_));
 sg13g2_xor2_1 _1375_ (.B(_0603_),
    .A(_0046_),
    .X(_0605_));
 sg13g2_o21ai_1 _1376_ (.B1(_0595_),
    .Y(_0606_),
    .A1(_0597_),
    .A2(_0602_));
 sg13g2_xor2_1 _1377_ (.B(_0606_),
    .A(_0605_),
    .X(\stop.syn.filt.m2.sum[13] ));
 sg13g2_nand2b_1 _1378_ (.Y(_0607_),
    .B(_0605_),
    .A_N(_0597_));
 sg13g2_a21oi_1 _1379_ (.A1(_0046_),
    .A2(_0603_),
    .Y(_0608_),
    .B1(_0595_));
 sg13g2_nor2_1 _1380_ (.A(_0604_),
    .B(_0608_),
    .Y(_0609_));
 sg13g2_o21ai_1 _1381_ (.B1(_0609_),
    .Y(_0610_),
    .A1(_0602_),
    .A2(_0607_));
 sg13g2_nand3_1 _1382_ (.B(net305),
    .C(\stop.syn.adsr_data_reg[14] ),
    .A(\stop.syn.filt.m2.sum_in2[14] ),
    .Y(_0611_));
 sg13g2_a21o_1 _1383_ (.A2(\stop.syn.adsr_data_reg[14] ),
    .A1(net305),
    .B1(\stop.syn.filt.m2.sum_in2[14] ),
    .X(_0612_));
 sg13g2_nand2_1 _1384_ (.Y(_0613_),
    .A(_0611_),
    .B(_0612_));
 sg13g2_nand2b_1 _1385_ (.Y(_0614_),
    .B(_0610_),
    .A_N(_0613_));
 sg13g2_xnor2_1 _1386_ (.Y(\stop.syn.filt.m2.sum[14] ),
    .A(_0610_),
    .B(_0613_));
 sg13g2_and3_1 _1387_ (.X(_0615_),
    .A(\stop.syn.filt.m2.sum_in2[15] ),
    .B(net305),
    .C(\stop.syn.adsr_data_reg[15] ));
 sg13g2_a21oi_1 _1388_ (.A1(net304),
    .A2(\stop.syn.adsr_data_reg[15] ),
    .Y(_0616_),
    .B1(\stop.syn.filt.m2.sum_in2[15] ));
 sg13g2_nor2_1 _1389_ (.A(_0615_),
    .B(_0616_),
    .Y(_0617_));
 sg13g2_nand2_1 _1390_ (.Y(_0618_),
    .A(_0611_),
    .B(_0614_));
 sg13g2_xor2_1 _1391_ (.B(_0618_),
    .A(_0617_),
    .X(\stop.syn.filt.m2.sum[15] ));
 sg13g2_a21oi_1 _1392_ (.A1(_0466_),
    .A2(_0469_),
    .Y(\stop.syn.filt.m1.sum[16] ),
    .B1(_0467_));
 sg13g2_nor4_1 _1393_ (.A(\stop.syn.adsr_data[12] ),
    .B(_0312_),
    .C(\stop.syn.adsr_data[14] ),
    .D(\stop.syn.adsr_data[15] ),
    .Y(_0619_));
 sg13g2_nor4_1 _1394_ (.A(\stop.syn.adsr_data[8] ),
    .B(\stop.syn.adsr_data[9] ),
    .C(\stop.syn.adsr_data[10] ),
    .D(_0311_),
    .Y(_0620_));
 sg13g2_a21oi_1 _1395_ (.A1(_0619_),
    .A2(_0620_),
    .Y(_0070_),
    .B1(_0534_));
 sg13g2_a21oi_1 _1396_ (.A1(_0611_),
    .A2(_0614_),
    .Y(_0621_),
    .B1(_0616_));
 sg13g2_or2_1 _1397_ (.X(\stop.syn.filt.m2.sum[16] ),
    .B(_0621_),
    .A(_0615_));
 sg13g2_nand2b_1 _1398_ (.Y(\stop.syn.clki.arstn ),
    .B(\stop.syn.rstn_fst_reg2 ),
    .A_N(\stop.syn.rstn_fst_reg1 ));
 sg13g2_o21ai_1 _1399_ (.B1(net362),
    .Y(_0622_),
    .A1(net2),
    .A2(\stop.ctrl.first_bit_reg ));
 sg13g2_inv_2 _1400_ (.Y(\stop.merge_rstn ),
    .A(_0622_));
 sg13g2_or2_1 _1401_ (.X(\stop.merge_trig ),
    .B(net1),
    .A(\stop.ctrl.trig ));
 sg13g2_nor2_1 _1402_ (.A(_0082_),
    .B(net2),
    .Y(_0623_));
 sg13g2_mux2_1 _1403_ (.A0(\stop.ctrl.trig ),
    .A1(net3),
    .S(_0623_),
    .X(_0135_));
 sg13g2_nand2_1 _1404_ (.Y(_0624_),
    .A(_0301_),
    .B(_0379_));
 sg13g2_o21ai_1 _1405_ (.B1(net281),
    .Y(_0625_),
    .A1(_0389_),
    .A2(_0624_));
 sg13g2_or4_2 _1406_ (.A(_0302_),
    .B(net283),
    .C(_0380_),
    .D(_0624_),
    .X(_0626_));
 sg13g2_a21oi_1 _1407_ (.A1(_0366_),
    .A2(_0626_),
    .Y(_0136_),
    .B1(_0625_));
 sg13g2_a21oi_1 _1408_ (.A1(_0364_),
    .A2(_0626_),
    .Y(_0137_),
    .B1(_0625_));
 sg13g2_a21oi_1 _1409_ (.A1(_0363_),
    .A2(_0626_),
    .Y(_0138_),
    .B1(_0625_));
 sg13g2_a21oi_1 _1410_ (.A1(_0362_),
    .A2(_0626_),
    .Y(_0139_),
    .B1(_0625_));
 sg13g2_a21oi_1 _1411_ (.A1(_0360_),
    .A2(_0626_),
    .Y(_0140_),
    .B1(_0625_));
 sg13g2_a21oi_1 _1412_ (.A1(_0359_),
    .A2(_0626_),
    .Y(_0141_),
    .B1(_0625_));
 sg13g2_a21oi_1 _1413_ (.A1(_0358_),
    .A2(_0626_),
    .Y(_0142_),
    .B1(_0625_));
 sg13g2_a21oi_1 _1414_ (.A1(_0356_),
    .A2(_0626_),
    .Y(_0143_),
    .B1(_0625_));
 sg13g2_xnor2_1 _1415_ (.Y(_0627_),
    .A(\stop.ctrl.cfg[35] ),
    .B(\stop.syn.osci.counter[3] ));
 sg13g2_xnor2_1 _1416_ (.Y(_0628_),
    .A(\stop.ctrl.cfg[43] ),
    .B(\stop.syn.osci.counter[11] ));
 sg13g2_xnor2_1 _1417_ (.Y(_0629_),
    .A(\stop.ctrl.cfg[32] ),
    .B(\stop.syn.osci.counter[0] ));
 sg13g2_xnor2_1 _1418_ (.Y(_0630_),
    .A(\stop.ctrl.cfg[37] ),
    .B(\stop.syn.osci.counter[5] ));
 sg13g2_xnor2_1 _1419_ (.Y(_0631_),
    .A(\stop.ctrl.cfg[33] ),
    .B(\stop.syn.osci.counter[1] ));
 sg13g2_xnor2_1 _1420_ (.Y(_0632_),
    .A(\stop.ctrl.cfg[42] ),
    .B(\stop.syn.osci.counter[10] ));
 sg13g2_xnor2_1 _1421_ (.Y(_0633_),
    .A(\stop.ctrl.cfg[39] ),
    .B(\stop.syn.osci.counter[7] ));
 sg13g2_xnor2_1 _1422_ (.Y(_0634_),
    .A(\stop.ctrl.cfg[38] ),
    .B(\stop.syn.osci.counter[6] ));
 sg13g2_xnor2_1 _1423_ (.Y(_0635_),
    .A(\stop.ctrl.cfg[36] ),
    .B(\stop.syn.osci.counter[4] ));
 sg13g2_xnor2_1 _1424_ (.Y(_0636_),
    .A(\stop.ctrl.cfg[40] ),
    .B(\stop.syn.osci.counter[8] ));
 sg13g2_xnor2_1 _1425_ (.Y(_0637_),
    .A(\stop.ctrl.cfg[41] ),
    .B(\stop.syn.osci.counter[9] ));
 sg13g2_xnor2_1 _1426_ (.Y(_0638_),
    .A(\stop.ctrl.cfg[34] ),
    .B(\stop.syn.osci.counter[2] ));
 sg13g2_nand4_1 _1427_ (.B(_0632_),
    .C(_0633_),
    .A(_0631_),
    .Y(_0639_),
    .D(_0636_));
 sg13g2_nand4_1 _1428_ (.B(_0628_),
    .C(_0634_),
    .A(_0627_),
    .Y(_0640_),
    .D(_0637_));
 sg13g2_nand4_1 _1429_ (.B(_0630_),
    .C(_0635_),
    .A(_0629_),
    .Y(_0641_),
    .D(_0638_));
 sg13g2_nor3_1 _1430_ (.A(_0639_),
    .B(_0640_),
    .C(_0641_),
    .Y(_0642_));
 sg13g2_or2_1 _1431_ (.X(_0643_),
    .B(_0642_),
    .A(_0047_));
 sg13g2_inv_2 _1432_ (.Y(_0644_),
    .A(net278));
 sg13g2_and2_1 _1433_ (.A(_0079_),
    .B(_0644_),
    .X(_0144_));
 sg13g2_xnor2_1 _1434_ (.Y(_0645_),
    .A(\stop.syn.osci.counter[0] ),
    .B(\stop.syn.osci.counter[1] ));
 sg13g2_nor2_1 _1435_ (.A(net278),
    .B(_0645_),
    .Y(_0145_));
 sg13g2_and3_1 _1436_ (.X(_0646_),
    .A(\stop.syn.osci.counter[0] ),
    .B(\stop.syn.osci.counter[1] ),
    .C(\stop.syn.osci.counter[2] ));
 sg13g2_a21oi_1 _1437_ (.A1(\stop.syn.osci.counter[0] ),
    .A2(\stop.syn.osci.counter[1] ),
    .Y(_0647_),
    .B1(\stop.syn.osci.counter[2] ));
 sg13g2_nor3_1 _1438_ (.A(net278),
    .B(_0646_),
    .C(_0647_),
    .Y(_0146_));
 sg13g2_nor2_1 _1439_ (.A(\stop.syn.osci.counter[3] ),
    .B(_0646_),
    .Y(_0648_));
 sg13g2_and2_1 _1440_ (.A(\stop.syn.osci.counter[3] ),
    .B(_0646_),
    .X(_0649_));
 sg13g2_nor3_1 _1441_ (.A(net278),
    .B(_0648_),
    .C(_0649_),
    .Y(_0147_));
 sg13g2_nor2_1 _1442_ (.A(\stop.syn.osci.counter[4] ),
    .B(_0649_),
    .Y(_0650_));
 sg13g2_and2_1 _1443_ (.A(\stop.syn.osci.counter[4] ),
    .B(_0649_),
    .X(_0651_));
 sg13g2_nor3_1 _1444_ (.A(net278),
    .B(_0650_),
    .C(_0651_),
    .Y(_0148_));
 sg13g2_nor2_1 _1445_ (.A(\stop.syn.osci.counter[5] ),
    .B(_0651_),
    .Y(_0652_));
 sg13g2_and2_1 _1446_ (.A(\stop.syn.osci.counter[5] ),
    .B(_0651_),
    .X(_0653_));
 sg13g2_nor3_1 _1447_ (.A(net278),
    .B(_0652_),
    .C(_0653_),
    .Y(_0149_));
 sg13g2_nor2_1 _1448_ (.A(\stop.syn.osci.counter[6] ),
    .B(_0653_),
    .Y(_0654_));
 sg13g2_and2_1 _1449_ (.A(\stop.syn.osci.counter[6] ),
    .B(_0653_),
    .X(_0655_));
 sg13g2_nor3_1 _1450_ (.A(net278),
    .B(_0654_),
    .C(_0655_),
    .Y(_0150_));
 sg13g2_and2_1 _1451_ (.A(\stop.syn.osci.counter[7] ),
    .B(_0655_),
    .X(_0656_));
 sg13g2_o21ai_1 _1452_ (.B1(_0644_),
    .Y(_0657_),
    .A1(\stop.syn.osci.counter[7] ),
    .A2(_0655_));
 sg13g2_nor2_1 _1453_ (.A(_0656_),
    .B(_0657_),
    .Y(_0151_));
 sg13g2_and2_1 _1454_ (.A(\stop.syn.osci.counter[8] ),
    .B(_0656_),
    .X(_0658_));
 sg13g2_o21ai_1 _1455_ (.B1(_0644_),
    .Y(_0659_),
    .A1(\stop.syn.osci.counter[8] ),
    .A2(_0656_));
 sg13g2_nor2_1 _1456_ (.A(_0658_),
    .B(_0659_),
    .Y(_0152_));
 sg13g2_and2_1 _1457_ (.A(\stop.syn.osci.counter[9] ),
    .B(_0658_),
    .X(_0660_));
 sg13g2_o21ai_1 _1458_ (.B1(_0644_),
    .Y(_0661_),
    .A1(\stop.syn.osci.counter[9] ),
    .A2(_0658_));
 sg13g2_nor2_1 _1459_ (.A(_0660_),
    .B(_0661_),
    .Y(_0153_));
 sg13g2_nor2_1 _1460_ (.A(\stop.syn.osci.counter[10] ),
    .B(_0660_),
    .Y(_0662_));
 sg13g2_and2_1 _1461_ (.A(\stop.syn.osci.counter[10] ),
    .B(_0660_),
    .X(_0663_));
 sg13g2_nor3_1 _1462_ (.A(_0643_),
    .B(_0662_),
    .C(_0663_),
    .Y(_0154_));
 sg13g2_a21oi_1 _1463_ (.A1(\stop.syn.osci.counter[11] ),
    .A2(_0663_),
    .Y(_0664_),
    .B1(net278));
 sg13g2_o21ai_1 _1464_ (.B1(_0664_),
    .Y(_0665_),
    .A1(\stop.syn.osci.counter[11] ),
    .A2(_0663_));
 sg13g2_inv_1 _1465_ (.Y(_0155_),
    .A(_0665_));
 sg13g2_a22oi_1 _1466_ (.Y(_0666_),
    .B1(_0644_),
    .B2(\stop.syn.osci.data_buf ),
    .A2(_0642_),
    .A1(_0042_));
 sg13g2_inv_1 _1467_ (.Y(_0157_),
    .A(_0666_));
 sg13g2_or2_1 _1468_ (.X(_0667_),
    .B(net119),
    .A(\stop.syn.daci.din[0] ));
 sg13g2_nand2_1 _1469_ (.Y(_0668_),
    .A(\stop.syn.daci.din[0] ),
    .B(net119));
 sg13g2_and3_1 _1470_ (.X(_0159_),
    .A(net281),
    .B(_0667_),
    .C(_0668_));
 sg13g2_nand2_1 _1471_ (.Y(_0669_),
    .A(\stop.syn.daci.din[1] ),
    .B(\stop.syn.daci.accumulator[1] ));
 sg13g2_xnor2_1 _1472_ (.Y(_0670_),
    .A(\stop.syn.daci.din[1] ),
    .B(\stop.syn.daci.accumulator[1] ));
 sg13g2_o21ai_1 _1473_ (.B1(net281),
    .Y(_0671_),
    .A1(_0668_),
    .A2(_0670_));
 sg13g2_a21oi_1 _1474_ (.A1(_0668_),
    .A2(_0670_),
    .Y(_0160_),
    .B1(_0671_));
 sg13g2_and2_1 _1475_ (.A(\stop.syn.daci.din[2] ),
    .B(\stop.syn.daci.accumulator[2] ),
    .X(_0672_));
 sg13g2_xor2_1 _1476_ (.B(net139),
    .A(\stop.syn.daci.din[2] ),
    .X(_0673_));
 sg13g2_o21ai_1 _1477_ (.B1(_0669_),
    .Y(_0674_),
    .A1(_0668_),
    .A2(_0670_));
 sg13g2_or2_1 _1478_ (.X(_0675_),
    .B(_0674_),
    .A(_0673_));
 sg13g2_nand2_1 _1479_ (.Y(_0676_),
    .A(_0673_),
    .B(_0674_));
 sg13g2_and3_1 _1480_ (.X(_0161_),
    .A(net280),
    .B(_0675_),
    .C(net140));
 sg13g2_nand2_1 _1481_ (.Y(_0677_),
    .A(\stop.syn.daci.din[3] ),
    .B(\stop.syn.daci.accumulator[3] ));
 sg13g2_xnor2_1 _1482_ (.Y(_0678_),
    .A(\stop.syn.daci.din[3] ),
    .B(net124));
 sg13g2_a21oi_1 _1483_ (.A1(_0673_),
    .A2(_0674_),
    .Y(_0679_),
    .B1(_0672_));
 sg13g2_o21ai_1 _1484_ (.B1(net280),
    .Y(_0680_),
    .A1(_0678_),
    .A2(_0679_));
 sg13g2_a21oi_1 _1485_ (.A1(_0678_),
    .A2(_0679_),
    .Y(_0162_),
    .B1(_0680_));
 sg13g2_o21ai_1 _1486_ (.B1(_0677_),
    .Y(_0681_),
    .A1(_0678_),
    .A2(_0679_));
 sg13g2_nand2_1 _1487_ (.Y(_0682_),
    .A(\stop.syn.daci.din[4] ),
    .B(\stop.syn.daci.accumulator[4] ));
 sg13g2_xnor2_1 _1488_ (.Y(_0683_),
    .A(\stop.syn.daci.din[4] ),
    .B(net141));
 sg13g2_nand2b_1 _1489_ (.Y(_0684_),
    .B(_0683_),
    .A_N(_0681_));
 sg13g2_nand2b_1 _1490_ (.Y(_0685_),
    .B(_0681_),
    .A_N(_0683_));
 sg13g2_and3_1 _1491_ (.X(_0163_),
    .A(net280),
    .B(_0684_),
    .C(_0685_));
 sg13g2_nor2_1 _1492_ (.A(\stop.syn.daci.din[5] ),
    .B(\stop.syn.daci.accumulator[5] ),
    .Y(_0686_));
 sg13g2_xnor2_1 _1493_ (.Y(_0687_),
    .A(\stop.syn.daci.din[5] ),
    .B(net134));
 sg13g2_and2_1 _1494_ (.A(_0682_),
    .B(_0685_),
    .X(_0688_));
 sg13g2_o21ai_1 _1495_ (.B1(net280),
    .Y(_0689_),
    .A1(_0687_),
    .A2(_0688_));
 sg13g2_a21oi_1 _1496_ (.A1(_0687_),
    .A2(_0688_),
    .Y(_0164_),
    .B1(_0689_));
 sg13g2_nand2_1 _1497_ (.Y(_0690_),
    .A(\stop.syn.daci.din[6] ),
    .B(net130));
 sg13g2_xnor2_1 _1498_ (.Y(_0691_),
    .A(\stop.syn.daci.din[6] ),
    .B(net130));
 sg13g2_nor2_1 _1499_ (.A(_0682_),
    .B(_0686_),
    .Y(_0692_));
 sg13g2_nor2_1 _1500_ (.A(_0683_),
    .B(_0687_),
    .Y(_0693_));
 sg13g2_a221oi_1 _1501_ (.B2(_0693_),
    .C1(_0692_),
    .B1(_0681_),
    .A1(\stop.syn.daci.din[5] ),
    .Y(_0694_),
    .A2(\stop.syn.daci.accumulator[5] ));
 sg13g2_o21ai_1 _1502_ (.B1(net279),
    .Y(_0695_),
    .A1(_0691_),
    .A2(_0694_));
 sg13g2_a21oi_1 _1503_ (.A1(_0691_),
    .A2(_0694_),
    .Y(_0165_),
    .B1(_0695_));
 sg13g2_o21ai_1 _1504_ (.B1(_0690_),
    .Y(_0236_),
    .A1(_0691_),
    .A2(_0694_));
 sg13g2_and2_1 _1505_ (.A(\stop.syn.daci.din[7] ),
    .B(\stop.syn.daci.accumulator[7] ),
    .X(_0237_));
 sg13g2_xor2_1 _1506_ (.B(net138),
    .A(\stop.syn.daci.din[7] ),
    .X(_0238_));
 sg13g2_o21ai_1 _1507_ (.B1(net279),
    .Y(_0239_),
    .A1(_0236_),
    .A2(_0238_));
 sg13g2_a21oi_1 _1508_ (.A1(_0236_),
    .A2(_0238_),
    .Y(_0166_),
    .B1(_0239_));
 sg13g2_a21oi_2 _1509_ (.B1(_0237_),
    .Y(_0240_),
    .A2(_0238_),
    .A1(_0236_));
 sg13g2_a21o_1 _1510_ (.A2(_0238_),
    .A1(_0236_),
    .B1(_0237_),
    .X(_0241_));
 sg13g2_nand2_1 _1511_ (.Y(_0242_),
    .A(\stop.syn.daci.din[8] ),
    .B(net132));
 sg13g2_xnor2_1 _1512_ (.Y(_0243_),
    .A(\stop.syn.daci.din[8] ),
    .B(net132));
 sg13g2_nand2b_1 _1513_ (.Y(_0244_),
    .B(_0241_),
    .A_N(_0243_));
 sg13g2_nand2_1 _1514_ (.Y(_0245_),
    .A(net279),
    .B(_0244_));
 sg13g2_a21oi_1 _1515_ (.A1(_0240_),
    .A2(_0243_),
    .Y(_0167_),
    .B1(_0245_));
 sg13g2_nor2_1 _1516_ (.A(\stop.syn.daci.din[9] ),
    .B(net136),
    .Y(_0246_));
 sg13g2_nand2_1 _1517_ (.Y(_0247_),
    .A(\stop.syn.daci.din[9] ),
    .B(net136));
 sg13g2_nand2b_1 _1518_ (.Y(_0248_),
    .B(_0247_),
    .A_N(_0246_));
 sg13g2_nand3_1 _1519_ (.B(_0244_),
    .C(_0248_),
    .A(_0242_),
    .Y(_0249_));
 sg13g2_a21oi_1 _1520_ (.A1(_0242_),
    .A2(_0244_),
    .Y(_0250_),
    .B1(_0248_));
 sg13g2_nand2_1 _1521_ (.Y(_0251_),
    .A(net279),
    .B(_0249_));
 sg13g2_nor2_1 _1522_ (.A(_0250_),
    .B(_0251_),
    .Y(_0168_));
 sg13g2_nand2_1 _1523_ (.Y(_0252_),
    .A(\stop.syn.daci.din[10] ),
    .B(net128));
 sg13g2_xnor2_1 _1524_ (.Y(_0253_),
    .A(\stop.syn.daci.din[10] ),
    .B(net128));
 sg13g2_o21ai_1 _1525_ (.B1(_0247_),
    .Y(_0254_),
    .A1(_0242_),
    .A2(_0246_));
 sg13g2_nor2_1 _1526_ (.A(_0243_),
    .B(_0248_),
    .Y(_0255_));
 sg13g2_a21oi_1 _1527_ (.A1(_0241_),
    .A2(_0255_),
    .Y(_0256_),
    .B1(_0254_));
 sg13g2_or2_1 _1528_ (.X(_0257_),
    .B(_0256_),
    .A(_0253_));
 sg13g2_nand2_1 _1529_ (.Y(_0258_),
    .A(net280),
    .B(_0257_));
 sg13g2_a21oi_1 _1530_ (.A1(_0253_),
    .A2(_0256_),
    .Y(_0169_),
    .B1(_0258_));
 sg13g2_nor2_1 _1531_ (.A(\stop.syn.daci.din[11] ),
    .B(\stop.syn.daci.accumulator[11] ),
    .Y(_0259_));
 sg13g2_xnor2_1 _1532_ (.Y(_0260_),
    .A(\stop.syn.daci.din[11] ),
    .B(net137));
 sg13g2_nand3_1 _1533_ (.B(_0257_),
    .C(_0260_),
    .A(_0252_),
    .Y(_0261_));
 sg13g2_a21oi_1 _1534_ (.A1(_0252_),
    .A2(_0257_),
    .Y(_0262_),
    .B1(_0260_));
 sg13g2_nand2_1 _1535_ (.Y(_0263_),
    .A(net280),
    .B(_0261_));
 sg13g2_nor2_1 _1536_ (.A(_0262_),
    .B(_0263_),
    .Y(_0170_));
 sg13g2_nor2_1 _1537_ (.A(_0253_),
    .B(_0260_),
    .Y(_0264_));
 sg13g2_nand2_1 _1538_ (.Y(_0265_),
    .A(_0255_),
    .B(_0264_));
 sg13g2_nor2_1 _1539_ (.A(_0240_),
    .B(_0265_),
    .Y(_0266_));
 sg13g2_nor2_1 _1540_ (.A(_0252_),
    .B(_0259_),
    .Y(_0267_));
 sg13g2_a221oi_1 _1541_ (.B2(_0264_),
    .C1(_0267_),
    .B1(_0254_),
    .A1(\stop.syn.daci.din[11] ),
    .Y(_0268_),
    .A2(\stop.syn.daci.accumulator[11] ));
 sg13g2_nor2b_1 _1542_ (.A(_0266_),
    .B_N(_0268_),
    .Y(_0269_));
 sg13g2_o21ai_1 _1543_ (.B1(_0268_),
    .Y(_0270_),
    .A1(_0240_),
    .A2(_0265_));
 sg13g2_nand2_1 _1544_ (.Y(_0271_),
    .A(\stop.syn.daci.din[12] ),
    .B(net123));
 sg13g2_xnor2_1 _1545_ (.Y(_0272_),
    .A(\stop.syn.daci.din[12] ),
    .B(net123));
 sg13g2_nand2b_1 _1546_ (.Y(_0273_),
    .B(_0270_),
    .A_N(_0272_));
 sg13g2_nand2_1 _1547_ (.Y(_0274_),
    .A(net279),
    .B(_0273_));
 sg13g2_a21oi_1 _1548_ (.A1(_0269_),
    .A2(_0272_),
    .Y(_0171_),
    .B1(_0274_));
 sg13g2_nor2_1 _1549_ (.A(\stop.syn.daci.din[13] ),
    .B(net127),
    .Y(_0275_));
 sg13g2_xnor2_1 _1550_ (.Y(_0276_),
    .A(\stop.syn.daci.din[13] ),
    .B(net127));
 sg13g2_nand3_1 _1551_ (.B(_0273_),
    .C(_0276_),
    .A(_0271_),
    .Y(_0277_));
 sg13g2_a21oi_1 _1552_ (.A1(_0271_),
    .A2(_0273_),
    .Y(_0278_),
    .B1(_0276_));
 sg13g2_nand2_1 _1553_ (.Y(_0279_),
    .A(net280),
    .B(_0277_));
 sg13g2_nor2_1 _1554_ (.A(_0278_),
    .B(_0279_),
    .Y(_0172_));
 sg13g2_nor2_1 _1555_ (.A(_0272_),
    .B(_0276_),
    .Y(_0280_));
 sg13g2_nor2_1 _1556_ (.A(_0271_),
    .B(_0275_),
    .Y(_0281_));
 sg13g2_a221oi_1 _1557_ (.B2(_0280_),
    .C1(_0281_),
    .B1(_0270_),
    .A1(\stop.syn.daci.din[13] ),
    .Y(_0282_),
    .A2(net127));
 sg13g2_nand2_1 _1558_ (.Y(_0283_),
    .A(\stop.syn.daci.din[14] ),
    .B(net126));
 sg13g2_xnor2_1 _1559_ (.Y(_0284_),
    .A(\stop.syn.daci.din[14] ),
    .B(net126));
 sg13g2_o21ai_1 _1560_ (.B1(net279),
    .Y(_0285_),
    .A1(_0282_),
    .A2(_0284_));
 sg13g2_a21oi_1 _1561_ (.A1(_0282_),
    .A2(_0284_),
    .Y(_0173_),
    .B1(_0285_));
 sg13g2_xor2_1 _1562_ (.B(net121),
    .A(\stop.syn.daci.din[15] ),
    .X(_0286_));
 sg13g2_o21ai_1 _1563_ (.B1(_0283_),
    .Y(_0287_),
    .A1(_0282_),
    .A2(_0284_));
 sg13g2_o21ai_1 _1564_ (.B1(net279),
    .Y(_0288_),
    .A1(_0286_),
    .A2(_0287_));
 sg13g2_a21oi_1 _1565_ (.A1(_0286_),
    .A2(_0287_),
    .Y(_0174_),
    .B1(_0288_));
 sg13g2_a21oi_1 _1566_ (.A1(\stop.syn.daci.din[15] ),
    .A2(net121),
    .Y(_0289_),
    .B1(_0287_));
 sg13g2_o21ai_1 _1567_ (.B1(net279),
    .Y(_0290_),
    .A1(\stop.syn.daci.din[15] ),
    .A2(net121));
 sg13g2_nor2_1 _1568_ (.A(_0289_),
    .B(_0290_),
    .Y(_0175_));
 sg13g2_nor2_1 _1569_ (.A(\stop.ctrl.first_bit ),
    .B(net2),
    .Y(_0291_));
 sg13g2_mux2_1 _1570_ (.A0(\stop.adsr_ai[0] ),
    .A1(\stop.adsr_ai[1] ),
    .S(net337),
    .X(_0176_));
 sg13g2_nor2_1 _1571_ (.A(\stop.adsr_ai[1] ),
    .B(net336),
    .Y(_0292_));
 sg13g2_a21oi_1 _1572_ (.A1(_0304_),
    .A2(net336),
    .Y(_0177_),
    .B1(_0292_));
 sg13g2_nor2_1 _1573_ (.A(\stop.adsr_ai[2] ),
    .B(net335),
    .Y(_0293_));
 sg13g2_a21oi_1 _1574_ (.A1(_0305_),
    .A2(net335),
    .Y(_0178_),
    .B1(_0293_));
 sg13g2_nor2_1 _1575_ (.A(\stop.adsr_ai[3] ),
    .B(net334),
    .Y(_0294_));
 sg13g2_a21oi_1 _1576_ (.A1(_0306_),
    .A2(net334),
    .Y(_0179_),
    .B1(_0294_));
 sg13g2_nor2_1 _1577_ (.A(\stop.adsr_ai[4] ),
    .B(net333),
    .Y(_0295_));
 sg13g2_a21oi_1 _1578_ (.A1(_0307_),
    .A2(net333),
    .Y(_0180_),
    .B1(_0295_));
 sg13g2_nor2_1 _1579_ (.A(\stop.adsr_ai[5] ),
    .B(net333),
    .Y(_0296_));
 sg13g2_a21oi_1 _1580_ (.A1(_0308_),
    .A2(net333),
    .Y(_0181_),
    .B1(_0296_));
 sg13g2_nor2_1 _1581_ (.A(\stop.adsr_ai[6] ),
    .B(net334),
    .Y(_0297_));
 sg13g2_a21oi_1 _1582_ (.A1(_0309_),
    .A2(net333),
    .Y(_0182_),
    .B1(_0297_));
 sg13g2_nand2_1 _1583_ (.Y(_0298_),
    .A(\stop.adsr_di[0] ),
    .B(net335));
 sg13g2_o21ai_1 _1584_ (.B1(_0298_),
    .Y(_0183_),
    .A1(_0309_),
    .A2(net335));
 sg13g2_mux2_1 _1585_ (.A0(\stop.adsr_di[0] ),
    .A1(\stop.adsr_di[1] ),
    .S(net336),
    .X(_0184_));
 sg13g2_mux2_1 _1586_ (.A0(\stop.adsr_di[1] ),
    .A1(\stop.adsr_di[2] ),
    .S(net336),
    .X(_0185_));
 sg13g2_mux2_1 _1587_ (.A0(\stop.adsr_di[2] ),
    .A1(\stop.adsr_di[3] ),
    .S(net335),
    .X(_0186_));
 sg13g2_mux2_1 _1588_ (.A0(\stop.adsr_di[3] ),
    .A1(\stop.adsr_di[4] ),
    .S(net334),
    .X(_0187_));
 sg13g2_mux2_1 _1589_ (.A0(\stop.adsr_di[4] ),
    .A1(\stop.adsr_di[5] ),
    .S(net333),
    .X(_0188_));
 sg13g2_mux2_1 _1590_ (.A0(\stop.adsr_di[5] ),
    .A1(\stop.adsr_di[6] ),
    .S(net333),
    .X(_0189_));
 sg13g2_mux2_1 _1591_ (.A0(\stop.adsr_di[6] ),
    .A1(\stop.adsr_di[7] ),
    .S(net332),
    .X(_0190_));
 sg13g2_mux2_1 _1592_ (.A0(\stop.adsr_di[7] ),
    .A1(\stop.adsr_s[0] ),
    .S(net332),
    .X(_0191_));
 sg13g2_mux2_1 _1593_ (.A0(\stop.adsr_s[0] ),
    .A1(\stop.adsr_s[1] ),
    .S(net331),
    .X(_0192_));
 sg13g2_mux2_1 _1594_ (.A0(\stop.adsr_s[1] ),
    .A1(\stop.adsr_s[2] ),
    .S(net331),
    .X(_0193_));
 sg13g2_mux2_1 _1595_ (.A0(\stop.adsr_s[2] ),
    .A1(\stop.adsr_s[3] ),
    .S(net331),
    .X(_0194_));
 sg13g2_mux2_1 _1596_ (.A0(\stop.adsr_s[3] ),
    .A1(\stop.adsr_s[4] ),
    .S(net331),
    .X(_0195_));
 sg13g2_mux2_1 _1597_ (.A0(\stop.adsr_s[4] ),
    .A1(\stop.adsr_s[5] ),
    .S(net331),
    .X(_0196_));
 sg13g2_mux2_1 _1598_ (.A0(\stop.adsr_s[5] ),
    .A1(\stop.adsr_s[6] ),
    .S(net329),
    .X(_0197_));
 sg13g2_mux2_1 _1599_ (.A0(\stop.adsr_s[6] ),
    .A1(\stop.adsr_s[7] ),
    .S(net330),
    .X(_0198_));
 sg13g2_mux2_1 _1600_ (.A0(\stop.adsr_s[7] ),
    .A1(\stop.adsr_ri[0] ),
    .S(net337),
    .X(_0199_));
 sg13g2_mux2_1 _1601_ (.A0(\stop.adsr_ri[0] ),
    .A1(\stop.adsr_ri[1] ),
    .S(net335),
    .X(_0200_));
 sg13g2_mux2_1 _1602_ (.A0(\stop.adsr_ri[1] ),
    .A1(\stop.adsr_ri[2] ),
    .S(net336),
    .X(_0201_));
 sg13g2_mux2_1 _1603_ (.A0(\stop.adsr_ri[2] ),
    .A1(\stop.adsr_ri[3] ),
    .S(net335),
    .X(_0202_));
 sg13g2_mux2_1 _1604_ (.A0(\stop.adsr_ri[3] ),
    .A1(\stop.adsr_ri[4] ),
    .S(net335),
    .X(_0203_));
 sg13g2_mux2_1 _1605_ (.A0(\stop.adsr_ri[4] ),
    .A1(\stop.adsr_ri[5] ),
    .S(net334),
    .X(_0204_));
 sg13g2_mux2_1 _1606_ (.A0(\stop.adsr_ri[5] ),
    .A1(\stop.adsr_ri[6] ),
    .S(net333),
    .X(_0205_));
 sg13g2_mux2_1 _1607_ (.A0(\stop.adsr_ri[6] ),
    .A1(\stop.adsr_ri[7] ),
    .S(net331),
    .X(_0206_));
 sg13g2_mux2_1 _1608_ (.A0(\stop.adsr_ri[7] ),
    .A1(\stop.ctrl.cfg[32] ),
    .S(net329),
    .X(_0207_));
 sg13g2_mux2_1 _1609_ (.A0(\stop.ctrl.cfg[32] ),
    .A1(\stop.ctrl.cfg[33] ),
    .S(net329),
    .X(_0208_));
 sg13g2_mux2_1 _1610_ (.A0(\stop.ctrl.cfg[33] ),
    .A1(\stop.ctrl.cfg[34] ),
    .S(net329),
    .X(_0209_));
 sg13g2_mux2_1 _1611_ (.A0(\stop.ctrl.cfg[34] ),
    .A1(\stop.ctrl.cfg[35] ),
    .S(net329),
    .X(_0210_));
 sg13g2_mux2_1 _1612_ (.A0(\stop.ctrl.cfg[35] ),
    .A1(\stop.ctrl.cfg[36] ),
    .S(net329),
    .X(_0211_));
 sg13g2_mux2_1 _1613_ (.A0(\stop.ctrl.cfg[36] ),
    .A1(\stop.ctrl.cfg[37] ),
    .S(net329),
    .X(_0212_));
 sg13g2_mux2_1 _1614_ (.A0(\stop.ctrl.cfg[37] ),
    .A1(\stop.ctrl.cfg[38] ),
    .S(net329),
    .X(_0213_));
 sg13g2_mux2_1 _1615_ (.A0(\stop.ctrl.cfg[38] ),
    .A1(\stop.ctrl.cfg[39] ),
    .S(net330),
    .X(_0214_));
 sg13g2_mux2_1 _1616_ (.A0(\stop.ctrl.cfg[39] ),
    .A1(\stop.ctrl.cfg[40] ),
    .S(net330),
    .X(_0215_));
 sg13g2_mux2_1 _1617_ (.A0(\stop.ctrl.cfg[40] ),
    .A1(\stop.ctrl.cfg[41] ),
    .S(net330),
    .X(_0216_));
 sg13g2_mux2_1 _1618_ (.A0(\stop.ctrl.cfg[41] ),
    .A1(\stop.ctrl.cfg[42] ),
    .S(net338),
    .X(_0217_));
 sg13g2_mux2_1 _1619_ (.A0(\stop.ctrl.cfg[42] ),
    .A1(\stop.ctrl.cfg[43] ),
    .S(net338),
    .X(_0218_));
 sg13g2_mux2_1 _1620_ (.A0(\stop.ctrl.cfg[43] ),
    .A1(\stop.ctrl.cfg[44] ),
    .S(net332),
    .X(_0219_));
 sg13g2_mux2_1 _1621_ (.A0(\stop.ctrl.cfg[44] ),
    .A1(\stop.ctrl.cfg[45] ),
    .S(net332),
    .X(_0220_));
 sg13g2_mux2_1 _1622_ (.A0(\stop.ctrl.cfg[45] ),
    .A1(\stop.ctrl.cfg[46] ),
    .S(net338),
    .X(_0221_));
 sg13g2_mux2_1 _1623_ (.A0(\stop.ctrl.cfg[46] ),
    .A1(\stop.ctrl.cfg[47] ),
    .S(net332),
    .X(_0222_));
 sg13g2_mux2_1 _1624_ (.A0(\stop.ctrl.cfg[47] ),
    .A1(\stop.ctrl.cfg[48] ),
    .S(net332),
    .X(_0223_));
 sg13g2_mux2_1 _1625_ (.A0(\stop.ctrl.cfg[48] ),
    .A1(\stop.ctrl.cfg[49] ),
    .S(net332),
    .X(_0224_));
 sg13g2_mux2_1 _1626_ (.A0(\stop.ctrl.cfg[49] ),
    .A1(\stop.ctrl.cfg[50] ),
    .S(net340),
    .X(_0225_));
 sg13g2_mux2_1 _1627_ (.A0(\stop.ctrl.cfg[50] ),
    .A1(\stop.ctrl.cfg[51] ),
    .S(net340),
    .X(_0226_));
 sg13g2_mux2_1 _1628_ (.A0(\stop.ctrl.cfg[51] ),
    .A1(\stop.ctrl.cfg[52] ),
    .S(net340),
    .X(_0227_));
 sg13g2_mux2_1 _1629_ (.A0(\stop.ctrl.cfg[52] ),
    .A1(\stop.ctrl.cfg[53] ),
    .S(net339),
    .X(_0228_));
 sg13g2_mux2_1 _1630_ (.A0(\stop.ctrl.cfg[53] ),
    .A1(\stop.ctrl.cfg[54] ),
    .S(net339),
    .X(_0229_));
 sg13g2_mux2_1 _1631_ (.A0(\stop.ctrl.cfg[54] ),
    .A1(\stop.ctrl.cfg[55] ),
    .S(net339),
    .X(_0230_));
 sg13g2_mux2_1 _1632_ (.A0(\stop.ctrl.cfg[55] ),
    .A1(\stop.ctrl.cfg[56] ),
    .S(net339),
    .X(_0231_));
 sg13g2_mux2_1 _1633_ (.A0(\stop.ctrl.cfg[56] ),
    .A1(\stop.ctrl.cfg[57] ),
    .S(net339),
    .X(_0232_));
 sg13g2_mux2_1 _1634_ (.A0(\stop.ctrl.cfg[57] ),
    .A1(\stop.ctrl.cfg[58] ),
    .S(net339),
    .X(_0233_));
 sg13g2_mux2_1 _1635_ (.A0(\stop.ctrl.cfg[58] ),
    .A1(\stop.ctrl.cfg[59] ),
    .S(net339),
    .X(_0234_));
 sg13g2_mux2_1 _1636_ (.A0(\stop.ctrl.cfg[59] ),
    .A1(net3),
    .S(net339),
    .X(_0235_));
 sg13g2_inv_1 _1637_ (.Y(_0132_),
    .A(net291));
 sg13g2_inv_1 _1638_ (.Y(_0131_),
    .A(net291));
 sg13g2_inv_1 _1639_ (.Y(_0130_),
    .A(net291));
 sg13g2_inv_1 _1640_ (.Y(_0129_),
    .A(net291));
 sg13g2_inv_1 _1641_ (.Y(_0128_),
    .A(net291));
 sg13g2_inv_1 _1642_ (.Y(_0127_),
    .A(net291));
 sg13g2_inv_1 _1643_ (.Y(_0126_),
    .A(net287));
 sg13g2_inv_1 _1644_ (.Y(_0125_),
    .A(net287));
 sg13g2_inv_1 _1645_ (.Y(_0124_),
    .A(net294));
 sg13g2_inv_1 _1646_ (.Y(_0123_),
    .A(net294));
 sg13g2_inv_1 _1647_ (.Y(_0122_),
    .A(net292));
 sg13g2_inv_1 _1648_ (.Y(_0121_),
    .A(net292));
 sg13g2_inv_1 _1649_ (.Y(_0120_),
    .A(net293));
 sg13g2_inv_1 _1650_ (.Y(_0119_),
    .A(net293));
 sg13g2_inv_1 _1651_ (.Y(_0118_),
    .A(net292));
 sg13g2_inv_1 _1652_ (.Y(_0117_),
    .A(net290));
 sg13g2_inv_1 _1653_ (.Y(_0116_),
    .A(net290));
 sg13g2_inv_1 _1654_ (.Y(_0115_),
    .A(net290));
 sg13g2_inv_1 _1655_ (.Y(_0114_),
    .A(net290));
 sg13g2_inv_1 _1656_ (.Y(_0113_),
    .A(net290));
 sg13g2_inv_1 _1657_ (.Y(_0112_),
    .A(net289));
 sg13g2_inv_1 _1658_ (.Y(_0111_),
    .A(net289));
 sg13g2_inv_1 _1659_ (.Y(_0110_),
    .A(net289));
 sg13g2_inv_1 _1660_ (.Y(_0109_),
    .A(net288));
 sg13g2_inv_1 _1661_ (.Y(_0108_),
    .A(net288));
 sg13g2_inv_1 _1662_ (.Y(_0107_),
    .A(net294));
 sg13g2_inv_1 _1663_ (.Y(_0106_),
    .A(net294));
 sg13g2_inv_1 _1664_ (.Y(_0105_),
    .A(net293));
 sg13g2_inv_1 _1665_ (.Y(_0104_),
    .A(net293));
 sg13g2_inv_1 _1666_ (.Y(_0103_),
    .A(net293));
 sg13g2_inv_1 _1667_ (.Y(_0102_),
    .A(net292));
 sg13g2_inv_1 _1668_ (.Y(_0101_),
    .A(net289));
 sg13g2_inv_1 _1669_ (.Y(_0100_),
    .A(net290));
 sg13g2_inv_1 _1670_ (.Y(_0099_),
    .A(net290));
 sg13g2_inv_1 _1671_ (.Y(_0098_),
    .A(net290));
 sg13g2_inv_1 _1672_ (.Y(_0097_),
    .A(net289));
 sg13g2_inv_1 _1673_ (.Y(_0096_),
    .A(net289));
 sg13g2_inv_1 _1674_ (.Y(_0095_),
    .A(net289));
 sg13g2_inv_1 _1675_ (.Y(_0094_),
    .A(net289));
 sg13g2_inv_1 _1676_ (.Y(_0093_),
    .A(net288));
 sg13g2_inv_1 _1677_ (.Y(_0092_),
    .A(net288));
 sg13g2_inv_1 _1678_ (.Y(_0091_),
    .A(net288));
 sg13g2_inv_1 _1679_ (.Y(_0090_),
    .A(net294));
 sg13g2_inv_1 _1680_ (.Y(_0089_),
    .A(net294));
 sg13g2_inv_1 _1681_ (.Y(_0088_),
    .A(net294));
 sg13g2_inv_1 _1682_ (.Y(_0087_),
    .A(net292));
 sg13g2_inv_1 _1683_ (.Y(_0086_),
    .A(net292));
 sg13g2_inv_1 _1684_ (.Y(_0085_),
    .A(net2));
 sg13g2_dfrbp_1 _1685_ (.CLK(net285),
    .RESET_B(net29),
    .D(_0000_),
    .Q_N(_0856_),
    .Q(\stop.syn.adsri.state[0] ));
 sg13g2_dfrbp_1 _1686_ (.CLK(net285),
    .RESET_B(net30),
    .D(_0001_),
    .Q_N(_0857_),
    .Q(\stop.syn.adsri.state[1] ));
 sg13g2_dfrbp_1 _1687_ (.CLK(\stop.syn.adsri.clk ),
    .RESET_B(net31),
    .D(_0002_),
    .Q_N(_0858_),
    .Q(\stop.syn.adsri.state[2] ));
 sg13g2_dfrbp_1 _1688_ (.CLK(net285),
    .RESET_B(net46),
    .D(_0003_),
    .Q_N(_0859_),
    .Q(\stop.syn.adsri.state[3] ));
 sg13g2_dfrbp_1 _1689_ (.CLK(net285),
    .RESET_B(net28),
    .D(_0004_),
    .Q_N(_0855_),
    .Q(\stop.syn.adsri.state[4] ));
 sg13g2_dfrbp_1 _1690_ (.CLK(net320),
    .RESET_B(net85),
    .D(_0134_),
    .Q_N(_0854_),
    .Q(\stop.syn.smul8.b_latched[7] ));
 sg13g2_dfrbp_1 _1691_ (.CLK(net314),
    .RESET_B(net83),
    .D(_0005_),
    .Q_N(_0853_),
    .Q(\stop.syn.filt.m1.b_bit ));
 sg13g2_dfrbp_1 _1692_ (.CLK(net315),
    .RESET_B(net82),
    .D(_0006_),
    .Q_N(_0852_),
    .Q(\stop.syn.filt.m1.b_latched[1] ));
 sg13g2_dfrbp_1 _1693_ (.CLK(net315),
    .RESET_B(net81),
    .D(_0007_),
    .Q_N(_0851_),
    .Q(\stop.syn.filt.m1.b_latched[2] ));
 sg13g2_dfrbp_1 _1694_ (.CLK(net315),
    .RESET_B(net80),
    .D(_0008_),
    .Q_N(_0850_),
    .Q(\stop.syn.filt.m1.b_latched[3] ));
 sg13g2_dfrbp_1 _1695_ (.CLK(net315),
    .RESET_B(net79),
    .D(_0009_),
    .Q_N(_0849_),
    .Q(\stop.syn.filt.m1.b_latched[4] ));
 sg13g2_dfrbp_1 _1696_ (.CLK(net314),
    .RESET_B(net78),
    .D(_0010_),
    .Q_N(_0848_),
    .Q(\stop.syn.filt.m1.b_latched[5] ));
 sg13g2_dfrbp_1 _1697_ (.CLK(net314),
    .RESET_B(net77),
    .D(_0011_),
    .Q_N(_0847_),
    .Q(\stop.syn.filt.m1.b_latched[6] ));
 sg13g2_dfrbp_1 _1698_ (.CLK(net326),
    .RESET_B(net76),
    .D(_0012_),
    .Q_N(_0846_),
    .Q(\stop.syn.filt.m2.b_bit ));
 sg13g2_dfrbp_1 _1699_ (.CLK(net325),
    .RESET_B(net75),
    .D(_0013_),
    .Q_N(_0845_),
    .Q(\stop.syn.filt.m2.b_latched[1] ));
 sg13g2_dfrbp_1 _1700_ (.CLK(net325),
    .RESET_B(net74),
    .D(_0014_),
    .Q_N(_0844_),
    .Q(\stop.syn.filt.m2.b_latched[2] ));
 sg13g2_dfrbp_1 _1701_ (.CLK(net325),
    .RESET_B(net73),
    .D(_0015_),
    .Q_N(_0843_),
    .Q(\stop.syn.filt.m2.b_latched[3] ));
 sg13g2_dfrbp_1 _1702_ (.CLK(net325),
    .RESET_B(net72),
    .D(_0016_),
    .Q_N(_0842_),
    .Q(\stop.syn.filt.m2.b_latched[4] ));
 sg13g2_dfrbp_1 _1703_ (.CLK(net326),
    .RESET_B(net71),
    .D(_0017_),
    .Q_N(_0841_),
    .Q(\stop.syn.filt.m2.b_latched[5] ));
 sg13g2_dfrbp_1 _1704_ (.CLK(net325),
    .RESET_B(net70),
    .D(_0018_),
    .Q_N(_0840_),
    .Q(\stop.syn.filt.m2.b_latched[6] ));
 sg13g2_dfrbp_1 _1705_ (.CLK(net314),
    .RESET_B(net69),
    .D(_0019_),
    .Q_N(_0839_),
    .Q(\stop.syn.smul8.b_bit ));
 sg13g2_dfrbp_1 _1706_ (.CLK(net322),
    .RESET_B(net45),
    .D(_0020_),
    .Q_N(_0838_),
    .Q(\stop.syn.smul8.b_latched[1] ));
 sg13g2_dfrbp_1 _1707_ (.CLK(net322),
    .RESET_B(net44),
    .D(_0021_),
    .Q_N(_0837_),
    .Q(\stop.syn.smul8.b_latched[2] ));
 sg13g2_dfrbp_1 _1708_ (.CLK(net322),
    .RESET_B(net43),
    .D(_0022_),
    .Q_N(_0836_),
    .Q(\stop.syn.smul8.b_latched[3] ));
 sg13g2_dfrbp_1 _1709_ (.CLK(net320),
    .RESET_B(net42),
    .D(_0023_),
    .Q_N(_0835_),
    .Q(\stop.syn.smul8.b_latched[4] ));
 sg13g2_dfrbp_1 _1710_ (.CLK(net320),
    .RESET_B(net41),
    .D(_0024_),
    .Q_N(_0834_),
    .Q(\stop.syn.smul8.b_latched[5] ));
 sg13g2_dfrbp_1 _1711_ (.CLK(net320),
    .RESET_B(net40),
    .D(_0025_),
    .Q_N(_0833_),
    .Q(\stop.syn.smul8.b_latched[6] ));
 sg13g2_dfrbp_1 _1712_ (.CLK(net351),
    .RESET_B(_0083_),
    .D(_0082_),
    .Q_N(\stop.ctrl.first_bit_reg ),
    .Q(_0080_));
 sg13g2_dfrbp_1 _1713_ (.CLK(net352),
    .RESET_B(net362),
    .D(_0135_),
    .Q_N(_0832_),
    .Q(\stop.ctrl.trig ));
 sg13g2_dfrbp_1 _1714_ (.CLK(net351),
    .RESET_B(_0085_),
    .D(net116),
    .Q_N(\stop.ctrl.first_bit ),
    .Q(_0081_));
 sg13g2_dfrbp_1 _1715_ (.CLK(net303),
    .RESET_B(net47),
    .D(\stop.syn.adsr_data[0] ),
    .Q_N(_0860_),
    .Q(\stop.syn.adsr_data_reg[0] ));
 sg13g2_dfrbp_1 _1716_ (.CLK(net303),
    .RESET_B(net48),
    .D(\stop.syn.adsr_data[1] ),
    .Q_N(_0861_),
    .Q(\stop.syn.adsr_data_reg[1] ));
 sg13g2_dfrbp_1 _1717_ (.CLK(net303),
    .RESET_B(net49),
    .D(\stop.syn.adsr_data[2] ),
    .Q_N(_0862_),
    .Q(\stop.syn.adsr_data_reg[2] ));
 sg13g2_dfrbp_1 _1718_ (.CLK(net303),
    .RESET_B(net50),
    .D(\stop.syn.adsr_data[3] ),
    .Q_N(_0863_),
    .Q(\stop.syn.adsr_data_reg[3] ));
 sg13g2_dfrbp_1 _1719_ (.CLK(net303),
    .RESET_B(net51),
    .D(\stop.syn.adsr_data[4] ),
    .Q_N(_0864_),
    .Q(\stop.syn.adsr_data_reg[4] ));
 sg13g2_dfrbp_1 _1720_ (.CLK(net302),
    .RESET_B(net52),
    .D(\stop.syn.adsr_data[5] ),
    .Q_N(_0865_),
    .Q(\stop.syn.adsr_data_reg[5] ));
 sg13g2_dfrbp_1 _1721_ (.CLK(net301),
    .RESET_B(net53),
    .D(\stop.syn.adsr_data[6] ),
    .Q_N(_0866_),
    .Q(\stop.syn.adsr_data_reg[6] ));
 sg13g2_dfrbp_1 _1722_ (.CLK(net299),
    .RESET_B(net54),
    .D(\stop.syn.adsr_data[7] ),
    .Q_N(_0867_),
    .Q(\stop.syn.adsr_data_reg[7] ));
 sg13g2_dfrbp_1 _1723_ (.CLK(net299),
    .RESET_B(net55),
    .D(\stop.syn.adsr_data[8] ),
    .Q_N(_0868_),
    .Q(\stop.syn.adsr_data_reg[8] ));
 sg13g2_dfrbp_1 _1724_ (.CLK(net299),
    .RESET_B(net56),
    .D(\stop.syn.adsr_data[9] ),
    .Q_N(_0869_),
    .Q(\stop.syn.adsr_data_reg[9] ));
 sg13g2_dfrbp_1 _1725_ (.CLK(net299),
    .RESET_B(net57),
    .D(\stop.syn.adsr_data[10] ),
    .Q_N(_0870_),
    .Q(\stop.syn.adsr_data_reg[10] ));
 sg13g2_dfrbp_1 _1726_ (.CLK(net300),
    .RESET_B(net58),
    .D(\stop.syn.adsr_data[11] ),
    .Q_N(_0871_),
    .Q(\stop.syn.adsr_data_reg[11] ));
 sg13g2_dfrbp_1 _1727_ (.CLK(net299),
    .RESET_B(net59),
    .D(\stop.syn.adsr_data[12] ),
    .Q_N(_0872_),
    .Q(\stop.syn.adsr_data_reg[12] ));
 sg13g2_dfrbp_1 _1728_ (.CLK(net299),
    .RESET_B(net60),
    .D(\stop.syn.adsr_data[13] ),
    .Q_N(_0873_),
    .Q(\stop.syn.adsr_data_reg[13] ));
 sg13g2_dfrbp_1 _1729_ (.CLK(net299),
    .RESET_B(net61),
    .D(\stop.syn.adsr_data[14] ),
    .Q_N(_0874_),
    .Q(\stop.syn.adsr_data_reg[14] ));
 sg13g2_dfrbp_1 _1730_ (.CLK(net299),
    .RESET_B(net62),
    .D(\stop.syn.adsr_data[15] ),
    .Q_N(_0875_),
    .Q(\stop.syn.adsr_data_reg[15] ));
 sg13g2_dfrbp_1 _1731_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net63),
    .D(net327),
    .Q_N(_0876_),
    .Q(\stop.syn.rstn_fst_reg1 ));
 sg13g2_dfrbp_1 _1732_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net64),
    .D(net118),
    .Q_N(_0877_),
    .Q(\stop.syn.rstn_fst_reg2 ));
 sg13g2_dfrbp_1 _1733_ (.CLK(net285),
    .RESET_B(net65),
    .D(\stop.merge_trig ),
    .Q_N(_0878_),
    .Q(\stop.syn.trig_reg1 ));
 sg13g2_dfrbp_1 _1734_ (.CLK(net285),
    .RESET_B(net66),
    .D(\stop.syn.trig_reg1 ),
    .Q_N(_0879_),
    .Q(\stop.syn.adsri.trig ));
 sg13g2_dfrbp_1 _1735_ (.CLK(net286),
    .RESET_B(net67),
    .D(net327),
    .Q_N(_0880_),
    .Q(\stop.syn.rstn_reg1 ));
 sg13g2_dfrbp_1 _1736_ (.CLK(net286),
    .RESET_B(net68),
    .D(\stop.syn.rstn_reg1 ),
    .Q_N(_0047_),
    .Q(\stop.syn.adsri.rstn ));
 sg13g2_dfrbp_1 _1737_ (.CLK(\stop.syn.clki.gen[14].inst.q ),
    .RESET_B(net342),
    .D(_0033_),
    .Q_N(_0033_),
    .Q(\stop.syn.adsri.clk ));
 sg13g2_dfrbp_1 _1738_ (.CLK(\stop.syn.clki.gen[13].inst.q ),
    .RESET_B(net342),
    .D(_0032_),
    .Q_N(_0032_),
    .Q(\stop.syn.clki.gen[14].inst.q ));
 sg13g2_dfrbp_1 _1739_ (.CLK(\stop.syn.clki.gen[12].inst.q ),
    .RESET_B(net342),
    .D(_0031_),
    .Q_N(_0031_),
    .Q(\stop.syn.clki.gen[13].inst.q ));
 sg13g2_dfrbp_1 _1740_ (.CLK(\stop.syn.clki.gen[11].inst.q ),
    .RESET_B(net341),
    .D(_0030_),
    .Q_N(_0030_),
    .Q(\stop.syn.clki.gen[12].inst.q ));
 sg13g2_dfrbp_1 _1741_ (.CLK(\stop.syn.clki.gen[10].inst.q ),
    .RESET_B(net341),
    .D(_0029_),
    .Q_N(_0029_),
    .Q(\stop.syn.clki.gen[11].inst.q ));
 sg13g2_dfrbp_1 _1742_ (.CLK(\stop.syn.clki.gen[10].inst.clk ),
    .RESET_B(net341),
    .D(_0028_),
    .Q_N(_0028_),
    .Q(\stop.syn.clki.gen[10].inst.q ));
 sg13g2_dfrbp_1 _1743_ (.CLK(net298),
    .RESET_B(net341),
    .D(_0041_),
    .Q_N(_0041_),
    .Q(\stop.syn.clki.gen[10].inst.clk ));
 sg13g2_dfrbp_1 _1744_ (.CLK(\stop.syn.clk_sample_x2 ),
    .RESET_B(\stop.syn.clki.arstn ),
    .D(_0040_),
    .Q_N(_0040_),
    .Q(\stop.syn.clk_sample ));
 sg13g2_dfrbp_1 _1745_ (.CLK(\stop.syn.clki.gen[6].inst.q ),
    .RESET_B(net342),
    .D(_0026_),
    .Q_N(_0026_),
    .Q(\stop.syn.clk_sample_x2 ));
 sg13g2_dfrbp_1 _1746_ (.CLK(\stop.syn.clki.gen[5].inst.q ),
    .RESET_B(net342),
    .D(_0039_),
    .Q_N(_0039_),
    .Q(\stop.syn.clki.gen[6].inst.q ));
 sg13g2_dfrbp_1 _1747_ (.CLK(\stop.syn.clk_mult ),
    .RESET_B(net342),
    .D(_0038_),
    .Q_N(_0038_),
    .Q(\stop.syn.clki.gen[5].inst.q ));
 sg13g2_dfrbp_1 _1748_ (.CLK(\stop.syn.clki.gen[3].inst.q ),
    .RESET_B(net341),
    .D(net314),
    .Q_N(_0037_),
    .Q(\stop.syn.clk_mult ));
 sg13g2_dfrbp_1 _1749_ (.CLK(\stop.syn.clki.gen[2].inst.q ),
    .RESET_B(net341),
    .D(_0036_),
    .Q_N(_0036_),
    .Q(\stop.syn.clki.gen[3].inst.q ));
 sg13g2_dfrbp_1 _1750_ (.CLK(\stop.syn.clki.gen[1].inst.q ),
    .RESET_B(net342),
    .D(_0035_),
    .Q_N(_0035_),
    .Q(\stop.syn.clki.gen[2].inst.q ));
 sg13g2_dfrbp_1 _1751_ (.CLK(\stop.syn.clki.gen[0].inst.q ),
    .RESET_B(net341),
    .D(_0034_),
    .Q_N(_0034_),
    .Q(\stop.syn.clki.gen[1].inst.q ));
 sg13g2_dfrbp_1 _1752_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net341),
    .D(net117),
    .Q_N(_0027_),
    .Q(\stop.syn.clki.gen[0].inst.q ));
 sg13g2_dfrbp_1 _1753_ (.CLK(net285),
    .RESET_B(net37),
    .D(_0136_),
    .Q_N(_0831_),
    .Q(\stop.syn.adsri.envelope[0] ));
 sg13g2_dfrbp_1 _1754_ (.CLK(\stop.syn.adsri.clk ),
    .RESET_B(net36),
    .D(_0137_),
    .Q_N(_0830_),
    .Q(\stop.syn.adsri.envelope[1] ));
 sg13g2_dfrbp_1 _1755_ (.CLK(net285),
    .RESET_B(net35),
    .D(_0138_),
    .Q_N(_0829_),
    .Q(\stop.syn.adsri.envelope[2] ));
 sg13g2_dfrbp_1 _1756_ (.CLK(net286),
    .RESET_B(net34),
    .D(_0139_),
    .Q_N(_0828_),
    .Q(\stop.syn.adsri.envelope[3] ));
 sg13g2_dfrbp_1 _1757_ (.CLK(net286),
    .RESET_B(net33),
    .D(_0140_),
    .Q_N(_0827_),
    .Q(\stop.syn.adsri.envelope[4] ));
 sg13g2_dfrbp_1 _1758_ (.CLK(net286),
    .RESET_B(net32),
    .D(_0141_),
    .Q_N(_0826_),
    .Q(\stop.syn.adsri.envelope[5] ));
 sg13g2_dfrbp_1 _1759_ (.CLK(net286),
    .RESET_B(net27),
    .D(_0142_),
    .Q_N(_0825_),
    .Q(\stop.syn.adsri.envelope[6] ));
 sg13g2_dfrbp_1 _1760_ (.CLK(net286),
    .RESET_B(net115),
    .D(_0143_),
    .Q_N(_0824_),
    .Q(\stop.syn.adsri.envelope[7] ));
 sg13g2_dfrbp_1 _1761_ (.CLK(net298),
    .RESET_B(net114),
    .D(_0144_),
    .Q_N(_0079_),
    .Q(\stop.syn.osci.counter[0] ));
 sg13g2_dfrbp_1 _1762_ (.CLK(net297),
    .RESET_B(net113),
    .D(_0145_),
    .Q_N(_0823_),
    .Q(\stop.syn.osci.counter[1] ));
 sg13g2_dfrbp_1 _1763_ (.CLK(net297),
    .RESET_B(net112),
    .D(_0146_),
    .Q_N(_0822_),
    .Q(\stop.syn.osci.counter[2] ));
 sg13g2_dfrbp_1 _1764_ (.CLK(net297),
    .RESET_B(net111),
    .D(_0147_),
    .Q_N(_0821_),
    .Q(\stop.syn.osci.counter[3] ));
 sg13g2_dfrbp_1 _1765_ (.CLK(net297),
    .RESET_B(net110),
    .D(_0148_),
    .Q_N(_0820_),
    .Q(\stop.syn.osci.counter[4] ));
 sg13g2_dfrbp_1 _1766_ (.CLK(net297),
    .RESET_B(net109),
    .D(_0149_),
    .Q_N(_0819_),
    .Q(\stop.syn.osci.counter[5] ));
 sg13g2_dfrbp_1 _1767_ (.CLK(net298),
    .RESET_B(net108),
    .D(_0150_),
    .Q_N(_0818_),
    .Q(\stop.syn.osci.counter[6] ));
 sg13g2_dfrbp_1 _1768_ (.CLK(net297),
    .RESET_B(net107),
    .D(_0151_),
    .Q_N(_0817_),
    .Q(\stop.syn.osci.counter[7] ));
 sg13g2_dfrbp_1 _1769_ (.CLK(net297),
    .RESET_B(net106),
    .D(_0152_),
    .Q_N(_0816_),
    .Q(\stop.syn.osci.counter[8] ));
 sg13g2_dfrbp_1 _1770_ (.CLK(net297),
    .RESET_B(net105),
    .D(_0153_),
    .Q_N(_0815_),
    .Q(\stop.syn.osci.counter[9] ));
 sg13g2_dfrbp_1 _1771_ (.CLK(net298),
    .RESET_B(net104),
    .D(_0154_),
    .Q_N(_0814_),
    .Q(\stop.syn.osci.counter[10] ));
 sg13g2_dfrbp_1 _1772_ (.CLK(net298),
    .RESET_B(net103),
    .D(_0155_),
    .Q_N(_0813_),
    .Q(\stop.syn.osci.counter[11] ));
 sg13g2_dfrbp_1 _1773_ (.CLK(net325),
    .RESET_B(net102),
    .D(_0156_),
    .Q_N(_0812_),
    .Q(\stop.syn.filt.m2.b_latched[7] ));
 sg13g2_dfrbp_1 _1774_ (.CLK(net298),
    .RESET_B(net101),
    .D(_0157_),
    .Q_N(_0042_),
    .Q(\stop.syn.osci.data_buf ));
 sg13g2_dfrbp_1 _1775_ (.CLK(net322),
    .RESET_B(_0086_),
    .D(\stop.syn.adsr_data[1] ),
    .Q_N(_0811_),
    .Q(\stop.syn.adsr_data[0] ));
 sg13g2_dfrbp_1 _1776_ (.CLK(net320),
    .RESET_B(_0087_),
    .D(\stop.syn.adsr_data[2] ),
    .Q_N(_0810_),
    .Q(\stop.syn.adsr_data[1] ));
 sg13g2_dfrbp_1 _1777_ (.CLK(net320),
    .RESET_B(_0088_),
    .D(\stop.syn.adsr_data[3] ),
    .Q_N(_0809_),
    .Q(\stop.syn.adsr_data[2] ));
 sg13g2_dfrbp_1 _1778_ (.CLK(net320),
    .RESET_B(_0089_),
    .D(\stop.syn.adsr_data[4] ),
    .Q_N(_0808_),
    .Q(\stop.syn.adsr_data[3] ));
 sg13g2_dfrbp_1 _1779_ (.CLK(net321),
    .RESET_B(_0090_),
    .D(\stop.syn.adsr_data[5] ),
    .Q_N(_0807_),
    .Q(\stop.syn.adsr_data[4] ));
 sg13g2_dfrbp_1 _1780_ (.CLK(net315),
    .RESET_B(_0091_),
    .D(\stop.syn.adsr_data[6] ),
    .Q_N(_0806_),
    .Q(\stop.syn.adsr_data[5] ));
 sg13g2_dfrbp_1 _1781_ (.CLK(net314),
    .RESET_B(_0092_),
    .D(\stop.syn.adsr_data[7] ),
    .Q_N(_0805_),
    .Q(\stop.syn.adsr_data[6] ));
 sg13g2_dfrbp_1 _1782_ (.CLK(net314),
    .RESET_B(_0093_),
    .D(_0071_),
    .Q_N(_0804_),
    .Q(\stop.syn.adsr_data[7] ));
 sg13g2_dfrbp_1 _1783_ (.CLK(net317),
    .RESET_B(_0094_),
    .D(_0072_),
    .Q_N(_0803_),
    .Q(\stop.syn.adsr_data[8] ));
 sg13g2_dfrbp_1 _1784_ (.CLK(net317),
    .RESET_B(_0095_),
    .D(_0073_),
    .Q_N(_0802_),
    .Q(\stop.syn.adsr_data[9] ));
 sg13g2_dfrbp_1 _1785_ (.CLK(net317),
    .RESET_B(_0096_),
    .D(_0074_),
    .Q_N(_0801_),
    .Q(\stop.syn.adsr_data[10] ));
 sg13g2_dfrbp_1 _1786_ (.CLK(net317),
    .RESET_B(_0097_),
    .D(_0075_),
    .Q_N(_0052_),
    .Q(\stop.syn.adsr_data[11] ));
 sg13g2_dfrbp_1 _1787_ (.CLK(net316),
    .RESET_B(_0098_),
    .D(_0076_),
    .Q_N(_0800_),
    .Q(\stop.syn.adsr_data[12] ));
 sg13g2_dfrbp_1 _1788_ (.CLK(net316),
    .RESET_B(_0099_),
    .D(_0077_),
    .Q_N(_0053_),
    .Q(\stop.syn.adsr_data[13] ));
 sg13g2_dfrbp_1 _1789_ (.CLK(net316),
    .RESET_B(_0100_),
    .D(_0078_),
    .Q_N(_0799_),
    .Q(\stop.syn.adsr_data[14] ));
 sg13g2_dfrbp_1 _1790_ (.CLK(net316),
    .RESET_B(_0101_),
    .D(_0070_),
    .Q_N(_0798_),
    .Q(\stop.syn.adsr_data[15] ));
 sg13g2_dfrbp_1 _1791_ (.CLK(net322),
    .RESET_B(_0102_),
    .D(\stop.syn.filt.m2.sum[1] ),
    .Q_N(_0797_),
    .Q(\stop.syn.filt.m2.sum_in2[0] ));
 sg13g2_dfrbp_1 _1792_ (.CLK(net323),
    .RESET_B(_0103_),
    .D(\stop.syn.filt.m2.sum[2] ),
    .Q_N(_0796_),
    .Q(\stop.syn.filt.m2.sum_in2[1] ));
 sg13g2_dfrbp_1 _1793_ (.CLK(net323),
    .RESET_B(_0104_),
    .D(\stop.syn.filt.m2.sum[3] ),
    .Q_N(_0795_),
    .Q(\stop.syn.filt.m2.sum_in2[2] ));
 sg13g2_dfrbp_1 _1794_ (.CLK(net321),
    .RESET_B(_0105_),
    .D(\stop.syn.filt.m2.sum[4] ),
    .Q_N(_0043_),
    .Q(\stop.syn.filt.m2.sum_in2[3] ));
 sg13g2_dfrbp_1 _1795_ (.CLK(net321),
    .RESET_B(_0106_),
    .D(\stop.syn.filt.m2.sum[5] ),
    .Q_N(_0794_),
    .Q(\stop.syn.filt.m2.sum_in2[4] ));
 sg13g2_dfrbp_1 _1796_ (.CLK(net321),
    .RESET_B(_0107_),
    .D(\stop.syn.filt.m2.sum[6] ),
    .Q_N(_0044_),
    .Q(\stop.syn.filt.m2.sum_in2[5] ));
 sg13g2_dfrbp_1 _1797_ (.CLK(net315),
    .RESET_B(_0108_),
    .D(\stop.syn.filt.m2.sum[7] ),
    .Q_N(_0793_),
    .Q(\stop.syn.filt.m2.sum_in2[6] ));
 sg13g2_dfrbp_1 _1798_ (.CLK(net317),
    .RESET_B(_0109_),
    .D(\stop.syn.filt.m2.sum[8] ),
    .Q_N(_0792_),
    .Q(\stop.syn.filt.m2.sum_in2[7] ));
 sg13g2_dfrbp_1 _1799_ (.CLK(net317),
    .RESET_B(_0110_),
    .D(\stop.syn.filt.m2.sum[9] ),
    .Q_N(_0791_),
    .Q(\stop.syn.filt.m2.sum_in2[8] ));
 sg13g2_dfrbp_1 _1800_ (.CLK(net317),
    .RESET_B(_0111_),
    .D(\stop.syn.filt.m2.sum[10] ),
    .Q_N(_0045_),
    .Q(\stop.syn.filt.m2.sum_in2[9] ));
 sg13g2_dfrbp_1 _1801_ (.CLK(net317),
    .RESET_B(_0112_),
    .D(\stop.syn.filt.m2.sum[11] ),
    .Q_N(_0790_),
    .Q(\stop.syn.filt.m2.sum_in2[10] ));
 sg13g2_dfrbp_1 _1802_ (.CLK(net318),
    .RESET_B(_0113_),
    .D(\stop.syn.filt.m2.sum[12] ),
    .Q_N(_0789_),
    .Q(\stop.syn.filt.m2.sum_in2[11] ));
 sg13g2_dfrbp_1 _1803_ (.CLK(net316),
    .RESET_B(_0114_),
    .D(\stop.syn.filt.m2.sum[13] ),
    .Q_N(_0788_),
    .Q(\stop.syn.filt.m2.sum_in2[12] ));
 sg13g2_dfrbp_1 _1804_ (.CLK(net316),
    .RESET_B(_0115_),
    .D(\stop.syn.filt.m2.sum[14] ),
    .Q_N(_0046_),
    .Q(\stop.syn.filt.m2.sum_in2[13] ));
 sg13g2_dfrbp_1 _1805_ (.CLK(net316),
    .RESET_B(_0116_),
    .D(\stop.syn.filt.m2.sum[15] ),
    .Q_N(_0787_),
    .Q(\stop.syn.filt.m2.sum_in2[14] ));
 sg13g2_dfrbp_1 _1806_ (.CLK(net316),
    .RESET_B(_0117_),
    .D(\stop.syn.filt.m2.sum[16] ),
    .Q_N(_0786_),
    .Q(\stop.syn.filt.m2.sum_in2[15] ));
 sg13g2_dfrbp_1 _1807_ (.CLK(net322),
    .RESET_B(_0118_),
    .D(\stop.syn.filt.m1.sum[1] ),
    .Q_N(_0785_),
    .Q(\stop.syn.filt.m1.sum_in2[0] ));
 sg13g2_dfrbp_1 _1808_ (.CLK(net323),
    .RESET_B(_0119_),
    .D(\stop.syn.filt.m1.sum[2] ),
    .Q_N(_0784_),
    .Q(\stop.syn.filt.m1.sum_in2[1] ));
 sg13g2_dfrbp_1 _1809_ (.CLK(net323),
    .RESET_B(_0120_),
    .D(\stop.syn.filt.m1.sum[3] ),
    .Q_N(_0783_),
    .Q(\stop.syn.filt.m1.sum_in2[2] ));
 sg13g2_dfrbp_1 _1810_ (.CLK(net322),
    .RESET_B(_0121_),
    .D(\stop.syn.filt.m1.sum[4] ),
    .Q_N(_0048_),
    .Q(\stop.syn.filt.m1.sum_in2[3] ));
 sg13g2_dfrbp_1 _1811_ (.CLK(net322),
    .RESET_B(_0122_),
    .D(\stop.syn.filt.m1.sum[5] ),
    .Q_N(_0782_),
    .Q(\stop.syn.filt.m1.sum_in2[4] ));
 sg13g2_dfrbp_1 _1812_ (.CLK(net325),
    .RESET_B(_0123_),
    .D(\stop.syn.filt.m1.sum[6] ),
    .Q_N(_0049_),
    .Q(\stop.syn.filt.m1.sum_in2[5] ));
 sg13g2_dfrbp_1 _1813_ (.CLK(net320),
    .RESET_B(_0124_),
    .D(\stop.syn.filt.m1.sum[7] ),
    .Q_N(_0781_),
    .Q(\stop.syn.filt.m1.sum_in2[6] ));
 sg13g2_dfrbp_1 _1814_ (.CLK(net319),
    .RESET_B(_0125_),
    .D(\stop.syn.filt.m1.sum[8] ),
    .Q_N(_0780_),
    .Q(\stop.syn.filt.m1.sum_in2[7] ));
 sg13g2_dfrbp_1 _1815_ (.CLK(net319),
    .RESET_B(_0126_),
    .D(\stop.syn.filt.m1.sum[9] ),
    .Q_N(_0779_),
    .Q(\stop.syn.filt.m1.sum_in2[8] ));
 sg13g2_dfrbp_1 _1816_ (.CLK(net319),
    .RESET_B(_0127_),
    .D(\stop.syn.filt.m1.sum[10] ),
    .Q_N(_0050_),
    .Q(\stop.syn.filt.m1.sum_in2[9] ));
 sg13g2_dfrbp_1 _1817_ (.CLK(net318),
    .RESET_B(_0128_),
    .D(\stop.syn.filt.m1.sum[11] ),
    .Q_N(_0778_),
    .Q(\stop.syn.filt.m1.sum_in2[10] ));
 sg13g2_dfrbp_1 _1818_ (.CLK(net318),
    .RESET_B(_0129_),
    .D(\stop.syn.filt.m1.sum[12] ),
    .Q_N(_0777_),
    .Q(\stop.syn.filt.m1.sum_in2[11] ));
 sg13g2_dfrbp_1 _1819_ (.CLK(net318),
    .RESET_B(_0130_),
    .D(\stop.syn.filt.m1.sum[13] ),
    .Q_N(_0776_),
    .Q(\stop.syn.filt.m1.sum_in2[12] ));
 sg13g2_dfrbp_1 _1820_ (.CLK(net318),
    .RESET_B(_0131_),
    .D(\stop.syn.filt.m1.sum[14] ),
    .Q_N(_0051_),
    .Q(\stop.syn.filt.m1.sum_in2[13] ));
 sg13g2_dfrbp_1 _1821_ (.CLK(net318),
    .RESET_B(_0132_),
    .D(\stop.syn.filt.m1.sum[15] ),
    .Q_N(_0775_),
    .Q(\stop.syn.filt.m1.sum_in2[14] ));
 sg13g2_dfrbp_1 _1822_ (.CLK(net325),
    .RESET_B(_0133_),
    .D(\stop.syn.filt.m1.sum[16] ),
    .Q_N(_0881_),
    .Q(\stop.syn.filt.m1.sum_in2[15] ));
 sg13g2_dfrbp_1 _1823_ (.CLK(net303),
    .RESET_B(\stop.merge_rstn ),
    .D(_0054_),
    .Q_N(_0882_),
    .Q(\stop.syn.daci.din[0] ));
 sg13g2_dfrbp_1 _1824_ (.CLK(net302),
    .RESET_B(net328),
    .D(_0061_),
    .Q_N(_0883_),
    .Q(\stop.syn.daci.din[1] ));
 sg13g2_dfrbp_1 _1825_ (.CLK(net302),
    .RESET_B(net328),
    .D(_0062_),
    .Q_N(_0884_),
    .Q(\stop.syn.daci.din[2] ));
 sg13g2_dfrbp_1 _1826_ (.CLK(net303),
    .RESET_B(net328),
    .D(_0063_),
    .Q_N(_0885_),
    .Q(\stop.syn.daci.din[3] ));
 sg13g2_dfrbp_1 _1827_ (.CLK(net302),
    .RESET_B(net328),
    .D(_0064_),
    .Q_N(_0886_),
    .Q(\stop.syn.daci.din[4] ));
 sg13g2_dfrbp_1 _1828_ (.CLK(net302),
    .RESET_B(\stop.merge_rstn ),
    .D(_0065_),
    .Q_N(_0887_),
    .Q(\stop.syn.daci.din[5] ));
 sg13g2_dfrbp_1 _1829_ (.CLK(net302),
    .RESET_B(\stop.merge_rstn ),
    .D(_0066_),
    .Q_N(_0888_),
    .Q(\stop.syn.daci.din[6] ));
 sg13g2_dfrbp_1 _1830_ (.CLK(net302),
    .RESET_B(net327),
    .D(_0067_),
    .Q_N(_0889_),
    .Q(\stop.syn.daci.din[7] ));
 sg13g2_dfrbp_1 _1831_ (.CLK(net300),
    .RESET_B(net327),
    .D(_0068_),
    .Q_N(_0890_),
    .Q(\stop.syn.daci.din[8] ));
 sg13g2_dfrbp_1 _1832_ (.CLK(net301),
    .RESET_B(net328),
    .D(_0069_),
    .Q_N(_0891_),
    .Q(\stop.syn.daci.din[9] ));
 sg13g2_dfrbp_1 _1833_ (.CLK(net300),
    .RESET_B(net328),
    .D(_0055_),
    .Q_N(_0892_),
    .Q(\stop.syn.daci.din[10] ));
 sg13g2_dfrbp_1 _1834_ (.CLK(net300),
    .RESET_B(net328),
    .D(_0056_),
    .Q_N(_0893_),
    .Q(\stop.syn.daci.din[11] ));
 sg13g2_dfrbp_1 _1835_ (.CLK(net300),
    .RESET_B(net327),
    .D(_0057_),
    .Q_N(_0894_),
    .Q(\stop.syn.daci.din[12] ));
 sg13g2_dfrbp_1 _1836_ (.CLK(net300),
    .RESET_B(net327),
    .D(_0058_),
    .Q_N(_0895_),
    .Q(\stop.syn.daci.din[13] ));
 sg13g2_dfrbp_1 _1837_ (.CLK(net300),
    .RESET_B(net327),
    .D(_0059_),
    .Q_N(_0896_),
    .Q(\stop.syn.daci.din[14] ));
 sg13g2_dfrbp_1 _1838_ (.CLK(net302),
    .RESET_B(net327),
    .D(_0060_),
    .Q_N(_0774_),
    .Q(\stop.syn.daci.din[15] ));
 sg13g2_dfrbp_1 _1839_ (.CLK(net314),
    .RESET_B(net100),
    .D(_0158_),
    .Q_N(_0773_),
    .Q(\stop.syn.filt.m1.b_latched[7] ));
 sg13g2_dfrbp_1 _1840_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net99),
    .D(_0159_),
    .Q_N(_0772_),
    .Q(\stop.syn.daci.accumulator[0] ));
 sg13g2_dfrbp_1 _1841_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net98),
    .D(net120),
    .Q_N(_0771_),
    .Q(\stop.syn.daci.accumulator[1] ));
 sg13g2_dfrbp_1 _1842_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net97),
    .D(_0161_),
    .Q_N(_0770_),
    .Q(\stop.syn.daci.accumulator[2] ));
 sg13g2_dfrbp_1 _1843_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net96),
    .D(net125),
    .Q_N(_0769_),
    .Q(\stop.syn.daci.accumulator[3] ));
 sg13g2_dfrbp_1 _1844_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net95),
    .D(_0163_),
    .Q_N(_0768_),
    .Q(\stop.syn.daci.accumulator[4] ));
 sg13g2_dfrbp_1 _1845_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net94),
    .D(net135),
    .Q_N(_0767_),
    .Q(\stop.syn.daci.accumulator[5] ));
 sg13g2_dfrbp_1 _1846_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net93),
    .D(net131),
    .Q_N(_0766_),
    .Q(\stop.syn.daci.accumulator[6] ));
 sg13g2_dfrbp_1 _1847_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net92),
    .D(_0166_),
    .Q_N(_0765_),
    .Q(\stop.syn.daci.accumulator[7] ));
 sg13g2_dfrbp_1 _1848_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net91),
    .D(net133),
    .Q_N(_0764_),
    .Q(\stop.syn.daci.accumulator[8] ));
 sg13g2_dfrbp_1 _1849_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net90),
    .D(_0168_),
    .Q_N(_0763_),
    .Q(\stop.syn.daci.accumulator[9] ));
 sg13g2_dfrbp_1 _1850_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net89),
    .D(net129),
    .Q_N(_0762_),
    .Q(\stop.syn.daci.accumulator[10] ));
 sg13g2_dfrbp_1 _1851_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net88),
    .D(_0170_),
    .Q_N(_0761_),
    .Q(\stop.syn.daci.accumulator[11] ));
 sg13g2_dfrbp_1 _1852_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net87),
    .D(_0171_),
    .Q_N(_0760_),
    .Q(\stop.syn.daci.accumulator[12] ));
 sg13g2_dfrbp_1 _1853_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net86),
    .D(_0172_),
    .Q_N(_0759_),
    .Q(\stop.syn.daci.accumulator[13] ));
 sg13g2_dfrbp_1 _1854_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net84),
    .D(_0173_),
    .Q_N(_0758_),
    .Q(\stop.syn.daci.accumulator[14] ));
 sg13g2_dfrbp_1 _1855_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net39),
    .D(_0174_),
    .Q_N(_0757_),
    .Q(\stop.syn.daci.accumulator[15] ));
 sg13g2_dfrbp_1 _1856_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net38),
    .D(net122),
    .Q_N(_0756_),
    .Q(data));
 sg13g2_dfrbp_1 _1857_ (.CLK(net349),
    .RESET_B(net360),
    .D(_0176_),
    .Q_N(_0755_),
    .Q(\stop.adsr_ai[0] ));
 sg13g2_dfrbp_1 _1858_ (.CLK(net348),
    .RESET_B(net359),
    .D(_0177_),
    .Q_N(_0754_),
    .Q(\stop.adsr_ai[1] ));
 sg13g2_dfrbp_1 _1859_ (.CLK(net350),
    .RESET_B(net361),
    .D(_0178_),
    .Q_N(_0753_),
    .Q(\stop.adsr_ai[2] ));
 sg13g2_dfrbp_1 _1860_ (.CLK(net350),
    .RESET_B(net361),
    .D(_0179_),
    .Q_N(_0752_),
    .Q(\stop.adsr_ai[3] ));
 sg13g2_dfrbp_1 _1861_ (.CLK(net350),
    .RESET_B(net361),
    .D(_0180_),
    .Q_N(_0751_),
    .Q(\stop.adsr_ai[4] ));
 sg13g2_dfrbp_1 _1862_ (.CLK(net345),
    .RESET_B(net356),
    .D(_0181_),
    .Q_N(_0750_),
    .Q(\stop.adsr_ai[5] ));
 sg13g2_dfrbp_1 _1863_ (.CLK(net345),
    .RESET_B(net356),
    .D(_0182_),
    .Q_N(_0749_),
    .Q(\stop.adsr_ai[6] ));
 sg13g2_dfrbp_1 _1864_ (.CLK(net348),
    .RESET_B(net359),
    .D(_0183_),
    .Q_N(_0748_),
    .Q(\stop.adsr_ai[7] ));
 sg13g2_dfrbp_1 _1865_ (.CLK(net348),
    .RESET_B(net359),
    .D(_0184_),
    .Q_N(_0747_),
    .Q(\stop.adsr_di[0] ));
 sg13g2_dfrbp_1 _1866_ (.CLK(net348),
    .RESET_B(net359),
    .D(_0185_),
    .Q_N(_0746_),
    .Q(\stop.adsr_di[1] ));
 sg13g2_dfrbp_1 _1867_ (.CLK(net348),
    .RESET_B(net359),
    .D(_0186_),
    .Q_N(_0745_),
    .Q(\stop.adsr_di[2] ));
 sg13g2_dfrbp_1 _1868_ (.CLK(net348),
    .RESET_B(net359),
    .D(_0187_),
    .Q_N(_0744_),
    .Q(\stop.adsr_di[3] ));
 sg13g2_dfrbp_1 _1869_ (.CLK(net350),
    .RESET_B(net361),
    .D(_0188_),
    .Q_N(_0743_),
    .Q(\stop.adsr_di[4] ));
 sg13g2_dfrbp_1 _1870_ (.CLK(net350),
    .RESET_B(net361),
    .D(_0189_),
    .Q_N(_0742_),
    .Q(\stop.adsr_di[5] ));
 sg13g2_dfrbp_1 _1871_ (.CLK(net345),
    .RESET_B(net356),
    .D(_0190_),
    .Q_N(_0741_),
    .Q(\stop.adsr_di[6] ));
 sg13g2_dfrbp_1 _1872_ (.CLK(net345),
    .RESET_B(net356),
    .D(_0191_),
    .Q_N(_0740_),
    .Q(\stop.adsr_di[7] ));
 sg13g2_dfrbp_1 _1873_ (.CLK(net345),
    .RESET_B(net356),
    .D(_0192_),
    .Q_N(_0739_),
    .Q(\stop.adsr_s[0] ));
 sg13g2_dfrbp_1 _1874_ (.CLK(net345),
    .RESET_B(net356),
    .D(_0193_),
    .Q_N(_0738_),
    .Q(\stop.adsr_s[1] ));
 sg13g2_dfrbp_1 _1875_ (.CLK(net345),
    .RESET_B(net356),
    .D(_0194_),
    .Q_N(_0737_),
    .Q(\stop.adsr_s[2] ));
 sg13g2_dfrbp_1 _1876_ (.CLK(net346),
    .RESET_B(net357),
    .D(_0195_),
    .Q_N(_0736_),
    .Q(\stop.adsr_s[3] ));
 sg13g2_dfrbp_1 _1877_ (.CLK(net346),
    .RESET_B(net357),
    .D(_0196_),
    .Q_N(_0735_),
    .Q(\stop.adsr_s[4] ));
 sg13g2_dfrbp_1 _1878_ (.CLK(net344),
    .RESET_B(net355),
    .D(_0197_),
    .Q_N(_0734_),
    .Q(\stop.adsr_s[5] ));
 sg13g2_dfrbp_1 _1879_ (.CLK(net343),
    .RESET_B(net354),
    .D(_0198_),
    .Q_N(_0733_),
    .Q(\stop.adsr_s[6] ));
 sg13g2_dfrbp_1 _1880_ (.CLK(net350),
    .RESET_B(net361),
    .D(_0199_),
    .Q_N(_0732_),
    .Q(\stop.adsr_s[7] ));
 sg13g2_dfrbp_1 _1881_ (.CLK(net349),
    .RESET_B(net360),
    .D(_0200_),
    .Q_N(_0731_),
    .Q(\stop.adsr_ri[0] ));
 sg13g2_dfrbp_1 _1882_ (.CLK(net348),
    .RESET_B(net359),
    .D(_0201_),
    .Q_N(_0730_),
    .Q(\stop.adsr_ri[1] ));
 sg13g2_dfrbp_1 _1883_ (.CLK(net349),
    .RESET_B(net360),
    .D(_0202_),
    .Q_N(_0729_),
    .Q(\stop.adsr_ri[2] ));
 sg13g2_dfrbp_1 _1884_ (.CLK(net348),
    .RESET_B(net359),
    .D(_0203_),
    .Q_N(_0728_),
    .Q(\stop.adsr_ri[3] ));
 sg13g2_dfrbp_1 _1885_ (.CLK(net350),
    .RESET_B(net361),
    .D(_0204_),
    .Q_N(_0727_),
    .Q(\stop.adsr_ri[4] ));
 sg13g2_dfrbp_1 _1886_ (.CLK(net350),
    .RESET_B(net361),
    .D(_0205_),
    .Q_N(_0726_),
    .Q(\stop.adsr_ri[5] ));
 sg13g2_dfrbp_1 _1887_ (.CLK(net345),
    .RESET_B(net356),
    .D(_0206_),
    .Q_N(_0725_),
    .Q(\stop.adsr_ri[6] ));
 sg13g2_dfrbp_1 _1888_ (.CLK(net343),
    .RESET_B(net354),
    .D(_0207_),
    .Q_N(_0724_),
    .Q(\stop.adsr_ri[7] ));
 sg13g2_dfrbp_1 _1889_ (.CLK(net343),
    .RESET_B(net354),
    .D(_0208_),
    .Q_N(_0723_),
    .Q(\stop.ctrl.cfg[32] ));
 sg13g2_dfrbp_1 _1890_ (.CLK(net343),
    .RESET_B(net354),
    .D(_0209_),
    .Q_N(_0722_),
    .Q(\stop.ctrl.cfg[33] ));
 sg13g2_dfrbp_1 _1891_ (.CLK(net343),
    .RESET_B(net354),
    .D(_0210_),
    .Q_N(_0721_),
    .Q(\stop.ctrl.cfg[34] ));
 sg13g2_dfrbp_1 _1892_ (.CLK(net343),
    .RESET_B(net354),
    .D(_0211_),
    .Q_N(_0720_),
    .Q(\stop.ctrl.cfg[35] ));
 sg13g2_dfrbp_1 _1893_ (.CLK(net343),
    .RESET_B(net354),
    .D(_0212_),
    .Q_N(_0719_),
    .Q(\stop.ctrl.cfg[36] ));
 sg13g2_dfrbp_1 _1894_ (.CLK(net343),
    .RESET_B(net354),
    .D(_0213_),
    .Q_N(_0718_),
    .Q(\stop.ctrl.cfg[37] ));
 sg13g2_dfrbp_1 _1895_ (.CLK(net344),
    .RESET_B(net355),
    .D(_0214_),
    .Q_N(_0717_),
    .Q(\stop.ctrl.cfg[38] ));
 sg13g2_dfrbp_1 _1896_ (.CLK(net344),
    .RESET_B(net355),
    .D(_0215_),
    .Q_N(_0716_),
    .Q(\stop.ctrl.cfg[39] ));
 sg13g2_dfrbp_1 _1897_ (.CLK(net344),
    .RESET_B(net355),
    .D(_0216_),
    .Q_N(_0715_),
    .Q(\stop.ctrl.cfg[40] ));
 sg13g2_dfrbp_1 _1898_ (.CLK(net344),
    .RESET_B(net355),
    .D(_0217_),
    .Q_N(_0714_),
    .Q(\stop.ctrl.cfg[41] ));
 sg13g2_dfrbp_1 _1899_ (.CLK(net347),
    .RESET_B(net358),
    .D(_0218_),
    .Q_N(_0713_),
    .Q(\stop.ctrl.cfg[42] ));
 sg13g2_dfrbp_1 _1900_ (.CLK(net347),
    .RESET_B(net358),
    .D(_0219_),
    .Q_N(_0712_),
    .Q(\stop.ctrl.cfg[43] ));
 sg13g2_dfrbp_1 _1901_ (.CLK(net347),
    .RESET_B(net358),
    .D(_0220_),
    .Q_N(_0711_),
    .Q(\stop.ctrl.cfg[44] ));
 sg13g2_dfrbp_1 _1902_ (.CLK(net347),
    .RESET_B(net358),
    .D(_0221_),
    .Q_N(_0710_),
    .Q(\stop.ctrl.cfg[45] ));
 sg13g2_dfrbp_1 _1903_ (.CLK(net347),
    .RESET_B(net358),
    .D(_0222_),
    .Q_N(_0709_),
    .Q(\stop.ctrl.cfg[46] ));
 sg13g2_dfrbp_1 _1904_ (.CLK(net347),
    .RESET_B(net358),
    .D(_0223_),
    .Q_N(_0708_),
    .Q(\stop.ctrl.cfg[47] ));
 sg13g2_dfrbp_1 _1905_ (.CLK(net347),
    .RESET_B(net358),
    .D(_0224_),
    .Q_N(_0707_),
    .Q(\stop.ctrl.cfg[48] ));
 sg13g2_dfrbp_1 _1906_ (.CLK(net353),
    .RESET_B(net364),
    .D(_0225_),
    .Q_N(_0706_),
    .Q(\stop.ctrl.cfg[49] ));
 sg13g2_dfrbp_1 _1907_ (.CLK(net353),
    .RESET_B(net364),
    .D(_0226_),
    .Q_N(_0705_),
    .Q(\stop.ctrl.cfg[50] ));
 sg13g2_dfrbp_1 _1908_ (.CLK(net352),
    .RESET_B(net363),
    .D(_0227_),
    .Q_N(_0704_),
    .Q(\stop.ctrl.cfg[51] ));
 sg13g2_dfrbp_1 _1909_ (.CLK(net351),
    .RESET_B(net363),
    .D(_0228_),
    .Q_N(_0703_),
    .Q(\stop.ctrl.cfg[52] ));
 sg13g2_dfrbp_1 _1910_ (.CLK(net351),
    .RESET_B(net363),
    .D(_0229_),
    .Q_N(_0702_),
    .Q(\stop.ctrl.cfg[53] ));
 sg13g2_dfrbp_1 _1911_ (.CLK(net352),
    .RESET_B(net362),
    .D(_0230_),
    .Q_N(_0701_),
    .Q(\stop.ctrl.cfg[54] ));
 sg13g2_dfrbp_1 _1912_ (.CLK(net352),
    .RESET_B(net362),
    .D(_0231_),
    .Q_N(_0700_),
    .Q(\stop.ctrl.cfg[55] ));
 sg13g2_dfrbp_1 _1913_ (.CLK(net351),
    .RESET_B(net362),
    .D(_0232_),
    .Q_N(_0699_),
    .Q(\stop.ctrl.cfg[56] ));
 sg13g2_dfrbp_1 _1914_ (.CLK(net351),
    .RESET_B(net362),
    .D(_0233_),
    .Q_N(_0698_),
    .Q(\stop.ctrl.cfg[57] ));
 sg13g2_dfrbp_1 _1915_ (.CLK(net351),
    .RESET_B(net362),
    .D(_0234_),
    .Q_N(_0697_),
    .Q(\stop.ctrl.cfg[58] ));
 sg13g2_dfrbp_1 _1916_ (.CLK(net351),
    .RESET_B(net362),
    .D(_0235_),
    .Q_N(_0696_),
    .Q(\stop.ctrl.cfg[59] ));
 sg13g2_tiehi _1689__28 (.L_HI(net28));
 sg13g2_tiehi _1685__29 (.L_HI(net29));
 sg13g2_tiehi _1686__30 (.L_HI(net30));
 sg13g2_tiehi _1687__31 (.L_HI(net31));
 sg13g2_tiehi _1758__32 (.L_HI(net32));
 sg13g2_tiehi _1757__33 (.L_HI(net33));
 sg13g2_tiehi _1756__34 (.L_HI(net34));
 sg13g2_tiehi _1755__35 (.L_HI(net35));
 sg13g2_tiehi _1754__36 (.L_HI(net36));
 sg13g2_tiehi _1753__37 (.L_HI(net37));
 sg13g2_tiehi _1856__38 (.L_HI(net38));
 sg13g2_tiehi _1855__39 (.L_HI(net39));
 sg13g2_tiehi _1711__40 (.L_HI(net40));
 sg13g2_tiehi _1710__41 (.L_HI(net41));
 sg13g2_tiehi _1709__42 (.L_HI(net42));
 sg13g2_tiehi _1708__43 (.L_HI(net43));
 sg13g2_tiehi _1707__44 (.L_HI(net44));
 sg13g2_tiehi _1706__45 (.L_HI(net45));
 sg13g2_tiehi _1688__46 (.L_HI(net46));
 sg13g2_tiehi _1715__47 (.L_HI(net47));
 sg13g2_tiehi _1716__48 (.L_HI(net48));
 sg13g2_tiehi _1717__49 (.L_HI(net49));
 sg13g2_tiehi _1718__50 (.L_HI(net50));
 sg13g2_tiehi _1719__51 (.L_HI(net51));
 sg13g2_tiehi _1720__52 (.L_HI(net52));
 sg13g2_tiehi _1721__53 (.L_HI(net53));
 sg13g2_tiehi _1722__54 (.L_HI(net54));
 sg13g2_tiehi _1723__55 (.L_HI(net55));
 sg13g2_tiehi _1724__56 (.L_HI(net56));
 sg13g2_tiehi _1725__57 (.L_HI(net57));
 sg13g2_tiehi _1726__58 (.L_HI(net58));
 sg13g2_tiehi _1727__59 (.L_HI(net59));
 sg13g2_tiehi _1728__60 (.L_HI(net60));
 sg13g2_tiehi _1729__61 (.L_HI(net61));
 sg13g2_tiehi _1730__62 (.L_HI(net62));
 sg13g2_tiehi _1731__63 (.L_HI(net63));
 sg13g2_tiehi _1732__64 (.L_HI(net64));
 sg13g2_tiehi _1733__65 (.L_HI(net65));
 sg13g2_tiehi _1734__66 (.L_HI(net66));
 sg13g2_tiehi _1735__67 (.L_HI(net67));
 sg13g2_tiehi _1736__68 (.L_HI(net68));
 sg13g2_tiehi _1705__69 (.L_HI(net69));
 sg13g2_tiehi _1704__70 (.L_HI(net70));
 sg13g2_tiehi _1703__71 (.L_HI(net71));
 sg13g2_tiehi _1702__72 (.L_HI(net72));
 sg13g2_tiehi _1701__73 (.L_HI(net73));
 sg13g2_tiehi _1700__74 (.L_HI(net74));
 sg13g2_tiehi _1699__75 (.L_HI(net75));
 sg13g2_tiehi _1698__76 (.L_HI(net76));
 sg13g2_tiehi _1697__77 (.L_HI(net77));
 sg13g2_tiehi _1696__78 (.L_HI(net78));
 sg13g2_tiehi _1695__79 (.L_HI(net79));
 sg13g2_tiehi _1694__80 (.L_HI(net80));
 sg13g2_tiehi _1693__81 (.L_HI(net81));
 sg13g2_tiehi _1692__82 (.L_HI(net82));
 sg13g2_tiehi _1691__83 (.L_HI(net83));
 sg13g2_tiehi _1854__84 (.L_HI(net84));
 sg13g2_tiehi _1690__85 (.L_HI(net85));
 sg13g2_tiehi _1853__86 (.L_HI(net86));
 sg13g2_tiehi _1852__87 (.L_HI(net87));
 sg13g2_tiehi _1851__88 (.L_HI(net88));
 sg13g2_tiehi _1850__89 (.L_HI(net89));
 sg13g2_tiehi _1849__90 (.L_HI(net90));
 sg13g2_tiehi _1848__91 (.L_HI(net91));
 sg13g2_tiehi _1847__92 (.L_HI(net92));
 sg13g2_tiehi _1846__93 (.L_HI(net93));
 sg13g2_tiehi _1845__94 (.L_HI(net94));
 sg13g2_tiehi _1844__95 (.L_HI(net95));
 sg13g2_tiehi _1843__96 (.L_HI(net96));
 sg13g2_tiehi _1842__97 (.L_HI(net97));
 sg13g2_tiehi _1841__98 (.L_HI(net98));
 sg13g2_tiehi _1840__99 (.L_HI(net99));
 sg13g2_tiehi _1839__100 (.L_HI(net100));
 sg13g2_tiehi _1774__101 (.L_HI(net101));
 sg13g2_tiehi _1773__102 (.L_HI(net102));
 sg13g2_tiehi _1772__103 (.L_HI(net103));
 sg13g2_tiehi _1771__104 (.L_HI(net104));
 sg13g2_tiehi _1770__105 (.L_HI(net105));
 sg13g2_tiehi _1769__106 (.L_HI(net106));
 sg13g2_tiehi _1768__107 (.L_HI(net107));
 sg13g2_tiehi _1767__108 (.L_HI(net108));
 sg13g2_tiehi _1766__109 (.L_HI(net109));
 sg13g2_tiehi _1765__110 (.L_HI(net110));
 sg13g2_tiehi _1764__111 (.L_HI(net111));
 sg13g2_tiehi _1763__112 (.L_HI(net112));
 sg13g2_tiehi _1762__113 (.L_HI(net113));
 sg13g2_tiehi _1761__114 (.L_HI(net114));
 sg13g2_tiehi _1760__115 (.L_HI(net115));
 sg13g2_tiehi _1714__116 (.L_HI(net116));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_kch_cd101_5 (.L_LO(net5));
 sg13g2_tielo tt_um_kch_cd101_6 (.L_LO(net6));
 sg13g2_tielo tt_um_kch_cd101_7 (.L_LO(net7));
 sg13g2_tielo tt_um_kch_cd101_8 (.L_LO(net8));
 sg13g2_tielo tt_um_kch_cd101_9 (.L_LO(net9));
 sg13g2_tielo tt_um_kch_cd101_10 (.L_LO(net10));
 sg13g2_tielo tt_um_kch_cd101_11 (.L_LO(net11));
 sg13g2_tielo tt_um_kch_cd101_12 (.L_LO(net12));
 sg13g2_tielo tt_um_kch_cd101_13 (.L_LO(net13));
 sg13g2_tielo tt_um_kch_cd101_14 (.L_LO(net14));
 sg13g2_tielo tt_um_kch_cd101_15 (.L_LO(net15));
 sg13g2_tielo tt_um_kch_cd101_16 (.L_LO(net16));
 sg13g2_tielo tt_um_kch_cd101_17 (.L_LO(net17));
 sg13g2_tielo tt_um_kch_cd101_18 (.L_LO(net18));
 sg13g2_tielo tt_um_kch_cd101_19 (.L_LO(net19));
 sg13g2_tielo tt_um_kch_cd101_20 (.L_LO(net20));
 sg13g2_tielo tt_um_kch_cd101_21 (.L_LO(net21));
 sg13g2_tielo tt_um_kch_cd101_22 (.L_LO(net22));
 sg13g2_tielo tt_um_kch_cd101_23 (.L_LO(net23));
 sg13g2_tielo tt_um_kch_cd101_24 (.L_LO(net24));
 sg13g2_tielo tt_um_kch_cd101_25 (.L_LO(net25));
 sg13g2_tielo tt_um_kch_cd101_26 (.L_LO(net26));
 sg13g2_tiehi _1759__27 (.L_HI(net27));
 sg13g2_buf_1 _2030_ (.A(data),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout278 (.A(_0643_),
    .X(net278));
 sg13g2_buf_2 fanout279 (.A(net280),
    .X(net279));
 sg13g2_buf_2 fanout280 (.A(net281),
    .X(net280));
 sg13g2_buf_2 fanout281 (.A(\stop.syn.adsri.rstn ),
    .X(net281));
 sg13g2_buf_4 fanout282 (.X(net282),
    .A(\stop.syn.adsri.state[2] ));
 sg13g2_buf_2 fanout283 (.A(\stop.syn.adsri.state[1] ),
    .X(net283));
 sg13g2_buf_1 fanout284 (.A(\stop.syn.adsri.state[1] ),
    .X(net284));
 sg13g2_buf_2 fanout285 (.A(net286),
    .X(net285));
 sg13g2_buf_2 fanout286 (.A(\stop.syn.adsri.clk ),
    .X(net286));
 sg13g2_buf_4 fanout287 (.X(net287),
    .A(net288));
 sg13g2_buf_2 fanout288 (.A(_0313_),
    .X(net288));
 sg13g2_buf_2 fanout289 (.A(net291),
    .X(net289));
 sg13g2_buf_2 fanout290 (.A(net291),
    .X(net290));
 sg13g2_buf_4 fanout291 (.X(net291),
    .A(_0313_));
 sg13g2_buf_2 fanout292 (.A(net296),
    .X(net292));
 sg13g2_buf_2 fanout293 (.A(net296),
    .X(net293));
 sg13g2_buf_2 fanout294 (.A(net296),
    .X(net294));
 sg13g2_buf_4 fanout295 (.X(net295),
    .A(net296));
 sg13g2_buf_2 fanout296 (.A(_0313_),
    .X(net296));
 sg13g2_buf_2 fanout297 (.A(net298),
    .X(net297));
 sg13g2_buf_4 fanout298 (.X(net298),
    .A(net301));
 sg13g2_buf_2 fanout299 (.A(net300),
    .X(net299));
 sg13g2_buf_4 fanout300 (.X(net300),
    .A(net301));
 sg13g2_buf_2 fanout301 (.A(\stop.syn.clk_sample ),
    .X(net301));
 sg13g2_buf_4 fanout302 (.X(net302),
    .A(net303));
 sg13g2_buf_4 fanout303 (.X(net303),
    .A(\stop.syn.clk_sample ));
 sg13g2_buf_2 fanout304 (.A(net305),
    .X(net304));
 sg13g2_buf_1 fanout305 (.A(net306),
    .X(net305));
 sg13g2_buf_2 fanout306 (.A(net308),
    .X(net306));
 sg13g2_buf_2 fanout307 (.A(net308),
    .X(net307));
 sg13g2_buf_2 fanout308 (.A(\stop.syn.filt.m2.b_bit ),
    .X(net308));
 sg13g2_buf_2 fanout309 (.A(net311),
    .X(net309));
 sg13g2_buf_1 fanout310 (.A(net311),
    .X(net310));
 sg13g2_buf_2 fanout311 (.A(\stop.syn.filt.m1.b_bit ),
    .X(net311));
 sg13g2_buf_2 fanout312 (.A(net313),
    .X(net312));
 sg13g2_buf_2 fanout313 (.A(\stop.syn.filt.m1.b_bit ),
    .X(net313));
 sg13g2_buf_2 fanout314 (.A(net319),
    .X(net314));
 sg13g2_buf_2 fanout315 (.A(net319),
    .X(net315));
 sg13g2_buf_2 fanout316 (.A(net318),
    .X(net316));
 sg13g2_buf_2 fanout317 (.A(net318),
    .X(net317));
 sg13g2_buf_2 fanout318 (.A(net319),
    .X(net318));
 sg13g2_buf_2 fanout319 (.A(_0037_),
    .X(net319));
 sg13g2_buf_2 fanout320 (.A(net324),
    .X(net320));
 sg13g2_buf_1 fanout321 (.A(net324),
    .X(net321));
 sg13g2_buf_2 fanout322 (.A(net324),
    .X(net322));
 sg13g2_buf_1 fanout323 (.A(net324),
    .X(net323));
 sg13g2_buf_1 fanout324 (.A(net326),
    .X(net324));
 sg13g2_buf_4 fanout325 (.X(net325),
    .A(net326));
 sg13g2_buf_2 fanout326 (.A(_0037_),
    .X(net326));
 sg13g2_buf_4 fanout327 (.X(net327),
    .A(net328));
 sg13g2_buf_4 fanout328 (.X(net328),
    .A(\stop.merge_rstn ));
 sg13g2_buf_4 fanout329 (.X(net329),
    .A(net331));
 sg13g2_buf_2 fanout330 (.A(net331),
    .X(net330));
 sg13g2_buf_4 fanout331 (.X(net331),
    .A(net332));
 sg13g2_buf_4 fanout332 (.X(net332),
    .A(net338));
 sg13g2_buf_2 fanout333 (.A(net334),
    .X(net333));
 sg13g2_buf_2 fanout334 (.A(net337),
    .X(net334));
 sg13g2_buf_4 fanout335 (.X(net335),
    .A(net337));
 sg13g2_buf_2 fanout336 (.A(net337),
    .X(net336));
 sg13g2_buf_2 fanout337 (.A(net338),
    .X(net337));
 sg13g2_buf_4 fanout338 (.X(net338),
    .A(_0291_));
 sg13g2_buf_4 fanout339 (.X(net339),
    .A(net340));
 sg13g2_buf_2 fanout340 (.A(_0291_),
    .X(net340));
 sg13g2_buf_4 fanout341 (.X(net341),
    .A(net342));
 sg13g2_buf_4 fanout342 (.X(net342),
    .A(\stop.syn.clki.arstn ));
 sg13g2_buf_2 fanout343 (.A(net346),
    .X(net343));
 sg13g2_buf_1 fanout344 (.A(net346),
    .X(net344));
 sg13g2_buf_2 fanout345 (.A(net346),
    .X(net345));
 sg13g2_buf_1 fanout346 (.A(net347),
    .X(net346));
 sg13g2_buf_2 fanout347 (.A(net353),
    .X(net347));
 sg13g2_buf_2 fanout348 (.A(net349),
    .X(net348));
 sg13g2_buf_1 fanout349 (.A(net353),
    .X(net349));
 sg13g2_buf_2 fanout350 (.A(net353),
    .X(net350));
 sg13g2_buf_2 fanout351 (.A(net352),
    .X(net351));
 sg13g2_buf_2 fanout352 (.A(net353),
    .X(net352));
 sg13g2_buf_4 fanout353 (.X(net353),
    .A(uio_in[3]));
 sg13g2_buf_4 fanout354 (.X(net354),
    .A(net357));
 sg13g2_buf_2 fanout355 (.A(net357),
    .X(net355));
 sg13g2_buf_4 fanout356 (.X(net356),
    .A(net357));
 sg13g2_buf_2 fanout357 (.A(net358),
    .X(net357));
 sg13g2_buf_4 fanout358 (.X(net358),
    .A(net364));
 sg13g2_buf_4 fanout359 (.X(net359),
    .A(net360));
 sg13g2_buf_2 fanout360 (.A(net364),
    .X(net360));
 sg13g2_buf_4 fanout361 (.X(net361),
    .A(net364));
 sg13g2_buf_4 fanout362 (.X(net362),
    .A(net363));
 sg13g2_buf_2 fanout363 (.A(net364),
    .X(net363));
 sg13g2_buf_4 fanout364 (.X(net364),
    .A(rst_n));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(uio_in[0]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(uio_in[1]),
    .X(net3));
 sg13g2_tielo tt_um_kch_cd101_4 (.L_LO(net4));
 sg13g2_buf_2 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .X(clknet_2_0__leaf_clk));
 sg13g2_buf_2 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .X(clknet_2_1__leaf_clk));
 sg13g2_buf_2 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .X(clknet_2_2__leaf_clk));
 sg13g2_buf_2 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .X(clknet_2_3__leaf_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(_0027_),
    .X(net117));
 sg13g2_dlygate4sd3_1 hold2 (.A(\stop.syn.rstn_fst_reg1 ),
    .X(net118));
 sg13g2_dlygate4sd3_1 hold3 (.A(\stop.syn.daci.accumulator[0] ),
    .X(net119));
 sg13g2_dlygate4sd3_1 hold4 (.A(_0160_),
    .X(net120));
 sg13g2_dlygate4sd3_1 hold5 (.A(\stop.syn.daci.accumulator[15] ),
    .X(net121));
 sg13g2_dlygate4sd3_1 hold6 (.A(_0175_),
    .X(net122));
 sg13g2_dlygate4sd3_1 hold7 (.A(\stop.syn.daci.accumulator[12] ),
    .X(net123));
 sg13g2_dlygate4sd3_1 hold8 (.A(\stop.syn.daci.accumulator[3] ),
    .X(net124));
 sg13g2_dlygate4sd3_1 hold9 (.A(_0162_),
    .X(net125));
 sg13g2_dlygate4sd3_1 hold10 (.A(\stop.syn.daci.accumulator[14] ),
    .X(net126));
 sg13g2_dlygate4sd3_1 hold11 (.A(\stop.syn.daci.accumulator[13] ),
    .X(net127));
 sg13g2_dlygate4sd3_1 hold12 (.A(\stop.syn.daci.accumulator[10] ),
    .X(net128));
 sg13g2_dlygate4sd3_1 hold13 (.A(_0169_),
    .X(net129));
 sg13g2_dlygate4sd3_1 hold14 (.A(\stop.syn.daci.accumulator[6] ),
    .X(net130));
 sg13g2_dlygate4sd3_1 hold15 (.A(_0165_),
    .X(net131));
 sg13g2_dlygate4sd3_1 hold16 (.A(\stop.syn.daci.accumulator[8] ),
    .X(net132));
 sg13g2_dlygate4sd3_1 hold17 (.A(_0167_),
    .X(net133));
 sg13g2_dlygate4sd3_1 hold18 (.A(\stop.syn.daci.accumulator[5] ),
    .X(net134));
 sg13g2_dlygate4sd3_1 hold19 (.A(_0164_),
    .X(net135));
 sg13g2_dlygate4sd3_1 hold20 (.A(\stop.syn.daci.accumulator[9] ),
    .X(net136));
 sg13g2_dlygate4sd3_1 hold21 (.A(\stop.syn.daci.accumulator[11] ),
    .X(net137));
 sg13g2_dlygate4sd3_1 hold22 (.A(\stop.syn.daci.accumulator[7] ),
    .X(net138));
 sg13g2_dlygate4sd3_1 hold23 (.A(\stop.syn.daci.accumulator[2] ),
    .X(net139));
 sg13g2_dlygate4sd3_1 hold24 (.A(_0676_),
    .X(net140));
 sg13g2_dlygate4sd3_1 hold25 (.A(\stop.syn.daci.accumulator[4] ),
    .X(net141));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_fill_2 FILLER_0_238 ();
 sg13g2_fill_1 FILLER_0_240 ();
 sg13g2_decap_4 FILLER_0_267 ();
 sg13g2_fill_1 FILLER_0_271 ();
 sg13g2_decap_4 FILLER_0_298 ();
 sg13g2_fill_2 FILLER_0_302 ();
 sg13g2_decap_8 FILLER_0_330 ();
 sg13g2_decap_8 FILLER_0_337 ();
 sg13g2_decap_8 FILLER_0_344 ();
 sg13g2_decap_8 FILLER_0_351 ();
 sg13g2_decap_4 FILLER_0_358 ();
 sg13g2_fill_2 FILLER_0_362 ();
 sg13g2_decap_8 FILLER_0_390 ();
 sg13g2_decap_8 FILLER_0_397 ();
 sg13g2_decap_4 FILLER_0_404 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_4 FILLER_1_70 ();
 sg13g2_fill_1 FILLER_1_74 ();
 sg13g2_decap_8 FILLER_1_83 ();
 sg13g2_decap_8 FILLER_1_90 ();
 sg13g2_decap_8 FILLER_1_97 ();
 sg13g2_decap_8 FILLER_1_104 ();
 sg13g2_decap_8 FILLER_1_121 ();
 sg13g2_decap_8 FILLER_1_128 ();
 sg13g2_fill_1 FILLER_1_135 ();
 sg13g2_decap_8 FILLER_1_146 ();
 sg13g2_decap_8 FILLER_1_153 ();
 sg13g2_fill_1 FILLER_1_160 ();
 sg13g2_decap_8 FILLER_1_171 ();
 sg13g2_decap_8 FILLER_1_178 ();
 sg13g2_decap_4 FILLER_1_185 ();
 sg13g2_decap_8 FILLER_1_215 ();
 sg13g2_fill_2 FILLER_1_222 ();
 sg13g2_fill_1 FILLER_1_224 ();
 sg13g2_fill_2 FILLER_1_243 ();
 sg13g2_fill_1 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_fill_2 FILLER_1_259 ();
 sg13g2_fill_1 FILLER_1_261 ();
 sg13g2_fill_1 FILLER_1_272 ();
 sg13g2_decap_8 FILLER_1_283 ();
 sg13g2_decap_4 FILLER_1_290 ();
 sg13g2_fill_2 FILLER_1_304 ();
 sg13g2_fill_1 FILLER_1_306 ();
 sg13g2_decap_8 FILLER_1_317 ();
 sg13g2_fill_2 FILLER_1_381 ();
 sg13g2_decap_8 FILLER_1_386 ();
 sg13g2_decap_8 FILLER_1_393 ();
 sg13g2_decap_8 FILLER_1_400 ();
 sg13g2_fill_2 FILLER_1_407 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_fill_2 FILLER_2_7 ();
 sg13g2_decap_4 FILLER_2_73 ();
 sg13g2_fill_1 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_192 ();
 sg13g2_decap_4 FILLER_2_199 ();
 sg13g2_fill_2 FILLER_2_229 ();
 sg13g2_fill_1 FILLER_2_240 ();
 sg13g2_decap_4 FILLER_2_277 ();
 sg13g2_fill_1 FILLER_2_281 ();
 sg13g2_decap_4 FILLER_2_308 ();
 sg13g2_fill_2 FILLER_2_312 ();
 sg13g2_fill_1 FILLER_2_340 ();
 sg13g2_fill_2 FILLER_2_351 ();
 sg13g2_fill_1 FILLER_2_353 ();
 sg13g2_decap_8 FILLER_2_394 ();
 sg13g2_decap_8 FILLER_2_401 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_fill_1 FILLER_3_0 ();
 sg13g2_decap_4 FILLER_3_31 ();
 sg13g2_fill_2 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_fill_2 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_88 ();
 sg13g2_decap_8 FILLER_3_121 ();
 sg13g2_decap_8 FILLER_3_128 ();
 sg13g2_decap_4 FILLER_3_135 ();
 sg13g2_fill_1 FILLER_3_139 ();
 sg13g2_decap_8 FILLER_3_148 ();
 sg13g2_decap_8 FILLER_3_155 ();
 sg13g2_decap_8 FILLER_3_162 ();
 sg13g2_decap_8 FILLER_3_169 ();
 sg13g2_fill_1 FILLER_3_176 ();
 sg13g2_decap_8 FILLER_3_213 ();
 sg13g2_decap_8 FILLER_3_220 ();
 sg13g2_fill_1 FILLER_3_227 ();
 sg13g2_fill_2 FILLER_3_250 ();
 sg13g2_decap_8 FILLER_3_256 ();
 sg13g2_decap_4 FILLER_3_263 ();
 sg13g2_fill_2 FILLER_3_270 ();
 sg13g2_decap_8 FILLER_3_278 ();
 sg13g2_fill_2 FILLER_3_285 ();
 sg13g2_decap_4 FILLER_3_292 ();
 sg13g2_decap_8 FILLER_3_306 ();
 sg13g2_decap_8 FILLER_3_313 ();
 sg13g2_decap_4 FILLER_3_333 ();
 sg13g2_decap_4 FILLER_3_343 ();
 sg13g2_fill_1 FILLER_3_347 ();
 sg13g2_decap_8 FILLER_3_353 ();
 sg13g2_fill_1 FILLER_3_360 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_4 FILLER_3_378 ();
 sg13g2_fill_1 FILLER_3_382 ();
 sg13g2_decap_4 FILLER_4_0 ();
 sg13g2_fill_1 FILLER_4_4 ();
 sg13g2_fill_2 FILLER_4_35 ();
 sg13g2_fill_1 FILLER_4_37 ();
 sg13g2_decap_4 FILLER_4_64 ();
 sg13g2_fill_2 FILLER_4_68 ();
 sg13g2_fill_1 FILLER_4_86 ();
 sg13g2_decap_8 FILLER_4_97 ();
 sg13g2_decap_8 FILLER_4_104 ();
 sg13g2_decap_8 FILLER_4_111 ();
 sg13g2_fill_2 FILLER_4_118 ();
 sg13g2_fill_1 FILLER_4_156 ();
 sg13g2_decap_8 FILLER_4_191 ();
 sg13g2_decap_4 FILLER_4_198 ();
 sg13g2_fill_1 FILLER_4_202 ();
 sg13g2_fill_2 FILLER_4_331 ();
 sg13g2_decap_4 FILLER_4_359 ();
 sg13g2_decap_8 FILLER_4_394 ();
 sg13g2_decap_8 FILLER_4_401 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_4 FILLER_5_14 ();
 sg13g2_fill_1 FILLER_5_18 ();
 sg13g2_decap_8 FILLER_5_23 ();
 sg13g2_decap_4 FILLER_5_30 ();
 sg13g2_fill_1 FILLER_5_75 ();
 sg13g2_decap_4 FILLER_5_90 ();
 sg13g2_fill_2 FILLER_5_94 ();
 sg13g2_decap_8 FILLER_5_132 ();
 sg13g2_decap_8 FILLER_5_139 ();
 sg13g2_fill_2 FILLER_5_146 ();
 sg13g2_decap_8 FILLER_5_156 ();
 sg13g2_fill_2 FILLER_5_163 ();
 sg13g2_decap_4 FILLER_5_175 ();
 sg13g2_fill_2 FILLER_5_179 ();
 sg13g2_decap_8 FILLER_5_191 ();
 sg13g2_decap_8 FILLER_5_198 ();
 sg13g2_decap_8 FILLER_5_205 ();
 sg13g2_decap_8 FILLER_5_212 ();
 sg13g2_decap_8 FILLER_5_219 ();
 sg13g2_fill_2 FILLER_5_226 ();
 sg13g2_decap_4 FILLER_5_239 ();
 sg13g2_fill_2 FILLER_5_243 ();
 sg13g2_decap_8 FILLER_5_250 ();
 sg13g2_decap_8 FILLER_5_257 ();
 sg13g2_decap_4 FILLER_5_264 ();
 sg13g2_fill_1 FILLER_5_268 ();
 sg13g2_decap_4 FILLER_5_279 ();
 sg13g2_fill_2 FILLER_5_283 ();
 sg13g2_decap_4 FILLER_5_289 ();
 sg13g2_fill_1 FILLER_5_293 ();
 sg13g2_decap_8 FILLER_5_297 ();
 sg13g2_decap_4 FILLER_5_304 ();
 sg13g2_decap_4 FILLER_5_312 ();
 sg13g2_fill_1 FILLER_5_316 ();
 sg13g2_fill_1 FILLER_5_322 ();
 sg13g2_fill_2 FILLER_5_331 ();
 sg13g2_fill_1 FILLER_5_333 ();
 sg13g2_fill_1 FILLER_5_344 ();
 sg13g2_decap_4 FILLER_5_349 ();
 sg13g2_decap_8 FILLER_5_373 ();
 sg13g2_decap_4 FILLER_5_380 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_4 FILLER_6_7 ();
 sg13g2_fill_2 FILLER_6_11 ();
 sg13g2_decap_8 FILLER_6_39 ();
 sg13g2_fill_2 FILLER_6_46 ();
 sg13g2_decap_8 FILLER_6_52 ();
 sg13g2_fill_2 FILLER_6_59 ();
 sg13g2_decap_8 FILLER_6_65 ();
 sg13g2_decap_8 FILLER_6_72 ();
 sg13g2_decap_8 FILLER_6_115 ();
 sg13g2_decap_8 FILLER_6_122 ();
 sg13g2_decap_4 FILLER_6_129 ();
 sg13g2_fill_2 FILLER_6_133 ();
 sg13g2_decap_4 FILLER_6_166 ();
 sg13g2_decap_4 FILLER_6_178 ();
 sg13g2_fill_2 FILLER_6_182 ();
 sg13g2_fill_2 FILLER_6_280 ();
 sg13g2_fill_1 FILLER_6_282 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_fill_2 FILLER_6_294 ();
 sg13g2_fill_1 FILLER_6_296 ();
 sg13g2_fill_1 FILLER_6_323 ();
 sg13g2_fill_2 FILLER_6_328 ();
 sg13g2_fill_1 FILLER_6_330 ();
 sg13g2_fill_2 FILLER_6_379 ();
 sg13g2_fill_2 FILLER_6_407 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_fill_1 FILLER_7_12 ();
 sg13g2_decap_8 FILLER_7_17 ();
 sg13g2_fill_2 FILLER_7_28 ();
 sg13g2_fill_2 FILLER_7_90 ();
 sg13g2_fill_1 FILLER_7_102 ();
 sg13g2_decap_4 FILLER_7_129 ();
 sg13g2_fill_2 FILLER_7_133 ();
 sg13g2_decap_4 FILLER_7_155 ();
 sg13g2_decap_4 FILLER_7_200 ();
 sg13g2_fill_2 FILLER_7_204 ();
 sg13g2_decap_8 FILLER_7_212 ();
 sg13g2_decap_4 FILLER_7_219 ();
 sg13g2_decap_8 FILLER_7_236 ();
 sg13g2_decap_8 FILLER_7_243 ();
 sg13g2_decap_4 FILLER_7_250 ();
 sg13g2_fill_1 FILLER_7_254 ();
 sg13g2_decap_4 FILLER_7_263 ();
 sg13g2_fill_1 FILLER_7_312 ();
 sg13g2_fill_1 FILLER_7_341 ();
 sg13g2_decap_8 FILLER_7_346 ();
 sg13g2_fill_1 FILLER_7_353 ();
 sg13g2_decap_4 FILLER_7_374 ();
 sg13g2_fill_2 FILLER_7_378 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_fill_2 FILLER_8_0 ();
 sg13g2_decap_4 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_50 ();
 sg13g2_decap_8 FILLER_8_57 ();
 sg13g2_decap_4 FILLER_8_64 ();
 sg13g2_fill_2 FILLER_8_68 ();
 sg13g2_decap_8 FILLER_8_127 ();
 sg13g2_fill_2 FILLER_8_134 ();
 sg13g2_decap_4 FILLER_8_162 ();
 sg13g2_fill_2 FILLER_8_166 ();
 sg13g2_decap_8 FILLER_8_178 ();
 sg13g2_decap_8 FILLER_8_185 ();
 sg13g2_fill_1 FILLER_8_200 ();
 sg13g2_fill_1 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_239 ();
 sg13g2_decap_8 FILLER_8_264 ();
 sg13g2_decap_8 FILLER_8_271 ();
 sg13g2_decap_8 FILLER_8_278 ();
 sg13g2_fill_1 FILLER_8_285 ();
 sg13g2_fill_2 FILLER_8_294 ();
 sg13g2_decap_4 FILLER_8_321 ();
 sg13g2_fill_2 FILLER_8_329 ();
 sg13g2_fill_1 FILLER_8_331 ();
 sg13g2_fill_1 FILLER_8_358 ();
 sg13g2_decap_4 FILLER_8_378 ();
 sg13g2_fill_2 FILLER_8_382 ();
 sg13g2_fill_2 FILLER_8_389 ();
 sg13g2_fill_1 FILLER_8_391 ();
 sg13g2_fill_2 FILLER_8_396 ();
 sg13g2_decap_8 FILLER_8_401 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_fill_2 FILLER_9_7 ();
 sg13g2_fill_2 FILLER_9_71 ();
 sg13g2_fill_1 FILLER_9_73 ();
 sg13g2_decap_8 FILLER_9_124 ();
 sg13g2_fill_2 FILLER_9_131 ();
 sg13g2_fill_1 FILLER_9_133 ();
 sg13g2_fill_2 FILLER_9_143 ();
 sg13g2_fill_1 FILLER_9_145 ();
 sg13g2_fill_2 FILLER_9_151 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_4 FILLER_9_220 ();
 sg13g2_fill_1 FILLER_9_224 ();
 sg13g2_decap_4 FILLER_9_233 ();
 sg13g2_fill_1 FILLER_9_237 ();
 sg13g2_decap_4 FILLER_9_261 ();
 sg13g2_fill_2 FILLER_9_278 ();
 sg13g2_fill_1 FILLER_9_300 ();
 sg13g2_fill_1 FILLER_9_330 ();
 sg13g2_decap_4 FILLER_9_336 ();
 sg13g2_decap_4 FILLER_9_352 ();
 sg13g2_fill_2 FILLER_9_356 ();
 sg13g2_decap_4 FILLER_9_378 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_4 FILLER_10_14 ();
 sg13g2_fill_2 FILLER_10_18 ();
 sg13g2_decap_8 FILLER_10_24 ();
 sg13g2_decap_4 FILLER_10_31 ();
 sg13g2_decap_4 FILLER_10_39 ();
 sg13g2_fill_1 FILLER_10_48 ();
 sg13g2_decap_8 FILLER_10_62 ();
 sg13g2_fill_2 FILLER_10_69 ();
 sg13g2_fill_1 FILLER_10_71 ();
 sg13g2_decap_8 FILLER_10_88 ();
 sg13g2_decap_8 FILLER_10_95 ();
 sg13g2_decap_4 FILLER_10_102 ();
 sg13g2_fill_2 FILLER_10_106 ();
 sg13g2_decap_8 FILLER_10_144 ();
 sg13g2_decap_8 FILLER_10_187 ();
 sg13g2_decap_4 FILLER_10_194 ();
 sg13g2_fill_1 FILLER_10_198 ();
 sg13g2_decap_4 FILLER_10_213 ();
 sg13g2_decap_4 FILLER_10_236 ();
 sg13g2_decap_4 FILLER_10_245 ();
 sg13g2_fill_2 FILLER_10_261 ();
 sg13g2_fill_1 FILLER_10_263 ();
 sg13g2_fill_2 FILLER_10_269 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_fill_1 FILLER_10_287 ();
 sg13g2_fill_2 FILLER_10_292 ();
 sg13g2_fill_1 FILLER_10_294 ();
 sg13g2_fill_2 FILLER_10_299 ();
 sg13g2_fill_1 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_307 ();
 sg13g2_fill_2 FILLER_10_314 ();
 sg13g2_decap_8 FILLER_10_321 ();
 sg13g2_decap_4 FILLER_10_328 ();
 sg13g2_decap_8 FILLER_10_353 ();
 sg13g2_fill_1 FILLER_10_360 ();
 sg13g2_decap_8 FILLER_10_376 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_fill_2 FILLER_11_21 ();
 sg13g2_decap_4 FILLER_11_27 ();
 sg13g2_fill_2 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_120 ();
 sg13g2_fill_1 FILLER_11_127 ();
 sg13g2_decap_4 FILLER_11_136 ();
 sg13g2_fill_2 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_146 ();
 sg13g2_fill_1 FILLER_11_153 ();
 sg13g2_decap_8 FILLER_11_159 ();
 sg13g2_decap_8 FILLER_11_166 ();
 sg13g2_decap_8 FILLER_11_173 ();
 sg13g2_decap_8 FILLER_11_180 ();
 sg13g2_fill_2 FILLER_11_187 ();
 sg13g2_decap_4 FILLER_11_215 ();
 sg13g2_fill_1 FILLER_11_219 ();
 sg13g2_fill_2 FILLER_11_324 ();
 sg13g2_fill_1 FILLER_11_326 ();
 sg13g2_decap_8 FILLER_11_331 ();
 sg13g2_decap_4 FILLER_11_343 ();
 sg13g2_fill_1 FILLER_11_347 ();
 sg13g2_decap_8 FILLER_11_352 ();
 sg13g2_decap_4 FILLER_11_359 ();
 sg13g2_decap_4 FILLER_11_389 ();
 sg13g2_fill_1 FILLER_11_393 ();
 sg13g2_decap_8 FILLER_11_398 ();
 sg13g2_decap_4 FILLER_11_405 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_fill_2 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_38 ();
 sg13g2_decap_8 FILLER_12_45 ();
 sg13g2_decap_4 FILLER_12_65 ();
 sg13g2_fill_1 FILLER_12_69 ();
 sg13g2_decap_8 FILLER_12_78 ();
 sg13g2_decap_8 FILLER_12_85 ();
 sg13g2_decap_8 FILLER_12_92 ();
 sg13g2_decap_8 FILLER_12_99 ();
 sg13g2_decap_8 FILLER_12_106 ();
 sg13g2_decap_8 FILLER_12_113 ();
 sg13g2_fill_2 FILLER_12_120 ();
 sg13g2_fill_1 FILLER_12_122 ();
 sg13g2_decap_8 FILLER_12_159 ();
 sg13g2_fill_2 FILLER_12_166 ();
 sg13g2_fill_1 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_fill_2 FILLER_12_189 ();
 sg13g2_fill_1 FILLER_12_191 ();
 sg13g2_decap_8 FILLER_12_223 ();
 sg13g2_fill_2 FILLER_12_230 ();
 sg13g2_decap_8 FILLER_12_236 ();
 sg13g2_decap_8 FILLER_12_243 ();
 sg13g2_fill_1 FILLER_12_250 ();
 sg13g2_decap_8 FILLER_12_255 ();
 sg13g2_decap_4 FILLER_12_262 ();
 sg13g2_fill_1 FILLER_12_292 ();
 sg13g2_fill_2 FILLER_12_298 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_fill_1 FILLER_12_315 ();
 sg13g2_fill_2 FILLER_12_372 ();
 sg13g2_decap_8 FILLER_12_381 ();
 sg13g2_decap_4 FILLER_12_388 ();
 sg13g2_fill_1 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_397 ();
 sg13g2_decap_4 FILLER_12_404 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_fill_2 FILLER_13_56 ();
 sg13g2_fill_1 FILLER_13_58 ();
 sg13g2_decap_8 FILLER_13_85 ();
 sg13g2_fill_1 FILLER_13_92 ();
 sg13g2_fill_2 FILLER_13_139 ();
 sg13g2_decap_4 FILLER_13_187 ();
 sg13g2_decap_4 FILLER_13_195 ();
 sg13g2_fill_1 FILLER_13_199 ();
 sg13g2_decap_4 FILLER_13_204 ();
 sg13g2_decap_8 FILLER_13_212 ();
 sg13g2_fill_2 FILLER_13_219 ();
 sg13g2_decap_8 FILLER_13_247 ();
 sg13g2_decap_8 FILLER_13_254 ();
 sg13g2_fill_2 FILLER_13_261 ();
 sg13g2_decap_4 FILLER_13_267 ();
 sg13g2_fill_1 FILLER_13_271 ();
 sg13g2_decap_8 FILLER_13_286 ();
 sg13g2_fill_2 FILLER_13_293 ();
 sg13g2_decap_4 FILLER_13_299 ();
 sg13g2_fill_1 FILLER_13_313 ();
 sg13g2_decap_4 FILLER_13_340 ();
 sg13g2_fill_1 FILLER_13_344 ();
 sg13g2_fill_2 FILLER_13_371 ();
 sg13g2_fill_2 FILLER_13_407 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_fill_2 FILLER_14_28 ();
 sg13g2_fill_1 FILLER_14_30 ();
 sg13g2_decap_8 FILLER_14_37 ();
 sg13g2_decap_8 FILLER_14_44 ();
 sg13g2_decap_8 FILLER_14_51 ();
 sg13g2_decap_8 FILLER_14_58 ();
 sg13g2_decap_8 FILLER_14_65 ();
 sg13g2_decap_8 FILLER_14_72 ();
 sg13g2_decap_8 FILLER_14_79 ();
 sg13g2_decap_4 FILLER_14_86 ();
 sg13g2_decap_8 FILLER_14_116 ();
 sg13g2_fill_1 FILLER_14_123 ();
 sg13g2_decap_4 FILLER_14_176 ();
 sg13g2_fill_1 FILLER_14_180 ();
 sg13g2_fill_2 FILLER_14_207 ();
 sg13g2_fill_2 FILLER_14_214 ();
 sg13g2_fill_1 FILLER_14_216 ();
 sg13g2_decap_4 FILLER_14_279 ();
 sg13g2_fill_2 FILLER_14_283 ();
 sg13g2_decap_4 FILLER_14_311 ();
 sg13g2_decap_8 FILLER_14_318 ();
 sg13g2_decap_4 FILLER_14_329 ();
 sg13g2_fill_2 FILLER_14_333 ();
 sg13g2_fill_1 FILLER_14_345 ();
 sg13g2_decap_8 FILLER_14_349 ();
 sg13g2_decap_8 FILLER_14_360 ();
 sg13g2_decap_8 FILLER_14_372 ();
 sg13g2_fill_2 FILLER_15_0 ();
 sg13g2_decap_4 FILLER_15_28 ();
 sg13g2_fill_2 FILLER_15_32 ();
 sg13g2_decap_8 FILLER_15_60 ();
 sg13g2_fill_1 FILLER_15_67 ();
 sg13g2_decap_8 FILLER_15_94 ();
 sg13g2_decap_8 FILLER_15_101 ();
 sg13g2_decap_8 FILLER_15_108 ();
 sg13g2_decap_8 FILLER_15_125 ();
 sg13g2_fill_1 FILLER_15_132 ();
 sg13g2_decap_8 FILLER_15_137 ();
 sg13g2_fill_2 FILLER_15_144 ();
 sg13g2_decap_4 FILLER_15_172 ();
 sg13g2_fill_1 FILLER_15_180 ();
 sg13g2_decap_8 FILLER_15_191 ();
 sg13g2_decap_4 FILLER_15_198 ();
 sg13g2_decap_8 FILLER_15_228 ();
 sg13g2_fill_2 FILLER_15_235 ();
 sg13g2_decap_4 FILLER_15_241 ();
 sg13g2_decap_8 FILLER_15_258 ();
 sg13g2_decap_4 FILLER_15_265 ();
 sg13g2_fill_2 FILLER_15_272 ();
 sg13g2_decap_8 FILLER_15_300 ();
 sg13g2_fill_1 FILLER_15_307 ();
 sg13g2_decap_4 FILLER_15_334 ();
 sg13g2_fill_1 FILLER_15_338 ();
 sg13g2_fill_1 FILLER_15_365 ();
 sg13g2_decap_8 FILLER_15_395 ();
 sg13g2_decap_8 FILLER_15_402 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_4 FILLER_16_14 ();
 sg13g2_fill_2 FILLER_16_18 ();
 sg13g2_decap_4 FILLER_16_46 ();
 sg13g2_fill_1 FILLER_16_50 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_fill_2 FILLER_16_110 ();
 sg13g2_decap_4 FILLER_16_148 ();
 sg13g2_decap_8 FILLER_16_221 ();
 sg13g2_fill_2 FILLER_16_228 ();
 sg13g2_decap_8 FILLER_16_308 ();
 sg13g2_decap_8 FILLER_16_341 ();
 sg13g2_fill_2 FILLER_16_348 ();
 sg13g2_fill_1 FILLER_16_376 ();
 sg13g2_decap_8 FILLER_16_381 ();
 sg13g2_decap_4 FILLER_16_388 ();
 sg13g2_fill_1 FILLER_16_392 ();
 sg13g2_decap_8 FILLER_16_398 ();
 sg13g2_decap_4 FILLER_16_405 ();
 sg13g2_decap_8 FILLER_17_26 ();
 sg13g2_decap_8 FILLER_17_33 ();
 sg13g2_fill_2 FILLER_17_40 ();
 sg13g2_fill_1 FILLER_17_42 ();
 sg13g2_decap_4 FILLER_17_51 ();
 sg13g2_decap_8 FILLER_17_81 ();
 sg13g2_decap_8 FILLER_17_88 ();
 sg13g2_decap_8 FILLER_17_131 ();
 sg13g2_fill_2 FILLER_17_138 ();
 sg13g2_decap_8 FILLER_17_150 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_fill_2 FILLER_17_168 ();
 sg13g2_fill_1 FILLER_17_170 ();
 sg13g2_decap_8 FILLER_17_181 ();
 sg13g2_decap_8 FILLER_17_188 ();
 sg13g2_decap_4 FILLER_17_195 ();
 sg13g2_decap_4 FILLER_17_203 ();
 sg13g2_fill_2 FILLER_17_207 ();
 sg13g2_decap_4 FILLER_17_235 ();
 sg13g2_fill_2 FILLER_17_239 ();
 sg13g2_decap_8 FILLER_17_245 ();
 sg13g2_decap_8 FILLER_17_252 ();
 sg13g2_fill_2 FILLER_17_272 ();
 sg13g2_decap_8 FILLER_17_279 ();
 sg13g2_fill_1 FILLER_17_286 ();
 sg13g2_fill_1 FILLER_17_294 ();
 sg13g2_decap_8 FILLER_17_311 ();
 sg13g2_decap_4 FILLER_17_318 ();
 sg13g2_decap_8 FILLER_17_329 ();
 sg13g2_fill_2 FILLER_17_336 ();
 sg13g2_fill_1 FILLER_17_338 ();
 sg13g2_fill_2 FILLER_17_358 ();
 sg13g2_fill_1 FILLER_17_360 ();
 sg13g2_decap_4 FILLER_17_365 ();
 sg13g2_decap_8 FILLER_17_372 ();
 sg13g2_decap_4 FILLER_17_379 ();
 sg13g2_fill_2 FILLER_17_383 ();
 sg13g2_fill_2 FILLER_17_407 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_4 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_44 ();
 sg13g2_decap_8 FILLER_18_51 ();
 sg13g2_decap_4 FILLER_18_58 ();
 sg13g2_fill_2 FILLER_18_62 ();
 sg13g2_decap_8 FILLER_18_99 ();
 sg13g2_fill_2 FILLER_18_106 ();
 sg13g2_fill_1 FILLER_18_108 ();
 sg13g2_fill_2 FILLER_18_117 ();
 sg13g2_fill_1 FILLER_18_119 ();
 sg13g2_decap_4 FILLER_18_172 ();
 sg13g2_fill_2 FILLER_18_202 ();
 sg13g2_fill_2 FILLER_18_230 ();
 sg13g2_fill_1 FILLER_18_232 ();
 sg13g2_fill_2 FILLER_18_246 ();
 sg13g2_fill_1 FILLER_18_248 ();
 sg13g2_fill_2 FILLER_18_265 ();
 sg13g2_fill_1 FILLER_18_267 ();
 sg13g2_fill_1 FILLER_18_276 ();
 sg13g2_fill_2 FILLER_18_311 ();
 sg13g2_fill_1 FILLER_18_313 ();
 sg13g2_decap_4 FILLER_18_347 ();
 sg13g2_fill_2 FILLER_18_351 ();
 sg13g2_fill_1 FILLER_18_361 ();
 sg13g2_fill_1 FILLER_18_388 ();
 sg13g2_decap_4 FILLER_18_405 ();
 sg13g2_fill_1 FILLER_19_35 ();
 sg13g2_decap_4 FILLER_19_62 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_4 FILLER_19_77 ();
 sg13g2_fill_2 FILLER_19_81 ();
 sg13g2_decap_4 FILLER_19_87 ();
 sg13g2_fill_1 FILLER_19_91 ();
 sg13g2_fill_1 FILLER_19_97 ();
 sg13g2_fill_1 FILLER_19_134 ();
 sg13g2_decap_4 FILLER_19_152 ();
 sg13g2_fill_1 FILLER_19_156 ();
 sg13g2_decap_4 FILLER_19_161 ();
 sg13g2_decap_8 FILLER_19_175 ();
 sg13g2_decap_8 FILLER_19_182 ();
 sg13g2_decap_8 FILLER_19_189 ();
 sg13g2_decap_8 FILLER_19_196 ();
 sg13g2_decap_4 FILLER_19_203 ();
 sg13g2_decap_4 FILLER_19_219 ();
 sg13g2_fill_1 FILLER_19_223 ();
 sg13g2_decap_8 FILLER_19_227 ();
 sg13g2_decap_8 FILLER_19_262 ();
 sg13g2_decap_8 FILLER_19_269 ();
 sg13g2_fill_2 FILLER_19_276 ();
 sg13g2_fill_1 FILLER_19_278 ();
 sg13g2_decap_4 FILLER_19_283 ();
 sg13g2_fill_2 FILLER_19_287 ();
 sg13g2_decap_4 FILLER_19_294 ();
 sg13g2_fill_2 FILLER_19_298 ();
 sg13g2_fill_2 FILLER_19_305 ();
 sg13g2_fill_1 FILLER_19_307 ();
 sg13g2_decap_8 FILLER_19_325 ();
 sg13g2_fill_1 FILLER_19_342 ();
 sg13g2_fill_2 FILLER_19_407 ();
 sg13g2_decap_4 FILLER_20_0 ();
 sg13g2_fill_1 FILLER_20_4 ();
 sg13g2_decap_8 FILLER_20_31 ();
 sg13g2_decap_8 FILLER_20_38 ();
 sg13g2_decap_8 FILLER_20_45 ();
 sg13g2_decap_4 FILLER_20_52 ();
 sg13g2_fill_2 FILLER_20_56 ();
 sg13g2_fill_2 FILLER_20_136 ();
 sg13g2_fill_1 FILLER_20_138 ();
 sg13g2_decap_4 FILLER_20_201 ();
 sg13g2_fill_1 FILLER_20_205 ();
 sg13g2_fill_1 FILLER_20_248 ();
 sg13g2_decap_4 FILLER_20_275 ();
 sg13g2_fill_2 FILLER_20_279 ();
 sg13g2_decap_4 FILLER_20_290 ();
 sg13g2_decap_4 FILLER_20_323 ();
 sg13g2_fill_2 FILLER_20_327 ();
 sg13g2_fill_2 FILLER_20_349 ();
 sg13g2_decap_4 FILLER_20_354 ();
 sg13g2_fill_1 FILLER_20_358 ();
 sg13g2_decap_8 FILLER_20_374 ();
 sg13g2_decap_8 FILLER_20_381 ();
 sg13g2_fill_1 FILLER_20_388 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_4 FILLER_21_14 ();
 sg13g2_fill_2 FILLER_21_18 ();
 sg13g2_decap_8 FILLER_21_75 ();
 sg13g2_decap_8 FILLER_21_82 ();
 sg13g2_fill_2 FILLER_21_89 ();
 sg13g2_fill_1 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_100 ();
 sg13g2_decap_4 FILLER_21_107 ();
 sg13g2_fill_1 FILLER_21_111 ();
 sg13g2_decap_8 FILLER_21_125 ();
 sg13g2_fill_2 FILLER_21_132 ();
 sg13g2_decap_4 FILLER_21_139 ();
 sg13g2_fill_2 FILLER_21_143 ();
 sg13g2_decap_4 FILLER_21_148 ();
 sg13g2_fill_1 FILLER_21_152 ();
 sg13g2_fill_2 FILLER_21_163 ();
 sg13g2_decap_4 FILLER_21_182 ();
 sg13g2_fill_2 FILLER_21_186 ();
 sg13g2_fill_1 FILLER_21_196 ();
 sg13g2_decap_8 FILLER_21_223 ();
 sg13g2_decap_8 FILLER_21_230 ();
 sg13g2_decap_4 FILLER_21_237 ();
 sg13g2_fill_2 FILLER_21_241 ();
 sg13g2_decap_8 FILLER_21_246 ();
 sg13g2_fill_2 FILLER_21_253 ();
 sg13g2_fill_1 FILLER_21_255 ();
 sg13g2_decap_8 FILLER_21_265 ();
 sg13g2_fill_1 FILLER_21_272 ();
 sg13g2_fill_2 FILLER_21_281 ();
 sg13g2_decap_8 FILLER_21_295 ();
 sg13g2_fill_2 FILLER_21_302 ();
 sg13g2_fill_1 FILLER_21_304 ();
 sg13g2_decap_4 FILLER_21_331 ();
 sg13g2_fill_2 FILLER_21_335 ();
 sg13g2_decap_8 FILLER_21_345 ();
 sg13g2_fill_2 FILLER_21_352 ();
 sg13g2_decap_8 FILLER_21_376 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_29 ();
 sg13g2_fill_2 FILLER_22_36 ();
 sg13g2_fill_1 FILLER_22_38 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_fill_2 FILLER_22_56 ();
 sg13g2_fill_1 FILLER_22_58 ();
 sg13g2_decap_8 FILLER_22_85 ();
 sg13g2_fill_1 FILLER_22_92 ();
 sg13g2_decap_4 FILLER_22_98 ();
 sg13g2_decap_8 FILLER_22_164 ();
 sg13g2_fill_2 FILLER_22_171 ();
 sg13g2_decap_8 FILLER_22_198 ();
 sg13g2_fill_2 FILLER_22_205 ();
 sg13g2_fill_1 FILLER_22_210 ();
 sg13g2_decap_4 FILLER_22_216 ();
 sg13g2_fill_2 FILLER_22_220 ();
 sg13g2_fill_1 FILLER_22_272 ();
 sg13g2_fill_2 FILLER_22_304 ();
 sg13g2_fill_1 FILLER_22_306 ();
 sg13g2_decap_8 FILLER_22_320 ();
 sg13g2_fill_1 FILLER_22_327 ();
 sg13g2_fill_2 FILLER_22_348 ();
 sg13g2_fill_1 FILLER_22_350 ();
 sg13g2_fill_2 FILLER_22_377 ();
 sg13g2_fill_1 FILLER_22_379 ();
 sg13g2_decap_4 FILLER_22_405 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_4 FILLER_23_14 ();
 sg13g2_fill_2 FILLER_23_18 ();
 sg13g2_decap_8 FILLER_23_72 ();
 sg13g2_fill_1 FILLER_23_79 ();
 sg13g2_fill_2 FILLER_23_107 ();
 sg13g2_fill_2 FILLER_23_112 ();
 sg13g2_decap_4 FILLER_23_135 ();
 sg13g2_fill_2 FILLER_23_139 ();
 sg13g2_decap_4 FILLER_23_179 ();
 sg13g2_fill_2 FILLER_23_183 ();
 sg13g2_fill_2 FILLER_23_201 ();
 sg13g2_fill_2 FILLER_23_208 ();
 sg13g2_fill_1 FILLER_23_210 ();
 sg13g2_fill_2 FILLER_23_239 ();
 sg13g2_fill_1 FILLER_23_241 ();
 sg13g2_fill_2 FILLER_23_255 ();
 sg13g2_fill_1 FILLER_23_257 ();
 sg13g2_fill_2 FILLER_23_266 ();
 sg13g2_fill_1 FILLER_23_268 ();
 sg13g2_fill_2 FILLER_23_277 ();
 sg13g2_fill_1 FILLER_23_289 ();
 sg13g2_fill_2 FILLER_23_301 ();
 sg13g2_fill_1 FILLER_23_303 ();
 sg13g2_decap_8 FILLER_23_322 ();
 sg13g2_decap_8 FILLER_23_329 ();
 sg13g2_decap_8 FILLER_23_366 ();
 sg13g2_decap_4 FILLER_23_373 ();
 sg13g2_fill_1 FILLER_23_395 ();
 sg13g2_decap_4 FILLER_23_404 ();
 sg13g2_fill_1 FILLER_23_408 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_4 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_4 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_50 ();
 sg13g2_decap_4 FILLER_24_61 ();
 sg13g2_fill_2 FILLER_24_65 ();
 sg13g2_decap_8 FILLER_24_101 ();
 sg13g2_fill_2 FILLER_24_108 ();
 sg13g2_fill_1 FILLER_24_110 ();
 sg13g2_decap_4 FILLER_24_124 ();
 sg13g2_decap_8 FILLER_24_168 ();
 sg13g2_decap_4 FILLER_24_175 ();
 sg13g2_fill_1 FILLER_24_179 ();
 sg13g2_fill_2 FILLER_24_188 ();
 sg13g2_fill_1 FILLER_24_190 ();
 sg13g2_fill_2 FILLER_24_205 ();
 sg13g2_fill_1 FILLER_24_220 ();
 sg13g2_decap_8 FILLER_24_246 ();
 sg13g2_fill_2 FILLER_24_313 ();
 sg13g2_decap_8 FILLER_24_341 ();
 sg13g2_decap_8 FILLER_24_348 ();
 sg13g2_decap_8 FILLER_24_355 ();
 sg13g2_decap_8 FILLER_24_362 ();
 sg13g2_fill_1 FILLER_24_369 ();
 sg13g2_fill_1 FILLER_24_377 ();
 sg13g2_decap_4 FILLER_24_404 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_decap_4 FILLER_25_0 ();
 sg13g2_fill_1 FILLER_25_61 ();
 sg13g2_decap_4 FILLER_25_82 ();
 sg13g2_fill_1 FILLER_25_86 ();
 sg13g2_decap_4 FILLER_25_113 ();
 sg13g2_fill_1 FILLER_25_117 ();
 sg13g2_fill_1 FILLER_25_126 ();
 sg13g2_decap_8 FILLER_25_144 ();
 sg13g2_fill_1 FILLER_25_151 ();
 sg13g2_decap_4 FILLER_25_178 ();
 sg13g2_fill_2 FILLER_25_182 ();
 sg13g2_decap_4 FILLER_25_197 ();
 sg13g2_fill_2 FILLER_25_201 ();
 sg13g2_decap_4 FILLER_25_234 ();
 sg13g2_decap_4 FILLER_25_246 ();
 sg13g2_fill_1 FILLER_25_250 ();
 sg13g2_decap_8 FILLER_25_281 ();
 sg13g2_decap_8 FILLER_25_288 ();
 sg13g2_decap_4 FILLER_25_295 ();
 sg13g2_fill_1 FILLER_25_299 ();
 sg13g2_decap_8 FILLER_25_319 ();
 sg13g2_fill_2 FILLER_25_326 ();
 sg13g2_fill_2 FILLER_25_380 ();
 sg13g2_fill_1 FILLER_25_382 ();
 sg13g2_decap_8 FILLER_26_40 ();
 sg13g2_decap_8 FILLER_26_51 ();
 sg13g2_decap_8 FILLER_26_58 ();
 sg13g2_fill_2 FILLER_26_65 ();
 sg13g2_fill_1 FILLER_26_71 ();
 sg13g2_decap_8 FILLER_26_85 ();
 sg13g2_fill_2 FILLER_26_92 ();
 sg13g2_fill_1 FILLER_26_94 ();
 sg13g2_decap_8 FILLER_26_101 ();
 sg13g2_decap_8 FILLER_26_108 ();
 sg13g2_fill_1 FILLER_26_115 ();
 sg13g2_decap_8 FILLER_26_137 ();
 sg13g2_decap_8 FILLER_26_144 ();
 sg13g2_decap_8 FILLER_26_151 ();
 sg13g2_decap_4 FILLER_26_158 ();
 sg13g2_fill_2 FILLER_26_162 ();
 sg13g2_decap_8 FILLER_26_167 ();
 sg13g2_fill_2 FILLER_26_174 ();
 sg13g2_fill_1 FILLER_26_176 ();
 sg13g2_decap_8 FILLER_26_201 ();
 sg13g2_decap_8 FILLER_26_208 ();
 sg13g2_decap_8 FILLER_26_215 ();
 sg13g2_decap_4 FILLER_26_222 ();
 sg13g2_fill_1 FILLER_26_226 ();
 sg13g2_fill_1 FILLER_26_244 ();
 sg13g2_decap_8 FILLER_26_249 ();
 sg13g2_decap_4 FILLER_26_256 ();
 sg13g2_fill_2 FILLER_26_260 ();
 sg13g2_decap_8 FILLER_26_266 ();
 sg13g2_fill_1 FILLER_26_273 ();
 sg13g2_decap_4 FILLER_26_279 ();
 sg13g2_fill_2 FILLER_26_283 ();
 sg13g2_decap_8 FILLER_26_340 ();
 sg13g2_fill_2 FILLER_26_347 ();
 sg13g2_decap_4 FILLER_26_354 ();
 sg13g2_fill_1 FILLER_26_358 ();
 sg13g2_fill_2 FILLER_26_368 ();
 sg13g2_decap_4 FILLER_26_380 ();
 sg13g2_fill_2 FILLER_26_407 ();
 sg13g2_decap_4 FILLER_27_0 ();
 sg13g2_fill_2 FILLER_27_4 ();
 sg13g2_fill_2 FILLER_27_20 ();
 sg13g2_decap_8 FILLER_27_25 ();
 sg13g2_decap_4 FILLER_27_32 ();
 sg13g2_fill_2 FILLER_27_62 ();
 sg13g2_decap_4 FILLER_27_198 ();
 sg13g2_fill_2 FILLER_27_228 ();
 sg13g2_fill_1 FILLER_27_260 ();
 sg13g2_fill_2 FILLER_27_275 ();
 sg13g2_fill_2 FILLER_27_289 ();
 sg13g2_fill_1 FILLER_27_291 ();
 sg13g2_fill_1 FILLER_27_332 ();
 sg13g2_decap_4 FILLER_27_364 ();
 sg13g2_fill_1 FILLER_28_0 ();
 sg13g2_fill_2 FILLER_28_61 ();
 sg13g2_fill_1 FILLER_28_63 ();
 sg13g2_fill_1 FILLER_28_78 ();
 sg13g2_decap_8 FILLER_28_87 ();
 sg13g2_decap_8 FILLER_28_94 ();
 sg13g2_fill_1 FILLER_28_101 ();
 sg13g2_decap_8 FILLER_28_107 ();
 sg13g2_decap_4 FILLER_28_114 ();
 sg13g2_decap_8 FILLER_28_131 ();
 sg13g2_decap_8 FILLER_28_138 ();
 sg13g2_decap_4 FILLER_28_145 ();
 sg13g2_decap_8 FILLER_28_159 ();
 sg13g2_decap_8 FILLER_28_166 ();
 sg13g2_decap_4 FILLER_28_173 ();
 sg13g2_fill_2 FILLER_28_177 ();
 sg13g2_fill_2 FILLER_28_210 ();
 sg13g2_fill_1 FILLER_28_212 ();
 sg13g2_fill_2 FILLER_28_217 ();
 sg13g2_fill_2 FILLER_28_223 ();
 sg13g2_decap_4 FILLER_28_247 ();
 sg13g2_fill_1 FILLER_28_277 ();
 sg13g2_fill_2 FILLER_28_287 ();
 sg13g2_decap_4 FILLER_28_364 ();
 sg13g2_fill_2 FILLER_28_368 ();
 sg13g2_fill_1 FILLER_28_380 ();
 sg13g2_fill_1 FILLER_28_408 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_fill_1 FILLER_29_19 ();
 sg13g2_decap_8 FILLER_29_29 ();
 sg13g2_decap_8 FILLER_29_36 ();
 sg13g2_fill_2 FILLER_29_43 ();
 sg13g2_fill_1 FILLER_29_45 ();
 sg13g2_decap_8 FILLER_29_50 ();
 sg13g2_decap_4 FILLER_29_57 ();
 sg13g2_fill_2 FILLER_29_61 ();
 sg13g2_fill_2 FILLER_29_93 ();
 sg13g2_fill_1 FILLER_29_95 ();
 sg13g2_decap_8 FILLER_29_101 ();
 sg13g2_decap_8 FILLER_29_108 ();
 sg13g2_fill_1 FILLER_29_115 ();
 sg13g2_fill_1 FILLER_29_136 ();
 sg13g2_fill_2 FILLER_29_163 ();
 sg13g2_decap_8 FILLER_29_168 ();
 sg13g2_decap_8 FILLER_29_175 ();
 sg13g2_fill_2 FILLER_29_182 ();
 sg13g2_fill_2 FILLER_29_196 ();
 sg13g2_decap_8 FILLER_29_212 ();
 sg13g2_decap_4 FILLER_29_219 ();
 sg13g2_fill_2 FILLER_29_252 ();
 sg13g2_fill_1 FILLER_29_254 ();
 sg13g2_decap_8 FILLER_29_281 ();
 sg13g2_decap_4 FILLER_29_288 ();
 sg13g2_fill_1 FILLER_29_292 ();
 sg13g2_fill_1 FILLER_29_324 ();
 sg13g2_fill_2 FILLER_29_351 ();
 sg13g2_decap_8 FILLER_29_368 ();
 sg13g2_decap_4 FILLER_29_405 ();
 sg13g2_decap_4 FILLER_30_0 ();
 sg13g2_fill_1 FILLER_30_4 ();
 sg13g2_fill_2 FILLER_30_36 ();
 sg13g2_fill_2 FILLER_30_64 ();
 sg13g2_fill_1 FILLER_30_66 ();
 sg13g2_fill_2 FILLER_30_87 ();
 sg13g2_fill_2 FILLER_30_115 ();
 sg13g2_fill_1 FILLER_30_117 ();
 sg13g2_decap_8 FILLER_30_144 ();
 sg13g2_decap_4 FILLER_30_151 ();
 sg13g2_fill_2 FILLER_30_155 ();
 sg13g2_fill_2 FILLER_30_183 ();
 sg13g2_fill_1 FILLER_30_193 ();
 sg13g2_fill_2 FILLER_30_230 ();
 sg13g2_fill_1 FILLER_30_232 ();
 sg13g2_decap_4 FILLER_30_246 ();
 sg13g2_fill_1 FILLER_30_250 ();
 sg13g2_fill_2 FILLER_30_266 ();
 sg13g2_fill_1 FILLER_30_268 ();
 sg13g2_decap_8 FILLER_30_303 ();
 sg13g2_fill_2 FILLER_30_310 ();
 sg13g2_decap_8 FILLER_30_330 ();
 sg13g2_decap_8 FILLER_30_337 ();
 sg13g2_fill_2 FILLER_30_344 ();
 sg13g2_fill_1 FILLER_30_346 ();
 sg13g2_fill_2 FILLER_31_0 ();
 sg13g2_fill_1 FILLER_31_2 ();
 sg13g2_decap_8 FILLER_31_37 ();
 sg13g2_decap_4 FILLER_31_44 ();
 sg13g2_fill_1 FILLER_31_48 ();
 sg13g2_decap_8 FILLER_31_53 ();
 sg13g2_decap_8 FILLER_31_60 ();
 sg13g2_decap_8 FILLER_31_87 ();
 sg13g2_fill_2 FILLER_31_94 ();
 sg13g2_fill_1 FILLER_31_96 ();
 sg13g2_decap_8 FILLER_31_103 ();
 sg13g2_decap_4 FILLER_31_110 ();
 sg13g2_fill_1 FILLER_31_128 ();
 sg13g2_fill_2 FILLER_31_137 ();
 sg13g2_decap_4 FILLER_31_165 ();
 sg13g2_fill_1 FILLER_31_169 ();
 sg13g2_decap_8 FILLER_31_173 ();
 sg13g2_decap_4 FILLER_31_180 ();
 sg13g2_fill_2 FILLER_31_184 ();
 sg13g2_fill_1 FILLER_31_198 ();
 sg13g2_fill_2 FILLER_31_217 ();
 sg13g2_fill_1 FILLER_31_228 ();
 sg13g2_fill_2 FILLER_31_245 ();
 sg13g2_fill_1 FILLER_31_247 ();
 sg13g2_fill_1 FILLER_31_257 ();
 sg13g2_fill_1 FILLER_31_263 ();
 sg13g2_fill_2 FILLER_31_274 ();
 sg13g2_fill_1 FILLER_31_276 ();
 sg13g2_decap_8 FILLER_31_290 ();
 sg13g2_fill_2 FILLER_31_297 ();
 sg13g2_fill_1 FILLER_31_299 ();
 sg13g2_fill_1 FILLER_31_303 ();
 sg13g2_fill_2 FILLER_31_313 ();
 sg13g2_fill_2 FILLER_31_327 ();
 sg13g2_fill_1 FILLER_31_373 ();
 sg13g2_decap_4 FILLER_31_384 ();
 sg13g2_fill_2 FILLER_31_388 ();
 sg13g2_decap_8 FILLER_31_398 ();
 sg13g2_decap_4 FILLER_31_405 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_fill_1 FILLER_32_7 ();
 sg13g2_fill_2 FILLER_32_19 ();
 sg13g2_fill_1 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_25 ();
 sg13g2_decap_8 FILLER_32_32 ();
 sg13g2_fill_1 FILLER_32_39 ();
 sg13g2_decap_4 FILLER_32_66 ();
 sg13g2_fill_2 FILLER_32_70 ();
 sg13g2_fill_2 FILLER_32_116 ();
 sg13g2_decap_8 FILLER_32_130 ();
 sg13g2_decap_8 FILLER_32_137 ();
 sg13g2_decap_8 FILLER_32_144 ();
 sg13g2_fill_2 FILLER_32_151 ();
 sg13g2_fill_1 FILLER_32_153 ();
 sg13g2_fill_2 FILLER_32_188 ();
 sg13g2_decap_8 FILLER_32_216 ();
 sg13g2_fill_2 FILLER_32_246 ();
 sg13g2_fill_1 FILLER_32_248 ();
 sg13g2_decap_4 FILLER_32_267 ();
 sg13g2_fill_2 FILLER_32_276 ();
 sg13g2_decap_4 FILLER_32_283 ();
 sg13g2_fill_1 FILLER_32_291 ();
 sg13g2_fill_1 FILLER_32_325 ();
 sg13g2_decap_8 FILLER_32_331 ();
 sg13g2_decap_8 FILLER_32_358 ();
 sg13g2_decap_8 FILLER_32_365 ();
 sg13g2_decap_8 FILLER_32_372 ();
 sg13g2_decap_4 FILLER_32_379 ();
 sg13g2_fill_2 FILLER_33_0 ();
 sg13g2_fill_1 FILLER_33_13 ();
 sg13g2_fill_2 FILLER_33_40 ();
 sg13g2_fill_1 FILLER_33_42 ();
 sg13g2_fill_2 FILLER_33_48 ();
 sg13g2_fill_1 FILLER_33_50 ();
 sg13g2_decap_8 FILLER_33_55 ();
 sg13g2_fill_1 FILLER_33_62 ();
 sg13g2_fill_2 FILLER_33_87 ();
 sg13g2_fill_1 FILLER_33_89 ();
 sg13g2_decap_4 FILLER_33_116 ();
 sg13g2_fill_1 FILLER_33_120 ();
 sg13g2_fill_1 FILLER_33_155 ();
 sg13g2_fill_2 FILLER_33_172 ();
 sg13g2_fill_1 FILLER_33_174 ();
 sg13g2_decap_4 FILLER_33_178 ();
 sg13g2_decap_8 FILLER_33_186 ();
 sg13g2_decap_4 FILLER_33_193 ();
 sg13g2_decap_8 FILLER_33_206 ();
 sg13g2_decap_4 FILLER_33_213 ();
 sg13g2_decap_4 FILLER_33_221 ();
 sg13g2_decap_4 FILLER_33_233 ();
 sg13g2_fill_1 FILLER_33_237 ();
 sg13g2_fill_1 FILLER_33_259 ();
 sg13g2_fill_2 FILLER_33_315 ();
 sg13g2_fill_1 FILLER_33_317 ();
 sg13g2_decap_4 FILLER_33_344 ();
 sg13g2_fill_1 FILLER_33_374 ();
 sg13g2_decap_8 FILLER_33_385 ();
 sg13g2_fill_1 FILLER_33_392 ();
 sg13g2_decap_8 FILLER_33_401 ();
 sg13g2_fill_1 FILLER_33_408 ();
 sg13g2_fill_1 FILLER_34_0 ();
 sg13g2_fill_1 FILLER_34_35 ();
 sg13g2_fill_1 FILLER_34_62 ();
 sg13g2_decap_8 FILLER_34_90 ();
 sg13g2_fill_2 FILLER_34_97 ();
 sg13g2_decap_8 FILLER_34_105 ();
 sg13g2_decap_4 FILLER_34_112 ();
 sg13g2_fill_2 FILLER_34_116 ();
 sg13g2_decap_8 FILLER_34_135 ();
 sg13g2_decap_8 FILLER_34_142 ();
 sg13g2_decap_4 FILLER_34_149 ();
 sg13g2_decap_8 FILLER_34_197 ();
 sg13g2_decap_8 FILLER_34_204 ();
 sg13g2_decap_4 FILLER_34_211 ();
 sg13g2_fill_2 FILLER_34_241 ();
 sg13g2_fill_1 FILLER_34_243 ();
 sg13g2_decap_8 FILLER_34_288 ();
 sg13g2_decap_8 FILLER_34_295 ();
 sg13g2_decap_8 FILLER_34_302 ();
 sg13g2_decap_8 FILLER_34_319 ();
 sg13g2_decap_8 FILLER_34_326 ();
 sg13g2_decap_4 FILLER_34_333 ();
 sg13g2_fill_2 FILLER_34_337 ();
 sg13g2_decap_8 FILLER_34_375 ();
 sg13g2_fill_1 FILLER_34_382 ();
 sg13g2_decap_4 FILLER_35_0 ();
 sg13g2_fill_1 FILLER_35_4 ();
 sg13g2_decap_8 FILLER_35_23 ();
 sg13g2_fill_1 FILLER_35_30 ();
 sg13g2_decap_4 FILLER_35_61 ();
 sg13g2_fill_2 FILLER_35_65 ();
 sg13g2_decap_4 FILLER_35_71 ();
 sg13g2_fill_1 FILLER_35_79 ();
 sg13g2_decap_4 FILLER_35_177 ();
 sg13g2_decap_8 FILLER_35_233 ();
 sg13g2_fill_1 FILLER_35_240 ();
 sg13g2_decap_8 FILLER_35_331 ();
 sg13g2_fill_1 FILLER_35_338 ();
 sg13g2_decap_8 FILLER_35_375 ();
 sg13g2_fill_1 FILLER_35_382 ();
 sg13g2_decap_4 FILLER_36_0 ();
 sg13g2_fill_2 FILLER_36_4 ();
 sg13g2_decap_8 FILLER_36_32 ();
 sg13g2_fill_2 FILLER_36_39 ();
 sg13g2_decap_4 FILLER_36_67 ();
 sg13g2_fill_2 FILLER_36_71 ();
 sg13g2_fill_2 FILLER_36_94 ();
 sg13g2_fill_1 FILLER_36_96 ();
 sg13g2_fill_1 FILLER_36_102 ();
 sg13g2_decap_4 FILLER_36_111 ();
 sg13g2_decap_4 FILLER_36_133 ();
 sg13g2_decap_8 FILLER_36_140 ();
 sg13g2_decap_8 FILLER_36_147 ();
 sg13g2_fill_1 FILLER_36_154 ();
 sg13g2_fill_2 FILLER_36_167 ();
 sg13g2_fill_2 FILLER_36_195 ();
 sg13g2_fill_1 FILLER_36_197 ();
 sg13g2_decap_8 FILLER_36_206 ();
 sg13g2_fill_2 FILLER_36_213 ();
 sg13g2_fill_1 FILLER_36_215 ();
 sg13g2_decap_8 FILLER_36_220 ();
 sg13g2_decap_4 FILLER_36_227 ();
 sg13g2_fill_1 FILLER_36_231 ();
 sg13g2_fill_1 FILLER_36_236 ();
 sg13g2_fill_2 FILLER_36_260 ();
 sg13g2_fill_1 FILLER_36_262 ();
 sg13g2_fill_2 FILLER_36_282 ();
 sg13g2_fill_2 FILLER_36_310 ();
 sg13g2_decap_8 FILLER_36_338 ();
 sg13g2_fill_1 FILLER_36_345 ();
 sg13g2_fill_2 FILLER_36_372 ();
 sg13g2_fill_1 FILLER_36_374 ();
 sg13g2_decap_8 FILLER_36_399 ();
 sg13g2_fill_2 FILLER_36_406 ();
 sg13g2_fill_1 FILLER_36_408 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_fill_2 FILLER_37_14 ();
 sg13g2_fill_1 FILLER_37_16 ();
 sg13g2_decap_8 FILLER_37_20 ();
 sg13g2_decap_8 FILLER_37_27 ();
 sg13g2_decap_8 FILLER_37_34 ();
 sg13g2_fill_1 FILLER_37_41 ();
 sg13g2_fill_2 FILLER_37_46 ();
 sg13g2_fill_1 FILLER_37_48 ();
 sg13g2_fill_1 FILLER_37_92 ();
 sg13g2_decap_8 FILLER_37_119 ();
 sg13g2_fill_2 FILLER_37_126 ();
 sg13g2_fill_1 FILLER_37_128 ();
 sg13g2_fill_2 FILLER_37_155 ();
 sg13g2_fill_1 FILLER_37_173 ();
 sg13g2_fill_1 FILLER_37_220 ();
 sg13g2_decap_4 FILLER_37_251 ();
 sg13g2_fill_1 FILLER_37_255 ();
 sg13g2_decap_8 FILLER_37_295 ();
 sg13g2_fill_2 FILLER_37_302 ();
 sg13g2_fill_1 FILLER_37_304 ();
 sg13g2_fill_1 FILLER_37_324 ();
 sg13g2_decap_8 FILLER_37_345 ();
 sg13g2_decap_8 FILLER_37_352 ();
 sg13g2_decap_4 FILLER_37_363 ();
 sg13g2_fill_1 FILLER_37_367 ();
 sg13g2_decap_4 FILLER_37_404 ();
 sg13g2_fill_1 FILLER_37_408 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_4 FILLER_38_42 ();
 sg13g2_fill_2 FILLER_38_46 ();
 sg13g2_fill_1 FILLER_38_74 ();
 sg13g2_fill_2 FILLER_38_93 ();
 sg13g2_fill_1 FILLER_38_95 ();
 sg13g2_decap_4 FILLER_38_108 ();
 sg13g2_decap_4 FILLER_38_116 ();
 sg13g2_decap_4 FILLER_38_124 ();
 sg13g2_decap_4 FILLER_38_132 ();
 sg13g2_fill_1 FILLER_38_196 ();
 sg13g2_fill_2 FILLER_38_245 ();
 sg13g2_decap_8 FILLER_38_260 ();
 sg13g2_fill_2 FILLER_38_310 ();
 sg13g2_fill_1 FILLER_38_312 ();
 sg13g2_decap_4 FILLER_38_343 ();
 sg13g2_fill_1 FILLER_38_347 ();
 sg13g2_decap_8 FILLER_38_378 ();
 sg13g2_decap_4 FILLER_38_385 ();
 sg13g2_decap_8 FILLER_38_393 ();
 sg13g2_decap_8 FILLER_38_400 ();
 sg13g2_fill_2 FILLER_38_407 ();
 assign uio_oe[0] = net4;
 assign uio_oe[1] = net5;
 assign uio_oe[2] = net6;
 assign uio_oe[3] = net7;
 assign uio_oe[4] = net8;
 assign uio_oe[5] = net9;
 assign uio_oe[6] = net10;
 assign uio_oe[7] = net11;
 assign uio_out[0] = net12;
 assign uio_out[1] = net13;
 assign uio_out[2] = net14;
 assign uio_out[3] = net15;
 assign uio_out[4] = net16;
 assign uio_out[5] = net17;
 assign uio_out[6] = net18;
 assign uio_out[7] = net19;
 assign uo_out[0] = net20;
 assign uo_out[1] = net21;
 assign uo_out[2] = net22;
 assign uo_out[3] = net23;
 assign uo_out[4] = net24;
 assign uo_out[5] = net25;
 assign uo_out[6] = net26;
endmodule

module tt_um_mroblesh (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire net49;
 wire net48;
 wire _011_;
 wire net47;
 wire net46;
 wire net45;
 wire net44;
 wire net43;
 wire net42;
 wire net41;
 wire net40;
 wire net39;
 wire net38;
 wire _022_;
 wire net37;
 wire net36;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire net35;
 wire net34;
 wire net33;
 wire net32;
 wire net31;
 wire net30;
 wire net29;
 wire net28;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire _297_;
 wire _298_;
 wire _299_;
 wire _300_;
 wire _301_;
 wire _302_;
 wire _303_;
 wire _304_;
 wire _305_;
 wire _306_;
 wire _307_;
 wire _308_;
 wire _309_;
 wire _310_;
 wire _311_;
 wire _312_;
 wire _313_;
 wire _314_;
 wire _315_;
 wire _316_;
 wire _317_;
 wire _318_;
 wire _319_;
 wire _320_;
 wire _321_;
 wire _322_;
 wire _323_;
 wire _324_;
 wire _325_;
 wire _326_;
 wire _327_;
 wire _328_;
 wire _329_;
 wire _330_;
 wire _331_;
 wire _332_;
 wire _333_;
 wire _334_;
 wire _335_;
 wire _336_;
 wire _337_;
 wire _338_;
 wire _339_;
 wire _340_;
 wire _341_;
 wire _342_;
 wire _343_;
 wire _344_;
 wire _345_;
 wire _346_;
 wire _347_;
 wire _348_;
 wire _349_;
 wire _350_;
 wire _351_;
 wire _352_;
 wire _353_;
 wire _354_;
 wire _355_;
 wire _356_;
 wire _357_;
 wire _358_;
 wire _359_;
 wire _360_;
 wire _361_;
 wire _362_;
 wire _363_;
 wire _364_;
 wire _365_;
 wire _366_;
 wire _367_;
 wire _368_;
 wire _369_;
 wire _370_;
 wire _371_;
 wire _372_;
 wire _373_;
 wire _374_;
 wire _375_;
 wire _376_;
 wire _377_;
 wire _378_;
 wire _379_;
 wire _380_;
 wire _381_;
 wire _382_;
 wire _383_;
 wire _384_;
 wire _385_;
 wire _386_;
 wire _387_;
 wire _388_;
 wire _389_;
 wire _390_;
 wire _391_;
 wire _392_;
 wire _393_;
 wire _394_;
 wire _395_;
 wire _396_;
 wire _397_;
 wire _398_;
 wire _399_;
 wire _400_;
 wire _401_;
 wire _402_;
 wire _403_;
 wire _404_;
 wire _405_;
 wire _406_;
 wire _407_;
 wire _408_;
 wire _409_;
 wire _410_;
 wire _411_;
 wire _412_;
 wire _413_;
 wire _414_;
 wire _415_;
 wire _416_;
 wire _417_;
 wire _418_;
 wire _419_;
 wire _420_;
 wire _421_;
 wire _422_;
 wire _423_;
 wire _424_;
 wire _425_;
 wire _426_;
 wire _427_;
 wire _428_;
 wire _429_;
 wire _430_;
 wire _431_;
 wire _432_;
 wire _433_;
 wire _434_;
 wire _435_;
 wire _436_;
 wire _437_;
 wire _438_;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire clknet_0_clk;
 wire \decoder_inst.counter[0] ;
 wire \decoder_inst.counter[10] ;
 wire \decoder_inst.counter[11] ;
 wire \decoder_inst.counter[12] ;
 wire \decoder_inst.counter[13] ;
 wire \decoder_inst.counter[14] ;
 wire \decoder_inst.counter[15] ;
 wire \decoder_inst.counter[16] ;
 wire \decoder_inst.counter[17] ;
 wire \decoder_inst.counter[18] ;
 wire \decoder_inst.counter[19] ;
 wire \decoder_inst.counter[1] ;
 wire \decoder_inst.counter[20] ;
 wire \decoder_inst.counter[21] ;
 wire \decoder_inst.counter[22] ;
 wire \decoder_inst.counter[23] ;
 wire \decoder_inst.counter[24] ;
 wire \decoder_inst.counter[25] ;
 wire \decoder_inst.counter[26] ;
 wire \decoder_inst.counter[27] ;
 wire \decoder_inst.counter[28] ;
 wire \decoder_inst.counter[29] ;
 wire \decoder_inst.counter[2] ;
 wire \decoder_inst.counter[30] ;
 wire \decoder_inst.counter[31] ;
 wire \decoder_inst.counter[3] ;
 wire \decoder_inst.counter[4] ;
 wire \decoder_inst.counter[5] ;
 wire \decoder_inst.counter[6] ;
 wire \decoder_inst.counter[7] ;
 wire \decoder_inst.counter[8] ;
 wire \decoder_inst.counter[9] ;
 wire \decoder_inst.freq_out[0] ;
 wire \decoder_inst.freq_out[1] ;
 wire \decoder_inst.freq_out[2] ;
 wire \decoder_inst.freq_out[3] ;
 wire \decoder_inst.freq_out[4] ;
 wire \decoder_inst.freq_out[5] ;
 wire \decoder_inst.freq_out[6] ;
 wire \decoder_inst.freq_out[7] ;
 wire \decoder_inst.frequency[0] ;
 wire \decoder_inst.frequency[10] ;
 wire \decoder_inst.frequency[11] ;
 wire \decoder_inst.frequency[12] ;
 wire \decoder_inst.frequency[13] ;
 wire \decoder_inst.frequency[14] ;
 wire \decoder_inst.frequency[15] ;
 wire \decoder_inst.frequency[16] ;
 wire \decoder_inst.frequency[17] ;
 wire \decoder_inst.frequency[18] ;
 wire \decoder_inst.frequency[19] ;
 wire \decoder_inst.frequency[1] ;
 wire \decoder_inst.frequency[20] ;
 wire \decoder_inst.frequency[21] ;
 wire \decoder_inst.frequency[22] ;
 wire \decoder_inst.frequency[23] ;
 wire \decoder_inst.frequency[24] ;
 wire \decoder_inst.frequency[25] ;
 wire \decoder_inst.frequency[26] ;
 wire \decoder_inst.frequency[27] ;
 wire \decoder_inst.frequency[28] ;
 wire \decoder_inst.frequency[29] ;
 wire \decoder_inst.frequency[2] ;
 wire \decoder_inst.frequency[30] ;
 wire \decoder_inst.frequency[31] ;
 wire \decoder_inst.frequency[3] ;
 wire \decoder_inst.frequency[4] ;
 wire \decoder_inst.frequency[5] ;
 wire \decoder_inst.frequency[6] ;
 wire \decoder_inst.frequency[7] ;
 wire \decoder_inst.frequency[8] ;
 wire \decoder_inst.frequency[9] ;
 wire \decoder_inst.signal_in_prev ;
 wire \encoder_inst.counter[0] ;
 wire \encoder_inst.counter[10] ;
 wire \encoder_inst.counter[11] ;
 wire \encoder_inst.counter[12] ;
 wire \encoder_inst.counter[13] ;
 wire \encoder_inst.counter[14] ;
 wire \encoder_inst.counter[15] ;
 wire \encoder_inst.counter[1] ;
 wire \encoder_inst.counter[2] ;
 wire \encoder_inst.counter[3] ;
 wire \encoder_inst.counter[4] ;
 wire \encoder_inst.counter[5] ;
 wire \encoder_inst.counter[6] ;
 wire \encoder_inst.counter[7] ;
 wire \encoder_inst.counter[8] ;
 wire \encoder_inst.counter[9] ;
 wire \encoder_inst.divide_value[0] ;
 wire \encoder_inst.divide_value[1] ;
 wire \encoder_inst.divide_value[2] ;
 wire \encoder_inst.divide_value[3] ;
 wire \encoder_inst.divide_value[4] ;
 wire \encoder_inst.divide_value[5] ;
 wire \encoder_inst.divide_value[6] ;
 wire \encoder_inst.divide_value[7] ;
 wire \encoder_inst.out ;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;

 sg13g2_inv_1 _465_ (.Y(_109_),
    .A(\encoder_inst.out ));
 sg13g2_inv_1 _466_ (.Y(_110_),
    .A(\encoder_inst.counter[0] ));
 sg13g2_inv_1 _467_ (.Y(_111_),
    .A(\decoder_inst.counter[7] ));
 sg13g2_inv_1 _468_ (.Y(_112_),
    .A(\decoder_inst.counter[6] ));
 sg13g2_inv_1 _469_ (.Y(_113_),
    .A(\encoder_inst.divide_value[1] ));
 sg13g2_inv_1 _470_ (.Y(_114_),
    .A(\encoder_inst.counter[1] ));
 sg13g2_inv_1 _471_ (.Y(_115_),
    .A(\encoder_inst.counter[3] ));
 sg13g2_inv_1 _472_ (.Y(_116_),
    .A(\encoder_inst.counter[2] ));
 sg13g2_inv_1 _473_ (.Y(_117_),
    .A(net241));
 sg13g2_inv_1 _474_ (.Y(_118_),
    .A(\encoder_inst.divide_value[6] ));
 sg13g2_inv_1 _475_ (.Y(_119_),
    .A(net247));
 sg13g2_inv_1 _476_ (.Y(_120_),
    .A(\encoder_inst.divide_value[5] ));
 sg13g2_inv_2 _477_ (.Y(_121_),
    .A(net116));
 sg13g2_inv_1 _478_ (.Y(_122_),
    .A(net188));
 sg13g2_inv_1 _479_ (.Y(_123_),
    .A(net163));
 sg13g2_inv_1 _480_ (.Y(_124_),
    .A(net249));
 sg13g2_inv_1 _481_ (.Y(_125_),
    .A(net191));
 sg13g2_inv_1 _482_ (.Y(_126_),
    .A(\decoder_inst.frequency[14] ));
 sg13g2_inv_1 _483_ (.Y(_127_),
    .A(net151));
 sg13g2_inv_1 _484_ (.Y(_128_),
    .A(net157));
 sg13g2_inv_1 _485_ (.Y(_129_),
    .A(net173));
 sg13g2_inv_1 _486_ (.Y(_130_),
    .A(net207));
 sg13g2_inv_1 _487_ (.Y(_131_),
    .A(net197));
 sg13g2_inv_1 _488_ (.Y(_132_),
    .A(net170));
 sg13g2_inv_1 _489_ (.Y(_133_),
    .A(net147));
 sg13g2_inv_1 _490_ (.Y(_134_),
    .A(net134));
 sg13g2_inv_1 _491_ (.Y(_135_),
    .A(net235));
 sg13g2_nor2_1 _492_ (.A(net100),
    .B(\decoder_inst.freq_out[0] ),
    .Y(_136_));
 sg13g2_a21oi_1 _493_ (.A1(_109_),
    .A2(net99),
    .Y(uo_out[0]),
    .B1(_136_));
 sg13g2_nor2b_1 _494_ (.A(net100),
    .B_N(\decoder_inst.freq_out[1] ),
    .Y(uo_out[1]));
 sg13g2_nor2b_1 _495_ (.A(net99),
    .B_N(\decoder_inst.freq_out[2] ),
    .Y(uo_out[2]));
 sg13g2_nor2b_1 _496_ (.A(net99),
    .B_N(\decoder_inst.freq_out[3] ),
    .Y(uo_out[3]));
 sg13g2_nor2b_1 _497_ (.A(net99),
    .B_N(\decoder_inst.freq_out[4] ),
    .Y(uo_out[4]));
 sg13g2_nor2b_1 _498_ (.A(net99),
    .B_N(\decoder_inst.freq_out[5] ),
    .Y(uo_out[5]));
 sg13g2_nor2b_1 _499_ (.A(net99),
    .B_N(\decoder_inst.freq_out[6] ),
    .Y(uo_out[6]));
 sg13g2_nor2b_1 _500_ (.A(net99),
    .B_N(\decoder_inst.freq_out[7] ),
    .Y(uo_out[7]));
 sg13g2_nor2b_2 _501_ (.A(net100),
    .B_N(net10),
    .Y(_137_));
 sg13g2_nand2b_2 _502_ (.Y(_138_),
    .B(net10),
    .A_N(net99));
 sg13g2_nand2b_2 _503_ (.Y(_139_),
    .B(net9),
    .A_N(net100));
 sg13g2_nand2_2 _504_ (.Y(_140_),
    .A(_138_),
    .B(_139_));
 sg13g2_o21ai_1 _505_ (.B1(_033_),
    .Y(_141_),
    .A1(\decoder_inst.counter[16] ),
    .A2(_140_));
 sg13g2_nor2_1 _506_ (.A(\decoder_inst.counter[15] ),
    .B(_140_),
    .Y(_142_));
 sg13g2_o21ai_1 _507_ (.B1(_140_),
    .Y(_143_),
    .A1(\decoder_inst.counter[16] ),
    .A2(\decoder_inst.counter[15] ));
 sg13g2_nor2_1 _508_ (.A(\decoder_inst.counter[14] ),
    .B(_142_),
    .Y(_144_));
 sg13g2_nand3b_1 _509_ (.B(_143_),
    .C(_144_),
    .Y(_145_),
    .A_N(_141_));
 sg13g2_nor2_1 _510_ (.A(net10),
    .B(_139_),
    .Y(_146_));
 sg13g2_nor3_1 _511_ (.A(net10),
    .B(\decoder_inst.counter[13] ),
    .C(_139_),
    .Y(_147_));
 sg13g2_nor2b_1 _512_ (.A(_146_),
    .B_N(\decoder_inst.counter[13] ),
    .Y(_148_));
 sg13g2_or3_1 _513_ (.A(\decoder_inst.counter[12] ),
    .B(_147_),
    .C(_148_),
    .X(_149_));
 sg13g2_a21oi_1 _514_ (.A1(_036_),
    .A2(_138_),
    .Y(_150_),
    .B1(\decoder_inst.counter[11] ));
 sg13g2_o21ai_1 _515_ (.B1(_150_),
    .Y(_151_),
    .A1(_036_),
    .A2(_138_));
 sg13g2_nand2_2 _516_ (.Y(_152_),
    .A(net9),
    .B(_137_));
 sg13g2_nand2_1 _517_ (.Y(_153_),
    .A(_140_),
    .B(_152_));
 sg13g2_xnor2_1 _518_ (.Y(_154_),
    .A(_037_),
    .B(_153_));
 sg13g2_nand2b_1 _519_ (.Y(_155_),
    .B(_152_),
    .A_N(\decoder_inst.counter[9] ));
 sg13g2_nand3_1 _520_ (.B(\decoder_inst.counter[9] ),
    .C(_137_),
    .A(net9),
    .Y(_156_));
 sg13g2_and3_1 _521_ (.X(_157_),
    .A(_154_),
    .B(_155_),
    .C(_156_));
 sg13g2_xor2_1 _522_ (.B(_139_),
    .A(_038_),
    .X(_158_));
 sg13g2_and2_1 _523_ (.A(_039_),
    .B(_137_),
    .X(_159_));
 sg13g2_a22oi_1 _524_ (.Y(_160_),
    .B1(_158_),
    .B2(_159_),
    .A2(_139_),
    .A1(_111_));
 sg13g2_xnor2_1 _525_ (.Y(_161_),
    .A(\decoder_inst.counter[6] ),
    .B(_137_));
 sg13g2_nand2_1 _526_ (.Y(_162_),
    .A(_158_),
    .B(_161_));
 sg13g2_xnor2_1 _527_ (.Y(_163_),
    .A(_040_),
    .B(_137_));
 sg13g2_nor2_1 _528_ (.A(\decoder_inst.counter[4] ),
    .B(_140_),
    .Y(_164_));
 sg13g2_xnor2_1 _529_ (.Y(_165_),
    .A(\decoder_inst.counter[4] ),
    .B(_140_));
 sg13g2_nor2_1 _530_ (.A(_163_),
    .B(_165_),
    .Y(_166_));
 sg13g2_nor2_1 _531_ (.A(_041_),
    .B(_152_),
    .Y(_167_));
 sg13g2_a21oi_1 _532_ (.A1(\decoder_inst.counter[3] ),
    .A2(_137_),
    .Y(_168_),
    .B1(_167_));
 sg13g2_nor2_1 _533_ (.A(\decoder_inst.counter[5] ),
    .B(_138_),
    .Y(_169_));
 sg13g2_a221oi_1 _534_ (.B2(_168_),
    .C1(_169_),
    .B1(_166_),
    .A1(_040_),
    .Y(_170_),
    .A2(_164_));
 sg13g2_o21ai_1 _535_ (.B1(_160_),
    .Y(_171_),
    .A1(_162_),
    .A2(_170_));
 sg13g2_o21ai_1 _536_ (.B1(_155_),
    .Y(_172_),
    .A1(\decoder_inst.counter[8] ),
    .A2(_153_));
 sg13g2_nand3_1 _537_ (.B(_158_),
    .C(_161_),
    .A(_157_),
    .Y(_173_));
 sg13g2_a21oi_1 _538_ (.A1(_157_),
    .A2(_171_),
    .Y(_174_),
    .B1(_172_));
 sg13g2_or2_1 _539_ (.X(_175_),
    .B(_151_),
    .A(_149_));
 sg13g2_nor3_1 _540_ (.A(\decoder_inst.counter[10] ),
    .B(_137_),
    .C(_149_),
    .Y(_176_));
 sg13g2_a22oi_1 _541_ (.Y(_177_),
    .B1(_176_),
    .B2(_035_),
    .A2(_146_),
    .A1(_034_));
 sg13g2_o21ai_1 _542_ (.B1(_177_),
    .Y(_178_),
    .A1(_174_),
    .A2(_175_));
 sg13g2_nor2b_1 _543_ (.A(_145_),
    .B_N(_178_),
    .Y(_179_));
 sg13g2_nor3_1 _544_ (.A(\decoder_inst.counter[16] ),
    .B(\decoder_inst.counter[17] ),
    .C(_140_),
    .Y(_180_));
 sg13g2_nor2b_1 _545_ (.A(_141_),
    .B_N(_142_),
    .Y(_181_));
 sg13g2_nor3_1 _546_ (.A(_179_),
    .B(_180_),
    .C(_181_),
    .Y(_182_));
 sg13g2_or4_1 _547_ (.A(\decoder_inst.counter[29] ),
    .B(\decoder_inst.counter[28] ),
    .C(\decoder_inst.counter[27] ),
    .D(\decoder_inst.counter[26] ),
    .X(_183_));
 sg13g2_nor3_1 _548_ (.A(\decoder_inst.counter[30] ),
    .B(\decoder_inst.counter[31] ),
    .C(_183_),
    .Y(_184_));
 sg13g2_nor4_1 _549_ (.A(\decoder_inst.counter[25] ),
    .B(\decoder_inst.counter[24] ),
    .C(\decoder_inst.counter[23] ),
    .D(\decoder_inst.counter[22] ),
    .Y(_185_));
 sg13g2_nor4_1 _550_ (.A(\decoder_inst.counter[21] ),
    .B(\decoder_inst.counter[20] ),
    .C(\decoder_inst.counter[19] ),
    .D(\decoder_inst.counter[18] ),
    .Y(_186_));
 sg13g2_nand3_1 _551_ (.B(_185_),
    .C(_186_),
    .A(_184_),
    .Y(_187_));
 sg13g2_nand2b_1 _552_ (.Y(_188_),
    .B(_138_),
    .A_N(\decoder_inst.counter[3] ));
 sg13g2_and2_1 _553_ (.A(net150),
    .B(net78),
    .X(_189_));
 sg13g2_nand2_1 _554_ (.Y(_190_),
    .A(\decoder_inst.counter[1] ),
    .B(net78));
 sg13g2_a21oi_1 _555_ (.A1(\decoder_inst.counter[3] ),
    .A2(_137_),
    .Y(_191_),
    .B1(_190_));
 sg13g2_xnor2_1 _556_ (.Y(_192_),
    .A(\decoder_inst.counter[2] ),
    .B(_152_));
 sg13g2_nand4_1 _557_ (.B(_188_),
    .C(_191_),
    .A(_166_),
    .Y(_193_),
    .D(_192_));
 sg13g2_nor4_1 _558_ (.A(_145_),
    .B(_173_),
    .C(_175_),
    .D(_193_),
    .Y(_194_));
 sg13g2_or3_2 _559_ (.A(_182_),
    .B(_187_),
    .C(_194_),
    .X(_195_));
 sg13g2_nor2_1 _560_ (.A(net78),
    .B(net94),
    .Y(_000_));
 sg13g2_nor2_1 _561_ (.A(net150),
    .B(net78),
    .Y(_196_));
 sg13g2_nor3_1 _562_ (.A(_189_),
    .B(net94),
    .C(_196_),
    .Y(_011_));
 sg13g2_xnor2_1 _563_ (.Y(_197_),
    .A(net125),
    .B(_190_));
 sg13g2_nor2_1 _564_ (.A(net94),
    .B(net126),
    .Y(_022_));
 sg13g2_and3_1 _565_ (.X(_198_),
    .A(net154),
    .B(\decoder_inst.counter[2] ),
    .C(_189_));
 sg13g2_a21oi_1 _566_ (.A1(\decoder_inst.counter[2] ),
    .A2(_189_),
    .Y(_199_),
    .B1(net154));
 sg13g2_nor3_1 _567_ (.A(net94),
    .B(_198_),
    .C(net155),
    .Y(_025_));
 sg13g2_and2_1 _568_ (.A(net225),
    .B(_198_),
    .X(_200_));
 sg13g2_nor2_1 _569_ (.A(net225),
    .B(_198_),
    .Y(_201_));
 sg13g2_nor3_1 _570_ (.A(net95),
    .B(_200_),
    .C(net226),
    .Y(_026_));
 sg13g2_xor2_1 _571_ (.B(_200_),
    .A(net202),
    .X(_202_));
 sg13g2_nor2_1 _572_ (.A(net94),
    .B(net203),
    .Y(_027_));
 sg13g2_nand2_1 _573_ (.Y(_203_),
    .A(\decoder_inst.counter[5] ),
    .B(_200_));
 sg13g2_nor2_1 _574_ (.A(net138),
    .B(_203_),
    .Y(_204_));
 sg13g2_and2_1 _575_ (.A(net138),
    .B(_203_),
    .X(_205_));
 sg13g2_nor3_1 _576_ (.A(net94),
    .B(_204_),
    .C(net139),
    .Y(_028_));
 sg13g2_xor2_1 _577_ (.B(_204_),
    .A(net184),
    .X(_206_));
 sg13g2_nor2_1 _578_ (.A(net95),
    .B(net185),
    .Y(_029_));
 sg13g2_nor3_1 _579_ (.A(_111_),
    .B(_112_),
    .C(_203_),
    .Y(_207_));
 sg13g2_nand4_1 _580_ (.B(\decoder_inst.counter[6] ),
    .C(\decoder_inst.counter[5] ),
    .A(\decoder_inst.counter[7] ),
    .Y(_208_),
    .D(_200_));
 sg13g2_xnor2_1 _581_ (.Y(_209_),
    .A(net145),
    .B(_208_));
 sg13g2_nor2_1 _582_ (.A(net94),
    .B(net146),
    .Y(_030_));
 sg13g2_a21oi_1 _583_ (.A1(\decoder_inst.counter[8] ),
    .A2(_207_),
    .Y(_210_),
    .B1(net238));
 sg13g2_nand3_1 _584_ (.B(\decoder_inst.counter[8] ),
    .C(_207_),
    .A(net238),
    .Y(_211_));
 sg13g2_nand2b_1 _585_ (.Y(_212_),
    .B(_211_),
    .A_N(net239));
 sg13g2_nor2_1 _586_ (.A(net94),
    .B(net240),
    .Y(_031_));
 sg13g2_and2_1 _587_ (.A(net210),
    .B(_211_),
    .X(_213_));
 sg13g2_nor2_1 _588_ (.A(net210),
    .B(_211_),
    .Y(_214_));
 sg13g2_nor3_1 _589_ (.A(net97),
    .B(net211),
    .C(_214_),
    .Y(_001_));
 sg13g2_xor2_1 _590_ (.B(_214_),
    .A(net143),
    .X(_215_));
 sg13g2_nor2_1 _591_ (.A(net97),
    .B(net144),
    .Y(_002_));
 sg13g2_nand4_1 _592_ (.B(\decoder_inst.counter[10] ),
    .C(\decoder_inst.counter[9] ),
    .A(\decoder_inst.counter[11] ),
    .Y(_216_),
    .D(\decoder_inst.counter[8] ));
 sg13g2_nor2_2 _593_ (.A(_208_),
    .B(_216_),
    .Y(_217_));
 sg13g2_nand2_1 _594_ (.Y(_218_),
    .A(\decoder_inst.counter[12] ),
    .B(_217_));
 sg13g2_xnor2_1 _595_ (.Y(_219_),
    .A(net218),
    .B(_217_));
 sg13g2_nor2_1 _596_ (.A(net98),
    .B(net219),
    .Y(_003_));
 sg13g2_xnor2_1 _597_ (.Y(_220_),
    .A(net82),
    .B(_218_));
 sg13g2_nor2_1 _598_ (.A(net98),
    .B(net83),
    .Y(_004_));
 sg13g2_and3_1 _599_ (.X(_221_),
    .A(\decoder_inst.counter[13] ),
    .B(\decoder_inst.counter[12] ),
    .C(_217_));
 sg13g2_xnor2_1 _600_ (.Y(_222_),
    .A(net200),
    .B(_221_));
 sg13g2_nor2_1 _601_ (.A(net95),
    .B(net201),
    .Y(_005_));
 sg13g2_a21oi_1 _602_ (.A1(\decoder_inst.counter[14] ),
    .A2(_221_),
    .Y(_223_),
    .B1(net160));
 sg13g2_and3_1 _603_ (.X(_224_),
    .A(net160),
    .B(net200),
    .C(_221_));
 sg13g2_nor3_1 _604_ (.A(net95),
    .B(net161),
    .C(_224_),
    .Y(_006_));
 sg13g2_xnor2_1 _605_ (.Y(_225_),
    .A(net222),
    .B(_224_));
 sg13g2_nor2_1 _606_ (.A(net95),
    .B(_225_),
    .Y(_007_));
 sg13g2_nor2_1 _607_ (.A(net75),
    .B(net95),
    .Y(_008_));
 sg13g2_a21oi_1 _608_ (.A1(net101),
    .A2(net1),
    .Y(_043_),
    .B1(_121_));
 sg13g2_a21oi_1 _609_ (.A1(net102),
    .A2(net2),
    .Y(_044_),
    .B1(_121_));
 sg13g2_a21oi_1 _610_ (.A1(net101),
    .A2(net3),
    .Y(_045_),
    .B1(_121_));
 sg13g2_a21oi_1 _611_ (.A1(net101),
    .A2(net4),
    .Y(_046_),
    .B1(_121_));
 sg13g2_a21oi_1 _612_ (.A1(net101),
    .A2(net5),
    .Y(_047_),
    .B1(_121_));
 sg13g2_a21oi_1 _613_ (.A1(net101),
    .A2(net6),
    .Y(_048_),
    .B1(_121_));
 sg13g2_a21oi_1 _614_ (.A1(net101),
    .A2(net7),
    .Y(_049_),
    .B1(_121_));
 sg13g2_a21oi_1 _615_ (.A1(net101),
    .A2(net8),
    .Y(_050_),
    .B1(_121_));
 sg13g2_nand2b_2 _616_ (.Y(_226_),
    .B(net1),
    .A_N(net101));
 sg13g2_nor2_1 _617_ (.A(\decoder_inst.signal_in_prev ),
    .B(_226_),
    .Y(_227_));
 sg13g2_nor2_1 _618_ (.A(net188),
    .B(_227_),
    .Y(_228_));
 sg13g2_nor3_1 _619_ (.A(\decoder_inst.signal_in_prev ),
    .B(_122_),
    .C(_226_),
    .Y(_229_));
 sg13g2_nor3_1 _620_ (.A(net96),
    .B(net189),
    .C(_229_),
    .Y(_051_));
 sg13g2_nor2_1 _621_ (.A(net163),
    .B(_229_),
    .Y(_230_));
 sg13g2_nor4_2 _622_ (.A(\decoder_inst.signal_in_prev ),
    .B(_122_),
    .C(_123_),
    .Y(_231_),
    .D(_226_));
 sg13g2_nor3_1 _623_ (.A(net97),
    .B(net164),
    .C(_231_),
    .Y(_052_));
 sg13g2_nor2_1 _624_ (.A(net176),
    .B(_231_),
    .Y(_232_));
 sg13g2_and2_1 _625_ (.A(net176),
    .B(_231_),
    .X(_233_));
 sg13g2_nor3_1 _626_ (.A(net96),
    .B(net177),
    .C(_233_),
    .Y(_053_));
 sg13g2_nor2_1 _627_ (.A(net196),
    .B(_233_),
    .Y(_234_));
 sg13g2_and2_1 _628_ (.A(net196),
    .B(_233_),
    .X(_235_));
 sg13g2_nor3_1 _629_ (.A(net91),
    .B(_234_),
    .C(_235_),
    .Y(_054_));
 sg13g2_nand4_1 _630_ (.B(net196),
    .C(net186),
    .A(net176),
    .Y(_236_),
    .D(_231_));
 sg13g2_xnor2_1 _631_ (.Y(_237_),
    .A(net186),
    .B(_235_));
 sg13g2_nor2_1 _632_ (.A(net92),
    .B(net187),
    .Y(_055_));
 sg13g2_nor2_2 _633_ (.A(_124_),
    .B(_236_),
    .Y(_238_));
 sg13g2_and2_1 _634_ (.A(_124_),
    .B(_236_),
    .X(_239_));
 sg13g2_nor3_1 _635_ (.A(net90),
    .B(_238_),
    .C(_239_),
    .Y(_056_));
 sg13g2_xnor2_1 _636_ (.Y(_240_),
    .A(net223),
    .B(_238_));
 sg13g2_nor2_1 _637_ (.A(net90),
    .B(net224),
    .Y(_057_));
 sg13g2_a21oi_1 _638_ (.A1(\decoder_inst.frequency[6] ),
    .A2(_238_),
    .Y(_241_),
    .B1(net129));
 sg13g2_nand2_1 _639_ (.Y(_242_),
    .A(net223),
    .B(net129));
 sg13g2_nor3_1 _640_ (.A(_124_),
    .B(_236_),
    .C(_242_),
    .Y(_243_));
 sg13g2_nor3_1 _641_ (.A(net89),
    .B(net130),
    .C(_243_),
    .Y(_058_));
 sg13g2_nor4_2 _642_ (.A(_124_),
    .B(_125_),
    .C(_236_),
    .Y(_244_),
    .D(_242_));
 sg13g2_nor2_1 _643_ (.A(net191),
    .B(_243_),
    .Y(_245_));
 sg13g2_nor3_1 _644_ (.A(net91),
    .B(_244_),
    .C(net192),
    .Y(_059_));
 sg13g2_xnor2_1 _645_ (.Y(_246_),
    .A(net233),
    .B(_244_));
 sg13g2_nor2_1 _646_ (.A(net91),
    .B(net234),
    .Y(_060_));
 sg13g2_a21oi_1 _647_ (.A1(net233),
    .A2(_244_),
    .Y(_247_),
    .B1(net244));
 sg13g2_nand3_1 _648_ (.B(net244),
    .C(_244_),
    .A(net233),
    .Y(_248_));
 sg13g2_nand2b_1 _649_ (.Y(_249_),
    .B(_248_),
    .A_N(_247_));
 sg13g2_nor2_1 _650_ (.A(net91),
    .B(_249_),
    .Y(_061_));
 sg13g2_nand4_1 _651_ (.B(\decoder_inst.frequency[10] ),
    .C(\decoder_inst.frequency[11] ),
    .A(\decoder_inst.frequency[9] ),
    .Y(_250_),
    .D(_244_));
 sg13g2_inv_1 _652_ (.Y(_251_),
    .A(_250_));
 sg13g2_xor2_1 _653_ (.B(_248_),
    .A(net229),
    .X(_252_));
 sg13g2_nor2_1 _654_ (.A(net91),
    .B(net230),
    .Y(_062_));
 sg13g2_xor2_1 _655_ (.B(_250_),
    .A(net236),
    .X(_253_));
 sg13g2_nor2_1 _656_ (.A(net89),
    .B(net237),
    .Y(_063_));
 sg13g2_a21oi_1 _657_ (.A1(\decoder_inst.frequency[12] ),
    .A2(_251_),
    .Y(_254_),
    .B1(net166));
 sg13g2_nand2_1 _658_ (.Y(_255_),
    .A(\decoder_inst.frequency[12] ),
    .B(net166));
 sg13g2_nor2_1 _659_ (.A(_250_),
    .B(_255_),
    .Y(_256_));
 sg13g2_nor3_1 _660_ (.A(net89),
    .B(net167),
    .C(_256_),
    .Y(_064_));
 sg13g2_xnor2_1 _661_ (.Y(_257_),
    .A(net231),
    .B(_256_));
 sg13g2_nor2_1 _662_ (.A(net90),
    .B(net232),
    .Y(_065_));
 sg13g2_nor4_2 _663_ (.A(_126_),
    .B(_127_),
    .C(_250_),
    .Y(_258_),
    .D(_255_));
 sg13g2_a21oi_1 _664_ (.A1(\decoder_inst.frequency[14] ),
    .A2(_256_),
    .Y(_259_),
    .B1(net151));
 sg13g2_nor3_1 _665_ (.A(net89),
    .B(_258_),
    .C(net152),
    .Y(_066_));
 sg13g2_nor2_1 _666_ (.A(net213),
    .B(_258_),
    .Y(_260_));
 sg13g2_and2_1 _667_ (.A(net213),
    .B(_258_),
    .X(_261_));
 sg13g2_nor3_1 _668_ (.A(net89),
    .B(net214),
    .C(_261_),
    .Y(_067_));
 sg13g2_and2_1 _669_ (.A(net215),
    .B(_261_),
    .X(_262_));
 sg13g2_nor2_1 _670_ (.A(net215),
    .B(_261_),
    .Y(_263_));
 sg13g2_nor3_1 _671_ (.A(net89),
    .B(_262_),
    .C(_263_),
    .Y(_068_));
 sg13g2_and2_1 _672_ (.A(net168),
    .B(_262_),
    .X(_264_));
 sg13g2_nand4_1 _673_ (.B(\decoder_inst.frequency[17] ),
    .C(net168),
    .A(\decoder_inst.frequency[16] ),
    .Y(_265_),
    .D(_258_));
 sg13g2_nor2_1 _674_ (.A(net168),
    .B(_262_),
    .Y(_266_));
 sg13g2_nor3_1 _675_ (.A(net87),
    .B(_264_),
    .C(net169),
    .Y(_069_));
 sg13g2_nor2_1 _676_ (.A(net157),
    .B(_264_),
    .Y(_267_));
 sg13g2_nor2_1 _677_ (.A(_128_),
    .B(_265_),
    .Y(_268_));
 sg13g2_nor3_1 _678_ (.A(net87),
    .B(net158),
    .C(_268_),
    .Y(_070_));
 sg13g2_nor2_1 _679_ (.A(net173),
    .B(_268_),
    .Y(_269_));
 sg13g2_nor3_1 _680_ (.A(_128_),
    .B(_129_),
    .C(_265_),
    .Y(_270_));
 sg13g2_nor3_1 _681_ (.A(net87),
    .B(net174),
    .C(_270_),
    .Y(_071_));
 sg13g2_nor2_1 _682_ (.A(net207),
    .B(_270_),
    .Y(_271_));
 sg13g2_nor4_2 _683_ (.A(_128_),
    .B(_129_),
    .C(_130_),
    .Y(_272_),
    .D(_265_));
 sg13g2_nor3_1 _684_ (.A(net87),
    .B(net208),
    .C(_272_),
    .Y(_072_));
 sg13g2_nor2_1 _685_ (.A(net193),
    .B(_272_),
    .Y(_273_));
 sg13g2_and2_1 _686_ (.A(net193),
    .B(_272_),
    .X(_274_));
 sg13g2_nor3_1 _687_ (.A(net87),
    .B(net194),
    .C(_274_),
    .Y(_073_));
 sg13g2_nor2_1 _688_ (.A(net195),
    .B(_274_),
    .Y(_275_));
 sg13g2_and2_1 _689_ (.A(net195),
    .B(_274_),
    .X(_276_));
 sg13g2_nor3_1 _690_ (.A(net87),
    .B(_275_),
    .C(_276_),
    .Y(_074_));
 sg13g2_nor2_1 _691_ (.A(net216),
    .B(_276_),
    .Y(_277_));
 sg13g2_and2_1 _692_ (.A(net216),
    .B(_276_),
    .X(_278_));
 sg13g2_nand4_1 _693_ (.B(\decoder_inst.frequency[23] ),
    .C(\decoder_inst.frequency[24] ),
    .A(net193),
    .Y(_279_),
    .D(_272_));
 sg13g2_nor3_1 _694_ (.A(net87),
    .B(_277_),
    .C(_278_),
    .Y(_075_));
 sg13g2_nor2_1 _695_ (.A(net197),
    .B(_278_),
    .Y(_280_));
 sg13g2_nor2_1 _696_ (.A(_131_),
    .B(_279_),
    .Y(_281_));
 sg13g2_nor3_1 _697_ (.A(net87),
    .B(net198),
    .C(_281_),
    .Y(_076_));
 sg13g2_nor2_1 _698_ (.A(net170),
    .B(_281_),
    .Y(_282_));
 sg13g2_nor3_1 _699_ (.A(_131_),
    .B(_132_),
    .C(_279_),
    .Y(_283_));
 sg13g2_nor3_1 _700_ (.A(net88),
    .B(net171),
    .C(_283_),
    .Y(_077_));
 sg13g2_nor2_1 _701_ (.A(net147),
    .B(_283_),
    .Y(_284_));
 sg13g2_nor4_2 _702_ (.A(_131_),
    .B(_132_),
    .C(_133_),
    .Y(_285_),
    .D(_279_));
 sg13g2_nor3_1 _703_ (.A(net88),
    .B(net148),
    .C(_285_),
    .Y(_078_));
 sg13g2_nor2_1 _704_ (.A(net220),
    .B(_285_),
    .Y(_286_));
 sg13g2_and2_1 _705_ (.A(net220),
    .B(_285_),
    .X(_287_));
 sg13g2_nor3_1 _706_ (.A(net88),
    .B(net221),
    .C(_287_),
    .Y(_079_));
 sg13g2_nor2_1 _707_ (.A(net178),
    .B(_287_),
    .Y(_288_));
 sg13g2_nand3_1 _708_ (.B(net178),
    .C(_285_),
    .A(\decoder_inst.frequency[28] ),
    .Y(_289_));
 sg13g2_nand2b_1 _709_ (.Y(_290_),
    .B(_289_),
    .A_N(net88));
 sg13g2_nor2_1 _710_ (.A(net179),
    .B(_290_),
    .Y(_080_));
 sg13g2_nand4_1 _711_ (.B(net178),
    .C(net134),
    .A(net220),
    .Y(_291_),
    .D(_285_));
 sg13g2_nand2b_1 _712_ (.Y(_292_),
    .B(_291_),
    .A_N(net88));
 sg13g2_a21oi_1 _713_ (.A1(_134_),
    .A2(_289_),
    .Y(_081_),
    .B1(_292_));
 sg13g2_and2_1 _714_ (.A(_135_),
    .B(_291_),
    .X(_293_));
 sg13g2_nor2_1 _715_ (.A(_135_),
    .B(_291_),
    .Y(_294_));
 sg13g2_nor3_1 _716_ (.A(net88),
    .B(_293_),
    .C(_294_),
    .Y(_082_));
 sg13g2_nor4_1 _717_ (.A(\decoder_inst.frequency[12] ),
    .B(\decoder_inst.frequency[13] ),
    .C(\decoder_inst.frequency[14] ),
    .D(\decoder_inst.frequency[15] ),
    .Y(_295_));
 sg13g2_nor4_1 _718_ (.A(\decoder_inst.frequency[8] ),
    .B(\decoder_inst.frequency[9] ),
    .C(\decoder_inst.frequency[10] ),
    .D(\decoder_inst.frequency[11] ),
    .Y(_296_));
 sg13g2_nand2_1 _719_ (.Y(_297_),
    .A(_295_),
    .B(_296_));
 sg13g2_nor4_1 _720_ (.A(\decoder_inst.frequency[20] ),
    .B(\decoder_inst.frequency[21] ),
    .C(\decoder_inst.frequency[22] ),
    .D(\decoder_inst.frequency[23] ),
    .Y(_298_));
 sg13g2_nor3_1 _721_ (.A(\decoder_inst.frequency[16] ),
    .B(\decoder_inst.frequency[17] ),
    .C(\decoder_inst.frequency[18] ),
    .Y(_299_));
 sg13g2_nand3_1 _722_ (.B(_298_),
    .C(_299_),
    .A(_128_),
    .Y(_300_));
 sg13g2_nor4_1 _723_ (.A(\decoder_inst.frequency[28] ),
    .B(\decoder_inst.frequency[29] ),
    .C(\decoder_inst.frequency[30] ),
    .D(\decoder_inst.frequency[31] ),
    .Y(_301_));
 sg13g2_nor3_1 _724_ (.A(\decoder_inst.frequency[24] ),
    .B(\decoder_inst.frequency[25] ),
    .C(\decoder_inst.frequency[26] ),
    .Y(_302_));
 sg13g2_nand3_1 _725_ (.B(_301_),
    .C(_302_),
    .A(_133_),
    .Y(_303_));
 sg13g2_nor3_2 _726_ (.A(_297_),
    .B(_300_),
    .C(_303_),
    .Y(_304_));
 sg13g2_a21oi_1 _727_ (.A1(\decoder_inst.frequency[0] ),
    .A2(_304_),
    .Y(_305_),
    .B1(\decoder_inst.frequency[8] ));
 sg13g2_nor2_1 _728_ (.A(net141),
    .B(net97),
    .Y(_306_));
 sg13g2_a21oi_1 _729_ (.A1(net96),
    .A2(_305_),
    .Y(_083_),
    .B1(_306_));
 sg13g2_nor2_1 _730_ (.A(net127),
    .B(net96),
    .Y(_307_));
 sg13g2_a21oi_1 _731_ (.A1(\decoder_inst.frequency[1] ),
    .A2(_304_),
    .Y(_308_),
    .B1(\decoder_inst.frequency[9] ));
 sg13g2_a21oi_1 _732_ (.A1(net96),
    .A2(_308_),
    .Y(_084_),
    .B1(_307_));
 sg13g2_a21oi_1 _733_ (.A1(\decoder_inst.frequency[2] ),
    .A2(_304_),
    .Y(_309_),
    .B1(\decoder_inst.frequency[10] ));
 sg13g2_nor2_1 _734_ (.A(net123),
    .B(net96),
    .Y(_310_));
 sg13g2_a21oi_1 _735_ (.A1(net96),
    .A2(_309_),
    .Y(_085_),
    .B1(_310_));
 sg13g2_nor2_1 _736_ (.A(net132),
    .B(net96),
    .Y(_311_));
 sg13g2_a21oi_1 _737_ (.A1(\decoder_inst.frequency[3] ),
    .A2(_304_),
    .Y(_312_),
    .B1(\decoder_inst.frequency[11] ));
 sg13g2_a21oi_1 _738_ (.A1(net91),
    .A2(_312_),
    .Y(_086_),
    .B1(_311_));
 sg13g2_nor2_1 _739_ (.A(net86),
    .B(net91),
    .Y(_313_));
 sg13g2_a21oi_1 _740_ (.A1(\decoder_inst.frequency[4] ),
    .A2(_304_),
    .Y(_314_),
    .B1(\decoder_inst.frequency[12] ));
 sg13g2_a21oi_1 _741_ (.A1(net92),
    .A2(_314_),
    .Y(_087_),
    .B1(_313_));
 sg13g2_a21oi_1 _742_ (.A1(\decoder_inst.frequency[5] ),
    .A2(_304_),
    .Y(_315_),
    .B1(\decoder_inst.frequency[13] ));
 sg13g2_nor2_1 _743_ (.A(net136),
    .B(net92),
    .Y(_316_));
 sg13g2_a21oi_1 _744_ (.A1(net92),
    .A2(_315_),
    .Y(_088_),
    .B1(_316_));
 sg13g2_a21oi_1 _745_ (.A1(\decoder_inst.frequency[6] ),
    .A2(_304_),
    .Y(_317_),
    .B1(\decoder_inst.frequency[14] ));
 sg13g2_nor2_1 _746_ (.A(net84),
    .B(net90),
    .Y(_318_));
 sg13g2_a21oi_1 _747_ (.A1(net89),
    .A2(_317_),
    .Y(_089_),
    .B1(_318_));
 sg13g2_a21oi_1 _748_ (.A1(\decoder_inst.frequency[7] ),
    .A2(_304_),
    .Y(_319_),
    .B1(\decoder_inst.frequency[15] ));
 sg13g2_nor2_1 _749_ (.A(net121),
    .B(net91),
    .Y(_320_));
 sg13g2_a21oi_1 _750_ (.A1(net89),
    .A2(_319_),
    .Y(_090_),
    .B1(_320_));
 sg13g2_a22oi_1 _751_ (.Y(_321_),
    .B1(\encoder_inst.divide_value[1] ),
    .B2(_114_),
    .A2(\encoder_inst.divide_value[0] ),
    .A1(_110_));
 sg13g2_a21oi_1 _752_ (.A1(_113_),
    .A2(\encoder_inst.counter[1] ),
    .Y(_322_),
    .B1(_321_));
 sg13g2_o21ai_1 _753_ (.B1(_322_),
    .Y(_323_),
    .A1(\encoder_inst.divide_value[2] ),
    .A2(_116_));
 sg13g2_a22oi_1 _754_ (.Y(_324_),
    .B1(\encoder_inst.divide_value[2] ),
    .B2(_116_),
    .A2(_115_),
    .A1(\encoder_inst.divide_value[3] ));
 sg13g2_nand2b_1 _755_ (.Y(_325_),
    .B(\encoder_inst.counter[4] ),
    .A_N(\encoder_inst.divide_value[4] ));
 sg13g2_o21ai_1 _756_ (.B1(_325_),
    .Y(_326_),
    .A1(\encoder_inst.divide_value[3] ),
    .A2(_115_));
 sg13g2_a21oi_1 _757_ (.A1(_323_),
    .A2(_324_),
    .Y(_327_),
    .B1(_326_));
 sg13g2_nand2b_1 _758_ (.Y(_328_),
    .B(\encoder_inst.divide_value[4] ),
    .A_N(\encoder_inst.counter[4] ));
 sg13g2_o21ai_1 _759_ (.B1(_328_),
    .Y(_329_),
    .A1(_120_),
    .A2(\encoder_inst.counter[5] ));
 sg13g2_a22oi_1 _760_ (.Y(_330_),
    .B1(_120_),
    .B2(\encoder_inst.counter[5] ),
    .A2(\encoder_inst.counter[6] ),
    .A1(_118_));
 sg13g2_o21ai_1 _761_ (.B1(_330_),
    .Y(_331_),
    .A1(_327_),
    .A2(_329_));
 sg13g2_a22oi_1 _762_ (.Y(_332_),
    .B1(\encoder_inst.divide_value[6] ),
    .B2(_119_),
    .A2(_117_),
    .A1(\encoder_inst.divide_value[7] ));
 sg13g2_nor4_1 _763_ (.A(\encoder_inst.counter[11] ),
    .B(\encoder_inst.counter[10] ),
    .C(\encoder_inst.counter[9] ),
    .D(\encoder_inst.counter[8] ),
    .Y(_333_));
 sg13g2_nand2b_1 _764_ (.Y(_334_),
    .B(net241),
    .A_N(\encoder_inst.divide_value[7] ));
 sg13g2_nor4_1 _765_ (.A(\encoder_inst.counter[15] ),
    .B(\encoder_inst.counter[14] ),
    .C(\encoder_inst.counter[12] ),
    .D(\encoder_inst.counter[13] ),
    .Y(_335_));
 sg13g2_nand3_1 _766_ (.B(_334_),
    .C(_335_),
    .A(_333_),
    .Y(_336_));
 sg13g2_a21oi_2 _767_ (.B1(_336_),
    .Y(_337_),
    .A2(_332_),
    .A1(_331_));
 sg13g2_nand2_2 _768_ (.Y(_338_),
    .A(net115),
    .B(_337_));
 sg13g2_and3_1 _769_ (.X(_091_),
    .A(net115),
    .B(net76),
    .C(_337_));
 sg13g2_xnor2_1 _770_ (.Y(_339_),
    .A(net204),
    .B(\encoder_inst.counter[1] ));
 sg13g2_nor2_1 _771_ (.A(_338_),
    .B(net205),
    .Y(_092_));
 sg13g2_and3_1 _772_ (.X(_340_),
    .A(\encoder_inst.counter[0] ),
    .B(\encoder_inst.counter[1] ),
    .C(net118));
 sg13g2_a21oi_1 _773_ (.A1(\encoder_inst.counter[0] ),
    .A2(\encoder_inst.counter[1] ),
    .Y(_341_),
    .B1(net118));
 sg13g2_nor3_1 _774_ (.A(_338_),
    .B(_340_),
    .C(net119),
    .Y(_093_));
 sg13g2_nor2_1 _775_ (.A(net181),
    .B(_340_),
    .Y(_342_));
 sg13g2_and2_1 _776_ (.A(net181),
    .B(_340_),
    .X(_343_));
 sg13g2_nor3_1 _777_ (.A(_338_),
    .B(net182),
    .C(_343_),
    .Y(_094_));
 sg13g2_xnor2_1 _778_ (.Y(_344_),
    .A(net227),
    .B(_343_));
 sg13g2_nor2_1 _779_ (.A(_338_),
    .B(_344_),
    .Y(_095_));
 sg13g2_a21o_1 _780_ (.A2(_343_),
    .A1(net227),
    .B1(net245),
    .X(_345_));
 sg13g2_nand3_1 _781_ (.B(net245),
    .C(_343_),
    .A(net227),
    .Y(_346_));
 sg13g2_and4_1 _782_ (.A(net115),
    .B(_337_),
    .C(_345_),
    .D(_346_),
    .X(_096_));
 sg13g2_nand2_1 _783_ (.Y(_347_),
    .A(_119_),
    .B(_346_));
 sg13g2_or2_1 _784_ (.X(_348_),
    .B(_346_),
    .A(_119_));
 sg13g2_and4_1 _785_ (.A(net115),
    .B(_337_),
    .C(_347_),
    .D(_348_),
    .X(_097_));
 sg13g2_xnor2_1 _786_ (.Y(_349_),
    .A(_117_),
    .B(_348_));
 sg13g2_nor2_1 _787_ (.A(_338_),
    .B(net242),
    .Y(_098_));
 sg13g2_nor2_1 _788_ (.A(net217),
    .B(net114),
    .Y(_350_));
 sg13g2_a21oi_1 _789_ (.A1(net114),
    .A2(_226_),
    .Y(_107_),
    .B1(_350_));
 sg13g2_o21ai_1 _790_ (.B1(net114),
    .Y(_351_),
    .A1(net79),
    .A2(_337_));
 sg13g2_a21oi_1 _791_ (.A1(_109_),
    .A2(_337_),
    .Y(_108_),
    .B1(net80));
 sg13g2_dfrbp_1 _792_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net61),
    .D(_043_),
    .Q_N(_415_),
    .Q(\encoder_inst.divide_value[0] ));
 sg13g2_dfrbp_1 _793_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net68),
    .D(_044_),
    .Q_N(_414_),
    .Q(\encoder_inst.divide_value[1] ));
 sg13g2_dfrbp_1 _794_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net67),
    .D(_045_),
    .Q_N(_413_),
    .Q(\encoder_inst.divide_value[2] ));
 sg13g2_dfrbp_1 _795_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net66),
    .D(_046_),
    .Q_N(_412_),
    .Q(\encoder_inst.divide_value[3] ));
 sg13g2_dfrbp_1 _796_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net65),
    .D(_047_),
    .Q_N(_411_),
    .Q(\encoder_inst.divide_value[4] ));
 sg13g2_dfrbp_1 _797_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net64),
    .D(_048_),
    .Q_N(_410_),
    .Q(\encoder_inst.divide_value[5] ));
 sg13g2_dfrbp_1 _798_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net63),
    .D(_049_),
    .Q_N(_409_),
    .Q(\encoder_inst.divide_value[6] ));
 sg13g2_dfrbp_1 _799_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net62),
    .D(_050_),
    .Q_N(_408_),
    .Q(\encoder_inst.divide_value[7] ));
 sg13g2_dfrbp_1 _800_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net115),
    .D(net190),
    .Q_N(_407_),
    .Q(\decoder_inst.frequency[0] ));
 sg13g2_dfrbp_1 _801_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net115),
    .D(net165),
    .Q_N(_406_),
    .Q(\decoder_inst.frequency[1] ));
 sg13g2_dfrbp_1 _802_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net108),
    .D(_053_),
    .Q_N(_405_),
    .Q(\decoder_inst.frequency[2] ));
 sg13g2_dfrbp_1 _803_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net107),
    .D(_054_),
    .Q_N(_404_),
    .Q(\decoder_inst.frequency[3] ));
 sg13g2_dfrbp_1 _804_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net107),
    .D(_055_),
    .Q_N(_403_),
    .Q(\decoder_inst.frequency[4] ));
 sg13g2_dfrbp_1 _805_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net106),
    .D(_056_),
    .Q_N(_402_),
    .Q(\decoder_inst.frequency[5] ));
 sg13g2_dfrbp_1 _806_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net106),
    .D(_057_),
    .Q_N(_401_),
    .Q(\decoder_inst.frequency[6] ));
 sg13g2_dfrbp_1 _807_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net106),
    .D(net131),
    .Q_N(_400_),
    .Q(\decoder_inst.frequency[7] ));
 sg13g2_dfrbp_1 _808_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net107),
    .D(_059_),
    .Q_N(_399_),
    .Q(\decoder_inst.frequency[8] ));
 sg13g2_dfrbp_1 _809_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net107),
    .D(_060_),
    .Q_N(_398_),
    .Q(\decoder_inst.frequency[9] ));
 sg13g2_dfrbp_1 _810_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net107),
    .D(_061_),
    .Q_N(_397_),
    .Q(\decoder_inst.frequency[10] ));
 sg13g2_dfrbp_1 _811_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net107),
    .D(_062_),
    .Q_N(_396_),
    .Q(\decoder_inst.frequency[11] ));
 sg13g2_dfrbp_1 _812_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net105),
    .D(_063_),
    .Q_N(_395_),
    .Q(\decoder_inst.frequency[12] ));
 sg13g2_dfrbp_1 _813_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net105),
    .D(_064_),
    .Q_N(_394_),
    .Q(\decoder_inst.frequency[13] ));
 sg13g2_dfrbp_1 _814_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net106),
    .D(_065_),
    .Q_N(_393_),
    .Q(\decoder_inst.frequency[14] ));
 sg13g2_dfrbp_1 _815_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net105),
    .D(net153),
    .Q_N(_392_),
    .Q(\decoder_inst.frequency[15] ));
 sg13g2_dfrbp_1 _816_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net105),
    .D(_067_),
    .Q_N(_391_),
    .Q(\decoder_inst.frequency[16] ));
 sg13g2_dfrbp_1 _817_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net105),
    .D(_068_),
    .Q_N(_390_),
    .Q(\decoder_inst.frequency[17] ));
 sg13g2_dfrbp_1 _818_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net105),
    .D(_069_),
    .Q_N(_389_),
    .Q(\decoder_inst.frequency[18] ));
 sg13g2_dfrbp_1 _819_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net104),
    .D(net159),
    .Q_N(_388_),
    .Q(\decoder_inst.frequency[19] ));
 sg13g2_dfrbp_1 _820_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net104),
    .D(net175),
    .Q_N(_387_),
    .Q(\decoder_inst.frequency[20] ));
 sg13g2_dfrbp_1 _821_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net104),
    .D(net209),
    .Q_N(_386_),
    .Q(\decoder_inst.frequency[21] ));
 sg13g2_dfrbp_1 _822_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net104),
    .D(_073_),
    .Q_N(_385_),
    .Q(\decoder_inst.frequency[22] ));
 sg13g2_dfrbp_1 _823_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net104),
    .D(_074_),
    .Q_N(_384_),
    .Q(\decoder_inst.frequency[23] ));
 sg13g2_dfrbp_1 _824_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net104),
    .D(_075_),
    .Q_N(_383_),
    .Q(\decoder_inst.frequency[24] ));
 sg13g2_dfrbp_1 _825_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net104),
    .D(net199),
    .Q_N(_382_),
    .Q(\decoder_inst.frequency[25] ));
 sg13g2_dfrbp_1 _826_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net104),
    .D(net172),
    .Q_N(_381_),
    .Q(\decoder_inst.frequency[26] ));
 sg13g2_dfrbp_1 _827_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net109),
    .D(net149),
    .Q_N(_380_),
    .Q(\decoder_inst.frequency[27] ));
 sg13g2_dfrbp_1 _828_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net103),
    .D(_079_),
    .Q_N(_379_),
    .Q(\decoder_inst.frequency[28] ));
 sg13g2_dfrbp_1 _829_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net103),
    .D(net180),
    .Q_N(_378_),
    .Q(\decoder_inst.frequency[29] ));
 sg13g2_dfrbp_1 _830_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net103),
    .D(net135),
    .Q_N(_377_),
    .Q(\decoder_inst.frequency[30] ));
 sg13g2_dfrbp_1 _831_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net109),
    .D(_082_),
    .Q_N(_416_),
    .Q(\decoder_inst.frequency[31] ));
 sg13g2_dfrbp_1 _832_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net103),
    .D(_000_),
    .Q_N(_417_),
    .Q(\decoder_inst.counter[0] ));
 sg13g2_dfrbp_1 _833_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net113),
    .D(_011_),
    .Q_N(_418_),
    .Q(\decoder_inst.counter[1] ));
 sg13g2_dfrbp_1 _834_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net113),
    .D(_022_),
    .Q_N(_041_),
    .Q(\decoder_inst.counter[2] ));
 sg13g2_dfrbp_1 _835_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net113),
    .D(net156),
    .Q_N(_419_),
    .Q(\decoder_inst.counter[3] ));
 sg13g2_dfrbp_1 _836_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net113),
    .D(_026_),
    .Q_N(_420_),
    .Q(\decoder_inst.counter[4] ));
 sg13g2_dfrbp_1 _837_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net113),
    .D(_027_),
    .Q_N(_040_),
    .Q(\decoder_inst.counter[5] ));
 sg13g2_dfrbp_1 _838_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net103),
    .D(net140),
    .Q_N(_039_),
    .Q(\decoder_inst.counter[6] ));
 sg13g2_dfrbp_1 _839_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net103),
    .D(_029_),
    .Q_N(_038_),
    .Q(\decoder_inst.counter[7] ));
 sg13g2_dfrbp_1 _840_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net103),
    .D(_030_),
    .Q_N(_037_),
    .Q(\decoder_inst.counter[8] ));
 sg13g2_dfrbp_1 _841_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net103),
    .D(_031_),
    .Q_N(_421_),
    .Q(\decoder_inst.counter[9] ));
 sg13g2_dfrbp_1 _842_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net114),
    .D(net212),
    .Q_N(_036_),
    .Q(\decoder_inst.counter[10] ));
 sg13g2_dfrbp_1 _843_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net114),
    .D(_002_),
    .Q_N(_035_),
    .Q(\decoder_inst.counter[11] ));
 sg13g2_dfrbp_1 _844_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net114),
    .D(_003_),
    .Q_N(_422_),
    .Q(\decoder_inst.counter[12] ));
 sg13g2_dfrbp_1 _845_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net114),
    .D(_004_),
    .Q_N(_034_),
    .Q(\decoder_inst.counter[13] ));
 sg13g2_dfrbp_1 _846_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net116),
    .D(_005_),
    .Q_N(_423_),
    .Q(\decoder_inst.counter[14] ));
 sg13g2_dfrbp_1 _847_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net112),
    .D(net162),
    .Q_N(_424_),
    .Q(\decoder_inst.counter[15] ));
 sg13g2_dfrbp_1 _848_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net112),
    .D(_007_),
    .Q_N(_425_),
    .Q(\decoder_inst.counter[16] ));
 sg13g2_dfrbp_1 _849_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net112),
    .D(_008_),
    .Q_N(_033_),
    .Q(\decoder_inst.counter[17] ));
 sg13g2_dfrbp_1 _850_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net110),
    .D(net48),
    .Q_N(_426_),
    .Q(\decoder_inst.counter[18] ));
 sg13g2_dfrbp_1 _851_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net110),
    .D(net47),
    .Q_N(_427_),
    .Q(\decoder_inst.counter[19] ));
 sg13g2_dfrbp_1 _852_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net111),
    .D(net46),
    .Q_N(_428_),
    .Q(\decoder_inst.counter[20] ));
 sg13g2_dfrbp_1 _853_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net111),
    .D(net45),
    .Q_N(_429_),
    .Q(\decoder_inst.counter[21] ));
 sg13g2_dfrbp_1 _854_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net110),
    .D(net44),
    .Q_N(_430_),
    .Q(\decoder_inst.counter[22] ));
 sg13g2_dfrbp_1 _855_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net110),
    .D(net43),
    .Q_N(_431_),
    .Q(\decoder_inst.counter[23] ));
 sg13g2_dfrbp_1 _856_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net111),
    .D(net42),
    .Q_N(_432_),
    .Q(\decoder_inst.counter[24] ));
 sg13g2_dfrbp_1 _857_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net111),
    .D(net41),
    .Q_N(_433_),
    .Q(\decoder_inst.counter[25] ));
 sg13g2_dfrbp_1 _858_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net113),
    .D(net40),
    .Q_N(_434_),
    .Q(\decoder_inst.counter[26] ));
 sg13g2_dfrbp_1 _859_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net113),
    .D(net39),
    .Q_N(_435_),
    .Q(\decoder_inst.counter[27] ));
 sg13g2_dfrbp_1 _860_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net110),
    .D(net38),
    .Q_N(_436_),
    .Q(\decoder_inst.counter[28] ));
 sg13g2_dfrbp_1 _861_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net110),
    .D(net37),
    .Q_N(_437_),
    .Q(\decoder_inst.counter[29] ));
 sg13g2_dfrbp_1 _862_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net110),
    .D(net36),
    .Q_N(_438_),
    .Q(\decoder_inst.counter[30] ));
 sg13g2_dfrbp_1 _863_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net110),
    .D(net35),
    .Q_N(_376_),
    .Q(\decoder_inst.counter[31] ));
 sg13g2_dfrbp_1 _864_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net114),
    .D(net142),
    .Q_N(_375_),
    .Q(\decoder_inst.freq_out[0] ));
 sg13g2_dfrbp_1 _865_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net115),
    .D(net128),
    .Q_N(_374_),
    .Q(\decoder_inst.freq_out[1] ));
 sg13g2_dfrbp_1 _866_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net107),
    .D(net124),
    .Q_N(_373_),
    .Q(\decoder_inst.freq_out[2] ));
 sg13g2_dfrbp_1 _867_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net107),
    .D(net133),
    .Q_N(_372_),
    .Q(\decoder_inst.freq_out[3] ));
 sg13g2_dfrbp_1 _868_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net108),
    .D(net117),
    .Q_N(_371_),
    .Q(\decoder_inst.freq_out[4] ));
 sg13g2_dfrbp_1 _869_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net108),
    .D(net137),
    .Q_N(_370_),
    .Q(\decoder_inst.freq_out[5] ));
 sg13g2_dfrbp_1 _870_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net105),
    .D(net85),
    .Q_N(_369_),
    .Q(\decoder_inst.freq_out[6] ));
 sg13g2_dfrbp_1 _871_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net105),
    .D(net122),
    .Q_N(_368_),
    .Q(\decoder_inst.freq_out[7] ));
 sg13g2_dfrbp_1 _872_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net60),
    .D(net77),
    .Q_N(_042_),
    .Q(\encoder_inst.counter[0] ));
 sg13g2_dfrbp_1 _873_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net59),
    .D(net206),
    .Q_N(_367_),
    .Q(\encoder_inst.counter[1] ));
 sg13g2_dfrbp_1 _874_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net58),
    .D(net120),
    .Q_N(_366_),
    .Q(\encoder_inst.counter[2] ));
 sg13g2_dfrbp_1 _875_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net57),
    .D(net183),
    .Q_N(_365_),
    .Q(\encoder_inst.counter[3] ));
 sg13g2_dfrbp_1 _876_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net56),
    .D(net228),
    .Q_N(_364_),
    .Q(\encoder_inst.counter[4] ));
 sg13g2_dfrbp_1 _877_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net55),
    .D(net246),
    .Q_N(_363_),
    .Q(\encoder_inst.counter[5] ));
 sg13g2_dfrbp_1 _878_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net54),
    .D(net248),
    .Q_N(_362_),
    .Q(\encoder_inst.counter[6] ));
 sg13g2_dfrbp_1 _879_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net53),
    .D(net243),
    .Q_N(_361_),
    .Q(\encoder_inst.counter[7] ));
 sg13g2_dfrbp_1 _880_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net52),
    .D(net34),
    .Q_N(_360_),
    .Q(\encoder_inst.counter[8] ));
 sg13g2_dfrbp_1 _881_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net51),
    .D(net33),
    .Q_N(_359_),
    .Q(\encoder_inst.counter[9] ));
 sg13g2_dfrbp_1 _882_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net50),
    .D(net32),
    .Q_N(_358_),
    .Q(\encoder_inst.counter[10] ));
 sg13g2_dfrbp_1 _883_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net49),
    .D(net31),
    .Q_N(_357_),
    .Q(\encoder_inst.counter[11] ));
 sg13g2_dfrbp_1 _884_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net74),
    .D(net30),
    .Q_N(_356_),
    .Q(\encoder_inst.counter[12] ));
 sg13g2_dfrbp_1 _885_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net73),
    .D(net29),
    .Q_N(_355_),
    .Q(\encoder_inst.counter[13] ));
 sg13g2_dfrbp_1 _886_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net72),
    .D(net28),
    .Q_N(_354_),
    .Q(\encoder_inst.counter[14] ));
 sg13g2_dfrbp_1 _887_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net71),
    .D(net27),
    .Q_N(_353_),
    .Q(\encoder_inst.counter[15] ));
 sg13g2_dfrbp_1 _888_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net70),
    .D(_107_),
    .Q_N(_352_),
    .Q(\decoder_inst.signal_in_prev ));
 sg13g2_dfrbp_1 _889_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net69),
    .D(net81),
    .Q_N(_032_),
    .Q(\encoder_inst.out ));
 sg13g2_tiehi _882__50 (.L_HI(net50));
 sg13g2_tiehi _881__51 (.L_HI(net51));
 sg13g2_tiehi _880__52 (.L_HI(net52));
 sg13g2_tiehi _879__53 (.L_HI(net53));
 sg13g2_tiehi _878__54 (.L_HI(net54));
 sg13g2_tiehi _877__55 (.L_HI(net55));
 sg13g2_tiehi _876__56 (.L_HI(net56));
 sg13g2_tiehi _875__57 (.L_HI(net57));
 sg13g2_tiehi _874__58 (.L_HI(net58));
 sg13g2_tiehi _873__59 (.L_HI(net59));
 sg13g2_tiehi _872__60 (.L_HI(net60));
 sg13g2_tiehi _792__61 (.L_HI(net61));
 sg13g2_tiehi _799__62 (.L_HI(net62));
 sg13g2_tiehi _798__63 (.L_HI(net63));
 sg13g2_tiehi _797__64 (.L_HI(net64));
 sg13g2_tiehi _796__65 (.L_HI(net65));
 sg13g2_tiehi _795__66 (.L_HI(net66));
 sg13g2_tiehi _794__67 (.L_HI(net67));
 sg13g2_tiehi _793__68 (.L_HI(net68));
 sg13g2_tiehi _889__69 (.L_HI(net69));
 sg13g2_tiehi _888__70 (.L_HI(net70));
 sg13g2_tiehi _887__71 (.L_HI(net71));
 sg13g2_tiehi _886__72 (.L_HI(net72));
 sg13g2_tiehi _885__73 (.L_HI(net73));
 sg13g2_tiehi _884__74 (.L_HI(net74));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_mroblesh_12 (.L_LO(net12));
 sg13g2_tielo tt_um_mroblesh_13 (.L_LO(net13));
 sg13g2_tielo tt_um_mroblesh_14 (.L_LO(net14));
 sg13g2_tielo tt_um_mroblesh_15 (.L_LO(net15));
 sg13g2_tielo tt_um_mroblesh_16 (.L_LO(net16));
 sg13g2_tielo tt_um_mroblesh_17 (.L_LO(net17));
 sg13g2_tielo tt_um_mroblesh_18 (.L_LO(net18));
 sg13g2_tielo tt_um_mroblesh_19 (.L_LO(net19));
 sg13g2_tielo tt_um_mroblesh_20 (.L_LO(net20));
 sg13g2_tielo tt_um_mroblesh_21 (.L_LO(net21));
 sg13g2_tielo tt_um_mroblesh_22 (.L_LO(net22));
 sg13g2_tielo tt_um_mroblesh_23 (.L_LO(net23));
 sg13g2_tielo tt_um_mroblesh_24 (.L_LO(net24));
 sg13g2_tielo tt_um_mroblesh_25 (.L_LO(net25));
 sg13g2_tielo tt_um_mroblesh_26 (.L_LO(net26));
 sg13g2_tielo _887__27 (.L_LO(net27));
 sg13g2_tielo _886__28 (.L_LO(net28));
 sg13g2_tielo _885__29 (.L_LO(net29));
 sg13g2_tielo _884__30 (.L_LO(net30));
 sg13g2_tielo _883__31 (.L_LO(net31));
 sg13g2_tielo _882__32 (.L_LO(net32));
 sg13g2_tielo _881__33 (.L_LO(net33));
 sg13g2_tielo _880__34 (.L_LO(net34));
 sg13g2_tielo _863__35 (.L_LO(net35));
 sg13g2_tielo _862__36 (.L_LO(net36));
 sg13g2_tielo _861__37 (.L_LO(net37));
 sg13g2_tielo _860__38 (.L_LO(net38));
 sg13g2_tielo _859__39 (.L_LO(net39));
 sg13g2_tielo _858__40 (.L_LO(net40));
 sg13g2_tielo _857__41 (.L_LO(net41));
 sg13g2_tielo _856__42 (.L_LO(net42));
 sg13g2_tielo _855__43 (.L_LO(net43));
 sg13g2_tielo _854__44 (.L_LO(net44));
 sg13g2_tielo _853__45 (.L_LO(net45));
 sg13g2_tielo _852__46 (.L_LO(net46));
 sg13g2_tielo _851__47 (.L_LO(net47));
 sg13g2_tielo _850__48 (.L_LO(net48));
 sg13g2_tiehi _883__49 (.L_HI(net49));
 sg13g2_buf_2 fanout87 (.A(net88),
    .X(net87));
 sg13g2_buf_2 fanout88 (.A(_195_),
    .X(net88));
 sg13g2_buf_2 fanout89 (.A(net93),
    .X(net89));
 sg13g2_buf_1 fanout90 (.A(net93),
    .X(net90));
 sg13g2_buf_2 fanout91 (.A(net93),
    .X(net91));
 sg13g2_buf_1 fanout92 (.A(net93),
    .X(net92));
 sg13g2_buf_1 fanout93 (.A(_195_),
    .X(net93));
 sg13g2_buf_2 fanout94 (.A(net95),
    .X(net94));
 sg13g2_buf_2 fanout95 (.A(net98),
    .X(net95));
 sg13g2_buf_2 fanout96 (.A(net97),
    .X(net96));
 sg13g2_buf_2 fanout97 (.A(net98),
    .X(net97));
 sg13g2_buf_1 fanout98 (.A(_195_),
    .X(net98));
 sg13g2_buf_2 fanout99 (.A(net102),
    .X(net99));
 sg13g2_buf_1 fanout100 (.A(net102),
    .X(net100));
 sg13g2_buf_2 fanout101 (.A(net102),
    .X(net101));
 sg13g2_buf_1 fanout102 (.A(uio_in[0]),
    .X(net102));
 sg13g2_buf_4 fanout103 (.X(net103),
    .A(net109));
 sg13g2_buf_4 fanout104 (.X(net104),
    .A(net109));
 sg13g2_buf_4 fanout105 (.X(net105),
    .A(net108));
 sg13g2_buf_2 fanout106 (.A(net108),
    .X(net106));
 sg13g2_buf_4 fanout107 (.X(net107),
    .A(net108));
 sg13g2_buf_4 fanout108 (.X(net108),
    .A(net109));
 sg13g2_buf_2 fanout109 (.A(rst_n),
    .X(net109));
 sg13g2_buf_4 fanout110 (.X(net110),
    .A(net112));
 sg13g2_buf_2 fanout111 (.A(net112),
    .X(net111));
 sg13g2_buf_2 fanout112 (.A(net113),
    .X(net112));
 sg13g2_buf_4 fanout113 (.X(net113),
    .A(net116));
 sg13g2_buf_4 fanout114 (.X(net114),
    .A(net115));
 sg13g2_buf_4 fanout115 (.X(net115),
    .A(net116));
 sg13g2_buf_2 fanout116 (.A(rst_n),
    .X(net116));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[5]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[6]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(ui_in[7]),
    .X(net8));
 sg13g2_buf_2 input9 (.A(uio_in[6]),
    .X(net9));
 sg13g2_buf_2 input10 (.A(uio_in[7]),
    .X(net10));
 sg13g2_tielo tt_um_mroblesh_11 (.L_LO(net11));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_4_1_0_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_4_2_0_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_4_3_0_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_4_4_0_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_4_5_0_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_4_6_0_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_4_7_0_clk));
 sg13g2_inv_1 clkload7 (.A(clknet_4_9_0_clk));
 sg13g2_inv_1 clkload8 (.A(clknet_4_10_0_clk));
 sg13g2_inv_1 clkload9 (.A(clknet_4_11_0_clk));
 sg13g2_inv_1 clkload10 (.A(clknet_4_12_0_clk));
 sg13g2_inv_1 clkload11 (.A(clknet_4_13_0_clk));
 sg13g2_inv_1 clkload12 (.A(clknet_4_14_0_clk));
 sg13g2_inv_1 clkload13 (.A(clknet_4_15_0_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(_033_),
    .X(net75));
 sg13g2_dlygate4sd3_1 hold2 (.A(_042_),
    .X(net76));
 sg13g2_dlygate4sd3_1 hold3 (.A(_091_),
    .X(net77));
 sg13g2_dlygate4sd3_1 hold4 (.A(\decoder_inst.counter[0] ),
    .X(net78));
 sg13g2_dlygate4sd3_1 hold5 (.A(_032_),
    .X(net79));
 sg13g2_dlygate4sd3_1 hold6 (.A(_351_),
    .X(net80));
 sg13g2_dlygate4sd3_1 hold7 (.A(_108_),
    .X(net81));
 sg13g2_dlygate4sd3_1 hold8 (.A(_034_),
    .X(net82));
 sg13g2_dlygate4sd3_1 hold9 (.A(_220_),
    .X(net83));
 sg13g2_dlygate4sd3_1 hold10 (.A(\decoder_inst.freq_out[6] ),
    .X(net84));
 sg13g2_dlygate4sd3_1 hold11 (.A(_089_),
    .X(net85));
 sg13g2_dlygate4sd3_1 hold12 (.A(\decoder_inst.freq_out[4] ),
    .X(net86));
 sg13g2_dlygate4sd3_1 hold13 (.A(_087_),
    .X(net117));
 sg13g2_dlygate4sd3_1 hold14 (.A(\encoder_inst.counter[2] ),
    .X(net118));
 sg13g2_dlygate4sd3_1 hold15 (.A(_341_),
    .X(net119));
 sg13g2_dlygate4sd3_1 hold16 (.A(_093_),
    .X(net120));
 sg13g2_dlygate4sd3_1 hold17 (.A(\decoder_inst.freq_out[7] ),
    .X(net121));
 sg13g2_dlygate4sd3_1 hold18 (.A(_090_),
    .X(net122));
 sg13g2_dlygate4sd3_1 hold19 (.A(\decoder_inst.freq_out[2] ),
    .X(net123));
 sg13g2_dlygate4sd3_1 hold20 (.A(_085_),
    .X(net124));
 sg13g2_dlygate4sd3_1 hold21 (.A(_041_),
    .X(net125));
 sg13g2_dlygate4sd3_1 hold22 (.A(_197_),
    .X(net126));
 sg13g2_dlygate4sd3_1 hold23 (.A(\decoder_inst.freq_out[1] ),
    .X(net127));
 sg13g2_dlygate4sd3_1 hold24 (.A(_084_),
    .X(net128));
 sg13g2_dlygate4sd3_1 hold25 (.A(\decoder_inst.frequency[7] ),
    .X(net129));
 sg13g2_dlygate4sd3_1 hold26 (.A(_241_),
    .X(net130));
 sg13g2_dlygate4sd3_1 hold27 (.A(_058_),
    .X(net131));
 sg13g2_dlygate4sd3_1 hold28 (.A(\decoder_inst.freq_out[3] ),
    .X(net132));
 sg13g2_dlygate4sd3_1 hold29 (.A(_086_),
    .X(net133));
 sg13g2_dlygate4sd3_1 hold30 (.A(\decoder_inst.frequency[30] ),
    .X(net134));
 sg13g2_dlygate4sd3_1 hold31 (.A(_081_),
    .X(net135));
 sg13g2_dlygate4sd3_1 hold32 (.A(\decoder_inst.freq_out[5] ),
    .X(net136));
 sg13g2_dlygate4sd3_1 hold33 (.A(_088_),
    .X(net137));
 sg13g2_dlygate4sd3_1 hold34 (.A(_039_),
    .X(net138));
 sg13g2_dlygate4sd3_1 hold35 (.A(_205_),
    .X(net139));
 sg13g2_dlygate4sd3_1 hold36 (.A(_028_),
    .X(net140));
 sg13g2_dlygate4sd3_1 hold37 (.A(\decoder_inst.freq_out[0] ),
    .X(net141));
 sg13g2_dlygate4sd3_1 hold38 (.A(_083_),
    .X(net142));
 sg13g2_dlygate4sd3_1 hold39 (.A(_035_),
    .X(net143));
 sg13g2_dlygate4sd3_1 hold40 (.A(_215_),
    .X(net144));
 sg13g2_dlygate4sd3_1 hold41 (.A(_037_),
    .X(net145));
 sg13g2_dlygate4sd3_1 hold42 (.A(_209_),
    .X(net146));
 sg13g2_dlygate4sd3_1 hold43 (.A(\decoder_inst.frequency[27] ),
    .X(net147));
 sg13g2_dlygate4sd3_1 hold44 (.A(_284_),
    .X(net148));
 sg13g2_dlygate4sd3_1 hold45 (.A(_078_),
    .X(net149));
 sg13g2_dlygate4sd3_1 hold46 (.A(\decoder_inst.counter[1] ),
    .X(net150));
 sg13g2_dlygate4sd3_1 hold47 (.A(\decoder_inst.frequency[15] ),
    .X(net151));
 sg13g2_dlygate4sd3_1 hold48 (.A(_259_),
    .X(net152));
 sg13g2_dlygate4sd3_1 hold49 (.A(_066_),
    .X(net153));
 sg13g2_dlygate4sd3_1 hold50 (.A(\decoder_inst.counter[3] ),
    .X(net154));
 sg13g2_dlygate4sd3_1 hold51 (.A(_199_),
    .X(net155));
 sg13g2_dlygate4sd3_1 hold52 (.A(_025_),
    .X(net156));
 sg13g2_dlygate4sd3_1 hold53 (.A(\decoder_inst.frequency[19] ),
    .X(net157));
 sg13g2_dlygate4sd3_1 hold54 (.A(_267_),
    .X(net158));
 sg13g2_dlygate4sd3_1 hold55 (.A(_070_),
    .X(net159));
 sg13g2_dlygate4sd3_1 hold56 (.A(\decoder_inst.counter[15] ),
    .X(net160));
 sg13g2_dlygate4sd3_1 hold57 (.A(_223_),
    .X(net161));
 sg13g2_dlygate4sd3_1 hold58 (.A(_006_),
    .X(net162));
 sg13g2_dlygate4sd3_1 hold59 (.A(\decoder_inst.frequency[1] ),
    .X(net163));
 sg13g2_dlygate4sd3_1 hold60 (.A(_230_),
    .X(net164));
 sg13g2_dlygate4sd3_1 hold61 (.A(_052_),
    .X(net165));
 sg13g2_dlygate4sd3_1 hold62 (.A(\decoder_inst.frequency[13] ),
    .X(net166));
 sg13g2_dlygate4sd3_1 hold63 (.A(_254_),
    .X(net167));
 sg13g2_dlygate4sd3_1 hold64 (.A(\decoder_inst.frequency[18] ),
    .X(net168));
 sg13g2_dlygate4sd3_1 hold65 (.A(_266_),
    .X(net169));
 sg13g2_dlygate4sd3_1 hold66 (.A(\decoder_inst.frequency[26] ),
    .X(net170));
 sg13g2_dlygate4sd3_1 hold67 (.A(_282_),
    .X(net171));
 sg13g2_dlygate4sd3_1 hold68 (.A(_077_),
    .X(net172));
 sg13g2_dlygate4sd3_1 hold69 (.A(\decoder_inst.frequency[20] ),
    .X(net173));
 sg13g2_dlygate4sd3_1 hold70 (.A(_269_),
    .X(net174));
 sg13g2_dlygate4sd3_1 hold71 (.A(_071_),
    .X(net175));
 sg13g2_dlygate4sd3_1 hold72 (.A(\decoder_inst.frequency[2] ),
    .X(net176));
 sg13g2_dlygate4sd3_1 hold73 (.A(_232_),
    .X(net177));
 sg13g2_dlygate4sd3_1 hold74 (.A(\decoder_inst.frequency[29] ),
    .X(net178));
 sg13g2_dlygate4sd3_1 hold75 (.A(_288_),
    .X(net179));
 sg13g2_dlygate4sd3_1 hold76 (.A(_080_),
    .X(net180));
 sg13g2_dlygate4sd3_1 hold77 (.A(\encoder_inst.counter[3] ),
    .X(net181));
 sg13g2_dlygate4sd3_1 hold78 (.A(_342_),
    .X(net182));
 sg13g2_dlygate4sd3_1 hold79 (.A(_094_),
    .X(net183));
 sg13g2_dlygate4sd3_1 hold80 (.A(_038_),
    .X(net184));
 sg13g2_dlygate4sd3_1 hold81 (.A(_206_),
    .X(net185));
 sg13g2_dlygate4sd3_1 hold82 (.A(\decoder_inst.frequency[4] ),
    .X(net186));
 sg13g2_dlygate4sd3_1 hold83 (.A(_237_),
    .X(net187));
 sg13g2_dlygate4sd3_1 hold84 (.A(\decoder_inst.frequency[0] ),
    .X(net188));
 sg13g2_dlygate4sd3_1 hold85 (.A(_228_),
    .X(net189));
 sg13g2_dlygate4sd3_1 hold86 (.A(_051_),
    .X(net190));
 sg13g2_dlygate4sd3_1 hold87 (.A(\decoder_inst.frequency[8] ),
    .X(net191));
 sg13g2_dlygate4sd3_1 hold88 (.A(_245_),
    .X(net192));
 sg13g2_dlygate4sd3_1 hold89 (.A(\decoder_inst.frequency[22] ),
    .X(net193));
 sg13g2_dlygate4sd3_1 hold90 (.A(_273_),
    .X(net194));
 sg13g2_dlygate4sd3_1 hold91 (.A(\decoder_inst.frequency[23] ),
    .X(net195));
 sg13g2_dlygate4sd3_1 hold92 (.A(\decoder_inst.frequency[3] ),
    .X(net196));
 sg13g2_dlygate4sd3_1 hold93 (.A(\decoder_inst.frequency[25] ),
    .X(net197));
 sg13g2_dlygate4sd3_1 hold94 (.A(_280_),
    .X(net198));
 sg13g2_dlygate4sd3_1 hold95 (.A(_076_),
    .X(net199));
 sg13g2_dlygate4sd3_1 hold96 (.A(\decoder_inst.counter[14] ),
    .X(net200));
 sg13g2_dlygate4sd3_1 hold97 (.A(_222_),
    .X(net201));
 sg13g2_dlygate4sd3_1 hold98 (.A(_040_),
    .X(net202));
 sg13g2_dlygate4sd3_1 hold99 (.A(_202_),
    .X(net203));
 sg13g2_dlygate4sd3_1 hold100 (.A(\encoder_inst.counter[0] ),
    .X(net204));
 sg13g2_dlygate4sd3_1 hold101 (.A(_339_),
    .X(net205));
 sg13g2_dlygate4sd3_1 hold102 (.A(_092_),
    .X(net206));
 sg13g2_dlygate4sd3_1 hold103 (.A(\decoder_inst.frequency[21] ),
    .X(net207));
 sg13g2_dlygate4sd3_1 hold104 (.A(_271_),
    .X(net208));
 sg13g2_dlygate4sd3_1 hold105 (.A(_072_),
    .X(net209));
 sg13g2_dlygate4sd3_1 hold106 (.A(_036_),
    .X(net210));
 sg13g2_dlygate4sd3_1 hold107 (.A(_213_),
    .X(net211));
 sg13g2_dlygate4sd3_1 hold108 (.A(_001_),
    .X(net212));
 sg13g2_dlygate4sd3_1 hold109 (.A(\decoder_inst.frequency[16] ),
    .X(net213));
 sg13g2_dlygate4sd3_1 hold110 (.A(_260_),
    .X(net214));
 sg13g2_dlygate4sd3_1 hold111 (.A(\decoder_inst.frequency[17] ),
    .X(net215));
 sg13g2_dlygate4sd3_1 hold112 (.A(\decoder_inst.frequency[24] ),
    .X(net216));
 sg13g2_dlygate4sd3_1 hold113 (.A(\decoder_inst.signal_in_prev ),
    .X(net217));
 sg13g2_dlygate4sd3_1 hold114 (.A(\decoder_inst.counter[12] ),
    .X(net218));
 sg13g2_dlygate4sd3_1 hold115 (.A(_219_),
    .X(net219));
 sg13g2_dlygate4sd3_1 hold116 (.A(\decoder_inst.frequency[28] ),
    .X(net220));
 sg13g2_dlygate4sd3_1 hold117 (.A(_286_),
    .X(net221));
 sg13g2_dlygate4sd3_1 hold118 (.A(\decoder_inst.counter[16] ),
    .X(net222));
 sg13g2_dlygate4sd3_1 hold119 (.A(\decoder_inst.frequency[6] ),
    .X(net223));
 sg13g2_dlygate4sd3_1 hold120 (.A(_240_),
    .X(net224));
 sg13g2_dlygate4sd3_1 hold121 (.A(\decoder_inst.counter[4] ),
    .X(net225));
 sg13g2_dlygate4sd3_1 hold122 (.A(_201_),
    .X(net226));
 sg13g2_dlygate4sd3_1 hold123 (.A(\encoder_inst.counter[4] ),
    .X(net227));
 sg13g2_dlygate4sd3_1 hold124 (.A(_095_),
    .X(net228));
 sg13g2_dlygate4sd3_1 hold125 (.A(\decoder_inst.frequency[11] ),
    .X(net229));
 sg13g2_dlygate4sd3_1 hold126 (.A(_252_),
    .X(net230));
 sg13g2_dlygate4sd3_1 hold127 (.A(\decoder_inst.frequency[14] ),
    .X(net231));
 sg13g2_dlygate4sd3_1 hold128 (.A(_257_),
    .X(net232));
 sg13g2_dlygate4sd3_1 hold129 (.A(\decoder_inst.frequency[9] ),
    .X(net233));
 sg13g2_dlygate4sd3_1 hold130 (.A(_246_),
    .X(net234));
 sg13g2_dlygate4sd3_1 hold131 (.A(\decoder_inst.frequency[31] ),
    .X(net235));
 sg13g2_dlygate4sd3_1 hold132 (.A(\decoder_inst.frequency[12] ),
    .X(net236));
 sg13g2_dlygate4sd3_1 hold133 (.A(_253_),
    .X(net237));
 sg13g2_dlygate4sd3_1 hold134 (.A(\decoder_inst.counter[9] ),
    .X(net238));
 sg13g2_dlygate4sd3_1 hold135 (.A(_210_),
    .X(net239));
 sg13g2_dlygate4sd3_1 hold136 (.A(_212_),
    .X(net240));
 sg13g2_dlygate4sd3_1 hold137 (.A(\encoder_inst.counter[7] ),
    .X(net241));
 sg13g2_dlygate4sd3_1 hold138 (.A(_349_),
    .X(net242));
 sg13g2_dlygate4sd3_1 hold139 (.A(_098_),
    .X(net243));
 sg13g2_dlygate4sd3_1 hold140 (.A(\decoder_inst.frequency[10] ),
    .X(net244));
 sg13g2_dlygate4sd3_1 hold141 (.A(\encoder_inst.counter[5] ),
    .X(net245));
 sg13g2_dlygate4sd3_1 hold142 (.A(_096_),
    .X(net246));
 sg13g2_dlygate4sd3_1 hold143 (.A(\encoder_inst.counter[6] ),
    .X(net247));
 sg13g2_dlygate4sd3_1 hold144 (.A(_097_),
    .X(net248));
 sg13g2_dlygate4sd3_1 hold145 (.A(\decoder_inst.frequency[5] ),
    .X(net249));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_fill_2 FILLER_14_406 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_252 ();
 sg13g2_decap_8 FILLER_15_259 ();
 sg13g2_decap_8 FILLER_15_266 ();
 sg13g2_decap_8 FILLER_15_273 ();
 sg13g2_decap_8 FILLER_15_280 ();
 sg13g2_decap_8 FILLER_15_287 ();
 sg13g2_decap_8 FILLER_15_294 ();
 sg13g2_decap_8 FILLER_15_301 ();
 sg13g2_decap_8 FILLER_15_308 ();
 sg13g2_decap_8 FILLER_15_315 ();
 sg13g2_decap_8 FILLER_15_322 ();
 sg13g2_decap_8 FILLER_15_329 ();
 sg13g2_decap_8 FILLER_15_336 ();
 sg13g2_decap_8 FILLER_15_343 ();
 sg13g2_decap_8 FILLER_15_350 ();
 sg13g2_decap_8 FILLER_15_357 ();
 sg13g2_decap_8 FILLER_15_364 ();
 sg13g2_decap_8 FILLER_15_371 ();
 sg13g2_decap_8 FILLER_15_378 ();
 sg13g2_decap_8 FILLER_15_385 ();
 sg13g2_decap_8 FILLER_15_392 ();
 sg13g2_decap_8 FILLER_15_399 ();
 sg13g2_fill_2 FILLER_15_406 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_decap_8 FILLER_16_217 ();
 sg13g2_decap_8 FILLER_16_224 ();
 sg13g2_decap_8 FILLER_16_231 ();
 sg13g2_decap_8 FILLER_16_238 ();
 sg13g2_decap_8 FILLER_16_245 ();
 sg13g2_decap_8 FILLER_16_252 ();
 sg13g2_decap_8 FILLER_16_259 ();
 sg13g2_decap_8 FILLER_16_266 ();
 sg13g2_decap_8 FILLER_16_273 ();
 sg13g2_decap_8 FILLER_16_280 ();
 sg13g2_decap_8 FILLER_16_287 ();
 sg13g2_decap_8 FILLER_16_294 ();
 sg13g2_decap_8 FILLER_16_301 ();
 sg13g2_decap_8 FILLER_16_308 ();
 sg13g2_decap_8 FILLER_16_315 ();
 sg13g2_decap_8 FILLER_16_322 ();
 sg13g2_decap_8 FILLER_16_329 ();
 sg13g2_decap_8 FILLER_16_336 ();
 sg13g2_decap_8 FILLER_16_343 ();
 sg13g2_decap_8 FILLER_16_350 ();
 sg13g2_decap_8 FILLER_16_357 ();
 sg13g2_decap_8 FILLER_16_364 ();
 sg13g2_decap_8 FILLER_16_371 ();
 sg13g2_decap_8 FILLER_16_378 ();
 sg13g2_decap_8 FILLER_16_385 ();
 sg13g2_decap_8 FILLER_16_392 ();
 sg13g2_decap_8 FILLER_16_399 ();
 sg13g2_fill_2 FILLER_16_406 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_decap_8 FILLER_17_168 ();
 sg13g2_decap_8 FILLER_17_175 ();
 sg13g2_decap_8 FILLER_17_182 ();
 sg13g2_decap_8 FILLER_17_189 ();
 sg13g2_decap_8 FILLER_17_196 ();
 sg13g2_decap_8 FILLER_17_203 ();
 sg13g2_decap_8 FILLER_17_210 ();
 sg13g2_decap_8 FILLER_17_217 ();
 sg13g2_decap_8 FILLER_17_224 ();
 sg13g2_decap_8 FILLER_17_231 ();
 sg13g2_decap_8 FILLER_17_238 ();
 sg13g2_decap_8 FILLER_17_245 ();
 sg13g2_decap_8 FILLER_17_252 ();
 sg13g2_decap_8 FILLER_17_259 ();
 sg13g2_decap_8 FILLER_17_266 ();
 sg13g2_decap_8 FILLER_17_273 ();
 sg13g2_decap_8 FILLER_17_280 ();
 sg13g2_decap_8 FILLER_17_287 ();
 sg13g2_decap_8 FILLER_17_294 ();
 sg13g2_decap_8 FILLER_17_301 ();
 sg13g2_decap_8 FILLER_17_308 ();
 sg13g2_decap_8 FILLER_17_315 ();
 sg13g2_decap_8 FILLER_17_322 ();
 sg13g2_decap_8 FILLER_17_329 ();
 sg13g2_decap_8 FILLER_17_336 ();
 sg13g2_decap_8 FILLER_17_343 ();
 sg13g2_decap_8 FILLER_17_350 ();
 sg13g2_decap_8 FILLER_17_357 ();
 sg13g2_decap_8 FILLER_17_364 ();
 sg13g2_decap_8 FILLER_17_371 ();
 sg13g2_decap_8 FILLER_17_378 ();
 sg13g2_decap_8 FILLER_17_385 ();
 sg13g2_decap_8 FILLER_17_392 ();
 sg13g2_decap_8 FILLER_17_399 ();
 sg13g2_fill_2 FILLER_17_406 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_decap_8 FILLER_18_147 ();
 sg13g2_decap_8 FILLER_18_154 ();
 sg13g2_decap_8 FILLER_18_161 ();
 sg13g2_decap_8 FILLER_18_168 ();
 sg13g2_decap_8 FILLER_18_175 ();
 sg13g2_decap_8 FILLER_18_182 ();
 sg13g2_decap_8 FILLER_18_189 ();
 sg13g2_decap_8 FILLER_18_196 ();
 sg13g2_decap_8 FILLER_18_203 ();
 sg13g2_decap_8 FILLER_18_210 ();
 sg13g2_decap_8 FILLER_18_217 ();
 sg13g2_decap_4 FILLER_18_224 ();
 sg13g2_fill_2 FILLER_18_228 ();
 sg13g2_decap_8 FILLER_18_238 ();
 sg13g2_decap_8 FILLER_18_245 ();
 sg13g2_decap_8 FILLER_18_252 ();
 sg13g2_decap_8 FILLER_18_264 ();
 sg13g2_decap_8 FILLER_18_271 ();
 sg13g2_decap_8 FILLER_18_278 ();
 sg13g2_decap_8 FILLER_18_285 ();
 sg13g2_decap_8 FILLER_18_292 ();
 sg13g2_fill_1 FILLER_18_299 ();
 sg13g2_fill_2 FILLER_18_326 ();
 sg13g2_decap_8 FILLER_18_362 ();
 sg13g2_decap_8 FILLER_18_369 ();
 sg13g2_decap_8 FILLER_18_376 ();
 sg13g2_decap_8 FILLER_18_383 ();
 sg13g2_decap_8 FILLER_18_390 ();
 sg13g2_decap_8 FILLER_18_397 ();
 sg13g2_decap_4 FILLER_18_404 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_decap_8 FILLER_19_140 ();
 sg13g2_decap_8 FILLER_19_147 ();
 sg13g2_decap_8 FILLER_19_154 ();
 sg13g2_decap_8 FILLER_19_161 ();
 sg13g2_decap_8 FILLER_19_168 ();
 sg13g2_decap_8 FILLER_19_175 ();
 sg13g2_decap_8 FILLER_19_182 ();
 sg13g2_decap_8 FILLER_19_189 ();
 sg13g2_fill_2 FILLER_19_196 ();
 sg13g2_decap_4 FILLER_19_224 ();
 sg13g2_fill_1 FILLER_19_228 ();
 sg13g2_fill_2 FILLER_19_238 ();
 sg13g2_fill_1 FILLER_19_240 ();
 sg13g2_decap_4 FILLER_19_250 ();
 sg13g2_fill_2 FILLER_19_259 ();
 sg13g2_fill_2 FILLER_19_270 ();
 sg13g2_decap_8 FILLER_19_281 ();
 sg13g2_decap_8 FILLER_19_288 ();
 sg13g2_decap_4 FILLER_19_295 ();
 sg13g2_fill_2 FILLER_19_299 ();
 sg13g2_fill_2 FILLER_19_327 ();
 sg13g2_decap_8 FILLER_19_363 ();
 sg13g2_decap_4 FILLER_19_370 ();
 sg13g2_fill_2 FILLER_19_374 ();
 sg13g2_decap_8 FILLER_19_402 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_fill_1 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_103 ();
 sg13g2_decap_8 FILLER_20_110 ();
 sg13g2_decap_8 FILLER_20_117 ();
 sg13g2_decap_8 FILLER_20_124 ();
 sg13g2_decap_8 FILLER_20_131 ();
 sg13g2_decap_8 FILLER_20_138 ();
 sg13g2_decap_8 FILLER_20_145 ();
 sg13g2_decap_8 FILLER_20_152 ();
 sg13g2_decap_8 FILLER_20_159 ();
 sg13g2_decap_8 FILLER_20_166 ();
 sg13g2_decap_8 FILLER_20_173 ();
 sg13g2_decap_8 FILLER_20_180 ();
 sg13g2_decap_4 FILLER_20_187 ();
 sg13g2_fill_2 FILLER_20_191 ();
 sg13g2_fill_1 FILLER_20_211 ();
 sg13g2_fill_2 FILLER_20_221 ();
 sg13g2_decap_4 FILLER_20_286 ();
 sg13g2_fill_1 FILLER_20_290 ();
 sg13g2_decap_8 FILLER_20_295 ();
 sg13g2_decap_8 FILLER_20_310 ();
 sg13g2_fill_1 FILLER_20_317 ();
 sg13g2_decap_8 FILLER_20_322 ();
 sg13g2_decap_8 FILLER_20_329 ();
 sg13g2_decap_4 FILLER_20_336 ();
 sg13g2_fill_1 FILLER_20_340 ();
 sg13g2_decap_4 FILLER_20_367 ();
 sg13g2_fill_1 FILLER_20_371 ();
 sg13g2_decap_8 FILLER_20_402 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_fill_1 FILLER_21_77 ();
 sg13g2_fill_2 FILLER_21_87 ();
 sg13g2_fill_1 FILLER_21_89 ();
 sg13g2_fill_2 FILLER_21_95 ();
 sg13g2_fill_2 FILLER_21_106 ();
 sg13g2_fill_2 FILLER_21_125 ();
 sg13g2_fill_1 FILLER_21_127 ();
 sg13g2_decap_8 FILLER_21_132 ();
 sg13g2_decap_8 FILLER_21_139 ();
 sg13g2_decap_8 FILLER_21_146 ();
 sg13g2_decap_8 FILLER_21_153 ();
 sg13g2_decap_8 FILLER_21_160 ();
 sg13g2_decap_8 FILLER_21_167 ();
 sg13g2_decap_4 FILLER_21_174 ();
 sg13g2_fill_1 FILLER_21_178 ();
 sg13g2_fill_2 FILLER_21_238 ();
 sg13g2_fill_2 FILLER_21_257 ();
 sg13g2_fill_2 FILLER_21_313 ();
 sg13g2_fill_1 FILLER_21_315 ();
 sg13g2_fill_1 FILLER_21_342 ();
 sg13g2_decap_8 FILLER_21_347 ();
 sg13g2_fill_2 FILLER_21_354 ();
 sg13g2_fill_1 FILLER_21_356 ();
 sg13g2_decap_8 FILLER_21_362 ();
 sg13g2_fill_2 FILLER_21_369 ();
 sg13g2_fill_1 FILLER_21_371 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_4 FILLER_22_49 ();
 sg13g2_fill_2 FILLER_22_53 ();
 sg13g2_fill_2 FILLER_22_143 ();
 sg13g2_fill_1 FILLER_22_145 ();
 sg13g2_decap_8 FILLER_22_159 ();
 sg13g2_decap_8 FILLER_22_166 ();
 sg13g2_decap_8 FILLER_22_173 ();
 sg13g2_decap_8 FILLER_22_180 ();
 sg13g2_decap_8 FILLER_22_187 ();
 sg13g2_decap_4 FILLER_22_194 ();
 sg13g2_fill_1 FILLER_22_198 ();
 sg13g2_fill_2 FILLER_22_247 ();
 sg13g2_fill_1 FILLER_22_265 ();
 sg13g2_fill_1 FILLER_22_294 ();
 sg13g2_fill_2 FILLER_22_330 ();
 sg13g2_fill_1 FILLER_22_340 ();
 sg13g2_fill_2 FILLER_22_372 ();
 sg13g2_decap_8 FILLER_22_400 ();
 sg13g2_fill_2 FILLER_22_407 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_fill_1 FILLER_23_63 ();
 sg13g2_fill_1 FILLER_23_77 ();
 sg13g2_fill_1 FILLER_23_94 ();
 sg13g2_fill_2 FILLER_23_254 ();
 sg13g2_fill_2 FILLER_23_272 ();
 sg13g2_fill_2 FILLER_23_325 ();
 sg13g2_decap_8 FILLER_23_353 ();
 sg13g2_decap_8 FILLER_23_366 ();
 sg13g2_fill_2 FILLER_23_373 ();
 sg13g2_decap_8 FILLER_23_383 ();
 sg13g2_decap_8 FILLER_23_390 ();
 sg13g2_decap_8 FILLER_23_397 ();
 sg13g2_decap_4 FILLER_23_404 ();
 sg13g2_fill_1 FILLER_23_408 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_4 FILLER_24_49 ();
 sg13g2_fill_1 FILLER_24_53 ();
 sg13g2_fill_1 FILLER_24_101 ();
 sg13g2_fill_1 FILLER_24_128 ();
 sg13g2_fill_2 FILLER_24_190 ();
 sg13g2_decap_4 FILLER_24_333 ();
 sg13g2_fill_1 FILLER_24_337 ();
 sg13g2_decap_8 FILLER_24_346 ();
 sg13g2_fill_2 FILLER_24_353 ();
 sg13g2_decap_8 FILLER_24_384 ();
 sg13g2_decap_8 FILLER_24_391 ();
 sg13g2_decap_8 FILLER_24_398 ();
 sg13g2_decap_4 FILLER_24_405 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_fill_2 FILLER_25_49 ();
 sg13g2_fill_2 FILLER_25_92 ();
 sg13g2_fill_1 FILLER_25_121 ();
 sg13g2_fill_1 FILLER_25_195 ();
 sg13g2_fill_1 FILLER_25_229 ();
 sg13g2_decap_4 FILLER_25_233 ();
 sg13g2_fill_1 FILLER_25_247 ();
 sg13g2_decap_4 FILLER_25_257 ();
 sg13g2_fill_1 FILLER_25_261 ();
 sg13g2_fill_2 FILLER_25_267 ();
 sg13g2_fill_1 FILLER_25_269 ();
 sg13g2_fill_2 FILLER_25_304 ();
 sg13g2_fill_2 FILLER_25_326 ();
 sg13g2_fill_1 FILLER_25_328 ();
 sg13g2_fill_1 FILLER_25_363 ();
 sg13g2_decap_8 FILLER_25_378 ();
 sg13g2_decap_8 FILLER_25_385 ();
 sg13g2_decap_8 FILLER_25_392 ();
 sg13g2_decap_8 FILLER_25_399 ();
 sg13g2_fill_2 FILLER_25_406 ();
 sg13g2_fill_1 FILLER_25_408 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_fill_1 FILLER_26_49 ();
 sg13g2_fill_1 FILLER_26_100 ();
 sg13g2_fill_1 FILLER_26_111 ();
 sg13g2_fill_2 FILLER_26_157 ();
 sg13g2_fill_1 FILLER_26_177 ();
 sg13g2_fill_2 FILLER_26_183 ();
 sg13g2_decap_4 FILLER_26_260 ();
 sg13g2_fill_1 FILLER_26_264 ();
 sg13g2_fill_1 FILLER_26_305 ();
 sg13g2_decap_8 FILLER_26_332 ();
 sg13g2_decap_8 FILLER_26_339 ();
 sg13g2_decap_8 FILLER_26_346 ();
 sg13g2_decap_8 FILLER_26_353 ();
 sg13g2_fill_2 FILLER_26_363 ();
 sg13g2_fill_1 FILLER_26_365 ();
 sg13g2_fill_1 FILLER_26_392 ();
 sg13g2_decap_8 FILLER_26_397 ();
 sg13g2_fill_1 FILLER_26_408 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_4 FILLER_27_35 ();
 sg13g2_fill_1 FILLER_27_39 ();
 sg13g2_fill_2 FILLER_27_107 ();
 sg13g2_fill_1 FILLER_27_135 ();
 sg13g2_fill_2 FILLER_27_180 ();
 sg13g2_fill_1 FILLER_27_182 ();
 sg13g2_fill_1 FILLER_27_188 ();
 sg13g2_fill_2 FILLER_27_253 ();
 sg13g2_fill_1 FILLER_27_255 ();
 sg13g2_decap_8 FILLER_27_278 ();
 sg13g2_decap_4 FILLER_27_285 ();
 sg13g2_fill_2 FILLER_27_289 ();
 sg13g2_fill_1 FILLER_27_312 ();
 sg13g2_fill_2 FILLER_27_348 ();
 sg13g2_decap_8 FILLER_27_354 ();
 sg13g2_decap_4 FILLER_27_361 ();
 sg13g2_fill_2 FILLER_27_365 ();
 sg13g2_fill_1 FILLER_27_371 ();
 sg13g2_fill_2 FILLER_27_406 ();
 sg13g2_fill_1 FILLER_27_408 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_fill_2 FILLER_28_42 ();
 sg13g2_fill_1 FILLER_28_44 ();
 sg13g2_fill_2 FILLER_28_114 ();
 sg13g2_fill_2 FILLER_28_125 ();
 sg13g2_decap_8 FILLER_28_183 ();
 sg13g2_decap_4 FILLER_28_190 ();
 sg13g2_fill_1 FILLER_28_194 ();
 sg13g2_decap_4 FILLER_28_199 ();
 sg13g2_fill_1 FILLER_28_217 ();
 sg13g2_fill_2 FILLER_28_257 ();
 sg13g2_decap_4 FILLER_28_278 ();
 sg13g2_fill_1 FILLER_28_282 ();
 sg13g2_decap_4 FILLER_28_300 ();
 sg13g2_fill_2 FILLER_28_304 ();
 sg13g2_fill_1 FILLER_28_366 ();
 sg13g2_fill_2 FILLER_28_375 ();
 sg13g2_fill_1 FILLER_28_377 ();
 sg13g2_fill_1 FILLER_28_408 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_fill_2 FILLER_29_49 ();
 sg13g2_fill_2 FILLER_29_252 ();
 sg13g2_fill_2 FILLER_29_259 ();
 sg13g2_fill_1 FILLER_29_277 ();
 sg13g2_decap_4 FILLER_29_312 ();
 sg13g2_fill_1 FILLER_29_316 ();
 sg13g2_decap_8 FILLER_29_321 ();
 sg13g2_decap_8 FILLER_29_328 ();
 sg13g2_fill_2 FILLER_29_339 ();
 sg13g2_fill_2 FILLER_29_345 ();
 sg13g2_fill_1 FILLER_29_347 ();
 sg13g2_fill_2 FILLER_29_354 ();
 sg13g2_fill_2 FILLER_29_407 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_fill_1 FILLER_30_42 ();
 sg13g2_fill_2 FILLER_30_111 ();
 sg13g2_fill_2 FILLER_30_127 ();
 sg13g2_fill_2 FILLER_30_160 ();
 sg13g2_fill_2 FILLER_30_175 ();
 sg13g2_fill_1 FILLER_30_191 ();
 sg13g2_fill_2 FILLER_30_201 ();
 sg13g2_fill_2 FILLER_30_284 ();
 sg13g2_fill_1 FILLER_30_286 ();
 sg13g2_decap_8 FILLER_30_304 ();
 sg13g2_decap_8 FILLER_30_311 ();
 sg13g2_fill_2 FILLER_30_318 ();
 sg13g2_fill_1 FILLER_30_350 ();
 sg13g2_fill_2 FILLER_30_378 ();
 sg13g2_fill_2 FILLER_30_406 ();
 sg13g2_fill_1 FILLER_30_408 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_4 FILLER_31_42 ();
 sg13g2_fill_2 FILLER_31_99 ();
 sg13g2_fill_1 FILLER_31_113 ();
 sg13g2_fill_1 FILLER_31_154 ();
 sg13g2_fill_1 FILLER_31_190 ();
 sg13g2_fill_1 FILLER_31_260 ();
 sg13g2_fill_1 FILLER_31_266 ();
 sg13g2_fill_2 FILLER_31_297 ();
 sg13g2_fill_1 FILLER_31_299 ();
 sg13g2_fill_1 FILLER_31_408 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_fill_2 FILLER_32_49 ();
 sg13g2_fill_1 FILLER_32_51 ();
 sg13g2_fill_2 FILLER_32_90 ();
 sg13g2_fill_1 FILLER_32_131 ();
 sg13g2_fill_1 FILLER_32_141 ();
 sg13g2_fill_2 FILLER_32_297 ();
 sg13g2_decap_8 FILLER_32_304 ();
 sg13g2_fill_2 FILLER_32_315 ();
 sg13g2_decap_4 FILLER_32_322 ();
 sg13g2_fill_1 FILLER_32_340 ();
 sg13g2_fill_1 FILLER_32_367 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_fill_1 FILLER_33_56 ();
 sg13g2_fill_2 FILLER_33_177 ();
 sg13g2_fill_1 FILLER_33_268 ();
 sg13g2_fill_2 FILLER_33_341 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_fill_2 FILLER_34_63 ();
 sg13g2_fill_2 FILLER_34_108 ();
 sg13g2_fill_2 FILLER_34_127 ();
 sg13g2_fill_2 FILLER_34_184 ();
 sg13g2_fill_2 FILLER_34_221 ();
 sg13g2_fill_1 FILLER_34_352 ();
 sg13g2_fill_2 FILLER_34_363 ();
 sg13g2_fill_1 FILLER_34_408 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_fill_2 FILLER_35_70 ();
 sg13g2_fill_1 FILLER_35_85 ();
 sg13g2_fill_1 FILLER_35_109 ();
 sg13g2_fill_1 FILLER_35_119 ();
 sg13g2_fill_1 FILLER_35_134 ();
 sg13g2_fill_2 FILLER_35_157 ();
 sg13g2_fill_1 FILLER_35_215 ();
 sg13g2_fill_1 FILLER_35_252 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_fill_2 FILLER_36_77 ();
 sg13g2_fill_1 FILLER_36_79 ();
 sg13g2_fill_2 FILLER_36_241 ();
 sg13g2_fill_2 FILLER_36_305 ();
 sg13g2_fill_2 FILLER_36_382 ();
 sg13g2_fill_2 FILLER_36_407 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_fill_2 FILLER_37_70 ();
 sg13g2_fill_1 FILLER_37_119 ();
 sg13g2_fill_2 FILLER_37_255 ();
 sg13g2_fill_1 FILLER_37_292 ();
 sg13g2_fill_1 FILLER_37_337 ();
 sg13g2_fill_1 FILLER_37_355 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_fill_2 FILLER_38_60 ();
 sg13g2_fill_1 FILLER_38_62 ();
 sg13g2_fill_1 FILLER_38_112 ();
 sg13g2_fill_2 FILLER_38_147 ();
 sg13g2_fill_2 FILLER_38_190 ();
 sg13g2_fill_2 FILLER_38_197 ();
 sg13g2_fill_2 FILLER_38_213 ();
 sg13g2_fill_1 FILLER_38_234 ();
 sg13g2_fill_2 FILLER_38_265 ();
 sg13g2_fill_1 FILLER_38_325 ();
 assign uio_oe[0] = net11;
 assign uio_oe[1] = net12;
 assign uio_oe[2] = net13;
 assign uio_oe[3] = net14;
 assign uio_oe[4] = net15;
 assign uio_oe[5] = net16;
 assign uio_oe[6] = net17;
 assign uio_oe[7] = net18;
 assign uio_out[0] = net19;
 assign uio_out[1] = net20;
 assign uio_out[2] = net21;
 assign uio_out[3] = net22;
 assign uio_out[4] = net23;
 assign uio_out[5] = net24;
 assign uio_out[6] = net25;
 assign uio_out[7] = net26;
endmodule

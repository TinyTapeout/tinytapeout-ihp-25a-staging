module tt_um_yuri_panchul_sea_battle_vga_game (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire clknet_leaf_0_clk;
 wire hsync;
 wire \i_game_and_vga.display_on ;
 wire \i_game_and_vga.i_game_top.collision ;
 wire \i_game_and_vga.i_game_top.end_of_game_timer_running ;
 wire \i_game_and_vga.i_game_top.end_of_game_timer_start ;
 wire \i_game_and_vga.i_game_top.game_won ;
 wire \i_game_and_vga.i_game_top.master_fsm.d_end_of_game_timer_start ;
 wire \i_game_and_vga.i_game_top.master_fsm.d_sprite_target_enable_update ;
 wire \i_game_and_vga.i_game_top.master_fsm.d_sprite_target_write_dxy ;
 wire \i_game_and_vga.i_game_top.master_fsm.d_sprite_torpedo_enable_update ;
 wire \i_game_and_vga.i_game_top.master_fsm.sprite_target_enable_update ;
 wire \i_game_and_vga.i_game_top.master_fsm.sprite_target_within_screen ;
 wire \i_game_and_vga.i_game_top.master_fsm.sprite_target_write_dxy ;
 wire \i_game_and_vga.i_game_top.master_fsm.sprite_torpedo_enable_update ;
 wire \i_game_and_vga.i_game_top.master_fsm.sprite_torpedo_within_screen ;
 wire \i_game_and_vga.i_game_top.master_fsm.state[0] ;
 wire \i_game_and_vga.i_game_top.master_fsm.state[1] ;
 wire \i_game_and_vga.i_game_top.mixer.random ;
 wire \i_game_and_vga.i_game_top.mixer.sprite_target_rgb[0] ;
 wire \i_game_and_vga.i_game_top.mixer.sprite_target_rgb[1] ;
 wire \i_game_and_vga.i_game_top.mixer.sprite_target_rgb[2] ;
 wire \i_game_and_vga.i_game_top.mixer.sprite_target_rgb_en ;
 wire \i_game_and_vga.i_game_top.mixer.sprite_torpedo_rgb[1] ;
 wire \i_game_and_vga.i_game_top.mixer.sprite_torpedo_rgb[2] ;
 wire \i_game_and_vga.i_game_top.mixer.sprite_torpedo_rgb_en ;
 wire \i_game_and_vga.i_game_top.overlap.bottom_1[0] ;
 wire \i_game_and_vga.i_game_top.overlap.bottom_1[1] ;
 wire \i_game_and_vga.i_game_top.overlap.bottom_1[2] ;
 wire \i_game_and_vga.i_game_top.overlap.bottom_1[3] ;
 wire \i_game_and_vga.i_game_top.overlap.bottom_1[4] ;
 wire \i_game_and_vga.i_game_top.overlap.bottom_1[5] ;
 wire \i_game_and_vga.i_game_top.overlap.bottom_1[6] ;
 wire \i_game_and_vga.i_game_top.overlap.bottom_1[7] ;
 wire \i_game_and_vga.i_game_top.overlap.bottom_2[0] ;
 wire \i_game_and_vga.i_game_top.overlap.bottom_2[1] ;
 wire \i_game_and_vga.i_game_top.overlap.bottom_2[2] ;
 wire \i_game_and_vga.i_game_top.overlap.bottom_2[3] ;
 wire \i_game_and_vga.i_game_top.overlap.bottom_2[4] ;
 wire \i_game_and_vga.i_game_top.overlap.bottom_2[5] ;
 wire \i_game_and_vga.i_game_top.overlap.bottom_2[6] ;
 wire \i_game_and_vga.i_game_top.overlap.bottom_2[7] ;
 wire \i_game_and_vga.i_game_top.overlap.bottom_2[8] ;
 wire \i_game_and_vga.i_game_top.overlap.left_1[0] ;
 wire \i_game_and_vga.i_game_top.overlap.left_1[1] ;
 wire \i_game_and_vga.i_game_top.overlap.left_1[2] ;
 wire \i_game_and_vga.i_game_top.overlap.left_1[3] ;
 wire \i_game_and_vga.i_game_top.overlap.left_1[4] ;
 wire \i_game_and_vga.i_game_top.overlap.left_1[5] ;
 wire \i_game_and_vga.i_game_top.overlap.left_1[6] ;
 wire \i_game_and_vga.i_game_top.overlap.left_1[7] ;
 wire \i_game_and_vga.i_game_top.overlap.left_1[8] ;
 wire \i_game_and_vga.i_game_top.overlap.left_1[9] ;
 wire \i_game_and_vga.i_game_top.overlap.left_2[0] ;
 wire \i_game_and_vga.i_game_top.overlap.left_2[1] ;
 wire \i_game_and_vga.i_game_top.overlap.left_2[2] ;
 wire \i_game_and_vga.i_game_top.overlap.left_2[3] ;
 wire \i_game_and_vga.i_game_top.overlap.left_2[4] ;
 wire \i_game_and_vga.i_game_top.overlap.left_2[5] ;
 wire \i_game_and_vga.i_game_top.overlap.left_2[6] ;
 wire \i_game_and_vga.i_game_top.overlap.left_2[7] ;
 wire \i_game_and_vga.i_game_top.overlap.left_2[8] ;
 wire \i_game_and_vga.i_game_top.overlap.left_2[9] ;
 wire \i_game_and_vga.i_game_top.overlap.right_1[0] ;
 wire \i_game_and_vga.i_game_top.overlap.right_1[1] ;
 wire \i_game_and_vga.i_game_top.overlap.right_1[2] ;
 wire \i_game_and_vga.i_game_top.overlap.right_1[3] ;
 wire \i_game_and_vga.i_game_top.overlap.right_1[4] ;
 wire \i_game_and_vga.i_game_top.overlap.right_1[5] ;
 wire \i_game_and_vga.i_game_top.overlap.right_1[6] ;
 wire \i_game_and_vga.i_game_top.overlap.right_1[7] ;
 wire \i_game_and_vga.i_game_top.overlap.right_1[8] ;
 wire \i_game_and_vga.i_game_top.overlap.right_1[9] ;
 wire \i_game_and_vga.i_game_top.overlap.right_2[0] ;
 wire \i_game_and_vga.i_game_top.overlap.right_2[1] ;
 wire \i_game_and_vga.i_game_top.overlap.right_2[2] ;
 wire \i_game_and_vga.i_game_top.overlap.right_2[3] ;
 wire \i_game_and_vga.i_game_top.overlap.right_2[4] ;
 wire \i_game_and_vga.i_game_top.overlap.right_2[5] ;
 wire \i_game_and_vga.i_game_top.overlap.right_2[6] ;
 wire \i_game_and_vga.i_game_top.overlap.right_2[7] ;
 wire \i_game_and_vga.i_game_top.overlap.right_2[8] ;
 wire \i_game_and_vga.i_game_top.overlap.right_2[9] ;
 wire \i_game_and_vga.i_game_top.overlap.top_1[0] ;
 wire \i_game_and_vga.i_game_top.overlap.top_1[1] ;
 wire \i_game_and_vga.i_game_top.overlap.top_1[2] ;
 wire \i_game_and_vga.i_game_top.overlap.top_1[3] ;
 wire \i_game_and_vga.i_game_top.overlap.top_1[4] ;
 wire \i_game_and_vga.i_game_top.overlap.top_1[5] ;
 wire \i_game_and_vga.i_game_top.overlap.top_1[6] ;
 wire \i_game_and_vga.i_game_top.overlap.top_2[0] ;
 wire \i_game_and_vga.i_game_top.overlap.top_2[1] ;
 wire \i_game_and_vga.i_game_top.overlap.top_2[2] ;
 wire \i_game_and_vga.i_game_top.overlap.top_2[3] ;
 wire \i_game_and_vga.i_game_top.overlap.top_2[4] ;
 wire \i_game_and_vga.i_game_top.overlap.top_2[5] ;
 wire \i_game_and_vga.i_game_top.overlap.top_2[6] ;
 wire \i_game_and_vga.i_game_top.overlap.top_2[7] ;
 wire \i_game_and_vga.i_game_top.overlap.top_2[8] ;
 wire \i_game_and_vga.i_game_top.random[10] ;
 wire \i_game_and_vga.i_game_top.random[11] ;
 wire \i_game_and_vga.i_game_top.random[12] ;
 wire \i_game_and_vga.i_game_top.random[13] ;
 wire \i_game_and_vga.i_game_top.random[14] ;
 wire \i_game_and_vga.i_game_top.random[15] ;
 wire \i_game_and_vga.i_game_top.random[1] ;
 wire \i_game_and_vga.i_game_top.random[2] ;
 wire \i_game_and_vga.i_game_top.random[3] ;
 wire \i_game_and_vga.i_game_top.random[4] ;
 wire \i_game_and_vga.i_game_top.random[5] ;
 wire \i_game_and_vga.i_game_top.random[6] ;
 wire \i_game_and_vga.i_game_top.random[7] ;
 wire \i_game_and_vga.i_game_top.random[8] ;
 wire \i_game_and_vga.i_game_top.random[9] ;
 wire \i_game_and_vga.i_game_top.sprite_target.pixel_x[0] ;
 wire \i_game_and_vga.i_game_top.sprite_target.pixel_x[1] ;
 wire \i_game_and_vga.i_game_top.sprite_target.pixel_x[2] ;
 wire \i_game_and_vga.i_game_top.sprite_target.pixel_x[3] ;
 wire \i_game_and_vga.i_game_top.sprite_target.pixel_x[4] ;
 wire \i_game_and_vga.i_game_top.sprite_target.pixel_x[5] ;
 wire \i_game_and_vga.i_game_top.sprite_target.pixel_x[6] ;
 wire \i_game_and_vga.i_game_top.sprite_target.pixel_x[7] ;
 wire \i_game_and_vga.i_game_top.sprite_target.pixel_x[8] ;
 wire \i_game_and_vga.i_game_top.sprite_target.pixel_x[9] ;
 wire \i_game_and_vga.i_game_top.sprite_target.pixel_y[0] ;
 wire \i_game_and_vga.i_game_top.sprite_target.pixel_y[1] ;
 wire \i_game_and_vga.i_game_top.sprite_target.pixel_y[2] ;
 wire \i_game_and_vga.i_game_top.sprite_target.pixel_y[3] ;
 wire \i_game_and_vga.i_game_top.sprite_target.pixel_y[4] ;
 wire \i_game_and_vga.i_game_top.sprite_target.pixel_y[5] ;
 wire \i_game_and_vga.i_game_top.sprite_target.pixel_y[6] ;
 wire \i_game_and_vga.i_game_top.sprite_target.pixel_y[7] ;
 wire \i_game_and_vga.i_game_top.sprite_target.pixel_y[8] ;
 wire \i_game_and_vga.i_game_top.sprite_target.sprite_control.dx[0] ;
 wire \i_game_and_vga.i_game_top.sprite_target.sprite_control.dx[1] ;
 wire \i_game_and_vga.i_game_top.sprite_target.sprite_control.sprite_x[0] ;
 wire \i_game_and_vga.i_game_top.sprite_target.sprite_control.sprite_x[1] ;
 wire \i_game_and_vga.i_game_top.sprite_target.sprite_control.sprite_x[2] ;
 wire \i_game_and_vga.i_game_top.sprite_target.sprite_control.sprite_x[3] ;
 wire \i_game_and_vga.i_game_top.sprite_target.sprite_control.sprite_x[4] ;
 wire \i_game_and_vga.i_game_top.sprite_target.sprite_control.sprite_x[5] ;
 wire \i_game_and_vga.i_game_top.sprite_target.sprite_control.sprite_x[6] ;
 wire \i_game_and_vga.i_game_top.sprite_target.sprite_control.sprite_x[7] ;
 wire \i_game_and_vga.i_game_top.sprite_target.sprite_control.sprite_x[8] ;
 wire \i_game_and_vga.i_game_top.sprite_target.sprite_control.sprite_x[9] ;
 wire \i_game_and_vga.i_game_top.sprite_target.sprite_control.sprite_y[0] ;
 wire \i_game_and_vga.i_game_top.sprite_target.sprite_control.sprite_y[1] ;
 wire \i_game_and_vga.i_game_top.sprite_target.sprite_control.sprite_y[2] ;
 wire \i_game_and_vga.i_game_top.sprite_target.sprite_control.sprite_y[3] ;
 wire \i_game_and_vga.i_game_top.sprite_target.sprite_control.sprite_y[4] ;
 wire \i_game_and_vga.i_game_top.sprite_target.sprite_control.sprite_y[5] ;
 wire \i_game_and_vga.i_game_top.sprite_target.sprite_control.sprite_y[6] ;
 wire \i_game_and_vga.i_game_top.sprite_target.sprite_control.strobe_generator.counter[0] ;
 wire \i_game_and_vga.i_game_top.sprite_target.sprite_control.strobe_generator.counter[10] ;
 wire \i_game_and_vga.i_game_top.sprite_target.sprite_control.strobe_generator.counter[11] ;
 wire \i_game_and_vga.i_game_top.sprite_target.sprite_control.strobe_generator.counter[12] ;
 wire \i_game_and_vga.i_game_top.sprite_target.sprite_control.strobe_generator.counter[13] ;
 wire \i_game_and_vga.i_game_top.sprite_target.sprite_control.strobe_generator.counter[14] ;
 wire \i_game_and_vga.i_game_top.sprite_target.sprite_control.strobe_generator.counter[15] ;
 wire \i_game_and_vga.i_game_top.sprite_target.sprite_control.strobe_generator.counter[16] ;
 wire \i_game_and_vga.i_game_top.sprite_target.sprite_control.strobe_generator.counter[17] ;
 wire \i_game_and_vga.i_game_top.sprite_target.sprite_control.strobe_generator.counter[18] ;
 wire \i_game_and_vga.i_game_top.sprite_target.sprite_control.strobe_generator.counter[1] ;
 wire \i_game_and_vga.i_game_top.sprite_target.sprite_control.strobe_generator.counter[2] ;
 wire \i_game_and_vga.i_game_top.sprite_target.sprite_control.strobe_generator.counter[3] ;
 wire \i_game_and_vga.i_game_top.sprite_target.sprite_control.strobe_generator.counter[4] ;
 wire \i_game_and_vga.i_game_top.sprite_target.sprite_control.strobe_generator.counter[5] ;
 wire \i_game_and_vga.i_game_top.sprite_target.sprite_control.strobe_generator.counter[6] ;
 wire \i_game_and_vga.i_game_top.sprite_target.sprite_control.strobe_generator.counter[7] ;
 wire \i_game_and_vga.i_game_top.sprite_target.sprite_control.strobe_generator.counter[8] ;
 wire \i_game_and_vga.i_game_top.sprite_target.sprite_control.strobe_generator.counter[9] ;
 wire \i_game_and_vga.i_game_top.sprite_target.sprite_control.strobe_generator.strobe ;
 wire \i_game_and_vga.i_game_top.sprite_target.sprite_display.x_sprite_plus_w_1[0] ;
 wire \i_game_and_vga.i_game_top.sprite_target.sprite_display.x_sprite_plus_w_1[1] ;
 wire \i_game_and_vga.i_game_top.sprite_target.sprite_display.x_sprite_plus_w_1[2] ;
 wire \i_game_and_vga.i_game_top.sprite_target.sprite_display.x_sprite_plus_w_1[3] ;
 wire \i_game_and_vga.i_game_top.sprite_target.sprite_display.x_sprite_plus_w_1[4] ;
 wire \i_game_and_vga.i_game_top.sprite_target.sprite_display.x_sprite_plus_w_1[5] ;
 wire \i_game_and_vga.i_game_top.sprite_target.sprite_display.x_sprite_plus_w_1[6] ;
 wire \i_game_and_vga.i_game_top.sprite_target.sprite_display.x_sprite_plus_w_1[7] ;
 wire \i_game_and_vga.i_game_top.sprite_target.sprite_display.x_sprite_plus_w_1[8] ;
 wire \i_game_and_vga.i_game_top.sprite_target.sprite_display.x_sprite_plus_w_1[9] ;
 wire \i_game_and_vga.i_game_top.sprite_target.sprite_display.x_sprite_within_screen ;
 wire \i_game_and_vga.i_game_top.sprite_target.sprite_display.y_sprite_plus_h_1[0] ;
 wire \i_game_and_vga.i_game_top.sprite_target.sprite_display.y_sprite_plus_h_1[1] ;
 wire \i_game_and_vga.i_game_top.sprite_target.sprite_display.y_sprite_plus_h_1[2] ;
 wire \i_game_and_vga.i_game_top.sprite_target.sprite_display.y_sprite_plus_h_1[3] ;
 wire \i_game_and_vga.i_game_top.sprite_target.sprite_display.y_sprite_plus_h_1[4] ;
 wire \i_game_and_vga.i_game_top.sprite_target.sprite_display.y_sprite_plus_h_1[5] ;
 wire \i_game_and_vga.i_game_top.sprite_target.sprite_display.y_sprite_plus_h_1[6] ;
 wire \i_game_and_vga.i_game_top.sprite_target.sprite_display.y_sprite_plus_h_1[7] ;
 wire \i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.dx[0] ;
 wire \i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.dx[1] ;
 wire \i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.dy[0] ;
 wire \i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.dy[1] ;
 wire \i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.sprite_x[0] ;
 wire \i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.sprite_x[1] ;
 wire \i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.sprite_x[2] ;
 wire \i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.sprite_x[3] ;
 wire \i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.sprite_x[4] ;
 wire \i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.sprite_x[5] ;
 wire \i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.sprite_x[6] ;
 wire \i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.sprite_x[7] ;
 wire \i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.sprite_x[8] ;
 wire \i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.sprite_x[9] ;
 wire \i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.sprite_y[0] ;
 wire \i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.sprite_y[1] ;
 wire \i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.sprite_y[2] ;
 wire \i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.sprite_y[3] ;
 wire \i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.sprite_y[4] ;
 wire \i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.sprite_y[5] ;
 wire \i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.sprite_y[6] ;
 wire \i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.sprite_y[7] ;
 wire \i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.sprite_y[8] ;
 wire \i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.strobe_generator.counter[0] ;
 wire \i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.strobe_generator.counter[10] ;
 wire \i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.strobe_generator.counter[11] ;
 wire \i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.strobe_generator.counter[12] ;
 wire \i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.strobe_generator.counter[13] ;
 wire \i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.strobe_generator.counter[14] ;
 wire \i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.strobe_generator.counter[15] ;
 wire \i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.strobe_generator.counter[16] ;
 wire \i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.strobe_generator.counter[17] ;
 wire \i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.strobe_generator.counter[18] ;
 wire \i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.strobe_generator.counter[1] ;
 wire \i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.strobe_generator.counter[2] ;
 wire \i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.strobe_generator.counter[3] ;
 wire \i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.strobe_generator.counter[4] ;
 wire \i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.strobe_generator.counter[5] ;
 wire \i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.strobe_generator.counter[6] ;
 wire \i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.strobe_generator.counter[7] ;
 wire \i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.strobe_generator.counter[8] ;
 wire \i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.strobe_generator.counter[9] ;
 wire \i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.strobe_generator.strobe ;
 wire \i_game_and_vga.i_game_top.sprite_torpedo.sprite_display.x_sprite_plus_w_1[0] ;
 wire \i_game_and_vga.i_game_top.sprite_torpedo.sprite_display.x_sprite_plus_w_1[1] ;
 wire \i_game_and_vga.i_game_top.sprite_torpedo.sprite_display.x_sprite_plus_w_1[2] ;
 wire \i_game_and_vga.i_game_top.sprite_torpedo.sprite_display.x_sprite_plus_w_1[3] ;
 wire \i_game_and_vga.i_game_top.sprite_torpedo.sprite_display.x_sprite_plus_w_1[4] ;
 wire \i_game_and_vga.i_game_top.sprite_torpedo.sprite_display.x_sprite_plus_w_1[5] ;
 wire \i_game_and_vga.i_game_top.sprite_torpedo.sprite_display.x_sprite_plus_w_1[6] ;
 wire \i_game_and_vga.i_game_top.sprite_torpedo.sprite_display.x_sprite_plus_w_1[7] ;
 wire \i_game_and_vga.i_game_top.sprite_torpedo.sprite_display.x_sprite_plus_w_1[8] ;
 wire \i_game_and_vga.i_game_top.sprite_torpedo.sprite_display.x_sprite_plus_w_1[9] ;
 wire \i_game_and_vga.i_game_top.sprite_torpedo.sprite_display.y_sprite_plus_h_1[0] ;
 wire \i_game_and_vga.i_game_top.sprite_torpedo.sprite_display.y_sprite_plus_h_1[1] ;
 wire \i_game_and_vga.i_game_top.sprite_torpedo.sprite_display.y_sprite_plus_h_1[2] ;
 wire \i_game_and_vga.i_game_top.sprite_torpedo.sprite_display.y_sprite_plus_h_1[3] ;
 wire \i_game_and_vga.i_game_top.sprite_torpedo.sprite_display.y_sprite_plus_h_1[4] ;
 wire \i_game_and_vga.i_game_top.sprite_torpedo.sprite_display.y_sprite_plus_h_1[5] ;
 wire \i_game_and_vga.i_game_top.sprite_torpedo.sprite_display.y_sprite_plus_h_1[6] ;
 wire \i_game_and_vga.i_game_top.sprite_torpedo.sprite_display.y_sprite_plus_h_1[7] ;
 wire \i_game_and_vga.i_game_top.sprite_torpedo.sprite_display.y_sprite_plus_h_1[8] ;
 wire \i_game_and_vga.i_game_top.timer.counter[0] ;
 wire \i_game_and_vga.i_game_top.timer.counter[10] ;
 wire \i_game_and_vga.i_game_top.timer.counter[11] ;
 wire \i_game_and_vga.i_game_top.timer.counter[12] ;
 wire \i_game_and_vga.i_game_top.timer.counter[13] ;
 wire \i_game_and_vga.i_game_top.timer.counter[14] ;
 wire \i_game_and_vga.i_game_top.timer.counter[15] ;
 wire \i_game_and_vga.i_game_top.timer.counter[16] ;
 wire \i_game_and_vga.i_game_top.timer.counter[17] ;
 wire \i_game_and_vga.i_game_top.timer.counter[18] ;
 wire \i_game_and_vga.i_game_top.timer.counter[19] ;
 wire \i_game_and_vga.i_game_top.timer.counter[1] ;
 wire \i_game_and_vga.i_game_top.timer.counter[20] ;
 wire \i_game_and_vga.i_game_top.timer.counter[21] ;
 wire \i_game_and_vga.i_game_top.timer.counter[22] ;
 wire \i_game_and_vga.i_game_top.timer.counter[23] ;
 wire \i_game_and_vga.i_game_top.timer.counter[24] ;
 wire \i_game_and_vga.i_game_top.timer.counter[2] ;
 wire \i_game_and_vga.i_game_top.timer.counter[3] ;
 wire \i_game_and_vga.i_game_top.timer.counter[4] ;
 wire \i_game_and_vga.i_game_top.timer.counter[5] ;
 wire \i_game_and_vga.i_game_top.timer.counter[6] ;
 wire \i_game_and_vga.i_game_top.timer.counter[7] ;
 wire \i_game_and_vga.i_game_top.timer.counter[8] ;
 wire \i_game_and_vga.i_game_top.timer.counter[9] ;
 wire \i_game_and_vga.i_vga.clk_en ;
 wire \i_game_and_vga.i_vga.clk_en_cnt[0] ;
 wire \i_game_and_vga.i_vga.clk_en_cnt[1] ;
 wire \i_game_and_vga.i_vga.clk_en_cnt[2] ;
 wire \i_game_and_vga.i_vga.clk_en_cnt[3] ;
 wire \i_game_and_vga.i_vga.vpos[9] ;
 wire \i_game_and_vga.i_vga.vsync ;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net1;
 wire net2;
 wire net3;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;

 sg13g2_inv_1 _1212_ (.Y(_0536_),
    .A(\i_game_and_vga.i_game_top.end_of_game_timer_start ));
 sg13g2_inv_1 _1213_ (.Y(_0097_),
    .A(net61));
 sg13g2_inv_1 _1214_ (.Y(_0096_),
    .A(net57));
 sg13g2_inv_1 _1215_ (.Y(_0095_),
    .A(net58));
 sg13g2_inv_1 _1216_ (.Y(_0094_),
    .A(net67));
 sg13g2_inv_1 _1217_ (.Y(_0093_),
    .A(net63));
 sg13g2_inv_1 _1218_ (.Y(_0092_),
    .A(net73));
 sg13g2_inv_1 _1219_ (.Y(_0091_),
    .A(net182));
 sg13g2_inv_1 _1220_ (.Y(_0090_),
    .A(net55));
 sg13g2_inv_1 _1221_ (.Y(_0088_),
    .A(net60));
 sg13g2_inv_1 _1222_ (.Y(_0537_),
    .A(net365));
 sg13g2_inv_1 _1223_ (.Y(_0538_),
    .A(net339));
 sg13g2_inv_4 _1224_ (.A(net278),
    .Y(_0539_));
 sg13g2_inv_1 _1225_ (.Y(_0540_),
    .A(net304));
 sg13g2_inv_1 _1226_ (.Y(_0541_),
    .A(net91));
 sg13g2_inv_1 _1227_ (.Y(_0542_),
    .A(net113));
 sg13g2_inv_1 _1228_ (.Y(_0543_),
    .A(net412));
 sg13g2_inv_1 _1229_ (.Y(_0544_),
    .A(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.sprite_x[7] ));
 sg13g2_inv_2 _1230_ (.Y(_0545_),
    .A(\i_game_and_vga.i_game_top.sprite_target.pixel_x[7] ));
 sg13g2_inv_1 _1231_ (.Y(_0546_),
    .A(net154));
 sg13g2_inv_2 _1232_ (.Y(_0547_),
    .A(\i_game_and_vga.i_game_top.sprite_target.pixel_x[6] ));
 sg13g2_inv_1 _1233_ (.Y(_0548_),
    .A(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.sprite_x[5] ));
 sg13g2_inv_1 _1234_ (.Y(_0549_),
    .A(\i_game_and_vga.i_game_top.sprite_target.pixel_x[5] ));
 sg13g2_inv_1 _1235_ (.Y(_0550_),
    .A(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.sprite_x[4] ));
 sg13g2_inv_1 _1236_ (.Y(_0551_),
    .A(net285));
 sg13g2_inv_2 _1237_ (.Y(_0552_),
    .A(\i_game_and_vga.i_game_top.sprite_target.pixel_x[3] ));
 sg13g2_inv_2 _1238_ (.Y(_0553_),
    .A(net373));
 sg13g2_inv_1 _1239_ (.Y(_0554_),
    .A(net82));
 sg13g2_inv_1 _1240_ (.Y(_0555_),
    .A(\i_game_and_vga.i_game_top.sprite_target.pixel_y[8] ));
 sg13g2_inv_1 _1241_ (.Y(_0556_),
    .A(net181));
 sg13g2_inv_1 _1242_ (.Y(_0557_),
    .A(net311));
 sg13g2_inv_1 _1243_ (.Y(_0558_),
    .A(net98));
 sg13g2_inv_1 _1244_ (.Y(_0559_),
    .A(\i_game_and_vga.i_game_top.sprite_target.pixel_y[6] ));
 sg13g2_inv_2 _1245_ (.Y(_0560_),
    .A(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.sprite_y[5] ));
 sg13g2_inv_2 _1246_ (.Y(_0561_),
    .A(\i_game_and_vga.i_game_top.sprite_target.pixel_y[5] ));
 sg13g2_inv_2 _1247_ (.Y(_0562_),
    .A(net368));
 sg13g2_inv_1 _1248_ (.Y(_0563_),
    .A(net289));
 sg13g2_inv_1 _1249_ (.Y(_0564_),
    .A(net290));
 sg13g2_inv_2 _1250_ (.Y(_0565_),
    .A(net312));
 sg13g2_inv_2 _1251_ (.Y(_0566_),
    .A(\i_game_and_vga.i_game_top.sprite_target.pixel_y[2] ));
 sg13g2_inv_1 _1252_ (.Y(_0567_),
    .A(net396));
 sg13g2_inv_1 _1253_ (.Y(_0568_),
    .A(net198));
 sg13g2_inv_1 _1254_ (.Y(_0569_),
    .A(\i_game_and_vga.i_game_top.sprite_target.sprite_control.sprite_x[7] ));
 sg13g2_inv_1 _1255_ (.Y(_0570_),
    .A(\i_game_and_vga.i_game_top.sprite_target.sprite_control.sprite_x[6] ));
 sg13g2_inv_1 _1256_ (.Y(_0571_),
    .A(\i_game_and_vga.i_game_top.sprite_target.sprite_control.sprite_x[5] ));
 sg13g2_inv_1 _1257_ (.Y(_0572_),
    .A(net258));
 sg13g2_inv_1 _1258_ (.Y(_0573_),
    .A(net246));
 sg13g2_inv_2 _1259_ (.Y(_0574_),
    .A(net66));
 sg13g2_inv_1 _1260_ (.Y(_0575_),
    .A(net79));
 sg13g2_inv_1 _1261_ (.Y(_0576_),
    .A(\i_game_and_vga.i_game_top.sprite_target.sprite_control.sprite_y[4] ));
 sg13g2_inv_1 _1262_ (.Y(_0577_),
    .A(net68));
 sg13g2_inv_1 _1263_ (.Y(_0578_),
    .A(_0034_));
 sg13g2_inv_1 _1264_ (.Y(_0579_),
    .A(net122));
 sg13g2_inv_1 _1265_ (.Y(_0580_),
    .A(net131));
 sg13g2_inv_1 _1266_ (.Y(_0581_),
    .A(net124));
 sg13g2_inv_1 _1267_ (.Y(_0582_),
    .A(net141));
 sg13g2_inv_1 _1268_ (.Y(_0583_),
    .A(net145));
 sg13g2_inv_1 _1269_ (.Y(_0584_),
    .A(net118));
 sg13g2_inv_1 _1270_ (.Y(_0585_),
    .A(net189));
 sg13g2_inv_1 _1271_ (.Y(_0586_),
    .A(_0036_));
 sg13g2_inv_1 _1272_ (.Y(_0587_),
    .A(\i_game_and_vga.i_game_top.overlap.left_2[8] ));
 sg13g2_inv_1 _1273_ (.Y(_0588_),
    .A(\i_game_and_vga.i_game_top.overlap.right_1[7] ));
 sg13g2_inv_1 _1274_ (.Y(_0589_),
    .A(\i_game_and_vga.i_game_top.overlap.right_1[6] ));
 sg13g2_inv_1 _1275_ (.Y(_0590_),
    .A(\i_game_and_vga.i_game_top.overlap.left_2[6] ));
 sg13g2_inv_1 _1276_ (.Y(_0591_),
    .A(\i_game_and_vga.i_game_top.overlap.left_2[5] ));
 sg13g2_inv_1 _1277_ (.Y(_0592_),
    .A(\i_game_and_vga.i_game_top.overlap.left_2[4] ));
 sg13g2_inv_1 _1278_ (.Y(_0593_),
    .A(\i_game_and_vga.i_game_top.overlap.right_1[4] ));
 sg13g2_inv_1 _1279_ (.Y(_0594_),
    .A(\i_game_and_vga.i_game_top.overlap.right_1[3] ));
 sg13g2_inv_1 _1280_ (.Y(_0595_),
    .A(\i_game_and_vga.i_game_top.overlap.right_1[1] ));
 sg13g2_inv_1 _1281_ (.Y(_0596_),
    .A(\i_game_and_vga.i_game_top.overlap.right_1[0] ));
 sg13g2_inv_1 _1282_ (.Y(_0597_),
    .A(\i_game_and_vga.i_game_top.overlap.left_1[8] ));
 sg13g2_inv_1 _1283_ (.Y(_0598_),
    .A(\i_game_and_vga.i_game_top.overlap.left_1[7] ));
 sg13g2_inv_1 _1284_ (.Y(_0599_),
    .A(\i_game_and_vga.i_game_top.overlap.left_1[5] ));
 sg13g2_inv_1 _1285_ (.Y(_0600_),
    .A(\i_game_and_vga.i_game_top.overlap.right_2[5] ));
 sg13g2_inv_1 _1286_ (.Y(_0601_),
    .A(\i_game_and_vga.i_game_top.overlap.right_2[4] ));
 sg13g2_inv_1 _1287_ (.Y(_0602_),
    .A(\i_game_and_vga.i_game_top.overlap.left_1[3] ));
 sg13g2_inv_1 _1288_ (.Y(_0603_),
    .A(\i_game_and_vga.i_game_top.overlap.right_2[2] ));
 sg13g2_inv_1 _1289_ (.Y(_0604_),
    .A(\i_game_and_vga.i_game_top.overlap.right_2[1] ));
 sg13g2_inv_1 _1290_ (.Y(_0605_),
    .A(\i_game_and_vga.i_game_top.overlap.top_2[6] ));
 sg13g2_inv_1 _1291_ (.Y(_0606_),
    .A(\i_game_and_vga.i_game_top.overlap.bottom_1[5] ));
 sg13g2_inv_1 _1292_ (.Y(_0607_),
    .A(\i_game_and_vga.i_game_top.overlap.top_2[4] ));
 sg13g2_inv_1 _1293_ (.Y(_0608_),
    .A(\i_game_and_vga.i_game_top.overlap.bottom_1[4] ));
 sg13g2_inv_1 _1294_ (.Y(_0609_),
    .A(\i_game_and_vga.i_game_top.overlap.top_2[3] ));
 sg13g2_inv_1 _1295_ (.Y(_0610_),
    .A(\i_game_and_vga.i_game_top.overlap.top_2[2] ));
 sg13g2_inv_1 _1296_ (.Y(_0611_),
    .A(\i_game_and_vga.i_game_top.overlap.bottom_2[6] ));
 sg13g2_inv_1 _1297_ (.Y(_0612_),
    .A(\i_game_and_vga.i_game_top.overlap.bottom_2[5] ));
 sg13g2_inv_1 _1298_ (.Y(_0613_),
    .A(\i_game_and_vga.i_game_top.overlap.bottom_2[4] ));
 sg13g2_inv_1 _1299_ (.Y(_0614_),
    .A(\i_game_and_vga.i_game_top.overlap.top_1[4] ));
 sg13g2_inv_1 _1300_ (.Y(_0615_),
    .A(\i_game_and_vga.i_game_top.overlap.bottom_2[3] ));
 sg13g2_inv_1 _1301_ (.Y(_0616_),
    .A(\i_game_and_vga.i_game_top.overlap.bottom_2[2] ));
 sg13g2_inv_1 _1302_ (.Y(_0617_),
    .A(net90));
 sg13g2_inv_1 _1303_ (.Y(_0618_),
    .A(net296));
 sg13g2_inv_1 _1304_ (.Y(_0619_),
    .A(net86));
 sg13g2_inv_1 _1305_ (.Y(_0620_),
    .A(_0016_));
 sg13g2_inv_1 _1306_ (.Y(_0621_),
    .A(net217));
 sg13g2_inv_1 _1307_ (.Y(_0622_),
    .A(_0017_));
 sg13g2_inv_1 _1308_ (.Y(_0623_),
    .A(net308));
 sg13g2_inv_1 _1309_ (.Y(_0624_),
    .A(net236));
 sg13g2_nand3_1 _1310_ (.B(net226),
    .C(net116),
    .A(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.strobe_generator.counter[0] ),
    .Y(_0625_));
 sg13g2_and4_2 _1311_ (.A(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.strobe_generator.counter[0] ),
    .B(net120),
    .C(net226),
    .D(net116),
    .X(_0626_));
 sg13g2_nand3_1 _1312_ (.B(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.strobe_generator.counter[4] ),
    .C(_0626_),
    .A(net210),
    .Y(_0627_));
 sg13g2_a21o_1 _1313_ (.A2(_0626_),
    .A1(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.strobe_generator.counter[4] ),
    .B1(net210),
    .X(_0628_));
 sg13g2_nand2_1 _1314_ (.Y(_0104_),
    .A(net211),
    .B(_0628_));
 sg13g2_a21o_1 _1315_ (.A2(net116),
    .A1(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.strobe_generator.counter[0] ),
    .B1(net226),
    .X(_0629_));
 sg13g2_nand2_1 _1316_ (.Y(_0103_),
    .A(net227),
    .B(_0629_));
 sg13g2_xnor2_1 _1317_ (.Y(_0102_),
    .A(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.strobe_generator.counter[0] ),
    .B(net116));
 sg13g2_nand3_1 _1318_ (.B(\i_game_and_vga.i_game_top.sprite_target.sprite_control.strobe_generator.counter[1] ),
    .C(\i_game_and_vga.i_game_top.sprite_target.sprite_control.strobe_generator.counter[0] ),
    .A(net138),
    .Y(_0630_));
 sg13g2_and4_2 _1319_ (.A(net126),
    .B(net138),
    .C(net147),
    .D(\i_game_and_vga.i_game_top.sprite_target.sprite_control.strobe_generator.counter[0] ),
    .X(_0631_));
 sg13g2_nand3_1 _1320_ (.B(\i_game_and_vga.i_game_top.sprite_target.sprite_control.strobe_generator.counter[4] ),
    .C(_0631_),
    .A(net172),
    .Y(_0632_));
 sg13g2_a21o_1 _1321_ (.A2(_0631_),
    .A1(\i_game_and_vga.i_game_top.sprite_target.sprite_control.strobe_generator.counter[4] ),
    .B1(net172),
    .X(_0633_));
 sg13g2_nand2_1 _1322_ (.Y(_0101_),
    .A(net173),
    .B(_0633_));
 sg13g2_a21o_1 _1323_ (.A2(\i_game_and_vga.i_game_top.sprite_target.sprite_control.strobe_generator.counter[0] ),
    .A1(\i_game_and_vga.i_game_top.sprite_target.sprite_control.strobe_generator.counter[1] ),
    .B1(net138),
    .X(_0634_));
 sg13g2_nand2_1 _1324_ (.Y(_0100_),
    .A(net139),
    .B(_0634_));
 sg13g2_xnor2_1 _1325_ (.Y(_0099_),
    .A(net147),
    .B(\i_game_and_vga.i_game_top.sprite_target.sprite_control.strobe_generator.counter[0] ));
 sg13g2_xnor2_1 _1326_ (.Y(_0098_),
    .A(\i_game_and_vga.i_game_top.random[15] ),
    .B(net64));
 sg13g2_xnor2_1 _1327_ (.Y(_0089_),
    .A(\i_game_and_vga.i_game_top.random[15] ),
    .B(net71));
 sg13g2_xnor2_1 _1328_ (.Y(_0087_),
    .A(\i_game_and_vga.i_game_top.random[15] ),
    .B(net223));
 sg13g2_nor2b_1 _1329_ (.A(net213),
    .B_N(\i_game_and_vga.i_game_top.master_fsm.state[1] ),
    .Y(\i_game_and_vga.i_game_top.master_fsm.d_sprite_torpedo_enable_update ));
 sg13g2_or3_2 _1330_ (.A(\i_game_and_vga.i_game_top.sprite_target.sprite_control.sprite_y[2] ),
    .B(net310),
    .C(net363),
    .X(_0635_));
 sg13g2_nand3_1 _1331_ (.B(net106),
    .C(_0635_),
    .A(net78),
    .Y(_0636_));
 sg13g2_or2_1 _1332_ (.X(_0637_),
    .B(_0636_),
    .A(_0575_));
 sg13g2_nor2_2 _1333_ (.A(_0574_),
    .B(_0637_),
    .Y(\i_game_and_vga.i_game_top.sprite_target.sprite_display.y_sprite_plus_h_1[7] ));
 sg13g2_nand4_1 _1334_ (.B(net172),
    .C(\i_game_and_vga.i_game_top.sprite_target.sprite_control.strobe_generator.counter[4] ),
    .A(net128),
    .Y(_0638_),
    .D(_0631_));
 sg13g2_nor2_2 _1335_ (.A(_0580_),
    .B(_0638_),
    .Y(_0639_));
 sg13g2_nand3_1 _1336_ (.B(net206),
    .C(_0639_),
    .A(net392),
    .Y(_0640_));
 sg13g2_and4_1 _1337_ (.A(net114),
    .B(\i_game_and_vga.i_game_top.sprite_target.sprite_control.strobe_generator.counter[9] ),
    .C(\i_game_and_vga.i_game_top.sprite_target.sprite_control.strobe_generator.counter[8] ),
    .D(_0639_),
    .X(_0641_));
 sg13g2_nand3_1 _1338_ (.B(net170),
    .C(_0641_),
    .A(net380),
    .Y(_0642_));
 sg13g2_nor2_1 _1339_ (.A(_0579_),
    .B(_0642_),
    .Y(_0643_));
 sg13g2_nand3_1 _1340_ (.B(net158),
    .C(_0643_),
    .A(net188),
    .Y(_0644_));
 sg13g2_nor2_1 _1341_ (.A(_0581_),
    .B(_0644_),
    .Y(_0645_));
 sg13g2_and3_1 _1342_ (.X(_0004_),
    .A(net111),
    .B(net103),
    .C(_0645_));
 sg13g2_nand4_1 _1343_ (.B(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.strobe_generator.counter[5] ),
    .C(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.strobe_generator.counter[4] ),
    .A(net133),
    .Y(_0646_),
    .D(_0626_));
 sg13g2_nor2_2 _1344_ (.A(_0583_),
    .B(_0646_),
    .Y(_0647_));
 sg13g2_nand3_1 _1345_ (.B(net196),
    .C(_0647_),
    .A(net388),
    .Y(_0648_));
 sg13g2_and4_1 _1346_ (.A(net162),
    .B(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.strobe_generator.counter[9] ),
    .C(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.strobe_generator.counter[8] ),
    .D(_0647_),
    .X(_0649_));
 sg13g2_nand3_1 _1347_ (.B(net183),
    .C(_0649_),
    .A(net370),
    .Y(_0650_));
 sg13g2_nor2_1 _1348_ (.A(_0582_),
    .B(_0650_),
    .Y(_0651_));
 sg13g2_nand3_1 _1349_ (.B(net415),
    .C(_0651_),
    .A(net143),
    .Y(_0652_));
 sg13g2_nor2_1 _1350_ (.A(_0584_),
    .B(_0652_),
    .Y(_0653_));
 sg13g2_and3_1 _1351_ (.X(_0006_),
    .A(net109),
    .B(net99),
    .C(_0653_));
 sg13g2_nor4_1 _1352_ (.A(\i_game_and_vga.i_vga.clk_en_cnt[1] ),
    .B(\i_game_and_vga.i_vga.clk_en_cnt[0] ),
    .C(\i_game_and_vga.i_vga.clk_en_cnt[3] ),
    .D(net92),
    .Y(_0010_));
 sg13g2_nor2_1 _1353_ (.A(_0597_),
    .B(\i_game_and_vga.i_game_top.overlap.right_2[8] ),
    .Y(_0654_));
 sg13g2_nor2_1 _1354_ (.A(_0602_),
    .B(\i_game_and_vga.i_game_top.overlap.right_2[3] ),
    .Y(_0655_));
 sg13g2_nor2b_1 _1355_ (.A(\i_game_and_vga.i_game_top.overlap.right_2[0] ),
    .B_N(\i_game_and_vga.i_game_top.overlap.left_1[0] ),
    .Y(_0656_));
 sg13g2_o21ai_1 _1356_ (.B1(_0656_),
    .Y(_0657_),
    .A1(\i_game_and_vga.i_game_top.overlap.left_1[1] ),
    .A2(_0604_));
 sg13g2_a22oi_1 _1357_ (.Y(_0658_),
    .B1(\i_game_and_vga.i_game_top.overlap.left_1[1] ),
    .B2(_0604_),
    .A2(_0603_),
    .A1(\i_game_and_vga.i_game_top.overlap.left_1[2] ));
 sg13g2_nor2_1 _1358_ (.A(\i_game_and_vga.i_game_top.overlap.left_1[2] ),
    .B(_0603_),
    .Y(_0659_));
 sg13g2_a221oi_1 _1359_ (.B2(_0658_),
    .C1(_0659_),
    .B1(_0657_),
    .A1(_0602_),
    .Y(_0660_),
    .A2(\i_game_and_vga.i_game_top.overlap.right_2[3] ));
 sg13g2_nand2b_1 _1360_ (.Y(_0661_),
    .B(\i_game_and_vga.i_game_top.overlap.right_2[4] ),
    .A_N(\i_game_and_vga.i_game_top.overlap.left_1[4] ));
 sg13g2_o21ai_1 _1361_ (.B1(_0661_),
    .Y(_0662_),
    .A1(_0655_),
    .A2(_0660_));
 sg13g2_a22oi_1 _1362_ (.Y(_0663_),
    .B1(_0601_),
    .B2(\i_game_and_vga.i_game_top.overlap.left_1[4] ),
    .A2(_0600_),
    .A1(\i_game_and_vga.i_game_top.overlap.left_1[5] ));
 sg13g2_nand2b_1 _1363_ (.Y(_0664_),
    .B(\i_game_and_vga.i_game_top.overlap.right_2[6] ),
    .A_N(\i_game_and_vga.i_game_top.overlap.left_1[6] ));
 sg13g2_a22oi_1 _1364_ (.Y(_0665_),
    .B1(_0662_),
    .B2(_0663_),
    .A2(\i_game_and_vga.i_game_top.overlap.right_2[5] ),
    .A1(_0599_));
 sg13g2_nand2b_1 _1365_ (.Y(_0666_),
    .B(\i_game_and_vga.i_game_top.overlap.left_1[6] ),
    .A_N(\i_game_and_vga.i_game_top.overlap.right_2[6] ));
 sg13g2_o21ai_1 _1366_ (.B1(_0666_),
    .Y(_0667_),
    .A1(_0598_),
    .A2(\i_game_and_vga.i_game_top.overlap.right_2[7] ));
 sg13g2_a21oi_1 _1367_ (.A1(_0664_),
    .A2(_0665_),
    .Y(_0668_),
    .B1(_0667_));
 sg13g2_a221oi_1 _1368_ (.B2(\i_game_and_vga.i_game_top.overlap.right_2[7] ),
    .C1(_0668_),
    .B1(_0598_),
    .A1(_0597_),
    .Y(_0669_),
    .A2(\i_game_and_vga.i_game_top.overlap.right_2[8] ));
 sg13g2_nand2b_1 _1369_ (.Y(_0670_),
    .B(\i_game_and_vga.i_game_top.overlap.right_2[9] ),
    .A_N(\i_game_and_vga.i_game_top.overlap.left_1[9] ));
 sg13g2_o21ai_1 _1370_ (.B1(_0670_),
    .Y(_0671_),
    .A1(_0654_),
    .A2(_0669_));
 sg13g2_nand2b_1 _1371_ (.Y(_0672_),
    .B(\i_game_and_vga.i_game_top.overlap.right_1[9] ),
    .A_N(\i_game_and_vga.i_game_top.overlap.left_2[9] ));
 sg13g2_a22oi_1 _1372_ (.Y(_0673_),
    .B1(_0596_),
    .B2(\i_game_and_vga.i_game_top.overlap.left_2[0] ),
    .A2(\i_game_and_vga.i_game_top.overlap.left_2[1] ),
    .A1(_0595_));
 sg13g2_nand2b_1 _1373_ (.Y(_0674_),
    .B(\i_game_and_vga.i_game_top.overlap.right_1[2] ),
    .A_N(\i_game_and_vga.i_game_top.overlap.left_2[2] ));
 sg13g2_o21ai_1 _1374_ (.B1(_0674_),
    .Y(_0675_),
    .A1(_0595_),
    .A2(\i_game_and_vga.i_game_top.overlap.left_2[1] ));
 sg13g2_nand2b_1 _1375_ (.Y(_0676_),
    .B(\i_game_and_vga.i_game_top.overlap.left_2[2] ),
    .A_N(\i_game_and_vga.i_game_top.overlap.right_1[2] ));
 sg13g2_nor2_1 _1376_ (.A(\i_game_and_vga.i_game_top.overlap.right_1[5] ),
    .B(_0591_),
    .Y(_0677_));
 sg13g2_o21ai_1 _1377_ (.B1(_0676_),
    .Y(_0678_),
    .A1(_0673_),
    .A2(_0675_));
 sg13g2_o21ai_1 _1378_ (.B1(_0678_),
    .Y(_0679_),
    .A1(_0594_),
    .A2(\i_game_and_vga.i_game_top.overlap.left_2[3] ));
 sg13g2_a22oi_1 _1379_ (.Y(_0680_),
    .B1(_0594_),
    .B2(\i_game_and_vga.i_game_top.overlap.left_2[3] ),
    .A2(_0593_),
    .A1(\i_game_and_vga.i_game_top.overlap.left_2[4] ));
 sg13g2_a22oi_1 _1380_ (.Y(_0681_),
    .B1(_0679_),
    .B2(_0680_),
    .A2(\i_game_and_vga.i_game_top.overlap.right_1[4] ),
    .A1(_0592_));
 sg13g2_a22oi_1 _1381_ (.Y(_0682_),
    .B1(\i_game_and_vga.i_game_top.overlap.right_1[5] ),
    .B2(_0591_),
    .A2(_0590_),
    .A1(\i_game_and_vga.i_game_top.overlap.right_1[6] ));
 sg13g2_o21ai_1 _1382_ (.B1(_0682_),
    .Y(_0683_),
    .A1(_0677_),
    .A2(_0681_));
 sg13g2_a22oi_1 _1383_ (.Y(_0684_),
    .B1(_0589_),
    .B2(\i_game_and_vga.i_game_top.overlap.left_2[6] ),
    .A2(\i_game_and_vga.i_game_top.overlap.left_2[7] ),
    .A1(_0588_));
 sg13g2_nor2_1 _1384_ (.A(_0588_),
    .B(\i_game_and_vga.i_game_top.overlap.left_2[7] ),
    .Y(_0685_));
 sg13g2_a221oi_1 _1385_ (.B2(_0684_),
    .C1(_0685_),
    .B1(_0683_),
    .A1(\i_game_and_vga.i_game_top.overlap.right_1[8] ),
    .Y(_0686_),
    .A2(_0587_));
 sg13g2_nand2b_1 _1386_ (.Y(_0687_),
    .B(\i_game_and_vga.i_game_top.overlap.top_1[1] ),
    .A_N(\i_game_and_vga.i_game_top.overlap.bottom_2[1] ));
 sg13g2_nand2b_1 _1387_ (.Y(_0688_),
    .B(\i_game_and_vga.i_game_top.overlap.top_1[0] ),
    .A_N(\i_game_and_vga.i_game_top.overlap.bottom_2[0] ));
 sg13g2_nor2b_1 _1388_ (.A(\i_game_and_vga.i_game_top.overlap.top_1[1] ),
    .B_N(\i_game_and_vga.i_game_top.overlap.bottom_2[1] ),
    .Y(_0689_));
 sg13g2_a21oi_1 _1389_ (.A1(_0687_),
    .A2(_0688_),
    .Y(_0690_),
    .B1(_0689_));
 sg13g2_o21ai_1 _1390_ (.B1(_0690_),
    .Y(_0691_),
    .A1(\i_game_and_vga.i_game_top.overlap.top_1[2] ),
    .A2(_0616_));
 sg13g2_a22oi_1 _1391_ (.Y(_0692_),
    .B1(\i_game_and_vga.i_game_top.overlap.top_1[2] ),
    .B2(_0616_),
    .A2(_0615_),
    .A1(\i_game_and_vga.i_game_top.overlap.top_1[3] ));
 sg13g2_nand2b_1 _1392_ (.Y(_0693_),
    .B(\i_game_and_vga.i_game_top.overlap.bottom_2[3] ),
    .A_N(\i_game_and_vga.i_game_top.overlap.top_1[3] ));
 sg13g2_a22oi_1 _1393_ (.Y(_0694_),
    .B1(_0691_),
    .B2(_0692_),
    .A2(_0614_),
    .A1(\i_game_and_vga.i_game_top.overlap.bottom_2[4] ));
 sg13g2_a22oi_1 _1394_ (.Y(_0695_),
    .B1(_0693_),
    .B2(_0694_),
    .A2(\i_game_and_vga.i_game_top.overlap.top_1[4] ),
    .A1(_0613_));
 sg13g2_nor2_1 _1395_ (.A(\i_game_and_vga.i_game_top.overlap.top_1[5] ),
    .B(_0612_),
    .Y(_0696_));
 sg13g2_a22oi_1 _1396_ (.Y(_0697_),
    .B1(\i_game_and_vga.i_game_top.overlap.top_1[5] ),
    .B2(_0612_),
    .A2(\i_game_and_vga.i_game_top.overlap.top_1[6] ),
    .A1(_0611_));
 sg13g2_o21ai_1 _1397_ (.B1(_0697_),
    .Y(_0698_),
    .A1(_0695_),
    .A2(_0696_));
 sg13g2_o21ai_1 _1398_ (.B1(_0698_),
    .Y(_0699_),
    .A1(_0611_),
    .A2(\i_game_and_vga.i_game_top.overlap.top_1[6] ));
 sg13g2_nor3_1 _1399_ (.A(\i_game_and_vga.i_game_top.overlap.bottom_2[7] ),
    .B(\i_game_and_vga.i_game_top.overlap.bottom_2[8] ),
    .C(_0699_),
    .Y(_0700_));
 sg13g2_nand2b_1 _1400_ (.Y(_0701_),
    .B(\i_game_and_vga.i_game_top.overlap.bottom_1[7] ),
    .A_N(\i_game_and_vga.i_game_top.overlap.top_2[7] ));
 sg13g2_nor2_1 _1401_ (.A(\i_game_and_vga.i_game_top.overlap.bottom_1[6] ),
    .B(_0605_),
    .Y(_0702_));
 sg13g2_nand2b_1 _1402_ (.Y(_0703_),
    .B(\i_game_and_vga.i_game_top.overlap.top_2[1] ),
    .A_N(\i_game_and_vga.i_game_top.overlap.bottom_1[1] ));
 sg13g2_nand2b_1 _1403_ (.Y(_0704_),
    .B(\i_game_and_vga.i_game_top.overlap.bottom_1[1] ),
    .A_N(\i_game_and_vga.i_game_top.overlap.top_2[1] ));
 sg13g2_nand3b_1 _1404_ (.B(_0704_),
    .C(\i_game_and_vga.i_game_top.overlap.top_2[0] ),
    .Y(_0705_),
    .A_N(\i_game_and_vga.i_game_top.overlap.bottom_1[0] ));
 sg13g2_a22oi_1 _1405_ (.Y(_0706_),
    .B1(_0703_),
    .B2(_0705_),
    .A2(_0610_),
    .A1(\i_game_and_vga.i_game_top.overlap.bottom_1[2] ));
 sg13g2_nand2b_1 _1406_ (.Y(_0707_),
    .B(\i_game_and_vga.i_game_top.overlap.top_2[3] ),
    .A_N(\i_game_and_vga.i_game_top.overlap.bottom_1[3] ));
 sg13g2_o21ai_1 _1407_ (.B1(_0707_),
    .Y(_0708_),
    .A1(\i_game_and_vga.i_game_top.overlap.bottom_1[2] ),
    .A2(_0610_));
 sg13g2_a22oi_1 _1408_ (.Y(_0709_),
    .B1(\i_game_and_vga.i_game_top.overlap.bottom_1[3] ),
    .B2(_0609_),
    .A2(\i_game_and_vga.i_game_top.overlap.bottom_1[4] ),
    .A1(_0607_));
 sg13g2_o21ai_1 _1409_ (.B1(_0709_),
    .Y(_0710_),
    .A1(_0706_),
    .A2(_0708_));
 sg13g2_a22oi_1 _1410_ (.Y(_0711_),
    .B1(\i_game_and_vga.i_game_top.overlap.top_2[4] ),
    .B2(_0608_),
    .A2(\i_game_and_vga.i_game_top.overlap.top_2[5] ),
    .A1(_0606_));
 sg13g2_nor2_1 _1411_ (.A(_0606_),
    .B(\i_game_and_vga.i_game_top.overlap.top_2[5] ),
    .Y(_0712_));
 sg13g2_a221oi_1 _1412_ (.B2(_0711_),
    .C1(_0712_),
    .B1(_0710_),
    .A1(\i_game_and_vga.i_game_top.overlap.bottom_1[6] ),
    .Y(_0713_),
    .A2(_0605_));
 sg13g2_o21ai_1 _1413_ (.B1(_0701_),
    .Y(_0714_),
    .A1(_0702_),
    .A2(_0713_));
 sg13g2_nor2b_1 _1414_ (.A(\i_game_and_vga.i_game_top.overlap.bottom_1[7] ),
    .B_N(\i_game_and_vga.i_game_top.overlap.top_2[7] ),
    .Y(_0715_));
 sg13g2_nor2b_1 _1415_ (.A(\i_game_and_vga.i_game_top.overlap.right_2[9] ),
    .B_N(\i_game_and_vga.i_game_top.overlap.left_1[9] ),
    .Y(_0716_));
 sg13g2_nand2b_1 _1416_ (.Y(_0717_),
    .B(\i_game_and_vga.i_game_top.overlap.left_2[9] ),
    .A_N(\i_game_and_vga.i_game_top.overlap.right_1[9] ));
 sg13g2_o21ai_1 _1417_ (.B1(_0717_),
    .Y(_0718_),
    .A1(\i_game_and_vga.i_game_top.overlap.right_1[8] ),
    .A2(_0587_));
 sg13g2_o21ai_1 _1418_ (.B1(_0672_),
    .Y(_0719_),
    .A1(_0686_),
    .A2(_0718_));
 sg13g2_nor4_1 _1419_ (.A(net231),
    .B(_0700_),
    .C(_0715_),
    .D(_0716_),
    .Y(_0720_));
 sg13g2_and4_1 _1420_ (.A(_0671_),
    .B(_0714_),
    .C(_0719_),
    .D(net232),
    .X(_0003_));
 sg13g2_o21ai_1 _1421_ (.B1(net298),
    .Y(\i_game_and_vga.i_game_top.sprite_target.sprite_display.x_sprite_within_screen ),
    .A1(net208),
    .A2(net192));
 sg13g2_nand2_1 _1422_ (.Y(_0721_),
    .A(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.sprite_y[7] ),
    .B(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.sprite_y[6] ));
 sg13g2_nor2_1 _1423_ (.A(net294),
    .B(net292),
    .Y(_0722_));
 sg13g2_nor3_2 _1424_ (.A(net294),
    .B(net291),
    .C(net293),
    .Y(_0723_));
 sg13g2_or3_1 _1425_ (.A(net294),
    .B(net291),
    .C(net292),
    .X(_0724_));
 sg13g2_nand3_1 _1426_ (.B(net290),
    .C(_0724_),
    .A(net289),
    .Y(_0725_));
 sg13g2_nand4_1 _1427_ (.B(net289),
    .C(net290),
    .A(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.sprite_y[5] ),
    .Y(_0726_),
    .D(_0724_));
 sg13g2_nor3_2 _1428_ (.A(net252),
    .B(_0721_),
    .C(_0726_),
    .Y(_0727_));
 sg13g2_inv_1 _1429_ (.Y(_0728_),
    .A(_0727_));
 sg13g2_a21oi_1 _1430_ (.A1(_0542_),
    .A2(_0544_),
    .Y(_0729_),
    .B1(_0541_));
 sg13g2_nor3_1 _1431_ (.A(_0554_),
    .B(_0560_),
    .C(_0721_),
    .Y(_0730_));
 sg13g2_nor3_1 _1432_ (.A(_0727_),
    .B(_0729_),
    .C(_0730_),
    .Y(_0008_));
 sg13g2_nor2_1 _1433_ (.A(net186),
    .B(net93),
    .Y(_0011_));
 sg13g2_xor2_1 _1434_ (.B(net186),
    .A(net225),
    .X(_0012_));
 sg13g2_nand3_1 _1435_ (.B(net186),
    .C(net92),
    .A(net225),
    .Y(_0731_));
 sg13g2_a21o_1 _1436_ (.A2(net186),
    .A1(net225),
    .B1(net92),
    .X(_0732_));
 sg13g2_and2_1 _1437_ (.A(_0731_),
    .B(_0732_),
    .X(_0013_));
 sg13g2_xnor2_1 _1438_ (.Y(_0014_),
    .A(net155),
    .B(_0731_));
 sg13g2_nor2b_1 _1439_ (.A(\i_game_and_vga.i_game_top.mixer.sprite_torpedo_rgb_en ),
    .B_N(\i_game_and_vga.i_game_top.mixer.sprite_target_rgb_en ),
    .Y(_0733_));
 sg13g2_a21oi_1 _1440_ (.A1(\i_game_and_vga.i_game_top.mixer.sprite_target_rgb[0] ),
    .A2(_0733_),
    .Y(_0734_),
    .B1(\i_game_and_vga.i_game_top.end_of_game_timer_running ));
 sg13g2_o21ai_1 _1441_ (.B1(net86),
    .Y(_0735_),
    .A1(_0537_),
    .A2(\i_game_and_vga.i_game_top.mixer.random ));
 sg13g2_nor2_1 _1442_ (.A(_0734_),
    .B(net87),
    .Y(_0000_));
 sg13g2_a221oi_1 _1443_ (.B2(net200),
    .C1(\i_game_and_vga.i_game_top.end_of_game_timer_running ),
    .B1(_0733_),
    .A1(\i_game_and_vga.i_game_top.mixer.sprite_torpedo_rgb_en ),
    .Y(_0736_),
    .A2(_0620_));
 sg13g2_nor2_1 _1444_ (.A(_0537_),
    .B(_0621_),
    .Y(_0737_));
 sg13g2_nor3_1 _1445_ (.A(_0619_),
    .B(_0736_),
    .C(net218),
    .Y(_0001_));
 sg13g2_a221oi_1 _1446_ (.B2(net178),
    .C1(_0568_),
    .B1(_0733_),
    .A1(\i_game_and_vga.i_game_top.mixer.sprite_torpedo_rgb_en ),
    .Y(_0738_),
    .A2(\i_game_and_vga.i_game_top.mixer.sprite_torpedo_rgb[2] ));
 sg13g2_nor2_1 _1447_ (.A(_0619_),
    .B(net199),
    .Y(_0002_));
 sg13g2_xor2_1 _1448_ (.B(net239),
    .A(net213),
    .X(\i_game_and_vga.i_game_top.master_fsm.d_sprite_target_enable_update ));
 sg13g2_nand3b_1 _1449_ (.B(\i_game_and_vga.i_game_top.master_fsm.sprite_target_within_screen ),
    .C(\i_game_and_vga.i_game_top.master_fsm.sprite_torpedo_within_screen ),
    .Y(_0739_),
    .A_N(\i_game_and_vga.i_game_top.collision ));
 sg13g2_and2_1 _1450_ (.A(\i_game_and_vga.i_game_top.master_fsm.d_sprite_target_enable_update ),
    .B(_0739_),
    .X(\i_game_and_vga.i_game_top.master_fsm.d_end_of_game_timer_start ));
 sg13g2_nor2_1 _1451_ (.A(net213),
    .B(net239),
    .Y(\i_game_and_vga.i_game_top.master_fsm.d_sprite_target_write_dxy ));
 sg13g2_or3_2 _1452_ (.A(net303),
    .B(\i_game_and_vga.i_game_top.sprite_target.sprite_control.sprite_x[2] ),
    .C(net302),
    .X(_0740_));
 sg13g2_nand3_1 _1453_ (.B(net301),
    .C(_0740_),
    .A(net300),
    .Y(_0741_));
 sg13g2_nand4_1 _1454_ (.B(net300),
    .C(net301),
    .A(\i_game_and_vga.i_game_top.sprite_target.sprite_control.sprite_x[5] ),
    .Y(_0742_),
    .D(_0740_));
 sg13g2_nor3_2 _1455_ (.A(_0569_),
    .B(_0570_),
    .C(_0742_),
    .Y(_0743_));
 sg13g2_and3_1 _1456_ (.X(_0744_),
    .A(net216),
    .B(net208),
    .C(_0743_));
 sg13g2_nand3_1 _1457_ (.B(\i_game_and_vga.i_game_top.sprite_target.sprite_control.sprite_x[8] ),
    .C(_0743_),
    .A(net298),
    .Y(_0745_));
 sg13g2_a21oi_1 _1458_ (.A1(net299),
    .A2(_0743_),
    .Y(_0746_),
    .B1(net298));
 sg13g2_nor2_1 _1459_ (.A(_0744_),
    .B(_0746_),
    .Y(\i_game_and_vga.i_game_top.sprite_target.sprite_display.x_sprite_plus_w_1[9] ));
 sg13g2_nand2b_1 _1460_ (.Y(_0747_),
    .B(net304),
    .A_N(\i_game_and_vga.i_game_top.sprite_target.sprite_display.x_sprite_plus_w_1[9] ));
 sg13g2_xor2_1 _1461_ (.B(_0743_),
    .A(net299),
    .X(\i_game_and_vga.i_game_top.sprite_target.sprite_display.x_sprite_plus_w_1[8] ));
 sg13g2_nand2_1 _1462_ (.Y(_0748_),
    .A(_0543_),
    .B(\i_game_and_vga.i_game_top.sprite_target.sprite_display.x_sprite_plus_w_1[8] ));
 sg13g2_o21ai_1 _1463_ (.B1(net89),
    .Y(_0749_),
    .A1(net303),
    .A2(net302));
 sg13g2_nand2_2 _1464_ (.Y(\i_game_and_vga.i_game_top.sprite_target.sprite_display.x_sprite_plus_w_1[2] ),
    .A(_0740_),
    .B(_0749_));
 sg13g2_nand2b_1 _1465_ (.Y(_0750_),
    .B(\i_game_and_vga.i_game_top.sprite_target.pixel_x[1] ),
    .A_N(\i_game_and_vga.i_game_top.sprite_target.sprite_control.sprite_x[1] ));
 sg13g2_nor2b_1 _1466_ (.A(\i_game_and_vga.i_game_top.sprite_target.pixel_x[1] ),
    .B_N(\i_game_and_vga.i_game_top.sprite_target.sprite_control.sprite_x[1] ),
    .Y(_0751_));
 sg13g2_nor2b_1 _1467_ (.A(\i_game_and_vga.i_game_top.sprite_target.pixel_x[0] ),
    .B_N(net303),
    .Y(_0752_));
 sg13g2_a21oi_2 _1468_ (.B1(_0751_),
    .Y(_0753_),
    .A2(_0752_),
    .A1(_0750_));
 sg13g2_o21ai_1 _1469_ (.B1(_0753_),
    .Y(_0754_),
    .A1(net303),
    .A2(net302));
 sg13g2_xor2_1 _1470_ (.B(\i_game_and_vga.i_game_top.sprite_target.sprite_display.x_sprite_plus_w_1[2] ),
    .A(_0024_),
    .X(_0755_));
 sg13g2_xnor2_1 _1471_ (.Y(\i_game_and_vga.i_game_top.sprite_target.sprite_display.x_sprite_plus_w_1[3] ),
    .A(_0573_),
    .B(_0740_));
 sg13g2_and2_1 _1472_ (.A(_0552_),
    .B(\i_game_and_vga.i_game_top.sprite_target.sprite_display.x_sprite_plus_w_1[3] ),
    .X(_0756_));
 sg13g2_a221oi_1 _1473_ (.B2(_0755_),
    .C1(_0756_),
    .B1(_0754_),
    .A1(_0553_),
    .Y(_0757_),
    .A2(\i_game_and_vga.i_game_top.sprite_target.sprite_display.x_sprite_plus_w_1[2] ));
 sg13g2_a21o_1 _1474_ (.A2(_0740_),
    .A1(net301),
    .B1(net300),
    .X(_0758_));
 sg13g2_and2_1 _1475_ (.A(_0741_),
    .B(_0758_),
    .X(\i_game_and_vga.i_game_top.sprite_target.sprite_display.x_sprite_plus_w_1[4] ));
 sg13g2_nand2b_1 _1476_ (.Y(_0759_),
    .B(\i_game_and_vga.i_game_top.sprite_target.pixel_x[3] ),
    .A_N(\i_game_and_vga.i_game_top.sprite_target.sprite_display.x_sprite_plus_w_1[3] ));
 sg13g2_o21ai_1 _1477_ (.B1(_0759_),
    .Y(_0760_),
    .A1(_0023_),
    .A2(\i_game_and_vga.i_game_top.sprite_target.sprite_display.x_sprite_plus_w_1[4] ));
 sg13g2_xnor2_1 _1478_ (.Y(\i_game_and_vga.i_game_top.sprite_target.sprite_display.x_sprite_plus_w_1[5] ),
    .A(net416),
    .B(_0741_));
 sg13g2_a22oi_1 _1479_ (.Y(_0761_),
    .B1(\i_game_and_vga.i_game_top.sprite_target.sprite_display.x_sprite_plus_w_1[5] ),
    .B2(_0549_),
    .A2(\i_game_and_vga.i_game_top.sprite_target.sprite_display.x_sprite_plus_w_1[4] ),
    .A1(_0023_));
 sg13g2_o21ai_1 _1480_ (.B1(_0761_),
    .Y(_0762_),
    .A1(_0757_),
    .A2(_0760_));
 sg13g2_nor2_1 _1481_ (.A(net215),
    .B(_0742_),
    .Y(_0763_));
 sg13g2_xor2_1 _1482_ (.B(_0742_),
    .A(net215),
    .X(\i_game_and_vga.i_game_top.sprite_target.sprite_display.x_sprite_plus_w_1[6] ));
 sg13g2_nor2_1 _1483_ (.A(_0022_),
    .B(\i_game_and_vga.i_game_top.sprite_target.sprite_display.x_sprite_plus_w_1[5] ),
    .Y(_0764_));
 sg13g2_and3_1 _1484_ (.X(_0765_),
    .A(\i_game_and_vga.i_game_top.sprite_target.pixel_x[5] ),
    .B(_0022_),
    .C(\i_game_and_vga.i_game_top.sprite_target.sprite_display.x_sprite_plus_w_1[5] ));
 sg13g2_xnor2_1 _1485_ (.Y(_0766_),
    .A(_0021_),
    .B(\i_game_and_vga.i_game_top.sprite_target.sprite_display.x_sprite_plus_w_1[6] ));
 sg13g2_nor3_1 _1486_ (.A(_0764_),
    .B(_0765_),
    .C(_0766_),
    .Y(_0767_));
 sg13g2_xnor2_1 _1487_ (.Y(_0768_),
    .A(net406),
    .B(_0763_));
 sg13g2_inv_1 _1488_ (.Y(\i_game_and_vga.i_game_top.sprite_target.sprite_display.x_sprite_plus_w_1[7] ),
    .A(_0768_));
 sg13g2_nor2_1 _1489_ (.A(\i_game_and_vga.i_game_top.sprite_target.pixel_x[7] ),
    .B(_0768_),
    .Y(_0769_));
 sg13g2_a221oi_1 _1490_ (.B2(_0762_),
    .C1(_0769_),
    .B1(_0767_),
    .A1(_0547_),
    .Y(_0770_),
    .A2(\i_game_and_vga.i_game_top.sprite_target.sprite_display.x_sprite_plus_w_1[6] ));
 sg13g2_a22oi_1 _1491_ (.Y(_0771_),
    .B1(_0768_),
    .B2(\i_game_and_vga.i_game_top.sprite_target.pixel_x[7] ),
    .A2(\i_game_and_vga.i_game_top.sprite_target.sprite_display.x_sprite_plus_w_1[8] ),
    .A1(_0019_));
 sg13g2_o21ai_1 _1492_ (.B1(_0771_),
    .Y(_0772_),
    .A1(_0019_),
    .A2(\i_game_and_vga.i_game_top.sprite_target.sprite_display.x_sprite_plus_w_1[8] ));
 sg13g2_o21ai_1 _1493_ (.B1(_0748_),
    .Y(_0773_),
    .A1(_0770_),
    .A2(_0772_));
 sg13g2_o21ai_1 _1494_ (.B1(_0745_),
    .Y(_0774_),
    .A1(net304),
    .A2(_0746_));
 sg13g2_a21oi_2 _1495_ (.B1(_0774_),
    .Y(_0775_),
    .A2(_0773_),
    .A1(_0747_));
 sg13g2_nand2_1 _1496_ (.Y(_0776_),
    .A(_0543_),
    .B(net299));
 sg13g2_nor2_1 _1497_ (.A(_0553_),
    .B(\i_game_and_vga.i_game_top.sprite_target.sprite_control.sprite_x[2] ),
    .Y(_0777_));
 sg13g2_nand2_1 _1498_ (.Y(_0778_),
    .A(_0553_),
    .B(\i_game_and_vga.i_game_top.sprite_target.sprite_control.sprite_x[2] ));
 sg13g2_nand2b_1 _1499_ (.Y(_0779_),
    .B(_0778_),
    .A_N(_0777_));
 sg13g2_a221oi_1 _1500_ (.B2(_0778_),
    .C1(_0777_),
    .B1(_0753_),
    .A1(\i_game_and_vga.i_game_top.sprite_target.pixel_x[3] ),
    .Y(_0780_),
    .A2(_0573_));
 sg13g2_nand2b_1 _1501_ (.Y(_0781_),
    .B(net300),
    .A_N(\i_game_and_vga.i_game_top.sprite_target.pixel_x[4] ));
 sg13g2_o21ai_1 _1502_ (.B1(_0781_),
    .Y(_0782_),
    .A1(\i_game_and_vga.i_game_top.sprite_target.pixel_x[3] ),
    .A2(_0573_));
 sg13g2_a22oi_1 _1503_ (.Y(_0783_),
    .B1(_0572_),
    .B2(\i_game_and_vga.i_game_top.sprite_target.pixel_x[4] ),
    .A2(_0571_),
    .A1(\i_game_and_vga.i_game_top.sprite_target.pixel_x[5] ));
 sg13g2_o21ai_1 _1504_ (.B1(_0783_),
    .Y(_0784_),
    .A1(_0780_),
    .A2(_0782_));
 sg13g2_a22oi_1 _1505_ (.Y(_0785_),
    .B1(\i_game_and_vga.i_game_top.sprite_target.sprite_control.sprite_x[5] ),
    .B2(_0549_),
    .A2(\i_game_and_vga.i_game_top.sprite_target.sprite_control.sprite_x[6] ),
    .A1(_0547_));
 sg13g2_a22oi_1 _1506_ (.Y(_0786_),
    .B1(_0784_),
    .B2(_0785_),
    .A2(_0570_),
    .A1(\i_game_and_vga.i_game_top.sprite_target.pixel_x[6] ));
 sg13g2_a21oi_1 _1507_ (.A1(_0545_),
    .A2(\i_game_and_vga.i_game_top.sprite_target.sprite_control.sprite_x[7] ),
    .Y(_0787_),
    .B1(_0786_));
 sg13g2_a21o_1 _1508_ (.A2(_0569_),
    .A1(\i_game_and_vga.i_game_top.sprite_target.pixel_x[7] ),
    .B1(_0787_),
    .X(_0788_));
 sg13g2_nand2b_1 _1509_ (.Y(_0789_),
    .B(\i_game_and_vga.i_game_top.sprite_target.pixel_x[8] ),
    .A_N(net299));
 sg13g2_o21ai_1 _1510_ (.B1(_0789_),
    .Y(_0790_),
    .A1(_0540_),
    .A2(net298));
 sg13g2_a21oi_2 _1511_ (.B1(_0790_),
    .Y(_0791_),
    .A2(_0788_),
    .A1(_0776_));
 sg13g2_xnor2_1 _1512_ (.Y(\i_game_and_vga.i_game_top.sprite_target.sprite_display.y_sprite_plus_h_1[5] ),
    .A(net79),
    .B(_0636_));
 sg13g2_o21ai_1 _1513_ (.B1(net80),
    .Y(_0792_),
    .A1(net310),
    .A2(net157));
 sg13g2_nand2_1 _1514_ (.Y(\i_game_and_vga.i_game_top.sprite_target.sprite_display.y_sprite_plus_h_1[2] ),
    .A(_0635_),
    .B(_0792_));
 sg13g2_nand2b_1 _1515_ (.Y(_0793_),
    .B(net313),
    .A_N(net310));
 sg13g2_nor2b_1 _1516_ (.A(net313),
    .B_N(net310),
    .Y(_0794_));
 sg13g2_nor2b_1 _1517_ (.A(\i_game_and_vga.i_game_top.sprite_target.pixel_y[0] ),
    .B_N(\i_game_and_vga.i_game_top.sprite_target.sprite_control.sprite_y[0] ),
    .Y(_0795_));
 sg13g2_o21ai_1 _1518_ (.B1(_0793_),
    .Y(_0796_),
    .A1(_0794_),
    .A2(_0795_));
 sg13g2_o21ai_1 _1519_ (.B1(_0796_),
    .Y(_0797_),
    .A1(net310),
    .A2(\i_game_and_vga.i_game_top.sprite_target.sprite_control.sprite_y[0] ));
 sg13g2_xor2_1 _1520_ (.B(\i_game_and_vga.i_game_top.sprite_target.sprite_display.y_sprite_plus_h_1[2] ),
    .A(_0030_),
    .X(_0798_));
 sg13g2_xnor2_1 _1521_ (.Y(\i_game_and_vga.i_game_top.sprite_target.sprite_display.y_sprite_plus_h_1[3] ),
    .A(_0577_),
    .B(_0635_));
 sg13g2_and2_1 _1522_ (.A(_0565_),
    .B(\i_game_and_vga.i_game_top.sprite_target.sprite_display.y_sprite_plus_h_1[3] ),
    .X(_0799_));
 sg13g2_a221oi_1 _1523_ (.B2(_0798_),
    .C1(_0799_),
    .B1(_0797_),
    .A1(_0566_),
    .Y(_0800_),
    .A2(\i_game_and_vga.i_game_top.sprite_target.sprite_display.y_sprite_plus_h_1[2] ));
 sg13g2_a21o_1 _1524_ (.A2(_0635_),
    .A1(net68),
    .B1(net78),
    .X(_0801_));
 sg13g2_and2_1 _1525_ (.A(_0636_),
    .B(_0801_),
    .X(\i_game_and_vga.i_game_top.sprite_target.sprite_display.y_sprite_plus_h_1[4] ));
 sg13g2_nand2b_1 _1526_ (.Y(_0802_),
    .B(net312),
    .A_N(\i_game_and_vga.i_game_top.sprite_target.sprite_display.y_sprite_plus_h_1[3] ));
 sg13g2_o21ai_1 _1527_ (.B1(_0802_),
    .Y(_0803_),
    .A1(_0029_),
    .A2(\i_game_and_vga.i_game_top.sprite_target.sprite_display.y_sprite_plus_h_1[4] ));
 sg13g2_nand2_1 _1528_ (.Y(_0804_),
    .A(_0029_),
    .B(\i_game_and_vga.i_game_top.sprite_target.sprite_display.y_sprite_plus_h_1[4] ));
 sg13g2_o21ai_1 _1529_ (.B1(_0804_),
    .Y(_0805_),
    .A1(_0800_),
    .A2(_0803_));
 sg13g2_xor2_1 _1530_ (.B(\i_game_and_vga.i_game_top.sprite_target.sprite_display.y_sprite_plus_h_1[5] ),
    .A(_0028_),
    .X(_0806_));
 sg13g2_a22oi_1 _1531_ (.Y(_0807_),
    .B1(_0805_),
    .B2(_0806_),
    .A2(\i_game_and_vga.i_game_top.sprite_target.sprite_display.y_sprite_plus_h_1[5] ),
    .A1(_0561_));
 sg13g2_nand2_1 _1532_ (.Y(_0808_),
    .A(_0574_),
    .B(_0637_));
 sg13g2_nand3_1 _1533_ (.B(_0035_),
    .C(_0808_),
    .A(_0027_),
    .Y(_0809_));
 sg13g2_nor2b_1 _1534_ (.A(\i_game_and_vga.i_game_top.sprite_target.sprite_display.y_sprite_plus_h_1[7] ),
    .B_N(_0808_),
    .Y(\i_game_and_vga.i_game_top.sprite_target.sprite_display.y_sprite_plus_h_1[6] ));
 sg13g2_o21ai_1 _1535_ (.B1(_0809_),
    .Y(_0810_),
    .A1(_0027_),
    .A2(\i_game_and_vga.i_game_top.sprite_target.sprite_display.y_sprite_plus_h_1[6] ));
 sg13g2_o21ai_1 _1536_ (.B1(_0637_),
    .Y(_0811_),
    .A1(\i_game_and_vga.i_game_top.sprite_target.pixel_y[6] ),
    .A2(_0574_));
 sg13g2_nand2_1 _1537_ (.Y(_0812_),
    .A(\i_game_and_vga.i_game_top.sprite_target.pixel_y[6] ),
    .B(_0574_));
 sg13g2_nand3_1 _1538_ (.B(_0811_),
    .C(_0812_),
    .A(_0035_),
    .Y(_0813_));
 sg13g2_o21ai_1 _1539_ (.B1(_0813_),
    .Y(_0814_),
    .A1(_0807_),
    .A2(_0810_));
 sg13g2_nor2_1 _1540_ (.A(_0566_),
    .B(\i_game_and_vga.i_game_top.sprite_target.sprite_control.sprite_y[2] ),
    .Y(_0815_));
 sg13g2_xnor2_1 _1541_ (.Y(_0816_),
    .A(\i_game_and_vga.i_game_top.sprite_target.pixel_y[2] ),
    .B(\i_game_and_vga.i_game_top.sprite_target.sprite_control.sprite_y[2] ));
 sg13g2_a221oi_1 _1542_ (.B2(_0816_),
    .C1(_0815_),
    .B1(_0796_),
    .A1(\i_game_and_vga.i_game_top.sprite_target.pixel_y[3] ),
    .Y(_0817_),
    .A2(_0577_));
 sg13g2_a221oi_1 _1543_ (.B2(_0565_),
    .C1(_0817_),
    .B1(\i_game_and_vga.i_game_top.sprite_target.sprite_control.sprite_y[3] ),
    .A1(_0562_),
    .Y(_0818_),
    .A2(\i_game_and_vga.i_game_top.sprite_target.sprite_control.sprite_y[4] ));
 sg13g2_a221oi_1 _1544_ (.B2(\i_game_and_vga.i_game_top.sprite_target.pixel_y[4] ),
    .C1(_0818_),
    .B1(_0576_),
    .A1(\i_game_and_vga.i_game_top.sprite_target.pixel_y[5] ),
    .Y(_0819_),
    .A2(_0575_));
 sg13g2_a22oi_1 _1545_ (.Y(_0820_),
    .B1(\i_game_and_vga.i_game_top.sprite_target.sprite_control.sprite_y[5] ),
    .B2(_0561_),
    .A2(\i_game_and_vga.i_game_top.sprite_target.sprite_control.sprite_y[6] ),
    .A1(_0559_));
 sg13g2_nand3b_1 _1546_ (.B(_0820_),
    .C(_0035_),
    .Y(_0821_),
    .A_N(_0819_));
 sg13g2_nand4_1 _1547_ (.B(_0034_),
    .C(_0812_),
    .A(_0557_),
    .Y(_0822_),
    .D(_0821_));
 sg13g2_nor2_1 _1548_ (.A(_0035_),
    .B(\i_game_and_vga.i_game_top.sprite_target.sprite_display.y_sprite_plus_h_1[7] ),
    .Y(_0823_));
 sg13g2_a21oi_1 _1549_ (.A1(_0540_),
    .A2(net298),
    .Y(_0824_),
    .B1(_0823_));
 sg13g2_nand4_1 _1550_ (.B(_0814_),
    .C(_0822_),
    .A(_0555_),
    .Y(_0825_),
    .D(_0824_));
 sg13g2_nor3_1 _1551_ (.A(_0775_),
    .B(_0791_),
    .C(_0825_),
    .Y(_0826_));
 sg13g2_xor2_1 _1552_ (.B(net302),
    .A(\i_game_and_vga.i_game_top.sprite_target.pixel_x[1] ),
    .X(_0827_));
 sg13g2_nor2b_1 _1553_ (.A(net303),
    .B_N(\i_game_and_vga.i_game_top.sprite_target.pixel_x[0] ),
    .Y(_0828_));
 sg13g2_xnor2_1 _1554_ (.Y(_0829_),
    .A(_0827_),
    .B(_0828_));
 sg13g2_nor2_1 _1555_ (.A(_0752_),
    .B(_0828_),
    .Y(_0830_));
 sg13g2_xnor2_1 _1556_ (.Y(_0831_),
    .A(_0753_),
    .B(_0779_));
 sg13g2_xnor2_1 _1557_ (.Y(_0832_),
    .A(_0830_),
    .B(_0831_));
 sg13g2_nand2_1 _1558_ (.Y(_0833_),
    .A(_0829_),
    .B(_0832_));
 sg13g2_xnor2_1 _1559_ (.Y(_0834_),
    .A(_0796_),
    .B(_0816_));
 sg13g2_xor2_1 _1560_ (.B(net310),
    .A(net313),
    .X(_0835_));
 sg13g2_nor2_1 _1561_ (.A(_0795_),
    .B(_0835_),
    .Y(_0836_));
 sg13g2_nand2b_1 _1562_ (.Y(_0837_),
    .B(\i_game_and_vga.i_game_top.sprite_target.pixel_y[0] ),
    .A_N(\i_game_and_vga.i_game_top.sprite_target.sprite_control.sprite_y[0] ));
 sg13g2_nand2_1 _1563_ (.Y(_0838_),
    .A(_0836_),
    .B(_0837_));
 sg13g2_a21o_1 _1564_ (.A2(_0837_),
    .A1(_0835_),
    .B1(_0836_),
    .X(_0839_));
 sg13g2_mux2_1 _1565_ (.A0(_0838_),
    .A1(_0839_),
    .S(_0834_),
    .X(_0840_));
 sg13g2_nand2_1 _1566_ (.Y(_0841_),
    .A(_0833_),
    .B(_0840_));
 sg13g2_and2_1 _1567_ (.A(_0826_),
    .B(_0841_),
    .X(_0005_));
 sg13g2_nor2b_1 _1568_ (.A(\i_game_and_vga.i_game_top.sprite_target.pixel_y[0] ),
    .B_N(net294),
    .Y(_0842_));
 sg13g2_nand2b_1 _1569_ (.Y(_0843_),
    .B(net313),
    .A_N(net292));
 sg13g2_nor2b_1 _1570_ (.A(net313),
    .B_N(net292),
    .Y(_0844_));
 sg13g2_xnor2_1 _1571_ (.Y(_0845_),
    .A(net292),
    .B(net313));
 sg13g2_or2_1 _1572_ (.X(_0846_),
    .B(_0845_),
    .A(_0842_));
 sg13g2_nor2_1 _1573_ (.A(net291),
    .B(_0566_),
    .Y(_0847_));
 sg13g2_a21oi_2 _1574_ (.B1(_0844_),
    .Y(_0848_),
    .A2(_0843_),
    .A1(_0842_));
 sg13g2_nand2_1 _1575_ (.Y(_0849_),
    .A(net291),
    .B(_0566_));
 sg13g2_nor2b_1 _1576_ (.A(_0847_),
    .B_N(_0849_),
    .Y(_0850_));
 sg13g2_mux2_1 _1577_ (.A0(_0844_),
    .A1(_0848_),
    .S(_0850_),
    .X(_0851_));
 sg13g2_nor2b_1 _1578_ (.A(\i_game_and_vga.i_game_top.sprite_target.pixel_x[0] ),
    .B_N(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.sprite_x[0] ),
    .Y(_0852_));
 sg13g2_xnor2_1 _1579_ (.Y(_0853_),
    .A(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.sprite_x[0] ),
    .B(\i_game_and_vga.i_game_top.sprite_target.pixel_x[0] ));
 sg13g2_nor2_1 _1580_ (.A(net286),
    .B(_0553_),
    .Y(_0854_));
 sg13g2_xnor2_1 _1581_ (.Y(_0855_),
    .A(net286),
    .B(\i_game_and_vga.i_game_top.sprite_target.pixel_x[2] ));
 sg13g2_nor2b_1 _1582_ (.A(\i_game_and_vga.i_game_top.sprite_target.pixel_x[1] ),
    .B_N(net287),
    .Y(_0856_));
 sg13g2_nand2b_1 _1583_ (.Y(_0857_),
    .B(\i_game_and_vga.i_game_top.sprite_target.pixel_x[1] ),
    .A_N(net287));
 sg13g2_o21ai_1 _1584_ (.B1(_0857_),
    .Y(_0858_),
    .A1(_0852_),
    .A2(_0856_));
 sg13g2_xnor2_1 _1585_ (.Y(_0859_),
    .A(_0855_),
    .B(_0858_));
 sg13g2_and2_1 _1586_ (.A(_0853_),
    .B(_0859_),
    .X(_0860_));
 sg13g2_nor2b_2 _1587_ (.A(_0856_),
    .B_N(_0857_),
    .Y(_0861_));
 sg13g2_inv_1 _1588_ (.Y(_0862_),
    .A(_0861_));
 sg13g2_xor2_1 _1589_ (.B(_0861_),
    .A(_0852_),
    .X(_0863_));
 sg13g2_inv_1 _1590_ (.Y(_0864_),
    .A(_0863_));
 sg13g2_nor2_1 _1591_ (.A(_0853_),
    .B(_0859_),
    .Y(_0865_));
 sg13g2_a22oi_1 _1592_ (.Y(_0866_),
    .B1(_0863_),
    .B2(_0865_),
    .A2(_0862_),
    .A1(_0860_));
 sg13g2_xnor2_1 _1593_ (.Y(_0867_),
    .A(net294),
    .B(\i_game_and_vga.i_game_top.sprite_target.pixel_y[0] ));
 sg13g2_xnor2_1 _1594_ (.Y(_0868_),
    .A(_0848_),
    .B(_0850_));
 sg13g2_nand2_1 _1595_ (.Y(_0869_),
    .A(_0867_),
    .B(_0868_));
 sg13g2_nand2_1 _1596_ (.Y(_0870_),
    .A(_0866_),
    .B(_0869_));
 sg13g2_a22oi_1 _1597_ (.Y(_0871_),
    .B1(_0864_),
    .B2(_0859_),
    .A2(_0861_),
    .A1(_0853_));
 sg13g2_nand2b_1 _1598_ (.Y(_0872_),
    .B(_0871_),
    .A_N(_0865_));
 sg13g2_a22oi_1 _1599_ (.Y(_0873_),
    .B1(_0870_),
    .B2(_0872_),
    .A2(_0851_),
    .A1(_0846_));
 sg13g2_or2_1 _1600_ (.X(_0874_),
    .B(_0871_),
    .A(_0860_));
 sg13g2_nand2_1 _1601_ (.Y(_0875_),
    .A(_0845_),
    .B(_0867_));
 sg13g2_nand2_1 _1602_ (.Y(_0876_),
    .A(_0868_),
    .B(_0875_));
 sg13g2_o21ai_1 _1603_ (.B1(_0874_),
    .Y(_0877_),
    .A1(_0866_),
    .A2(_0876_));
 sg13g2_or2_1 _1604_ (.X(_0878_),
    .B(_0877_),
    .A(_0873_));
 sg13g2_nor2_1 _1605_ (.A(net287),
    .B(net288),
    .Y(_0879_));
 sg13g2_nor3_1 _1606_ (.A(net286),
    .B(net287),
    .C(net288),
    .Y(_0880_));
 sg13g2_or3_1 _1607_ (.A(net286),
    .B(net287),
    .C(net288),
    .X(_0881_));
 sg13g2_nand3_1 _1608_ (.B(net285),
    .C(_0881_),
    .A(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.sprite_x[4] ),
    .Y(_0882_));
 sg13g2_nand4_1 _1609_ (.B(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.sprite_x[4] ),
    .C(net285),
    .A(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.sprite_x[5] ),
    .Y(_0883_),
    .D(_0881_));
 sg13g2_nand2_1 _1610_ (.Y(_0884_),
    .A(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.sprite_x[7] ),
    .B(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.sprite_x[6] ));
 sg13g2_nor2_1 _1611_ (.A(_0883_),
    .B(_0884_),
    .Y(_0885_));
 sg13g2_nor3_1 _1612_ (.A(_0542_),
    .B(_0883_),
    .C(_0884_),
    .Y(_0886_));
 sg13g2_nand2_1 _1613_ (.Y(_0887_),
    .A(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.sprite_x[9] ),
    .B(_0886_));
 sg13g2_xnor2_1 _1614_ (.Y(_0888_),
    .A(_0548_),
    .B(_0882_));
 sg13g2_inv_1 _1615_ (.Y(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_display.x_sprite_plus_w_1[5] ),
    .A(_0888_));
 sg13g2_xnor2_1 _1616_ (.Y(_0889_),
    .A(_0022_),
    .B(_0888_));
 sg13g2_xor2_1 _1617_ (.B(_0879_),
    .A(net286),
    .X(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_display.x_sprite_plus_w_1[2] ));
 sg13g2_nor2b_1 _1618_ (.A(_0879_),
    .B_N(_0858_),
    .Y(_0890_));
 sg13g2_xnor2_1 _1619_ (.Y(_0891_),
    .A(_0024_),
    .B(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_display.x_sprite_plus_w_1[2] ));
 sg13g2_xnor2_1 _1620_ (.Y(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_display.x_sprite_plus_w_1[3] ),
    .A(net285),
    .B(_0880_));
 sg13g2_a22oi_1 _1621_ (.Y(_0892_),
    .B1(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_display.x_sprite_plus_w_1[3] ),
    .B2(_0552_),
    .A2(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_display.x_sprite_plus_w_1[2] ),
    .A1(_0553_));
 sg13g2_o21ai_1 _1622_ (.B1(_0892_),
    .Y(_0893_),
    .A1(_0890_),
    .A2(_0891_));
 sg13g2_o21ai_1 _1623_ (.B1(_0550_),
    .Y(_0894_),
    .A1(_0551_),
    .A2(_0880_));
 sg13g2_and2_2 _1624_ (.A(_0882_),
    .B(_0894_),
    .X(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_display.x_sprite_plus_w_1[4] ));
 sg13g2_nand2b_1 _1625_ (.Y(_0895_),
    .B(\i_game_and_vga.i_game_top.sprite_target.pixel_x[3] ),
    .A_N(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_display.x_sprite_plus_w_1[3] ));
 sg13g2_and2_1 _1626_ (.A(_0023_),
    .B(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_display.x_sprite_plus_w_1[4] ),
    .X(_0896_));
 sg13g2_xor2_1 _1627_ (.B(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_display.x_sprite_plus_w_1[4] ),
    .A(_0023_),
    .X(_0897_));
 sg13g2_nand4_1 _1628_ (.B(_0893_),
    .C(_0895_),
    .A(_0889_),
    .Y(_0898_),
    .D(_0897_));
 sg13g2_a22oi_1 _1629_ (.Y(_0899_),
    .B1(_0889_),
    .B2(_0896_),
    .A2(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_display.x_sprite_plus_w_1[5] ),
    .A1(_0549_));
 sg13g2_nor2_1 _1630_ (.A(net391),
    .B(_0883_),
    .Y(_0900_));
 sg13g2_xor2_1 _1631_ (.B(_0883_),
    .A(net391),
    .X(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_display.x_sprite_plus_w_1[6] ));
 sg13g2_nand2b_1 _1632_ (.Y(_0901_),
    .B(_0021_),
    .A_N(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_display.x_sprite_plus_w_1[6] ));
 sg13g2_nand2b_1 _1633_ (.Y(_0902_),
    .B(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_display.x_sprite_plus_w_1[6] ),
    .A_N(_0021_));
 sg13g2_xnor2_1 _1634_ (.Y(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_display.x_sprite_plus_w_1[7] ),
    .A(_0544_),
    .B(_0900_));
 sg13g2_nor2_1 _1635_ (.A(_0545_),
    .B(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_display.x_sprite_plus_w_1[7] ),
    .Y(_0903_));
 sg13g2_xnor2_1 _1636_ (.Y(_0904_),
    .A(_0545_),
    .B(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_display.x_sprite_plus_w_1[7] ));
 sg13g2_a221oi_1 _1637_ (.B2(_0902_),
    .C1(_0904_),
    .B1(_0901_),
    .A1(_0898_),
    .Y(_0905_),
    .A2(_0899_));
 sg13g2_a22oi_1 _1638_ (.Y(_0906_),
    .B1(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_display.x_sprite_plus_w_1[7] ),
    .B2(_0545_),
    .A2(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_display.x_sprite_plus_w_1[6] ),
    .A1(_0547_));
 sg13g2_nor2_1 _1639_ (.A(_0903_),
    .B(_0906_),
    .Y(_0907_));
 sg13g2_xnor2_1 _1640_ (.Y(_0908_),
    .A(net91),
    .B(_0886_));
 sg13g2_inv_1 _1641_ (.Y(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_display.x_sprite_plus_w_1[9] ),
    .A(_0908_));
 sg13g2_nand2_1 _1642_ (.Y(_0909_),
    .A(\i_game_and_vga.i_game_top.sprite_target.pixel_x[9] ),
    .B(_0908_));
 sg13g2_xnor2_1 _1643_ (.Y(_0910_),
    .A(net417),
    .B(_0885_));
 sg13g2_inv_1 _1644_ (.Y(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_display.x_sprite_plus_w_1[8] ),
    .A(_0910_));
 sg13g2_xnor2_1 _1645_ (.Y(_0911_),
    .A(_0019_),
    .B(_0910_));
 sg13g2_and2_1 _1646_ (.A(_0909_),
    .B(_0911_),
    .X(_0912_));
 sg13g2_o21ai_1 _1647_ (.B1(_0912_),
    .Y(_0913_),
    .A1(_0905_),
    .A2(_0907_));
 sg13g2_nor2_1 _1648_ (.A(\i_game_and_vga.i_game_top.sprite_target.pixel_x[9] ),
    .B(_0908_),
    .Y(_0914_));
 sg13g2_nor2_1 _1649_ (.A(\i_game_and_vga.i_game_top.sprite_target.pixel_x[8] ),
    .B(_0910_),
    .Y(_0915_));
 sg13g2_o21ai_1 _1650_ (.B1(_0909_),
    .Y(_0916_),
    .A1(_0914_),
    .A2(_0915_));
 sg13g2_nand3_1 _1651_ (.B(_0913_),
    .C(_0916_),
    .A(_0887_),
    .Y(_0917_));
 sg13g2_a21o_2 _1652_ (.A2(_0916_),
    .A1(_0913_),
    .B1(_0887_),
    .X(_0918_));
 sg13g2_xnor2_1 _1653_ (.Y(_0919_),
    .A(_0560_),
    .B(_0725_));
 sg13g2_inv_1 _1654_ (.Y(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_display.y_sprite_plus_h_1[5] ),
    .A(_0919_));
 sg13g2_xnor2_1 _1655_ (.Y(_0920_),
    .A(_0028_),
    .B(_0919_));
 sg13g2_xor2_1 _1656_ (.B(_0722_),
    .A(net291),
    .X(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_display.y_sprite_plus_h_1[2] ));
 sg13g2_nor2b_1 _1657_ (.A(_0722_),
    .B_N(_0848_),
    .Y(_0921_));
 sg13g2_xnor2_1 _1658_ (.Y(_0922_),
    .A(_0030_),
    .B(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_display.y_sprite_plus_h_1[2] ));
 sg13g2_xnor2_1 _1659_ (.Y(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_display.y_sprite_plus_h_1[3] ),
    .A(net290),
    .B(_0723_));
 sg13g2_a22oi_1 _1660_ (.Y(_0923_),
    .B1(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_display.y_sprite_plus_h_1[3] ),
    .B2(_0565_),
    .A2(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_display.y_sprite_plus_h_1[2] ),
    .A1(_0566_));
 sg13g2_o21ai_1 _1661_ (.B1(_0923_),
    .Y(_0924_),
    .A1(_0921_),
    .A2(_0922_));
 sg13g2_o21ai_1 _1662_ (.B1(_0563_),
    .Y(_0925_),
    .A1(_0564_),
    .A2(_0723_));
 sg13g2_and2_1 _1663_ (.A(_0725_),
    .B(_0925_),
    .X(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_display.y_sprite_plus_h_1[4] ));
 sg13g2_and2_1 _1664_ (.A(_0029_),
    .B(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_display.y_sprite_plus_h_1[4] ),
    .X(_0926_));
 sg13g2_nand2b_1 _1665_ (.Y(_0927_),
    .B(net312),
    .A_N(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_display.y_sprite_plus_h_1[3] ));
 sg13g2_xor2_1 _1666_ (.B(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_display.y_sprite_plus_h_1[4] ),
    .A(_0029_),
    .X(_0928_));
 sg13g2_nand4_1 _1667_ (.B(_0924_),
    .C(_0927_),
    .A(_0920_),
    .Y(_0929_),
    .D(_0928_));
 sg13g2_a22oi_1 _1668_ (.Y(_0930_),
    .B1(_0920_),
    .B2(_0926_),
    .A2(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_display.y_sprite_plus_h_1[5] ),
    .A1(_0561_));
 sg13g2_nor2_1 _1669_ (.A(net185),
    .B(_0726_),
    .Y(_0931_));
 sg13g2_xnor2_1 _1670_ (.Y(_0932_),
    .A(net409),
    .B(_0931_));
 sg13g2_inv_1 _1671_ (.Y(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_display.y_sprite_plus_h_1[7] ),
    .A(_0932_));
 sg13g2_xor2_1 _1672_ (.B(_0726_),
    .A(net185),
    .X(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_display.y_sprite_plus_h_1[6] ));
 sg13g2_xnor2_1 _1673_ (.Y(_0933_),
    .A(_0027_),
    .B(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_display.y_sprite_plus_h_1[6] ));
 sg13g2_a21o_1 _1674_ (.A2(_0932_),
    .A1(net311),
    .B1(_0933_),
    .X(_0934_));
 sg13g2_nor2_1 _1675_ (.A(net311),
    .B(_0932_),
    .Y(_0935_));
 sg13g2_a221oi_1 _1676_ (.B2(_0557_),
    .C1(_0934_),
    .B1(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_display.y_sprite_plus_h_1[7] ),
    .A1(_0929_),
    .Y(_0936_),
    .A2(_0930_));
 sg13g2_nand2_1 _1677_ (.Y(_0937_),
    .A(_0559_),
    .B(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_display.y_sprite_plus_h_1[6] ));
 sg13g2_a21oi_1 _1678_ (.A1(net311),
    .A2(_0932_),
    .Y(_0938_),
    .B1(_0937_));
 sg13g2_o21ai_1 _1679_ (.B1(net252),
    .Y(_0939_),
    .A1(_0721_),
    .A2(_0726_));
 sg13g2_nand2b_1 _1680_ (.Y(_0940_),
    .B(_0939_),
    .A_N(_0727_));
 sg13g2_inv_1 _1681_ (.Y(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_display.y_sprite_plus_h_1[8] ),
    .A(_0940_));
 sg13g2_nor2_1 _1682_ (.A(\i_game_and_vga.i_game_top.sprite_target.pixel_y[8] ),
    .B(_0940_),
    .Y(_0941_));
 sg13g2_or3_1 _1683_ (.A(_0935_),
    .B(_0938_),
    .C(_0941_),
    .X(_0942_));
 sg13g2_nand2_1 _1684_ (.Y(_0943_),
    .A(\i_game_and_vga.i_game_top.sprite_target.pixel_y[8] ),
    .B(_0940_));
 sg13g2_o21ai_1 _1685_ (.B1(_0943_),
    .Y(_0944_),
    .A1(_0936_),
    .A2(_0942_));
 sg13g2_nor2_1 _1686_ (.A(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.sprite_x[7] ),
    .B(_0545_),
    .Y(_0945_));
 sg13g2_a22oi_1 _1687_ (.Y(_0946_),
    .B1(net286),
    .B2(_0553_),
    .A2(_0552_),
    .A1(net285));
 sg13g2_o21ai_1 _1688_ (.B1(_0946_),
    .Y(_0947_),
    .A1(_0854_),
    .A2(_0858_));
 sg13g2_a22oi_1 _1689_ (.Y(_0948_),
    .B1(_0551_),
    .B2(\i_game_and_vga.i_game_top.sprite_target.pixel_x[3] ),
    .A2(_0550_),
    .A1(\i_game_and_vga.i_game_top.sprite_target.pixel_x[4] ));
 sg13g2_nand2_1 _1690_ (.Y(_0949_),
    .A(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.sprite_x[5] ),
    .B(_0549_));
 sg13g2_o21ai_1 _1691_ (.B1(_0949_),
    .Y(_0950_),
    .A1(\i_game_and_vga.i_game_top.sprite_target.pixel_x[4] ),
    .A2(_0550_));
 sg13g2_a21o_1 _1692_ (.A2(_0948_),
    .A1(_0947_),
    .B1(_0950_),
    .X(_0951_));
 sg13g2_a22oi_1 _1693_ (.Y(_0952_),
    .B1(_0548_),
    .B2(\i_game_and_vga.i_game_top.sprite_target.pixel_x[5] ),
    .A2(\i_game_and_vga.i_game_top.sprite_target.pixel_x[6] ),
    .A1(_0546_));
 sg13g2_a22oi_1 _1694_ (.Y(_0953_),
    .B1(_0951_),
    .B2(_0952_),
    .A2(_0547_),
    .A1(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.sprite_x[6] ));
 sg13g2_a22oi_1 _1695_ (.Y(_0954_),
    .B1(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.sprite_x[7] ),
    .B2(_0545_),
    .A2(_0543_),
    .A1(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.sprite_x[8] ));
 sg13g2_o21ai_1 _1696_ (.B1(_0954_),
    .Y(_0955_),
    .A1(_0945_),
    .A2(_0953_));
 sg13g2_a22oi_1 _1697_ (.Y(_0956_),
    .B1(_0542_),
    .B2(\i_game_and_vga.i_game_top.sprite_target.pixel_x[8] ),
    .A2(_0541_),
    .A1(net304));
 sg13g2_nand2_1 _1698_ (.Y(_0957_),
    .A(_0554_),
    .B(\i_game_and_vga.i_game_top.sprite_target.pixel_y[8] ));
 sg13g2_nor2_1 _1699_ (.A(_0562_),
    .B(net289),
    .Y(_0958_));
 sg13g2_a221oi_1 _1700_ (.B2(_0849_),
    .C1(_0847_),
    .B1(_0848_),
    .A1(_0564_),
    .Y(_0959_),
    .A2(net312));
 sg13g2_a21oi_1 _1701_ (.A1(net290),
    .A2(_0565_),
    .Y(_0960_),
    .B1(_0959_));
 sg13g2_a22oi_1 _1702_ (.Y(_0961_),
    .B1(_0562_),
    .B2(net289),
    .A2(_0561_),
    .A1(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.sprite_y[5] ));
 sg13g2_o21ai_1 _1703_ (.B1(_0961_),
    .Y(_0962_),
    .A1(_0958_),
    .A2(_0960_));
 sg13g2_a22oi_1 _1704_ (.Y(_0963_),
    .B1(_0560_),
    .B2(\i_game_and_vga.i_game_top.sprite_target.pixel_y[5] ),
    .A2(\i_game_and_vga.i_game_top.sprite_target.pixel_y[6] ),
    .A1(_0558_));
 sg13g2_a22oi_1 _1705_ (.Y(_0964_),
    .B1(_0962_),
    .B2(_0963_),
    .A2(_0559_),
    .A1(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.sprite_y[6] ));
 sg13g2_nor2_1 _1706_ (.A(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.sprite_y[7] ),
    .B(_0557_),
    .Y(_0965_));
 sg13g2_a22oi_1 _1707_ (.Y(_0966_),
    .B1(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.sprite_y[7] ),
    .B2(_0557_),
    .A2(_0555_),
    .A1(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.sprite_y[8] ));
 sg13g2_o21ai_1 _1708_ (.B1(_0966_),
    .Y(_0967_),
    .A1(_0964_),
    .A2(_0965_));
 sg13g2_nor2_1 _1709_ (.A(net304),
    .B(_0541_),
    .Y(_0968_));
 sg13g2_a21o_1 _1710_ (.A2(_0956_),
    .A1(_0955_),
    .B1(_0968_),
    .X(_0969_));
 sg13g2_a221oi_1 _1711_ (.B2(_0967_),
    .C1(_0969_),
    .B1(_0957_),
    .A1(_0728_),
    .Y(_0970_),
    .A2(_0944_));
 sg13g2_and4_1 _1712_ (.A(_0878_),
    .B(_0917_),
    .C(_0918_),
    .D(_0970_),
    .X(_0007_));
 sg13g2_or2_1 _1713_ (.X(_0971_),
    .B(net201),
    .A(\i_game_and_vga.i_game_top.timer.counter[11] ));
 sg13g2_nor4_2 _1714_ (.A(\i_game_and_vga.i_game_top.timer.counter[13] ),
    .B(\i_game_and_vga.i_game_top.timer.counter[14] ),
    .C(net164),
    .Y(_0972_),
    .D(_0971_));
 sg13g2_nor2_1 _1715_ (.A(\i_game_and_vga.i_game_top.timer.counter[7] ),
    .B(net243),
    .Y(_0973_));
 sg13g2_nor4_2 _1716_ (.A(net255),
    .B(\i_game_and_vga.i_game_top.timer.counter[7] ),
    .C(net243),
    .Y(_0974_),
    .D(\i_game_and_vga.i_game_top.timer.counter[9] ));
 sg13g2_nor2_1 _1717_ (.A(\i_game_and_vga.i_game_top.timer.counter[16] ),
    .B(net248),
    .Y(_0975_));
 sg13g2_nor3_1 _1718_ (.A(\i_game_and_vga.i_game_top.timer.counter[16] ),
    .B(\i_game_and_vga.i_game_top.timer.counter[17] ),
    .C(\i_game_and_vga.i_game_top.timer.counter[20] ),
    .Y(_0976_));
 sg13g2_nor4_1 _1719_ (.A(\i_game_and_vga.i_game_top.timer.counter[10] ),
    .B(\i_game_and_vga.i_game_top.timer.counter[18] ),
    .C(\i_game_and_vga.i_game_top.timer.counter[19] ),
    .D(net152),
    .Y(_0977_));
 sg13g2_nand4_1 _1720_ (.B(_0974_),
    .C(_0976_),
    .A(_0972_),
    .Y(_0978_),
    .D(_0977_));
 sg13g2_nor3_1 _1721_ (.A(net190),
    .B(net160),
    .C(_0978_),
    .Y(_0979_));
 sg13g2_nor2b_1 _1722_ (.A(net149),
    .B_N(\i_game_and_vga.i_game_top.timer.counter[5] ),
    .Y(_0980_));
 sg13g2_nand4_1 _1723_ (.B(\i_game_and_vga.i_game_top.timer.counter[1] ),
    .C(net361),
    .A(_0536_),
    .Y(_0981_),
    .D(_0980_));
 sg13g2_nor4_1 _1724_ (.A(\i_game_and_vga.i_game_top.timer.counter[0] ),
    .B(net263),
    .C(net175),
    .D(_0981_),
    .Y(_0982_));
 sg13g2_a22oi_1 _1725_ (.Y(_0009_),
    .B1(_0979_),
    .B2(_0982_),
    .A2(_0537_),
    .A1(_0536_));
 sg13g2_xnor2_1 _1726_ (.Y(_0061_),
    .A(net120),
    .B(_0625_));
 sg13g2_xor2_1 _1727_ (.B(_0626_),
    .A(net234),
    .X(_0062_));
 sg13g2_xnor2_1 _1728_ (.Y(_0063_),
    .A(net133),
    .B(_0627_));
 sg13g2_xnor2_1 _1729_ (.Y(_0064_),
    .A(net145),
    .B(_0646_));
 sg13g2_xor2_1 _1730_ (.B(_0647_),
    .A(net196),
    .X(_0065_));
 sg13g2_a21o_1 _1731_ (.A2(_0647_),
    .A1(net196),
    .B1(net388),
    .X(_0203_));
 sg13g2_and2_1 _1732_ (.A(_0648_),
    .B(_0203_),
    .X(_0066_));
 sg13g2_xnor2_1 _1733_ (.Y(_0052_),
    .A(net162),
    .B(_0648_));
 sg13g2_xor2_1 _1734_ (.B(_0649_),
    .A(net183),
    .X(_0053_));
 sg13g2_a21o_1 _1735_ (.A2(_0649_),
    .A1(net183),
    .B1(net370),
    .X(_0204_));
 sg13g2_and2_1 _1736_ (.A(_0650_),
    .B(_0204_),
    .X(_0054_));
 sg13g2_xnor2_1 _1737_ (.Y(_0055_),
    .A(net141),
    .B(_0650_));
 sg13g2_xor2_1 _1738_ (.B(_0651_),
    .A(net179),
    .X(_0056_));
 sg13g2_a21o_1 _1739_ (.A2(_0651_),
    .A1(net179),
    .B1(net143),
    .X(_0205_));
 sg13g2_and2_1 _1740_ (.A(net144),
    .B(_0205_),
    .X(_0057_));
 sg13g2_xnor2_1 _1741_ (.Y(_0058_),
    .A(net118),
    .B(_0652_));
 sg13g2_xor2_1 _1742_ (.B(_0653_),
    .A(net109),
    .X(_0059_));
 sg13g2_a21oi_1 _1743_ (.A1(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.strobe_generator.counter[17] ),
    .A2(_0653_),
    .Y(_0206_),
    .B1(net99));
 sg13g2_nor2_1 _1744_ (.A(_0006_),
    .B(net100),
    .Y(_0060_));
 sg13g2_xnor2_1 _1745_ (.Y(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_display.y_sprite_plus_h_1[1] ),
    .A(net294),
    .B(net293));
 sg13g2_xnor2_1 _1746_ (.Y(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_display.x_sprite_plus_w_1[1] ),
    .A(net287),
    .B(net288));
 sg13g2_xnor2_1 _1747_ (.Y(\i_game_and_vga.i_game_top.sprite_target.sprite_display.y_sprite_plus_h_1[1] ),
    .A(net310),
    .B(net157));
 sg13g2_xnor2_1 _1748_ (.Y(\i_game_and_vga.i_game_top.sprite_target.sprite_display.x_sprite_plus_w_1[1] ),
    .A(net135),
    .B(\i_game_and_vga.i_game_top.sprite_target.sprite_control.sprite_x[1] ));
 sg13g2_xnor2_1 _1749_ (.Y(_0046_),
    .A(net126),
    .B(_0630_));
 sg13g2_xor2_1 _1750_ (.B(_0631_),
    .A(net220),
    .X(_0047_));
 sg13g2_xnor2_1 _1751_ (.Y(_0048_),
    .A(net128),
    .B(_0632_));
 sg13g2_xnor2_1 _1752_ (.Y(_0049_),
    .A(net131),
    .B(_0638_));
 sg13g2_xor2_1 _1753_ (.B(_0639_),
    .A(net206),
    .X(_0050_));
 sg13g2_a21o_1 _1754_ (.A2(_0639_),
    .A1(net206),
    .B1(net392),
    .X(_0207_));
 sg13g2_and2_1 _1755_ (.A(_0640_),
    .B(_0207_),
    .X(_0051_));
 sg13g2_xnor2_1 _1756_ (.Y(_0037_),
    .A(net114),
    .B(_0640_));
 sg13g2_xor2_1 _1757_ (.B(_0641_),
    .A(net170),
    .X(_0038_));
 sg13g2_a21o_1 _1758_ (.A2(_0641_),
    .A1(net170),
    .B1(net380),
    .X(_0208_));
 sg13g2_and2_1 _1759_ (.A(_0642_),
    .B(_0208_),
    .X(_0039_));
 sg13g2_xnor2_1 _1760_ (.Y(_0040_),
    .A(net122),
    .B(_0642_));
 sg13g2_xor2_1 _1761_ (.B(_0643_),
    .A(net158),
    .X(_0041_));
 sg13g2_a21o_1 _1762_ (.A2(_0643_),
    .A1(net158),
    .B1(net188),
    .X(_0209_));
 sg13g2_and2_1 _1763_ (.A(_0644_),
    .B(_0209_),
    .X(_0042_));
 sg13g2_xnor2_1 _1764_ (.Y(_0043_),
    .A(net124),
    .B(_0644_));
 sg13g2_xor2_1 _1765_ (.B(_0645_),
    .A(net111),
    .X(_0044_));
 sg13g2_a21oi_1 _1766_ (.A1(\i_game_and_vga.i_game_top.sprite_target.sprite_control.strobe_generator.counter[17] ),
    .A2(_0645_),
    .Y(_0210_),
    .B1(net103));
 sg13g2_nor2_1 _1767_ (.A(_0004_),
    .B(net104),
    .Y(_0045_));
 sg13g2_nand2_1 _1768_ (.Y(_0211_),
    .A(net304),
    .B(\i_game_and_vga.i_game_top.sprite_target.pixel_x[8] ));
 sg13g2_nor4_1 _1769_ (.A(\i_game_and_vga.i_game_top.sprite_target.pixel_x[7] ),
    .B(\i_game_and_vga.i_game_top.sprite_target.pixel_x[6] ),
    .C(\i_game_and_vga.i_game_top.sprite_target.pixel_x[5] ),
    .D(_0211_),
    .Y(_0212_));
 sg13g2_nand2_1 _1770_ (.Y(_0213_),
    .A(net393),
    .B(net309));
 sg13g2_nand2_1 _1771_ (.Y(_0214_),
    .A(\i_game_and_vga.i_game_top.sprite_target.pixel_x[1] ),
    .B(\i_game_and_vga.i_game_top.sprite_target.pixel_x[0] ));
 sg13g2_nor3_2 _1772_ (.A(_0552_),
    .B(_0553_),
    .C(_0214_),
    .Y(_0215_));
 sg13g2_and2_2 _1773_ (.A(\i_game_and_vga.i_game_top.sprite_target.pixel_x[4] ),
    .B(_0215_),
    .X(_0216_));
 sg13g2_and2_1 _1774_ (.A(_0212_),
    .B(_0216_),
    .X(_0217_));
 sg13g2_nand2_1 _1775_ (.Y(_0218_),
    .A(_0212_),
    .B(_0216_));
 sg13g2_nand2_2 _1776_ (.Y(_0219_),
    .A(net307),
    .B(_0217_));
 sg13g2_nor4_1 _1777_ (.A(\i_game_and_vga.i_game_top.sprite_target.pixel_y[6] ),
    .B(\i_game_and_vga.i_game_top.sprite_target.pixel_y[5] ),
    .C(\i_game_and_vga.i_game_top.sprite_target.pixel_y[4] ),
    .D(_0585_),
    .Y(_0220_));
 sg13g2_nor2_1 _1778_ (.A(net194),
    .B(\i_game_and_vga.i_game_top.sprite_target.pixel_y[0] ),
    .Y(_0221_));
 sg13g2_nor4_1 _1779_ (.A(\i_game_and_vga.i_game_top.sprite_target.pixel_y[8] ),
    .B(\i_game_and_vga.i_game_top.sprite_target.pixel_y[7] ),
    .C(net313),
    .D(\i_game_and_vga.i_game_top.sprite_target.pixel_y[0] ),
    .Y(_0222_));
 sg13g2_nand4_1 _1780_ (.B(\i_game_and_vga.i_game_top.sprite_target.pixel_y[2] ),
    .C(_0220_),
    .A(net312),
    .Y(_0223_),
    .D(_0222_));
 sg13g2_a21oi_1 _1781_ (.A1(_0567_),
    .A2(_0223_),
    .Y(_0224_),
    .B1(_0219_));
 sg13g2_a21oi_1 _1782_ (.A1(_0567_),
    .A2(_0219_),
    .Y(_0105_),
    .B1(_0224_));
 sg13g2_and2_1 _1783_ (.A(net313),
    .B(\i_game_and_vga.i_game_top.sprite_target.pixel_y[0] ),
    .X(_0225_));
 sg13g2_nor3_1 _1784_ (.A(net268),
    .B(_0221_),
    .C(_0225_),
    .Y(_0226_));
 sg13g2_a21oi_1 _1785_ (.A1(_0586_),
    .A2(net267),
    .Y(_0227_),
    .B1(_0226_));
 sg13g2_nor2_1 _1786_ (.A(net194),
    .B(net308),
    .Y(_0228_));
 sg13g2_a21oi_1 _1787_ (.A1(net308),
    .A2(_0227_),
    .Y(_0106_),
    .B1(_0228_));
 sg13g2_nand2_1 _1788_ (.Y(_0229_),
    .A(net376),
    .B(_0219_));
 sg13g2_and2_2 _1789_ (.A(_0217_),
    .B(_0223_),
    .X(_0230_));
 sg13g2_xnor2_1 _1790_ (.Y(_0231_),
    .A(_0566_),
    .B(_0225_));
 sg13g2_nand3_1 _1791_ (.B(_0230_),
    .C(_0231_),
    .A(net308),
    .Y(_0232_));
 sg13g2_nand2_1 _1792_ (.Y(_0107_),
    .A(_0229_),
    .B(_0232_));
 sg13g2_nand2_1 _1793_ (.Y(_0233_),
    .A(net312),
    .B(_0219_));
 sg13g2_nor2b_1 _1794_ (.A(_0030_),
    .B_N(_0225_),
    .Y(_0234_));
 sg13g2_xnor2_1 _1795_ (.Y(_0235_),
    .A(_0565_),
    .B(_0234_));
 sg13g2_nand2_1 _1796_ (.Y(_0236_),
    .A(_0230_),
    .B(_0235_));
 sg13g2_o21ai_1 _1797_ (.B1(_0233_),
    .Y(_0108_),
    .A1(_0623_),
    .A2(_0236_));
 sg13g2_nand3_1 _1798_ (.B(\i_game_and_vga.i_game_top.sprite_target.pixel_y[2] ),
    .C(_0225_),
    .A(net312),
    .Y(_0237_));
 sg13g2_nor2_1 _1799_ (.A(net267),
    .B(_0237_),
    .Y(_0238_));
 sg13g2_xnor2_1 _1800_ (.Y(_0239_),
    .A(_0562_),
    .B(_0238_));
 sg13g2_nor2_1 _1801_ (.A(_0623_),
    .B(_0239_),
    .Y(_0240_));
 sg13g2_a21oi_1 _1802_ (.A1(_0562_),
    .A2(_0623_),
    .Y(_0109_),
    .B1(_0240_));
 sg13g2_nand2_1 _1803_ (.Y(_0241_),
    .A(net359),
    .B(_0219_));
 sg13g2_or2_1 _1804_ (.X(_0242_),
    .B(_0237_),
    .A(_0562_));
 sg13g2_xor2_1 _1805_ (.B(_0242_),
    .A(_0028_),
    .X(_0243_));
 sg13g2_nand3_1 _1806_ (.B(_0230_),
    .C(_0243_),
    .A(net308),
    .Y(_0244_));
 sg13g2_nand2_1 _1807_ (.Y(_0110_),
    .A(_0241_),
    .B(_0244_));
 sg13g2_or2_1 _1808_ (.X(_0245_),
    .B(_0223_),
    .A(net267));
 sg13g2_or2_1 _1809_ (.X(_0246_),
    .B(_0242_),
    .A(_0561_));
 sg13g2_nor2_1 _1810_ (.A(net267),
    .B(_0246_),
    .Y(_0247_));
 sg13g2_xnor2_1 _1811_ (.Y(_0248_),
    .A(_0027_),
    .B(_0247_));
 sg13g2_nor2_1 _1812_ (.A(_0027_),
    .B(_0246_),
    .Y(_0249_));
 sg13g2_nand2_1 _1813_ (.Y(_0250_),
    .A(_0245_),
    .B(_0248_));
 sg13g2_nor2_1 _1814_ (.A(net398),
    .B(net307),
    .Y(_0251_));
 sg13g2_a21oi_1 _1815_ (.A1(net307),
    .A2(_0250_),
    .Y(_0111_),
    .B1(_0251_));
 sg13g2_nand2_1 _1816_ (.Y(_0252_),
    .A(net311),
    .B(_0219_));
 sg13g2_xnor2_1 _1817_ (.Y(_0253_),
    .A(_0035_),
    .B(_0249_));
 sg13g2_nand3_1 _1818_ (.B(_0230_),
    .C(_0253_),
    .A(net307),
    .Y(_0254_));
 sg13g2_nand2_1 _1819_ (.Y(_0112_),
    .A(_0252_),
    .B(_0254_));
 sg13g2_nor2_1 _1820_ (.A(net384),
    .B(net307),
    .Y(_0255_));
 sg13g2_nand3_1 _1821_ (.B(\i_game_and_vga.i_game_top.sprite_target.pixel_y[6] ),
    .C(_0247_),
    .A(net311),
    .Y(_0256_));
 sg13g2_xnor2_1 _1822_ (.Y(_0257_),
    .A(_0555_),
    .B(_0256_));
 sg13g2_a21oi_1 _1823_ (.A1(net307),
    .A2(_0257_),
    .Y(_0113_),
    .B1(_0255_));
 sg13g2_nand4_1 _1824_ (.B(\i_game_and_vga.i_game_top.sprite_target.pixel_y[6] ),
    .C(_0578_),
    .A(net311),
    .Y(_0258_),
    .D(_0247_));
 sg13g2_o21ai_1 _1825_ (.B1(_0245_),
    .Y(_0259_),
    .A1(_0585_),
    .A2(_0258_));
 sg13g2_a21o_1 _1826_ (.A2(_0258_),
    .A1(_0585_),
    .B1(_0259_),
    .X(_0260_));
 sg13g2_nor2_1 _1827_ (.A(net189),
    .B(net308),
    .Y(_0261_));
 sg13g2_a21oi_1 _1828_ (.A1(net308),
    .A2(_0260_),
    .Y(_0114_),
    .B1(_0261_));
 sg13g2_mux2_1 _1829_ (.A0(net157),
    .A1(net223),
    .S(net130),
    .X(_0115_));
 sg13g2_nor2_1 _1830_ (.A(net279),
    .B(net83),
    .Y(_0262_));
 sg13g2_a21oi_1 _1831_ (.A1(_0088_),
    .A2(net279),
    .Y(_0116_),
    .B1(net84));
 sg13g2_mux2_1 _1832_ (.A0(net80),
    .A1(net71),
    .S(net279),
    .X(_0117_));
 sg13g2_nor2_1 _1833_ (.A(net279),
    .B(net68),
    .Y(_0263_));
 sg13g2_a21oi_1 _1834_ (.A1(_0090_),
    .A2(net279),
    .Y(_0118_),
    .B1(net69));
 sg13g2_nor2_1 _1835_ (.A(net279),
    .B(net78),
    .Y(_0264_));
 sg13g2_a21oi_1 _1836_ (.A1(net182),
    .A2(net279),
    .Y(_0119_),
    .B1(_0264_));
 sg13g2_o21ai_1 _1837_ (.B1(net278),
    .Y(_0265_),
    .A1(net73),
    .A2(net182));
 sg13g2_a21oi_1 _1838_ (.A1(net73),
    .A2(net182),
    .Y(_0266_),
    .B1(_0265_));
 sg13g2_a21oi_1 _1839_ (.A1(_0539_),
    .A2(_0575_),
    .Y(_0120_),
    .B1(_0266_));
 sg13g2_o21ai_1 _1840_ (.B1(_0265_),
    .Y(_0121_),
    .A1(net278),
    .A2(_0574_));
 sg13g2_a22oi_1 _1841_ (.Y(_0267_),
    .B1(_0230_),
    .B2(_0253_),
    .A2(net267),
    .A1(net311));
 sg13g2_a22oi_1 _1842_ (.Y(_0268_),
    .B1(_0230_),
    .B2(_0243_),
    .A2(net267),
    .A1(\i_game_and_vga.i_game_top.sprite_target.pixel_y[5] ));
 sg13g2_or4_1 _1843_ (.A(_0250_),
    .B(_0257_),
    .C(_0267_),
    .D(_0268_),
    .X(_0269_));
 sg13g2_nand2_1 _1844_ (.Y(_0270_),
    .A(\i_game_and_vga.i_game_top.sprite_target.pixel_x[5] ),
    .B(_0216_));
 sg13g2_nand4_1 _1845_ (.B(\i_game_and_vga.i_game_top.sprite_target.pixel_x[6] ),
    .C(\i_game_and_vga.i_game_top.sprite_target.pixel_x[5] ),
    .A(\i_game_and_vga.i_game_top.sprite_target.pixel_x[7] ),
    .Y(_0271_),
    .D(_0216_));
 sg13g2_inv_1 _1846_ (.Y(_0272_),
    .A(_0271_));
 sg13g2_a21oi_1 _1847_ (.A1(\i_game_and_vga.i_game_top.sprite_target.pixel_x[8] ),
    .A2(_0272_),
    .Y(_0273_),
    .B1(net304));
 sg13g2_o21ai_1 _1848_ (.B1(net268),
    .Y(_0274_),
    .A1(_0211_),
    .A2(_0271_));
 sg13g2_nor2_1 _1849_ (.A(_0273_),
    .B(_0274_),
    .Y(_0275_));
 sg13g2_o21ai_1 _1850_ (.B1(net268),
    .Y(_0276_),
    .A1(_0019_),
    .A2(_0271_));
 sg13g2_a21oi_1 _1851_ (.A1(_0019_),
    .A2(_0271_),
    .Y(_0277_),
    .B1(_0276_));
 sg13g2_nor2_1 _1852_ (.A(_0021_),
    .B(_0270_),
    .Y(_0278_));
 sg13g2_xnor2_1 _1853_ (.Y(_0279_),
    .A(\i_game_and_vga.i_game_top.sprite_target.pixel_x[7] ),
    .B(_0278_));
 sg13g2_inv_1 _1854_ (.Y(_0280_),
    .A(_0279_));
 sg13g2_o21ai_1 _1855_ (.B1(_0275_),
    .Y(_0281_),
    .A1(_0277_),
    .A2(_0280_));
 sg13g2_nand4_1 _1856_ (.B(_0260_),
    .C(_0269_),
    .A(net308),
    .Y(_0282_),
    .D(_0281_));
 sg13g2_o21ai_1 _1857_ (.B1(_0282_),
    .Y(_0122_),
    .A1(_0619_),
    .A2(net309));
 sg13g2_xnor2_1 _1858_ (.Y(_0283_),
    .A(_0022_),
    .B(_0216_));
 sg13g2_nand2_1 _1859_ (.Y(_0284_),
    .A(net268),
    .B(_0283_));
 sg13g2_xnor2_1 _1860_ (.Y(_0285_),
    .A(_0547_),
    .B(_0270_));
 sg13g2_xnor2_1 _1861_ (.Y(_0286_),
    .A(\i_game_and_vga.i_game_top.sprite_target.pixel_x[4] ),
    .B(_0215_));
 sg13g2_and3_1 _1862_ (.X(_0287_),
    .A(_0284_),
    .B(_0285_),
    .C(_0286_));
 sg13g2_nor4_1 _1863_ (.A(_0545_),
    .B(_0547_),
    .C(_0284_),
    .D(_0286_),
    .Y(_0288_));
 sg13g2_nor4_1 _1864_ (.A(_0277_),
    .B(_0279_),
    .C(_0287_),
    .D(_0288_),
    .Y(_0289_));
 sg13g2_nand3_1 _1865_ (.B(_0275_),
    .C(_0289_),
    .A(net306),
    .Y(_0290_));
 sg13g2_o21ai_1 _1866_ (.B1(_0290_),
    .Y(_0291_),
    .A1(net309),
    .A2(net229));
 sg13g2_inv_1 _1867_ (.Y(_0123_),
    .A(net230));
 sg13g2_a21oi_1 _1868_ (.A1(\i_game_and_vga.i_game_top.sprite_target.pixel_y[2] ),
    .A2(net267),
    .Y(_0292_),
    .B1(_0227_));
 sg13g2_nand2_1 _1869_ (.Y(_0293_),
    .A(net312),
    .B(net267));
 sg13g2_a22oi_1 _1870_ (.Y(_0294_),
    .B1(_0236_),
    .B2(_0293_),
    .A2(_0231_),
    .A1(_0230_));
 sg13g2_nand3_1 _1871_ (.B(_0292_),
    .C(_0294_),
    .A(_0240_),
    .Y(_0295_));
 sg13g2_nor2_1 _1872_ (.A(_0269_),
    .B(_0295_),
    .Y(_0296_));
 sg13g2_a22oi_1 _1873_ (.Y(_0124_),
    .B1(_0260_),
    .B2(_0296_),
    .A2(_0624_),
    .A1(_0623_));
 sg13g2_xor2_1 _1874_ (.B(net309),
    .A(net393),
    .X(_0125_));
 sg13g2_xnor2_1 _1875_ (.Y(_0126_),
    .A(net397),
    .B(_0213_));
 sg13g2_xor2_1 _1876_ (.B(_0214_),
    .A(net407),
    .X(_0297_));
 sg13g2_nand3_1 _1877_ (.B(net268),
    .C(_0297_),
    .A(net305),
    .Y(_0298_));
 sg13g2_o21ai_1 _1878_ (.B1(_0298_),
    .Y(_0127_),
    .A1(_0553_),
    .A2(net306));
 sg13g2_nand4_1 _1879_ (.B(\i_game_and_vga.i_game_top.sprite_target.pixel_x[1] ),
    .C(\i_game_and_vga.i_game_top.sprite_target.pixel_x[0] ),
    .A(net373),
    .Y(_0299_),
    .D(net305));
 sg13g2_a22oi_1 _1880_ (.Y(_0128_),
    .B1(net374),
    .B2(_0552_),
    .A2(_0215_),
    .A1(net305));
 sg13g2_a21oi_1 _1881_ (.A1(net305),
    .A2(_0215_),
    .Y(_0300_),
    .B1(net367));
 sg13g2_a21oi_1 _1882_ (.A1(net305),
    .A2(_0216_),
    .Y(_0129_),
    .B1(_0300_));
 sg13g2_nor2_1 _1883_ (.A(net385),
    .B(net305),
    .Y(_0301_));
 sg13g2_a21oi_1 _1884_ (.A1(net305),
    .A2(_0284_),
    .Y(_0130_),
    .B1(_0301_));
 sg13g2_nor2_1 _1885_ (.A(net383),
    .B(net306),
    .Y(_0302_));
 sg13g2_a21oi_1 _1886_ (.A1(net305),
    .A2(_0285_),
    .Y(_0131_),
    .B1(_0302_));
 sg13g2_nor2_1 _1887_ (.A(net404),
    .B(net306),
    .Y(_0303_));
 sg13g2_a21oi_1 _1888_ (.A1(net307),
    .A2(_0279_),
    .Y(_0132_),
    .B1(_0303_));
 sg13g2_nand2_1 _1889_ (.Y(_0304_),
    .A(net306),
    .B(_0277_));
 sg13g2_o21ai_1 _1890_ (.B1(_0304_),
    .Y(_0133_),
    .A1(_0543_),
    .A2(net306));
 sg13g2_mux2_1 _1891_ (.A0(net304),
    .A1(_0275_),
    .S(net306),
    .X(_0134_));
 sg13g2_a21oi_2 _1892_ (.B1(net277),
    .Y(_0305_),
    .A2(\i_game_and_vga.i_game_top.master_fsm.sprite_target_enable_update ),
    .A1(\i_game_and_vga.i_game_top.sprite_target.sprite_control.strobe_generator.strobe ));
 sg13g2_inv_1 _1893_ (.Y(_0306_),
    .A(net276));
 sg13g2_nand2_2 _1894_ (.Y(_0307_),
    .A(net303),
    .B(net90));
 sg13g2_a21oi_1 _1895_ (.A1(net238),
    .A2(_0307_),
    .Y(_0308_),
    .B1(net276));
 sg13g2_a21oi_1 _1896_ (.A1(net90),
    .A2(_0306_),
    .Y(_0309_),
    .B1(net303));
 sg13g2_nor2_1 _1897_ (.A(_0308_),
    .B(_0309_),
    .Y(_0135_));
 sg13g2_nor2_1 _1898_ (.A(net302),
    .B(net297),
    .Y(_0310_));
 sg13g2_nand2_1 _1899_ (.Y(_0311_),
    .A(net302),
    .B(net297));
 sg13g2_nor2b_1 _1900_ (.A(_0310_),
    .B_N(_0311_),
    .Y(_0312_));
 sg13g2_nor2b_2 _1901_ (.A(net276),
    .B_N(_0015_),
    .Y(_0313_));
 sg13g2_inv_1 _1902_ (.Y(_0314_),
    .A(_0313_));
 sg13g2_xnor2_1 _1903_ (.Y(_0315_),
    .A(_0307_),
    .B(_0312_));
 sg13g2_a22oi_1 _1904_ (.Y(_0316_),
    .B1(_0313_),
    .B2(_0315_),
    .A2(net276),
    .A1(net302));
 sg13g2_inv_1 _1905_ (.Y(_0136_),
    .A(_0316_));
 sg13g2_and2_1 _1906_ (.A(\i_game_and_vga.i_game_top.sprite_target.sprite_control.sprite_x[2] ),
    .B(net297),
    .X(_0317_));
 sg13g2_xor2_1 _1907_ (.B(net297),
    .A(\i_game_and_vga.i_game_top.sprite_target.sprite_control.sprite_x[2] ),
    .X(_0318_));
 sg13g2_o21ai_1 _1908_ (.B1(_0311_),
    .Y(_0319_),
    .A1(_0307_),
    .A2(_0310_));
 sg13g2_o21ai_1 _1909_ (.B1(_0313_),
    .Y(_0320_),
    .A1(_0318_),
    .A2(_0319_));
 sg13g2_a21oi_1 _1910_ (.A1(_0318_),
    .A2(_0319_),
    .Y(_0321_),
    .B1(_0320_));
 sg13g2_a21o_1 _1911_ (.A2(net275),
    .A1(net89),
    .B1(_0321_),
    .X(_0137_));
 sg13g2_a21oi_1 _1912_ (.A1(_0318_),
    .A2(_0319_),
    .Y(_0322_),
    .B1(_0317_));
 sg13g2_nor2_1 _1913_ (.A(net301),
    .B(net296),
    .Y(_0323_));
 sg13g2_xnor2_1 _1914_ (.Y(_0324_),
    .A(net301),
    .B(net296));
 sg13g2_nand3_1 _1915_ (.B(net377),
    .C(net387),
    .A(_0539_),
    .Y(_0325_));
 sg13g2_xnor2_1 _1916_ (.Y(_0326_),
    .A(_0322_),
    .B(_0324_));
 sg13g2_nor2_2 _1917_ (.A(net67),
    .B(_0539_),
    .Y(_0327_));
 sg13g2_a21oi_1 _1918_ (.A1(net301),
    .A2(net275),
    .Y(_0328_),
    .B1(_0327_));
 sg13g2_o21ai_1 _1919_ (.B1(_0328_),
    .Y(_0138_),
    .A1(net378),
    .A2(_0326_));
 sg13g2_xnor2_1 _1920_ (.Y(_0329_),
    .A(net300),
    .B(net296));
 sg13g2_a221oi_1 _1921_ (.B2(_0319_),
    .C1(_0317_),
    .B1(_0318_),
    .A1(net301),
    .Y(_0330_),
    .A2(net296));
 sg13g2_or3_1 _1922_ (.A(_0323_),
    .B(_0329_),
    .C(_0330_),
    .X(_0331_));
 sg13g2_o21ai_1 _1923_ (.B1(_0329_),
    .Y(_0332_),
    .A1(_0323_),
    .A2(_0330_));
 sg13g2_nand2_1 _1924_ (.Y(_0333_),
    .A(_0331_),
    .B(_0332_));
 sg13g2_a21oi_1 _1925_ (.A1(net300),
    .A2(net275),
    .Y(_0334_),
    .B1(_0327_));
 sg13g2_o21ai_1 _1926_ (.B1(_0334_),
    .Y(_0139_),
    .A1(_0325_),
    .A2(_0333_));
 sg13g2_xor2_1 _1927_ (.B(net296),
    .A(\i_game_and_vga.i_game_top.sprite_target.sprite_control.sprite_x[5] ),
    .X(_0335_));
 sg13g2_o21ai_1 _1928_ (.B1(_0331_),
    .Y(_0336_),
    .A1(_0572_),
    .A2(_0618_));
 sg13g2_xnor2_1 _1929_ (.Y(_0337_),
    .A(_0335_),
    .B(_0336_));
 sg13g2_a21oi_1 _1930_ (.A1(net222),
    .A2(net275),
    .Y(_0338_),
    .B1(_0327_));
 sg13g2_o21ai_1 _1931_ (.B1(_0338_),
    .Y(_0140_),
    .A1(net378),
    .A2(_0337_));
 sg13g2_xnor2_1 _1932_ (.Y(_0339_),
    .A(\i_game_and_vga.i_game_top.sprite_target.sprite_control.sprite_x[6] ),
    .B(net295));
 sg13g2_nand2b_1 _1933_ (.Y(_0340_),
    .B(_0335_),
    .A_N(_0331_));
 sg13g2_o21ai_1 _1934_ (.B1(net295),
    .Y(_0341_),
    .A1(\i_game_and_vga.i_game_top.sprite_target.sprite_control.sprite_x[5] ),
    .A2(net300));
 sg13g2_and3_1 _1935_ (.X(_0342_),
    .A(_0339_),
    .B(_0340_),
    .C(_0341_));
 sg13g2_a21oi_1 _1936_ (.A1(_0340_),
    .A2(_0341_),
    .Y(_0343_),
    .B1(_0339_));
 sg13g2_or2_1 _1937_ (.X(_0344_),
    .B(_0343_),
    .A(_0325_));
 sg13g2_a21oi_1 _1938_ (.A1(net97),
    .A2(net275),
    .Y(_0345_),
    .B1(_0327_));
 sg13g2_o21ai_1 _1939_ (.B1(_0345_),
    .Y(_0141_),
    .A1(_0342_),
    .A2(_0344_));
 sg13g2_xor2_1 _1940_ (.B(net295),
    .A(\i_game_and_vga.i_game_top.sprite_target.sprite_control.sprite_x[7] ),
    .X(_0346_));
 sg13g2_a21oi_1 _1941_ (.A1(\i_game_and_vga.i_game_top.sprite_target.sprite_control.sprite_x[6] ),
    .A2(net295),
    .Y(_0347_),
    .B1(_0343_));
 sg13g2_xnor2_1 _1942_ (.Y(_0348_),
    .A(_0346_),
    .B(_0347_));
 sg13g2_a22oi_1 _1943_ (.Y(_0349_),
    .B1(_0313_),
    .B2(_0348_),
    .A2(net275),
    .A1(net192));
 sg13g2_inv_1 _1944_ (.Y(_0142_),
    .A(_0349_));
 sg13g2_nand2_1 _1945_ (.Y(_0350_),
    .A(net299),
    .B(net275));
 sg13g2_nor2_1 _1946_ (.A(_0339_),
    .B(_0340_),
    .Y(_0351_));
 sg13g2_o21ai_1 _1947_ (.B1(net295),
    .Y(_0352_),
    .A1(\i_game_and_vga.i_game_top.sprite_target.sprite_control.sprite_x[7] ),
    .A2(\i_game_and_vga.i_game_top.sprite_target.sprite_control.sprite_x[6] ));
 sg13g2_nand2_1 _1948_ (.Y(_0353_),
    .A(_0341_),
    .B(_0352_));
 sg13g2_a21oi_1 _1949_ (.A1(_0346_),
    .A2(_0351_),
    .Y(_0354_),
    .B1(_0353_));
 sg13g2_nand2_1 _1950_ (.Y(_0355_),
    .A(net299),
    .B(net295));
 sg13g2_xnor2_1 _1951_ (.Y(_0356_),
    .A(net299),
    .B(net295));
 sg13g2_xnor2_1 _1952_ (.Y(_0357_),
    .A(_0354_),
    .B(_0356_));
 sg13g2_o21ai_1 _1953_ (.B1(_0350_),
    .Y(_0143_),
    .A1(_0314_),
    .A2(_0357_));
 sg13g2_o21ai_1 _1954_ (.B1(_0355_),
    .Y(_0358_),
    .A1(_0354_),
    .A2(_0356_));
 sg13g2_xor2_1 _1955_ (.B(net295),
    .A(net298),
    .X(_0359_));
 sg13g2_xnor2_1 _1956_ (.Y(_0360_),
    .A(_0358_),
    .B(_0359_));
 sg13g2_a21oi_1 _1957_ (.A1(net298),
    .A2(net275),
    .Y(_0361_),
    .B1(_0327_));
 sg13g2_o21ai_1 _1958_ (.B1(_0361_),
    .Y(_0144_),
    .A1(net378),
    .A2(_0360_));
 sg13g2_o21ai_1 _1959_ (.B1(\i_game_and_vga.i_game_top.master_fsm.state[1] ),
    .Y(_0362_),
    .A1(\i_game_and_vga.i_game_top.collision ),
    .A2(\i_game_and_vga.i_game_top.game_won ));
 sg13g2_o21ai_1 _1960_ (.B1(_0362_),
    .Y(_0145_),
    .A1(net76),
    .A2(_0621_));
 sg13g2_a22oi_1 _1961_ (.Y(_0146_),
    .B1(_0327_),
    .B2(_0093_),
    .A2(_0617_),
    .A1(_0539_));
 sg13g2_a21o_1 _1962_ (.A2(net297),
    .A1(_0539_),
    .B1(_0327_),
    .X(_0147_));
 sg13g2_nand2_1 _1963_ (.Y(_0363_),
    .A(net107),
    .B(\i_game_and_vga.i_game_top.master_fsm.sprite_torpedo_enable_update ));
 sg13g2_a21oi_1 _1964_ (.A1(net107),
    .A2(\i_game_and_vga.i_game_top.master_fsm.sprite_torpedo_enable_update ),
    .Y(_0364_),
    .B1(net278));
 sg13g2_inv_2 _1965_ (.Y(_0365_),
    .A(net272));
 sg13g2_nand2_2 _1966_ (.Y(_0366_),
    .A(net294),
    .B(net259));
 sg13g2_a21oi_1 _1967_ (.A1(_0015_),
    .A2(_0366_),
    .Y(_0367_),
    .B1(net274));
 sg13g2_a21oi_1 _1968_ (.A1(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.dy[0] ),
    .A2(_0365_),
    .Y(_0368_),
    .B1(net94));
 sg13g2_nor2_1 _1969_ (.A(_0367_),
    .B(net95),
    .Y(_0148_));
 sg13g2_nand2_1 _1970_ (.Y(_0369_),
    .A(net292),
    .B(net273));
 sg13g2_nand2_1 _1971_ (.Y(_0370_),
    .A(net292),
    .B(net283));
 sg13g2_xnor2_1 _1972_ (.Y(_0371_),
    .A(net292),
    .B(net283));
 sg13g2_nand2_2 _1973_ (.Y(_0372_),
    .A(_0015_),
    .B(_0365_));
 sg13g2_xnor2_1 _1974_ (.Y(_0373_),
    .A(_0366_),
    .B(_0371_));
 sg13g2_o21ai_1 _1975_ (.B1(_0369_),
    .Y(_0149_),
    .A1(_0372_),
    .A2(_0373_));
 sg13g2_and2_1 _1976_ (.A(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.sprite_y[2] ),
    .B(net283),
    .X(_0374_));
 sg13g2_xor2_1 _1977_ (.B(net283),
    .A(net291),
    .X(_0375_));
 sg13g2_o21ai_1 _1978_ (.B1(_0370_),
    .Y(_0376_),
    .A1(_0366_),
    .A2(_0371_));
 sg13g2_and2_1 _1979_ (.A(_0375_),
    .B(_0376_),
    .X(_0377_));
 sg13g2_nor2_1 _1980_ (.A(_0375_),
    .B(_0376_),
    .Y(_0378_));
 sg13g2_nor3_1 _1981_ (.A(_0372_),
    .B(_0377_),
    .C(_0378_),
    .Y(_0379_));
 sg13g2_a21o_1 _1982_ (.A2(net273),
    .A1(net291),
    .B1(_0379_),
    .X(_0150_));
 sg13g2_nor2_1 _1983_ (.A(_0374_),
    .B(_0377_),
    .Y(_0380_));
 sg13g2_nor2_2 _1984_ (.A(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.sprite_y[3] ),
    .B(net283),
    .Y(_0381_));
 sg13g2_and2_1 _1985_ (.A(net290),
    .B(net283),
    .X(_0382_));
 sg13g2_nor3_1 _1986_ (.A(_0380_),
    .B(_0381_),
    .C(_0382_),
    .Y(_0383_));
 sg13g2_o21ai_1 _1987_ (.B1(_0380_),
    .Y(_0384_),
    .A1(_0381_),
    .A2(_0382_));
 sg13g2_nor2_1 _1988_ (.A(_0372_),
    .B(_0383_),
    .Y(_0385_));
 sg13g2_a22oi_1 _1989_ (.Y(_0386_),
    .B1(_0384_),
    .B2(_0385_),
    .A2(net273),
    .A1(net290));
 sg13g2_inv_1 _1990_ (.Y(_0151_),
    .A(_0386_));
 sg13g2_nor2_2 _1991_ (.A(net277),
    .B(_0363_),
    .Y(_0387_));
 sg13g2_nand2b_2 _1992_ (.Y(_0388_),
    .B(_0539_),
    .A_N(_0363_));
 sg13g2_xnor2_1 _1993_ (.Y(_0389_),
    .A(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.sprite_y[4] ),
    .B(net283));
 sg13g2_a221oi_1 _1994_ (.B2(_0376_),
    .C1(_0374_),
    .B1(_0375_),
    .A1(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.sprite_y[3] ),
    .Y(_0390_),
    .A2(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.dy[1] ));
 sg13g2_nor2_1 _1995_ (.A(_0381_),
    .B(_0390_),
    .Y(_0391_));
 sg13g2_nor3_2 _1996_ (.A(_0381_),
    .B(_0389_),
    .C(_0390_),
    .Y(_0392_));
 sg13g2_xor2_1 _1997_ (.B(_0391_),
    .A(_0389_),
    .X(_0393_));
 sg13g2_a22oi_1 _1998_ (.Y(_0152_),
    .B1(_0387_),
    .B2(_0393_),
    .A2(net274),
    .A1(_0563_));
 sg13g2_xor2_1 _1999_ (.B(net284),
    .A(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.sprite_y[5] ),
    .X(_0394_));
 sg13g2_a21oi_1 _2000_ (.A1(net289),
    .A2(net284),
    .Y(_0395_),
    .B1(_0392_));
 sg13g2_xor2_1 _2001_ (.B(_0395_),
    .A(_0394_),
    .X(_0396_));
 sg13g2_nand2_1 _2002_ (.Y(_0397_),
    .A(net102),
    .B(net274));
 sg13g2_o21ai_1 _2003_ (.B1(_0397_),
    .Y(_0153_),
    .A1(_0372_),
    .A2(_0396_));
 sg13g2_xnor2_1 _2004_ (.Y(_0398_),
    .A(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.sprite_y[6] ),
    .B(net284));
 sg13g2_nand2_2 _2005_ (.Y(_0399_),
    .A(_0392_),
    .B(_0394_));
 sg13g2_o21ai_1 _2006_ (.B1(net284),
    .Y(_0400_),
    .A1(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.sprite_y[5] ),
    .A2(net289));
 sg13g2_a21oi_1 _2007_ (.A1(_0399_),
    .A2(_0400_),
    .Y(_0401_),
    .B1(_0398_));
 sg13g2_nand3_1 _2008_ (.B(_0399_),
    .C(_0400_),
    .A(_0398_),
    .Y(_0402_));
 sg13g2_nand2b_1 _2009_ (.Y(_0403_),
    .B(_0402_),
    .A_N(_0401_));
 sg13g2_a22oi_1 _2010_ (.Y(_0154_),
    .B1(_0387_),
    .B2(_0403_),
    .A2(net272),
    .A1(_0558_));
 sg13g2_xor2_1 _2011_ (.B(net284),
    .A(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.sprite_y[7] ),
    .X(_0404_));
 sg13g2_a21oi_1 _2012_ (.A1(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.sprite_y[6] ),
    .A2(net284),
    .Y(_0405_),
    .B1(_0401_));
 sg13g2_o21ai_1 _2013_ (.B1(_0387_),
    .Y(_0406_),
    .A1(_0404_),
    .A2(_0405_));
 sg13g2_a21oi_1 _2014_ (.A1(_0404_),
    .A2(_0405_),
    .Y(_0407_),
    .B1(_0406_));
 sg13g2_a21oi_1 _2015_ (.A1(_0556_),
    .A2(net272),
    .Y(_0155_),
    .B1(_0407_));
 sg13g2_nand2b_1 _2016_ (.Y(_0408_),
    .B(_0404_),
    .A_N(_0398_));
 sg13g2_o21ai_1 _2017_ (.B1(net284),
    .Y(_0409_),
    .A1(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.sprite_y[7] ),
    .A2(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.sprite_y[6] ));
 sg13g2_and2_1 _2018_ (.A(_0400_),
    .B(_0409_),
    .X(_0410_));
 sg13g2_o21ai_1 _2019_ (.B1(_0410_),
    .Y(_0411_),
    .A1(_0399_),
    .A2(_0408_));
 sg13g2_xor2_1 _2020_ (.B(net284),
    .A(net82),
    .X(_0412_));
 sg13g2_xnor2_1 _2021_ (.Y(_0413_),
    .A(_0411_),
    .B(_0412_));
 sg13g2_a22oi_1 _2022_ (.Y(_0156_),
    .B1(_0387_),
    .B2(_0413_),
    .A2(net272),
    .A1(_0554_));
 sg13g2_nand2_1 _2023_ (.Y(_0414_),
    .A(net288),
    .B(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.dx[0] ));
 sg13g2_xnor2_1 _2024_ (.Y(_0415_),
    .A(net288),
    .B(net167));
 sg13g2_a22oi_1 _2025_ (.Y(_0416_),
    .B1(net288),
    .B2(net273),
    .A2(net277),
    .A1(net61));
 sg13g2_o21ai_1 _2026_ (.B1(_0416_),
    .Y(_0157_),
    .A1(_0388_),
    .A2(net168));
 sg13g2_nand2_1 _2027_ (.Y(_0417_),
    .A(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.sprite_x[1] ),
    .B(net282));
 sg13g2_xnor2_1 _2028_ (.Y(_0418_),
    .A(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.sprite_x[1] ),
    .B(net282));
 sg13g2_xnor2_1 _2029_ (.Y(_0419_),
    .A(_0414_),
    .B(_0418_));
 sg13g2_a22oi_1 _2030_ (.Y(_0420_),
    .B1(net273),
    .B2(net287),
    .A2(net64),
    .A1(net277));
 sg13g2_o21ai_1 _2031_ (.B1(_0420_),
    .Y(_0158_),
    .A1(_0388_),
    .A2(_0419_));
 sg13g2_and2_1 _2032_ (.A(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.sprite_x[2] ),
    .B(net280),
    .X(_0421_));
 sg13g2_or2_1 _2033_ (.X(_0422_),
    .B(net280),
    .A(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.sprite_x[2] ));
 sg13g2_nor2b_1 _2034_ (.A(_0421_),
    .B_N(_0422_),
    .Y(_0423_));
 sg13g2_o21ai_1 _2035_ (.B1(_0417_),
    .Y(_0424_),
    .A1(_0414_),
    .A2(_0418_));
 sg13g2_xnor2_1 _2036_ (.Y(_0425_),
    .A(_0423_),
    .B(_0424_));
 sg13g2_a22oi_1 _2037_ (.Y(_0426_),
    .B1(net273),
    .B2(net286),
    .A2(net62),
    .A1(net277));
 sg13g2_o21ai_1 _2038_ (.B1(_0426_),
    .Y(_0159_),
    .A1(_0388_),
    .A2(_0425_));
 sg13g2_a21oi_1 _2039_ (.A1(_0422_),
    .A2(_0424_),
    .Y(_0427_),
    .B1(_0421_));
 sg13g2_nor2_1 _2040_ (.A(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.sprite_x[3] ),
    .B(net280),
    .Y(_0428_));
 sg13g2_xnor2_1 _2041_ (.Y(_0429_),
    .A(net193),
    .B(net280));
 sg13g2_xnor2_1 _2042_ (.Y(_0430_),
    .A(_0427_),
    .B(_0429_));
 sg13g2_a22oi_1 _2043_ (.Y(_0431_),
    .B1(net273),
    .B2(net285),
    .A2(net59),
    .A1(net277));
 sg13g2_o21ai_1 _2044_ (.B1(_0431_),
    .Y(_0160_),
    .A1(_0388_),
    .A2(_0430_));
 sg13g2_xnor2_1 _2045_ (.Y(_0432_),
    .A(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.sprite_x[4] ),
    .B(net280));
 sg13g2_a221oi_1 _2046_ (.B2(_0424_),
    .C1(_0421_),
    .B1(_0423_),
    .A1(net285),
    .Y(_0433_),
    .A2(net280));
 sg13g2_nor3_1 _2047_ (.A(_0428_),
    .B(_0432_),
    .C(_0433_),
    .Y(_0434_));
 sg13g2_o21ai_1 _2048_ (.B1(_0432_),
    .Y(_0435_),
    .A1(_0428_),
    .A2(_0433_));
 sg13g2_nand2_1 _2049_ (.Y(_0436_),
    .A(_0387_),
    .B(_0435_));
 sg13g2_a22oi_1 _2050_ (.Y(_0437_),
    .B1(net272),
    .B2(net166),
    .A2(net81),
    .A1(net277));
 sg13g2_o21ai_1 _2051_ (.B1(_0437_),
    .Y(_0161_),
    .A1(_0434_),
    .A2(_0436_));
 sg13g2_xnor2_1 _2052_ (.Y(_0438_),
    .A(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.sprite_x[5] ),
    .B(net280));
 sg13g2_a21oi_1 _2053_ (.A1(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.sprite_x[4] ),
    .A2(net280),
    .Y(_0439_),
    .B1(_0434_));
 sg13g2_xnor2_1 _2054_ (.Y(_0440_),
    .A(_0438_),
    .B(_0439_));
 sg13g2_a22oi_1 _2055_ (.Y(_0441_),
    .B1(net251),
    .B2(net273),
    .A2(net277),
    .A1(net403));
 sg13g2_o21ai_1 _2056_ (.B1(_0441_),
    .Y(_0162_),
    .A1(_0388_),
    .A2(_0440_));
 sg13g2_nand2_1 _2057_ (.Y(_0442_),
    .A(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.sprite_x[6] ),
    .B(net281));
 sg13g2_xor2_1 _2058_ (.B(net281),
    .A(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.sprite_x[6] ),
    .X(_0443_));
 sg13g2_o21ai_1 _2059_ (.B1(net281),
    .Y(_0444_),
    .A1(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.sprite_x[5] ),
    .A2(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.sprite_x[4] ));
 sg13g2_inv_1 _2060_ (.Y(_0445_),
    .A(_0444_));
 sg13g2_nor4_2 _2061_ (.A(_0428_),
    .B(_0432_),
    .C(_0433_),
    .Y(_0446_),
    .D(_0438_));
 sg13g2_o21ai_1 _2062_ (.B1(_0443_),
    .Y(_0447_),
    .A1(_0445_),
    .A2(_0446_));
 sg13g2_or3_1 _2063_ (.A(_0443_),
    .B(_0445_),
    .C(_0446_),
    .X(_0448_));
 sg13g2_nand2_1 _2064_ (.Y(_0449_),
    .A(_0447_),
    .B(_0448_));
 sg13g2_a22oi_1 _2065_ (.Y(_0163_),
    .B1(_0387_),
    .B2(_0449_),
    .A2(net272),
    .A1(_0546_));
 sg13g2_xnor2_1 _2066_ (.Y(_0450_),
    .A(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.sprite_x[7] ),
    .B(net281));
 sg13g2_a21oi_1 _2067_ (.A1(_0442_),
    .A2(_0447_),
    .Y(_0451_),
    .B1(_0450_));
 sg13g2_nand3_1 _2068_ (.B(_0447_),
    .C(_0450_),
    .A(_0442_),
    .Y(_0452_));
 sg13g2_nor2_1 _2069_ (.A(_0372_),
    .B(_0451_),
    .Y(_0453_));
 sg13g2_a22oi_1 _2070_ (.Y(_0454_),
    .B1(_0452_),
    .B2(_0453_),
    .A2(net272),
    .A1(net151));
 sg13g2_inv_1 _2071_ (.Y(_0164_),
    .A(_0454_));
 sg13g2_and2_1 _2072_ (.A(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.sprite_x[8] ),
    .B(net281),
    .X(_0455_));
 sg13g2_xor2_1 _2073_ (.B(net281),
    .A(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.sprite_x[8] ),
    .X(_0456_));
 sg13g2_nand2_1 _2074_ (.Y(_0457_),
    .A(_0443_),
    .B(_0446_));
 sg13g2_nand2_1 _2075_ (.Y(_0458_),
    .A(_0442_),
    .B(_0444_));
 sg13g2_a21oi_1 _2076_ (.A1(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.sprite_x[7] ),
    .A2(net281),
    .Y(_0459_),
    .B1(_0458_));
 sg13g2_o21ai_1 _2077_ (.B1(_0459_),
    .Y(_0460_),
    .A1(_0450_),
    .A2(_0457_));
 sg13g2_xnor2_1 _2078_ (.Y(_0461_),
    .A(_0456_),
    .B(_0460_));
 sg13g2_a22oi_1 _2079_ (.Y(_0165_),
    .B1(_0387_),
    .B2(_0461_),
    .A2(net272),
    .A1(_0542_));
 sg13g2_a21oi_1 _2080_ (.A1(_0456_),
    .A2(_0460_),
    .Y(_0462_),
    .B1(_0455_));
 sg13g2_xnor2_1 _2081_ (.Y(_0463_),
    .A(net411),
    .B(net281));
 sg13g2_a21oi_1 _2082_ (.A1(_0462_),
    .A2(_0463_),
    .Y(_0464_),
    .B1(_0372_));
 sg13g2_o21ai_1 _2083_ (.B1(_0464_),
    .Y(_0465_),
    .A1(_0462_),
    .A2(_0463_));
 sg13g2_o21ai_1 _2084_ (.B1(_0465_),
    .Y(_0166_),
    .A1(_0541_),
    .A2(_0365_));
 sg13g2_nor4_2 _2085_ (.A(_0538_),
    .B(_0775_),
    .C(_0791_),
    .Y(_0466_),
    .D(_0825_));
 sg13g2_mux2_1 _2086_ (.A0(net187),
    .A1(_0841_),
    .S(_0466_),
    .X(_0167_));
 sg13g2_nand2b_1 _2087_ (.Y(_0467_),
    .B(_0840_),
    .A_N(_0832_));
 sg13g2_nand2_1 _2088_ (.Y(_0468_),
    .A(_0838_),
    .B(_0839_));
 sg13g2_and3_1 _2089_ (.X(_0469_),
    .A(_0829_),
    .B(_0467_),
    .C(_0468_));
 sg13g2_mux2_1 _2090_ (.A0(net200),
    .A1(_0469_),
    .S(_0466_),
    .X(_0168_));
 sg13g2_o21ai_1 _2091_ (.B1(net382),
    .Y(_0470_),
    .A1(net2),
    .A2(net1));
 sg13g2_o21ai_1 _2092_ (.B1(_0470_),
    .Y(_0471_),
    .A1(\i_game_and_vga.i_game_top.master_fsm.sprite_torpedo_enable_update ),
    .A2(net259));
 sg13g2_inv_1 _2093_ (.Y(_0169_),
    .A(net260));
 sg13g2_or2_1 _2094_ (.X(_0170_),
    .B(net283),
    .A(net382));
 sg13g2_and2_1 _2095_ (.A(net2),
    .B(net1),
    .X(_0472_));
 sg13g2_nand2b_1 _2096_ (.Y(_0473_),
    .B(net167),
    .A_N(net382));
 sg13g2_o21ai_1 _2097_ (.B1(_0473_),
    .Y(_0171_),
    .A1(_0470_),
    .A2(_0472_));
 sg13g2_nand2_1 _2098_ (.Y(_0474_),
    .A(net382),
    .B(net2));
 sg13g2_nand2b_1 _2099_ (.Y(_0475_),
    .B(net282),
    .A_N(net382));
 sg13g2_o21ai_1 _2100_ (.B1(_0475_),
    .Y(_0172_),
    .A1(net1),
    .A2(_0474_));
 sg13g2_o21ai_1 _2101_ (.B1(net339),
    .Y(_0476_),
    .A1(\i_game_and_vga.i_game_top.end_of_game_timer_start ),
    .A2(\i_game_and_vga.i_game_top.end_of_game_timer_running ));
 sg13g2_nor2_2 _2102_ (.A(\i_game_and_vga.i_game_top.end_of_game_timer_start ),
    .B(net271),
    .Y(_0477_));
 sg13g2_a22oi_1 _2103_ (.Y(_0478_),
    .B1(_0477_),
    .B2(net74),
    .A2(net271),
    .A1(\i_game_and_vga.i_game_top.timer.counter[0] ));
 sg13g2_inv_1 _2104_ (.Y(_0173_),
    .A(net75));
 sg13g2_nor2_1 _2105_ (.A(_0536_),
    .B(_0538_),
    .Y(_0479_));
 sg13g2_nand2_2 _2106_ (.Y(_0480_),
    .A(\i_game_and_vga.i_game_top.end_of_game_timer_start ),
    .B(net339));
 sg13g2_nor3_2 _2107_ (.A(\i_game_and_vga.i_game_top.timer.counter[0] ),
    .B(net400),
    .C(net271),
    .Y(_0481_));
 sg13g2_o21ai_1 _2108_ (.B1(net400),
    .Y(_0482_),
    .A1(\i_game_and_vga.i_game_top.timer.counter[0] ),
    .A2(_0476_));
 sg13g2_nor2b_1 _2109_ (.A(net401),
    .B_N(_0482_),
    .Y(_0483_));
 sg13g2_nor2_1 _2110_ (.A(_0479_),
    .B(net402),
    .Y(_0174_));
 sg13g2_nor2b_1 _2111_ (.A(\i_game_and_vga.i_game_top.timer.counter[2] ),
    .B_N(_0481_),
    .Y(_0484_));
 sg13g2_xnor2_1 _2112_ (.Y(_0485_),
    .A(net263),
    .B(_0481_));
 sg13g2_nor2_1 _2113_ (.A(_0479_),
    .B(net264),
    .Y(_0175_));
 sg13g2_o21ai_1 _2114_ (.B1(_0480_),
    .Y(_0486_),
    .A1(net175),
    .A2(_0484_));
 sg13g2_a21oi_1 _2115_ (.A1(net175),
    .A2(_0484_),
    .Y(_0176_),
    .B1(_0486_));
 sg13g2_or4_2 _2116_ (.A(\i_game_and_vga.i_game_top.timer.counter[0] ),
    .B(\i_game_and_vga.i_game_top.timer.counter[1] ),
    .C(\i_game_and_vga.i_game_top.timer.counter[2] ),
    .D(\i_game_and_vga.i_game_top.timer.counter[3] ),
    .X(_0487_));
 sg13g2_xnor2_1 _2117_ (.Y(_0488_),
    .A(_0622_),
    .B(_0487_));
 sg13g2_a22oi_1 _2118_ (.Y(_0489_),
    .B1(_0477_),
    .B2(_0488_),
    .A2(net271),
    .A1(net361));
 sg13g2_inv_1 _2119_ (.Y(_0177_),
    .A(net362));
 sg13g2_nor3_1 _2120_ (.A(_0622_),
    .B(net271),
    .C(_0487_),
    .Y(_0490_));
 sg13g2_o21ai_1 _2121_ (.B1(_0480_),
    .Y(_0491_),
    .A1(net357),
    .A2(_0490_));
 sg13g2_a21oi_1 _2122_ (.A1(net357),
    .A2(_0490_),
    .Y(_0178_),
    .B1(_0491_));
 sg13g2_nor4_2 _2123_ (.A(\i_game_and_vga.i_game_top.timer.counter[4] ),
    .B(\i_game_and_vga.i_game_top.timer.counter[5] ),
    .C(net271),
    .Y(_0492_),
    .D(_0487_));
 sg13g2_nand2b_1 _2124_ (.Y(_0493_),
    .B(_0492_),
    .A_N(net255));
 sg13g2_nand2b_1 _2125_ (.Y(_0494_),
    .B(net255),
    .A_N(_0492_));
 sg13g2_a21oi_1 _2126_ (.A1(_0493_),
    .A2(_0494_),
    .Y(_0179_),
    .B1(net270));
 sg13g2_xor2_1 _2127_ (.B(_0493_),
    .A(net390),
    .X(_0495_));
 sg13g2_nor2_1 _2128_ (.A(net269),
    .B(_0495_),
    .Y(_0180_));
 sg13g2_o21ai_1 _2129_ (.B1(net243),
    .Y(_0496_),
    .A1(\i_game_and_vga.i_game_top.timer.counter[7] ),
    .A2(_0493_));
 sg13g2_nand3b_1 _2130_ (.B(_0973_),
    .C(_0492_),
    .Y(_0497_),
    .A_N(\i_game_and_vga.i_game_top.timer.counter[6] ));
 sg13g2_a21oi_1 _2131_ (.A1(net244),
    .A2(_0497_),
    .Y(_0181_),
    .B1(net269));
 sg13g2_xor2_1 _2132_ (.B(_0497_),
    .A(net389),
    .X(_0498_));
 sg13g2_nor2_1 _2133_ (.A(net269),
    .B(_0498_),
    .Y(_0182_));
 sg13g2_o21ai_1 _2134_ (.B1(net265),
    .Y(_0499_),
    .A1(\i_game_and_vga.i_game_top.timer.counter[9] ),
    .A2(_0497_));
 sg13g2_nor3_2 _2135_ (.A(\i_game_and_vga.i_game_top.timer.counter[9] ),
    .B(\i_game_and_vga.i_game_top.timer.counter[10] ),
    .C(_0497_),
    .Y(_0500_));
 sg13g2_nand3b_1 _2136_ (.B(_0974_),
    .C(_0492_),
    .Y(_0501_),
    .A_N(net265));
 sg13g2_a21oi_1 _2137_ (.A1(net266),
    .A2(_0501_),
    .Y(_0183_),
    .B1(net269));
 sg13g2_xnor2_1 _2138_ (.Y(_0502_),
    .A(net261),
    .B(_0500_));
 sg13g2_nor2_1 _2139_ (.A(net269),
    .B(net262),
    .Y(_0184_));
 sg13g2_o21ai_1 _2140_ (.B1(net201),
    .Y(_0503_),
    .A1(\i_game_and_vga.i_game_top.timer.counter[11] ),
    .A2(_0501_));
 sg13g2_nand2b_2 _2141_ (.Y(_0504_),
    .B(_0500_),
    .A_N(_0971_));
 sg13g2_a21oi_1 _2142_ (.A1(net202),
    .A2(_0504_),
    .Y(_0185_),
    .B1(net269));
 sg13g2_nor2_1 _2143_ (.A(\i_game_and_vga.i_game_top.timer.counter[13] ),
    .B(_0504_),
    .Y(_0505_));
 sg13g2_xor2_1 _2144_ (.B(_0504_),
    .A(net381),
    .X(_0506_));
 sg13g2_nor2_1 _2145_ (.A(net269),
    .B(_0506_),
    .Y(_0186_));
 sg13g2_nor3_1 _2146_ (.A(\i_game_and_vga.i_game_top.timer.counter[13] ),
    .B(\i_game_and_vga.i_game_top.timer.counter[14] ),
    .C(_0504_),
    .Y(_0507_));
 sg13g2_xnor2_1 _2147_ (.Y(_0508_),
    .A(net253),
    .B(_0505_));
 sg13g2_nor2_1 _2148_ (.A(net269),
    .B(net254),
    .Y(_0187_));
 sg13g2_o21ai_1 _2149_ (.B1(_0480_),
    .Y(_0509_),
    .A1(net164),
    .A2(_0507_));
 sg13g2_a21oi_1 _2150_ (.A1(net164),
    .A2(_0507_),
    .Y(_0188_),
    .B1(_0509_));
 sg13g2_nand2_1 _2151_ (.Y(_0510_),
    .A(_0972_),
    .B(_0500_));
 sg13g2_xor2_1 _2152_ (.B(_0510_),
    .A(net369),
    .X(_0511_));
 sg13g2_nor2_1 _2153_ (.A(net270),
    .B(_0511_),
    .Y(_0189_));
 sg13g2_o21ai_1 _2154_ (.B1(net248),
    .Y(_0512_),
    .A1(\i_game_and_vga.i_game_top.timer.counter[16] ),
    .A2(_0510_));
 sg13g2_nand3_1 _2155_ (.B(_0975_),
    .C(_0500_),
    .A(_0972_),
    .Y(_0513_));
 sg13g2_a21oi_1 _2156_ (.A1(net249),
    .A2(_0513_),
    .Y(_0190_),
    .B1(net270));
 sg13g2_nand2_1 _2157_ (.Y(_0514_),
    .A(net204),
    .B(_0513_));
 sg13g2_or2_1 _2158_ (.X(_0515_),
    .B(_0513_),
    .A(net204));
 sg13g2_a21oi_1 _2159_ (.A1(_0514_),
    .A2(_0515_),
    .Y(_0191_),
    .B1(net270));
 sg13g2_nand2_1 _2160_ (.Y(_0516_),
    .A(net205),
    .B(_0515_));
 sg13g2_or2_1 _2161_ (.X(_0517_),
    .B(_0515_),
    .A(net205));
 sg13g2_a21oi_1 _2162_ (.A1(_0516_),
    .A2(_0517_),
    .Y(_0192_),
    .B1(net270));
 sg13g2_nor2_1 _2163_ (.A(\i_game_and_vga.i_game_top.timer.counter[20] ),
    .B(_0517_),
    .Y(_0518_));
 sg13g2_xor2_1 _2164_ (.B(_0517_),
    .A(net364),
    .X(_0519_));
 sg13g2_nor2_1 _2165_ (.A(net270),
    .B(_0519_),
    .Y(_0193_));
 sg13g2_nor2_1 _2166_ (.A(net152),
    .B(_0518_),
    .Y(_0520_));
 sg13g2_a221oi_1 _2167_ (.B2(_0518_),
    .C1(_0520_),
    .B1(net152),
    .A1(\i_game_and_vga.i_game_top.end_of_game_timer_start ),
    .Y(_0194_),
    .A2(net341));
 sg13g2_nor4_2 _2168_ (.A(\i_game_and_vga.i_game_top.timer.counter[4] ),
    .B(\i_game_and_vga.i_game_top.timer.counter[5] ),
    .C(_0978_),
    .Y(_0521_),
    .D(_0487_));
 sg13g2_nand2_1 _2169_ (.Y(_0522_),
    .A(_0018_),
    .B(_0521_));
 sg13g2_xnor2_1 _2170_ (.Y(_0523_),
    .A(_0018_),
    .B(_0521_));
 sg13g2_a22oi_1 _2171_ (.Y(_0524_),
    .B1(_0477_),
    .B2(_0523_),
    .A2(net271),
    .A1(net190));
 sg13g2_inv_1 _2172_ (.Y(_0195_),
    .A(net191));
 sg13g2_nor2_1 _2173_ (.A(net271),
    .B(_0522_),
    .Y(_0525_));
 sg13g2_o21ai_1 _2174_ (.B1(_0480_),
    .Y(_0526_),
    .A1(net160),
    .A2(_0525_));
 sg13g2_a21oi_1 _2175_ (.A1(net160),
    .A2(_0525_),
    .Y(_0196_),
    .B1(_0526_));
 sg13g2_nand2_1 _2176_ (.Y(_0527_),
    .A(_0979_),
    .B(_0492_));
 sg13g2_a21oi_1 _2177_ (.A1(net149),
    .A2(_0527_),
    .Y(_0528_),
    .B1(net270));
 sg13g2_o21ai_1 _2178_ (.B1(_0528_),
    .Y(_0197_),
    .A1(net149),
    .A2(_0527_));
 sg13g2_and3_1 _2179_ (.X(_0529_),
    .A(net213),
    .B(net239),
    .C(net198));
 sg13g2_nor3_1 _2180_ (.A(net2),
    .B(net1),
    .C(\i_game_and_vga.i_game_top.master_fsm.d_sprite_torpedo_enable_update ),
    .Y(_0530_));
 sg13g2_nor2_1 _2181_ (.A(_0739_),
    .B(_0530_),
    .Y(_0531_));
 sg13g2_a21oi_1 _2182_ (.A1(\i_game_and_vga.i_game_top.master_fsm.d_sprite_target_enable_update ),
    .A2(_0531_),
    .Y(_0198_),
    .B1(_0529_));
 sg13g2_nor4_1 _2183_ (.A(net239),
    .B(net2),
    .C(net1),
    .D(_0739_),
    .Y(_0532_));
 sg13g2_nor3_1 _2184_ (.A(\i_game_and_vga.i_game_top.master_fsm.d_sprite_target_write_dxy ),
    .B(_0529_),
    .C(_0532_),
    .Y(_0199_));
 sg13g2_nand4_1 _2185_ (.B(_0917_),
    .C(_0918_),
    .A(net342),
    .Y(_0533_),
    .D(_0970_));
 sg13g2_mux2_1 _2186_ (.A0(_0878_),
    .A1(net247),
    .S(_0533_),
    .X(_0200_));
 sg13g2_nor3_1 _2187_ (.A(_0845_),
    .B(_0869_),
    .C(_0874_),
    .Y(_0534_));
 sg13g2_mux2_1 _2188_ (.A0(_0534_),
    .A1(net177),
    .S(_0533_),
    .X(_0201_));
 sg13g2_nor2_1 _2189_ (.A(_0833_),
    .B(_0840_),
    .Y(_0535_));
 sg13g2_mux2_1 _2190_ (.A0(net178),
    .A1(_0535_),
    .S(_0466_),
    .X(_0202_));
 sg13g2_dfrbp_1 _2191_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net343),
    .D(_0105_),
    .Q_N(_1059_),
    .Q(\i_game_and_vga.i_game_top.sprite_target.pixel_y[0] ));
 sg13g2_dfrbp_1 _2192_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net343),
    .D(net195),
    .Q_N(_0036_),
    .Q(\i_game_and_vga.i_game_top.sprite_target.pixel_y[1] ));
 sg13g2_dfrbp_1 _2193_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net342),
    .D(_0107_),
    .Q_N(_0030_),
    .Q(\i_game_and_vga.i_game_top.sprite_target.pixel_y[2] ));
 sg13g2_dfrbp_1 _2194_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net343),
    .D(_0108_),
    .Q_N(_1058_),
    .Q(\i_game_and_vga.i_game_top.sprite_target.pixel_y[3] ));
 sg13g2_dfrbp_1 _2195_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net343),
    .D(_0109_),
    .Q_N(_0029_),
    .Q(\i_game_and_vga.i_game_top.sprite_target.pixel_y[4] ));
 sg13g2_dfrbp_1 _2196_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net342),
    .D(net360),
    .Q_N(_0028_),
    .Q(\i_game_and_vga.i_game_top.sprite_target.pixel_y[5] ));
 sg13g2_dfrbp_1 _2197_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net342),
    .D(net399),
    .Q_N(_0027_),
    .Q(\i_game_and_vga.i_game_top.sprite_target.pixel_y[6] ));
 sg13g2_dfrbp_1 _2198_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net342),
    .D(_0112_),
    .Q_N(_0035_),
    .Q(\i_game_and_vga.i_game_top.sprite_target.pixel_y[7] ));
 sg13g2_dfrbp_1 _2199_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net332),
    .D(_0113_),
    .Q_N(_0034_),
    .Q(\i_game_and_vga.i_game_top.sprite_target.pixel_y[8] ));
 sg13g2_dfrbp_1 _2200_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net342),
    .D(_0114_),
    .Q_N(_1057_),
    .Q(\i_game_and_vga.i_vga.vpos[9] ));
 sg13g2_dfrbp_1 _2201_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net350),
    .D(_0115_),
    .Q_N(\i_game_and_vga.i_game_top.sprite_target.sprite_display.y_sprite_plus_h_1[0] ),
    .Q(\i_game_and_vga.i_game_top.sprite_target.sprite_control.sprite_y[0] ));
 sg13g2_dfrbp_1 _2202_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net347),
    .D(net85),
    .Q_N(_1056_),
    .Q(\i_game_and_vga.i_game_top.sprite_target.sprite_control.sprite_y[1] ));
 sg13g2_dfrbp_1 _2203_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net350),
    .D(_0117_),
    .Q_N(_1055_),
    .Q(\i_game_and_vga.i_game_top.sprite_target.sprite_control.sprite_y[2] ));
 sg13g2_dfrbp_1 _2204_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net350),
    .D(net70),
    .Q_N(_1054_),
    .Q(\i_game_and_vga.i_game_top.sprite_target.sprite_control.sprite_y[3] ));
 sg13g2_dfrbp_1 _2205_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net349),
    .D(_0119_),
    .Q_N(_1053_),
    .Q(\i_game_and_vga.i_game_top.sprite_target.sprite_control.sprite_y[4] ));
 sg13g2_dfrbp_1 _2206_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net342),
    .D(_0120_),
    .Q_N(_1052_),
    .Q(\i_game_and_vga.i_game_top.sprite_target.sprite_control.sprite_y[5] ));
 sg13g2_dfrbp_1 _2207_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net330),
    .D(_0121_),
    .Q_N(_1060_),
    .Q(\i_game_and_vga.i_game_top.sprite_target.sprite_control.sprite_y[6] ));
 sg13g2_dfrbp_1 _2208_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net335),
    .D(net93),
    .Q_N(_1061_),
    .Q(\i_game_and_vga.i_vga.clk_en ));
 sg13g2_dfrbp_1 _2209_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net350),
    .D(net157),
    .Q_N(_1062_),
    .Q(\i_game_and_vga.i_game_top.overlap.top_1[0] ));
 sg13g2_dfrbp_1 _2210_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net350),
    .D(net310),
    .Q_N(_1063_),
    .Q(\i_game_and_vga.i_game_top.overlap.top_1[1] ));
 sg13g2_dfrbp_1 _2211_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net349),
    .D(net80),
    .Q_N(_1064_),
    .Q(\i_game_and_vga.i_game_top.overlap.top_1[2] ));
 sg13g2_dfrbp_1 _2212_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net349),
    .D(net68),
    .Q_N(_1065_),
    .Q(\i_game_and_vga.i_game_top.overlap.top_1[3] ));
 sg13g2_dfrbp_1 _2213_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net351),
    .D(net78),
    .Q_N(_1066_),
    .Q(\i_game_and_vga.i_game_top.overlap.top_1[4] ));
 sg13g2_dfrbp_1 _2214_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net330),
    .D(net79),
    .Q_N(_1067_),
    .Q(\i_game_and_vga.i_game_top.overlap.top_1[5] ));
 sg13g2_dfrbp_1 _2215_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net330),
    .D(net66),
    .Q_N(_1051_),
    .Q(\i_game_and_vga.i_game_top.overlap.top_1[6] ));
 sg13g2_dfrbp_1 _2216_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net339),
    .D(_0122_),
    .Q_N(_1050_),
    .Q(\i_game_and_vga.display_on ));
 sg13g2_dfrbp_1 _2217_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net340),
    .D(_0123_),
    .Q_N(_1068_),
    .Q(hsync));
 sg13g2_dfrbp_1 _2218_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net335),
    .D(_0011_),
    .Q_N(_1069_),
    .Q(\i_game_and_vga.i_vga.clk_en_cnt[0] ));
 sg13g2_dfrbp_1 _2219_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net334),
    .D(_0012_),
    .Q_N(_1070_),
    .Q(\i_game_and_vga.i_vga.clk_en_cnt[1] ));
 sg13g2_dfrbp_1 _2220_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net335),
    .D(_0013_),
    .Q_N(_1071_),
    .Q(\i_game_and_vga.i_vga.clk_en_cnt[2] ));
 sg13g2_dfrbp_1 _2221_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net335),
    .D(net156),
    .Q_N(_1049_),
    .Q(\i_game_and_vga.i_vga.clk_en_cnt[3] ));
 sg13g2_dfrbp_1 _2222_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net346),
    .D(net237),
    .Q_N(_1048_),
    .Q(\i_game_and_vga.i_vga.vsync ));
 sg13g2_dfrbp_1 _2223_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net322),
    .D(_0125_),
    .Q_N(_1047_),
    .Q(\i_game_and_vga.i_game_top.sprite_target.pixel_x[0] ));
 sg13g2_dfrbp_1 _2224_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net322),
    .D(_0126_),
    .Q_N(_1046_),
    .Q(\i_game_and_vga.i_game_top.sprite_target.pixel_x[1] ));
 sg13g2_dfrbp_1 _2225_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net322),
    .D(_0127_),
    .Q_N(_0024_),
    .Q(\i_game_and_vga.i_game_top.sprite_target.pixel_x[2] ));
 sg13g2_dfrbp_1 _2226_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net322),
    .D(net375),
    .Q_N(_1045_),
    .Q(\i_game_and_vga.i_game_top.sprite_target.pixel_x[3] ));
 sg13g2_dfrbp_1 _2227_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net317),
    .D(_0129_),
    .Q_N(_0023_),
    .Q(\i_game_and_vga.i_game_top.sprite_target.pixel_x[4] ));
 sg13g2_dfrbp_1 _2228_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net317),
    .D(net386),
    .Q_N(_0022_),
    .Q(\i_game_and_vga.i_game_top.sprite_target.pixel_x[5] ));
 sg13g2_dfrbp_1 _2229_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net328),
    .D(_0131_),
    .Q_N(_0021_),
    .Q(\i_game_and_vga.i_game_top.sprite_target.pixel_x[6] ));
 sg13g2_dfrbp_1 _2230_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net328),
    .D(net405),
    .Q_N(_1044_),
    .Q(\i_game_and_vga.i_game_top.sprite_target.pixel_x[7] ));
 sg13g2_dfrbp_1 _2231_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net328),
    .D(net413),
    .Q_N(_0019_),
    .Q(\i_game_and_vga.i_game_top.sprite_target.pixel_x[8] ));
 sg13g2_dfrbp_1 _2232_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net328),
    .D(_0134_),
    .Q_N(_1043_),
    .Q(\i_game_and_vga.i_game_top.sprite_target.pixel_x[9] ));
 sg13g2_dfrbp_1 _2233_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net348),
    .D(net49),
    .Q_N(\i_game_and_vga.i_game_top.mixer.random ),
    .Q(_0068_));
 sg13g2_dfrbp_1 _2234_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net346),
    .D(net224),
    .Q_N(\i_game_and_vga.i_game_top.random[1] ),
    .Q(_0069_));
 sg13g2_dfrbp_1 _2235_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net346),
    .D(_0088_),
    .Q_N(\i_game_and_vga.i_game_top.random[2] ),
    .Q(_0070_));
 sg13g2_dfrbp_1 _2236_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net347),
    .D(net72),
    .Q_N(\i_game_and_vga.i_game_top.random[3] ),
    .Q(_0071_));
 sg13g2_dfrbp_1 _2237_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net348),
    .D(_0090_),
    .Q_N(\i_game_and_vga.i_game_top.random[4] ),
    .Q(_0072_));
 sg13g2_dfrbp_1 _2238_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net332),
    .D(_0091_),
    .Q_N(\i_game_and_vga.i_game_top.random[5] ),
    .Q(_0073_));
 sg13g2_dfrbp_1 _2239_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net319),
    .D(_0092_),
    .Q_N(\i_game_and_vga.i_game_top.random[6] ),
    .Q(_0074_));
 sg13g2_dfrbp_1 _2240_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net319),
    .D(_0093_),
    .Q_N(\i_game_and_vga.i_game_top.random[7] ),
    .Q(_0075_));
 sg13g2_dfrbp_1 _2241_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net319),
    .D(_0094_),
    .Q_N(\i_game_and_vga.i_game_top.random[8] ),
    .Q(_0076_));
 sg13g2_dfrbp_1 _2242_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net337),
    .D(_0095_),
    .Q_N(\i_game_and_vga.i_game_top.random[9] ),
    .Q(_0077_));
 sg13g2_dfrbp_1 _2243_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net337),
    .D(_0096_),
    .Q_N(\i_game_and_vga.i_game_top.random[10] ),
    .Q(_0078_));
 sg13g2_dfrbp_1 _2244_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net338),
    .D(_0097_),
    .Q_N(\i_game_and_vga.i_game_top.random[11] ),
    .Q(_0079_));
 sg13g2_dfrbp_1 _2245_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net338),
    .D(net65),
    .Q_N(\i_game_and_vga.i_game_top.random[12] ),
    .Q(_0080_));
 sg13g2_dfrbp_1 _2246_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net338),
    .D(net62),
    .Q_N(_1072_),
    .Q(\i_game_and_vga.i_game_top.random[13] ));
 sg13g2_dfrbp_1 _2247_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net337),
    .D(net59),
    .Q_N(_1073_),
    .Q(\i_game_and_vga.i_game_top.random[14] ));
 sg13g2_dfrbp_1 _2248_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net348),
    .D(net81),
    .Q_N(_1074_),
    .Q(\i_game_and_vga.i_game_top.random[15] ));
 sg13g2_dfrbp_1 _2249_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net339),
    .D(_0005_),
    .Q_N(_1075_),
    .Q(\i_game_and_vga.i_game_top.mixer.sprite_target_rgb_en ));
 sg13g2_dfrbp_1 _2250_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net328),
    .D(net209),
    .Q_N(_1076_),
    .Q(\i_game_and_vga.i_game_top.master_fsm.sprite_target_within_screen ));
 sg13g2_dfrbp_1 _2251_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net350),
    .D(net52),
    .Q_N(_1077_),
    .Q(\i_game_and_vga.i_game_top.overlap.bottom_1[0] ));
 sg13g2_dfrbp_1 _2252_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net351),
    .D(\i_game_and_vga.i_game_top.sprite_target.sprite_display.y_sprite_plus_h_1[1] ),
    .Q_N(_1078_),
    .Q(\i_game_and_vga.i_game_top.overlap.bottom_1[1] ));
 sg13g2_dfrbp_1 _2253_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net344),
    .D(\i_game_and_vga.i_game_top.sprite_target.sprite_display.y_sprite_plus_h_1[2] ),
    .Q_N(_1079_),
    .Q(\i_game_and_vga.i_game_top.overlap.bottom_1[2] ));
 sg13g2_dfrbp_1 _2254_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net344),
    .D(\i_game_and_vga.i_game_top.sprite_target.sprite_display.y_sprite_plus_h_1[3] ),
    .Q_N(_1080_),
    .Q(\i_game_and_vga.i_game_top.overlap.bottom_1[3] ));
 sg13g2_dfrbp_1 _2255_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net344),
    .D(\i_game_and_vga.i_game_top.sprite_target.sprite_display.y_sprite_plus_h_1[4] ),
    .Q_N(_1081_),
    .Q(\i_game_and_vga.i_game_top.overlap.bottom_1[4] ));
 sg13g2_dfrbp_1 _2256_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net345),
    .D(\i_game_and_vga.i_game_top.sprite_target.sprite_display.y_sprite_plus_h_1[5] ),
    .Q_N(_1082_),
    .Q(\i_game_and_vga.i_game_top.overlap.bottom_1[5] ));
 sg13g2_dfrbp_1 _2257_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net333),
    .D(\i_game_and_vga.i_game_top.sprite_target.sprite_display.y_sprite_plus_h_1[6] ),
    .Q_N(_1083_),
    .Q(\i_game_and_vga.i_game_top.overlap.bottom_1[6] ));
 sg13g2_dfrbp_1 _2258_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net331),
    .D(\i_game_and_vga.i_game_top.sprite_target.sprite_display.y_sprite_plus_h_1[7] ),
    .Q_N(_1084_),
    .Q(\i_game_and_vga.i_game_top.overlap.bottom_1[7] ));
 sg13g2_dfrbp_1 _2259_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net322),
    .D(net303),
    .Q_N(_1085_),
    .Q(\i_game_and_vga.i_game_top.overlap.left_1[0] ));
 sg13g2_dfrbp_1 _2260_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net317),
    .D(net302),
    .Q_N(_1086_),
    .Q(\i_game_and_vga.i_game_top.overlap.left_1[1] ));
 sg13g2_dfrbp_1 _2261_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net317),
    .D(net89),
    .Q_N(_1087_),
    .Q(\i_game_and_vga.i_game_top.overlap.left_1[2] ));
 sg13g2_dfrbp_1 _2262_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net317),
    .D(net301),
    .Q_N(_1088_),
    .Q(\i_game_and_vga.i_game_top.overlap.left_1[3] ));
 sg13g2_dfrbp_1 _2263_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net318),
    .D(net300),
    .Q_N(_1089_),
    .Q(\i_game_and_vga.i_game_top.overlap.left_1[4] ));
 sg13g2_dfrbp_1 _2264_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net316),
    .D(net222),
    .Q_N(_1090_),
    .Q(\i_game_and_vga.i_game_top.overlap.left_1[5] ));
 sg13g2_dfrbp_1 _2265_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net327),
    .D(net97),
    .Q_N(_1091_),
    .Q(\i_game_and_vga.i_game_top.overlap.left_1[6] ));
 sg13g2_dfrbp_1 _2266_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net326),
    .D(net192),
    .Q_N(_1092_),
    .Q(\i_game_and_vga.i_game_top.overlap.left_1[7] ));
 sg13g2_dfrbp_1 _2267_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net326),
    .D(net299),
    .Q_N(_1093_),
    .Q(\i_game_and_vga.i_game_top.overlap.left_1[8] ));
 sg13g2_dfrbp_1 _2268_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net329),
    .D(net298),
    .Q_N(_1094_),
    .Q(\i_game_and_vga.i_game_top.overlap.left_1[9] ));
 sg13g2_dfrbp_1 _2269_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net323),
    .D(net54),
    .Q_N(_1095_),
    .Q(\i_game_and_vga.i_game_top.overlap.right_1[0] ));
 sg13g2_dfrbp_1 _2270_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net323),
    .D(net136),
    .Q_N(_1096_),
    .Q(\i_game_and_vga.i_game_top.overlap.right_1[1] ));
 sg13g2_dfrbp_1 _2271_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net322),
    .D(\i_game_and_vga.i_game_top.sprite_target.sprite_display.x_sprite_plus_w_1[2] ),
    .Q_N(_1097_),
    .Q(\i_game_and_vga.i_game_top.overlap.right_1[2] ));
 sg13g2_dfrbp_1 _2272_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net317),
    .D(\i_game_and_vga.i_game_top.sprite_target.sprite_display.x_sprite_plus_w_1[3] ),
    .Q_N(_1098_),
    .Q(\i_game_and_vga.i_game_top.overlap.right_1[3] ));
 sg13g2_dfrbp_1 _2273_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net317),
    .D(\i_game_and_vga.i_game_top.sprite_target.sprite_display.x_sprite_plus_w_1[4] ),
    .Q_N(_1099_),
    .Q(\i_game_and_vga.i_game_top.overlap.right_1[4] ));
 sg13g2_dfrbp_1 _2274_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net327),
    .D(\i_game_and_vga.i_game_top.sprite_target.sprite_display.x_sprite_plus_w_1[5] ),
    .Q_N(_1100_),
    .Q(\i_game_and_vga.i_game_top.overlap.right_1[5] ));
 sg13g2_dfrbp_1 _2275_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net326),
    .D(\i_game_and_vga.i_game_top.sprite_target.sprite_display.x_sprite_plus_w_1[6] ),
    .Q_N(_1101_),
    .Q(\i_game_and_vga.i_game_top.overlap.right_1[6] ));
 sg13g2_dfrbp_1 _2276_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net326),
    .D(\i_game_and_vga.i_game_top.sprite_target.sprite_display.x_sprite_plus_w_1[7] ),
    .Q_N(_1102_),
    .Q(\i_game_and_vga.i_game_top.overlap.right_1[7] ));
 sg13g2_dfrbp_1 _2277_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net326),
    .D(\i_game_and_vga.i_game_top.sprite_target.sprite_display.x_sprite_plus_w_1[8] ),
    .Q_N(_1103_),
    .Q(\i_game_and_vga.i_game_top.overlap.right_1[8] ));
 sg13g2_dfrbp_1 _2278_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net326),
    .D(\i_game_and_vga.i_game_top.sprite_target.sprite_display.x_sprite_plus_w_1[9] ),
    .Q_N(_1042_),
    .Q(\i_game_and_vga.i_game_top.overlap.right_1[9] ));
 sg13g2_dfrbp_1 _2279_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net323),
    .D(_0135_),
    .Q_N(\i_game_and_vga.i_game_top.sprite_target.sprite_display.x_sprite_plus_w_1[0] ),
    .Q(\i_game_and_vga.i_game_top.sprite_target.sprite_control.sprite_x[0] ));
 sg13g2_dfrbp_1 _2280_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net321),
    .D(_0136_),
    .Q_N(_1041_),
    .Q(\i_game_and_vga.i_game_top.sprite_target.sprite_control.sprite_x[1] ));
 sg13g2_dfrbp_1 _2281_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net314),
    .D(_0137_),
    .Q_N(_1040_),
    .Q(\i_game_and_vga.i_game_top.sprite_target.sprite_control.sprite_x[2] ));
 sg13g2_dfrbp_1 _2282_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net316),
    .D(_0138_),
    .Q_N(_1039_),
    .Q(\i_game_and_vga.i_game_top.sprite_target.sprite_control.sprite_x[3] ));
 sg13g2_dfrbp_1 _2283_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net316),
    .D(_0139_),
    .Q_N(_1038_),
    .Q(\i_game_and_vga.i_game_top.sprite_target.sprite_control.sprite_x[4] ));
 sg13g2_dfrbp_1 _2284_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net316),
    .D(_0140_),
    .Q_N(_1037_),
    .Q(\i_game_and_vga.i_game_top.sprite_target.sprite_control.sprite_x[5] ));
 sg13g2_dfrbp_1 _2285_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net318),
    .D(_0141_),
    .Q_N(_0033_),
    .Q(\i_game_and_vga.i_game_top.sprite_target.sprite_control.sprite_x[6] ));
 sg13g2_dfrbp_1 _2286_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net316),
    .D(_0142_),
    .Q_N(_1036_),
    .Q(\i_game_and_vga.i_game_top.sprite_target.sprite_control.sprite_x[7] ));
 sg13g2_dfrbp_1 _2287_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net316),
    .D(_0143_),
    .Q_N(_1035_),
    .Q(\i_game_and_vga.i_game_top.sprite_target.sprite_control.sprite_x[8] ));
 sg13g2_dfrbp_1 _2288_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net316),
    .D(_0144_),
    .Q_N(_1034_),
    .Q(\i_game_and_vga.i_game_top.sprite_target.sprite_control.sprite_x[9] ));
 sg13g2_dfrbp_1 _2289_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net346),
    .D(net77),
    .Q_N(_1033_),
    .Q(\i_game_and_vga.i_game_top.game_won ));
 sg13g2_dfrbp_1 _2290_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net320),
    .D(_0146_),
    .Q_N(_1032_),
    .Q(\i_game_and_vga.i_game_top.sprite_target.sprite_control.dx[0] ));
 sg13g2_dfrbp_1 _2291_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net321),
    .D(_0147_),
    .Q_N(_1104_),
    .Q(\i_game_and_vga.i_game_top.sprite_target.sprite_control.dx[1] ));
 sg13g2_dfrbp_1 _2292_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net315),
    .D(net51),
    .Q_N(_0983_),
    .Q(\i_game_and_vga.i_game_top.sprite_target.sprite_control.strobe_generator.counter[0] ));
 sg13g2_dfrbp_1 _2293_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net315),
    .D(net148),
    .Q_N(\i_game_and_vga.i_game_top.sprite_target.sprite_control.strobe_generator.counter[1] ),
    .Q(_0081_));
 sg13g2_dfrbp_1 _2294_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net315),
    .D(net140),
    .Q_N(\i_game_and_vga.i_game_top.sprite_target.sprite_control.strobe_generator.counter[2] ),
    .Q(_0082_));
 sg13g2_dfrbp_1 _2295_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net321),
    .D(net127),
    .Q_N(_1105_),
    .Q(\i_game_and_vga.i_game_top.sprite_target.sprite_control.strobe_generator.counter[3] ));
 sg13g2_dfrbp_1 _2296_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net321),
    .D(net221),
    .Q_N(_1031_),
    .Q(\i_game_and_vga.i_game_top.sprite_target.sprite_control.strobe_generator.counter[4] ));
 sg13g2_dfrbp_1 _2297_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net321),
    .D(net174),
    .Q_N(\i_game_and_vga.i_game_top.sprite_target.sprite_control.strobe_generator.counter[5] ),
    .Q(_0083_));
 sg13g2_dfrbp_1 _2298_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net319),
    .D(net129),
    .Q_N(_1106_),
    .Q(\i_game_and_vga.i_game_top.sprite_target.sprite_control.strobe_generator.counter[6] ));
 sg13g2_dfrbp_1 _2299_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net319),
    .D(net132),
    .Q_N(_1107_),
    .Q(\i_game_and_vga.i_game_top.sprite_target.sprite_control.strobe_generator.counter[7] ));
 sg13g2_dfrbp_1 _2300_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net319),
    .D(net207),
    .Q_N(_1108_),
    .Q(\i_game_and_vga.i_game_top.sprite_target.sprite_control.strobe_generator.counter[8] ));
 sg13g2_dfrbp_1 _2301_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net319),
    .D(_0051_),
    .Q_N(_1109_),
    .Q(\i_game_and_vga.i_game_top.sprite_target.sprite_control.strobe_generator.counter[9] ));
 sg13g2_dfrbp_1 _2302_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net319),
    .D(net115),
    .Q_N(_1110_),
    .Q(\i_game_and_vga.i_game_top.sprite_target.sprite_control.strobe_generator.counter[10] ));
 sg13g2_dfrbp_1 _2303_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net334),
    .D(net171),
    .Q_N(_1111_),
    .Q(\i_game_and_vga.i_game_top.sprite_target.sprite_control.strobe_generator.counter[11] ));
 sg13g2_dfrbp_1 _2304_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net334),
    .D(_0039_),
    .Q_N(_1112_),
    .Q(\i_game_and_vga.i_game_top.sprite_target.sprite_control.strobe_generator.counter[12] ));
 sg13g2_dfrbp_1 _2305_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net334),
    .D(net123),
    .Q_N(_1113_),
    .Q(\i_game_and_vga.i_game_top.sprite_target.sprite_control.strobe_generator.counter[13] ));
 sg13g2_dfrbp_1 _2306_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net336),
    .D(net159),
    .Q_N(_1114_),
    .Q(\i_game_and_vga.i_game_top.sprite_target.sprite_control.strobe_generator.counter[14] ));
 sg13g2_dfrbp_1 _2307_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net336),
    .D(_0042_),
    .Q_N(_1115_),
    .Q(\i_game_and_vga.i_game_top.sprite_target.sprite_control.strobe_generator.counter[15] ));
 sg13g2_dfrbp_1 _2308_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net336),
    .D(net125),
    .Q_N(_1116_),
    .Q(\i_game_and_vga.i_game_top.sprite_target.sprite_control.strobe_generator.counter[16] ));
 sg13g2_dfrbp_1 _2309_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net336),
    .D(_0044_),
    .Q_N(_1117_),
    .Q(\i_game_and_vga.i_game_top.sprite_target.sprite_control.strobe_generator.counter[17] ));
 sg13g2_dfrbp_1 _2310_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net334),
    .D(net105),
    .Q_N(_1118_),
    .Q(\i_game_and_vga.i_game_top.sprite_target.sprite_control.strobe_generator.counter[18] ));
 sg13g2_dfrbp_1 _2311_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net334),
    .D(net112),
    .Q_N(_1119_),
    .Q(\i_game_and_vga.i_game_top.sprite_target.sprite_control.strobe_generator.strobe ));
 sg13g2_dfrbp_1 _2312_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net348),
    .D(_0007_),
    .Q_N(_1120_),
    .Q(\i_game_and_vga.i_game_top.mixer.sprite_torpedo_rgb_en ));
 sg13g2_dfrbp_1 _2313_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net331),
    .D(_0008_),
    .Q_N(_1121_),
    .Q(\i_game_and_vga.i_game_top.master_fsm.sprite_torpedo_within_screen ));
 sg13g2_dfrbp_1 _2314_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net351),
    .D(net56),
    .Q_N(_1122_),
    .Q(\i_game_and_vga.i_game_top.overlap.bottom_2[0] ));
 sg13g2_dfrbp_1 _2315_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net350),
    .D(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_display.y_sprite_plus_h_1[1] ),
    .Q_N(_1123_),
    .Q(\i_game_and_vga.i_game_top.overlap.bottom_2[1] ));
 sg13g2_dfrbp_1 _2316_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net349),
    .D(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_display.y_sprite_plus_h_1[2] ),
    .Q_N(_1124_),
    .Q(\i_game_and_vga.i_game_top.overlap.bottom_2[2] ));
 sg13g2_dfrbp_1 _2317_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net344),
    .D(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_display.y_sprite_plus_h_1[3] ),
    .Q_N(_1125_),
    .Q(\i_game_and_vga.i_game_top.overlap.bottom_2[3] ));
 sg13g2_dfrbp_1 _2318_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net344),
    .D(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_display.y_sprite_plus_h_1[4] ),
    .Q_N(_1126_),
    .Q(\i_game_and_vga.i_game_top.overlap.bottom_2[4] ));
 sg13g2_dfrbp_1 _2319_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net345),
    .D(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_display.y_sprite_plus_h_1[5] ),
    .Q_N(_1127_),
    .Q(\i_game_and_vga.i_game_top.overlap.bottom_2[5] ));
 sg13g2_dfrbp_1 _2320_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net330),
    .D(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_display.y_sprite_plus_h_1[6] ),
    .Q_N(_1128_),
    .Q(\i_game_and_vga.i_game_top.overlap.bottom_2[6] ));
 sg13g2_dfrbp_1 _2321_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net330),
    .D(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_display.y_sprite_plus_h_1[7] ),
    .Q_N(_1129_),
    .Q(\i_game_and_vga.i_game_top.overlap.bottom_2[7] ));
 sg13g2_dfrbp_1 _2322_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net330),
    .D(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_display.y_sprite_plus_h_1[8] ),
    .Q_N(_1130_),
    .Q(\i_game_and_vga.i_game_top.overlap.bottom_2[8] ));
 sg13g2_dfrbp_1 _2323_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net323),
    .D(net288),
    .Q_N(_1131_),
    .Q(\i_game_and_vga.i_game_top.overlap.left_2[0] ));
 sg13g2_dfrbp_1 _2324_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net323),
    .D(net287),
    .Q_N(_1132_),
    .Q(\i_game_and_vga.i_game_top.overlap.left_2[1] ));
 sg13g2_dfrbp_1 _2325_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net323),
    .D(net286),
    .Q_N(_1133_),
    .Q(\i_game_and_vga.i_game_top.overlap.left_2[2] ));
 sg13g2_dfrbp_1 _2326_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net322),
    .D(net285),
    .Q_N(_1134_),
    .Q(\i_game_and_vga.i_game_top.overlap.left_2[3] ));
 sg13g2_dfrbp_1 _2327_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net332),
    .D(net166),
    .Q_N(_1135_),
    .Q(\i_game_and_vga.i_game_top.overlap.left_2[4] ));
 sg13g2_dfrbp_1 _2328_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net328),
    .D(net251),
    .Q_N(_1136_),
    .Q(\i_game_and_vga.i_game_top.overlap.left_2[5] ));
 sg13g2_dfrbp_1 _2329_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net328),
    .D(net154),
    .Q_N(_1137_),
    .Q(\i_game_and_vga.i_game_top.overlap.left_2[6] ));
 sg13g2_dfrbp_1 _2330_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net329),
    .D(net151),
    .Q_N(_1138_),
    .Q(\i_game_and_vga.i_game_top.overlap.left_2[7] ));
 sg13g2_dfrbp_1 _2331_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net329),
    .D(net113),
    .Q_N(_1139_),
    .Q(\i_game_and_vga.i_game_top.overlap.left_2[8] ));
 sg13g2_dfrbp_1 _2332_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net329),
    .D(net91),
    .Q_N(_1030_),
    .Q(\i_game_and_vga.i_game_top.overlap.left_2[9] ));
 sg13g2_dfrbp_1 _2333_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net350),
    .D(net96),
    .Q_N(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_display.y_sprite_plus_h_1[0] ),
    .Q(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.sprite_y[0] ));
 sg13g2_dfrbp_1 _2334_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net349),
    .D(_0149_),
    .Q_N(_1029_),
    .Q(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.sprite_y[1] ));
 sg13g2_dfrbp_1 _2335_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net345),
    .D(_0150_),
    .Q_N(_1028_),
    .Q(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.sprite_y[2] ));
 sg13g2_dfrbp_1 _2336_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net344),
    .D(_0151_),
    .Q_N(_1027_),
    .Q(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.sprite_y[3] ));
 sg13g2_dfrbp_1 _2337_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net345),
    .D(_0152_),
    .Q_N(_1026_),
    .Q(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.sprite_y[4] ));
 sg13g2_dfrbp_1 _2338_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net345),
    .D(_0153_),
    .Q_N(_1025_),
    .Q(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.sprite_y[5] ));
 sg13g2_dfrbp_1 _2339_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net330),
    .D(_0154_),
    .Q_N(_0026_),
    .Q(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.sprite_y[6] ));
 sg13g2_dfrbp_1 _2340_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net331),
    .D(_0155_),
    .Q_N(_1024_),
    .Q(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.sprite_y[7] ));
 sg13g2_dfrbp_1 _2341_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net331),
    .D(_0156_),
    .Q_N(_0025_),
    .Q(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.sprite_y[8] ));
 sg13g2_dfrbp_1 _2342_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net337),
    .D(net50),
    .Q_N(_1140_),
    .Q(\i_game_and_vga.i_game_top.overlap.right_2[0] ));
 sg13g2_dfrbp_1 _2343_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net322),
    .D(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_display.x_sprite_plus_w_1[1] ),
    .Q_N(_1141_),
    .Q(\i_game_and_vga.i_game_top.overlap.right_2[1] ));
 sg13g2_dfrbp_1 _2344_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net317),
    .D(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_display.x_sprite_plus_w_1[2] ),
    .Q_N(_1142_),
    .Q(\i_game_and_vga.i_game_top.overlap.right_2[2] ));
 sg13g2_dfrbp_1 _2345_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net318),
    .D(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_display.x_sprite_plus_w_1[3] ),
    .Q_N(_1143_),
    .Q(\i_game_and_vga.i_game_top.overlap.right_2[3] ));
 sg13g2_dfrbp_1 _2346_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net316),
    .D(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_display.x_sprite_plus_w_1[4] ),
    .Q_N(_1144_),
    .Q(\i_game_and_vga.i_game_top.overlap.right_2[4] ));
 sg13g2_dfrbp_1 _2347_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net327),
    .D(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_display.x_sprite_plus_w_1[5] ),
    .Q_N(_1145_),
    .Q(\i_game_and_vga.i_game_top.overlap.right_2[5] ));
 sg13g2_dfrbp_1 _2348_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net326),
    .D(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_display.x_sprite_plus_w_1[6] ),
    .Q_N(_1146_),
    .Q(\i_game_and_vga.i_game_top.overlap.right_2[6] ));
 sg13g2_dfrbp_1 _2349_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net326),
    .D(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_display.x_sprite_plus_w_1[7] ),
    .Q_N(_1147_),
    .Q(\i_game_and_vga.i_game_top.overlap.right_2[7] ));
 sg13g2_dfrbp_1 _2350_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net327),
    .D(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_display.x_sprite_plus_w_1[8] ),
    .Q_N(_1148_),
    .Q(\i_game_and_vga.i_game_top.overlap.right_2[8] ));
 sg13g2_dfrbp_1 _2351_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net329),
    .D(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_display.x_sprite_plus_w_1[9] ),
    .Q_N(_1149_),
    .Q(\i_game_and_vga.i_game_top.overlap.right_2[9] ));
 sg13g2_dfrbp_1 _2352_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net349),
    .D(net294),
    .Q_N(_1150_),
    .Q(\i_game_and_vga.i_game_top.overlap.top_2[0] ));
 sg13g2_dfrbp_1 _2353_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net349),
    .D(net293),
    .Q_N(_1151_),
    .Q(\i_game_and_vga.i_game_top.overlap.top_2[1] ));
 sg13g2_dfrbp_1 _2354_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net344),
    .D(net291),
    .Q_N(_1152_),
    .Q(\i_game_and_vga.i_game_top.overlap.top_2[2] ));
 sg13g2_dfrbp_1 _2355_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net344),
    .D(net290),
    .Q_N(_1153_),
    .Q(\i_game_and_vga.i_game_top.overlap.top_2[3] ));
 sg13g2_dfrbp_1 _2356_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net345),
    .D(net289),
    .Q_N(_1154_),
    .Q(\i_game_and_vga.i_game_top.overlap.top_2[4] ));
 sg13g2_dfrbp_1 _2357_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net345),
    .D(net102),
    .Q_N(_1155_),
    .Q(\i_game_and_vga.i_game_top.overlap.top_2[5] ));
 sg13g2_dfrbp_1 _2358_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net330),
    .D(net98),
    .Q_N(_1156_),
    .Q(\i_game_and_vga.i_game_top.overlap.top_2[6] ));
 sg13g2_dfrbp_1 _2359_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net331),
    .D(net181),
    .Q_N(_1157_),
    .Q(\i_game_and_vga.i_game_top.overlap.top_2[7] ));
 sg13g2_dfrbp_1 _2360_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net331),
    .D(net82),
    .Q_N(_1023_),
    .Q(\i_game_and_vga.i_game_top.overlap.top_2[8] ));
 sg13g2_dfrbp_1 _2361_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net337),
    .D(net169),
    .Q_N(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_display.x_sprite_plus_w_1[0] ),
    .Q(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.sprite_x[0] ));
 sg13g2_dfrbp_1 _2362_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net337),
    .D(net108),
    .Q_N(_1022_),
    .Q(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.sprite_x[1] ));
 sg13g2_dfrbp_1 _2363_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net337),
    .D(_0159_),
    .Q_N(_1021_),
    .Q(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.sprite_x[2] ));
 sg13g2_dfrbp_1 _2364_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net337),
    .D(_0160_),
    .Q_N(_1020_),
    .Q(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.sprite_x[3] ));
 sg13g2_dfrbp_1 _2365_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net332),
    .D(_0161_),
    .Q_N(_1019_),
    .Q(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.sprite_x[4] ));
 sg13g2_dfrbp_1 _2366_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net342),
    .D(_0162_),
    .Q_N(_1018_),
    .Q(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.sprite_x[5] ));
 sg13g2_dfrbp_1 _2367_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net332),
    .D(_0163_),
    .Q_N(_0020_),
    .Q(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.sprite_x[6] ));
 sg13g2_dfrbp_1 _2368_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net332),
    .D(_0164_),
    .Q_N(_1017_),
    .Q(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.sprite_x[7] ));
 sg13g2_dfrbp_1 _2369_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net332),
    .D(_0165_),
    .Q_N(_1016_),
    .Q(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.sprite_x[8] ));
 sg13g2_dfrbp_1 _2370_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net332),
    .D(_0166_),
    .Q_N(_1015_),
    .Q(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.sprite_x[9] ));
 sg13g2_dfrbp_1 _2371_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net47),
    .D(_0167_),
    .Q_N(_1014_),
    .Q(\i_game_and_vga.i_game_top.mixer.sprite_target_rgb[0] ));
 sg13g2_dfrbp_1 _2372_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net46),
    .D(_0168_),
    .Q_N(_1013_),
    .Q(\i_game_and_vga.i_game_top.mixer.sprite_target_rgb[1] ));
 sg13g2_dfrbp_1 _2373_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net346),
    .D(_0169_),
    .Q_N(_1012_),
    .Q(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.dy[0] ));
 sg13g2_dfrbp_1 _2374_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net349),
    .D(_0170_),
    .Q_N(_1011_),
    .Q(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.dy[1] ));
 sg13g2_dfrbp_1 _2375_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net347),
    .D(_0171_),
    .Q_N(_1010_),
    .Q(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.dx[0] ));
 sg13g2_dfrbp_1 _2376_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net347),
    .D(_0172_),
    .Q_N(_1158_),
    .Q(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.dx[1] ));
 sg13g2_dfrbp_1 _2377_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net314),
    .D(net53),
    .Q_N(_0984_),
    .Q(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.strobe_generator.counter[0] ));
 sg13g2_dfrbp_1 _2378_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net314),
    .D(net117),
    .Q_N(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.strobe_generator.counter[1] ),
    .Q(_0084_));
 sg13g2_dfrbp_1 _2379_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net314),
    .D(net228),
    .Q_N(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.strobe_generator.counter[2] ),
    .Q(_0085_));
 sg13g2_dfrbp_1 _2380_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net314),
    .D(net121),
    .Q_N(_1159_),
    .Q(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.strobe_generator.counter[3] ));
 sg13g2_dfrbp_1 _2381_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net314),
    .D(net235),
    .Q_N(_1009_),
    .Q(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.strobe_generator.counter[4] ));
 sg13g2_dfrbp_1 _2382_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net314),
    .D(net212),
    .Q_N(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.strobe_generator.counter[5] ),
    .Q(_0086_));
 sg13g2_dfrbp_1 _2383_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net314),
    .D(net134),
    .Q_N(_1160_),
    .Q(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.strobe_generator.counter[6] ));
 sg13g2_dfrbp_1 _2384_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net315),
    .D(net146),
    .Q_N(_1161_),
    .Q(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.strobe_generator.counter[7] ));
 sg13g2_dfrbp_1 _2385_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net315),
    .D(net197),
    .Q_N(_1162_),
    .Q(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.strobe_generator.counter[8] ));
 sg13g2_dfrbp_1 _2386_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net315),
    .D(_0066_),
    .Q_N(_1163_),
    .Q(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.strobe_generator.counter[9] ));
 sg13g2_dfrbp_1 _2387_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net315),
    .D(net163),
    .Q_N(_1164_),
    .Q(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.strobe_generator.counter[10] ));
 sg13g2_dfrbp_1 _2388_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net321),
    .D(net184),
    .Q_N(_1165_),
    .Q(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.strobe_generator.counter[11] ));
 sg13g2_dfrbp_1 _2389_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net321),
    .D(_0054_),
    .Q_N(_1166_),
    .Q(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.strobe_generator.counter[12] ));
 sg13g2_dfrbp_1 _2390_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net321),
    .D(net142),
    .Q_N(_1167_),
    .Q(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.strobe_generator.counter[13] ));
 sg13g2_dfrbp_1 _2391_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net320),
    .D(net180),
    .Q_N(_1168_),
    .Q(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.strobe_generator.counter[14] ));
 sg13g2_dfrbp_1 _2392_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net320),
    .D(_0057_),
    .Q_N(_1169_),
    .Q(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.strobe_generator.counter[15] ));
 sg13g2_dfrbp_1 _2393_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net320),
    .D(net119),
    .Q_N(_1170_),
    .Q(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.strobe_generator.counter[16] ));
 sg13g2_dfrbp_1 _2394_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net334),
    .D(_0059_),
    .Q_N(_1171_),
    .Q(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.strobe_generator.counter[17] ));
 sg13g2_dfrbp_1 _2395_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net334),
    .D(net101),
    .Q_N(_1172_),
    .Q(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.strobe_generator.counter[18] ));
 sg13g2_dfrbp_1 _2396_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net338),
    .D(net110),
    .Q_N(_1173_),
    .Q(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.strobe_generator.strobe ));
 sg13g2_dfrbp_1 _2397_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net331),
    .D(net233),
    .Q_N(_1174_),
    .Q(\i_game_and_vga.i_game_top.collision ));
 sg13g2_dfrbp_1 _2398_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net339),
    .D(net366),
    .Q_N(_0031_),
    .Q(\i_game_and_vga.i_game_top.end_of_game_timer_running ));
 sg13g2_dfrbp_1 _2399_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net42),
    .D(_0173_),
    .Q_N(_0067_),
    .Q(\i_game_and_vga.i_game_top.timer.counter[0] ));
 sg13g2_dfrbp_1 _2400_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net40),
    .D(_0174_),
    .Q_N(_1008_),
    .Q(\i_game_and_vga.i_game_top.timer.counter[1] ));
 sg13g2_dfrbp_1 _2401_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net38),
    .D(_0175_),
    .Q_N(_1007_),
    .Q(\i_game_and_vga.i_game_top.timer.counter[2] ));
 sg13g2_dfrbp_1 _2402_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net37),
    .D(net176),
    .Q_N(_1006_),
    .Q(\i_game_and_vga.i_game_top.timer.counter[3] ));
 sg13g2_dfrbp_1 _2403_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net35),
    .D(_0177_),
    .Q_N(_0017_),
    .Q(\i_game_and_vga.i_game_top.timer.counter[4] ));
 sg13g2_dfrbp_1 _2404_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net34),
    .D(net358),
    .Q_N(_1005_),
    .Q(\i_game_and_vga.i_game_top.timer.counter[5] ));
 sg13g2_dfrbp_1 _2405_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net32),
    .D(net256),
    .Q_N(_1004_),
    .Q(\i_game_and_vga.i_game_top.timer.counter[6] ));
 sg13g2_dfrbp_1 _2406_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net30),
    .D(_0180_),
    .Q_N(_1003_),
    .Q(\i_game_and_vga.i_game_top.timer.counter[7] ));
 sg13g2_dfrbp_1 _2407_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net28),
    .D(net245),
    .Q_N(_1002_),
    .Q(\i_game_and_vga.i_game_top.timer.counter[8] ));
 sg13g2_dfrbp_1 _2408_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net27),
    .D(_0182_),
    .Q_N(_1001_),
    .Q(\i_game_and_vga.i_game_top.timer.counter[9] ));
 sg13g2_dfrbp_1 _2409_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net25),
    .D(net354),
    .Q_N(_1000_),
    .Q(\i_game_and_vga.i_game_top.timer.counter[10] ));
 sg13g2_dfrbp_1 _2410_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net24),
    .D(_0184_),
    .Q_N(_0999_),
    .Q(\i_game_and_vga.i_game_top.timer.counter[11] ));
 sg13g2_dfrbp_1 _2411_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net22),
    .D(net203),
    .Q_N(_0998_),
    .Q(\i_game_and_vga.i_game_top.timer.counter[12] ));
 sg13g2_dfrbp_1 _2412_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net20),
    .D(_0186_),
    .Q_N(_0997_),
    .Q(\i_game_and_vga.i_game_top.timer.counter[13] ));
 sg13g2_dfrbp_1 _2413_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net45),
    .D(_0187_),
    .Q_N(_0996_),
    .Q(\i_game_and_vga.i_game_top.timer.counter[14] ));
 sg13g2_dfrbp_1 _2414_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net43),
    .D(net165),
    .Q_N(_0995_),
    .Q(\i_game_and_vga.i_game_top.timer.counter[15] ));
 sg13g2_dfrbp_1 _2415_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net39),
    .D(_0189_),
    .Q_N(_0994_),
    .Q(\i_game_and_vga.i_game_top.timer.counter[16] ));
 sg13g2_dfrbp_1 _2416_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net36),
    .D(net250),
    .Q_N(_0993_),
    .Q(\i_game_and_vga.i_game_top.timer.counter[17] ));
 sg13g2_dfrbp_1 _2417_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net33),
    .D(_0191_),
    .Q_N(_0992_),
    .Q(\i_game_and_vga.i_game_top.timer.counter[18] ));
 sg13g2_dfrbp_1 _2418_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net29),
    .D(_0192_),
    .Q_N(_0991_),
    .Q(\i_game_and_vga.i_game_top.timer.counter[19] ));
 sg13g2_dfrbp_1 _2419_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net26),
    .D(_0193_),
    .Q_N(_0990_),
    .Q(\i_game_and_vga.i_game_top.timer.counter[20] ));
 sg13g2_dfrbp_1 _2420_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net23),
    .D(net153),
    .Q_N(_0989_),
    .Q(\i_game_and_vga.i_game_top.timer.counter[21] ));
 sg13g2_dfrbp_1 _2421_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net19),
    .D(_0195_),
    .Q_N(_0018_),
    .Q(\i_game_and_vga.i_game_top.timer.counter[22] ));
 sg13g2_dfrbp_1 _2422_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net41),
    .D(net161),
    .Q_N(_0988_),
    .Q(\i_game_and_vga.i_game_top.timer.counter[23] ));
 sg13g2_dfrbp_1 _2423_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net48),
    .D(net150),
    .Q_N(_1175_),
    .Q(\i_game_and_vga.i_game_top.timer.counter[24] ));
 sg13g2_dfrbp_1 _2424_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net340),
    .D(net88),
    .Q_N(_1176_),
    .Q(uo_out[6]));
 sg13g2_dfrbp_1 _2425_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net340),
    .D(net219),
    .Q_N(_1177_),
    .Q(uo_out[5]));
 sg13g2_dfrbp_1 _2426_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net340),
    .D(_0002_),
    .Q_N(_1178_),
    .Q(uo_out[4]));
 sg13g2_dfrbp_1 _2427_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net339),
    .D(\i_game_and_vga.i_game_top.master_fsm.d_sprite_target_enable_update ),
    .Q_N(_1179_),
    .Q(\i_game_and_vga.i_game_top.master_fsm.sprite_target_enable_update ));
 sg13g2_dfrbp_1 _2428_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net346),
    .D(net214),
    .Q_N(_1180_),
    .Q(\i_game_and_vga.i_game_top.master_fsm.sprite_torpedo_enable_update ));
 sg13g2_dfrbp_1 _2429_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net339),
    .D(\i_game_and_vga.i_game_top.master_fsm.d_end_of_game_timer_start ),
    .Q_N(_1181_),
    .Q(\i_game_and_vga.i_game_top.end_of_game_timer_start ));
 sg13g2_dfrbp_1 _2430_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net348),
    .D(\i_game_and_vga.i_game_top.master_fsm.d_sprite_target_write_dxy ),
    .Q_N(_0015_),
    .Q(\i_game_and_vga.i_game_top.master_fsm.sprite_target_write_dxy ));
 sg13g2_dfrbp_1 _2431_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net346),
    .D(_0198_),
    .Q_N(_0032_),
    .Q(\i_game_and_vga.i_game_top.master_fsm.state[0] ));
 sg13g2_dfrbp_1 _2432_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net346),
    .D(_0199_),
    .Q_N(_0987_),
    .Q(\i_game_and_vga.i_game_top.master_fsm.state[1] ));
 sg13g2_dfrbp_1 _2433_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net21),
    .D(_0200_),
    .Q_N(_0986_),
    .Q(\i_game_and_vga.i_game_top.mixer.sprite_torpedo_rgb[2] ));
 sg13g2_dfrbp_1 _2434_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net44),
    .D(_0201_),
    .Q_N(_0016_),
    .Q(\i_game_and_vga.i_game_top.mixer.sprite_torpedo_rgb[1] ));
 sg13g2_dfrbp_1 _2435_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net31),
    .D(_0202_),
    .Q_N(_0985_),
    .Q(\i_game_and_vga.i_game_top.mixer.sprite_target_rgb[2] ));
 sg13g2_tiehi _2412__20 (.L_HI(net20));
 sg13g2_tiehi _2433__21 (.L_HI(net21));
 sg13g2_tiehi _2411__22 (.L_HI(net22));
 sg13g2_tiehi _2420__23 (.L_HI(net23));
 sg13g2_tiehi _2410__24 (.L_HI(net24));
 sg13g2_tiehi _2409__25 (.L_HI(net25));
 sg13g2_tiehi _2419__26 (.L_HI(net26));
 sg13g2_tiehi _2408__27 (.L_HI(net27));
 sg13g2_tiehi _2407__28 (.L_HI(net28));
 sg13g2_tiehi _2418__29 (.L_HI(net29));
 sg13g2_tiehi _2406__30 (.L_HI(net30));
 sg13g2_tiehi _2435__31 (.L_HI(net31));
 sg13g2_tiehi _2405__32 (.L_HI(net32));
 sg13g2_tiehi _2417__33 (.L_HI(net33));
 sg13g2_tiehi _2404__34 (.L_HI(net34));
 sg13g2_tiehi _2403__35 (.L_HI(net35));
 sg13g2_tiehi _2416__36 (.L_HI(net36));
 sg13g2_tiehi _2402__37 (.L_HI(net37));
 sg13g2_tiehi _2401__38 (.L_HI(net38));
 sg13g2_tiehi _2415__39 (.L_HI(net39));
 sg13g2_tiehi _2400__40 (.L_HI(net40));
 sg13g2_tiehi _2422__41 (.L_HI(net41));
 sg13g2_tiehi _2399__42 (.L_HI(net42));
 sg13g2_tiehi _2414__43 (.L_HI(net43));
 sg13g2_tiehi _2434__44 (.L_HI(net44));
 sg13g2_tiehi _2413__45 (.L_HI(net45));
 sg13g2_tiehi _2372__46 (.L_HI(net46));
 sg13g2_tiehi _2371__47 (.L_HI(net47));
 sg13g2_tiehi _2423__48 (.L_HI(net48));
 sg13g2_buf_2 clkbuf_leaf_0_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_tielo tt_um_yuri_panchul_sea_battle_vga_game_4 (.L_LO(net4));
 sg13g2_tielo tt_um_yuri_panchul_sea_battle_vga_game_5 (.L_LO(net5));
 sg13g2_tielo tt_um_yuri_panchul_sea_battle_vga_game_6 (.L_LO(net6));
 sg13g2_tielo tt_um_yuri_panchul_sea_battle_vga_game_7 (.L_LO(net7));
 sg13g2_tielo tt_um_yuri_panchul_sea_battle_vga_game_8 (.L_LO(net8));
 sg13g2_tielo tt_um_yuri_panchul_sea_battle_vga_game_9 (.L_LO(net9));
 sg13g2_tielo tt_um_yuri_panchul_sea_battle_vga_game_10 (.L_LO(net10));
 sg13g2_tielo tt_um_yuri_panchul_sea_battle_vga_game_11 (.L_LO(net11));
 sg13g2_tielo tt_um_yuri_panchul_sea_battle_vga_game_12 (.L_LO(net12));
 sg13g2_tielo tt_um_yuri_panchul_sea_battle_vga_game_13 (.L_LO(net13));
 sg13g2_tielo tt_um_yuri_panchul_sea_battle_vga_game_14 (.L_LO(net14));
 sg13g2_tielo tt_um_yuri_panchul_sea_battle_vga_game_15 (.L_LO(net15));
 sg13g2_tielo tt_um_yuri_panchul_sea_battle_vga_game_16 (.L_LO(net16));
 sg13g2_tielo tt_um_yuri_panchul_sea_battle_vga_game_17 (.L_LO(net17));
 sg13g2_tielo tt_um_yuri_panchul_sea_battle_vga_game_18 (.L_LO(net18));
 sg13g2_tiehi _2421__19 (.L_HI(net19));
 sg13g2_buf_1 _2482_ (.A(uo_out[4]),
    .X(uo_out[0]));
 sg13g2_buf_1 _2483_ (.A(uo_out[5]),
    .X(uo_out[1]));
 sg13g2_buf_1 _2484_ (.A(uo_out[6]),
    .X(uo_out[2]));
 sg13g2_buf_2 _2485_ (.A(\i_game_and_vga.i_vga.vsync ),
    .X(uo_out[3]));
 sg13g2_buf_2 _2486_ (.A(hsync),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout267 (.A(net268),
    .X(net267));
 sg13g2_buf_2 fanout268 (.A(_0218_),
    .X(net268));
 sg13g2_buf_2 fanout269 (.A(net270),
    .X(net269));
 sg13g2_buf_2 fanout270 (.A(_0479_),
    .X(net270));
 sg13g2_buf_2 fanout271 (.A(_0476_),
    .X(net271));
 sg13g2_buf_4 fanout272 (.X(net272),
    .A(net274));
 sg13g2_buf_4 fanout273 (.X(net273),
    .A(net274));
 sg13g2_buf_2 fanout274 (.A(_0364_),
    .X(net274));
 sg13g2_buf_2 fanout275 (.A(_0305_),
    .X(net275));
 sg13g2_buf_1 fanout276 (.A(_0305_),
    .X(net276));
 sg13g2_buf_4 fanout277 (.X(net277),
    .A(net278));
 sg13g2_buf_4 fanout278 (.X(net278),
    .A(net279));
 sg13g2_buf_2 fanout279 (.A(net130),
    .X(net279));
 sg13g2_buf_2 fanout280 (.A(net282),
    .X(net280));
 sg13g2_buf_2 fanout281 (.A(net282),
    .X(net281));
 sg13g2_buf_4 fanout282 (.X(net282),
    .A(net394));
 sg13g2_buf_2 fanout283 (.A(net395),
    .X(net283));
 sg13g2_buf_4 fanout284 (.X(net284),
    .A(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.dy[1] ));
 sg13g2_buf_4 fanout285 (.X(net285),
    .A(net193));
 sg13g2_buf_4 fanout286 (.X(net286),
    .A(net240));
 sg13g2_buf_2 fanout287 (.A(net242),
    .X(net287));
 sg13g2_buf_4 fanout288 (.X(net288),
    .A(net241));
 sg13g2_buf_2 fanout289 (.A(net355),
    .X(net289));
 sg13g2_buf_2 fanout290 (.A(net356),
    .X(net290));
 sg13g2_buf_2 fanout291 (.A(net257),
    .X(net291));
 sg13g2_buf_2 fanout292 (.A(net293),
    .X(net292));
 sg13g2_buf_2 fanout293 (.A(net137),
    .X(net293));
 sg13g2_buf_4 fanout294 (.X(net294),
    .A(net94));
 sg13g2_buf_2 fanout295 (.A(net296),
    .X(net295));
 sg13g2_buf_2 fanout296 (.A(net297),
    .X(net296));
 sg13g2_buf_2 fanout297 (.A(net371),
    .X(net297));
 sg13g2_buf_4 fanout298 (.X(net298),
    .A(net216));
 sg13g2_buf_2 fanout299 (.A(net208),
    .X(net299));
 sg13g2_buf_2 fanout300 (.A(net258),
    .X(net300));
 sg13g2_buf_2 fanout301 (.A(net246),
    .X(net301));
 sg13g2_buf_2 fanout302 (.A(net379),
    .X(net302));
 sg13g2_buf_2 fanout303 (.A(net135),
    .X(net303));
 sg13g2_buf_2 fanout304 (.A(net414),
    .X(net304));
 sg13g2_buf_2 fanout305 (.A(net306),
    .X(net305));
 sg13g2_buf_2 fanout306 (.A(net307),
    .X(net306));
 sg13g2_buf_4 fanout307 (.X(net307),
    .A(net309));
 sg13g2_buf_2 fanout308 (.A(net309),
    .X(net308));
 sg13g2_buf_4 fanout309 (.X(net309),
    .A(net372));
 sg13g2_buf_4 fanout310 (.X(net310),
    .A(net83));
 sg13g2_buf_2 fanout311 (.A(net408),
    .X(net311));
 sg13g2_buf_2 fanout312 (.A(net410),
    .X(net312));
 sg13g2_buf_2 fanout313 (.A(\i_game_and_vga.i_game_top.sprite_target.pixel_y[1] ),
    .X(net313));
 sg13g2_buf_4 fanout314 (.X(net314),
    .A(net325));
 sg13g2_buf_4 fanout315 (.X(net315),
    .A(net325));
 sg13g2_buf_4 fanout316 (.X(net316),
    .A(net318));
 sg13g2_buf_4 fanout317 (.X(net317),
    .A(net318));
 sg13g2_buf_2 fanout318 (.A(net325),
    .X(net318));
 sg13g2_buf_4 fanout319 (.X(net319),
    .A(net324));
 sg13g2_buf_2 fanout320 (.A(net324),
    .X(net320));
 sg13g2_buf_4 fanout321 (.X(net321),
    .A(net324));
 sg13g2_buf_4 fanout322 (.X(net322),
    .A(net324));
 sg13g2_buf_4 fanout323 (.X(net323),
    .A(net324));
 sg13g2_buf_2 fanout324 (.A(net325),
    .X(net324));
 sg13g2_buf_2 fanout325 (.A(net353),
    .X(net325));
 sg13g2_buf_4 fanout326 (.X(net326),
    .A(net327));
 sg13g2_buf_2 fanout327 (.A(net328),
    .X(net327));
 sg13g2_buf_4 fanout328 (.X(net328),
    .A(net329));
 sg13g2_buf_2 fanout329 (.A(net333),
    .X(net329));
 sg13g2_buf_4 fanout330 (.X(net330),
    .A(net331));
 sg13g2_buf_4 fanout331 (.X(net331),
    .A(net333));
 sg13g2_buf_4 fanout332 (.X(net332),
    .A(net333));
 sg13g2_buf_2 fanout333 (.A(net353),
    .X(net333));
 sg13g2_buf_4 fanout334 (.X(net334),
    .A(net336));
 sg13g2_buf_2 fanout335 (.A(net336),
    .X(net335));
 sg13g2_buf_2 fanout336 (.A(net341),
    .X(net336));
 sg13g2_buf_4 fanout337 (.X(net337),
    .A(net341));
 sg13g2_buf_2 fanout338 (.A(net341),
    .X(net338));
 sg13g2_buf_4 fanout339 (.X(net339),
    .A(net341));
 sg13g2_buf_2 fanout340 (.A(net341),
    .X(net340));
 sg13g2_buf_2 fanout341 (.A(net353),
    .X(net341));
 sg13g2_buf_4 fanout342 (.X(net342),
    .A(net352));
 sg13g2_buf_2 fanout343 (.A(net352),
    .X(net343));
 sg13g2_buf_4 fanout344 (.X(net344),
    .A(net345));
 sg13g2_buf_4 fanout345 (.X(net345),
    .A(net352));
 sg13g2_buf_4 fanout346 (.X(net346),
    .A(net348));
 sg13g2_buf_2 fanout347 (.A(net348),
    .X(net347));
 sg13g2_buf_4 fanout348 (.X(net348),
    .A(net352));
 sg13g2_buf_4 fanout349 (.X(net349),
    .A(net351));
 sg13g2_buf_4 fanout350 (.X(net350),
    .A(net351));
 sg13g2_buf_2 fanout351 (.A(net352),
    .X(net351));
 sg13g2_buf_2 fanout352 (.A(net353),
    .X(net352));
 sg13g2_buf_4 fanout353 (.X(net353),
    .A(rst_n));
 sg13g2_buf_2 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_2 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_tielo tt_um_yuri_panchul_sea_battle_vga_game_3 (.L_LO(net3));
 sg13g2_buf_2 clkbuf_leaf_1_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_2 clkbuf_leaf_2_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_2 clkbuf_leaf_3_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_2 clkbuf_leaf_4_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_2 clkbuf_leaf_5_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_2 clkbuf_leaf_6_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_2 clkbuf_leaf_7_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_2 clkbuf_leaf_8_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_2 clkbuf_leaf_9_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_2 clkbuf_leaf_10_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_2 clkbuf_leaf_11_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_2 clkbuf_leaf_12_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_2 clkbuf_leaf_13_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_2 clkbuf_leaf_14_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_2 clkbuf_leaf_15_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_2 clkbuf_leaf_16_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_2 clkbuf_leaf_17_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_2 clkbuf_leaf_18_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_2 clkbuf_leaf_19_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_2 clkbuf_leaf_20_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_2 clkbuf_leaf_21_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_2 clkbuf_leaf_22_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_2 clkbuf_leaf_23_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_2 clkbuf_leaf_24_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_2 clkbuf_leaf_25_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_2 clkbuf_leaf_26_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_2 clkbuf_leaf_27_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_2 clkbuf_leaf_28_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_2 clkbuf_leaf_29_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_2 clkbuf_leaf_30_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_2 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sg13g2_buf_2 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sg13g2_buf_2 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sg13g2_buf_2 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sg13g2_buf_2 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sg13g2_buf_2 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sg13g2_buf_2 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sg13g2_buf_2 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sg13g2_buf_2 clkload0 (.A(clknet_3_7__leaf_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_leaf_8_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_leaf_20_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_leaf_14_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(_1074_),
    .X(net49));
 sg13g2_dlygate4sd3_1 hold2 (.A(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_display.x_sprite_plus_w_1[0] ),
    .X(net50));
 sg13g2_dlygate4sd3_1 hold3 (.A(_0983_),
    .X(net51));
 sg13g2_dlygate4sd3_1 hold4 (.A(\i_game_and_vga.i_game_top.sprite_target.sprite_display.y_sprite_plus_h_1[0] ),
    .X(net52));
 sg13g2_dlygate4sd3_1 hold5 (.A(_0984_),
    .X(net53));
 sg13g2_dlygate4sd3_1 hold6 (.A(\i_game_and_vga.i_game_top.sprite_target.sprite_display.x_sprite_plus_w_1[0] ),
    .X(net54));
 sg13g2_dlygate4sd3_1 hold7 (.A(\i_game_and_vga.i_game_top.random[3] ),
    .X(net55));
 sg13g2_dlygate4sd3_1 hold8 (.A(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_display.y_sprite_plus_h_1[0] ),
    .X(net56));
 sg13g2_dlygate4sd3_1 hold9 (.A(\i_game_and_vga.i_game_top.random[9] ),
    .X(net57));
 sg13g2_dlygate4sd3_1 hold10 (.A(\i_game_and_vga.i_game_top.random[8] ),
    .X(net58));
 sg13g2_dlygate4sd3_1 hold11 (.A(\i_game_and_vga.i_game_top.random[13] ),
    .X(net59));
 sg13g2_dlygate4sd3_1 hold12 (.A(\i_game_and_vga.i_game_top.random[1] ),
    .X(net60));
 sg13g2_dlygate4sd3_1 hold13 (.A(\i_game_and_vga.i_game_top.random[10] ),
    .X(net61));
 sg13g2_dlygate4sd3_1 hold14 (.A(\i_game_and_vga.i_game_top.random[12] ),
    .X(net62));
 sg13g2_dlygate4sd3_1 hold15 (.A(\i_game_and_vga.i_game_top.random[6] ),
    .X(net63));
 sg13g2_dlygate4sd3_1 hold16 (.A(\i_game_and_vga.i_game_top.random[11] ),
    .X(net64));
 sg13g2_dlygate4sd3_1 hold17 (.A(_0098_),
    .X(net65));
 sg13g2_dlygate4sd3_1 hold18 (.A(\i_game_and_vga.i_game_top.sprite_target.sprite_control.sprite_y[6] ),
    .X(net66));
 sg13g2_dlygate4sd3_1 hold19 (.A(\i_game_and_vga.i_game_top.random[7] ),
    .X(net67));
 sg13g2_dlygate4sd3_1 hold20 (.A(\i_game_and_vga.i_game_top.sprite_target.sprite_control.sprite_y[3] ),
    .X(net68));
 sg13g2_dlygate4sd3_1 hold21 (.A(_0263_),
    .X(net69));
 sg13g2_dlygate4sd3_1 hold22 (.A(_0118_),
    .X(net70));
 sg13g2_dlygate4sd3_1 hold23 (.A(\i_game_and_vga.i_game_top.random[2] ),
    .X(net71));
 sg13g2_dlygate4sd3_1 hold24 (.A(_0089_),
    .X(net72));
 sg13g2_dlygate4sd3_1 hold25 (.A(\i_game_and_vga.i_game_top.random[5] ),
    .X(net73));
 sg13g2_dlygate4sd3_1 hold26 (.A(_0067_),
    .X(net74));
 sg13g2_dlygate4sd3_1 hold27 (.A(_0478_),
    .X(net75));
 sg13g2_dlygate4sd3_1 hold28 (.A(_0032_),
    .X(net76));
 sg13g2_dlygate4sd3_1 hold29 (.A(_0145_),
    .X(net77));
 sg13g2_dlygate4sd3_1 hold30 (.A(\i_game_and_vga.i_game_top.sprite_target.sprite_control.sprite_y[4] ),
    .X(net78));
 sg13g2_dlygate4sd3_1 hold31 (.A(\i_game_and_vga.i_game_top.sprite_target.sprite_control.sprite_y[5] ),
    .X(net79));
 sg13g2_dlygate4sd3_1 hold32 (.A(\i_game_and_vga.i_game_top.sprite_target.sprite_control.sprite_y[2] ),
    .X(net80));
 sg13g2_dlygate4sd3_1 hold33 (.A(\i_game_and_vga.i_game_top.random[14] ),
    .X(net81));
 sg13g2_dlygate4sd3_1 hold34 (.A(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.sprite_y[8] ),
    .X(net82));
 sg13g2_dlygate4sd3_1 hold35 (.A(\i_game_and_vga.i_game_top.sprite_target.sprite_control.sprite_y[1] ),
    .X(net83));
 sg13g2_dlygate4sd3_1 hold36 (.A(_0262_),
    .X(net84));
 sg13g2_dlygate4sd3_1 hold37 (.A(_0116_),
    .X(net85));
 sg13g2_dlygate4sd3_1 hold38 (.A(\i_game_and_vga.display_on ),
    .X(net86));
 sg13g2_dlygate4sd3_1 hold39 (.A(_0735_),
    .X(net87));
 sg13g2_dlygate4sd3_1 hold40 (.A(_0000_),
    .X(net88));
 sg13g2_dlygate4sd3_1 hold41 (.A(\i_game_and_vga.i_game_top.sprite_target.sprite_control.sprite_x[2] ),
    .X(net89));
 sg13g2_dlygate4sd3_1 hold42 (.A(\i_game_and_vga.i_game_top.sprite_target.sprite_control.dx[0] ),
    .X(net90));
 sg13g2_dlygate4sd3_1 hold43 (.A(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.sprite_x[9] ),
    .X(net91));
 sg13g2_dlygate4sd3_1 hold44 (.A(\i_game_and_vga.i_vga.clk_en_cnt[2] ),
    .X(net92));
 sg13g2_dlygate4sd3_1 hold45 (.A(_0010_),
    .X(net93));
 sg13g2_dlygate4sd3_1 hold46 (.A(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.sprite_y[0] ),
    .X(net94));
 sg13g2_dlygate4sd3_1 hold47 (.A(_0368_),
    .X(net95));
 sg13g2_dlygate4sd3_1 hold48 (.A(_0148_),
    .X(net96));
 sg13g2_dlygate4sd3_1 hold49 (.A(\i_game_and_vga.i_game_top.sprite_target.sprite_control.sprite_x[6] ),
    .X(net97));
 sg13g2_dlygate4sd3_1 hold50 (.A(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.sprite_y[6] ),
    .X(net98));
 sg13g2_dlygate4sd3_1 hold51 (.A(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.strobe_generator.counter[18] ),
    .X(net99));
 sg13g2_dlygate4sd3_1 hold52 (.A(_0206_),
    .X(net100));
 sg13g2_dlygate4sd3_1 hold53 (.A(_0060_),
    .X(net101));
 sg13g2_dlygate4sd3_1 hold54 (.A(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.sprite_y[5] ),
    .X(net102));
 sg13g2_dlygate4sd3_1 hold55 (.A(\i_game_and_vga.i_game_top.sprite_target.sprite_control.strobe_generator.counter[18] ),
    .X(net103));
 sg13g2_dlygate4sd3_1 hold56 (.A(_0210_),
    .X(net104));
 sg13g2_dlygate4sd3_1 hold57 (.A(_0045_),
    .X(net105));
 sg13g2_dlygate4sd3_1 hold58 (.A(\i_game_and_vga.i_game_top.sprite_target.sprite_control.sprite_y[3] ),
    .X(net106));
 sg13g2_dlygate4sd3_1 hold59 (.A(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.strobe_generator.strobe ),
    .X(net107));
 sg13g2_dlygate4sd3_1 hold60 (.A(_0158_),
    .X(net108));
 sg13g2_dlygate4sd3_1 hold61 (.A(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.strobe_generator.counter[17] ),
    .X(net109));
 sg13g2_dlygate4sd3_1 hold62 (.A(_0006_),
    .X(net110));
 sg13g2_dlygate4sd3_1 hold63 (.A(\i_game_and_vga.i_game_top.sprite_target.sprite_control.strobe_generator.counter[17] ),
    .X(net111));
 sg13g2_dlygate4sd3_1 hold64 (.A(_0004_),
    .X(net112));
 sg13g2_dlygate4sd3_1 hold65 (.A(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.sprite_x[8] ),
    .X(net113));
 sg13g2_dlygate4sd3_1 hold66 (.A(\i_game_and_vga.i_game_top.sprite_target.sprite_control.strobe_generator.counter[10] ),
    .X(net114));
 sg13g2_dlygate4sd3_1 hold67 (.A(_0037_),
    .X(net115));
 sg13g2_dlygate4sd3_1 hold68 (.A(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.strobe_generator.counter[1] ),
    .X(net116));
 sg13g2_dlygate4sd3_1 hold69 (.A(_0102_),
    .X(net117));
 sg13g2_dlygate4sd3_1 hold70 (.A(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.strobe_generator.counter[16] ),
    .X(net118));
 sg13g2_dlygate4sd3_1 hold71 (.A(_0058_),
    .X(net119));
 sg13g2_dlygate4sd3_1 hold72 (.A(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.strobe_generator.counter[3] ),
    .X(net120));
 sg13g2_dlygate4sd3_1 hold73 (.A(_0061_),
    .X(net121));
 sg13g2_dlygate4sd3_1 hold74 (.A(\i_game_and_vga.i_game_top.sprite_target.sprite_control.strobe_generator.counter[13] ),
    .X(net122));
 sg13g2_dlygate4sd3_1 hold75 (.A(_0040_),
    .X(net123));
 sg13g2_dlygate4sd3_1 hold76 (.A(\i_game_and_vga.i_game_top.sprite_target.sprite_control.strobe_generator.counter[16] ),
    .X(net124));
 sg13g2_dlygate4sd3_1 hold77 (.A(_0043_),
    .X(net125));
 sg13g2_dlygate4sd3_1 hold78 (.A(\i_game_and_vga.i_game_top.sprite_target.sprite_control.strobe_generator.counter[3] ),
    .X(net126));
 sg13g2_dlygate4sd3_1 hold79 (.A(_0046_),
    .X(net127));
 sg13g2_dlygate4sd3_1 hold80 (.A(\i_game_and_vga.i_game_top.sprite_target.sprite_control.strobe_generator.counter[6] ),
    .X(net128));
 sg13g2_dlygate4sd3_1 hold81 (.A(_0048_),
    .X(net129));
 sg13g2_dlygate4sd3_1 hold82 (.A(\i_game_and_vga.i_game_top.master_fsm.sprite_target_write_dxy ),
    .X(net130));
 sg13g2_dlygate4sd3_1 hold83 (.A(\i_game_and_vga.i_game_top.sprite_target.sprite_control.strobe_generator.counter[7] ),
    .X(net131));
 sg13g2_dlygate4sd3_1 hold84 (.A(_0049_),
    .X(net132));
 sg13g2_dlygate4sd3_1 hold85 (.A(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.strobe_generator.counter[6] ),
    .X(net133));
 sg13g2_dlygate4sd3_1 hold86 (.A(_0063_),
    .X(net134));
 sg13g2_dlygate4sd3_1 hold87 (.A(\i_game_and_vga.i_game_top.sprite_target.sprite_control.sprite_x[0] ),
    .X(net135));
 sg13g2_dlygate4sd3_1 hold88 (.A(\i_game_and_vga.i_game_top.sprite_target.sprite_display.x_sprite_plus_w_1[1] ),
    .X(net136));
 sg13g2_dlygate4sd3_1 hold89 (.A(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.sprite_y[1] ),
    .X(net137));
 sg13g2_dlygate4sd3_1 hold90 (.A(\i_game_and_vga.i_game_top.sprite_target.sprite_control.strobe_generator.counter[2] ),
    .X(net138));
 sg13g2_dlygate4sd3_1 hold91 (.A(_0630_),
    .X(net139));
 sg13g2_dlygate4sd3_1 hold92 (.A(_0100_),
    .X(net140));
 sg13g2_dlygate4sd3_1 hold93 (.A(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.strobe_generator.counter[13] ),
    .X(net141));
 sg13g2_dlygate4sd3_1 hold94 (.A(_0055_),
    .X(net142));
 sg13g2_dlygate4sd3_1 hold95 (.A(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.strobe_generator.counter[15] ),
    .X(net143));
 sg13g2_dlygate4sd3_1 hold96 (.A(_0652_),
    .X(net144));
 sg13g2_dlygate4sd3_1 hold97 (.A(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.strobe_generator.counter[7] ),
    .X(net145));
 sg13g2_dlygate4sd3_1 hold98 (.A(_0064_),
    .X(net146));
 sg13g2_dlygate4sd3_1 hold99 (.A(\i_game_and_vga.i_game_top.sprite_target.sprite_control.strobe_generator.counter[1] ),
    .X(net147));
 sg13g2_dlygate4sd3_1 hold100 (.A(_0099_),
    .X(net148));
 sg13g2_dlygate4sd3_1 hold101 (.A(\i_game_and_vga.i_game_top.timer.counter[24] ),
    .X(net149));
 sg13g2_dlygate4sd3_1 hold102 (.A(_0197_),
    .X(net150));
 sg13g2_dlygate4sd3_1 hold103 (.A(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.sprite_x[7] ),
    .X(net151));
 sg13g2_dlygate4sd3_1 hold104 (.A(\i_game_and_vga.i_game_top.timer.counter[21] ),
    .X(net152));
 sg13g2_dlygate4sd3_1 hold105 (.A(_0194_),
    .X(net153));
 sg13g2_dlygate4sd3_1 hold106 (.A(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.sprite_x[6] ),
    .X(net154));
 sg13g2_dlygate4sd3_1 hold107 (.A(\i_game_and_vga.i_vga.clk_en_cnt[3] ),
    .X(net155));
 sg13g2_dlygate4sd3_1 hold108 (.A(_0014_),
    .X(net156));
 sg13g2_dlygate4sd3_1 hold109 (.A(\i_game_and_vga.i_game_top.sprite_target.sprite_control.sprite_y[0] ),
    .X(net157));
 sg13g2_dlygate4sd3_1 hold110 (.A(\i_game_and_vga.i_game_top.sprite_target.sprite_control.strobe_generator.counter[14] ),
    .X(net158));
 sg13g2_dlygate4sd3_1 hold111 (.A(_0041_),
    .X(net159));
 sg13g2_dlygate4sd3_1 hold112 (.A(\i_game_and_vga.i_game_top.timer.counter[23] ),
    .X(net160));
 sg13g2_dlygate4sd3_1 hold113 (.A(_0196_),
    .X(net161));
 sg13g2_dlygate4sd3_1 hold114 (.A(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.strobe_generator.counter[10] ),
    .X(net162));
 sg13g2_dlygate4sd3_1 hold115 (.A(_0052_),
    .X(net163));
 sg13g2_dlygate4sd3_1 hold116 (.A(\i_game_and_vga.i_game_top.timer.counter[15] ),
    .X(net164));
 sg13g2_dlygate4sd3_1 hold117 (.A(_0188_),
    .X(net165));
 sg13g2_dlygate4sd3_1 hold118 (.A(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.sprite_x[4] ),
    .X(net166));
 sg13g2_dlygate4sd3_1 hold119 (.A(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.dx[0] ),
    .X(net167));
 sg13g2_dlygate4sd3_1 hold120 (.A(_0415_),
    .X(net168));
 sg13g2_dlygate4sd3_1 hold121 (.A(_0157_),
    .X(net169));
 sg13g2_dlygate4sd3_1 hold122 (.A(\i_game_and_vga.i_game_top.sprite_target.sprite_control.strobe_generator.counter[11] ),
    .X(net170));
 sg13g2_dlygate4sd3_1 hold123 (.A(_0038_),
    .X(net171));
 sg13g2_dlygate4sd3_1 hold124 (.A(\i_game_and_vga.i_game_top.sprite_target.sprite_control.strobe_generator.counter[5] ),
    .X(net172));
 sg13g2_dlygate4sd3_1 hold125 (.A(_0632_),
    .X(net173));
 sg13g2_dlygate4sd3_1 hold126 (.A(_0101_),
    .X(net174));
 sg13g2_dlygate4sd3_1 hold127 (.A(\i_game_and_vga.i_game_top.timer.counter[3] ),
    .X(net175));
 sg13g2_dlygate4sd3_1 hold128 (.A(_0176_),
    .X(net176));
 sg13g2_dlygate4sd3_1 hold129 (.A(\i_game_and_vga.i_game_top.mixer.sprite_torpedo_rgb[1] ),
    .X(net177));
 sg13g2_dlygate4sd3_1 hold130 (.A(\i_game_and_vga.i_game_top.mixer.sprite_target_rgb[2] ),
    .X(net178));
 sg13g2_dlygate4sd3_1 hold131 (.A(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.strobe_generator.counter[14] ),
    .X(net179));
 sg13g2_dlygate4sd3_1 hold132 (.A(_0056_),
    .X(net180));
 sg13g2_dlygate4sd3_1 hold133 (.A(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.sprite_y[7] ),
    .X(net181));
 sg13g2_dlygate4sd3_1 hold134 (.A(\i_game_and_vga.i_game_top.random[4] ),
    .X(net182));
 sg13g2_dlygate4sd3_1 hold135 (.A(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.strobe_generator.counter[11] ),
    .X(net183));
 sg13g2_dlygate4sd3_1 hold136 (.A(_0053_),
    .X(net184));
 sg13g2_dlygate4sd3_1 hold137 (.A(_0026_),
    .X(net185));
 sg13g2_dlygate4sd3_1 hold138 (.A(\i_game_and_vga.i_vga.clk_en_cnt[0] ),
    .X(net186));
 sg13g2_dlygate4sd3_1 hold139 (.A(\i_game_and_vga.i_game_top.mixer.sprite_target_rgb[0] ),
    .X(net187));
 sg13g2_dlygate4sd3_1 hold140 (.A(\i_game_and_vga.i_game_top.sprite_target.sprite_control.strobe_generator.counter[15] ),
    .X(net188));
 sg13g2_dlygate4sd3_1 hold141 (.A(\i_game_and_vga.i_vga.vpos[9] ),
    .X(net189));
 sg13g2_dlygate4sd3_1 hold142 (.A(\i_game_and_vga.i_game_top.timer.counter[22] ),
    .X(net190));
 sg13g2_dlygate4sd3_1 hold143 (.A(_0524_),
    .X(net191));
 sg13g2_dlygate4sd3_1 hold144 (.A(\i_game_and_vga.i_game_top.sprite_target.sprite_control.sprite_x[7] ),
    .X(net192));
 sg13g2_dlygate4sd3_1 hold145 (.A(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.sprite_x[3] ),
    .X(net193));
 sg13g2_dlygate4sd3_1 hold146 (.A(\i_game_and_vga.i_game_top.sprite_target.pixel_y[1] ),
    .X(net194));
 sg13g2_dlygate4sd3_1 hold147 (.A(_0106_),
    .X(net195));
 sg13g2_dlygate4sd3_1 hold148 (.A(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.strobe_generator.counter[8] ),
    .X(net196));
 sg13g2_dlygate4sd3_1 hold149 (.A(_0065_),
    .X(net197));
 sg13g2_dlygate4sd3_1 hold150 (.A(_0031_),
    .X(net198));
 sg13g2_dlygate4sd3_1 hold151 (.A(_0738_),
    .X(net199));
 sg13g2_dlygate4sd3_1 hold152 (.A(\i_game_and_vga.i_game_top.mixer.sprite_target_rgb[1] ),
    .X(net200));
 sg13g2_dlygate4sd3_1 hold153 (.A(\i_game_and_vga.i_game_top.timer.counter[12] ),
    .X(net201));
 sg13g2_dlygate4sd3_1 hold154 (.A(_0503_),
    .X(net202));
 sg13g2_dlygate4sd3_1 hold155 (.A(_0185_),
    .X(net203));
 sg13g2_dlygate4sd3_1 hold156 (.A(\i_game_and_vga.i_game_top.timer.counter[18] ),
    .X(net204));
 sg13g2_dlygate4sd3_1 hold157 (.A(\i_game_and_vga.i_game_top.timer.counter[19] ),
    .X(net205));
 sg13g2_dlygate4sd3_1 hold158 (.A(\i_game_and_vga.i_game_top.sprite_target.sprite_control.strobe_generator.counter[8] ),
    .X(net206));
 sg13g2_dlygate4sd3_1 hold159 (.A(_0050_),
    .X(net207));
 sg13g2_dlygate4sd3_1 hold160 (.A(\i_game_and_vga.i_game_top.sprite_target.sprite_control.sprite_x[8] ),
    .X(net208));
 sg13g2_dlygate4sd3_1 hold161 (.A(\i_game_and_vga.i_game_top.sprite_target.sprite_display.x_sprite_within_screen ),
    .X(net209));
 sg13g2_dlygate4sd3_1 hold162 (.A(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.strobe_generator.counter[5] ),
    .X(net210));
 sg13g2_dlygate4sd3_1 hold163 (.A(_0627_),
    .X(net211));
 sg13g2_dlygate4sd3_1 hold164 (.A(_0104_),
    .X(net212));
 sg13g2_dlygate4sd3_1 hold165 (.A(\i_game_and_vga.i_game_top.master_fsm.state[0] ),
    .X(net213));
 sg13g2_dlygate4sd3_1 hold166 (.A(\i_game_and_vga.i_game_top.master_fsm.d_sprite_torpedo_enable_update ),
    .X(net214));
 sg13g2_dlygate4sd3_1 hold167 (.A(_0033_),
    .X(net215));
 sg13g2_dlygate4sd3_1 hold168 (.A(\i_game_and_vga.i_game_top.sprite_target.sprite_control.sprite_x[9] ),
    .X(net216));
 sg13g2_dlygate4sd3_1 hold169 (.A(\i_game_and_vga.i_game_top.game_won ),
    .X(net217));
 sg13g2_dlygate4sd3_1 hold170 (.A(_0737_),
    .X(net218));
 sg13g2_dlygate4sd3_1 hold171 (.A(_0001_),
    .X(net219));
 sg13g2_dlygate4sd3_1 hold172 (.A(\i_game_and_vga.i_game_top.sprite_target.sprite_control.strobe_generator.counter[4] ),
    .X(net220));
 sg13g2_dlygate4sd3_1 hold173 (.A(_0047_),
    .X(net221));
 sg13g2_dlygate4sd3_1 hold174 (.A(\i_game_and_vga.i_game_top.sprite_target.sprite_control.sprite_x[5] ),
    .X(net222));
 sg13g2_dlygate4sd3_1 hold175 (.A(\i_game_and_vga.i_game_top.mixer.random ),
    .X(net223));
 sg13g2_dlygate4sd3_1 hold176 (.A(_0087_),
    .X(net224));
 sg13g2_dlygate4sd3_1 hold177 (.A(\i_game_and_vga.i_vga.clk_en_cnt[1] ),
    .X(net225));
 sg13g2_dlygate4sd3_1 hold178 (.A(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.strobe_generator.counter[2] ),
    .X(net226));
 sg13g2_dlygate4sd3_1 hold179 (.A(_0625_),
    .X(net227));
 sg13g2_dlygate4sd3_1 hold180 (.A(_0103_),
    .X(net228));
 sg13g2_dlygate4sd3_1 hold181 (.A(hsync),
    .X(net229));
 sg13g2_dlygate4sd3_1 hold182 (.A(_0291_),
    .X(net230));
 sg13g2_dlygate4sd3_1 hold183 (.A(\i_game_and_vga.i_game_top.overlap.top_2[8] ),
    .X(net231));
 sg13g2_dlygate4sd3_1 hold184 (.A(_0720_),
    .X(net232));
 sg13g2_dlygate4sd3_1 hold185 (.A(_0003_),
    .X(net233));
 sg13g2_dlygate4sd3_1 hold186 (.A(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.strobe_generator.counter[4] ),
    .X(net234));
 sg13g2_dlygate4sd3_1 hold187 (.A(_0062_),
    .X(net235));
 sg13g2_dlygate4sd3_1 hold188 (.A(\i_game_and_vga.i_vga.vsync ),
    .X(net236));
 sg13g2_dlygate4sd3_1 hold189 (.A(_0124_),
    .X(net237));
 sg13g2_dlygate4sd3_1 hold190 (.A(_0015_),
    .X(net238));
 sg13g2_dlygate4sd3_1 hold191 (.A(\i_game_and_vga.i_game_top.master_fsm.state[1] ),
    .X(net239));
 sg13g2_dlygate4sd3_1 hold192 (.A(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.sprite_x[2] ),
    .X(net240));
 sg13g2_dlygate4sd3_1 hold193 (.A(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.sprite_x[0] ),
    .X(net241));
 sg13g2_dlygate4sd3_1 hold194 (.A(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.sprite_x[1] ),
    .X(net242));
 sg13g2_dlygate4sd3_1 hold195 (.A(\i_game_and_vga.i_game_top.timer.counter[8] ),
    .X(net243));
 sg13g2_dlygate4sd3_1 hold196 (.A(_0496_),
    .X(net244));
 sg13g2_dlygate4sd3_1 hold197 (.A(_0181_),
    .X(net245));
 sg13g2_dlygate4sd3_1 hold198 (.A(\i_game_and_vga.i_game_top.sprite_target.sprite_control.sprite_x[3] ),
    .X(net246));
 sg13g2_dlygate4sd3_1 hold199 (.A(\i_game_and_vga.i_game_top.mixer.sprite_torpedo_rgb[2] ),
    .X(net247));
 sg13g2_dlygate4sd3_1 hold200 (.A(\i_game_and_vga.i_game_top.timer.counter[17] ),
    .X(net248));
 sg13g2_dlygate4sd3_1 hold201 (.A(_0512_),
    .X(net249));
 sg13g2_dlygate4sd3_1 hold202 (.A(_0190_),
    .X(net250));
 sg13g2_dlygate4sd3_1 hold203 (.A(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.sprite_x[5] ),
    .X(net251));
 sg13g2_dlygate4sd3_1 hold204 (.A(_0025_),
    .X(net252));
 sg13g2_dlygate4sd3_1 hold205 (.A(\i_game_and_vga.i_game_top.timer.counter[14] ),
    .X(net253));
 sg13g2_dlygate4sd3_1 hold206 (.A(_0508_),
    .X(net254));
 sg13g2_dlygate4sd3_1 hold207 (.A(\i_game_and_vga.i_game_top.timer.counter[6] ),
    .X(net255));
 sg13g2_dlygate4sd3_1 hold208 (.A(_0179_),
    .X(net256));
 sg13g2_dlygate4sd3_1 hold209 (.A(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.sprite_y[2] ),
    .X(net257));
 sg13g2_dlygate4sd3_1 hold210 (.A(\i_game_and_vga.i_game_top.sprite_target.sprite_control.sprite_x[4] ),
    .X(net258));
 sg13g2_dlygate4sd3_1 hold211 (.A(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.dy[0] ),
    .X(net259));
 sg13g2_dlygate4sd3_1 hold212 (.A(_0471_),
    .X(net260));
 sg13g2_dlygate4sd3_1 hold213 (.A(\i_game_and_vga.i_game_top.timer.counter[11] ),
    .X(net261));
 sg13g2_dlygate4sd3_1 hold214 (.A(_0502_),
    .X(net262));
 sg13g2_dlygate4sd3_1 hold215 (.A(\i_game_and_vga.i_game_top.timer.counter[2] ),
    .X(net263));
 sg13g2_dlygate4sd3_1 hold216 (.A(_0485_),
    .X(net264));
 sg13g2_dlygate4sd3_1 hold217 (.A(\i_game_and_vga.i_game_top.timer.counter[10] ),
    .X(net265));
 sg13g2_dlygate4sd3_1 hold218 (.A(_0499_),
    .X(net266));
 sg13g2_dlygate4sd3_1 hold219 (.A(_0183_),
    .X(net354));
 sg13g2_dlygate4sd3_1 hold220 (.A(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.sprite_y[4] ),
    .X(net355));
 sg13g2_dlygate4sd3_1 hold221 (.A(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.sprite_y[3] ),
    .X(net356));
 sg13g2_dlygate4sd3_1 hold222 (.A(\i_game_and_vga.i_game_top.timer.counter[5] ),
    .X(net357));
 sg13g2_dlygate4sd3_1 hold223 (.A(_0178_),
    .X(net358));
 sg13g2_dlygate4sd3_1 hold224 (.A(\i_game_and_vga.i_game_top.sprite_target.pixel_y[5] ),
    .X(net359));
 sg13g2_dlygate4sd3_1 hold225 (.A(_0110_),
    .X(net360));
 sg13g2_dlygate4sd3_1 hold226 (.A(\i_game_and_vga.i_game_top.timer.counter[4] ),
    .X(net361));
 sg13g2_dlygate4sd3_1 hold227 (.A(_0489_),
    .X(net362));
 sg13g2_dlygate4sd3_1 hold228 (.A(\i_game_and_vga.i_game_top.sprite_target.sprite_control.sprite_y[0] ),
    .X(net363));
 sg13g2_dlygate4sd3_1 hold229 (.A(\i_game_and_vga.i_game_top.timer.counter[20] ),
    .X(net364));
 sg13g2_dlygate4sd3_1 hold230 (.A(\i_game_and_vga.i_game_top.end_of_game_timer_running ),
    .X(net365));
 sg13g2_dlygate4sd3_1 hold231 (.A(_0009_),
    .X(net366));
 sg13g2_dlygate4sd3_1 hold232 (.A(\i_game_and_vga.i_game_top.sprite_target.pixel_x[4] ),
    .X(net367));
 sg13g2_dlygate4sd3_1 hold233 (.A(\i_game_and_vga.i_game_top.sprite_target.pixel_y[4] ),
    .X(net368));
 sg13g2_dlygate4sd3_1 hold234 (.A(\i_game_and_vga.i_game_top.timer.counter[16] ),
    .X(net369));
 sg13g2_dlygate4sd3_1 hold235 (.A(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.strobe_generator.counter[12] ),
    .X(net370));
 sg13g2_dlygate4sd3_1 hold236 (.A(\i_game_and_vga.i_game_top.sprite_target.sprite_control.dx[1] ),
    .X(net371));
 sg13g2_dlygate4sd3_1 hold237 (.A(\i_game_and_vga.i_vga.clk_en ),
    .X(net372));
 sg13g2_dlygate4sd3_1 hold238 (.A(\i_game_and_vga.i_game_top.sprite_target.pixel_x[2] ),
    .X(net373));
 sg13g2_dlygate4sd3_1 hold239 (.A(_0299_),
    .X(net374));
 sg13g2_dlygate4sd3_1 hold240 (.A(_0128_),
    .X(net375));
 sg13g2_dlygate4sd3_1 hold241 (.A(\i_game_and_vga.i_game_top.sprite_target.pixel_y[2] ),
    .X(net376));
 sg13g2_dlygate4sd3_1 hold242 (.A(\i_game_and_vga.i_game_top.sprite_target.sprite_control.strobe_generator.strobe ),
    .X(net377));
 sg13g2_dlygate4sd3_1 hold243 (.A(_0325_),
    .X(net378));
 sg13g2_dlygate4sd3_1 hold244 (.A(\i_game_and_vga.i_game_top.sprite_target.sprite_control.sprite_x[1] ),
    .X(net379));
 sg13g2_dlygate4sd3_1 hold245 (.A(\i_game_and_vga.i_game_top.sprite_target.sprite_control.strobe_generator.counter[12] ),
    .X(net380));
 sg13g2_dlygate4sd3_1 hold246 (.A(\i_game_and_vga.i_game_top.timer.counter[13] ),
    .X(net381));
 sg13g2_dlygate4sd3_1 hold247 (.A(\i_game_and_vga.i_game_top.master_fsm.sprite_torpedo_enable_update ),
    .X(net382));
 sg13g2_dlygate4sd3_1 hold248 (.A(\i_game_and_vga.i_game_top.sprite_target.pixel_x[6] ),
    .X(net383));
 sg13g2_dlygate4sd3_1 hold249 (.A(\i_game_and_vga.i_game_top.sprite_target.pixel_y[8] ),
    .X(net384));
 sg13g2_dlygate4sd3_1 hold250 (.A(\i_game_and_vga.i_game_top.sprite_target.pixel_x[5] ),
    .X(net385));
 sg13g2_dlygate4sd3_1 hold251 (.A(_0130_),
    .X(net386));
 sg13g2_dlygate4sd3_1 hold252 (.A(\i_game_and_vga.i_game_top.master_fsm.sprite_target_enable_update ),
    .X(net387));
 sg13g2_dlygate4sd3_1 hold253 (.A(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.strobe_generator.counter[9] ),
    .X(net388));
 sg13g2_dlygate4sd3_1 hold254 (.A(\i_game_and_vga.i_game_top.timer.counter[9] ),
    .X(net389));
 sg13g2_dlygate4sd3_1 hold255 (.A(\i_game_and_vga.i_game_top.timer.counter[7] ),
    .X(net390));
 sg13g2_dlygate4sd3_1 hold256 (.A(_0020_),
    .X(net391));
 sg13g2_dlygate4sd3_1 hold257 (.A(\i_game_and_vga.i_game_top.sprite_target.sprite_control.strobe_generator.counter[9] ),
    .X(net392));
 sg13g2_dlygate4sd3_1 hold258 (.A(\i_game_and_vga.i_game_top.sprite_target.pixel_x[0] ),
    .X(net393));
 sg13g2_dlygate4sd3_1 hold259 (.A(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.dx[1] ),
    .X(net394));
 sg13g2_dlygate4sd3_1 hold260 (.A(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.dy[1] ),
    .X(net395));
 sg13g2_dlygate4sd3_1 hold261 (.A(\i_game_and_vga.i_game_top.sprite_target.pixel_y[0] ),
    .X(net396));
 sg13g2_dlygate4sd3_1 hold262 (.A(\i_game_and_vga.i_game_top.sprite_target.pixel_x[1] ),
    .X(net397));
 sg13g2_dlygate4sd3_1 hold263 (.A(\i_game_and_vga.i_game_top.sprite_target.pixel_y[6] ),
    .X(net398));
 sg13g2_dlygate4sd3_1 hold264 (.A(_0111_),
    .X(net399));
 sg13g2_dlygate4sd3_1 hold265 (.A(\i_game_and_vga.i_game_top.timer.counter[1] ),
    .X(net400));
 sg13g2_dlygate4sd3_1 hold266 (.A(_0481_),
    .X(net401));
 sg13g2_dlygate4sd3_1 hold267 (.A(_0483_),
    .X(net402));
 sg13g2_dlygate4sd3_1 hold268 (.A(\i_game_and_vga.i_game_top.random[15] ),
    .X(net403));
 sg13g2_dlygate4sd3_1 hold269 (.A(\i_game_and_vga.i_game_top.sprite_target.pixel_x[7] ),
    .X(net404));
 sg13g2_dlygate4sd3_1 hold270 (.A(_0132_),
    .X(net405));
 sg13g2_dlygate4sd3_1 hold271 (.A(\i_game_and_vga.i_game_top.sprite_target.sprite_control.sprite_x[7] ),
    .X(net406));
 sg13g2_dlygate4sd3_1 hold272 (.A(_0024_),
    .X(net407));
 sg13g2_dlygate4sd3_1 hold273 (.A(\i_game_and_vga.i_game_top.sprite_target.pixel_y[7] ),
    .X(net408));
 sg13g2_dlygate4sd3_1 hold274 (.A(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.sprite_y[7] ),
    .X(net409));
 sg13g2_dlygate4sd3_1 hold275 (.A(\i_game_and_vga.i_game_top.sprite_target.pixel_y[3] ),
    .X(net410));
 sg13g2_dlygate4sd3_1 hold276 (.A(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.sprite_x[9] ),
    .X(net411));
 sg13g2_dlygate4sd3_1 hold277 (.A(\i_game_and_vga.i_game_top.sprite_target.pixel_x[8] ),
    .X(net412));
 sg13g2_dlygate4sd3_1 hold278 (.A(_0133_),
    .X(net413));
 sg13g2_dlygate4sd3_1 hold279 (.A(\i_game_and_vga.i_game_top.sprite_target.pixel_x[9] ),
    .X(net414));
 sg13g2_dlygate4sd3_1 hold280 (.A(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.strobe_generator.counter[14] ),
    .X(net415));
 sg13g2_dlygate4sd3_1 hold281 (.A(\i_game_and_vga.i_game_top.sprite_target.sprite_control.sprite_x[5] ),
    .X(net416));
 sg13g2_dlygate4sd3_1 hold282 (.A(\i_game_and_vga.i_game_top.sprite_torpedo.sprite_control.sprite_x[8] ),
    .X(net417));
 sg13g2_antennanp ANTENNA_1 (.A(clk));
 sg13g2_antennanp ANTENNA_2 (.A(clk));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_fill_2 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_4 FILLER_13_147 ();
 sg13g2_fill_2 FILLER_13_151 ();
 sg13g2_decap_4 FILLER_13_182 ();
 sg13g2_fill_1 FILLER_13_224 ();
 sg13g2_decap_4 FILLER_13_251 ();
 sg13g2_fill_2 FILLER_13_263 ();
 sg13g2_decap_8 FILLER_13_283 ();
 sg13g2_decap_8 FILLER_13_290 ();
 sg13g2_decap_8 FILLER_13_297 ();
 sg13g2_decap_8 FILLER_13_304 ();
 sg13g2_decap_8 FILLER_13_311 ();
 sg13g2_decap_8 FILLER_13_318 ();
 sg13g2_decap_8 FILLER_13_325 ();
 sg13g2_decap_8 FILLER_13_332 ();
 sg13g2_decap_8 FILLER_13_339 ();
 sg13g2_decap_8 FILLER_13_346 ();
 sg13g2_decap_8 FILLER_13_353 ();
 sg13g2_decap_8 FILLER_13_360 ();
 sg13g2_decap_8 FILLER_13_367 ();
 sg13g2_decap_8 FILLER_13_374 ();
 sg13g2_decap_8 FILLER_13_381 ();
 sg13g2_decap_8 FILLER_13_388 ();
 sg13g2_decap_8 FILLER_13_395 ();
 sg13g2_decap_8 FILLER_13_402 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_4 FILLER_14_140 ();
 sg13g2_fill_1 FILLER_14_144 ();
 sg13g2_fill_2 FILLER_14_156 ();
 sg13g2_decap_8 FILLER_14_293 ();
 sg13g2_decap_8 FILLER_14_300 ();
 sg13g2_decap_8 FILLER_14_307 ();
 sg13g2_decap_8 FILLER_14_314 ();
 sg13g2_decap_8 FILLER_14_321 ();
 sg13g2_decap_8 FILLER_14_328 ();
 sg13g2_decap_8 FILLER_14_335 ();
 sg13g2_decap_8 FILLER_14_342 ();
 sg13g2_decap_8 FILLER_14_349 ();
 sg13g2_decap_8 FILLER_14_356 ();
 sg13g2_decap_8 FILLER_14_363 ();
 sg13g2_decap_8 FILLER_14_370 ();
 sg13g2_decap_8 FILLER_14_377 ();
 sg13g2_decap_8 FILLER_14_384 ();
 sg13g2_decap_8 FILLER_14_391 ();
 sg13g2_decap_8 FILLER_14_398 ();
 sg13g2_decap_4 FILLER_14_405 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_fill_2 FILLER_15_174 ();
 sg13g2_fill_2 FILLER_15_202 ();
 sg13g2_fill_1 FILLER_15_204 ();
 sg13g2_fill_2 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_223 ();
 sg13g2_decap_8 FILLER_15_230 ();
 sg13g2_decap_8 FILLER_15_237 ();
 sg13g2_fill_1 FILLER_15_244 ();
 sg13g2_decap_8 FILLER_15_301 ();
 sg13g2_decap_8 FILLER_15_308 ();
 sg13g2_decap_8 FILLER_15_315 ();
 sg13g2_decap_8 FILLER_15_322 ();
 sg13g2_decap_8 FILLER_15_329 ();
 sg13g2_decap_8 FILLER_15_336 ();
 sg13g2_decap_8 FILLER_15_343 ();
 sg13g2_decap_8 FILLER_15_350 ();
 sg13g2_decap_8 FILLER_15_357 ();
 sg13g2_decap_8 FILLER_15_364 ();
 sg13g2_decap_8 FILLER_15_371 ();
 sg13g2_decap_8 FILLER_15_378 ();
 sg13g2_decap_8 FILLER_15_385 ();
 sg13g2_decap_8 FILLER_15_392 ();
 sg13g2_decap_8 FILLER_15_399 ();
 sg13g2_fill_2 FILLER_15_406 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_4 FILLER_16_126 ();
 sg13g2_fill_2 FILLER_16_130 ();
 sg13g2_decap_4 FILLER_16_185 ();
 sg13g2_fill_2 FILLER_16_221 ();
 sg13g2_fill_1 FILLER_16_223 ();
 sg13g2_fill_2 FILLER_16_228 ();
 sg13g2_decap_8 FILLER_16_239 ();
 sg13g2_decap_4 FILLER_16_246 ();
 sg13g2_fill_2 FILLER_16_250 ();
 sg13g2_fill_2 FILLER_16_278 ();
 sg13g2_fill_1 FILLER_16_280 ();
 sg13g2_decap_8 FILLER_16_292 ();
 sg13g2_decap_4 FILLER_16_299 ();
 sg13g2_decap_8 FILLER_16_308 ();
 sg13g2_decap_8 FILLER_16_315 ();
 sg13g2_decap_8 FILLER_16_322 ();
 sg13g2_decap_8 FILLER_16_329 ();
 sg13g2_decap_8 FILLER_16_336 ();
 sg13g2_decap_8 FILLER_16_343 ();
 sg13g2_decap_8 FILLER_16_350 ();
 sg13g2_decap_8 FILLER_16_357 ();
 sg13g2_decap_8 FILLER_16_364 ();
 sg13g2_decap_8 FILLER_16_371 ();
 sg13g2_decap_8 FILLER_16_378 ();
 sg13g2_decap_8 FILLER_16_385 ();
 sg13g2_decap_8 FILLER_16_392 ();
 sg13g2_decap_8 FILLER_16_399 ();
 sg13g2_fill_2 FILLER_16_406 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_4 FILLER_17_133 ();
 sg13g2_fill_2 FILLER_17_162 ();
 sg13g2_fill_1 FILLER_17_177 ();
 sg13g2_decap_4 FILLER_17_204 ();
 sg13g2_fill_2 FILLER_17_216 ();
 sg13g2_decap_4 FILLER_17_256 ();
 sg13g2_fill_1 FILLER_17_265 ();
 sg13g2_decap_4 FILLER_17_269 ();
 sg13g2_decap_8 FILLER_17_278 ();
 sg13g2_decap_8 FILLER_17_285 ();
 sg13g2_decap_8 FILLER_17_292 ();
 sg13g2_decap_8 FILLER_17_299 ();
 sg13g2_decap_8 FILLER_17_306 ();
 sg13g2_decap_8 FILLER_17_313 ();
 sg13g2_decap_8 FILLER_17_320 ();
 sg13g2_decap_8 FILLER_17_327 ();
 sg13g2_decap_8 FILLER_17_334 ();
 sg13g2_decap_8 FILLER_17_341 ();
 sg13g2_decap_8 FILLER_17_348 ();
 sg13g2_decap_8 FILLER_17_355 ();
 sg13g2_decap_8 FILLER_17_362 ();
 sg13g2_decap_8 FILLER_17_369 ();
 sg13g2_decap_8 FILLER_17_376 ();
 sg13g2_decap_8 FILLER_17_383 ();
 sg13g2_decap_8 FILLER_17_390 ();
 sg13g2_decap_8 FILLER_17_397 ();
 sg13g2_decap_4 FILLER_17_404 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_4 FILLER_18_105 ();
 sg13g2_fill_1 FILLER_18_109 ();
 sg13g2_decap_8 FILLER_18_128 ();
 sg13g2_decap_8 FILLER_18_135 ();
 sg13g2_decap_4 FILLER_18_142 ();
 sg13g2_fill_2 FILLER_18_161 ();
 sg13g2_decap_4 FILLER_18_168 ();
 sg13g2_decap_8 FILLER_18_198 ();
 sg13g2_fill_1 FILLER_18_205 ();
 sg13g2_fill_2 FILLER_18_226 ();
 sg13g2_decap_8 FILLER_18_249 ();
 sg13g2_decap_8 FILLER_18_256 ();
 sg13g2_decap_8 FILLER_18_294 ();
 sg13g2_decap_8 FILLER_18_301 ();
 sg13g2_decap_8 FILLER_18_308 ();
 sg13g2_decap_8 FILLER_18_315 ();
 sg13g2_decap_8 FILLER_18_322 ();
 sg13g2_decap_8 FILLER_18_329 ();
 sg13g2_decap_8 FILLER_18_336 ();
 sg13g2_decap_8 FILLER_18_343 ();
 sg13g2_decap_8 FILLER_18_350 ();
 sg13g2_decap_8 FILLER_18_357 ();
 sg13g2_decap_8 FILLER_18_364 ();
 sg13g2_decap_8 FILLER_18_371 ();
 sg13g2_decap_8 FILLER_18_378 ();
 sg13g2_decap_8 FILLER_18_385 ();
 sg13g2_decap_8 FILLER_18_392 ();
 sg13g2_decap_8 FILLER_18_399 ();
 sg13g2_fill_2 FILLER_18_406 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_fill_1 FILLER_19_98 ();
 sg13g2_decap_4 FILLER_19_116 ();
 sg13g2_decap_8 FILLER_19_129 ();
 sg13g2_fill_2 FILLER_19_136 ();
 sg13g2_decap_8 FILLER_19_143 ();
 sg13g2_fill_2 FILLER_19_150 ();
 sg13g2_fill_1 FILLER_19_152 ();
 sg13g2_decap_8 FILLER_19_163 ();
 sg13g2_decap_8 FILLER_19_170 ();
 sg13g2_decap_4 FILLER_19_177 ();
 sg13g2_fill_1 FILLER_19_195 ();
 sg13g2_fill_2 FILLER_19_214 ();
 sg13g2_fill_2 FILLER_19_230 ();
 sg13g2_fill_1 FILLER_19_237 ();
 sg13g2_decap_8 FILLER_19_306 ();
 sg13g2_decap_8 FILLER_19_313 ();
 sg13g2_decap_8 FILLER_19_320 ();
 sg13g2_decap_8 FILLER_19_327 ();
 sg13g2_decap_8 FILLER_19_334 ();
 sg13g2_decap_8 FILLER_19_341 ();
 sg13g2_decap_8 FILLER_19_348 ();
 sg13g2_decap_8 FILLER_19_355 ();
 sg13g2_decap_8 FILLER_19_362 ();
 sg13g2_decap_8 FILLER_19_369 ();
 sg13g2_decap_8 FILLER_19_376 ();
 sg13g2_decap_8 FILLER_19_383 ();
 sg13g2_decap_8 FILLER_19_390 ();
 sg13g2_decap_8 FILLER_19_397 ();
 sg13g2_decap_4 FILLER_19_404 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_4 FILLER_20_91 ();
 sg13g2_fill_1 FILLER_20_185 ();
 sg13g2_fill_2 FILLER_20_216 ();
 sg13g2_fill_2 FILLER_20_252 ();
 sg13g2_fill_1 FILLER_20_254 ();
 sg13g2_fill_1 FILLER_20_281 ();
 sg13g2_decap_8 FILLER_20_308 ();
 sg13g2_decap_8 FILLER_20_315 ();
 sg13g2_decap_8 FILLER_20_322 ();
 sg13g2_decap_8 FILLER_20_329 ();
 sg13g2_decap_8 FILLER_20_336 ();
 sg13g2_decap_8 FILLER_20_343 ();
 sg13g2_decap_8 FILLER_20_350 ();
 sg13g2_decap_8 FILLER_20_357 ();
 sg13g2_decap_8 FILLER_20_364 ();
 sg13g2_decap_8 FILLER_20_371 ();
 sg13g2_decap_8 FILLER_20_378 ();
 sg13g2_decap_8 FILLER_20_385 ();
 sg13g2_decap_8 FILLER_20_392 ();
 sg13g2_decap_8 FILLER_20_399 ();
 sg13g2_fill_2 FILLER_20_406 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_fill_1 FILLER_21_91 ();
 sg13g2_fill_1 FILLER_21_159 ();
 sg13g2_fill_1 FILLER_21_208 ();
 sg13g2_fill_1 FILLER_21_244 ();
 sg13g2_decap_8 FILLER_21_254 ();
 sg13g2_fill_1 FILLER_21_261 ();
 sg13g2_decap_8 FILLER_21_267 ();
 sg13g2_decap_8 FILLER_21_274 ();
 sg13g2_decap_8 FILLER_21_281 ();
 sg13g2_fill_2 FILLER_21_288 ();
 sg13g2_fill_1 FILLER_21_293 ();
 sg13g2_decap_8 FILLER_21_297 ();
 sg13g2_decap_8 FILLER_21_304 ();
 sg13g2_decap_8 FILLER_21_311 ();
 sg13g2_decap_8 FILLER_21_318 ();
 sg13g2_decap_8 FILLER_21_325 ();
 sg13g2_decap_8 FILLER_21_332 ();
 sg13g2_decap_8 FILLER_21_339 ();
 sg13g2_decap_8 FILLER_21_346 ();
 sg13g2_decap_8 FILLER_21_353 ();
 sg13g2_decap_8 FILLER_21_360 ();
 sg13g2_decap_8 FILLER_21_367 ();
 sg13g2_decap_8 FILLER_21_374 ();
 sg13g2_decap_8 FILLER_21_381 ();
 sg13g2_decap_8 FILLER_21_388 ();
 sg13g2_decap_8 FILLER_21_395 ();
 sg13g2_decap_8 FILLER_21_402 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_fill_1 FILLER_22_105 ();
 sg13g2_fill_2 FILLER_22_141 ();
 sg13g2_fill_1 FILLER_22_143 ();
 sg13g2_decap_4 FILLER_22_171 ();
 sg13g2_fill_1 FILLER_22_175 ();
 sg13g2_fill_2 FILLER_22_201 ();
 sg13g2_fill_2 FILLER_22_214 ();
 sg13g2_decap_8 FILLER_22_230 ();
 sg13g2_fill_2 FILLER_22_237 ();
 sg13g2_fill_1 FILLER_22_239 ();
 sg13g2_decap_4 FILLER_22_245 ();
 sg13g2_fill_1 FILLER_22_249 ();
 sg13g2_decap_4 FILLER_22_253 ();
 sg13g2_fill_2 FILLER_22_257 ();
 sg13g2_decap_4 FILLER_22_276 ();
 sg13g2_fill_2 FILLER_22_280 ();
 sg13g2_fill_1 FILLER_22_297 ();
 sg13g2_decap_8 FILLER_22_302 ();
 sg13g2_fill_1 FILLER_22_309 ();
 sg13g2_decap_8 FILLER_22_315 ();
 sg13g2_decap_8 FILLER_22_322 ();
 sg13g2_decap_8 FILLER_22_329 ();
 sg13g2_decap_8 FILLER_22_336 ();
 sg13g2_decap_8 FILLER_22_343 ();
 sg13g2_decap_8 FILLER_22_350 ();
 sg13g2_decap_8 FILLER_22_357 ();
 sg13g2_decap_8 FILLER_22_364 ();
 sg13g2_decap_8 FILLER_22_371 ();
 sg13g2_decap_8 FILLER_22_378 ();
 sg13g2_decap_8 FILLER_22_385 ();
 sg13g2_decap_8 FILLER_22_392 ();
 sg13g2_decap_8 FILLER_22_399 ();
 sg13g2_fill_2 FILLER_22_406 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_98 ();
 sg13g2_decap_8 FILLER_23_105 ();
 sg13g2_fill_2 FILLER_23_129 ();
 sg13g2_decap_4 FILLER_23_149 ();
 sg13g2_fill_1 FILLER_23_153 ();
 sg13g2_decap_8 FILLER_23_159 ();
 sg13g2_decap_8 FILLER_23_166 ();
 sg13g2_decap_8 FILLER_23_173 ();
 sg13g2_fill_1 FILLER_23_180 ();
 sg13g2_fill_1 FILLER_23_189 ();
 sg13g2_fill_2 FILLER_23_198 ();
 sg13g2_fill_1 FILLER_23_200 ();
 sg13g2_decap_8 FILLER_23_220 ();
 sg13g2_decap_4 FILLER_23_227 ();
 sg13g2_fill_2 FILLER_23_231 ();
 sg13g2_fill_2 FILLER_23_309 ();
 sg13g2_decap_8 FILLER_23_321 ();
 sg13g2_decap_8 FILLER_23_328 ();
 sg13g2_decap_8 FILLER_23_335 ();
 sg13g2_decap_8 FILLER_23_342 ();
 sg13g2_decap_8 FILLER_23_349 ();
 sg13g2_decap_8 FILLER_23_356 ();
 sg13g2_decap_8 FILLER_23_363 ();
 sg13g2_decap_8 FILLER_23_370 ();
 sg13g2_decap_8 FILLER_23_377 ();
 sg13g2_decap_8 FILLER_23_384 ();
 sg13g2_decap_8 FILLER_23_391 ();
 sg13g2_decap_8 FILLER_23_398 ();
 sg13g2_decap_4 FILLER_23_405 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_decap_8 FILLER_24_98 ();
 sg13g2_fill_1 FILLER_24_105 ();
 sg13g2_fill_2 FILLER_24_120 ();
 sg13g2_fill_1 FILLER_24_122 ();
 sg13g2_decap_8 FILLER_24_130 ();
 sg13g2_decap_8 FILLER_24_137 ();
 sg13g2_decap_8 FILLER_24_144 ();
 sg13g2_decap_8 FILLER_24_151 ();
 sg13g2_fill_2 FILLER_24_184 ();
 sg13g2_fill_2 FILLER_24_225 ();
 sg13g2_fill_1 FILLER_24_227 ();
 sg13g2_fill_2 FILLER_24_266 ();
 sg13g2_decap_4 FILLER_24_305 ();
 sg13g2_fill_1 FILLER_24_309 ();
 sg13g2_decap_8 FILLER_24_318 ();
 sg13g2_decap_8 FILLER_24_325 ();
 sg13g2_decap_8 FILLER_24_332 ();
 sg13g2_decap_8 FILLER_24_339 ();
 sg13g2_decap_8 FILLER_24_346 ();
 sg13g2_decap_8 FILLER_24_353 ();
 sg13g2_decap_8 FILLER_24_360 ();
 sg13g2_decap_8 FILLER_24_367 ();
 sg13g2_decap_8 FILLER_24_374 ();
 sg13g2_decap_8 FILLER_24_381 ();
 sg13g2_decap_8 FILLER_24_388 ();
 sg13g2_decap_8 FILLER_24_395 ();
 sg13g2_decap_8 FILLER_24_402 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_fill_2 FILLER_25_91 ();
 sg13g2_fill_1 FILLER_25_93 ();
 sg13g2_fill_2 FILLER_25_129 ();
 sg13g2_fill_1 FILLER_25_131 ();
 sg13g2_fill_1 FILLER_25_153 ();
 sg13g2_fill_2 FILLER_25_198 ();
 sg13g2_decap_4 FILLER_25_211 ();
 sg13g2_fill_1 FILLER_25_215 ();
 sg13g2_decap_4 FILLER_25_242 ();
 sg13g2_fill_1 FILLER_25_246 ();
 sg13g2_fill_2 FILLER_25_279 ();
 sg13g2_decap_8 FILLER_25_315 ();
 sg13g2_decap_8 FILLER_25_322 ();
 sg13g2_decap_8 FILLER_25_329 ();
 sg13g2_decap_8 FILLER_25_336 ();
 sg13g2_decap_8 FILLER_25_343 ();
 sg13g2_decap_8 FILLER_25_350 ();
 sg13g2_decap_8 FILLER_25_357 ();
 sg13g2_decap_8 FILLER_25_364 ();
 sg13g2_decap_8 FILLER_25_371 ();
 sg13g2_decap_8 FILLER_25_378 ();
 sg13g2_decap_8 FILLER_25_385 ();
 sg13g2_decap_8 FILLER_25_392 ();
 sg13g2_decap_8 FILLER_25_399 ();
 sg13g2_fill_2 FILLER_25_406 ();
 sg13g2_fill_1 FILLER_25_408 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_fill_1 FILLER_26_84 ();
 sg13g2_decap_4 FILLER_26_162 ();
 sg13g2_decap_4 FILLER_26_171 ();
 sg13g2_decap_4 FILLER_26_213 ();
 sg13g2_fill_1 FILLER_26_217 ();
 sg13g2_fill_2 FILLER_26_235 ();
 sg13g2_fill_1 FILLER_26_237 ();
 sg13g2_decap_4 FILLER_26_250 ();
 sg13g2_fill_1 FILLER_26_289 ();
 sg13g2_decap_8 FILLER_26_316 ();
 sg13g2_decap_8 FILLER_26_323 ();
 sg13g2_decap_8 FILLER_26_330 ();
 sg13g2_decap_8 FILLER_26_337 ();
 sg13g2_decap_8 FILLER_26_344 ();
 sg13g2_decap_8 FILLER_26_351 ();
 sg13g2_decap_8 FILLER_26_358 ();
 sg13g2_decap_8 FILLER_26_365 ();
 sg13g2_decap_8 FILLER_26_372 ();
 sg13g2_decap_8 FILLER_26_379 ();
 sg13g2_decap_8 FILLER_26_386 ();
 sg13g2_decap_8 FILLER_26_393 ();
 sg13g2_decap_8 FILLER_26_400 ();
 sg13g2_fill_2 FILLER_26_407 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_decap_8 FILLER_27_84 ();
 sg13g2_fill_2 FILLER_27_91 ();
 sg13g2_fill_2 FILLER_27_128 ();
 sg13g2_fill_1 FILLER_27_130 ();
 sg13g2_fill_2 FILLER_27_139 ();
 sg13g2_fill_2 FILLER_27_149 ();
 sg13g2_fill_2 FILLER_27_185 ();
 sg13g2_fill_1 FILLER_27_209 ();
 sg13g2_fill_1 FILLER_27_248 ();
 sg13g2_fill_2 FILLER_27_268 ();
 sg13g2_fill_2 FILLER_27_275 ();
 sg13g2_fill_2 FILLER_27_286 ();
 sg13g2_fill_1 FILLER_27_319 ();
 sg13g2_decap_8 FILLER_27_346 ();
 sg13g2_decap_8 FILLER_27_353 ();
 sg13g2_decap_8 FILLER_27_360 ();
 sg13g2_decap_8 FILLER_27_367 ();
 sg13g2_decap_8 FILLER_27_374 ();
 sg13g2_decap_8 FILLER_27_381 ();
 sg13g2_decap_8 FILLER_27_388 ();
 sg13g2_decap_8 FILLER_27_395 ();
 sg13g2_decap_8 FILLER_27_402 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_decap_8 FILLER_28_84 ();
 sg13g2_decap_8 FILLER_28_91 ();
 sg13g2_decap_4 FILLER_28_102 ();
 sg13g2_decap_8 FILLER_28_160 ();
 sg13g2_decap_8 FILLER_28_167 ();
 sg13g2_fill_2 FILLER_28_174 ();
 sg13g2_fill_2 FILLER_28_184 ();
 sg13g2_fill_2 FILLER_28_262 ();
 sg13g2_fill_1 FILLER_28_264 ();
 sg13g2_decap_8 FILLER_28_347 ();
 sg13g2_decap_8 FILLER_28_354 ();
 sg13g2_decap_8 FILLER_28_361 ();
 sg13g2_decap_8 FILLER_28_368 ();
 sg13g2_decap_8 FILLER_28_375 ();
 sg13g2_decap_8 FILLER_28_382 ();
 sg13g2_decap_8 FILLER_28_389 ();
 sg13g2_decap_8 FILLER_28_396 ();
 sg13g2_decap_4 FILLER_28_403 ();
 sg13g2_fill_2 FILLER_28_407 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_decap_8 FILLER_29_84 ();
 sg13g2_decap_8 FILLER_29_91 ();
 sg13g2_decap_8 FILLER_29_98 ();
 sg13g2_fill_2 FILLER_29_105 ();
 sg13g2_fill_2 FILLER_29_115 ();
 sg13g2_fill_2 FILLER_29_123 ();
 sg13g2_fill_2 FILLER_29_136 ();
 sg13g2_fill_1 FILLER_29_138 ();
 sg13g2_fill_1 FILLER_29_146 ();
 sg13g2_decap_8 FILLER_29_161 ();
 sg13g2_fill_2 FILLER_29_168 ();
 sg13g2_fill_1 FILLER_29_170 ();
 sg13g2_decap_8 FILLER_29_175 ();
 sg13g2_decap_8 FILLER_29_182 ();
 sg13g2_decap_8 FILLER_29_189 ();
 sg13g2_fill_1 FILLER_29_196 ();
 sg13g2_fill_2 FILLER_29_211 ();
 sg13g2_fill_1 FILLER_29_213 ();
 sg13g2_fill_1 FILLER_29_218 ();
 sg13g2_fill_2 FILLER_29_249 ();
 sg13g2_decap_4 FILLER_29_304 ();
 sg13g2_fill_2 FILLER_29_308 ();
 sg13g2_fill_1 FILLER_29_341 ();
 sg13g2_decap_8 FILLER_29_351 ();
 sg13g2_decap_8 FILLER_29_358 ();
 sg13g2_decap_8 FILLER_29_365 ();
 sg13g2_decap_8 FILLER_29_372 ();
 sg13g2_decap_8 FILLER_29_379 ();
 sg13g2_decap_8 FILLER_29_386 ();
 sg13g2_decap_8 FILLER_29_393 ();
 sg13g2_decap_8 FILLER_29_400 ();
 sg13g2_fill_2 FILLER_29_407 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_77 ();
 sg13g2_decap_8 FILLER_30_84 ();
 sg13g2_decap_8 FILLER_30_91 ();
 sg13g2_decap_8 FILLER_30_98 ();
 sg13g2_fill_2 FILLER_30_105 ();
 sg13g2_fill_1 FILLER_30_107 ();
 sg13g2_decap_4 FILLER_30_128 ();
 sg13g2_fill_2 FILLER_30_141 ();
 sg13g2_fill_1 FILLER_30_169 ();
 sg13g2_decap_8 FILLER_30_189 ();
 sg13g2_decap_8 FILLER_30_196 ();
 sg13g2_decap_8 FILLER_30_203 ();
 sg13g2_fill_1 FILLER_30_210 ();
 sg13g2_decap_8 FILLER_30_216 ();
 sg13g2_decap_8 FILLER_30_223 ();
 sg13g2_fill_1 FILLER_30_255 ();
 sg13g2_fill_2 FILLER_30_264 ();
 sg13g2_fill_1 FILLER_30_266 ();
 sg13g2_fill_1 FILLER_30_284 ();
 sg13g2_fill_2 FILLER_30_290 ();
 sg13g2_fill_2 FILLER_30_323 ();
 sg13g2_decap_8 FILLER_30_356 ();
 sg13g2_decap_8 FILLER_30_363 ();
 sg13g2_decap_8 FILLER_30_370 ();
 sg13g2_decap_8 FILLER_30_377 ();
 sg13g2_decap_8 FILLER_30_384 ();
 sg13g2_decap_8 FILLER_30_391 ();
 sg13g2_decap_8 FILLER_30_398 ();
 sg13g2_decap_4 FILLER_30_405 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_decap_8 FILLER_31_84 ();
 sg13g2_decap_8 FILLER_31_91 ();
 sg13g2_fill_1 FILLER_31_98 ();
 sg13g2_fill_2 FILLER_31_142 ();
 sg13g2_fill_1 FILLER_31_170 ();
 sg13g2_fill_1 FILLER_31_188 ();
 sg13g2_decap_8 FILLER_31_200 ();
 sg13g2_fill_1 FILLER_31_207 ();
 sg13g2_fill_1 FILLER_31_213 ();
 sg13g2_fill_1 FILLER_31_225 ();
 sg13g2_decap_4 FILLER_31_238 ();
 sg13g2_fill_2 FILLER_31_242 ();
 sg13g2_fill_2 FILLER_31_251 ();
 sg13g2_fill_2 FILLER_31_263 ();
 sg13g2_fill_1 FILLER_31_265 ();
 sg13g2_fill_1 FILLER_31_279 ();
 sg13g2_decap_4 FILLER_31_284 ();
 sg13g2_decap_8 FILLER_31_363 ();
 sg13g2_decap_8 FILLER_31_370 ();
 sg13g2_decap_8 FILLER_31_377 ();
 sg13g2_decap_8 FILLER_31_384 ();
 sg13g2_decap_8 FILLER_31_391 ();
 sg13g2_decap_8 FILLER_31_398 ();
 sg13g2_decap_4 FILLER_31_405 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_fill_2 FILLER_32_70 ();
 sg13g2_fill_2 FILLER_32_98 ();
 sg13g2_fill_2 FILLER_32_143 ();
 sg13g2_fill_1 FILLER_32_202 ();
 sg13g2_decap_8 FILLER_32_225 ();
 sg13g2_fill_1 FILLER_32_232 ();
 sg13g2_fill_1 FILLER_32_237 ();
 sg13g2_fill_2 FILLER_32_243 ();
 sg13g2_decap_8 FILLER_32_257 ();
 sg13g2_decap_4 FILLER_32_264 ();
 sg13g2_fill_1 FILLER_32_271 ();
 sg13g2_decap_4 FILLER_32_275 ();
 sg13g2_fill_2 FILLER_32_279 ();
 sg13g2_fill_1 FILLER_32_316 ();
 sg13g2_decap_4 FILLER_32_343 ();
 sg13g2_fill_1 FILLER_32_347 ();
 sg13g2_decap_8 FILLER_32_353 ();
 sg13g2_decap_8 FILLER_32_360 ();
 sg13g2_decap_8 FILLER_32_367 ();
 sg13g2_decap_8 FILLER_32_374 ();
 sg13g2_decap_8 FILLER_32_381 ();
 sg13g2_decap_8 FILLER_32_388 ();
 sg13g2_decap_8 FILLER_32_395 ();
 sg13g2_decap_8 FILLER_32_402 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_fill_2 FILLER_33_63 ();
 sg13g2_fill_1 FILLER_33_65 ();
 sg13g2_decap_8 FILLER_33_149 ();
 sg13g2_decap_8 FILLER_33_156 ();
 sg13g2_decap_4 FILLER_33_163 ();
 sg13g2_fill_2 FILLER_33_194 ();
 sg13g2_fill_1 FILLER_33_196 ();
 sg13g2_fill_1 FILLER_33_211 ();
 sg13g2_decap_4 FILLER_33_226 ();
 sg13g2_decap_4 FILLER_33_235 ();
 sg13g2_decap_4 FILLER_33_259 ();
 sg13g2_decap_8 FILLER_33_297 ();
 sg13g2_decap_8 FILLER_33_304 ();
 sg13g2_fill_2 FILLER_33_311 ();
 sg13g2_fill_1 FILLER_33_313 ();
 sg13g2_decap_8 FILLER_33_331 ();
 sg13g2_decap_8 FILLER_33_338 ();
 sg13g2_decap_4 FILLER_33_345 ();
 sg13g2_fill_1 FILLER_33_349 ();
 sg13g2_decap_8 FILLER_33_354 ();
 sg13g2_decap_8 FILLER_33_361 ();
 sg13g2_decap_8 FILLER_33_368 ();
 sg13g2_decap_8 FILLER_33_375 ();
 sg13g2_decap_8 FILLER_33_382 ();
 sg13g2_decap_8 FILLER_33_389 ();
 sg13g2_decap_8 FILLER_33_396 ();
 sg13g2_decap_4 FILLER_33_403 ();
 sg13g2_fill_2 FILLER_33_407 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_4 FILLER_34_63 ();
 sg13g2_fill_1 FILLER_34_67 ();
 sg13g2_fill_1 FILLER_34_103 ();
 sg13g2_fill_2 FILLER_34_127 ();
 sg13g2_fill_2 FILLER_34_178 ();
 sg13g2_decap_8 FILLER_34_216 ();
 sg13g2_fill_1 FILLER_34_223 ();
 sg13g2_fill_2 FILLER_34_267 ();
 sg13g2_decap_8 FILLER_34_303 ();
 sg13g2_decap_4 FILLER_34_310 ();
 sg13g2_fill_1 FILLER_34_314 ();
 sg13g2_fill_1 FILLER_34_333 ();
 sg13g2_decap_8 FILLER_34_342 ();
 sg13g2_fill_2 FILLER_34_349 ();
 sg13g2_decap_8 FILLER_34_362 ();
 sg13g2_decap_8 FILLER_34_369 ();
 sg13g2_decap_8 FILLER_34_376 ();
 sg13g2_decap_8 FILLER_34_383 ();
 sg13g2_decap_8 FILLER_34_390 ();
 sg13g2_decap_8 FILLER_34_397 ();
 sg13g2_decap_4 FILLER_34_404 ();
 sg13g2_fill_1 FILLER_34_408 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_fill_1 FILLER_35_110 ();
 sg13g2_fill_2 FILLER_35_208 ();
 sg13g2_fill_1 FILLER_35_210 ();
 sg13g2_decap_4 FILLER_35_225 ();
 sg13g2_fill_1 FILLER_35_229 ();
 sg13g2_decap_8 FILLER_35_236 ();
 sg13g2_decap_8 FILLER_35_243 ();
 sg13g2_fill_2 FILLER_35_250 ();
 sg13g2_decap_4 FILLER_35_273 ();
 sg13g2_fill_1 FILLER_35_291 ();
 sg13g2_fill_1 FILLER_35_318 ();
 sg13g2_fill_1 FILLER_35_335 ();
 sg13g2_decap_8 FILLER_35_362 ();
 sg13g2_decap_8 FILLER_35_369 ();
 sg13g2_decap_8 FILLER_35_376 ();
 sg13g2_decap_8 FILLER_35_383 ();
 sg13g2_decap_8 FILLER_35_390 ();
 sg13g2_decap_8 FILLER_35_397 ();
 sg13g2_decap_4 FILLER_35_404 ();
 sg13g2_fill_1 FILLER_35_408 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_fill_2 FILLER_36_63 ();
 sg13g2_decap_4 FILLER_36_121 ();
 sg13g2_fill_2 FILLER_36_125 ();
 sg13g2_decap_4 FILLER_36_167 ();
 sg13g2_fill_1 FILLER_36_176 ();
 sg13g2_fill_2 FILLER_36_230 ();
 sg13g2_fill_1 FILLER_36_232 ();
 sg13g2_decap_8 FILLER_36_238 ();
 sg13g2_decap_4 FILLER_36_245 ();
 sg13g2_decap_8 FILLER_36_253 ();
 sg13g2_fill_2 FILLER_36_260 ();
 sg13g2_fill_2 FILLER_36_270 ();
 sg13g2_fill_1 FILLER_36_272 ();
 sg13g2_fill_2 FILLER_36_279 ();
 sg13g2_fill_1 FILLER_36_298 ();
 sg13g2_decap_4 FILLER_36_327 ();
 sg13g2_fill_2 FILLER_36_331 ();
 sg13g2_decap_8 FILLER_36_357 ();
 sg13g2_decap_8 FILLER_36_364 ();
 sg13g2_decap_8 FILLER_36_371 ();
 sg13g2_decap_8 FILLER_36_378 ();
 sg13g2_decap_8 FILLER_36_385 ();
 sg13g2_decap_8 FILLER_36_392 ();
 sg13g2_decap_8 FILLER_36_399 ();
 sg13g2_fill_2 FILLER_36_406 ();
 sg13g2_fill_1 FILLER_36_408 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_4 FILLER_37_70 ();
 sg13g2_fill_2 FILLER_37_134 ();
 sg13g2_fill_1 FILLER_37_136 ();
 sg13g2_decap_4 FILLER_37_149 ();
 sg13g2_decap_8 FILLER_37_158 ();
 sg13g2_fill_2 FILLER_37_165 ();
 sg13g2_fill_1 FILLER_37_167 ();
 sg13g2_decap_4 FILLER_37_290 ();
 sg13g2_fill_1 FILLER_37_302 ();
 sg13g2_fill_2 FILLER_37_308 ();
 sg13g2_fill_2 FILLER_37_320 ();
 sg13g2_fill_1 FILLER_37_322 ();
 sg13g2_decap_8 FILLER_37_351 ();
 sg13g2_decap_8 FILLER_37_358 ();
 sg13g2_decap_8 FILLER_37_365 ();
 sg13g2_decap_8 FILLER_37_372 ();
 sg13g2_decap_8 FILLER_37_379 ();
 sg13g2_decap_8 FILLER_37_386 ();
 sg13g2_decap_8 FILLER_37_393 ();
 sg13g2_decap_8 FILLER_37_400 ();
 sg13g2_fill_2 FILLER_37_407 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_8 FILLER_38_56 ();
 sg13g2_decap_8 FILLER_38_63 ();
 sg13g2_decap_8 FILLER_38_70 ();
 sg13g2_decap_8 FILLER_38_77 ();
 sg13g2_decap_8 FILLER_38_84 ();
 sg13g2_decap_4 FILLER_38_91 ();
 sg13g2_fill_2 FILLER_38_95 ();
 sg13g2_fill_2 FILLER_38_142 ();
 sg13g2_fill_2 FILLER_38_182 ();
 sg13g2_decap_8 FILLER_38_216 ();
 sg13g2_decap_8 FILLER_38_223 ();
 sg13g2_fill_1 FILLER_38_230 ();
 sg13g2_fill_2 FILLER_38_266 ();
 sg13g2_decap_4 FILLER_38_283 ();
 sg13g2_fill_2 FILLER_38_320 ();
 sg13g2_fill_1 FILLER_38_322 ();
 sg13g2_fill_2 FILLER_38_331 ();
 sg13g2_fill_1 FILLER_38_333 ();
 sg13g2_decap_8 FILLER_38_360 ();
 sg13g2_decap_8 FILLER_38_367 ();
 sg13g2_decap_8 FILLER_38_374 ();
 sg13g2_decap_8 FILLER_38_381 ();
 sg13g2_decap_8 FILLER_38_388 ();
 sg13g2_decap_8 FILLER_38_395 ();
 sg13g2_decap_8 FILLER_38_402 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_14 ();
 sg13g2_decap_8 FILLER_39_21 ();
 sg13g2_decap_8 FILLER_39_28 ();
 sg13g2_decap_8 FILLER_39_35 ();
 sg13g2_decap_8 FILLER_39_42 ();
 sg13g2_decap_8 FILLER_39_49 ();
 sg13g2_decap_8 FILLER_39_56 ();
 sg13g2_decap_8 FILLER_39_63 ();
 sg13g2_decap_8 FILLER_39_70 ();
 sg13g2_decap_8 FILLER_39_77 ();
 sg13g2_fill_2 FILLER_39_84 ();
 sg13g2_fill_1 FILLER_39_112 ();
 sg13g2_fill_1 FILLER_39_122 ();
 sg13g2_fill_2 FILLER_39_175 ();
 sg13g2_fill_2 FILLER_39_185 ();
 sg13g2_decap_8 FILLER_39_200 ();
 sg13g2_decap_8 FILLER_39_207 ();
 sg13g2_decap_8 FILLER_39_214 ();
 sg13g2_decap_8 FILLER_39_221 ();
 sg13g2_fill_2 FILLER_39_237 ();
 sg13g2_fill_1 FILLER_39_244 ();
 sg13g2_fill_1 FILLER_39_313 ();
 sg13g2_decap_4 FILLER_39_327 ();
 sg13g2_fill_1 FILLER_39_331 ();
 sg13g2_decap_8 FILLER_39_363 ();
 sg13g2_decap_8 FILLER_39_370 ();
 sg13g2_decap_8 FILLER_39_377 ();
 sg13g2_decap_8 FILLER_39_384 ();
 sg13g2_decap_8 FILLER_39_391 ();
 sg13g2_decap_8 FILLER_39_398 ();
 sg13g2_decap_4 FILLER_39_405 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_14 ();
 sg13g2_decap_8 FILLER_40_21 ();
 sg13g2_decap_8 FILLER_40_28 ();
 sg13g2_decap_8 FILLER_40_35 ();
 sg13g2_decap_8 FILLER_40_42 ();
 sg13g2_decap_8 FILLER_40_49 ();
 sg13g2_decap_8 FILLER_40_56 ();
 sg13g2_decap_8 FILLER_40_63 ();
 sg13g2_fill_2 FILLER_40_70 ();
 sg13g2_fill_1 FILLER_40_110 ();
 sg13g2_fill_2 FILLER_40_152 ();
 sg13g2_fill_1 FILLER_40_173 ();
 sg13g2_fill_1 FILLER_40_190 ();
 sg13g2_fill_1 FILLER_40_217 ();
 sg13g2_decap_8 FILLER_40_261 ();
 sg13g2_fill_1 FILLER_40_268 ();
 sg13g2_fill_2 FILLER_40_274 ();
 sg13g2_fill_1 FILLER_40_276 ();
 sg13g2_decap_4 FILLER_40_285 ();
 sg13g2_fill_1 FILLER_40_289 ();
 sg13g2_fill_2 FILLER_40_293 ();
 sg13g2_decap_4 FILLER_40_299 ();
 sg13g2_fill_1 FILLER_40_306 ();
 sg13g2_fill_2 FILLER_40_318 ();
 sg13g2_fill_2 FILLER_40_332 ();
 sg13g2_fill_1 FILLER_40_339 ();
 sg13g2_decap_8 FILLER_40_349 ();
 sg13g2_decap_8 FILLER_40_356 ();
 sg13g2_decap_8 FILLER_40_363 ();
 sg13g2_decap_8 FILLER_40_370 ();
 sg13g2_decap_8 FILLER_40_377 ();
 sg13g2_decap_8 FILLER_40_384 ();
 sg13g2_decap_8 FILLER_40_391 ();
 sg13g2_decap_8 FILLER_40_398 ();
 sg13g2_decap_4 FILLER_40_405 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_8 FILLER_41_14 ();
 sg13g2_decap_8 FILLER_41_21 ();
 sg13g2_decap_8 FILLER_41_28 ();
 sg13g2_decap_8 FILLER_41_35 ();
 sg13g2_decap_8 FILLER_41_42 ();
 sg13g2_decap_8 FILLER_41_49 ();
 sg13g2_decap_8 FILLER_41_56 ();
 sg13g2_fill_2 FILLER_41_63 ();
 sg13g2_fill_1 FILLER_41_65 ();
 sg13g2_fill_2 FILLER_41_150 ();
 sg13g2_fill_1 FILLER_41_152 ();
 sg13g2_fill_1 FILLER_41_176 ();
 sg13g2_decap_4 FILLER_41_190 ();
 sg13g2_fill_2 FILLER_41_194 ();
 sg13g2_decap_8 FILLER_41_199 ();
 sg13g2_decap_8 FILLER_41_244 ();
 sg13g2_decap_4 FILLER_41_251 ();
 sg13g2_decap_8 FILLER_41_259 ();
 sg13g2_fill_2 FILLER_41_266 ();
 sg13g2_decap_8 FILLER_41_273 ();
 sg13g2_decap_4 FILLER_41_280 ();
 sg13g2_fill_2 FILLER_41_287 ();
 sg13g2_fill_2 FILLER_41_321 ();
 sg13g2_fill_2 FILLER_41_331 ();
 sg13g2_decap_8 FILLER_41_359 ();
 sg13g2_decap_8 FILLER_41_366 ();
 sg13g2_decap_8 FILLER_41_373 ();
 sg13g2_decap_8 FILLER_41_380 ();
 sg13g2_decap_8 FILLER_41_387 ();
 sg13g2_decap_8 FILLER_41_394 ();
 sg13g2_decap_8 FILLER_41_401 ();
 sg13g2_fill_1 FILLER_41_408 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_decap_8 FILLER_42_14 ();
 sg13g2_decap_8 FILLER_42_21 ();
 sg13g2_decap_8 FILLER_42_28 ();
 sg13g2_decap_8 FILLER_42_35 ();
 sg13g2_decap_8 FILLER_42_42 ();
 sg13g2_decap_8 FILLER_42_49 ();
 sg13g2_decap_8 FILLER_42_56 ();
 sg13g2_decap_8 FILLER_42_63 ();
 sg13g2_decap_4 FILLER_42_70 ();
 sg13g2_decap_4 FILLER_42_113 ();
 sg13g2_fill_2 FILLER_42_117 ();
 sg13g2_fill_1 FILLER_42_126 ();
 sg13g2_fill_1 FILLER_42_168 ();
 sg13g2_fill_2 FILLER_42_178 ();
 sg13g2_decap_8 FILLER_42_206 ();
 sg13g2_fill_1 FILLER_42_213 ();
 sg13g2_fill_1 FILLER_42_219 ();
 sg13g2_decap_8 FILLER_42_229 ();
 sg13g2_decap_8 FILLER_42_236 ();
 sg13g2_fill_2 FILLER_42_243 ();
 sg13g2_fill_1 FILLER_42_245 ();
 sg13g2_fill_1 FILLER_42_272 ();
 sg13g2_fill_1 FILLER_42_286 ();
 sg13g2_fill_1 FILLER_42_308 ();
 sg13g2_decap_4 FILLER_42_352 ();
 sg13g2_decap_8 FILLER_42_359 ();
 sg13g2_decap_8 FILLER_42_366 ();
 sg13g2_decap_8 FILLER_42_373 ();
 sg13g2_decap_8 FILLER_42_380 ();
 sg13g2_decap_8 FILLER_42_387 ();
 sg13g2_decap_8 FILLER_42_394 ();
 sg13g2_decap_8 FILLER_42_401 ();
 sg13g2_fill_1 FILLER_42_408 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_decap_8 FILLER_43_14 ();
 sg13g2_decap_8 FILLER_43_21 ();
 sg13g2_decap_8 FILLER_43_28 ();
 sg13g2_decap_8 FILLER_43_35 ();
 sg13g2_decap_8 FILLER_43_42 ();
 sg13g2_decap_8 FILLER_43_49 ();
 sg13g2_decap_8 FILLER_43_56 ();
 sg13g2_decap_8 FILLER_43_63 ();
 sg13g2_decap_8 FILLER_43_70 ();
 sg13g2_decap_4 FILLER_43_77 ();
 sg13g2_fill_1 FILLER_43_81 ();
 sg13g2_fill_1 FILLER_43_108 ();
 sg13g2_decap_4 FILLER_43_122 ();
 sg13g2_fill_2 FILLER_43_227 ();
 sg13g2_fill_1 FILLER_43_229 ();
 sg13g2_fill_1 FILLER_43_312 ();
 sg13g2_decap_8 FILLER_43_326 ();
 sg13g2_decap_4 FILLER_43_333 ();
 sg13g2_decap_8 FILLER_43_368 ();
 sg13g2_decap_8 FILLER_43_375 ();
 sg13g2_decap_8 FILLER_43_382 ();
 sg13g2_decap_8 FILLER_43_389 ();
 sg13g2_decap_8 FILLER_43_396 ();
 sg13g2_decap_4 FILLER_43_403 ();
 sg13g2_fill_2 FILLER_43_407 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_decap_8 FILLER_44_14 ();
 sg13g2_decap_8 FILLER_44_21 ();
 sg13g2_decap_8 FILLER_44_28 ();
 sg13g2_decap_8 FILLER_44_35 ();
 sg13g2_decap_8 FILLER_44_42 ();
 sg13g2_decap_8 FILLER_44_49 ();
 sg13g2_decap_8 FILLER_44_56 ();
 sg13g2_decap_8 FILLER_44_63 ();
 sg13g2_decap_8 FILLER_44_70 ();
 sg13g2_decap_4 FILLER_44_94 ();
 sg13g2_fill_2 FILLER_44_110 ();
 sg13g2_fill_1 FILLER_44_112 ();
 sg13g2_fill_1 FILLER_44_160 ();
 sg13g2_fill_2 FILLER_44_187 ();
 sg13g2_fill_1 FILLER_44_256 ();
 sg13g2_fill_2 FILLER_44_293 ();
 sg13g2_decap_8 FILLER_44_320 ();
 sg13g2_fill_2 FILLER_44_327 ();
 sg13g2_fill_1 FILLER_44_329 ();
 sg13g2_decap_8 FILLER_44_367 ();
 sg13g2_decap_8 FILLER_44_374 ();
 sg13g2_decap_8 FILLER_44_381 ();
 sg13g2_decap_8 FILLER_44_388 ();
 sg13g2_decap_8 FILLER_44_395 ();
 sg13g2_decap_8 FILLER_44_402 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_7 ();
 sg13g2_decap_8 FILLER_45_14 ();
 sg13g2_decap_8 FILLER_45_21 ();
 sg13g2_decap_8 FILLER_45_28 ();
 sg13g2_decap_8 FILLER_45_35 ();
 sg13g2_decap_8 FILLER_45_42 ();
 sg13g2_decap_8 FILLER_45_49 ();
 sg13g2_decap_8 FILLER_45_56 ();
 sg13g2_decap_8 FILLER_45_63 ();
 sg13g2_decap_8 FILLER_45_70 ();
 sg13g2_decap_4 FILLER_45_77 ();
 sg13g2_fill_2 FILLER_45_81 ();
 sg13g2_fill_1 FILLER_45_162 ();
 sg13g2_decap_8 FILLER_45_178 ();
 sg13g2_decap_4 FILLER_45_190 ();
 sg13g2_decap_8 FILLER_45_197 ();
 sg13g2_decap_8 FILLER_45_204 ();
 sg13g2_decap_4 FILLER_45_211 ();
 sg13g2_fill_1 FILLER_45_215 ();
 sg13g2_decap_8 FILLER_45_219 ();
 sg13g2_decap_8 FILLER_45_226 ();
 sg13g2_fill_1 FILLER_45_233 ();
 sg13g2_decap_4 FILLER_45_245 ();
 sg13g2_fill_1 FILLER_45_249 ();
 sg13g2_fill_1 FILLER_45_275 ();
 sg13g2_fill_2 FILLER_45_282 ();
 sg13g2_decap_4 FILLER_45_310 ();
 sg13g2_decap_8 FILLER_45_349 ();
 sg13g2_decap_8 FILLER_45_360 ();
 sg13g2_decap_8 FILLER_45_367 ();
 sg13g2_decap_8 FILLER_45_374 ();
 sg13g2_decap_8 FILLER_45_381 ();
 sg13g2_decap_8 FILLER_45_388 ();
 sg13g2_decap_8 FILLER_45_395 ();
 sg13g2_decap_8 FILLER_45_402 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_7 ();
 sg13g2_decap_8 FILLER_46_14 ();
 sg13g2_decap_8 FILLER_46_21 ();
 sg13g2_decap_8 FILLER_46_28 ();
 sg13g2_decap_8 FILLER_46_35 ();
 sg13g2_decap_8 FILLER_46_42 ();
 sg13g2_decap_8 FILLER_46_49 ();
 sg13g2_decap_8 FILLER_46_56 ();
 sg13g2_decap_8 FILLER_46_63 ();
 sg13g2_decap_8 FILLER_46_70 ();
 sg13g2_decap_8 FILLER_46_77 ();
 sg13g2_decap_4 FILLER_46_84 ();
 sg13g2_fill_2 FILLER_46_103 ();
 sg13g2_fill_2 FILLER_46_157 ();
 sg13g2_fill_2 FILLER_46_185 ();
 sg13g2_decap_8 FILLER_46_195 ();
 sg13g2_fill_1 FILLER_46_212 ();
 sg13g2_fill_2 FILLER_46_221 ();
 sg13g2_decap_4 FILLER_46_236 ();
 sg13g2_decap_8 FILLER_46_249 ();
 sg13g2_decap_8 FILLER_46_256 ();
 sg13g2_decap_4 FILLER_46_263 ();
 sg13g2_decap_8 FILLER_46_307 ();
 sg13g2_decap_4 FILLER_46_314 ();
 sg13g2_fill_1 FILLER_46_318 ();
 sg13g2_decap_8 FILLER_46_328 ();
 sg13g2_decap_8 FILLER_46_335 ();
 sg13g2_decap_8 FILLER_46_342 ();
 sg13g2_decap_8 FILLER_46_349 ();
 sg13g2_fill_1 FILLER_46_356 ();
 sg13g2_decap_8 FILLER_46_360 ();
 sg13g2_decap_8 FILLER_46_367 ();
 sg13g2_decap_8 FILLER_46_374 ();
 sg13g2_decap_8 FILLER_46_381 ();
 sg13g2_decap_8 FILLER_46_388 ();
 sg13g2_decap_8 FILLER_46_395 ();
 sg13g2_decap_8 FILLER_46_402 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_7 ();
 sg13g2_decap_8 FILLER_47_14 ();
 sg13g2_decap_8 FILLER_47_21 ();
 sg13g2_decap_8 FILLER_47_28 ();
 sg13g2_decap_8 FILLER_47_35 ();
 sg13g2_decap_8 FILLER_47_42 ();
 sg13g2_decap_8 FILLER_47_49 ();
 sg13g2_decap_8 FILLER_47_56 ();
 sg13g2_decap_8 FILLER_47_63 ();
 sg13g2_decap_8 FILLER_47_70 ();
 sg13g2_fill_2 FILLER_47_77 ();
 sg13g2_fill_1 FILLER_47_109 ();
 sg13g2_fill_2 FILLER_47_205 ();
 sg13g2_fill_2 FILLER_47_212 ();
 sg13g2_fill_1 FILLER_47_219 ();
 sg13g2_decap_8 FILLER_47_243 ();
 sg13g2_fill_2 FILLER_47_254 ();
 sg13g2_fill_2 FILLER_47_280 ();
 sg13g2_fill_2 FILLER_47_311 ();
 sg13g2_fill_2 FILLER_47_330 ();
 sg13g2_decap_8 FILLER_47_358 ();
 sg13g2_decap_8 FILLER_47_365 ();
 sg13g2_decap_8 FILLER_47_372 ();
 sg13g2_decap_8 FILLER_47_379 ();
 sg13g2_decap_8 FILLER_47_386 ();
 sg13g2_decap_8 FILLER_47_393 ();
 sg13g2_decap_8 FILLER_47_400 ();
 sg13g2_fill_2 FILLER_47_407 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_decap_8 FILLER_48_14 ();
 sg13g2_decap_8 FILLER_48_21 ();
 sg13g2_decap_8 FILLER_48_28 ();
 sg13g2_decap_8 FILLER_48_35 ();
 sg13g2_decap_8 FILLER_48_42 ();
 sg13g2_decap_8 FILLER_48_49 ();
 sg13g2_decap_8 FILLER_48_56 ();
 sg13g2_decap_8 FILLER_48_63 ();
 sg13g2_decap_8 FILLER_48_70 ();
 sg13g2_decap_4 FILLER_48_77 ();
 sg13g2_fill_2 FILLER_48_81 ();
 sg13g2_fill_1 FILLER_48_130 ();
 sg13g2_decap_8 FILLER_48_172 ();
 sg13g2_decap_8 FILLER_48_188 ();
 sg13g2_fill_2 FILLER_48_203 ();
 sg13g2_fill_1 FILLER_48_205 ();
 sg13g2_fill_1 FILLER_48_214 ();
 sg13g2_fill_1 FILLER_48_300 ();
 sg13g2_fill_1 FILLER_48_305 ();
 sg13g2_fill_1 FILLER_48_326 ();
 sg13g2_fill_2 FILLER_48_353 ();
 sg13g2_decap_8 FILLER_48_362 ();
 sg13g2_decap_8 FILLER_48_369 ();
 sg13g2_decap_8 FILLER_48_376 ();
 sg13g2_decap_8 FILLER_48_383 ();
 sg13g2_decap_8 FILLER_48_390 ();
 sg13g2_decap_8 FILLER_48_397 ();
 sg13g2_decap_4 FILLER_48_404 ();
 sg13g2_fill_1 FILLER_48_408 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_7 ();
 sg13g2_decap_8 FILLER_49_14 ();
 sg13g2_decap_8 FILLER_49_21 ();
 sg13g2_decap_8 FILLER_49_28 ();
 sg13g2_decap_8 FILLER_49_35 ();
 sg13g2_decap_8 FILLER_49_42 ();
 sg13g2_decap_8 FILLER_49_49 ();
 sg13g2_decap_8 FILLER_49_56 ();
 sg13g2_decap_8 FILLER_49_63 ();
 sg13g2_decap_4 FILLER_49_70 ();
 sg13g2_fill_1 FILLER_49_117 ();
 sg13g2_decap_8 FILLER_49_156 ();
 sg13g2_decap_8 FILLER_49_163 ();
 sg13g2_decap_4 FILLER_49_218 ();
 sg13g2_fill_2 FILLER_49_241 ();
 sg13g2_fill_2 FILLER_49_275 ();
 sg13g2_fill_2 FILLER_49_311 ();
 sg13g2_fill_1 FILLER_49_313 ();
 sg13g2_decap_8 FILLER_49_370 ();
 sg13g2_decap_8 FILLER_49_377 ();
 sg13g2_decap_8 FILLER_49_384 ();
 sg13g2_decap_8 FILLER_49_391 ();
 sg13g2_decap_8 FILLER_49_398 ();
 sg13g2_decap_4 FILLER_49_405 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_8 FILLER_50_7 ();
 sg13g2_decap_8 FILLER_50_14 ();
 sg13g2_decap_8 FILLER_50_21 ();
 sg13g2_decap_8 FILLER_50_28 ();
 sg13g2_decap_8 FILLER_50_35 ();
 sg13g2_decap_8 FILLER_50_42 ();
 sg13g2_decap_8 FILLER_50_49 ();
 sg13g2_decap_8 FILLER_50_56 ();
 sg13g2_decap_8 FILLER_50_63 ();
 sg13g2_decap_8 FILLER_50_70 ();
 sg13g2_fill_2 FILLER_50_77 ();
 sg13g2_fill_1 FILLER_50_79 ();
 sg13g2_decap_4 FILLER_50_106 ();
 sg13g2_fill_2 FILLER_50_110 ();
 sg13g2_decap_4 FILLER_50_138 ();
 sg13g2_fill_2 FILLER_50_142 ();
 sg13g2_fill_2 FILLER_50_179 ();
 sg13g2_fill_1 FILLER_50_192 ();
 sg13g2_fill_2 FILLER_50_214 ();
 sg13g2_decap_4 FILLER_50_224 ();
 sg13g2_fill_2 FILLER_50_259 ();
 sg13g2_decap_8 FILLER_50_282 ();
 sg13g2_decap_8 FILLER_50_289 ();
 sg13g2_decap_8 FILLER_50_296 ();
 sg13g2_fill_1 FILLER_50_303 ();
 sg13g2_fill_2 FILLER_50_343 ();
 sg13g2_fill_1 FILLER_50_345 ();
 sg13g2_decap_8 FILLER_50_355 ();
 sg13g2_decap_8 FILLER_50_362 ();
 sg13g2_decap_8 FILLER_50_369 ();
 sg13g2_decap_8 FILLER_50_376 ();
 sg13g2_decap_8 FILLER_50_383 ();
 sg13g2_decap_8 FILLER_50_390 ();
 sg13g2_decap_8 FILLER_50_397 ();
 sg13g2_decap_4 FILLER_50_404 ();
 sg13g2_fill_1 FILLER_50_408 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_decap_8 FILLER_51_7 ();
 sg13g2_decap_8 FILLER_51_14 ();
 sg13g2_decap_8 FILLER_51_21 ();
 sg13g2_decap_8 FILLER_51_28 ();
 sg13g2_decap_8 FILLER_51_35 ();
 sg13g2_decap_8 FILLER_51_42 ();
 sg13g2_decap_8 FILLER_51_49 ();
 sg13g2_decap_8 FILLER_51_56 ();
 sg13g2_decap_8 FILLER_51_63 ();
 sg13g2_decap_8 FILLER_51_70 ();
 sg13g2_decap_4 FILLER_51_77 ();
 sg13g2_fill_1 FILLER_51_90 ();
 sg13g2_fill_2 FILLER_51_100 ();
 sg13g2_fill_1 FILLER_51_102 ();
 sg13g2_fill_1 FILLER_51_167 ();
 sg13g2_fill_2 FILLER_51_183 ();
 sg13g2_fill_1 FILLER_51_185 ();
 sg13g2_decap_8 FILLER_51_247 ();
 sg13g2_decap_4 FILLER_51_254 ();
 sg13g2_fill_1 FILLER_51_258 ();
 sg13g2_fill_2 FILLER_51_272 ();
 sg13g2_fill_1 FILLER_51_274 ();
 sg13g2_fill_2 FILLER_51_283 ();
 sg13g2_decap_8 FILLER_51_297 ();
 sg13g2_decap_8 FILLER_51_304 ();
 sg13g2_fill_2 FILLER_51_311 ();
 sg13g2_decap_8 FILLER_51_362 ();
 sg13g2_decap_8 FILLER_51_369 ();
 sg13g2_decap_8 FILLER_51_376 ();
 sg13g2_decap_8 FILLER_51_383 ();
 sg13g2_decap_8 FILLER_51_390 ();
 sg13g2_decap_8 FILLER_51_397 ();
 sg13g2_decap_4 FILLER_51_404 ();
 sg13g2_fill_1 FILLER_51_408 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_decap_8 FILLER_52_7 ();
 sg13g2_decap_8 FILLER_52_14 ();
 sg13g2_decap_8 FILLER_52_21 ();
 sg13g2_decap_8 FILLER_52_28 ();
 sg13g2_decap_8 FILLER_52_35 ();
 sg13g2_decap_8 FILLER_52_42 ();
 sg13g2_decap_8 FILLER_52_49 ();
 sg13g2_decap_8 FILLER_52_56 ();
 sg13g2_decap_8 FILLER_52_63 ();
 sg13g2_decap_8 FILLER_52_70 ();
 sg13g2_decap_8 FILLER_52_77 ();
 sg13g2_decap_8 FILLER_52_84 ();
 sg13g2_fill_2 FILLER_52_148 ();
 sg13g2_fill_1 FILLER_52_190 ();
 sg13g2_fill_2 FILLER_52_204 ();
 sg13g2_fill_2 FILLER_52_211 ();
 sg13g2_fill_1 FILLER_52_213 ();
 sg13g2_decap_8 FILLER_52_228 ();
 sg13g2_fill_2 FILLER_52_235 ();
 sg13g2_fill_1 FILLER_52_237 ();
 sg13g2_fill_1 FILLER_52_270 ();
 sg13g2_decap_8 FILLER_52_353 ();
 sg13g2_decap_8 FILLER_52_360 ();
 sg13g2_decap_8 FILLER_52_367 ();
 sg13g2_decap_8 FILLER_52_374 ();
 sg13g2_decap_8 FILLER_52_381 ();
 sg13g2_decap_8 FILLER_52_388 ();
 sg13g2_decap_8 FILLER_52_395 ();
 sg13g2_decap_8 FILLER_52_402 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_decap_8 FILLER_53_7 ();
 sg13g2_decap_8 FILLER_53_14 ();
 sg13g2_decap_8 FILLER_53_21 ();
 sg13g2_decap_8 FILLER_53_28 ();
 sg13g2_decap_8 FILLER_53_35 ();
 sg13g2_decap_8 FILLER_53_42 ();
 sg13g2_decap_8 FILLER_53_49 ();
 sg13g2_decap_8 FILLER_53_56 ();
 sg13g2_decap_8 FILLER_53_63 ();
 sg13g2_decap_8 FILLER_53_70 ();
 sg13g2_decap_8 FILLER_53_77 ();
 sg13g2_fill_2 FILLER_53_84 ();
 sg13g2_fill_1 FILLER_53_200 ();
 sg13g2_fill_1 FILLER_53_214 ();
 sg13g2_decap_4 FILLER_53_232 ();
 sg13g2_fill_1 FILLER_53_236 ();
 sg13g2_fill_2 FILLER_53_288 ();
 sg13g2_fill_1 FILLER_53_298 ();
 sg13g2_decap_8 FILLER_53_333 ();
 sg13g2_decap_8 FILLER_53_340 ();
 sg13g2_decap_8 FILLER_53_347 ();
 sg13g2_fill_2 FILLER_53_354 ();
 sg13g2_fill_1 FILLER_53_356 ();
 sg13g2_decap_8 FILLER_53_363 ();
 sg13g2_decap_8 FILLER_53_370 ();
 sg13g2_decap_8 FILLER_53_377 ();
 sg13g2_decap_8 FILLER_53_384 ();
 sg13g2_decap_8 FILLER_53_391 ();
 sg13g2_decap_8 FILLER_53_398 ();
 sg13g2_decap_4 FILLER_53_405 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_decap_8 FILLER_54_7 ();
 sg13g2_decap_8 FILLER_54_14 ();
 sg13g2_decap_8 FILLER_54_21 ();
 sg13g2_decap_8 FILLER_54_28 ();
 sg13g2_decap_8 FILLER_54_35 ();
 sg13g2_decap_8 FILLER_54_42 ();
 sg13g2_decap_8 FILLER_54_49 ();
 sg13g2_decap_8 FILLER_54_56 ();
 sg13g2_decap_8 FILLER_54_63 ();
 sg13g2_decap_8 FILLER_54_70 ();
 sg13g2_decap_4 FILLER_54_77 ();
 sg13g2_fill_2 FILLER_54_81 ();
 sg13g2_fill_1 FILLER_54_183 ();
 sg13g2_decap_4 FILLER_54_218 ();
 sg13g2_fill_1 FILLER_54_262 ();
 sg13g2_fill_1 FILLER_54_291 ();
 sg13g2_fill_2 FILLER_54_297 ();
 sg13g2_fill_2 FILLER_54_306 ();
 sg13g2_fill_1 FILLER_54_308 ();
 sg13g2_fill_2 FILLER_54_314 ();
 sg13g2_decap_4 FILLER_54_326 ();
 sg13g2_fill_1 FILLER_54_330 ();
 sg13g2_decap_8 FILLER_54_357 ();
 sg13g2_decap_8 FILLER_54_364 ();
 sg13g2_decap_8 FILLER_54_371 ();
 sg13g2_decap_8 FILLER_54_378 ();
 sg13g2_decap_8 FILLER_54_385 ();
 sg13g2_decap_8 FILLER_54_392 ();
 sg13g2_decap_8 FILLER_54_399 ();
 sg13g2_fill_2 FILLER_54_406 ();
 sg13g2_fill_1 FILLER_54_408 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_decap_8 FILLER_55_7 ();
 sg13g2_decap_8 FILLER_55_14 ();
 sg13g2_decap_8 FILLER_55_21 ();
 sg13g2_decap_8 FILLER_55_28 ();
 sg13g2_decap_8 FILLER_55_35 ();
 sg13g2_decap_8 FILLER_55_42 ();
 sg13g2_decap_8 FILLER_55_49 ();
 sg13g2_decap_8 FILLER_55_56 ();
 sg13g2_decap_8 FILLER_55_63 ();
 sg13g2_decap_8 FILLER_55_70 ();
 sg13g2_decap_8 FILLER_55_77 ();
 sg13g2_decap_8 FILLER_55_84 ();
 sg13g2_fill_2 FILLER_55_170 ();
 sg13g2_fill_1 FILLER_55_188 ();
 sg13g2_fill_2 FILLER_55_222 ();
 sg13g2_fill_1 FILLER_55_243 ();
 sg13g2_fill_2 FILLER_55_271 ();
 sg13g2_fill_1 FILLER_55_273 ();
 sg13g2_fill_2 FILLER_55_282 ();
 sg13g2_fill_1 FILLER_55_292 ();
 sg13g2_fill_2 FILLER_55_306 ();
 sg13g2_fill_2 FILLER_55_327 ();
 sg13g2_decap_8 FILLER_55_364 ();
 sg13g2_decap_8 FILLER_55_371 ();
 sg13g2_decap_8 FILLER_55_378 ();
 sg13g2_decap_8 FILLER_55_385 ();
 sg13g2_decap_8 FILLER_55_392 ();
 sg13g2_decap_8 FILLER_55_399 ();
 sg13g2_fill_2 FILLER_55_406 ();
 sg13g2_fill_1 FILLER_55_408 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_decap_8 FILLER_56_7 ();
 sg13g2_decap_8 FILLER_56_14 ();
 sg13g2_decap_8 FILLER_56_21 ();
 sg13g2_decap_8 FILLER_56_28 ();
 sg13g2_decap_8 FILLER_56_35 ();
 sg13g2_decap_8 FILLER_56_42 ();
 sg13g2_decap_8 FILLER_56_49 ();
 sg13g2_decap_8 FILLER_56_56 ();
 sg13g2_decap_8 FILLER_56_63 ();
 sg13g2_decap_8 FILLER_56_70 ();
 sg13g2_decap_8 FILLER_56_77 ();
 sg13g2_decap_8 FILLER_56_84 ();
 sg13g2_fill_2 FILLER_56_174 ();
 sg13g2_fill_2 FILLER_56_199 ();
 sg13g2_decap_8 FILLER_56_235 ();
 sg13g2_decap_8 FILLER_56_242 ();
 sg13g2_fill_2 FILLER_56_249 ();
 sg13g2_fill_2 FILLER_56_298 ();
 sg13g2_fill_2 FILLER_56_329 ();
 sg13g2_decap_8 FILLER_56_367 ();
 sg13g2_decap_8 FILLER_56_374 ();
 sg13g2_decap_8 FILLER_56_381 ();
 sg13g2_decap_8 FILLER_56_388 ();
 sg13g2_decap_8 FILLER_56_395 ();
 sg13g2_decap_8 FILLER_56_402 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_decap_8 FILLER_57_7 ();
 sg13g2_decap_8 FILLER_57_14 ();
 sg13g2_decap_8 FILLER_57_21 ();
 sg13g2_decap_8 FILLER_57_28 ();
 sg13g2_decap_8 FILLER_57_35 ();
 sg13g2_decap_8 FILLER_57_42 ();
 sg13g2_decap_8 FILLER_57_49 ();
 sg13g2_decap_8 FILLER_57_56 ();
 sg13g2_decap_8 FILLER_57_63 ();
 sg13g2_decap_8 FILLER_57_70 ();
 sg13g2_decap_8 FILLER_57_77 ();
 sg13g2_decap_8 FILLER_57_84 ();
 sg13g2_fill_2 FILLER_57_91 ();
 sg13g2_fill_2 FILLER_57_114 ();
 sg13g2_fill_1 FILLER_57_148 ();
 sg13g2_decap_4 FILLER_57_154 ();
 sg13g2_fill_1 FILLER_57_195 ();
 sg13g2_fill_2 FILLER_57_231 ();
 sg13g2_decap_8 FILLER_57_252 ();
 sg13g2_decap_4 FILLER_57_259 ();
 sg13g2_fill_1 FILLER_57_263 ();
 sg13g2_decap_8 FILLER_57_268 ();
 sg13g2_decap_8 FILLER_57_275 ();
 sg13g2_decap_4 FILLER_57_282 ();
 sg13g2_fill_1 FILLER_57_286 ();
 sg13g2_decap_8 FILLER_57_292 ();
 sg13g2_fill_1 FILLER_57_299 ();
 sg13g2_fill_2 FILLER_57_316 ();
 sg13g2_decap_8 FILLER_57_331 ();
 sg13g2_decap_8 FILLER_57_338 ();
 sg13g2_decap_8 FILLER_57_345 ();
 sg13g2_fill_1 FILLER_57_352 ();
 sg13g2_decap_8 FILLER_57_358 ();
 sg13g2_decap_8 FILLER_57_365 ();
 sg13g2_decap_8 FILLER_57_372 ();
 sg13g2_decap_8 FILLER_57_379 ();
 sg13g2_decap_8 FILLER_57_386 ();
 sg13g2_decap_8 FILLER_57_393 ();
 sg13g2_decap_8 FILLER_57_400 ();
 sg13g2_fill_2 FILLER_57_407 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_decap_8 FILLER_58_7 ();
 sg13g2_decap_8 FILLER_58_14 ();
 sg13g2_decap_8 FILLER_58_21 ();
 sg13g2_decap_8 FILLER_58_28 ();
 sg13g2_decap_8 FILLER_58_35 ();
 sg13g2_decap_8 FILLER_58_42 ();
 sg13g2_decap_8 FILLER_58_49 ();
 sg13g2_decap_8 FILLER_58_56 ();
 sg13g2_decap_8 FILLER_58_63 ();
 sg13g2_decap_8 FILLER_58_70 ();
 sg13g2_decap_8 FILLER_58_77 ();
 sg13g2_decap_4 FILLER_58_84 ();
 sg13g2_fill_1 FILLER_58_88 ();
 sg13g2_decap_4 FILLER_58_154 ();
 sg13g2_fill_2 FILLER_58_173 ();
 sg13g2_fill_2 FILLER_58_201 ();
 sg13g2_fill_1 FILLER_58_212 ();
 sg13g2_decap_8 FILLER_58_229 ();
 sg13g2_fill_1 FILLER_58_236 ();
 sg13g2_fill_1 FILLER_58_265 ();
 sg13g2_fill_1 FILLER_58_320 ();
 sg13g2_decap_8 FILLER_58_359 ();
 sg13g2_decap_8 FILLER_58_366 ();
 sg13g2_decap_8 FILLER_58_373 ();
 sg13g2_decap_8 FILLER_58_380 ();
 sg13g2_decap_8 FILLER_58_387 ();
 sg13g2_decap_8 FILLER_58_394 ();
 sg13g2_decap_8 FILLER_58_401 ();
 sg13g2_fill_1 FILLER_58_408 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_decap_8 FILLER_59_7 ();
 sg13g2_decap_8 FILLER_59_14 ();
 sg13g2_decap_8 FILLER_59_21 ();
 sg13g2_decap_8 FILLER_59_28 ();
 sg13g2_decap_8 FILLER_59_35 ();
 sg13g2_decap_8 FILLER_59_42 ();
 sg13g2_decap_8 FILLER_59_49 ();
 sg13g2_decap_8 FILLER_59_56 ();
 sg13g2_decap_8 FILLER_59_63 ();
 sg13g2_decap_8 FILLER_59_70 ();
 sg13g2_decap_8 FILLER_59_77 ();
 sg13g2_fill_2 FILLER_59_84 ();
 sg13g2_fill_1 FILLER_59_86 ();
 sg13g2_fill_1 FILLER_59_163 ();
 sg13g2_decap_4 FILLER_59_199 ();
 sg13g2_decap_8 FILLER_59_213 ();
 sg13g2_fill_1 FILLER_59_220 ();
 sg13g2_fill_2 FILLER_59_274 ();
 sg13g2_fill_1 FILLER_59_276 ();
 sg13g2_fill_2 FILLER_59_314 ();
 sg13g2_decap_8 FILLER_59_358 ();
 sg13g2_decap_8 FILLER_59_365 ();
 sg13g2_decap_8 FILLER_59_372 ();
 sg13g2_decap_8 FILLER_59_379 ();
 sg13g2_decap_8 FILLER_59_386 ();
 sg13g2_decap_8 FILLER_59_393 ();
 sg13g2_decap_8 FILLER_59_400 ();
 sg13g2_fill_2 FILLER_59_407 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_decap_8 FILLER_60_7 ();
 sg13g2_decap_8 FILLER_60_14 ();
 sg13g2_decap_8 FILLER_60_21 ();
 sg13g2_decap_8 FILLER_60_28 ();
 sg13g2_decap_8 FILLER_60_35 ();
 sg13g2_decap_8 FILLER_60_42 ();
 sg13g2_decap_8 FILLER_60_49 ();
 sg13g2_decap_8 FILLER_60_56 ();
 sg13g2_decap_8 FILLER_60_63 ();
 sg13g2_decap_8 FILLER_60_70 ();
 sg13g2_decap_8 FILLER_60_77 ();
 sg13g2_decap_4 FILLER_60_84 ();
 sg13g2_fill_1 FILLER_60_88 ();
 sg13g2_fill_1 FILLER_60_141 ();
 sg13g2_fill_1 FILLER_60_168 ();
 sg13g2_fill_1 FILLER_60_182 ();
 sg13g2_fill_1 FILLER_60_192 ();
 sg13g2_decap_8 FILLER_60_198 ();
 sg13g2_fill_1 FILLER_60_205 ();
 sg13g2_fill_2 FILLER_60_210 ();
 sg13g2_fill_1 FILLER_60_212 ();
 sg13g2_decap_4 FILLER_60_274 ();
 sg13g2_fill_2 FILLER_60_286 ();
 sg13g2_fill_1 FILLER_60_288 ();
 sg13g2_fill_2 FILLER_60_308 ();
 sg13g2_decap_8 FILLER_60_321 ();
 sg13g2_decap_4 FILLER_60_328 ();
 sg13g2_decap_8 FILLER_60_367 ();
 sg13g2_decap_8 FILLER_60_374 ();
 sg13g2_decap_8 FILLER_60_381 ();
 sg13g2_decap_8 FILLER_60_388 ();
 sg13g2_decap_8 FILLER_60_395 ();
 sg13g2_decap_8 FILLER_60_402 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_decap_8 FILLER_61_7 ();
 sg13g2_decap_8 FILLER_61_14 ();
 sg13g2_decap_8 FILLER_61_21 ();
 sg13g2_decap_8 FILLER_61_28 ();
 sg13g2_decap_8 FILLER_61_35 ();
 sg13g2_decap_8 FILLER_61_42 ();
 sg13g2_decap_8 FILLER_61_49 ();
 sg13g2_decap_8 FILLER_61_56 ();
 sg13g2_decap_8 FILLER_61_63 ();
 sg13g2_decap_8 FILLER_61_70 ();
 sg13g2_decap_8 FILLER_61_77 ();
 sg13g2_decap_8 FILLER_61_84 ();
 sg13g2_decap_4 FILLER_61_91 ();
 sg13g2_fill_1 FILLER_61_95 ();
 sg13g2_fill_2 FILLER_61_134 ();
 sg13g2_decap_8 FILLER_61_225 ();
 sg13g2_fill_2 FILLER_61_232 ();
 sg13g2_fill_1 FILLER_61_234 ();
 sg13g2_fill_2 FILLER_61_244 ();
 sg13g2_fill_1 FILLER_61_246 ();
 sg13g2_fill_2 FILLER_61_258 ();
 sg13g2_fill_1 FILLER_61_260 ();
 sg13g2_fill_2 FILLER_61_266 ();
 sg13g2_fill_2 FILLER_61_278 ();
 sg13g2_fill_1 FILLER_61_280 ();
 sg13g2_decap_4 FILLER_61_314 ();
 sg13g2_decap_8 FILLER_61_343 ();
 sg13g2_decap_8 FILLER_61_350 ();
 sg13g2_decap_8 FILLER_61_357 ();
 sg13g2_decap_8 FILLER_61_364 ();
 sg13g2_decap_8 FILLER_61_371 ();
 sg13g2_decap_8 FILLER_61_378 ();
 sg13g2_decap_8 FILLER_61_385 ();
 sg13g2_decap_8 FILLER_61_392 ();
 sg13g2_decap_8 FILLER_61_399 ();
 sg13g2_fill_2 FILLER_61_406 ();
 sg13g2_fill_1 FILLER_61_408 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_decap_8 FILLER_62_7 ();
 sg13g2_decap_8 FILLER_62_14 ();
 sg13g2_decap_8 FILLER_62_21 ();
 sg13g2_decap_8 FILLER_62_28 ();
 sg13g2_decap_8 FILLER_62_35 ();
 sg13g2_decap_8 FILLER_62_42 ();
 sg13g2_decap_8 FILLER_62_49 ();
 sg13g2_decap_8 FILLER_62_56 ();
 sg13g2_decap_8 FILLER_62_63 ();
 sg13g2_decap_8 FILLER_62_70 ();
 sg13g2_decap_8 FILLER_62_77 ();
 sg13g2_decap_8 FILLER_62_84 ();
 sg13g2_decap_8 FILLER_62_91 ();
 sg13g2_fill_2 FILLER_62_98 ();
 sg13g2_fill_1 FILLER_62_100 ();
 sg13g2_fill_1 FILLER_62_127 ();
 sg13g2_fill_1 FILLER_62_171 ();
 sg13g2_fill_2 FILLER_62_203 ();
 sg13g2_fill_2 FILLER_62_228 ();
 sg13g2_fill_1 FILLER_62_239 ();
 sg13g2_fill_2 FILLER_62_272 ();
 sg13g2_fill_1 FILLER_62_274 ();
 sg13g2_decap_8 FILLER_62_293 ();
 sg13g2_decap_4 FILLER_62_300 ();
 sg13g2_decap_4 FILLER_62_308 ();
 sg13g2_fill_1 FILLER_62_342 ();
 sg13g2_decap_8 FILLER_62_351 ();
 sg13g2_decap_8 FILLER_62_358 ();
 sg13g2_decap_8 FILLER_62_365 ();
 sg13g2_decap_8 FILLER_62_372 ();
 sg13g2_decap_8 FILLER_62_379 ();
 sg13g2_decap_8 FILLER_62_386 ();
 sg13g2_decap_8 FILLER_62_393 ();
 sg13g2_decap_8 FILLER_62_400 ();
 sg13g2_fill_2 FILLER_62_407 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_decap_8 FILLER_63_7 ();
 sg13g2_decap_8 FILLER_63_14 ();
 sg13g2_decap_8 FILLER_63_21 ();
 sg13g2_decap_8 FILLER_63_28 ();
 sg13g2_decap_8 FILLER_63_35 ();
 sg13g2_decap_8 FILLER_63_42 ();
 sg13g2_decap_8 FILLER_63_49 ();
 sg13g2_decap_8 FILLER_63_56 ();
 sg13g2_decap_8 FILLER_63_63 ();
 sg13g2_decap_8 FILLER_63_70 ();
 sg13g2_decap_8 FILLER_63_77 ();
 sg13g2_decap_8 FILLER_63_84 ();
 sg13g2_decap_8 FILLER_63_91 ();
 sg13g2_decap_8 FILLER_63_98 ();
 sg13g2_decap_4 FILLER_63_105 ();
 sg13g2_fill_1 FILLER_63_109 ();
 sg13g2_fill_2 FILLER_63_126 ();
 sg13g2_fill_2 FILLER_63_180 ();
 sg13g2_fill_1 FILLER_63_182 ();
 sg13g2_fill_1 FILLER_63_219 ();
 sg13g2_fill_2 FILLER_63_256 ();
 sg13g2_decap_8 FILLER_63_287 ();
 sg13g2_fill_2 FILLER_63_310 ();
 sg13g2_fill_1 FILLER_63_312 ();
 sg13g2_decap_8 FILLER_63_365 ();
 sg13g2_decap_8 FILLER_63_372 ();
 sg13g2_decap_8 FILLER_63_379 ();
 sg13g2_decap_8 FILLER_63_386 ();
 sg13g2_decap_8 FILLER_63_393 ();
 sg13g2_decap_8 FILLER_63_400 ();
 sg13g2_fill_2 FILLER_63_407 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_8 FILLER_64_7 ();
 sg13g2_decap_8 FILLER_64_14 ();
 sg13g2_decap_8 FILLER_64_21 ();
 sg13g2_decap_8 FILLER_64_28 ();
 sg13g2_decap_8 FILLER_64_35 ();
 sg13g2_decap_8 FILLER_64_42 ();
 sg13g2_decap_8 FILLER_64_49 ();
 sg13g2_decap_8 FILLER_64_56 ();
 sg13g2_decap_8 FILLER_64_63 ();
 sg13g2_decap_8 FILLER_64_70 ();
 sg13g2_decap_8 FILLER_64_77 ();
 sg13g2_decap_8 FILLER_64_84 ();
 sg13g2_decap_8 FILLER_64_91 ();
 sg13g2_decap_8 FILLER_64_98 ();
 sg13g2_fill_2 FILLER_64_139 ();
 sg13g2_fill_2 FILLER_64_153 ();
 sg13g2_fill_2 FILLER_64_173 ();
 sg13g2_fill_1 FILLER_64_232 ();
 sg13g2_decap_8 FILLER_64_279 ();
 sg13g2_fill_2 FILLER_64_286 ();
 sg13g2_decap_8 FILLER_64_354 ();
 sg13g2_decap_8 FILLER_64_361 ();
 sg13g2_decap_8 FILLER_64_368 ();
 sg13g2_decap_8 FILLER_64_375 ();
 sg13g2_decap_8 FILLER_64_382 ();
 sg13g2_decap_8 FILLER_64_389 ();
 sg13g2_decap_8 FILLER_64_396 ();
 sg13g2_decap_4 FILLER_64_403 ();
 sg13g2_fill_2 FILLER_64_407 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_8 FILLER_65_7 ();
 sg13g2_decap_8 FILLER_65_14 ();
 sg13g2_decap_8 FILLER_65_21 ();
 sg13g2_decap_8 FILLER_65_28 ();
 sg13g2_decap_8 FILLER_65_35 ();
 sg13g2_decap_8 FILLER_65_42 ();
 sg13g2_decap_8 FILLER_65_49 ();
 sg13g2_decap_8 FILLER_65_56 ();
 sg13g2_decap_8 FILLER_65_63 ();
 sg13g2_decap_8 FILLER_65_70 ();
 sg13g2_decap_8 FILLER_65_77 ();
 sg13g2_decap_8 FILLER_65_84 ();
 sg13g2_decap_8 FILLER_65_91 ();
 sg13g2_fill_2 FILLER_65_98 ();
 sg13g2_fill_2 FILLER_65_142 ();
 sg13g2_fill_2 FILLER_65_149 ();
 sg13g2_fill_1 FILLER_65_151 ();
 sg13g2_decap_8 FILLER_65_158 ();
 sg13g2_decap_4 FILLER_65_165 ();
 sg13g2_fill_1 FILLER_65_169 ();
 sg13g2_decap_8 FILLER_65_175 ();
 sg13g2_fill_2 FILLER_65_201 ();
 sg13g2_decap_8 FILLER_65_264 ();
 sg13g2_decap_4 FILLER_65_271 ();
 sg13g2_fill_1 FILLER_65_275 ();
 sg13g2_fill_2 FILLER_65_293 ();
 sg13g2_fill_1 FILLER_65_307 ();
 sg13g2_fill_1 FILLER_65_327 ();
 sg13g2_decap_8 FILLER_65_354 ();
 sg13g2_decap_8 FILLER_65_361 ();
 sg13g2_decap_8 FILLER_65_368 ();
 sg13g2_decap_8 FILLER_65_375 ();
 sg13g2_decap_8 FILLER_65_382 ();
 sg13g2_decap_8 FILLER_65_389 ();
 sg13g2_decap_8 FILLER_65_396 ();
 sg13g2_decap_4 FILLER_65_403 ();
 sg13g2_fill_2 FILLER_65_407 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_8 FILLER_66_7 ();
 sg13g2_decap_8 FILLER_66_14 ();
 sg13g2_decap_8 FILLER_66_21 ();
 sg13g2_decap_8 FILLER_66_28 ();
 sg13g2_decap_8 FILLER_66_35 ();
 sg13g2_decap_8 FILLER_66_42 ();
 sg13g2_decap_8 FILLER_66_49 ();
 sg13g2_decap_8 FILLER_66_56 ();
 sg13g2_decap_8 FILLER_66_63 ();
 sg13g2_decap_8 FILLER_66_70 ();
 sg13g2_decap_8 FILLER_66_77 ();
 sg13g2_decap_8 FILLER_66_84 ();
 sg13g2_fill_2 FILLER_66_91 ();
 sg13g2_fill_1 FILLER_66_93 ();
 sg13g2_fill_2 FILLER_66_154 ();
 sg13g2_fill_1 FILLER_66_156 ();
 sg13g2_decap_8 FILLER_66_161 ();
 sg13g2_decap_8 FILLER_66_168 ();
 sg13g2_decap_8 FILLER_66_175 ();
 sg13g2_fill_2 FILLER_66_182 ();
 sg13g2_fill_1 FILLER_66_197 ();
 sg13g2_decap_8 FILLER_66_254 ();
 sg13g2_decap_8 FILLER_66_261 ();
 sg13g2_decap_4 FILLER_66_268 ();
 sg13g2_fill_2 FILLER_66_272 ();
 sg13g2_decap_8 FILLER_66_295 ();
 sg13g2_fill_2 FILLER_66_302 ();
 sg13g2_decap_8 FILLER_66_331 ();
 sg13g2_decap_8 FILLER_66_338 ();
 sg13g2_decap_8 FILLER_66_345 ();
 sg13g2_decap_8 FILLER_66_352 ();
 sg13g2_decap_8 FILLER_66_359 ();
 sg13g2_decap_8 FILLER_66_366 ();
 sg13g2_decap_8 FILLER_66_373 ();
 sg13g2_decap_8 FILLER_66_380 ();
 sg13g2_decap_8 FILLER_66_387 ();
 sg13g2_decap_8 FILLER_66_394 ();
 sg13g2_decap_8 FILLER_66_401 ();
 sg13g2_fill_1 FILLER_66_408 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_8 FILLER_67_7 ();
 sg13g2_decap_8 FILLER_67_14 ();
 sg13g2_decap_8 FILLER_67_21 ();
 sg13g2_decap_8 FILLER_67_28 ();
 sg13g2_decap_8 FILLER_67_35 ();
 sg13g2_decap_8 FILLER_67_42 ();
 sg13g2_decap_8 FILLER_67_49 ();
 sg13g2_decap_8 FILLER_67_56 ();
 sg13g2_decap_8 FILLER_67_63 ();
 sg13g2_decap_8 FILLER_67_70 ();
 sg13g2_decap_8 FILLER_67_77 ();
 sg13g2_decap_4 FILLER_67_84 ();
 sg13g2_fill_2 FILLER_67_132 ();
 sg13g2_fill_2 FILLER_67_286 ();
 sg13g2_decap_8 FILLER_67_328 ();
 sg13g2_decap_8 FILLER_67_335 ();
 sg13g2_decap_8 FILLER_67_342 ();
 sg13g2_decap_8 FILLER_67_355 ();
 sg13g2_decap_8 FILLER_67_362 ();
 sg13g2_decap_8 FILLER_67_369 ();
 sg13g2_decap_8 FILLER_67_376 ();
 sg13g2_decap_8 FILLER_67_383 ();
 sg13g2_decap_8 FILLER_67_390 ();
 sg13g2_decap_8 FILLER_67_397 ();
 sg13g2_decap_4 FILLER_67_404 ();
 sg13g2_fill_1 FILLER_67_408 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_8 FILLER_68_7 ();
 sg13g2_decap_8 FILLER_68_14 ();
 sg13g2_decap_8 FILLER_68_21 ();
 sg13g2_decap_8 FILLER_68_28 ();
 sg13g2_decap_8 FILLER_68_35 ();
 sg13g2_decap_8 FILLER_68_42 ();
 sg13g2_decap_8 FILLER_68_49 ();
 sg13g2_decap_8 FILLER_68_56 ();
 sg13g2_decap_8 FILLER_68_63 ();
 sg13g2_decap_8 FILLER_68_70 ();
 sg13g2_decap_8 FILLER_68_77 ();
 sg13g2_decap_4 FILLER_68_84 ();
 sg13g2_fill_1 FILLER_68_88 ();
 sg13g2_fill_1 FILLER_68_126 ();
 sg13g2_fill_1 FILLER_68_267 ();
 sg13g2_fill_2 FILLER_68_281 ();
 sg13g2_fill_2 FILLER_68_314 ();
 sg13g2_fill_1 FILLER_68_316 ();
 sg13g2_decap_8 FILLER_68_363 ();
 sg13g2_decap_8 FILLER_68_370 ();
 sg13g2_decap_8 FILLER_68_377 ();
 sg13g2_decap_8 FILLER_68_384 ();
 sg13g2_decap_8 FILLER_68_391 ();
 sg13g2_decap_8 FILLER_68_398 ();
 sg13g2_decap_4 FILLER_68_405 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_8 FILLER_69_7 ();
 sg13g2_decap_8 FILLER_69_14 ();
 sg13g2_decap_8 FILLER_69_21 ();
 sg13g2_decap_8 FILLER_69_28 ();
 sg13g2_decap_8 FILLER_69_35 ();
 sg13g2_decap_8 FILLER_69_42 ();
 sg13g2_decap_8 FILLER_69_49 ();
 sg13g2_decap_8 FILLER_69_56 ();
 sg13g2_decap_8 FILLER_69_63 ();
 sg13g2_decap_8 FILLER_69_70 ();
 sg13g2_decap_8 FILLER_69_77 ();
 sg13g2_fill_2 FILLER_69_84 ();
 sg13g2_fill_2 FILLER_69_123 ();
 sg13g2_fill_1 FILLER_69_141 ();
 sg13g2_fill_2 FILLER_69_186 ();
 sg13g2_fill_1 FILLER_69_188 ();
 sg13g2_decap_4 FILLER_69_197 ();
 sg13g2_fill_1 FILLER_69_201 ();
 sg13g2_fill_2 FILLER_69_248 ();
 sg13g2_fill_2 FILLER_69_276 ();
 sg13g2_fill_1 FILLER_69_278 ();
 sg13g2_decap_4 FILLER_69_336 ();
 sg13g2_fill_1 FILLER_69_340 ();
 sg13g2_decap_8 FILLER_69_355 ();
 sg13g2_decap_8 FILLER_69_362 ();
 sg13g2_decap_8 FILLER_69_369 ();
 sg13g2_decap_8 FILLER_69_376 ();
 sg13g2_decap_8 FILLER_69_383 ();
 sg13g2_decap_8 FILLER_69_390 ();
 sg13g2_decap_8 FILLER_69_397 ();
 sg13g2_decap_4 FILLER_69_404 ();
 sg13g2_fill_1 FILLER_69_408 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_decap_8 FILLER_70_14 ();
 sg13g2_decap_8 FILLER_70_21 ();
 sg13g2_decap_8 FILLER_70_28 ();
 sg13g2_decap_8 FILLER_70_35 ();
 sg13g2_decap_8 FILLER_70_42 ();
 sg13g2_decap_8 FILLER_70_49 ();
 sg13g2_decap_8 FILLER_70_56 ();
 sg13g2_decap_8 FILLER_70_63 ();
 sg13g2_decap_8 FILLER_70_70 ();
 sg13g2_decap_8 FILLER_70_77 ();
 sg13g2_fill_2 FILLER_70_133 ();
 sg13g2_fill_1 FILLER_70_139 ();
 sg13g2_decap_4 FILLER_70_144 ();
 sg13g2_fill_1 FILLER_70_148 ();
 sg13g2_fill_1 FILLER_70_158 ();
 sg13g2_fill_2 FILLER_70_189 ();
 sg13g2_decap_8 FILLER_70_197 ();
 sg13g2_fill_2 FILLER_70_204 ();
 sg13g2_fill_2 FILLER_70_220 ();
 sg13g2_fill_2 FILLER_70_266 ();
 sg13g2_fill_2 FILLER_70_277 ();
 sg13g2_fill_1 FILLER_70_298 ();
 sg13g2_decap_8 FILLER_70_343 ();
 sg13g2_decap_8 FILLER_70_350 ();
 sg13g2_decap_8 FILLER_70_357 ();
 sg13g2_decap_8 FILLER_70_364 ();
 sg13g2_decap_8 FILLER_70_371 ();
 sg13g2_decap_8 FILLER_70_378 ();
 sg13g2_decap_8 FILLER_70_385 ();
 sg13g2_decap_8 FILLER_70_392 ();
 sg13g2_decap_8 FILLER_70_399 ();
 sg13g2_fill_2 FILLER_70_406 ();
 sg13g2_fill_1 FILLER_70_408 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_decap_8 FILLER_71_7 ();
 sg13g2_decap_8 FILLER_71_14 ();
 sg13g2_decap_8 FILLER_71_21 ();
 sg13g2_decap_8 FILLER_71_28 ();
 sg13g2_decap_8 FILLER_71_35 ();
 sg13g2_decap_8 FILLER_71_42 ();
 sg13g2_decap_8 FILLER_71_49 ();
 sg13g2_decap_8 FILLER_71_56 ();
 sg13g2_decap_8 FILLER_71_63 ();
 sg13g2_decap_8 FILLER_71_70 ();
 sg13g2_decap_4 FILLER_71_77 ();
 sg13g2_fill_1 FILLER_71_107 ();
 sg13g2_decap_4 FILLER_71_143 ();
 sg13g2_fill_2 FILLER_71_147 ();
 sg13g2_fill_2 FILLER_71_181 ();
 sg13g2_fill_1 FILLER_71_183 ();
 sg13g2_fill_1 FILLER_71_235 ();
 sg13g2_fill_1 FILLER_71_253 ();
 sg13g2_fill_1 FILLER_71_285 ();
 sg13g2_fill_2 FILLER_71_300 ();
 sg13g2_decap_8 FILLER_71_341 ();
 sg13g2_decap_8 FILLER_71_348 ();
 sg13g2_decap_8 FILLER_71_355 ();
 sg13g2_decap_8 FILLER_71_362 ();
 sg13g2_decap_8 FILLER_71_369 ();
 sg13g2_decap_8 FILLER_71_376 ();
 sg13g2_decap_8 FILLER_71_383 ();
 sg13g2_decap_8 FILLER_71_390 ();
 sg13g2_decap_8 FILLER_71_397 ();
 sg13g2_decap_4 FILLER_71_404 ();
 sg13g2_fill_1 FILLER_71_408 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_decap_8 FILLER_72_14 ();
 sg13g2_decap_8 FILLER_72_21 ();
 sg13g2_decap_8 FILLER_72_28 ();
 sg13g2_decap_8 FILLER_72_35 ();
 sg13g2_decap_8 FILLER_72_42 ();
 sg13g2_decap_8 FILLER_72_49 ();
 sg13g2_decap_8 FILLER_72_56 ();
 sg13g2_decap_8 FILLER_72_63 ();
 sg13g2_decap_8 FILLER_72_70 ();
 sg13g2_fill_1 FILLER_72_133 ();
 sg13g2_fill_2 FILLER_72_146 ();
 sg13g2_fill_1 FILLER_72_148 ();
 sg13g2_fill_2 FILLER_72_158 ();
 sg13g2_fill_2 FILLER_72_165 ();
 sg13g2_fill_1 FILLER_72_173 ();
 sg13g2_fill_1 FILLER_72_234 ();
 sg13g2_decap_8 FILLER_72_331 ();
 sg13g2_fill_2 FILLER_72_338 ();
 sg13g2_decap_8 FILLER_72_345 ();
 sg13g2_decap_8 FILLER_72_352 ();
 sg13g2_decap_8 FILLER_72_359 ();
 sg13g2_decap_8 FILLER_72_366 ();
 sg13g2_decap_8 FILLER_72_373 ();
 sg13g2_decap_8 FILLER_72_380 ();
 sg13g2_decap_8 FILLER_72_387 ();
 sg13g2_decap_8 FILLER_72_394 ();
 sg13g2_decap_8 FILLER_72_401 ();
 sg13g2_fill_1 FILLER_72_408 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_decap_8 FILLER_73_14 ();
 sg13g2_decap_8 FILLER_73_21 ();
 sg13g2_decap_8 FILLER_73_28 ();
 sg13g2_decap_8 FILLER_73_35 ();
 sg13g2_decap_8 FILLER_73_42 ();
 sg13g2_decap_8 FILLER_73_49 ();
 sg13g2_decap_8 FILLER_73_56 ();
 sg13g2_decap_8 FILLER_73_63 ();
 sg13g2_decap_8 FILLER_73_70 ();
 sg13g2_fill_1 FILLER_73_77 ();
 sg13g2_fill_1 FILLER_73_189 ();
 sg13g2_fill_2 FILLER_73_230 ();
 sg13g2_fill_1 FILLER_73_293 ();
 sg13g2_decap_8 FILLER_73_353 ();
 sg13g2_decap_8 FILLER_73_360 ();
 sg13g2_decap_8 FILLER_73_367 ();
 sg13g2_decap_8 FILLER_73_374 ();
 sg13g2_decap_8 FILLER_73_381 ();
 sg13g2_decap_8 FILLER_73_388 ();
 sg13g2_decap_8 FILLER_73_395 ();
 sg13g2_decap_8 FILLER_73_402 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_decap_8 FILLER_74_14 ();
 sg13g2_decap_8 FILLER_74_21 ();
 sg13g2_decap_8 FILLER_74_28 ();
 sg13g2_decap_8 FILLER_74_35 ();
 sg13g2_decap_8 FILLER_74_42 ();
 sg13g2_decap_8 FILLER_74_49 ();
 sg13g2_decap_8 FILLER_74_56 ();
 sg13g2_decap_8 FILLER_74_63 ();
 sg13g2_decap_4 FILLER_74_70 ();
 sg13g2_fill_2 FILLER_74_74 ();
 sg13g2_fill_1 FILLER_74_167 ();
 sg13g2_fill_1 FILLER_74_214 ();
 sg13g2_fill_1 FILLER_74_315 ();
 sg13g2_decap_8 FILLER_74_347 ();
 sg13g2_decap_8 FILLER_74_354 ();
 sg13g2_decap_8 FILLER_74_361 ();
 sg13g2_decap_8 FILLER_74_368 ();
 sg13g2_decap_8 FILLER_74_375 ();
 sg13g2_decap_8 FILLER_74_382 ();
 sg13g2_decap_8 FILLER_74_389 ();
 sg13g2_decap_8 FILLER_74_396 ();
 sg13g2_decap_4 FILLER_74_403 ();
 sg13g2_fill_2 FILLER_74_407 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_14 ();
 sg13g2_decap_8 FILLER_75_21 ();
 sg13g2_decap_8 FILLER_75_28 ();
 sg13g2_decap_8 FILLER_75_35 ();
 sg13g2_decap_8 FILLER_75_42 ();
 sg13g2_decap_8 FILLER_75_49 ();
 sg13g2_decap_8 FILLER_75_56 ();
 sg13g2_decap_8 FILLER_75_63 ();
 sg13g2_decap_8 FILLER_75_70 ();
 sg13g2_fill_2 FILLER_75_77 ();
 sg13g2_fill_2 FILLER_75_96 ();
 sg13g2_fill_1 FILLER_75_98 ();
 sg13g2_fill_1 FILLER_75_155 ();
 sg13g2_fill_2 FILLER_75_206 ();
 sg13g2_fill_2 FILLER_75_221 ();
 sg13g2_fill_2 FILLER_75_253 ();
 sg13g2_decap_8 FILLER_75_327 ();
 sg13g2_decap_8 FILLER_75_334 ();
 sg13g2_decap_8 FILLER_75_341 ();
 sg13g2_decap_8 FILLER_75_348 ();
 sg13g2_decap_8 FILLER_75_355 ();
 sg13g2_decap_8 FILLER_75_362 ();
 sg13g2_decap_8 FILLER_75_369 ();
 sg13g2_decap_8 FILLER_75_376 ();
 sg13g2_decap_8 FILLER_75_383 ();
 sg13g2_decap_8 FILLER_75_390 ();
 sg13g2_decap_8 FILLER_75_397 ();
 sg13g2_decap_4 FILLER_75_404 ();
 sg13g2_fill_1 FILLER_75_408 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_8 FILLER_76_21 ();
 sg13g2_decap_8 FILLER_76_28 ();
 sg13g2_decap_8 FILLER_76_35 ();
 sg13g2_decap_8 FILLER_76_42 ();
 sg13g2_decap_8 FILLER_76_49 ();
 sg13g2_decap_8 FILLER_76_56 ();
 sg13g2_decap_8 FILLER_76_63 ();
 sg13g2_fill_1 FILLER_76_246 ();
 sg13g2_decap_8 FILLER_76_329 ();
 sg13g2_decap_8 FILLER_76_336 ();
 sg13g2_decap_8 FILLER_76_343 ();
 sg13g2_decap_8 FILLER_76_350 ();
 sg13g2_decap_8 FILLER_76_357 ();
 sg13g2_decap_8 FILLER_76_364 ();
 sg13g2_decap_8 FILLER_76_371 ();
 sg13g2_decap_8 FILLER_76_378 ();
 sg13g2_decap_8 FILLER_76_385 ();
 sg13g2_decap_8 FILLER_76_392 ();
 sg13g2_decap_8 FILLER_76_399 ();
 sg13g2_fill_2 FILLER_76_406 ();
 sg13g2_fill_1 FILLER_76_408 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_decap_8 FILLER_77_28 ();
 sg13g2_decap_8 FILLER_77_35 ();
 sg13g2_decap_8 FILLER_77_42 ();
 sg13g2_decap_8 FILLER_77_49 ();
 sg13g2_decap_8 FILLER_77_56 ();
 sg13g2_fill_2 FILLER_77_182 ();
 sg13g2_fill_1 FILLER_77_216 ();
 sg13g2_fill_1 FILLER_77_292 ();
 sg13g2_decap_8 FILLER_77_334 ();
 sg13g2_decap_8 FILLER_77_341 ();
 sg13g2_decap_8 FILLER_77_348 ();
 sg13g2_decap_8 FILLER_77_355 ();
 sg13g2_decap_8 FILLER_77_362 ();
 sg13g2_decap_8 FILLER_77_369 ();
 sg13g2_decap_8 FILLER_77_376 ();
 sg13g2_decap_8 FILLER_77_383 ();
 sg13g2_decap_8 FILLER_77_390 ();
 sg13g2_decap_8 FILLER_77_397 ();
 sg13g2_decap_4 FILLER_77_404 ();
 sg13g2_fill_1 FILLER_77_408 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_decap_8 FILLER_78_28 ();
 sg13g2_decap_8 FILLER_78_35 ();
 sg13g2_decap_8 FILLER_78_42 ();
 sg13g2_decap_8 FILLER_78_49 ();
 sg13g2_decap_8 FILLER_78_56 ();
 sg13g2_decap_8 FILLER_78_63 ();
 sg13g2_fill_2 FILLER_78_70 ();
 sg13g2_fill_1 FILLER_78_72 ();
 sg13g2_fill_1 FILLER_78_107 ();
 sg13g2_fill_1 FILLER_78_242 ();
 sg13g2_decap_8 FILLER_78_340 ();
 sg13g2_decap_8 FILLER_78_347 ();
 sg13g2_decap_8 FILLER_78_354 ();
 sg13g2_decap_8 FILLER_78_361 ();
 sg13g2_decap_8 FILLER_78_368 ();
 sg13g2_decap_8 FILLER_78_375 ();
 sg13g2_decap_8 FILLER_78_382 ();
 sg13g2_decap_8 FILLER_78_389 ();
 sg13g2_decap_8 FILLER_78_396 ();
 sg13g2_decap_4 FILLER_78_403 ();
 sg13g2_fill_2 FILLER_78_407 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_decap_8 FILLER_79_35 ();
 sg13g2_decap_8 FILLER_79_42 ();
 sg13g2_decap_8 FILLER_79_49 ();
 sg13g2_decap_4 FILLER_79_56 ();
 sg13g2_fill_2 FILLER_79_119 ();
 sg13g2_fill_1 FILLER_79_121 ();
 sg13g2_fill_2 FILLER_79_214 ();
 sg13g2_decap_8 FILLER_79_330 ();
 sg13g2_decap_8 FILLER_79_337 ();
 sg13g2_decap_8 FILLER_79_344 ();
 sg13g2_decap_8 FILLER_79_351 ();
 sg13g2_decap_8 FILLER_79_358 ();
 sg13g2_decap_8 FILLER_79_365 ();
 sg13g2_decap_8 FILLER_79_372 ();
 sg13g2_decap_8 FILLER_79_379 ();
 sg13g2_decap_8 FILLER_79_386 ();
 sg13g2_decap_8 FILLER_79_393 ();
 sg13g2_decap_8 FILLER_79_400 ();
 sg13g2_fill_2 FILLER_79_407 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_42 ();
 sg13g2_fill_1 FILLER_80_49 ();
 sg13g2_fill_2 FILLER_80_122 ();
 sg13g2_fill_1 FILLER_80_124 ();
 sg13g2_fill_1 FILLER_80_148 ();
 sg13g2_fill_2 FILLER_80_154 ();
 sg13g2_fill_1 FILLER_80_232 ();
 sg13g2_fill_1 FILLER_80_238 ();
 sg13g2_fill_1 FILLER_80_298 ();
 sg13g2_decap_8 FILLER_80_317 ();
 sg13g2_decap_8 FILLER_80_324 ();
 sg13g2_decap_8 FILLER_80_331 ();
 sg13g2_decap_8 FILLER_80_338 ();
 sg13g2_decap_8 FILLER_80_345 ();
 sg13g2_decap_8 FILLER_80_352 ();
 sg13g2_fill_1 FILLER_80_359 ();
 sg13g2_fill_2 FILLER_80_365 ();
 sg13g2_fill_1 FILLER_80_367 ();
 sg13g2_decap_8 FILLER_80_373 ();
 sg13g2_decap_8 FILLER_80_380 ();
 sg13g2_decap_8 FILLER_80_387 ();
 sg13g2_decap_8 FILLER_80_394 ();
 sg13g2_decap_8 FILLER_80_401 ();
 sg13g2_fill_1 FILLER_80_408 ();
 assign uio_oe[0] = net3;
 assign uio_oe[1] = net4;
 assign uio_oe[2] = net5;
 assign uio_oe[3] = net6;
 assign uio_oe[4] = net7;
 assign uio_oe[5] = net8;
 assign uio_oe[6] = net9;
 assign uio_oe[7] = net10;
 assign uio_out[0] = net11;
 assign uio_out[1] = net12;
 assign uio_out[2] = net13;
 assign uio_out[3] = net14;
 assign uio_out[4] = net15;
 assign uio_out[5] = net16;
 assign uio_out[6] = net17;
 assign uio_out[7] = net18;
endmodule

module tt_um_uart_bgdtanasa (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire clk_out;
 wire \clk_out_cnt[0] ;
 wire \clk_out_cnt[1] ;
 wire \clk_out_cnt[2] ;
 wire \clk_out_cnt[3] ;
 wire \fifo_d[0][0] ;
 wire \fifo_d[0][1] ;
 wire \fifo_d[0][2] ;
 wire \fifo_d[0][3] ;
 wire \fifo_d[0][4] ;
 wire \fifo_d[0][5] ;
 wire \fifo_d[0][6] ;
 wire \fifo_d[0][7] ;
 wire \fifo_d[10][0] ;
 wire \fifo_d[10][1] ;
 wire \fifo_d[10][2] ;
 wire \fifo_d[10][3] ;
 wire \fifo_d[10][4] ;
 wire \fifo_d[10][5] ;
 wire \fifo_d[10][6] ;
 wire \fifo_d[10][7] ;
 wire \fifo_d[11][0] ;
 wire \fifo_d[11][1] ;
 wire \fifo_d[11][2] ;
 wire \fifo_d[11][3] ;
 wire \fifo_d[11][4] ;
 wire \fifo_d[11][5] ;
 wire \fifo_d[11][6] ;
 wire \fifo_d[11][7] ;
 wire \fifo_d[12][0] ;
 wire \fifo_d[12][1] ;
 wire \fifo_d[12][2] ;
 wire \fifo_d[12][3] ;
 wire \fifo_d[12][4] ;
 wire \fifo_d[12][5] ;
 wire \fifo_d[12][6] ;
 wire \fifo_d[12][7] ;
 wire \fifo_d[13][0] ;
 wire \fifo_d[13][1] ;
 wire \fifo_d[13][2] ;
 wire \fifo_d[13][3] ;
 wire \fifo_d[13][4] ;
 wire \fifo_d[13][5] ;
 wire \fifo_d[13][6] ;
 wire \fifo_d[13][7] ;
 wire \fifo_d[14][0] ;
 wire \fifo_d[14][1] ;
 wire \fifo_d[14][2] ;
 wire \fifo_d[14][3] ;
 wire \fifo_d[14][4] ;
 wire \fifo_d[14][5] ;
 wire \fifo_d[14][6] ;
 wire \fifo_d[14][7] ;
 wire \fifo_d[15][0] ;
 wire \fifo_d[15][1] ;
 wire \fifo_d[15][2] ;
 wire \fifo_d[15][3] ;
 wire \fifo_d[15][4] ;
 wire \fifo_d[15][5] ;
 wire \fifo_d[15][6] ;
 wire \fifo_d[15][7] ;
 wire \fifo_d[1][0] ;
 wire \fifo_d[1][1] ;
 wire \fifo_d[1][2] ;
 wire \fifo_d[1][3] ;
 wire \fifo_d[1][4] ;
 wire \fifo_d[1][5] ;
 wire \fifo_d[1][6] ;
 wire \fifo_d[1][7] ;
 wire \fifo_d[2][0] ;
 wire \fifo_d[2][1] ;
 wire \fifo_d[2][2] ;
 wire \fifo_d[2][3] ;
 wire \fifo_d[2][4] ;
 wire \fifo_d[2][5] ;
 wire \fifo_d[2][6] ;
 wire \fifo_d[2][7] ;
 wire \fifo_d[3][0] ;
 wire \fifo_d[3][1] ;
 wire \fifo_d[3][2] ;
 wire \fifo_d[3][3] ;
 wire \fifo_d[3][4] ;
 wire \fifo_d[3][5] ;
 wire \fifo_d[3][6] ;
 wire \fifo_d[3][7] ;
 wire \fifo_d[4][0] ;
 wire \fifo_d[4][1] ;
 wire \fifo_d[4][2] ;
 wire \fifo_d[4][3] ;
 wire \fifo_d[4][4] ;
 wire \fifo_d[4][5] ;
 wire \fifo_d[4][6] ;
 wire \fifo_d[4][7] ;
 wire \fifo_d[5][0] ;
 wire \fifo_d[5][1] ;
 wire \fifo_d[5][2] ;
 wire \fifo_d[5][3] ;
 wire \fifo_d[5][4] ;
 wire \fifo_d[5][5] ;
 wire \fifo_d[5][6] ;
 wire \fifo_d[5][7] ;
 wire \fifo_d[6][0] ;
 wire \fifo_d[6][1] ;
 wire \fifo_d[6][2] ;
 wire \fifo_d[6][3] ;
 wire \fifo_d[6][4] ;
 wire \fifo_d[6][5] ;
 wire \fifo_d[6][6] ;
 wire \fifo_d[6][7] ;
 wire \fifo_d[7][0] ;
 wire \fifo_d[7][1] ;
 wire \fifo_d[7][2] ;
 wire \fifo_d[7][3] ;
 wire \fifo_d[7][4] ;
 wire \fifo_d[7][5] ;
 wire \fifo_d[7][6] ;
 wire \fifo_d[7][7] ;
 wire \fifo_d[8][0] ;
 wire \fifo_d[8][1] ;
 wire \fifo_d[8][2] ;
 wire \fifo_d[8][3] ;
 wire \fifo_d[8][4] ;
 wire \fifo_d[8][5] ;
 wire \fifo_d[8][6] ;
 wire \fifo_d[8][7] ;
 wire \fifo_d[9][0] ;
 wire \fifo_d[9][1] ;
 wire \fifo_d[9][2] ;
 wire \fifo_d[9][3] ;
 wire \fifo_d[9][4] ;
 wire \fifo_d[9][5] ;
 wire \fifo_d[9][6] ;
 wire \fifo_d[9][7] ;
 wire \fifo_h[0] ;
 wire \fifo_h[1] ;
 wire \fifo_h[2] ;
 wire \fifo_h[3] ;
 wire \fifo_t[0] ;
 wire \fifo_t[1] ;
 wire \fifo_t[2] ;
 wire \fifo_t[3] ;
 wire rx_data_ready;
 wire rx_sample_clk;
 wire \tx_data[0] ;
 wire \tx_data[1] ;
 wire \tx_data[2] ;
 wire \tx_data[3] ;
 wire \tx_data[4] ;
 wire \tx_data[5] ;
 wire \tx_data[6] ;
 wire \tx_data[7] ;
 wire tx_data_done;
 wire tx_data_out;
 wire tx_do;
 wire \uart_0.rx.rx_data_in ;
 wire \uart_0.rx.rx_marker[0] ;
 wire \uart_0.rx.rx_marker[1] ;
 wire \uart_0.rx.rx_marker[2] ;
 wire \uart_0.rx.rx_marker[3] ;
 wire \uart_0.rx.rx_marker[4] ;
 wire \uart_0.rx.rx_marker[5] ;
 wire \uart_0.rx.rx_marker[6] ;
 wire \uart_0.rx.rx_sample_clk_cnt[0] ;
 wire \uart_0.rx.rx_sample_clk_cnt[1] ;
 wire \uart_0.rx.rx_sample_clk_cnt[2] ;
 wire \uart_0.rx.rx_sample_clk_cnt[3] ;
 wire \uart_0.rx.rx_sample_clk_cnt[4] ;
 wire \uart_0.rx.rx_sample_clk_cnt[5] ;
 wire \uart_0.rx.rx_sample_clk_cnt[6] ;
 wire \uart_0.rx.rx_sample_cnt[0] ;
 wire \uart_0.rx.rx_sample_cnt[1] ;
 wire \uart_0.rx.rx_sample_cnt[2] ;
 wire \uart_0.rx.rx_sample_cnt[3] ;
 wire \uart_0.rx.rx_sample_cnt[4] ;
 wire \uart_0.rx.rx_sample_cnt[5] ;
 wire \uart_0.rx.rx_sample_cnt[6] ;
 wire \uart_0.rx.rx_sample_wrap[0] ;
 wire \uart_0.rx.rx_sample_wrap[3] ;
 wire \uart_0.rx.rx_samples[0] ;
 wire \uart_0.rx.rx_samples[10] ;
 wire \uart_0.rx.rx_samples[11] ;
 wire \uart_0.rx.rx_samples[12] ;
 wire \uart_0.rx.rx_samples[13] ;
 wire \uart_0.rx.rx_samples[14] ;
 wire \uart_0.rx.rx_samples[15] ;
 wire \uart_0.rx.rx_samples[16] ;
 wire \uart_0.rx.rx_samples[17] ;
 wire \uart_0.rx.rx_samples[18] ;
 wire \uart_0.rx.rx_samples[19] ;
 wire \uart_0.rx.rx_samples[1] ;
 wire \uart_0.rx.rx_samples[20] ;
 wire \uart_0.rx.rx_samples[21] ;
 wire \uart_0.rx.rx_samples[22] ;
 wire \uart_0.rx.rx_samples[23] ;
 wire \uart_0.rx.rx_samples[24] ;
 wire \uart_0.rx.rx_samples[25] ;
 wire \uart_0.rx.rx_samples[26] ;
 wire \uart_0.rx.rx_samples[27] ;
 wire \uart_0.rx.rx_samples[28] ;
 wire \uart_0.rx.rx_samples[29] ;
 wire \uart_0.rx.rx_samples[2] ;
 wire \uart_0.rx.rx_samples[30] ;
 wire \uart_0.rx.rx_samples[31] ;
 wire \uart_0.rx.rx_samples[32] ;
 wire \uart_0.rx.rx_samples[33] ;
 wire \uart_0.rx.rx_samples[34] ;
 wire \uart_0.rx.rx_samples[35] ;
 wire \uart_0.rx.rx_samples[36] ;
 wire \uart_0.rx.rx_samples[37] ;
 wire \uart_0.rx.rx_samples[38] ;
 wire \uart_0.rx.rx_samples[39] ;
 wire \uart_0.rx.rx_samples[3] ;
 wire \uart_0.rx.rx_samples[40] ;
 wire \uart_0.rx.rx_samples[41] ;
 wire \uart_0.rx.rx_samples[42] ;
 wire \uart_0.rx.rx_samples[43] ;
 wire \uart_0.rx.rx_samples[44] ;
 wire \uart_0.rx.rx_samples[45] ;
 wire \uart_0.rx.rx_samples[46] ;
 wire \uart_0.rx.rx_samples[47] ;
 wire \uart_0.rx.rx_samples[48] ;
 wire \uart_0.rx.rx_samples[49] ;
 wire \uart_0.rx.rx_samples[4] ;
 wire \uart_0.rx.rx_samples[50] ;
 wire \uart_0.rx.rx_samples[51] ;
 wire \uart_0.rx.rx_samples[52] ;
 wire \uart_0.rx.rx_samples[53] ;
 wire \uart_0.rx.rx_samples[54] ;
 wire \uart_0.rx.rx_samples[55] ;
 wire \uart_0.rx.rx_samples[56] ;
 wire \uart_0.rx.rx_samples[57] ;
 wire \uart_0.rx.rx_samples[58] ;
 wire \uart_0.rx.rx_samples[59] ;
 wire \uart_0.rx.rx_samples[5] ;
 wire \uart_0.rx.rx_samples[60] ;
 wire \uart_0.rx.rx_samples[61] ;
 wire \uart_0.rx.rx_samples[62] ;
 wire \uart_0.rx.rx_samples[63] ;
 wire \uart_0.rx.rx_samples[64] ;
 wire \uart_0.rx.rx_samples[65] ;
 wire \uart_0.rx.rx_samples[66] ;
 wire \uart_0.rx.rx_samples[67] ;
 wire \uart_0.rx.rx_samples[68] ;
 wire \uart_0.rx.rx_samples[69] ;
 wire \uart_0.rx.rx_samples[6] ;
 wire \uart_0.rx.rx_samples[70] ;
 wire \uart_0.rx.rx_samples[71] ;
 wire \uart_0.rx.rx_samples[72] ;
 wire \uart_0.rx.rx_samples[73] ;
 wire \uart_0.rx.rx_samples[74] ;
 wire \uart_0.rx.rx_samples[75] ;
 wire \uart_0.rx.rx_samples[76] ;
 wire \uart_0.rx.rx_samples[77] ;
 wire \uart_0.rx.rx_samples[78] ;
 wire \uart_0.rx.rx_samples[79] ;
 wire \uart_0.rx.rx_samples[7] ;
 wire \uart_0.rx.rx_samples[80] ;
 wire \uart_0.rx.rx_samples[81] ;
 wire \uart_0.rx.rx_samples[82] ;
 wire \uart_0.rx.rx_samples[83] ;
 wire \uart_0.rx.rx_samples[84] ;
 wire \uart_0.rx.rx_samples[85] ;
 wire \uart_0.rx.rx_samples[86] ;
 wire \uart_0.rx.rx_samples[87] ;
 wire \uart_0.rx.rx_samples[88] ;
 wire \uart_0.rx.rx_samples[89] ;
 wire \uart_0.rx.rx_samples[8] ;
 wire \uart_0.rx.rx_samples[9] ;
 wire \uart_0.rx.rx_stop_zeros[0] ;
 wire \uart_0.rx.rx_stop_zeros[1] ;
 wire \uart_0.rx.rx_stop_zeros[2] ;
 wire \uart_0.rx.rx_stop_zeros[3] ;
 wire \uart_0.rx.rx_stop_zeros[4] ;
 wire \uart_0.rx.rx_stop_zeros[5] ;
 wire \uart_0.rx.rx_stop_zeros[6] ;
 wire \uart_0.tx.tx_baudrate_cnt[0] ;
 wire \uart_0.tx.tx_baudrate_cnt[1] ;
 wire \uart_0.tx.tx_baudrate_cnt[2] ;
 wire \uart_0.tx.tx_baudrate_cnt[3] ;
 wire \uart_0.tx.tx_baudrate_cnt[4] ;
 wire \uart_0.tx.tx_baudrate_cnt[5] ;
 wire \uart_0.tx.tx_baudrate_cnt[6] ;
 wire \uart_0.tx.tx_baudrate_cnt[7] ;
 wire \uart_0.tx.tx_bit_cnt[0] ;
 wire \uart_0.tx.tx_bit_cnt[1] ;
 wire \uart_0.tx.tx_bit_cnt[2] ;
 wire \uart_0.tx.tx_bit_cnt[3] ;
 wire \uart_0.tx.tx_data_tmp[2] ;
 wire \uart_0.tx.tx_data_tmp[3] ;
 wire \uart_0.tx.tx_data_tmp[4] ;
 wire \uart_0.tx.tx_data_tmp[5] ;
 wire \uart_0.tx.tx_data_tmp[6] ;
 wire \uart_0.tx.tx_data_tmp[7] ;
 wire \uart_0.tx.tx_data_tmp[8] ;
 wire \uart_0.tx.tx_data_tmp[9] ;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire clknet_0_clk;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net1;
 wire net2;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;

 sg13g2_inv_1 _1579_ (.Y(_0137_),
    .A(net1));
 sg13g2_inv_1 _1580_ (.Y(_1124_),
    .A(_0125_));
 sg13g2_inv_1 _1581_ (.Y(_1125_),
    .A(_0106_));
 sg13g2_inv_1 _1582_ (.Y(_1126_),
    .A(_0071_));
 sg13g2_inv_1 _1583_ (.Y(_1127_),
    .A(_0063_));
 sg13g2_inv_1 _1584_ (.Y(_1128_),
    .A(\uart_0.rx.rx_samples[86] ));
 sg13g2_inv_1 _1585_ (.Y(_1129_),
    .A(\uart_0.rx.rx_samples[87] ));
 sg13g2_inv_1 _1586_ (.Y(_1130_),
    .A(\uart_0.rx.rx_samples[88] ));
 sg13g2_inv_1 _1587_ (.Y(_1131_),
    .A(\uart_0.rx.rx_samples[8] ));
 sg13g2_inv_1 _1588_ (.Y(_1132_),
    .A(\uart_0.rx.rx_samples[7] ));
 sg13g2_inv_1 _1589_ (.Y(_1133_),
    .A(\uart_0.rx.rx_marker[0] ));
 sg13g2_inv_1 _1590_ (.Y(_1134_),
    .A(\uart_0.rx.rx_marker[6] ));
 sg13g2_inv_1 _1591_ (.Y(_1135_),
    .A(\uart_0.rx.rx_marker[5] ));
 sg13g2_inv_1 _1592_ (.Y(_1136_),
    .A(\fifo_t[2] ));
 sg13g2_inv_1 _1593_ (.Y(_1137_),
    .A(\uart_0.tx.tx_bit_cnt[1] ));
 sg13g2_inv_1 _1594_ (.Y(_1138_),
    .A(\uart_0.tx.tx_bit_cnt[2] ));
 sg13g2_inv_1 _1595_ (.Y(_1139_),
    .A(\uart_0.tx.tx_baudrate_cnt[3] ));
 sg13g2_inv_1 _1596_ (.Y(_1140_),
    .A(\uart_0.rx.rx_sample_clk_cnt[1] ));
 sg13g2_inv_1 _1597_ (.Y(_1141_),
    .A(\uart_0.rx.rx_sample_clk_cnt[4] ));
 sg13g2_inv_1 _1598_ (.Y(_1142_),
    .A(\uart_0.rx.rx_sample_cnt[2] ));
 sg13g2_inv_1 _1599_ (.Y(_1143_),
    .A(\uart_0.rx.rx_sample_cnt[0] ));
 sg13g2_inv_1 _1600_ (.Y(_1144_),
    .A(\fifo_d[0][0] ));
 sg13g2_inv_1 _1601_ (.Y(_1145_),
    .A(\fifo_d[0][1] ));
 sg13g2_inv_1 _1602_ (.Y(_1146_),
    .A(\fifo_d[0][2] ));
 sg13g2_inv_1 _1603_ (.Y(_1147_),
    .A(\fifo_d[0][3] ));
 sg13g2_inv_1 _1604_ (.Y(_1148_),
    .A(\fifo_d[0][4] ));
 sg13g2_inv_1 _1605_ (.Y(_1149_),
    .A(\fifo_d[0][5] ));
 sg13g2_inv_1 _1606_ (.Y(_1150_),
    .A(\fifo_d[0][6] ));
 sg13g2_inv_1 _1607_ (.Y(_1151_),
    .A(\fifo_d[0][7] ));
 sg13g2_inv_1 _1608_ (.Y(_1152_),
    .A(\uart_0.rx.rx_samples[77] ));
 sg13g2_inv_1 _1609_ (.Y(_1153_),
    .A(\uart_0.rx.rx_samples[68] ));
 sg13g2_inv_1 _1610_ (.Y(_1154_),
    .A(\uart_0.rx.rx_samples[62] ));
 sg13g2_inv_1 _1611_ (.Y(_1155_),
    .A(\uart_0.rx.rx_samples[58] ));
 sg13g2_inv_1 _1612_ (.Y(_1156_),
    .A(\uart_0.rx.rx_samples[53] ));
 sg13g2_inv_1 _1613_ (.Y(_1157_),
    .A(\uart_0.rx.rx_samples[51] ));
 sg13g2_inv_1 _1614_ (.Y(_1158_),
    .A(\uart_0.rx.rx_samples[44] ));
 sg13g2_inv_1 _1615_ (.Y(_1159_),
    .A(\uart_0.rx.rx_samples[40] ));
 sg13g2_inv_1 _1616_ (.Y(_1160_),
    .A(\uart_0.rx.rx_samples[35] ));
 sg13g2_inv_1 _1617_ (.Y(_1161_),
    .A(\uart_0.rx.rx_samples[31] ));
 sg13g2_inv_1 _1618_ (.Y(_1162_),
    .A(\uart_0.rx.rx_samples[23] ));
 sg13g2_inv_1 _1619_ (.Y(_1163_),
    .A(\uart_0.rx.rx_samples[15] ));
 sg13g2_inv_1 _1620_ (.Y(_1164_),
    .A(\uart_0.rx.rx_samples[13] ));
 sg13g2_inv_1 _1621_ (.Y(_1165_),
    .A(net851));
 sg13g2_inv_2 _1622_ (.Y(_1166_),
    .A(_0028_));
 sg13g2_inv_2 _1623_ (.Y(_1167_),
    .A(_0029_));
 sg13g2_inv_1 _1624_ (.Y(_1168_),
    .A(\uart_0.rx.rx_stop_zeros[6] ));
 sg13g2_inv_1 _1625_ (.Y(_1169_),
    .A(_0032_));
 sg13g2_and2_1 _1626_ (.A(\uart_0.rx.rx_samples[1] ),
    .B(\uart_0.rx.rx_samples[0] ),
    .X(_1170_));
 sg13g2_xor2_1 _1627_ (.B(\uart_0.rx.rx_samples[0] ),
    .A(\uart_0.rx.rx_samples[1] ),
    .X(_1171_));
 sg13g2_xnor2_1 _1628_ (.Y(_1172_),
    .A(\uart_0.rx.rx_samples[3] ),
    .B(_1171_));
 sg13g2_nor2_1 _1629_ (.A(_1131_),
    .B(_1172_),
    .Y(_1173_));
 sg13g2_nand2_1 _1630_ (.Y(_1174_),
    .A(_1131_),
    .B(_1172_));
 sg13g2_xnor2_1 _1631_ (.Y(_1175_),
    .A(_1131_),
    .B(_1172_));
 sg13g2_xnor2_1 _1632_ (.Y(_1176_),
    .A(\uart_0.rx.rx_samples[5] ),
    .B(_1175_));
 sg13g2_nand2_1 _1633_ (.Y(_1177_),
    .A(\uart_0.rx.rx_samples[6] ),
    .B(_1176_));
 sg13g2_xnor2_1 _1634_ (.Y(_1178_),
    .A(\uart_0.rx.rx_samples[6] ),
    .B(_1176_));
 sg13g2_xnor2_1 _1635_ (.Y(_1179_),
    .A(\uart_0.rx.rx_samples[7] ),
    .B(_1178_));
 sg13g2_nand3_1 _1636_ (.B(\uart_0.rx.rx_samples[2] ),
    .C(_1179_),
    .A(\uart_0.rx.rx_samples[4] ),
    .Y(_1180_));
 sg13g2_o21ai_1 _1637_ (.B1(_1177_),
    .Y(_1181_),
    .A1(_1132_),
    .A2(_1178_));
 sg13g2_or2_1 _1638_ (.X(_1182_),
    .B(\uart_0.rx.rx_samples[2] ),
    .A(\uart_0.rx.rx_samples[4] ));
 sg13g2_o21ai_1 _1639_ (.B1(_1181_),
    .Y(_1183_),
    .A1(_1179_),
    .A2(_1182_));
 sg13g2_a21oi_1 _1640_ (.A1(\uart_0.rx.rx_samples[5] ),
    .A2(_1174_),
    .Y(_1184_),
    .B1(_1173_));
 sg13g2_a21oi_1 _1641_ (.A1(\uart_0.rx.rx_samples[3] ),
    .A2(_1171_),
    .Y(_1185_),
    .B1(_1170_));
 sg13g2_xnor2_1 _1642_ (.Y(_1186_),
    .A(_1184_),
    .B(_1185_));
 sg13g2_a21oi_1 _1643_ (.A1(_1180_),
    .A2(_1183_),
    .Y(_1187_),
    .B1(_1186_));
 sg13g2_nor3_1 _1644_ (.A(_1179_),
    .B(_1181_),
    .C(_1182_),
    .Y(_1188_));
 sg13g2_or3_1 _1645_ (.A(_1184_),
    .B(_1185_),
    .C(_1188_),
    .X(_1189_));
 sg13g2_nand2b_1 _1646_ (.Y(_1190_),
    .B(_1181_),
    .A_N(_1180_));
 sg13g2_nand3b_1 _1647_ (.B(_1189_),
    .C(_1190_),
    .Y(_1191_),
    .A_N(_1187_));
 sg13g2_and2_1 _1648_ (.A(\uart_0.rx.rx_samples[81] ),
    .B(\uart_0.rx.rx_samples[82] ),
    .X(_1192_));
 sg13g2_xor2_1 _1649_ (.B(\uart_0.rx.rx_samples[82] ),
    .A(\uart_0.rx.rx_samples[81] ),
    .X(_1193_));
 sg13g2_xnor2_1 _1650_ (.Y(_1194_),
    .A(\uart_0.rx.rx_samples[84] ),
    .B(_1193_));
 sg13g2_inv_1 _1651_ (.Y(_1195_),
    .A(_1194_));
 sg13g2_nand2_1 _1652_ (.Y(_1196_),
    .A(\uart_0.rx.rx_samples[89] ),
    .B(_1195_));
 sg13g2_xor2_1 _1653_ (.B(_1194_),
    .A(\uart_0.rx.rx_samples[89] ),
    .X(_1197_));
 sg13g2_or2_1 _1654_ (.X(_1198_),
    .B(_1197_),
    .A(_1128_));
 sg13g2_xnor2_1 _1655_ (.Y(_1199_),
    .A(_1128_),
    .B(_1197_));
 sg13g2_or2_1 _1656_ (.X(_1200_),
    .B(_1199_),
    .A(_1129_));
 sg13g2_xnor2_1 _1657_ (.Y(_1201_),
    .A(_1129_),
    .B(_1199_));
 sg13g2_o21ai_1 _1658_ (.B1(_1200_),
    .Y(_1202_),
    .A1(_1130_),
    .A2(_1201_));
 sg13g2_xnor2_1 _1659_ (.Y(_1203_),
    .A(_1130_),
    .B(_1201_));
 sg13g2_nand2_1 _1660_ (.Y(_1204_),
    .A(\uart_0.rx.rx_samples[85] ),
    .B(\uart_0.rx.rx_samples[83] ));
 sg13g2_nor2_1 _1661_ (.A(_1203_),
    .B(_1204_),
    .Y(_1205_));
 sg13g2_a21oi_1 _1662_ (.A1(\uart_0.rx.rx_samples[84] ),
    .A2(_1193_),
    .Y(_1206_),
    .B1(_1192_));
 sg13g2_a21oi_1 _1663_ (.A1(_1196_),
    .A2(_1198_),
    .Y(_1207_),
    .B1(_1206_));
 sg13g2_o21ai_1 _1664_ (.B1(_1202_),
    .Y(_1208_),
    .A1(_1205_),
    .A2(_1207_));
 sg13g2_nor2_1 _1665_ (.A(\uart_0.rx.rx_samples[85] ),
    .B(\uart_0.rx.rx_samples[83] ),
    .Y(_1209_));
 sg13g2_nand2_1 _1666_ (.Y(_1210_),
    .A(_1203_),
    .B(_1209_));
 sg13g2_nand3_1 _1667_ (.B(_1198_),
    .C(_1206_),
    .A(_1196_),
    .Y(_1211_));
 sg13g2_nand2b_1 _1668_ (.Y(_1212_),
    .B(_1211_),
    .A_N(_1207_));
 sg13g2_a21oi_1 _1669_ (.A1(_1203_),
    .A2(_1209_),
    .Y(_1213_),
    .B1(_1212_));
 sg13g2_o21ai_1 _1670_ (.B1(_1213_),
    .Y(_1214_),
    .A1(_1202_),
    .A2(_1205_));
 sg13g2_nand2b_2 _1671_ (.Y(_1215_),
    .B(\uart_0.rx.rx_marker[4] ),
    .A_N(\uart_0.rx.rx_marker[5] ));
 sg13g2_or2_1 _1672_ (.X(_1216_),
    .B(_1215_),
    .A(net848));
 sg13g2_nand2_1 _1673_ (.Y(_1217_),
    .A(\uart_0.rx.rx_marker[3] ),
    .B(\uart_0.rx.rx_marker[6] ));
 sg13g2_nor3_1 _1674_ (.A(net848),
    .B(_1215_),
    .C(_1217_),
    .Y(_1218_));
 sg13g2_nor4_1 _1675_ (.A(_1133_),
    .B(\uart_0.rx.rx_marker[1] ),
    .C(_1216_),
    .D(_1217_),
    .Y(_1219_));
 sg13g2_inv_1 _1676_ (.Y(_1220_),
    .A(_1219_));
 sg13g2_a21oi_1 _1677_ (.A1(_1207_),
    .A2(_1210_),
    .Y(_1221_),
    .B1(_1220_));
 sg13g2_and4_1 _1678_ (.A(net720),
    .B(_1208_),
    .C(_1214_),
    .D(_1221_),
    .X(rx_data_ready));
 sg13g2_or2_1 _1679_ (.X(_1222_),
    .B(\uart_0.tx.tx_bit_cnt[0] ),
    .A(\uart_0.tx.tx_bit_cnt[1] ));
 sg13g2_or3_2 _1680_ (.A(\uart_0.tx.tx_bit_cnt[2] ),
    .B(\uart_0.tx.tx_bit_cnt[3] ),
    .C(_1222_),
    .X(_1223_));
 sg13g2_inv_4 _1681_ (.A(_1223_),
    .Y(tx_data_done));
 sg13g2_xor2_1 _1682_ (.B(\fifo_h[3] ),
    .A(net820),
    .X(_1224_));
 sg13g2_xor2_1 _1683_ (.B(net856),
    .A(\fifo_t[0] ),
    .X(_1225_));
 sg13g2_xnor2_1 _1684_ (.Y(_1226_),
    .A(\fifo_t[1] ),
    .B(net855));
 sg13g2_xnor2_1 _1685_ (.Y(_1227_),
    .A(\fifo_t[2] ),
    .B(\fifo_h[2] ));
 sg13g2_nand3b_1 _1686_ (.B(_1226_),
    .C(_1227_),
    .Y(_1228_),
    .A_N(_1225_));
 sg13g2_o21ai_1 _1687_ (.B1(tx_data_done),
    .Y(_1229_),
    .A1(_1224_),
    .A2(_1228_));
 sg13g2_inv_1 _1688_ (.Y(_0012_),
    .A(_1229_));
 sg13g2_mux2_1 _1689_ (.A0(\uart_0.tx.tx_data_tmp[8] ),
    .A1(\uart_0.tx.tx_data_tmp[9] ),
    .S(\uart_0.tx.tx_bit_cnt[0] ),
    .X(_1230_));
 sg13g2_nor2_1 _1690_ (.A(\uart_0.tx.tx_bit_cnt[1] ),
    .B(_1230_),
    .Y(_1231_));
 sg13g2_nor2b_1 _1691_ (.A(\uart_0.tx.tx_bit_cnt[2] ),
    .B_N(\uart_0.tx.tx_bit_cnt[3] ),
    .Y(_1232_));
 sg13g2_o21ai_1 _1692_ (.B1(_1232_),
    .Y(_1233_),
    .A1(_1137_),
    .A2(_0037_));
 sg13g2_nor2_1 _1693_ (.A(_1137_),
    .B(\uart_0.tx.tx_bit_cnt[0] ),
    .Y(_1234_));
 sg13g2_nand2_2 _1694_ (.Y(_1235_),
    .A(\uart_0.tx.tx_bit_cnt[1] ),
    .B(\uart_0.tx.tx_bit_cnt[0] ));
 sg13g2_mux4_1 _1695_ (.S0(\uart_0.tx.tx_bit_cnt[0] ),
    .A0(\uart_0.tx.tx_data_tmp[4] ),
    .A1(\uart_0.tx.tx_data_tmp[5] ),
    .A2(\uart_0.tx.tx_data_tmp[6] ),
    .A3(\uart_0.tx.tx_data_tmp[7] ),
    .S1(\uart_0.tx.tx_bit_cnt[1] ),
    .X(_1236_));
 sg13g2_nand3_1 _1696_ (.B(\uart_0.tx.tx_bit_cnt[0] ),
    .C(\uart_0.tx.tx_data_tmp[3] ),
    .A(\uart_0.tx.tx_bit_cnt[1] ),
    .Y(_1237_));
 sg13g2_a221oi_1 _1697_ (.B2(\uart_0.tx.tx_data_tmp[2] ),
    .C1(\uart_0.tx.tx_bit_cnt[2] ),
    .B1(_1234_),
    .A1(_1137_),
    .Y(_1238_),
    .A2(_0037_));
 sg13g2_a21oi_1 _1698_ (.A1(_1237_),
    .A2(_1238_),
    .Y(_1239_),
    .B1(\uart_0.tx.tx_bit_cnt[3] ));
 sg13g2_o21ai_1 _1699_ (.B1(_1239_),
    .Y(_1240_),
    .A1(_1138_),
    .A2(_1236_));
 sg13g2_o21ai_1 _1700_ (.B1(_1240_),
    .Y(tx_data_out),
    .A1(_1231_),
    .A2(_1233_));
 sg13g2_nand2_2 _1701_ (.Y(_1241_),
    .A(net856),
    .B(net855));
 sg13g2_nor3_2 _1702_ (.A(net854),
    .B(net853),
    .C(_1241_),
    .Y(_1242_));
 sg13g2_nand2_2 _1703_ (.Y(_1243_),
    .A(net854),
    .B(net853));
 sg13g2_nor3_2 _1704_ (.A(net856),
    .B(net855),
    .C(_1243_),
    .Y(_1244_));
 sg13g2_nor2_2 _1705_ (.A(_1241_),
    .B(_1243_),
    .Y(_1245_));
 sg13g2_nand2b_2 _1706_ (.Y(_1246_),
    .B(net855),
    .A_N(net856));
 sg13g2_nor2_2 _1707_ (.A(_1243_),
    .B(_1246_),
    .Y(_1247_));
 sg13g2_nor4_2 _1708_ (.A(\fifo_h[0] ),
    .B(\fifo_h[1] ),
    .C(\fifo_h[2] ),
    .Y(_1248_),
    .D(net853));
 sg13g2_nand2b_2 _1709_ (.Y(_1249_),
    .B(net853),
    .A_N(net854));
 sg13g2_nand2b_2 _1710_ (.Y(_1250_),
    .B(net856),
    .A_N(net855));
 sg13g2_nor2_2 _1711_ (.A(_1249_),
    .B(_1250_),
    .Y(_1251_));
 sg13g2_nand2b_2 _1712_ (.Y(_1252_),
    .B(net854),
    .A_N(net853));
 sg13g2_inv_1 _1713_ (.Y(_1253_),
    .A(_1252_));
 sg13g2_nor2_2 _1714_ (.A(_1250_),
    .B(_1252_),
    .Y(_1254_));
 sg13g2_nor2_2 _1715_ (.A(_1243_),
    .B(_1250_),
    .Y(_1255_));
 sg13g2_nor3_2 _1716_ (.A(net856),
    .B(net855),
    .C(_1249_),
    .Y(_1256_));
 sg13g2_nor3_2 _1717_ (.A(net854),
    .B(net853),
    .C(_1250_),
    .Y(_1257_));
 sg13g2_nor2_2 _1718_ (.A(_1246_),
    .B(_1252_),
    .Y(_1258_));
 sg13g2_nor3_2 _1719_ (.A(net856),
    .B(net855),
    .C(_1252_),
    .Y(_1259_));
 sg13g2_nor2_2 _1720_ (.A(_1246_),
    .B(_1249_),
    .Y(_1260_));
 sg13g2_nor3_2 _1721_ (.A(net854),
    .B(net853),
    .C(_1246_),
    .Y(_1261_));
 sg13g2_nor2_2 _1722_ (.A(_1241_),
    .B(_1252_),
    .Y(_1262_));
 sg13g2_nor2_2 _1723_ (.A(_1241_),
    .B(_1249_),
    .Y(_1263_));
 sg13g2_a21oi_1 _1724_ (.A1(\fifo_d[7][0] ),
    .A2(_1262_),
    .Y(_1264_),
    .B1(_1248_));
 sg13g2_a22oi_1 _1725_ (.Y(_1265_),
    .B1(_1258_),
    .B2(\fifo_d[6][0] ),
    .A2(_1242_),
    .A1(\fifo_d[3][0] ));
 sg13g2_a22oi_1 _1726_ (.Y(_1266_),
    .B1(_1260_),
    .B2(\fifo_d[10][0] ),
    .A2(_1245_),
    .A1(\fifo_d[15][0] ));
 sg13g2_a22oi_1 _1727_ (.Y(_1267_),
    .B1(_1263_),
    .B2(\fifo_d[11][0] ),
    .A2(_1256_),
    .A1(\fifo_d[8][0] ));
 sg13g2_nand4_1 _1728_ (.B(_1265_),
    .C(_1266_),
    .A(_1264_),
    .Y(_1268_),
    .D(_1267_));
 sg13g2_a22oi_1 _1729_ (.Y(_1269_),
    .B1(_1261_),
    .B2(\fifo_d[2][0] ),
    .A2(_1257_),
    .A1(\fifo_d[1][0] ));
 sg13g2_a22oi_1 _1730_ (.Y(_1270_),
    .B1(_1259_),
    .B2(\fifo_d[4][0] ),
    .A2(_1247_),
    .A1(\fifo_d[14][0] ));
 sg13g2_a22oi_1 _1731_ (.Y(_1271_),
    .B1(_1254_),
    .B2(\fifo_d[5][0] ),
    .A2(_1244_),
    .A1(\fifo_d[12][0] ));
 sg13g2_a22oi_1 _1732_ (.Y(_1272_),
    .B1(_1255_),
    .B2(\fifo_d[13][0] ),
    .A2(_1251_),
    .A1(\fifo_d[9][0] ));
 sg13g2_nand4_1 _1733_ (.B(_1270_),
    .C(_1271_),
    .A(_1269_),
    .Y(_1273_),
    .D(_1272_));
 sg13g2_o21ai_1 _1734_ (.B1(_0012_),
    .Y(_1274_),
    .A1(_1268_),
    .A2(_1273_));
 sg13g2_a21oi_1 _1735_ (.A1(_1144_),
    .A2(net822),
    .Y(_0004_),
    .B1(_1274_));
 sg13g2_a22oi_1 _1736_ (.Y(_1275_),
    .B1(_1262_),
    .B2(\fifo_d[7][1] ),
    .A2(_1251_),
    .A1(\fifo_d[9][1] ));
 sg13g2_a22oi_1 _1737_ (.Y(_1276_),
    .B1(_1257_),
    .B2(\fifo_d[1][1] ),
    .A2(_1256_),
    .A1(\fifo_d[8][1] ));
 sg13g2_a21oi_1 _1738_ (.A1(\fifo_d[11][1] ),
    .A2(_1263_),
    .Y(_1277_),
    .B1(net822));
 sg13g2_a22oi_1 _1739_ (.Y(_1278_),
    .B1(_1260_),
    .B2(\fifo_d[10][1] ),
    .A2(_1254_),
    .A1(\fifo_d[5][1] ));
 sg13g2_a22oi_1 _1740_ (.Y(_1279_),
    .B1(_1261_),
    .B2(\fifo_d[2][1] ),
    .A2(_1258_),
    .A1(\fifo_d[6][1] ));
 sg13g2_nand4_1 _1741_ (.B(_1277_),
    .C(_1278_),
    .A(_1275_),
    .Y(_1280_),
    .D(_1279_));
 sg13g2_a22oi_1 _1742_ (.Y(_1281_),
    .B1(_1255_),
    .B2(\fifo_d[13][1] ),
    .A2(_1245_),
    .A1(\fifo_d[15][1] ));
 sg13g2_a22oi_1 _1743_ (.Y(_1282_),
    .B1(_1247_),
    .B2(\fifo_d[14][1] ),
    .A2(_1242_),
    .A1(\fifo_d[3][1] ));
 sg13g2_a22oi_1 _1744_ (.Y(_1283_),
    .B1(_1259_),
    .B2(\fifo_d[4][1] ),
    .A2(_1244_),
    .A1(\fifo_d[12][1] ));
 sg13g2_nand4_1 _1745_ (.B(_1281_),
    .C(_1282_),
    .A(_1276_),
    .Y(_1284_),
    .D(_1283_));
 sg13g2_o21ai_1 _1746_ (.B1(net754),
    .Y(_1285_),
    .A1(_1280_),
    .A2(_1284_));
 sg13g2_a21oi_1 _1747_ (.A1(_1145_),
    .A2(net822),
    .Y(_0005_),
    .B1(_1285_));
 sg13g2_a22oi_1 _1748_ (.Y(_1286_),
    .B1(_1261_),
    .B2(\fifo_d[2][2] ),
    .A2(_1254_),
    .A1(\fifo_d[5][2] ));
 sg13g2_a22oi_1 _1749_ (.Y(_1287_),
    .B1(_1255_),
    .B2(\fifo_d[13][2] ),
    .A2(_1244_),
    .A1(\fifo_d[12][2] ));
 sg13g2_a22oi_1 _1750_ (.Y(_1288_),
    .B1(_1256_),
    .B2(\fifo_d[8][2] ),
    .A2(_1251_),
    .A1(\fifo_d[9][2] ));
 sg13g2_a22oi_1 _1751_ (.Y(_1289_),
    .B1(_1259_),
    .B2(\fifo_d[4][2] ),
    .A2(_1257_),
    .A1(\fifo_d[1][2] ));
 sg13g2_a22oi_1 _1752_ (.Y(_1290_),
    .B1(_1263_),
    .B2(\fifo_d[11][2] ),
    .A2(_1262_),
    .A1(\fifo_d[7][2] ));
 sg13g2_a21oi_1 _1753_ (.A1(\fifo_d[15][2] ),
    .A2(_1245_),
    .Y(_1291_),
    .B1(net822));
 sg13g2_a22oi_1 _1754_ (.Y(_1292_),
    .B1(_1260_),
    .B2(\fifo_d[10][2] ),
    .A2(_1258_),
    .A1(\fifo_d[6][2] ));
 sg13g2_nand4_1 _1755_ (.B(_1290_),
    .C(_1291_),
    .A(_1286_),
    .Y(_1293_),
    .D(_1292_));
 sg13g2_a22oi_1 _1756_ (.Y(_1294_),
    .B1(_1247_),
    .B2(\fifo_d[14][2] ),
    .A2(_1242_),
    .A1(\fifo_d[3][2] ));
 sg13g2_nand4_1 _1757_ (.B(_1288_),
    .C(_1289_),
    .A(_1287_),
    .Y(_1295_),
    .D(_1294_));
 sg13g2_o21ai_1 _1758_ (.B1(net754),
    .Y(_1296_),
    .A1(_1293_),
    .A2(_1295_));
 sg13g2_a21oi_1 _1759_ (.A1(_1146_),
    .A2(net822),
    .Y(_0006_),
    .B1(_1296_));
 sg13g2_a21oi_1 _1760_ (.A1(\fifo_d[8][3] ),
    .A2(_1256_),
    .Y(_1297_),
    .B1(net823));
 sg13g2_a22oi_1 _1761_ (.Y(_1298_),
    .B1(_1260_),
    .B2(\fifo_d[10][3] ),
    .A2(_1251_),
    .A1(\fifo_d[9][3] ));
 sg13g2_a22oi_1 _1762_ (.Y(_1299_),
    .B1(_1263_),
    .B2(\fifo_d[11][3] ),
    .A2(_1259_),
    .A1(\fifo_d[4][3] ));
 sg13g2_a22oi_1 _1763_ (.Y(_1300_),
    .B1(_1254_),
    .B2(\fifo_d[5][3] ),
    .A2(_1244_),
    .A1(\fifo_d[12][3] ));
 sg13g2_nand4_1 _1764_ (.B(_1298_),
    .C(_1299_),
    .A(_1297_),
    .Y(_1301_),
    .D(_1300_));
 sg13g2_a22oi_1 _1765_ (.Y(_1302_),
    .B1(_1255_),
    .B2(\fifo_d[13][3] ),
    .A2(_1247_),
    .A1(\fifo_d[14][3] ));
 sg13g2_a22oi_1 _1766_ (.Y(_1303_),
    .B1(_1262_),
    .B2(\fifo_d[7][3] ),
    .A2(_1258_),
    .A1(\fifo_d[6][3] ));
 sg13g2_a22oi_1 _1767_ (.Y(_1304_),
    .B1(_1261_),
    .B2(\fifo_d[2][3] ),
    .A2(_1257_),
    .A1(\fifo_d[1][3] ));
 sg13g2_a22oi_1 _1768_ (.Y(_1305_),
    .B1(_1245_),
    .B2(\fifo_d[15][3] ),
    .A2(_1242_),
    .A1(\fifo_d[3][3] ));
 sg13g2_nand4_1 _1769_ (.B(_1303_),
    .C(_1304_),
    .A(_1302_),
    .Y(_1306_),
    .D(_1305_));
 sg13g2_o21ai_1 _1770_ (.B1(net754),
    .Y(_1307_),
    .A1(_1301_),
    .A2(_1306_));
 sg13g2_a21oi_1 _1771_ (.A1(_1147_),
    .A2(net823),
    .Y(_0007_),
    .B1(_1307_));
 sg13g2_a22oi_1 _1772_ (.Y(_1308_),
    .B1(_1254_),
    .B2(\fifo_d[5][4] ),
    .A2(_1247_),
    .A1(\fifo_d[14][4] ));
 sg13g2_a22oi_1 _1773_ (.Y(_1309_),
    .B1(_1257_),
    .B2(\fifo_d[1][4] ),
    .A2(_1251_),
    .A1(\fifo_d[9][4] ));
 sg13g2_a22oi_1 _1774_ (.Y(_1310_),
    .B1(_1260_),
    .B2(\fifo_d[10][4] ),
    .A2(_1245_),
    .A1(\fifo_d[15][4] ));
 sg13g2_a22oi_1 _1775_ (.Y(_1311_),
    .B1(_1261_),
    .B2(\fifo_d[2][4] ),
    .A2(_1244_),
    .A1(\fifo_d[12][4] ));
 sg13g2_a21oi_2 _1776_ (.B1(net823),
    .Y(_1312_),
    .A2(_1255_),
    .A1(\fifo_d[13][4] ));
 sg13g2_a22oi_1 _1777_ (.Y(_1313_),
    .B1(_1262_),
    .B2(\fifo_d[7][4] ),
    .A2(_1256_),
    .A1(\fifo_d[8][4] ));
 sg13g2_nand4_1 _1778_ (.B(_1310_),
    .C(_1312_),
    .A(_1309_),
    .Y(_1314_),
    .D(_1313_));
 sg13g2_a22oi_1 _1779_ (.Y(_1315_),
    .B1(_1263_),
    .B2(\fifo_d[11][4] ),
    .A2(_1258_),
    .A1(\fifo_d[6][4] ));
 sg13g2_a22oi_1 _1780_ (.Y(_1316_),
    .B1(_1259_),
    .B2(\fifo_d[4][4] ),
    .A2(_1242_),
    .A1(\fifo_d[3][4] ));
 sg13g2_nand4_1 _1781_ (.B(_1311_),
    .C(_1315_),
    .A(_1308_),
    .Y(_1317_),
    .D(_1316_));
 sg13g2_o21ai_1 _1782_ (.B1(net754),
    .Y(_1318_),
    .A1(_1314_),
    .A2(_1317_));
 sg13g2_a21oi_1 _1783_ (.A1(_1148_),
    .A2(net822),
    .Y(_0008_),
    .B1(_1318_));
 sg13g2_a22oi_1 _1784_ (.Y(_1319_),
    .B1(_1256_),
    .B2(\fifo_d[8][5] ),
    .A2(_1251_),
    .A1(\fifo_d[9][5] ));
 sg13g2_a22oi_1 _1785_ (.Y(_1320_),
    .B1(_1261_),
    .B2(\fifo_d[2][5] ),
    .A2(_1244_),
    .A1(\fifo_d[12][5] ));
 sg13g2_a22oi_1 _1786_ (.Y(_1321_),
    .B1(_1258_),
    .B2(\fifo_d[6][5] ),
    .A2(_1254_),
    .A1(\fifo_d[5][5] ));
 sg13g2_a22oi_1 _1787_ (.Y(_1322_),
    .B1(_1260_),
    .B2(\fifo_d[10][5] ),
    .A2(_1257_),
    .A1(\fifo_d[1][5] ));
 sg13g2_a21oi_1 _1788_ (.A1(\fifo_d[14][5] ),
    .A2(_1247_),
    .Y(_1323_),
    .B1(net823));
 sg13g2_a22oi_1 _1789_ (.Y(_1324_),
    .B1(_1262_),
    .B2(\fifo_d[7][5] ),
    .A2(_1245_),
    .A1(\fifo_d[15][5] ));
 sg13g2_nand4_1 _1790_ (.B(_1322_),
    .C(_1323_),
    .A(_1319_),
    .Y(_1325_),
    .D(_1324_));
 sg13g2_a22oi_1 _1791_ (.Y(_1326_),
    .B1(_1263_),
    .B2(\fifo_d[11][5] ),
    .A2(_1259_),
    .A1(\fifo_d[4][5] ));
 sg13g2_a22oi_1 _1792_ (.Y(_1327_),
    .B1(_1255_),
    .B2(\fifo_d[13][5] ),
    .A2(_1242_),
    .A1(\fifo_d[3][5] ));
 sg13g2_nand4_1 _1793_ (.B(_1321_),
    .C(_1326_),
    .A(_1320_),
    .Y(_1328_),
    .D(_1327_));
 sg13g2_o21ai_1 _1794_ (.B1(net754),
    .Y(_1329_),
    .A1(_1325_),
    .A2(_1328_));
 sg13g2_a21oi_1 _1795_ (.A1(_1149_),
    .A2(net823),
    .Y(_0009_),
    .B1(_1329_));
 sg13g2_a22oi_1 _1796_ (.Y(_1330_),
    .B1(_1260_),
    .B2(\fifo_d[10][6] ),
    .A2(_1256_),
    .A1(\fifo_d[8][6] ));
 sg13g2_a21oi_1 _1797_ (.A1(\fifo_d[9][6] ),
    .A2(_1251_),
    .Y(_1331_),
    .B1(net823));
 sg13g2_a22oi_1 _1798_ (.Y(_1332_),
    .B1(_1263_),
    .B2(\fifo_d[11][6] ),
    .A2(_1255_),
    .A1(\fifo_d[13][6] ));
 sg13g2_a22oi_1 _1799_ (.Y(_1333_),
    .B1(_1254_),
    .B2(\fifo_d[5][6] ),
    .A2(_1244_),
    .A1(\fifo_d[12][6] ));
 sg13g2_nand4_1 _1800_ (.B(_1331_),
    .C(_1332_),
    .A(_1330_),
    .Y(_1334_),
    .D(_1333_));
 sg13g2_a22oi_1 _1801_ (.Y(_1335_),
    .B1(_1259_),
    .B2(\fifo_d[4][6] ),
    .A2(_1247_),
    .A1(\fifo_d[14][6] ));
 sg13g2_a22oi_1 _1802_ (.Y(_1336_),
    .B1(_1262_),
    .B2(\fifo_d[7][6] ),
    .A2(_1258_),
    .A1(\fifo_d[6][6] ));
 sg13g2_a22oi_1 _1803_ (.Y(_1337_),
    .B1(_1261_),
    .B2(\fifo_d[2][6] ),
    .A2(_1245_),
    .A1(\fifo_d[15][6] ));
 sg13g2_a22oi_1 _1804_ (.Y(_1338_),
    .B1(_1257_),
    .B2(\fifo_d[1][6] ),
    .A2(_1242_),
    .A1(\fifo_d[3][6] ));
 sg13g2_nand4_1 _1805_ (.B(_1336_),
    .C(_1337_),
    .A(_1335_),
    .Y(_1339_),
    .D(_1338_));
 sg13g2_o21ai_1 _1806_ (.B1(net754),
    .Y(_1340_),
    .A1(_1334_),
    .A2(_1339_));
 sg13g2_a21oi_1 _1807_ (.A1(_1150_),
    .A2(net823),
    .Y(_0010_),
    .B1(_1340_));
 sg13g2_a22oi_1 _1808_ (.Y(_1341_),
    .B1(_1258_),
    .B2(\fifo_d[6][7] ),
    .A2(_1251_),
    .A1(\fifo_d[9][7] ));
 sg13g2_a22oi_1 _1809_ (.Y(_1342_),
    .B1(_1257_),
    .B2(\fifo_d[1][7] ),
    .A2(_1254_),
    .A1(\fifo_d[5][7] ));
 sg13g2_a21oi_1 _1810_ (.A1(\fifo_d[15][7] ),
    .A2(_1245_),
    .Y(_1343_),
    .B1(net822));
 sg13g2_a22oi_1 _1811_ (.Y(_1344_),
    .B1(_1263_),
    .B2(\fifo_d[11][7] ),
    .A2(_1261_),
    .A1(\fifo_d[2][7] ));
 sg13g2_a22oi_1 _1812_ (.Y(_1345_),
    .B1(_1256_),
    .B2(\fifo_d[8][7] ),
    .A2(_1242_),
    .A1(\fifo_d[3][7] ));
 sg13g2_nand4_1 _1813_ (.B(_1343_),
    .C(_1344_),
    .A(_1341_),
    .Y(_1346_),
    .D(_1345_));
 sg13g2_a22oi_1 _1814_ (.Y(_1347_),
    .B1(_1259_),
    .B2(\fifo_d[4][7] ),
    .A2(_1244_),
    .A1(\fifo_d[12][7] ));
 sg13g2_a22oi_1 _1815_ (.Y(_1348_),
    .B1(_1262_),
    .B2(\fifo_d[7][7] ),
    .A2(_1247_),
    .A1(\fifo_d[14][7] ));
 sg13g2_a22oi_1 _1816_ (.Y(_1349_),
    .B1(_1260_),
    .B2(\fifo_d[10][7] ),
    .A2(_1255_),
    .A1(\fifo_d[13][7] ));
 sg13g2_nand4_1 _1817_ (.B(_1347_),
    .C(_1348_),
    .A(_1342_),
    .Y(_1350_),
    .D(_1349_));
 sg13g2_o21ai_1 _1818_ (.B1(net754),
    .Y(_1351_),
    .A1(_1346_),
    .A2(_1350_));
 sg13g2_a21oi_1 _1819_ (.A1(_1151_),
    .A2(net822),
    .Y(_0011_),
    .B1(_1351_));
 sg13g2_nor4_2 _1820_ (.A(\clk_out_cnt[1] ),
    .B(net26),
    .C(net24),
    .Y(_1352_),
    .D(\clk_out_cnt[2] ));
 sg13g2_nor2_1 _1821_ (.A(net26),
    .B(_1352_),
    .Y(_0000_));
 sg13g2_xor2_1 _1822_ (.B(net26),
    .A(net28),
    .X(_0001_));
 sg13g2_nand3_1 _1823_ (.B(net26),
    .C(net29),
    .A(net28),
    .Y(_1353_));
 sg13g2_a21o_1 _1824_ (.A2(net26),
    .A1(net28),
    .B1(net29),
    .X(_1354_));
 sg13g2_and2_1 _1825_ (.A(_1353_),
    .B(_1354_),
    .X(_0002_));
 sg13g2_xnor2_1 _1826_ (.Y(_0003_),
    .A(net24),
    .B(_1353_));
 sg13g2_nor2b_1 _1827_ (.A(\uart_0.tx.tx_baudrate_cnt[5] ),
    .B_N(\uart_0.tx.tx_baudrate_cnt[4] ),
    .Y(_1355_));
 sg13g2_nor4_1 _1828_ (.A(\uart_0.tx.tx_baudrate_cnt[1] ),
    .B(\uart_0.tx.tx_baudrate_cnt[0] ),
    .C(\uart_0.tx.tx_baudrate_cnt[2] ),
    .D(_1139_),
    .Y(_1356_));
 sg13g2_nand4_1 _1829_ (.B(\uart_0.tx.tx_baudrate_cnt[7] ),
    .C(_1355_),
    .A(\uart_0.tx.tx_baudrate_cnt[6] ),
    .Y(_1357_),
    .D(_1356_));
 sg13g2_nand2_2 _1830_ (.Y(_1358_),
    .A(net818),
    .B(_1357_));
 sg13g2_inv_1 _1831_ (.Y(_1359_),
    .A(_1358_));
 sg13g2_nor2_1 _1832_ (.A(\uart_0.tx.tx_baudrate_cnt[0] ),
    .B(_1358_),
    .Y(_0020_));
 sg13g2_xnor2_1 _1833_ (.Y(_1360_),
    .A(\uart_0.tx.tx_baudrate_cnt[1] ),
    .B(\uart_0.tx.tx_baudrate_cnt[0] ));
 sg13g2_nor2_1 _1834_ (.A(tx_data_done),
    .B(_1360_),
    .Y(_0021_));
 sg13g2_a21oi_1 _1835_ (.A1(\uart_0.tx.tx_baudrate_cnt[1] ),
    .A2(\uart_0.tx.tx_baudrate_cnt[0] ),
    .Y(_1361_),
    .B1(\uart_0.tx.tx_baudrate_cnt[2] ));
 sg13g2_and3_1 _1836_ (.X(_1362_),
    .A(\uart_0.tx.tx_baudrate_cnt[1] ),
    .B(\uart_0.tx.tx_baudrate_cnt[0] ),
    .C(\uart_0.tx.tx_baudrate_cnt[2] ));
 sg13g2_nor3_1 _1837_ (.A(tx_data_done),
    .B(_1361_),
    .C(_1362_),
    .Y(_0022_));
 sg13g2_and2_1 _1838_ (.A(\uart_0.tx.tx_baudrate_cnt[3] ),
    .B(_1362_),
    .X(_1363_));
 sg13g2_nor2_1 _1839_ (.A(\uart_0.tx.tx_baudrate_cnt[3] ),
    .B(_1362_),
    .Y(_1364_));
 sg13g2_nor3_1 _1840_ (.A(_1358_),
    .B(_1363_),
    .C(_1364_),
    .Y(_0023_));
 sg13g2_a21oi_1 _1841_ (.A1(\uart_0.tx.tx_baudrate_cnt[4] ),
    .A2(_1363_),
    .Y(_1365_),
    .B1(_1358_));
 sg13g2_o21ai_1 _1842_ (.B1(_1365_),
    .Y(_1366_),
    .A1(\uart_0.tx.tx_baudrate_cnt[4] ),
    .A2(_1363_));
 sg13g2_inv_1 _1843_ (.Y(_0024_),
    .A(_1366_));
 sg13g2_a21oi_1 _1844_ (.A1(\uart_0.tx.tx_baudrate_cnt[4] ),
    .A2(_1363_),
    .Y(_1367_),
    .B1(\uart_0.tx.tx_baudrate_cnt[5] ));
 sg13g2_and3_1 _1845_ (.X(_1368_),
    .A(\uart_0.tx.tx_baudrate_cnt[5] ),
    .B(\uart_0.tx.tx_baudrate_cnt[4] ),
    .C(_1363_));
 sg13g2_nor3_1 _1846_ (.A(tx_data_done),
    .B(_1367_),
    .C(_1368_),
    .Y(_0025_));
 sg13g2_nand2_1 _1847_ (.Y(_1369_),
    .A(\uart_0.tx.tx_baudrate_cnt[6] ),
    .B(_1368_));
 sg13g2_o21ai_1 _1848_ (.B1(_1359_),
    .Y(_1370_),
    .A1(\uart_0.tx.tx_baudrate_cnt[6] ),
    .A2(_1368_));
 sg13g2_nor2b_1 _1849_ (.A(_1370_),
    .B_N(_1369_),
    .Y(_0026_));
 sg13g2_xor2_1 _1850_ (.B(_1369_),
    .A(\uart_0.tx.tx_baudrate_cnt[7] ),
    .X(_1371_));
 sg13g2_nor2_1 _1851_ (.A(_1358_),
    .B(_1371_),
    .Y(_0027_));
 sg13g2_a21oi_1 _1852_ (.A1(\uart_0.rx.rx_marker[3] ),
    .A2(\uart_0.rx.rx_marker[4] ),
    .Y(_1372_),
    .B1(\uart_0.rx.rx_marker[5] ));
 sg13g2_nor2_1 _1853_ (.A(_1134_),
    .B(_1372_),
    .Y(_1373_));
 sg13g2_and2_2 _1854_ (.A(\uart_0.rx.rx_marker[0] ),
    .B(\uart_0.rx.rx_marker[1] ),
    .X(_1374_));
 sg13g2_nand2_1 _1855_ (.Y(_1375_),
    .A(\uart_0.rx.rx_marker[0] ),
    .B(\uart_0.rx.rx_marker[1] ));
 sg13g2_or3_1 _1856_ (.A(net848),
    .B(_1215_),
    .C(_1374_),
    .X(_1376_));
 sg13g2_and2_1 _1857_ (.A(_1373_),
    .B(_1376_),
    .X(_1377_));
 sg13g2_nor2b_1 _1858_ (.A(\uart_0.rx.rx_marker[0] ),
    .B_N(\uart_0.rx.rx_marker[1] ),
    .Y(_1378_));
 sg13g2_a22oi_1 _1859_ (.Y(_1379_),
    .B1(_1378_),
    .B2(_1218_),
    .A2(_1376_),
    .A1(_1373_));
 sg13g2_a21o_1 _1860_ (.A2(_1378_),
    .A1(_1218_),
    .B1(_1377_),
    .X(_1380_));
 sg13g2_nor2_1 _1861_ (.A(\uart_0.rx.rx_sample_clk_cnt[0] ),
    .B(\uart_0.rx.rx_sample_clk_cnt[1] ),
    .Y(_1381_));
 sg13g2_and2_1 _1862_ (.A(\uart_0.rx.rx_sample_clk_cnt[0] ),
    .B(\uart_0.rx.rx_sample_clk_cnt[1] ),
    .X(_1382_));
 sg13g2_and3_1 _1863_ (.X(_1383_),
    .A(\uart_0.rx.rx_sample_clk_cnt[0] ),
    .B(\uart_0.rx.rx_sample_clk_cnt[1] ),
    .C(\uart_0.rx.rx_sample_clk_cnt[2] ));
 sg13g2_a21o_1 _1864_ (.A2(_1383_),
    .A1(\uart_0.rx.rx_sample_wrap[0] ),
    .B1(_1381_),
    .X(_1384_));
 sg13g2_o21ai_1 _1865_ (.B1(_1140_),
    .Y(_1385_),
    .A1(\uart_0.rx.rx_sample_wrap[0] ),
    .A2(\uart_0.rx.rx_sample_clk_cnt[2] ));
 sg13g2_xor2_1 _1866_ (.B(\uart_0.rx.rx_sample_clk_cnt[3] ),
    .A(\uart_0.rx.rx_sample_wrap[3] ),
    .X(_1386_));
 sg13g2_nor4_1 _1867_ (.A(\uart_0.rx.rx_sample_clk_cnt[5] ),
    .B(_1141_),
    .C(\uart_0.rx.rx_sample_clk_cnt[6] ),
    .D(_1386_),
    .Y(_1387_));
 sg13g2_nand3_1 _1868_ (.B(_1385_),
    .C(_1387_),
    .A(_1384_),
    .Y(_1388_));
 sg13g2_and2_1 _1869_ (.A(net816),
    .B(_1388_),
    .X(_1389_));
 sg13g2_nand2_2 _1870_ (.Y(_1390_),
    .A(net816),
    .B(_1388_));
 sg13g2_nor2_1 _1871_ (.A(\uart_0.rx.rx_sample_clk_cnt[0] ),
    .B(_1390_),
    .Y(_0013_));
 sg13g2_nor3_1 _1872_ (.A(net784),
    .B(_1381_),
    .C(_1382_),
    .Y(_0014_));
 sg13g2_o21ai_1 _1873_ (.B1(net816),
    .Y(_1391_),
    .A1(\uart_0.rx.rx_sample_clk_cnt[2] ),
    .A2(_1382_));
 sg13g2_nor2_1 _1874_ (.A(_1383_),
    .B(_1391_),
    .Y(_0015_));
 sg13g2_and2_1 _1875_ (.A(\uart_0.rx.rx_sample_clk_cnt[3] ),
    .B(_1383_),
    .X(_1392_));
 sg13g2_nor2_1 _1876_ (.A(\uart_0.rx.rx_sample_clk_cnt[3] ),
    .B(_1383_),
    .Y(_1393_));
 sg13g2_nor3_1 _1877_ (.A(_1390_),
    .B(_1392_),
    .C(_1393_),
    .Y(_0016_));
 sg13g2_and2_1 _1878_ (.A(\uart_0.rx.rx_sample_clk_cnt[4] ),
    .B(_1392_),
    .X(_1394_));
 sg13g2_nor2_1 _1879_ (.A(\uart_0.rx.rx_sample_clk_cnt[4] ),
    .B(_1392_),
    .Y(_1395_));
 sg13g2_nor3_1 _1880_ (.A(_1390_),
    .B(_1394_),
    .C(_1395_),
    .Y(_0017_));
 sg13g2_and2_1 _1881_ (.A(\uart_0.rx.rx_sample_clk_cnt[5] ),
    .B(_1394_),
    .X(_0401_));
 sg13g2_nor2_1 _1882_ (.A(\uart_0.rx.rx_sample_clk_cnt[5] ),
    .B(_1394_),
    .Y(_0402_));
 sg13g2_nor3_1 _1883_ (.A(_1390_),
    .B(_0401_),
    .C(_0402_),
    .Y(_0018_));
 sg13g2_a21oi_1 _1884_ (.A1(\uart_0.rx.rx_sample_clk_cnt[6] ),
    .A2(_0401_),
    .Y(_0403_),
    .B1(net784));
 sg13g2_o21ai_1 _1885_ (.B1(_0403_),
    .Y(_0404_),
    .A1(\uart_0.rx.rx_sample_clk_cnt[6] ),
    .A2(_0401_));
 sg13g2_inv_1 _1886_ (.Y(_0019_),
    .A(_0404_));
 sg13g2_mux2_1 _1887_ (.A0(net881),
    .A1(net22),
    .S(_1352_),
    .X(_0138_));
 sg13g2_mux2_1 _1888_ (.A0(_0040_),
    .A1(net856),
    .S(_1229_),
    .X(_0139_));
 sg13g2_a21oi_1 _1889_ (.A1(_1246_),
    .A2(_1250_),
    .Y(_0405_),
    .B1(_1229_));
 sg13g2_a21o_1 _1890_ (.A2(_1229_),
    .A1(net855),
    .B1(_0405_),
    .X(_0140_));
 sg13g2_nor2_1 _1891_ (.A(_1229_),
    .B(_1241_),
    .Y(_0406_));
 sg13g2_nand2_1 _1892_ (.Y(_0407_),
    .A(net854),
    .B(_0406_));
 sg13g2_xor2_1 _1893_ (.B(_0406_),
    .A(net854),
    .X(_0141_));
 sg13g2_a22oi_1 _1894_ (.Y(_0408_),
    .B1(_0407_),
    .B2(net853),
    .A2(_0406_),
    .A1(_1253_));
 sg13g2_inv_1 _1895_ (.Y(_0142_),
    .A(_0408_));
 sg13g2_and2_2 _1896_ (.A(\fifo_t[0] ),
    .B(\fifo_t[1] ),
    .X(_0409_));
 sg13g2_nor2_2 _1897_ (.A(\fifo_t[0] ),
    .B(\fifo_t[1] ),
    .Y(_0410_));
 sg13g2_nor2b_2 _1898_ (.A(\fifo_t[1] ),
    .B_N(\fifo_t[0] ),
    .Y(_0411_));
 sg13g2_nor2b_2 _1899_ (.A(\fifo_t[0] ),
    .B_N(\fifo_t[1] ),
    .Y(_0412_));
 sg13g2_nor2_1 _1900_ (.A(_0409_),
    .B(_0410_),
    .Y(_0413_));
 sg13g2_nand2_1 _1901_ (.Y(_0414_),
    .A(\fifo_t[2] ),
    .B(_0409_));
 sg13g2_inv_1 _1902_ (.Y(_0415_),
    .A(_0414_));
 sg13g2_xor2_1 _1903_ (.B(_0409_),
    .A(_1227_),
    .X(_0416_));
 sg13g2_or2_1 _1904_ (.X(_0417_),
    .B(_1226_),
    .A(\fifo_t[0] ));
 sg13g2_xnor2_1 _1905_ (.Y(_0418_),
    .A(_1224_),
    .B(_0414_));
 sg13g2_a21oi_1 _1906_ (.A1(\fifo_t[0] ),
    .A2(_1226_),
    .Y(_0419_),
    .B1(_0418_));
 sg13g2_nand4_1 _1907_ (.B(_0416_),
    .C(_0417_),
    .A(_1225_),
    .Y(_0420_),
    .D(_0419_));
 sg13g2_and3_2 _1908_ (.X(_0421_),
    .A(_1208_),
    .B(_1214_),
    .C(_1221_));
 sg13g2_and3_1 _1909_ (.X(_0422_),
    .A(net719),
    .B(_0420_),
    .C(_0421_));
 sg13g2_mux2_1 _1910_ (.A0(\fifo_t[0] ),
    .A1(_0039_),
    .S(_0422_),
    .X(_0143_));
 sg13g2_mux2_1 _1911_ (.A0(\fifo_t[1] ),
    .A1(_0413_),
    .S(_0422_),
    .X(_0144_));
 sg13g2_nand4_1 _1912_ (.B(_0409_),
    .C(net731),
    .A(net719),
    .Y(_0423_),
    .D(net718));
 sg13g2_nand4_1 _1913_ (.B(_0415_),
    .C(net731),
    .A(net719),
    .Y(_0424_),
    .D(net718));
 sg13g2_a22oi_1 _1914_ (.Y(_0145_),
    .B1(_0423_),
    .B2(_1136_),
    .A2(_0422_),
    .A1(_0415_));
 sg13g2_xnor2_1 _1915_ (.Y(_0146_),
    .A(net819),
    .B(_0424_));
 sg13g2_nor2_2 _1916_ (.A(net821),
    .B(net819),
    .Y(_0425_));
 sg13g2_and2_1 _1917_ (.A(_0410_),
    .B(_0425_),
    .X(_0426_));
 sg13g2_and2_1 _1918_ (.A(\uart_0.rx.rx_samples[72] ),
    .B(\uart_0.rx.rx_samples[73] ),
    .X(_0427_));
 sg13g2_xor2_1 _1919_ (.B(\uart_0.rx.rx_samples[73] ),
    .A(\uart_0.rx.rx_samples[72] ),
    .X(_0428_));
 sg13g2_a21oi_1 _1920_ (.A1(\uart_0.rx.rx_samples[75] ),
    .A2(_0428_),
    .Y(_0429_),
    .B1(_0427_));
 sg13g2_xnor2_1 _1921_ (.Y(_0430_),
    .A(\uart_0.rx.rx_samples[75] ),
    .B(_0428_));
 sg13g2_inv_1 _1922_ (.Y(_0431_),
    .A(_0430_));
 sg13g2_xor2_1 _1923_ (.B(_0430_),
    .A(\uart_0.rx.rx_samples[80] ),
    .X(_0432_));
 sg13g2_nor2_1 _1924_ (.A(_1152_),
    .B(_0432_),
    .Y(_0433_));
 sg13g2_a21oi_1 _1925_ (.A1(\uart_0.rx.rx_samples[80] ),
    .A2(_0431_),
    .Y(_0434_),
    .B1(_0433_));
 sg13g2_nand2_1 _1926_ (.Y(_0435_),
    .A(_0429_),
    .B(_0434_));
 sg13g2_nand2_1 _1927_ (.Y(_0436_),
    .A(\uart_0.rx.rx_samples[79] ),
    .B(\uart_0.rx.rx_samples[74] ));
 sg13g2_or2_1 _1928_ (.X(_0437_),
    .B(_0434_),
    .A(_0429_));
 sg13g2_nand2b_1 _1929_ (.Y(_0438_),
    .B(_0437_),
    .A_N(\uart_0.rx.rx_samples[76] ));
 sg13g2_xnor2_1 _1930_ (.Y(_0439_),
    .A(\uart_0.rx.rx_samples[77] ),
    .B(_0432_));
 sg13g2_and2_1 _1931_ (.A(\uart_0.rx.rx_samples[78] ),
    .B(_0439_),
    .X(_0440_));
 sg13g2_nor2_1 _1932_ (.A(\uart_0.rx.rx_samples[79] ),
    .B(\uart_0.rx.rx_samples[74] ),
    .Y(_0441_));
 sg13g2_or2_1 _1933_ (.X(_0442_),
    .B(_0439_),
    .A(\uart_0.rx.rx_samples[78] ));
 sg13g2_o21ai_1 _1934_ (.B1(_0442_),
    .Y(_0443_),
    .A1(\uart_0.rx.rx_samples[76] ),
    .A2(_0440_));
 sg13g2_a21oi_1 _1935_ (.A1(_0437_),
    .A2(_0443_),
    .Y(_0444_),
    .B1(_0441_));
 sg13g2_nor2_1 _1936_ (.A(\uart_0.rx.rx_samples[76] ),
    .B(_0442_),
    .Y(_0445_));
 sg13g2_a21oi_1 _1937_ (.A1(_0436_),
    .A2(_0437_),
    .Y(_0446_),
    .B1(_0445_));
 sg13g2_nand3_1 _1938_ (.B(_0434_),
    .C(_0436_),
    .A(_0429_),
    .Y(_0447_));
 sg13g2_nand3_1 _1939_ (.B(_0440_),
    .C(_0447_),
    .A(_0438_),
    .Y(_0448_));
 sg13g2_o21ai_1 _1940_ (.B1(_0435_),
    .Y(_0449_),
    .A1(_0444_),
    .A2(_0446_));
 sg13g2_nand2_1 _1941_ (.Y(_0450_),
    .A(_0448_),
    .B(_0449_));
 sg13g2_nand4_1 _1942_ (.B(_0420_),
    .C(_0421_),
    .A(net720),
    .Y(_0451_),
    .D(_0450_));
 sg13g2_nor2_1 _1943_ (.A(\fifo_d[0][0] ),
    .B(net814),
    .Y(_0452_));
 sg13g2_a21oi_1 _1944_ (.A1(net814),
    .A2(net717),
    .Y(_0147_),
    .B1(_0452_));
 sg13g2_and2_1 _1945_ (.A(\uart_0.rx.rx_samples[63] ),
    .B(\uart_0.rx.rx_samples[64] ),
    .X(_0453_));
 sg13g2_xor2_1 _1946_ (.B(\uart_0.rx.rx_samples[64] ),
    .A(\uart_0.rx.rx_samples[63] ),
    .X(_0454_));
 sg13g2_xnor2_1 _1947_ (.Y(_0455_),
    .A(\uart_0.rx.rx_samples[66] ),
    .B(_0454_));
 sg13g2_inv_1 _1948_ (.Y(_0456_),
    .A(_0455_));
 sg13g2_xor2_1 _1949_ (.B(_0455_),
    .A(\uart_0.rx.rx_samples[71] ),
    .X(_0457_));
 sg13g2_nor2_1 _1950_ (.A(_1153_),
    .B(_0457_),
    .Y(_0458_));
 sg13g2_a21oi_1 _1951_ (.A1(\uart_0.rx.rx_samples[71] ),
    .A2(_0456_),
    .Y(_0459_),
    .B1(_0458_));
 sg13g2_a21oi_1 _1952_ (.A1(\uart_0.rx.rx_samples[66] ),
    .A2(_0454_),
    .Y(_0460_),
    .B1(_0453_));
 sg13g2_nand2_1 _1953_ (.Y(_0461_),
    .A(_0459_),
    .B(_0460_));
 sg13g2_nand2_1 _1954_ (.Y(_0462_),
    .A(\uart_0.rx.rx_samples[70] ),
    .B(\uart_0.rx.rx_samples[65] ));
 sg13g2_xnor2_1 _1955_ (.Y(_0463_),
    .A(\uart_0.rx.rx_samples[68] ),
    .B(_0457_));
 sg13g2_and2_1 _1956_ (.A(\uart_0.rx.rx_samples[69] ),
    .B(_0463_),
    .X(_0464_));
 sg13g2_or2_1 _1957_ (.X(_0465_),
    .B(_0460_),
    .A(_0459_));
 sg13g2_inv_1 _1958_ (.Y(_0466_),
    .A(_0465_));
 sg13g2_o21ai_1 _1959_ (.B1(_0464_),
    .Y(_0467_),
    .A1(\uart_0.rx.rx_samples[67] ),
    .A2(_0466_));
 sg13g2_nor2_1 _1960_ (.A(\uart_0.rx.rx_samples[70] ),
    .B(\uart_0.rx.rx_samples[65] ),
    .Y(_0468_));
 sg13g2_or2_1 _1961_ (.X(_0469_),
    .B(_0463_),
    .A(\uart_0.rx.rx_samples[69] ));
 sg13g2_o21ai_1 _1962_ (.B1(_0469_),
    .Y(_0470_),
    .A1(\uart_0.rx.rx_samples[67] ),
    .A2(_0464_));
 sg13g2_a21oi_1 _1963_ (.A1(_0465_),
    .A2(_0470_),
    .Y(_0471_),
    .B1(_0468_));
 sg13g2_nor2_1 _1964_ (.A(\uart_0.rx.rx_samples[67] ),
    .B(_0469_),
    .Y(_0472_));
 sg13g2_a21oi_1 _1965_ (.A1(_0462_),
    .A2(_0465_),
    .Y(_0473_),
    .B1(_0472_));
 sg13g2_o21ai_1 _1966_ (.B1(_0461_),
    .Y(_0474_),
    .A1(_0471_),
    .A2(_0473_));
 sg13g2_nor2b_1 _1967_ (.A(_0461_),
    .B_N(_0462_),
    .Y(_0475_));
 sg13g2_o21ai_1 _1968_ (.B1(_0474_),
    .Y(_0476_),
    .A1(_0467_),
    .A2(_0475_));
 sg13g2_nand4_1 _1969_ (.B(_0420_),
    .C(_0421_),
    .A(net720),
    .Y(_0477_),
    .D(_0476_));
 sg13g2_nor2_1 _1970_ (.A(\fifo_d[0][1] ),
    .B(net814),
    .Y(_0478_));
 sg13g2_a21oi_1 _1971_ (.A1(net814),
    .A2(net715),
    .Y(_0148_),
    .B1(_0478_));
 sg13g2_and2_1 _1972_ (.A(\uart_0.rx.rx_samples[54] ),
    .B(\uart_0.rx.rx_samples[55] ),
    .X(_0479_));
 sg13g2_xor2_1 _1973_ (.B(\uart_0.rx.rx_samples[55] ),
    .A(\uart_0.rx.rx_samples[54] ),
    .X(_0480_));
 sg13g2_and2_1 _1974_ (.A(\uart_0.rx.rx_samples[57] ),
    .B(_0480_),
    .X(_0481_));
 sg13g2_xnor2_1 _1975_ (.Y(_0482_),
    .A(\uart_0.rx.rx_samples[57] ),
    .B(_0480_));
 sg13g2_nor2_1 _1976_ (.A(_1154_),
    .B(_0482_),
    .Y(_0483_));
 sg13g2_nand2_1 _1977_ (.Y(_0484_),
    .A(_1154_),
    .B(_0482_));
 sg13g2_nand2b_1 _1978_ (.Y(_0485_),
    .B(_0484_),
    .A_N(_0483_));
 sg13g2_xnor2_1 _1979_ (.Y(_0486_),
    .A(\uart_0.rx.rx_samples[59] ),
    .B(_0485_));
 sg13g2_nand2_1 _1980_ (.Y(_0487_),
    .A(\uart_0.rx.rx_samples[60] ),
    .B(_0486_));
 sg13g2_a21o_1 _1981_ (.A2(_0484_),
    .A1(\uart_0.rx.rx_samples[59] ),
    .B1(_0483_),
    .X(_0488_));
 sg13g2_nor2_1 _1982_ (.A(_0479_),
    .B(_0481_),
    .Y(_0489_));
 sg13g2_o21ai_1 _1983_ (.B1(_0488_),
    .Y(_0490_),
    .A1(_0479_),
    .A2(_0481_));
 sg13g2_a21oi_1 _1984_ (.A1(_1155_),
    .A2(_0490_),
    .Y(_0491_),
    .B1(_0487_));
 sg13g2_and2_1 _1985_ (.A(\uart_0.rx.rx_samples[61] ),
    .B(\uart_0.rx.rx_samples[56] ),
    .X(_0492_));
 sg13g2_nand2_1 _1986_ (.Y(_0493_),
    .A(\uart_0.rx.rx_samples[61] ),
    .B(\uart_0.rx.rx_samples[56] ));
 sg13g2_a21oi_1 _1987_ (.A1(_0491_),
    .A2(_0492_),
    .Y(_0494_),
    .B1(_0488_));
 sg13g2_nor2_1 _1988_ (.A(\uart_0.rx.rx_samples[60] ),
    .B(_0486_),
    .Y(_0495_));
 sg13g2_o21ai_1 _1989_ (.B1(\uart_0.rx.rx_samples[58] ),
    .Y(_0496_),
    .A1(\uart_0.rx.rx_samples[60] ),
    .A2(_0486_));
 sg13g2_nand3_1 _1990_ (.B(_0490_),
    .C(_0496_),
    .A(_0487_),
    .Y(_0497_));
 sg13g2_o21ai_1 _1991_ (.B1(_0497_),
    .Y(_0498_),
    .A1(\uart_0.rx.rx_samples[61] ),
    .A2(\uart_0.rx.rx_samples[56] ));
 sg13g2_a22oi_1 _1992_ (.Y(_0499_),
    .B1(_0495_),
    .B2(_1155_),
    .A2(_0493_),
    .A1(_0490_));
 sg13g2_nor2_1 _1993_ (.A(_0491_),
    .B(_0499_),
    .Y(_0500_));
 sg13g2_a22oi_1 _1994_ (.Y(_0501_),
    .B1(_0498_),
    .B2(_0500_),
    .A2(_0494_),
    .A1(_0489_));
 sg13g2_nand4_1 _1995_ (.B(net731),
    .C(net718),
    .A(net719),
    .Y(_0502_),
    .D(_0501_));
 sg13g2_nor2_1 _1996_ (.A(\fifo_d[0][2] ),
    .B(net814),
    .Y(_0503_));
 sg13g2_a21oi_1 _1997_ (.A1(net814),
    .A2(net713),
    .Y(_0149_),
    .B1(_0503_));
 sg13g2_and2_1 _1998_ (.A(\uart_0.rx.rx_samples[45] ),
    .B(\uart_0.rx.rx_samples[46] ),
    .X(_0504_));
 sg13g2_xor2_1 _1999_ (.B(\uart_0.rx.rx_samples[46] ),
    .A(\uart_0.rx.rx_samples[45] ),
    .X(_0505_));
 sg13g2_xnor2_1 _2000_ (.Y(_0506_),
    .A(\uart_0.rx.rx_samples[48] ),
    .B(_0505_));
 sg13g2_nor2_1 _2001_ (.A(_1156_),
    .B(_0506_),
    .Y(_0507_));
 sg13g2_xnor2_1 _2002_ (.Y(_0508_),
    .A(\uart_0.rx.rx_samples[53] ),
    .B(_0506_));
 sg13g2_a21oi_1 _2003_ (.A1(\uart_0.rx.rx_samples[50] ),
    .A2(_0508_),
    .Y(_0509_),
    .B1(_0507_));
 sg13g2_a21oi_1 _2004_ (.A1(\uart_0.rx.rx_samples[48] ),
    .A2(_0505_),
    .Y(_0510_),
    .B1(_0504_));
 sg13g2_nor2_1 _2005_ (.A(\uart_0.rx.rx_samples[52] ),
    .B(\uart_0.rx.rx_samples[47] ),
    .Y(_0511_));
 sg13g2_xnor2_1 _2006_ (.Y(_0512_),
    .A(\uart_0.rx.rx_samples[50] ),
    .B(_0508_));
 sg13g2_nand2_1 _2007_ (.Y(_0513_),
    .A(_1157_),
    .B(_0512_));
 sg13g2_or2_1 _2008_ (.X(_0514_),
    .B(_0510_),
    .A(_0509_));
 sg13g2_nor2_1 _2009_ (.A(_1157_),
    .B(_0512_),
    .Y(_0515_));
 sg13g2_o21ai_1 _2010_ (.B1(_0513_),
    .Y(_0516_),
    .A1(\uart_0.rx.rx_samples[49] ),
    .A2(_0515_));
 sg13g2_a21o_1 _2011_ (.A2(_0516_),
    .A1(_0514_),
    .B1(_0511_),
    .X(_0517_));
 sg13g2_nand2_1 _2012_ (.Y(_0518_),
    .A(\uart_0.rx.rx_samples[52] ),
    .B(\uart_0.rx.rx_samples[47] ));
 sg13g2_nand2_1 _2013_ (.Y(_0519_),
    .A(_0514_),
    .B(_0518_));
 sg13g2_o21ai_1 _2014_ (.B1(_0519_),
    .Y(_0520_),
    .A1(\uart_0.rx.rx_samples[49] ),
    .A2(_0513_));
 sg13g2_a22oi_1 _2015_ (.Y(_0521_),
    .B1(_0517_),
    .B2(_0520_),
    .A2(_0510_),
    .A1(_0509_));
 sg13g2_nand2b_1 _2016_ (.Y(_0522_),
    .B(_0514_),
    .A_N(\uart_0.rx.rx_samples[49] ));
 sg13g2_nand3_1 _2017_ (.B(_0510_),
    .C(_0518_),
    .A(_0509_),
    .Y(_0523_));
 sg13g2_nand3_1 _2018_ (.B(_0522_),
    .C(_0523_),
    .A(_0515_),
    .Y(_0524_));
 sg13g2_nand2b_1 _2019_ (.Y(_0525_),
    .B(_0524_),
    .A_N(_0521_));
 sg13g2_nand4_1 _2020_ (.B(net731),
    .C(net718),
    .A(net719),
    .Y(_0526_),
    .D(_0525_));
 sg13g2_nor2_1 _2021_ (.A(\fifo_d[0][3] ),
    .B(net813),
    .Y(_0527_));
 sg13g2_a21oi_1 _2022_ (.A1(net813),
    .A2(net710),
    .Y(_0150_),
    .B1(_0527_));
 sg13g2_and2_1 _2023_ (.A(\uart_0.rx.rx_samples[36] ),
    .B(\uart_0.rx.rx_samples[37] ),
    .X(_0528_));
 sg13g2_xor2_1 _2024_ (.B(\uart_0.rx.rx_samples[37] ),
    .A(\uart_0.rx.rx_samples[36] ),
    .X(_0529_));
 sg13g2_a21oi_1 _2025_ (.A1(\uart_0.rx.rx_samples[39] ),
    .A2(_0529_),
    .Y(_0530_),
    .B1(_0528_));
 sg13g2_xnor2_1 _2026_ (.Y(_0531_),
    .A(\uart_0.rx.rx_samples[39] ),
    .B(_0529_));
 sg13g2_nor2_1 _2027_ (.A(_1158_),
    .B(_0531_),
    .Y(_0532_));
 sg13g2_nand2_1 _2028_ (.Y(_0533_),
    .A(_1158_),
    .B(_0531_));
 sg13g2_nand2b_1 _2029_ (.Y(_0534_),
    .B(_0533_),
    .A_N(_0532_));
 sg13g2_a21oi_1 _2030_ (.A1(\uart_0.rx.rx_samples[41] ),
    .A2(_0533_),
    .Y(_0535_),
    .B1(_0532_));
 sg13g2_and2_1 _2031_ (.A(_0530_),
    .B(_0535_),
    .X(_0536_));
 sg13g2_nand2_1 _2032_ (.Y(_0537_),
    .A(\uart_0.rx.rx_samples[43] ),
    .B(\uart_0.rx.rx_samples[38] ));
 sg13g2_xnor2_1 _2033_ (.Y(_0538_),
    .A(\uart_0.rx.rx_samples[41] ),
    .B(_0534_));
 sg13g2_nand2_1 _2034_ (.Y(_0539_),
    .A(\uart_0.rx.rx_samples[42] ),
    .B(_0538_));
 sg13g2_or2_1 _2035_ (.X(_0540_),
    .B(_0535_),
    .A(_0530_));
 sg13g2_a21oi_1 _2036_ (.A1(_1159_),
    .A2(_0540_),
    .Y(_0541_),
    .B1(_0539_));
 sg13g2_nand2b_1 _2037_ (.Y(_0542_),
    .B(_0541_),
    .A_N(_0537_));
 sg13g2_nor2_1 _2038_ (.A(\uart_0.rx.rx_samples[42] ),
    .B(_0538_),
    .Y(_0543_));
 sg13g2_o21ai_1 _2039_ (.B1(\uart_0.rx.rx_samples[40] ),
    .Y(_0544_),
    .A1(\uart_0.rx.rx_samples[42] ),
    .A2(_0538_));
 sg13g2_nand3_1 _2040_ (.B(_0540_),
    .C(_0544_),
    .A(_0539_),
    .Y(_0545_));
 sg13g2_o21ai_1 _2041_ (.B1(_0545_),
    .Y(_0546_),
    .A1(\uart_0.rx.rx_samples[43] ),
    .A2(\uart_0.rx.rx_samples[38] ));
 sg13g2_a22oi_1 _2042_ (.Y(_0547_),
    .B1(_0543_),
    .B2(_1159_),
    .A2(_0540_),
    .A1(_0537_));
 sg13g2_nor2_1 _2043_ (.A(_0541_),
    .B(_0547_),
    .Y(_0548_));
 sg13g2_a22oi_1 _2044_ (.Y(_0549_),
    .B1(_0546_),
    .B2(_0548_),
    .A2(_0542_),
    .A1(_0536_));
 sg13g2_nand4_1 _2045_ (.B(net731),
    .C(net718),
    .A(net719),
    .Y(_0550_),
    .D(_0549_));
 sg13g2_nor2_1 _2046_ (.A(\fifo_d[0][4] ),
    .B(net814),
    .Y(_0551_));
 sg13g2_a21oi_1 _2047_ (.A1(net814),
    .A2(_0550_),
    .Y(_0151_),
    .B1(_0551_));
 sg13g2_and2_1 _2048_ (.A(\uart_0.rx.rx_samples[27] ),
    .B(\uart_0.rx.rx_samples[28] ),
    .X(_0552_));
 sg13g2_xor2_1 _2049_ (.B(\uart_0.rx.rx_samples[28] ),
    .A(\uart_0.rx.rx_samples[27] ),
    .X(_0553_));
 sg13g2_a21oi_1 _2050_ (.A1(\uart_0.rx.rx_samples[30] ),
    .A2(_0553_),
    .Y(_0554_),
    .B1(_0552_));
 sg13g2_xnor2_1 _2051_ (.Y(_0555_),
    .A(\uart_0.rx.rx_samples[30] ),
    .B(_0553_));
 sg13g2_nor2_1 _2052_ (.A(_1160_),
    .B(_0555_),
    .Y(_0556_));
 sg13g2_nand2_1 _2053_ (.Y(_0557_),
    .A(_1160_),
    .B(_0555_));
 sg13g2_nand2b_1 _2054_ (.Y(_0558_),
    .B(_0557_),
    .A_N(_0556_));
 sg13g2_a21oi_1 _2055_ (.A1(\uart_0.rx.rx_samples[32] ),
    .A2(_0557_),
    .Y(_0559_),
    .B1(_0556_));
 sg13g2_and2_1 _2056_ (.A(_0554_),
    .B(_0559_),
    .X(_0560_));
 sg13g2_nand2_1 _2057_ (.Y(_0561_),
    .A(\uart_0.rx.rx_samples[34] ),
    .B(\uart_0.rx.rx_samples[29] ));
 sg13g2_xnor2_1 _2058_ (.Y(_0562_),
    .A(\uart_0.rx.rx_samples[32] ),
    .B(_0558_));
 sg13g2_nand2_1 _2059_ (.Y(_0563_),
    .A(\uart_0.rx.rx_samples[33] ),
    .B(_0562_));
 sg13g2_or2_1 _2060_ (.X(_0564_),
    .B(_0559_),
    .A(_0554_));
 sg13g2_a21oi_1 _2061_ (.A1(_1161_),
    .A2(_0564_),
    .Y(_0565_),
    .B1(_0563_));
 sg13g2_nand2b_1 _2062_ (.Y(_0566_),
    .B(_0565_),
    .A_N(_0561_));
 sg13g2_nor2_1 _2063_ (.A(\uart_0.rx.rx_samples[33] ),
    .B(_0562_),
    .Y(_0567_));
 sg13g2_o21ai_1 _2064_ (.B1(\uart_0.rx.rx_samples[31] ),
    .Y(_0568_),
    .A1(\uart_0.rx.rx_samples[33] ),
    .A2(_0562_));
 sg13g2_nand3_1 _2065_ (.B(_0564_),
    .C(_0568_),
    .A(_0563_),
    .Y(_0569_));
 sg13g2_o21ai_1 _2066_ (.B1(_0569_),
    .Y(_0570_),
    .A1(\uart_0.rx.rx_samples[34] ),
    .A2(\uart_0.rx.rx_samples[29] ));
 sg13g2_a22oi_1 _2067_ (.Y(_0571_),
    .B1(_0567_),
    .B2(_1161_),
    .A2(_0564_),
    .A1(_0561_));
 sg13g2_nor2_1 _2068_ (.A(_0565_),
    .B(_0571_),
    .Y(_0572_));
 sg13g2_a22oi_1 _2069_ (.Y(_0573_),
    .B1(_0570_),
    .B2(_0572_),
    .A2(_0566_),
    .A1(_0560_));
 sg13g2_nand4_1 _2070_ (.B(net731),
    .C(net718),
    .A(net719),
    .Y(_0574_),
    .D(_0573_));
 sg13g2_nor2_1 _2071_ (.A(\fifo_d[0][5] ),
    .B(net813),
    .Y(_0575_));
 sg13g2_a21oi_1 _2072_ (.A1(net813),
    .A2(net706),
    .Y(_0152_),
    .B1(_0575_));
 sg13g2_and2_1 _2073_ (.A(\uart_0.rx.rx_samples[18] ),
    .B(\uart_0.rx.rx_samples[19] ),
    .X(_0576_));
 sg13g2_xor2_1 _2074_ (.B(\uart_0.rx.rx_samples[19] ),
    .A(\uart_0.rx.rx_samples[18] ),
    .X(_0577_));
 sg13g2_a21oi_1 _2075_ (.A1(\uart_0.rx.rx_samples[21] ),
    .A2(_0577_),
    .Y(_0578_),
    .B1(_0576_));
 sg13g2_xnor2_1 _2076_ (.Y(_0579_),
    .A(\uart_0.rx.rx_samples[21] ),
    .B(_0577_));
 sg13g2_inv_1 _2077_ (.Y(_0580_),
    .A(_0579_));
 sg13g2_xor2_1 _2078_ (.B(_0579_),
    .A(\uart_0.rx.rx_samples[26] ),
    .X(_0581_));
 sg13g2_nor2_1 _2079_ (.A(_1162_),
    .B(_0581_),
    .Y(_0582_));
 sg13g2_a21oi_1 _2080_ (.A1(\uart_0.rx.rx_samples[26] ),
    .A2(_0580_),
    .Y(_0583_),
    .B1(_0582_));
 sg13g2_nand2_1 _2081_ (.Y(_0584_),
    .A(_0578_),
    .B(_0583_));
 sg13g2_nand2_1 _2082_ (.Y(_0585_),
    .A(\uart_0.rx.rx_samples[25] ),
    .B(\uart_0.rx.rx_samples[20] ));
 sg13g2_xnor2_1 _2083_ (.Y(_0586_),
    .A(\uart_0.rx.rx_samples[23] ),
    .B(_0581_));
 sg13g2_and2_1 _2084_ (.A(\uart_0.rx.rx_samples[24] ),
    .B(_0586_),
    .X(_0587_));
 sg13g2_or2_1 _2085_ (.X(_0588_),
    .B(_0583_),
    .A(_0578_));
 sg13g2_inv_1 _2086_ (.Y(_0589_),
    .A(_0588_));
 sg13g2_o21ai_1 _2087_ (.B1(_0587_),
    .Y(_0590_),
    .A1(\uart_0.rx.rx_samples[22] ),
    .A2(_0589_));
 sg13g2_nor2_1 _2088_ (.A(\uart_0.rx.rx_samples[25] ),
    .B(\uart_0.rx.rx_samples[20] ),
    .Y(_0591_));
 sg13g2_or2_1 _2089_ (.X(_0592_),
    .B(_0586_),
    .A(\uart_0.rx.rx_samples[24] ));
 sg13g2_o21ai_1 _2090_ (.B1(_0592_),
    .Y(_0593_),
    .A1(\uart_0.rx.rx_samples[22] ),
    .A2(_0587_));
 sg13g2_a21oi_1 _2091_ (.A1(_0588_),
    .A2(_0593_),
    .Y(_0594_),
    .B1(_0591_));
 sg13g2_nor2_1 _2092_ (.A(\uart_0.rx.rx_samples[22] ),
    .B(_0592_),
    .Y(_0595_));
 sg13g2_a21oi_1 _2093_ (.A1(_0585_),
    .A2(_0588_),
    .Y(_0596_),
    .B1(_0595_));
 sg13g2_nor2b_1 _2094_ (.A(_0584_),
    .B_N(_0585_),
    .Y(_0597_));
 sg13g2_o21ai_1 _2095_ (.B1(_0584_),
    .Y(_0598_),
    .A1(_0594_),
    .A2(_0596_));
 sg13g2_o21ai_1 _2096_ (.B1(_0598_),
    .Y(_0599_),
    .A1(_0590_),
    .A2(_0597_));
 sg13g2_nand4_1 _2097_ (.B(net731),
    .C(net718),
    .A(net720),
    .Y(_0600_),
    .D(_0599_));
 sg13g2_nor2_1 _2098_ (.A(\fifo_d[0][6] ),
    .B(net813),
    .Y(_0601_));
 sg13g2_a21oi_1 _2099_ (.A1(net813),
    .A2(net704),
    .Y(_0153_),
    .B1(_0601_));
 sg13g2_nor2_1 _2100_ (.A(\uart_0.rx.rx_samples[16] ),
    .B(\uart_0.rx.rx_samples[11] ),
    .Y(_0602_));
 sg13g2_and2_1 _2101_ (.A(\uart_0.rx.rx_samples[9] ),
    .B(\uart_0.rx.rx_samples[10] ),
    .X(_0603_));
 sg13g2_xor2_1 _2102_ (.B(\uart_0.rx.rx_samples[10] ),
    .A(\uart_0.rx.rx_samples[9] ),
    .X(_0604_));
 sg13g2_xor2_1 _2103_ (.B(_0604_),
    .A(\uart_0.rx.rx_samples[12] ),
    .X(_0605_));
 sg13g2_and2_1 _2104_ (.A(\uart_0.rx.rx_samples[17] ),
    .B(_0605_),
    .X(_0606_));
 sg13g2_xor2_1 _2105_ (.B(_0605_),
    .A(\uart_0.rx.rx_samples[17] ),
    .X(_0607_));
 sg13g2_xnor2_1 _2106_ (.Y(_0608_),
    .A(\uart_0.rx.rx_samples[14] ),
    .B(_0607_));
 sg13g2_and2_1 _2107_ (.A(_1163_),
    .B(_0608_),
    .X(_0609_));
 sg13g2_or2_1 _2108_ (.X(_0610_),
    .B(_0608_),
    .A(_1163_));
 sg13g2_a21o_1 _2109_ (.A2(_0607_),
    .A1(\uart_0.rx.rx_samples[14] ),
    .B1(_0606_),
    .X(_0611_));
 sg13g2_a21o_1 _2110_ (.A2(_0604_),
    .A1(\uart_0.rx.rx_samples[12] ),
    .B1(_0603_),
    .X(_0612_));
 sg13g2_nand2_1 _2111_ (.Y(_0613_),
    .A(_0611_),
    .B(_0612_));
 sg13g2_a21o_1 _2112_ (.A2(_0610_),
    .A1(_1164_),
    .B1(_0609_),
    .X(_0614_));
 sg13g2_a21oi_1 _2113_ (.A1(_0613_),
    .A2(_0614_),
    .Y(_0615_),
    .B1(_0602_));
 sg13g2_a21o_1 _2114_ (.A2(_0613_),
    .A1(_1164_),
    .B1(_0610_),
    .X(_0616_));
 sg13g2_nand2_1 _2115_ (.Y(_0617_),
    .A(\uart_0.rx.rx_samples[16] ),
    .B(\uart_0.rx.rx_samples[11] ));
 sg13g2_a22oi_1 _2116_ (.Y(_0618_),
    .B1(_0613_),
    .B2(_0617_),
    .A2(_0609_),
    .A1(_1164_));
 sg13g2_nor2_1 _2117_ (.A(_0615_),
    .B(_0618_),
    .Y(_0619_));
 sg13g2_nor2_1 _2118_ (.A(_0616_),
    .B(_0617_),
    .Y(_0620_));
 sg13g2_nor3_1 _2119_ (.A(_0611_),
    .B(_0612_),
    .C(_0620_),
    .Y(_0621_));
 sg13g2_a21oi_2 _2120_ (.B1(_0621_),
    .Y(_0622_),
    .A2(_0619_),
    .A1(_0616_));
 sg13g2_nand4_1 _2121_ (.B(net731),
    .C(net718),
    .A(net719),
    .Y(_0623_),
    .D(_0622_));
 sg13g2_nor2_1 _2122_ (.A(\fifo_d[0][7] ),
    .B(net813),
    .Y(_0624_));
 sg13g2_a21oi_1 _2123_ (.A1(net813),
    .A2(net702),
    .Y(_0154_),
    .B1(_0624_));
 sg13g2_nand2_1 _2124_ (.Y(_0625_),
    .A(_0411_),
    .B(_0425_));
 sg13g2_nand2_1 _2125_ (.Y(_0626_),
    .A(\fifo_d[1][0] ),
    .B(net811));
 sg13g2_o21ai_1 _2126_ (.B1(_0626_),
    .Y(_0155_),
    .A1(net716),
    .A2(net811));
 sg13g2_nand2_1 _2127_ (.Y(_0627_),
    .A(\fifo_d[1][1] ),
    .B(net811));
 sg13g2_o21ai_1 _2128_ (.B1(_0627_),
    .Y(_0156_),
    .A1(net714),
    .A2(net811));
 sg13g2_nand2_1 _2129_ (.Y(_0628_),
    .A(\fifo_d[1][2] ),
    .B(net811));
 sg13g2_o21ai_1 _2130_ (.B1(_0628_),
    .Y(_0157_),
    .A1(net712),
    .A2(net811));
 sg13g2_nand2_1 _2131_ (.Y(_0629_),
    .A(\fifo_d[1][3] ),
    .B(net812));
 sg13g2_o21ai_1 _2132_ (.B1(_0629_),
    .Y(_0158_),
    .A1(net711),
    .A2(net812));
 sg13g2_nand2_1 _2133_ (.Y(_0630_),
    .A(\fifo_d[1][4] ),
    .B(net812));
 sg13g2_o21ai_1 _2134_ (.B1(_0630_),
    .Y(_0159_),
    .A1(net708),
    .A2(_0625_));
 sg13g2_nand2_1 _2135_ (.Y(_0631_),
    .A(\fifo_d[1][5] ),
    .B(net812));
 sg13g2_o21ai_1 _2136_ (.B1(_0631_),
    .Y(_0160_),
    .A1(_0574_),
    .A2(net812));
 sg13g2_nand2_1 _2137_ (.Y(_0632_),
    .A(\fifo_d[1][6] ),
    .B(net811));
 sg13g2_o21ai_1 _2138_ (.B1(_0632_),
    .Y(_0161_),
    .A1(net705),
    .A2(net811));
 sg13g2_nand2_1 _2139_ (.Y(_0633_),
    .A(\fifo_d[1][7] ),
    .B(net812));
 sg13g2_o21ai_1 _2140_ (.B1(_0633_),
    .Y(_0162_),
    .A1(net701),
    .A2(net812));
 sg13g2_nand2_1 _2141_ (.Y(_0634_),
    .A(_0412_),
    .B(_0425_));
 sg13g2_nand2_1 _2142_ (.Y(_0635_),
    .A(\fifo_d[2][0] ),
    .B(net809));
 sg13g2_o21ai_1 _2143_ (.B1(_0635_),
    .Y(_0163_),
    .A1(net716),
    .A2(net809));
 sg13g2_nand2_1 _2144_ (.Y(_0636_),
    .A(\fifo_d[2][1] ),
    .B(net810));
 sg13g2_o21ai_1 _2145_ (.B1(_0636_),
    .Y(_0164_),
    .A1(net715),
    .A2(net810));
 sg13g2_nand2_1 _2146_ (.Y(_0637_),
    .A(\fifo_d[2][2] ),
    .B(net810));
 sg13g2_o21ai_1 _2147_ (.B1(_0637_),
    .Y(_0165_),
    .A1(net713),
    .A2(net810));
 sg13g2_nand2_1 _2148_ (.Y(_0638_),
    .A(\fifo_d[2][3] ),
    .B(net809));
 sg13g2_o21ai_1 _2149_ (.B1(_0638_),
    .Y(_0166_),
    .A1(net711),
    .A2(net809));
 sg13g2_nand2_1 _2150_ (.Y(_0639_),
    .A(\fifo_d[2][4] ),
    .B(net809));
 sg13g2_o21ai_1 _2151_ (.B1(_0639_),
    .Y(_0167_),
    .A1(net709),
    .A2(net809));
 sg13g2_nand2_1 _2152_ (.Y(_0640_),
    .A(\fifo_d[2][5] ),
    .B(net809));
 sg13g2_o21ai_1 _2153_ (.B1(_0640_),
    .Y(_0168_),
    .A1(net707),
    .A2(net809));
 sg13g2_nand2_1 _2154_ (.Y(_0641_),
    .A(\fifo_d[2][6] ),
    .B(net810));
 sg13g2_o21ai_1 _2155_ (.B1(_0641_),
    .Y(_0169_),
    .A1(net704),
    .A2(net810));
 sg13g2_nand2_1 _2156_ (.Y(_0642_),
    .A(\fifo_d[2][7] ),
    .B(net810));
 sg13g2_o21ai_1 _2157_ (.B1(_0642_),
    .Y(_0170_),
    .A1(net702),
    .A2(net810));
 sg13g2_nand2_2 _2158_ (.Y(_0643_),
    .A(_0409_),
    .B(_0425_));
 sg13g2_nand2_1 _2159_ (.Y(_0644_),
    .A(\fifo_d[3][0] ),
    .B(_0643_));
 sg13g2_o21ai_1 _2160_ (.B1(_0644_),
    .Y(_0171_),
    .A1(net717),
    .A2(net808));
 sg13g2_nand2_1 _2161_ (.Y(_0645_),
    .A(\fifo_d[3][1] ),
    .B(net807));
 sg13g2_o21ai_1 _2162_ (.B1(_0645_),
    .Y(_0172_),
    .A1(net714),
    .A2(net807));
 sg13g2_nand2_1 _2163_ (.Y(_0646_),
    .A(\fifo_d[3][2] ),
    .B(net807));
 sg13g2_o21ai_1 _2164_ (.B1(_0646_),
    .Y(_0173_),
    .A1(net712),
    .A2(net807));
 sg13g2_nand2_1 _2165_ (.Y(_0647_),
    .A(\fifo_d[3][3] ),
    .B(net808));
 sg13g2_o21ai_1 _2166_ (.B1(_0647_),
    .Y(_0174_),
    .A1(net710),
    .A2(net808));
 sg13g2_nand2_1 _2167_ (.Y(_0648_),
    .A(\fifo_d[3][4] ),
    .B(net807));
 sg13g2_o21ai_1 _2168_ (.B1(_0648_),
    .Y(_0175_),
    .A1(net709),
    .A2(net807));
 sg13g2_nand2_1 _2169_ (.Y(_0649_),
    .A(\fifo_d[3][5] ),
    .B(net808));
 sg13g2_o21ai_1 _2170_ (.B1(_0649_),
    .Y(_0176_),
    .A1(net707),
    .A2(net808));
 sg13g2_nand2_1 _2171_ (.Y(_0650_),
    .A(\fifo_d[3][6] ),
    .B(net807));
 sg13g2_o21ai_1 _2172_ (.B1(_0650_),
    .Y(_0177_),
    .A1(net705),
    .A2(net807));
 sg13g2_nand2_1 _2173_ (.Y(_0651_),
    .A(\fifo_d[3][7] ),
    .B(net808));
 sg13g2_o21ai_1 _2174_ (.B1(_0651_),
    .Y(_0178_),
    .A1(net702),
    .A2(net808));
 sg13g2_nand3b_1 _2175_ (.B(_0410_),
    .C(net821),
    .Y(_0652_),
    .A_N(net819));
 sg13g2_nand2_1 _2176_ (.Y(_0653_),
    .A(\fifo_d[4][0] ),
    .B(net805));
 sg13g2_o21ai_1 _2177_ (.B1(_0653_),
    .Y(_0179_),
    .A1(net716),
    .A2(net805));
 sg13g2_nand2_1 _2178_ (.Y(_0654_),
    .A(\fifo_d[4][1] ),
    .B(net805));
 sg13g2_o21ai_1 _2179_ (.B1(_0654_),
    .Y(_0180_),
    .A1(net714),
    .A2(net805));
 sg13g2_nand2_1 _2180_ (.Y(_0655_),
    .A(\fifo_d[4][2] ),
    .B(net804));
 sg13g2_o21ai_1 _2181_ (.B1(_0655_),
    .Y(_0181_),
    .A1(net712),
    .A2(net804));
 sg13g2_nand2_1 _2182_ (.Y(_0656_),
    .A(\fifo_d[4][3] ),
    .B(net806));
 sg13g2_o21ai_1 _2183_ (.B1(_0656_),
    .Y(_0182_),
    .A1(net711),
    .A2(net806));
 sg13g2_nand2_1 _2184_ (.Y(_0657_),
    .A(\fifo_d[4][4] ),
    .B(net804));
 sg13g2_o21ai_1 _2185_ (.B1(_0657_),
    .Y(_0183_),
    .A1(net709),
    .A2(net804));
 sg13g2_nand2_1 _2186_ (.Y(_0658_),
    .A(\fifo_d[4][5] ),
    .B(net806));
 sg13g2_o21ai_1 _2187_ (.B1(_0658_),
    .Y(_0184_),
    .A1(net707),
    .A2(net806));
 sg13g2_nand2_1 _2188_ (.Y(_0659_),
    .A(\fifo_d[4][6] ),
    .B(net804));
 sg13g2_o21ai_1 _2189_ (.B1(_0659_),
    .Y(_0185_),
    .A1(net705),
    .A2(net804));
 sg13g2_nand2_1 _2190_ (.Y(_0660_),
    .A(\fifo_d[4][7] ),
    .B(net804));
 sg13g2_o21ai_1 _2191_ (.B1(_0660_),
    .Y(_0186_),
    .A1(net701),
    .A2(net804));
 sg13g2_nand2_1 _2192_ (.Y(_0661_),
    .A(net821),
    .B(_0411_));
 sg13g2_nor2_1 _2193_ (.A(net819),
    .B(_0661_),
    .Y(_0662_));
 sg13g2_nor2_1 _2194_ (.A(\fifo_d[5][0] ),
    .B(net780),
    .Y(_0663_));
 sg13g2_a21oi_1 _2195_ (.A1(net716),
    .A2(net780),
    .Y(_0187_),
    .B1(_0663_));
 sg13g2_nor2_1 _2196_ (.A(\fifo_d[5][1] ),
    .B(net781),
    .Y(_0664_));
 sg13g2_a21oi_1 _2197_ (.A1(net715),
    .A2(net781),
    .Y(_0188_),
    .B1(_0664_));
 sg13g2_nor2_1 _2198_ (.A(\fifo_d[5][2] ),
    .B(net781),
    .Y(_0665_));
 sg13g2_a21oi_1 _2199_ (.A1(net713),
    .A2(net781),
    .Y(_0189_),
    .B1(_0665_));
 sg13g2_nor2_1 _2200_ (.A(\fifo_d[5][3] ),
    .B(net781),
    .Y(_0666_));
 sg13g2_a21oi_1 _2201_ (.A1(net711),
    .A2(net781),
    .Y(_0190_),
    .B1(_0666_));
 sg13g2_nor2_1 _2202_ (.A(\fifo_d[5][4] ),
    .B(net780),
    .Y(_0667_));
 sg13g2_a21oi_1 _2203_ (.A1(net709),
    .A2(net780),
    .Y(_0191_),
    .B1(_0667_));
 sg13g2_nor2_1 _2204_ (.A(\fifo_d[5][5] ),
    .B(_0662_),
    .Y(_0668_));
 sg13g2_a21oi_1 _2205_ (.A1(net706),
    .A2(net781),
    .Y(_0192_),
    .B1(_0668_));
 sg13g2_nor2_1 _2206_ (.A(\fifo_d[5][6] ),
    .B(net780),
    .Y(_0669_));
 sg13g2_a21oi_1 _2207_ (.A1(net703),
    .A2(net780),
    .Y(_0193_),
    .B1(_0669_));
 sg13g2_nor2_1 _2208_ (.A(\fifo_d[5][7] ),
    .B(net780),
    .Y(_0670_));
 sg13g2_a21oi_1 _2209_ (.A1(net701),
    .A2(net780),
    .Y(_0194_),
    .B1(_0670_));
 sg13g2_nand2_1 _2210_ (.Y(_0671_),
    .A(net821),
    .B(_0412_));
 sg13g2_nor2_2 _2211_ (.A(net820),
    .B(_0671_),
    .Y(_0672_));
 sg13g2_nor2_1 _2212_ (.A(\fifo_d[6][0] ),
    .B(net778),
    .Y(_0673_));
 sg13g2_a21oi_1 _2213_ (.A1(net717),
    .A2(net778),
    .Y(_0195_),
    .B1(_0673_));
 sg13g2_nor2_1 _2214_ (.A(\fifo_d[6][1] ),
    .B(net778),
    .Y(_0674_));
 sg13g2_a21oi_1 _2215_ (.A1(net715),
    .A2(net778),
    .Y(_0196_),
    .B1(_0674_));
 sg13g2_nor2_1 _2216_ (.A(\fifo_d[6][2] ),
    .B(net778),
    .Y(_0675_));
 sg13g2_a21oi_1 _2217_ (.A1(net713),
    .A2(_0672_),
    .Y(_0197_),
    .B1(_0675_));
 sg13g2_nor2_1 _2218_ (.A(\fifo_d[6][3] ),
    .B(net778),
    .Y(_0676_));
 sg13g2_a21oi_1 _2219_ (.A1(net710),
    .A2(net779),
    .Y(_0198_),
    .B1(_0676_));
 sg13g2_nor2_1 _2220_ (.A(\fifo_d[6][4] ),
    .B(net779),
    .Y(_0677_));
 sg13g2_a21oi_1 _2221_ (.A1(net708),
    .A2(net779),
    .Y(_0199_),
    .B1(_0677_));
 sg13g2_nor2_1 _2222_ (.A(\fifo_d[6][5] ),
    .B(net779),
    .Y(_0678_));
 sg13g2_a21oi_1 _2223_ (.A1(net706),
    .A2(net779),
    .Y(_0200_),
    .B1(_0678_));
 sg13g2_nor2_1 _2224_ (.A(\fifo_d[6][6] ),
    .B(net779),
    .Y(_0679_));
 sg13g2_a21oi_1 _2225_ (.A1(net704),
    .A2(net779),
    .Y(_0201_),
    .B1(_0679_));
 sg13g2_nor2_1 _2226_ (.A(\fifo_d[6][7] ),
    .B(net778),
    .Y(_0680_));
 sg13g2_a21oi_1 _2227_ (.A1(net702),
    .A2(net778),
    .Y(_0202_),
    .B1(_0680_));
 sg13g2_nor2_1 _2228_ (.A(net819),
    .B(_0414_),
    .Y(_0681_));
 sg13g2_nor2_1 _2229_ (.A(\fifo_d[7][0] ),
    .B(net776),
    .Y(_0682_));
 sg13g2_a21oi_1 _2230_ (.A1(net717),
    .A2(net775),
    .Y(_0203_),
    .B1(_0682_));
 sg13g2_nor2_1 _2231_ (.A(\fifo_d[7][1] ),
    .B(net776),
    .Y(_0683_));
 sg13g2_a21oi_1 _2232_ (.A1(net715),
    .A2(net775),
    .Y(_0204_),
    .B1(_0683_));
 sg13g2_nor2_1 _2233_ (.A(\fifo_d[7][2] ),
    .B(net776),
    .Y(_0684_));
 sg13g2_a21oi_1 _2234_ (.A1(net713),
    .A2(net776),
    .Y(_0205_),
    .B1(_0684_));
 sg13g2_nor2_1 _2235_ (.A(\fifo_d[7][3] ),
    .B(net775),
    .Y(_0685_));
 sg13g2_a21oi_1 _2236_ (.A1(net710),
    .A2(net775),
    .Y(_0206_),
    .B1(_0685_));
 sg13g2_nor2_1 _2237_ (.A(\fifo_d[7][4] ),
    .B(net775),
    .Y(_0686_));
 sg13g2_a21oi_1 _2238_ (.A1(net708),
    .A2(net775),
    .Y(_0207_),
    .B1(_0686_));
 sg13g2_nor2_1 _2239_ (.A(\fifo_d[7][5] ),
    .B(net775),
    .Y(_0687_));
 sg13g2_a21oi_1 _2240_ (.A1(net706),
    .A2(net775),
    .Y(_0208_),
    .B1(_0687_));
 sg13g2_nor2_1 _2241_ (.A(\fifo_d[7][6] ),
    .B(net777),
    .Y(_0688_));
 sg13g2_a21oi_1 _2242_ (.A1(net703),
    .A2(net777),
    .Y(_0209_),
    .B1(_0688_));
 sg13g2_nor2_1 _2243_ (.A(\fifo_d[7][7] ),
    .B(net777),
    .Y(_0689_));
 sg13g2_a21oi_1 _2244_ (.A1(net701),
    .A2(net777),
    .Y(_0210_),
    .B1(_0689_));
 sg13g2_nor2b_2 _2245_ (.A(net821),
    .B_N(net820),
    .Y(_0690_));
 sg13g2_nand2_1 _2246_ (.Y(_0691_),
    .A(_0410_),
    .B(_0690_));
 sg13g2_nand2_1 _2247_ (.Y(_0692_),
    .A(\fifo_d[8][0] ),
    .B(net802));
 sg13g2_o21ai_1 _2248_ (.B1(_0692_),
    .Y(_0211_),
    .A1(net717),
    .A2(net801));
 sg13g2_nand2_1 _2249_ (.Y(_0693_),
    .A(\fifo_d[8][1] ),
    .B(net803));
 sg13g2_o21ai_1 _2250_ (.B1(_0693_),
    .Y(_0212_),
    .A1(net714),
    .A2(net803));
 sg13g2_nand2_1 _2251_ (.Y(_0694_),
    .A(\fifo_d[8][2] ),
    .B(net803));
 sg13g2_o21ai_1 _2252_ (.B1(_0694_),
    .Y(_0213_),
    .A1(net712),
    .A2(net803));
 sg13g2_nand2_1 _2253_ (.Y(_0695_),
    .A(\fifo_d[8][3] ),
    .B(net801));
 sg13g2_o21ai_1 _2254_ (.B1(_0695_),
    .Y(_0214_),
    .A1(_0526_),
    .A2(net801));
 sg13g2_nand2_1 _2255_ (.Y(_0696_),
    .A(\fifo_d[8][4] ),
    .B(net802));
 sg13g2_o21ai_1 _2256_ (.B1(_0696_),
    .Y(_0215_),
    .A1(net708),
    .A2(net802));
 sg13g2_nand2_1 _2257_ (.Y(_0697_),
    .A(\fifo_d[8][5] ),
    .B(net801));
 sg13g2_o21ai_1 _2258_ (.B1(_0697_),
    .Y(_0216_),
    .A1(net706),
    .A2(net801));
 sg13g2_nand2_1 _2259_ (.Y(_0698_),
    .A(\fifo_d[8][6] ),
    .B(net801));
 sg13g2_o21ai_1 _2260_ (.B1(_0698_),
    .Y(_0217_),
    .A1(net704),
    .A2(net801));
 sg13g2_nand2_1 _2261_ (.Y(_0699_),
    .A(\fifo_d[8][7] ),
    .B(net802));
 sg13g2_o21ai_1 _2262_ (.B1(_0699_),
    .Y(_0218_),
    .A1(net702),
    .A2(net801));
 sg13g2_nand2_1 _2263_ (.Y(_0700_),
    .A(_0411_),
    .B(_0690_));
 sg13g2_nand2_1 _2264_ (.Y(_0701_),
    .A(\fifo_d[9][0] ),
    .B(net800));
 sg13g2_o21ai_1 _2265_ (.B1(_0701_),
    .Y(_0219_),
    .A1(net716),
    .A2(net800));
 sg13g2_nand2_1 _2266_ (.Y(_0702_),
    .A(\fifo_d[9][1] ),
    .B(net799));
 sg13g2_o21ai_1 _2267_ (.B1(_0702_),
    .Y(_0220_),
    .A1(net715),
    .A2(net799));
 sg13g2_nand2_1 _2268_ (.Y(_0703_),
    .A(\fifo_d[9][2] ),
    .B(net800));
 sg13g2_o21ai_1 _2269_ (.B1(_0703_),
    .Y(_0221_),
    .A1(net712),
    .A2(net800));
 sg13g2_nand2_1 _2270_ (.Y(_0704_),
    .A(\fifo_d[9][3] ),
    .B(net798));
 sg13g2_o21ai_1 _2271_ (.B1(_0704_),
    .Y(_0222_),
    .A1(net710),
    .A2(net798));
 sg13g2_nand2_1 _2272_ (.Y(_0705_),
    .A(\fifo_d[9][4] ),
    .B(net798));
 sg13g2_o21ai_1 _2273_ (.B1(_0705_),
    .Y(_0223_),
    .A1(net708),
    .A2(net798));
 sg13g2_nand2_1 _2274_ (.Y(_0706_),
    .A(\fifo_d[9][5] ),
    .B(net798));
 sg13g2_o21ai_1 _2275_ (.B1(_0706_),
    .Y(_0224_),
    .A1(net706),
    .A2(net798));
 sg13g2_nand2_1 _2276_ (.Y(_0707_),
    .A(\fifo_d[9][6] ),
    .B(net799));
 sg13g2_o21ai_1 _2277_ (.B1(_0707_),
    .Y(_0225_),
    .A1(net703),
    .A2(net799));
 sg13g2_nand2_1 _2278_ (.Y(_0708_),
    .A(\fifo_d[9][7] ),
    .B(net798));
 sg13g2_o21ai_1 _2279_ (.B1(_0708_),
    .Y(_0226_),
    .A1(net702),
    .A2(net798));
 sg13g2_nand2_2 _2280_ (.Y(_0709_),
    .A(_0412_),
    .B(_0690_));
 sg13g2_nand2_1 _2281_ (.Y(_0710_),
    .A(\fifo_d[10][0] ),
    .B(net797));
 sg13g2_o21ai_1 _2282_ (.B1(_0710_),
    .Y(_0227_),
    .A1(net717),
    .A2(net797));
 sg13g2_nand2_1 _2283_ (.Y(_0711_),
    .A(\fifo_d[10][1] ),
    .B(net797));
 sg13g2_o21ai_1 _2284_ (.B1(_0711_),
    .Y(_0228_),
    .A1(net715),
    .A2(net797));
 sg13g2_nand2_1 _2285_ (.Y(_0712_),
    .A(\fifo_d[10][2] ),
    .B(net797));
 sg13g2_o21ai_1 _2286_ (.B1(_0712_),
    .Y(_0229_),
    .A1(net713),
    .A2(net797));
 sg13g2_nand2_1 _2287_ (.Y(_0713_),
    .A(\fifo_d[10][3] ),
    .B(net796));
 sg13g2_o21ai_1 _2288_ (.B1(_0713_),
    .Y(_0230_),
    .A1(net710),
    .A2(net796));
 sg13g2_nand2_1 _2289_ (.Y(_0714_),
    .A(\fifo_d[10][4] ),
    .B(net797));
 sg13g2_o21ai_1 _2290_ (.B1(_0714_),
    .Y(_0231_),
    .A1(net708),
    .A2(net797));
 sg13g2_nand2_1 _2291_ (.Y(_0715_),
    .A(\fifo_d[10][5] ),
    .B(net796));
 sg13g2_o21ai_1 _2292_ (.B1(_0715_),
    .Y(_0232_),
    .A1(net706),
    .A2(net796));
 sg13g2_nand2_1 _2293_ (.Y(_0716_),
    .A(\fifo_d[10][6] ),
    .B(net796));
 sg13g2_o21ai_1 _2294_ (.B1(_0716_),
    .Y(_0233_),
    .A1(net703),
    .A2(net796));
 sg13g2_nand2_1 _2295_ (.Y(_0717_),
    .A(\fifo_d[10][7] ),
    .B(net796));
 sg13g2_o21ai_1 _2296_ (.B1(_0717_),
    .Y(_0234_),
    .A1(net701),
    .A2(net796));
 sg13g2_nand2_1 _2297_ (.Y(_0718_),
    .A(_0409_),
    .B(_0690_));
 sg13g2_nand2_1 _2298_ (.Y(_0719_),
    .A(\fifo_d[11][0] ),
    .B(net795));
 sg13g2_o21ai_1 _2299_ (.B1(_0719_),
    .Y(_0235_),
    .A1(net717),
    .A2(net795));
 sg13g2_nand2_1 _2300_ (.Y(_0720_),
    .A(\fifo_d[11][1] ),
    .B(net795));
 sg13g2_o21ai_1 _2301_ (.B1(_0720_),
    .Y(_0236_),
    .A1(net715),
    .A2(net795));
 sg13g2_nand2_1 _2302_ (.Y(_0721_),
    .A(\fifo_d[11][2] ),
    .B(net795));
 sg13g2_o21ai_1 _2303_ (.B1(_0721_),
    .Y(_0237_),
    .A1(net713),
    .A2(net795));
 sg13g2_nand2_1 _2304_ (.Y(_0722_),
    .A(\fifo_d[11][3] ),
    .B(net794));
 sg13g2_o21ai_1 _2305_ (.B1(_0722_),
    .Y(_0238_),
    .A1(net710),
    .A2(net794));
 sg13g2_nand2_1 _2306_ (.Y(_0723_),
    .A(\fifo_d[11][4] ),
    .B(net794));
 sg13g2_o21ai_1 _2307_ (.B1(_0723_),
    .Y(_0239_),
    .A1(net708),
    .A2(net794));
 sg13g2_nand2_1 _2308_ (.Y(_0724_),
    .A(\fifo_d[11][5] ),
    .B(net794));
 sg13g2_o21ai_1 _2309_ (.B1(_0724_),
    .Y(_0240_),
    .A1(net707),
    .A2(net794));
 sg13g2_nand2_1 _2310_ (.Y(_0725_),
    .A(\fifo_d[11][6] ),
    .B(net794));
 sg13g2_o21ai_1 _2311_ (.B1(_0725_),
    .Y(_0241_),
    .A1(net703),
    .A2(net794));
 sg13g2_nand2_1 _2312_ (.Y(_0726_),
    .A(\fifo_d[11][7] ),
    .B(net795));
 sg13g2_o21ai_1 _2313_ (.B1(_0726_),
    .Y(_0242_),
    .A1(net702),
    .A2(net795));
 sg13g2_nand3_1 _2314_ (.B(net819),
    .C(_0410_),
    .A(net821),
    .Y(_0727_));
 sg13g2_nand2_1 _2315_ (.Y(_0728_),
    .A(\fifo_d[12][0] ),
    .B(net793));
 sg13g2_o21ai_1 _2316_ (.B1(_0728_),
    .Y(_0243_),
    .A1(net716),
    .A2(net793));
 sg13g2_nand2_1 _2317_ (.Y(_0729_),
    .A(\fifo_d[12][1] ),
    .B(net792));
 sg13g2_o21ai_1 _2318_ (.B1(_0729_),
    .Y(_0244_),
    .A1(net714),
    .A2(net792));
 sg13g2_nand2_1 _2319_ (.Y(_0730_),
    .A(\fifo_d[12][2] ),
    .B(net792));
 sg13g2_o21ai_1 _2320_ (.B1(_0730_),
    .Y(_0245_),
    .A1(net712),
    .A2(net792));
 sg13g2_nand2_1 _2321_ (.Y(_0731_),
    .A(\fifo_d[12][3] ),
    .B(net793));
 sg13g2_o21ai_1 _2322_ (.B1(_0731_),
    .Y(_0246_),
    .A1(net711),
    .A2(net793));
 sg13g2_nand2_1 _2323_ (.Y(_0732_),
    .A(\fifo_d[12][4] ),
    .B(net792));
 sg13g2_o21ai_1 _2324_ (.B1(_0732_),
    .Y(_0247_),
    .A1(net709),
    .A2(net792));
 sg13g2_nand2_1 _2325_ (.Y(_0733_),
    .A(\fifo_d[12][5] ),
    .B(net793));
 sg13g2_o21ai_1 _2326_ (.B1(_0733_),
    .Y(_0248_),
    .A1(net707),
    .A2(net793));
 sg13g2_nand2_1 _2327_ (.Y(_0734_),
    .A(\fifo_d[12][6] ),
    .B(_0727_));
 sg13g2_o21ai_1 _2328_ (.B1(_0734_),
    .Y(_0249_),
    .A1(net703),
    .A2(net793));
 sg13g2_nand2_1 _2329_ (.Y(_0735_),
    .A(\fifo_d[12][7] ),
    .B(net792));
 sg13g2_o21ai_1 _2330_ (.B1(_0735_),
    .Y(_0250_),
    .A1(net701),
    .A2(net792));
 sg13g2_and3_1 _2331_ (.X(_0736_),
    .A(net821),
    .B(net819),
    .C(_0411_));
 sg13g2_nor2_1 _2332_ (.A(\fifo_d[13][0] ),
    .B(net791),
    .Y(_0737_));
 sg13g2_a21oi_1 _2333_ (.A1(net716),
    .A2(net791),
    .Y(_0251_),
    .B1(_0737_));
 sg13g2_nor2_1 _2334_ (.A(\fifo_d[13][1] ),
    .B(net790),
    .Y(_0738_));
 sg13g2_a21oi_1 _2335_ (.A1(net714),
    .A2(net790),
    .Y(_0252_),
    .B1(_0738_));
 sg13g2_nor2_1 _2336_ (.A(\fifo_d[13][2] ),
    .B(net790),
    .Y(_0739_));
 sg13g2_a21oi_1 _2337_ (.A1(net712),
    .A2(net790),
    .Y(_0253_),
    .B1(_0739_));
 sg13g2_nor2_1 _2338_ (.A(\fifo_d[13][3] ),
    .B(net790),
    .Y(_0740_));
 sg13g2_a21oi_1 _2339_ (.A1(net711),
    .A2(net790),
    .Y(_0254_),
    .B1(_0740_));
 sg13g2_nor2_1 _2340_ (.A(\fifo_d[13][4] ),
    .B(net791),
    .Y(_0741_));
 sg13g2_a21oi_1 _2341_ (.A1(net709),
    .A2(net791),
    .Y(_0255_),
    .B1(_0741_));
 sg13g2_nor2_1 _2342_ (.A(\fifo_d[13][5] ),
    .B(net790),
    .Y(_0742_));
 sg13g2_a21oi_1 _2343_ (.A1(net707),
    .A2(net790),
    .Y(_0256_),
    .B1(_0742_));
 sg13g2_nor2_1 _2344_ (.A(\fifo_d[13][6] ),
    .B(_0736_),
    .Y(_0743_));
 sg13g2_a21oi_1 _2345_ (.A1(net703),
    .A2(net791),
    .Y(_0257_),
    .B1(_0743_));
 sg13g2_nor2_1 _2346_ (.A(\fifo_d[13][7] ),
    .B(net791),
    .Y(_0744_));
 sg13g2_a21oi_1 _2347_ (.A1(net701),
    .A2(net791),
    .Y(_0258_),
    .B1(_0744_));
 sg13g2_nand3_1 _2348_ (.B(net820),
    .C(_0412_),
    .A(net821),
    .Y(_0745_));
 sg13g2_nand2_1 _2349_ (.Y(_0746_),
    .A(\fifo_d[14][0] ),
    .B(net788));
 sg13g2_o21ai_1 _2350_ (.B1(_0746_),
    .Y(_0259_),
    .A1(net716),
    .A2(net788));
 sg13g2_nand2_1 _2351_ (.Y(_0747_),
    .A(\fifo_d[14][1] ),
    .B(net788));
 sg13g2_o21ai_1 _2352_ (.B1(_0747_),
    .Y(_0260_),
    .A1(net714),
    .A2(net788));
 sg13g2_nand2_1 _2353_ (.Y(_0748_),
    .A(\fifo_d[14][2] ),
    .B(net788));
 sg13g2_o21ai_1 _2354_ (.B1(_0748_),
    .Y(_0261_),
    .A1(net712),
    .A2(net788));
 sg13g2_nand2_1 _2355_ (.Y(_0749_),
    .A(\fifo_d[14][3] ),
    .B(_0745_));
 sg13g2_o21ai_1 _2356_ (.B1(_0749_),
    .Y(_0262_),
    .A1(net711),
    .A2(net789));
 sg13g2_nand2_1 _2357_ (.Y(_0750_),
    .A(\fifo_d[14][4] ),
    .B(net789));
 sg13g2_o21ai_1 _2358_ (.B1(_0750_),
    .Y(_0263_),
    .A1(net709),
    .A2(net789));
 sg13g2_nand2_1 _2359_ (.Y(_0751_),
    .A(\fifo_d[14][5] ),
    .B(net789));
 sg13g2_o21ai_1 _2360_ (.B1(_0751_),
    .Y(_0264_),
    .A1(net707),
    .A2(net789));
 sg13g2_nand2_1 _2361_ (.Y(_0752_),
    .A(\fifo_d[14][6] ),
    .B(net788));
 sg13g2_o21ai_1 _2362_ (.B1(_0752_),
    .Y(_0265_),
    .A1(net705),
    .A2(net788));
 sg13g2_nand2_1 _2363_ (.Y(_0753_),
    .A(\fifo_d[14][7] ),
    .B(net789));
 sg13g2_o21ai_1 _2364_ (.B1(_0753_),
    .Y(_0266_),
    .A1(net701),
    .A2(net789));
 sg13g2_nand2_1 _2365_ (.Y(_0754_),
    .A(net819),
    .B(_0415_));
 sg13g2_nand2_1 _2366_ (.Y(_0755_),
    .A(\fifo_d[15][0] ),
    .B(net751));
 sg13g2_o21ai_1 _2367_ (.B1(_0755_),
    .Y(_0267_),
    .A1(net717),
    .A2(net751));
 sg13g2_nand2_1 _2368_ (.Y(_0756_),
    .A(\fifo_d[15][1] ),
    .B(net753));
 sg13g2_o21ai_1 _2369_ (.B1(_0756_),
    .Y(_0268_),
    .A1(net714),
    .A2(net753));
 sg13g2_nand2_1 _2370_ (.Y(_0757_),
    .A(\fifo_d[15][2] ),
    .B(net751));
 sg13g2_o21ai_1 _2371_ (.B1(_0757_),
    .Y(_0269_),
    .A1(net713),
    .A2(net751));
 sg13g2_nand2_1 _2372_ (.Y(_0758_),
    .A(\fifo_d[15][3] ),
    .B(net751));
 sg13g2_o21ai_1 _2373_ (.B1(_0758_),
    .Y(_0270_),
    .A1(net710),
    .A2(net751));
 sg13g2_nand2_1 _2374_ (.Y(_0759_),
    .A(\fifo_d[15][4] ),
    .B(net752));
 sg13g2_o21ai_1 _2375_ (.B1(_0759_),
    .Y(_0271_),
    .A1(net708),
    .A2(net752));
 sg13g2_nand2_1 _2376_ (.Y(_0760_),
    .A(\fifo_d[15][5] ),
    .B(net751));
 sg13g2_o21ai_1 _2377_ (.B1(_0760_),
    .Y(_0272_),
    .A1(net706),
    .A2(net751));
 sg13g2_nand2_1 _2378_ (.Y(_0761_),
    .A(\fifo_d[15][6] ),
    .B(net753));
 sg13g2_o21ai_1 _2379_ (.B1(_0761_),
    .Y(_0273_),
    .A1(net703),
    .A2(net753));
 sg13g2_nand2_1 _2380_ (.Y(_0762_),
    .A(\fifo_d[15][7] ),
    .B(net752));
 sg13g2_o21ai_1 _2381_ (.B1(_0762_),
    .Y(_0274_),
    .A1(net702),
    .A2(net752));
 sg13g2_nor2_1 _2382_ (.A(\uart_0.rx.rx_sample_cnt[5] ),
    .B(\uart_0.rx.rx_sample_cnt[4] ),
    .Y(_0763_));
 sg13g2_nand2_1 _2383_ (.Y(_0764_),
    .A(_0034_),
    .B(_0763_));
 sg13g2_nor3_1 _2384_ (.A(\uart_0.rx.rx_sample_cnt[2] ),
    .B(\uart_0.rx.rx_sample_cnt[0] ),
    .C(\uart_0.rx.rx_sample_cnt[1] ),
    .Y(_0765_));
 sg13g2_nor2b_1 _2385_ (.A(_0765_),
    .B_N(\uart_0.rx.rx_sample_cnt[3] ),
    .Y(_0766_));
 sg13g2_nor3_1 _2386_ (.A(_1388_),
    .B(_0764_),
    .C(_0766_),
    .Y(_0767_));
 sg13g2_nor2_2 _2387_ (.A(net784),
    .B(_0767_),
    .Y(_0768_));
 sg13g2_nand2_1 _2388_ (.Y(_0769_),
    .A(_0041_),
    .B(_0768_));
 sg13g2_nand3_1 _2389_ (.B(\uart_0.rx.rx_sample_cnt[0] ),
    .C(\uart_0.rx.rx_sample_cnt[1] ),
    .A(\uart_0.rx.rx_sample_cnt[2] ),
    .Y(_0770_));
 sg13g2_nand3b_1 _2390_ (.B(net816),
    .C(_0767_),
    .Y(_0771_),
    .A_N(\uart_0.rx.rx_sample_cnt[3] ));
 sg13g2_or2_1 _2391_ (.X(_0772_),
    .B(_0771_),
    .A(_0770_));
 sg13g2_nand2_1 _2392_ (.Y(_0275_),
    .A(_0769_),
    .B(_0772_));
 sg13g2_nand2_1 _2393_ (.Y(_0773_),
    .A(\uart_0.rx.rx_sample_wrap[3] ),
    .B(_0768_));
 sg13g2_nand2_1 _2394_ (.Y(_0276_),
    .A(_0772_),
    .B(_0773_));
 sg13g2_nand2_1 _2395_ (.Y(_0774_),
    .A(_1232_),
    .B(_1234_));
 sg13g2_and2_1 _2396_ (.A(tx_do),
    .B(tx_data_done),
    .X(_0775_));
 sg13g2_nand3b_1 _2397_ (.B(_0774_),
    .C(net818),
    .Y(_0776_),
    .A_N(_1357_));
 sg13g2_inv_1 _2398_ (.Y(_0777_),
    .A(_0776_));
 sg13g2_a221oi_1 _2399_ (.B2(_0037_),
    .C1(net774),
    .B1(_0777_),
    .A1(\uart_0.tx.tx_bit_cnt[0] ),
    .Y(_0778_),
    .A2(_1357_));
 sg13g2_inv_1 _2400_ (.Y(_0277_),
    .A(_0778_));
 sg13g2_nand4_1 _2401_ (.B(_1235_),
    .C(_1358_),
    .A(_1222_),
    .Y(_0779_),
    .D(_0774_));
 sg13g2_o21ai_1 _2402_ (.B1(_0779_),
    .Y(_0278_),
    .A1(_1137_),
    .A2(_1358_));
 sg13g2_nand2_1 _2403_ (.Y(_0780_),
    .A(\uart_0.tx.tx_bit_cnt[2] ),
    .B(_1357_));
 sg13g2_nor2_1 _2404_ (.A(_0036_),
    .B(_1235_),
    .Y(_0781_));
 sg13g2_xnor2_1 _2405_ (.Y(_0782_),
    .A(_0036_),
    .B(_1235_));
 sg13g2_o21ai_1 _2406_ (.B1(_0780_),
    .Y(_0279_),
    .A1(_0776_),
    .A2(_0782_));
 sg13g2_nand2_1 _2407_ (.Y(_0783_),
    .A(\uart_0.tx.tx_bit_cnt[3] ),
    .B(_1357_));
 sg13g2_xor2_1 _2408_ (.B(_0781_),
    .A(_0035_),
    .X(_0784_));
 sg13g2_o21ai_1 _2409_ (.B1(_0783_),
    .Y(_0280_),
    .A1(_0776_),
    .A2(_0784_));
 sg13g2_nand2_1 _2410_ (.Y(_0785_),
    .A(_1220_),
    .B(_1390_));
 sg13g2_inv_4 _2411_ (.A(net738),
    .Y(_0786_));
 sg13g2_nor3_1 _2412_ (.A(\uart_0.rx.rx_marker[3] ),
    .B(net848),
    .C(_1374_),
    .Y(_0787_));
 sg13g2_o21ai_1 _2413_ (.B1(_0033_),
    .Y(_0788_),
    .A1(_1215_),
    .A2(_0787_));
 sg13g2_nor3_1 _2414_ (.A(\uart_0.rx.rx_marker[3] ),
    .B(_1216_),
    .C(_1375_),
    .Y(_0789_));
 sg13g2_nor3_1 _2415_ (.A(_1134_),
    .B(\uart_0.rx.rx_data_in ),
    .C(_0789_),
    .Y(_0790_));
 sg13g2_and2_1 _2416_ (.A(_0788_),
    .B(_0790_),
    .X(_0791_));
 sg13g2_nor2_1 _2417_ (.A(\uart_0.rx.rx_marker[0] ),
    .B(\uart_0.rx.rx_marker[1] ),
    .Y(_0792_));
 sg13g2_or2_1 _2418_ (.X(_0793_),
    .B(\uart_0.rx.rx_marker[1] ),
    .A(\uart_0.rx.rx_marker[0] ));
 sg13g2_nand3_1 _2419_ (.B(\uart_0.rx.rx_marker[6] ),
    .C(_0792_),
    .A(net848),
    .Y(_0794_));
 sg13g2_nor3_1 _2420_ (.A(\uart_0.rx.rx_marker[3] ),
    .B(_1215_),
    .C(_0794_),
    .Y(_0795_));
 sg13g2_nor2_1 _2421_ (.A(\uart_0.rx.rx_samples[0] ),
    .B(_0795_),
    .Y(_0796_));
 sg13g2_a21oi_1 _2422_ (.A1(net852),
    .A2(_0796_),
    .Y(_0797_),
    .B1(net783));
 sg13g2_a21oi_1 _2423_ (.A1(_0791_),
    .A2(_0797_),
    .Y(_0798_),
    .B1(net749));
 sg13g2_a21oi_1 _2424_ (.A1(_1165_),
    .A2(net749),
    .Y(_0281_),
    .B1(_0798_));
 sg13g2_nand2_1 _2425_ (.Y(_0799_),
    .A(\uart_0.rx.rx_stop_zeros[1] ),
    .B(net747));
 sg13g2_and2_2 _2426_ (.A(net851),
    .B(\uart_0.rx.rx_stop_zeros[1] ),
    .X(_0800_));
 sg13g2_nand2_2 _2427_ (.Y(_0801_),
    .A(net851),
    .B(\uart_0.rx.rx_stop_zeros[1] ));
 sg13g2_xnor2_1 _2428_ (.Y(_0802_),
    .A(net851),
    .B(\uart_0.rx.rx_stop_zeros[1] ));
 sg13g2_nor2_1 _2429_ (.A(\uart_0.rx.rx_data_in ),
    .B(net816),
    .Y(_0803_));
 sg13g2_or2_2 _2430_ (.X(_0804_),
    .B(net816),
    .A(\uart_0.rx.rx_data_in ));
 sg13g2_nand4_1 _2431_ (.B(_0791_),
    .C(_0796_),
    .A(_0786_),
    .Y(_0805_),
    .D(net770));
 sg13g2_o21ai_1 _2432_ (.B1(_0799_),
    .Y(_0282_),
    .A1(_0802_),
    .A2(_0805_));
 sg13g2_nand2_1 _2433_ (.Y(_0806_),
    .A(\uart_0.rx.rx_stop_zeros[2] ),
    .B(net747));
 sg13g2_nor2_2 _2434_ (.A(_0028_),
    .B(_0801_),
    .Y(_0807_));
 sg13g2_xnor2_1 _2435_ (.Y(_0808_),
    .A(_0028_),
    .B(_0800_));
 sg13g2_xnor2_1 _2436_ (.Y(_0809_),
    .A(_1166_),
    .B(_0800_));
 sg13g2_o21ai_1 _2437_ (.B1(_0806_),
    .Y(_0283_),
    .A1(_0805_),
    .A2(_0809_));
 sg13g2_nand2_1 _2438_ (.Y(_0810_),
    .A(net850),
    .B(net747));
 sg13g2_nor2b_2 _2439_ (.A(_0807_),
    .B_N(net849),
    .Y(_0811_));
 sg13g2_inv_1 _2440_ (.Y(_0812_),
    .A(_0811_));
 sg13g2_nor3_2 _2441_ (.A(_0028_),
    .B(net849),
    .C(_0801_),
    .Y(_0813_));
 sg13g2_nor2_2 _2442_ (.A(_0811_),
    .B(_0813_),
    .Y(_0814_));
 sg13g2_or2_1 _2443_ (.X(_0815_),
    .B(_0813_),
    .A(_0811_));
 sg13g2_o21ai_1 _2444_ (.B1(_0810_),
    .Y(_0284_),
    .A1(_0805_),
    .A2(_0814_));
 sg13g2_nand2_1 _2445_ (.Y(_0816_),
    .A(\uart_0.rx.rx_stop_zeros[4] ),
    .B(net749));
 sg13g2_nand3_1 _2446_ (.B(net850),
    .C(_0800_),
    .A(\uart_0.rx.rx_stop_zeros[2] ),
    .Y(_0817_));
 sg13g2_nor2_1 _2447_ (.A(_0030_),
    .B(_0817_),
    .Y(_0818_));
 sg13g2_xor2_1 _2448_ (.B(_0817_),
    .A(_0030_),
    .X(_0819_));
 sg13g2_xnor2_1 _2449_ (.Y(_0820_),
    .A(_0030_),
    .B(_0817_));
 sg13g2_o21ai_1 _2450_ (.B1(_0816_),
    .Y(_0285_),
    .A1(_0805_),
    .A2(_0820_));
 sg13g2_xnor2_1 _2451_ (.Y(_0821_),
    .A(_0029_),
    .B(_0818_));
 sg13g2_nor2b_1 _2452_ (.A(_0805_),
    .B_N(_0821_),
    .Y(_0822_));
 sg13g2_a21o_1 _2453_ (.A2(net747),
    .A1(\uart_0.rx.rx_stop_zeros[5] ),
    .B1(_0822_),
    .X(_0286_));
 sg13g2_nand2_1 _2454_ (.Y(_0823_),
    .A(\uart_0.rx.rx_stop_zeros[6] ),
    .B(net749));
 sg13g2_nand2_1 _2455_ (.Y(_0824_),
    .A(\uart_0.rx.rx_stop_zeros[4] ),
    .B(\uart_0.rx.rx_stop_zeros[5] ));
 sg13g2_o21ai_1 _2456_ (.B1(_0031_),
    .Y(_0825_),
    .A1(_0817_),
    .A2(_0824_));
 sg13g2_nor3_2 _2457_ (.A(_0031_),
    .B(_0817_),
    .C(_0824_),
    .Y(_0826_));
 sg13g2_inv_1 _2458_ (.Y(_0827_),
    .A(_0826_));
 sg13g2_nand2_2 _2459_ (.Y(_0828_),
    .A(_0825_),
    .B(_0827_));
 sg13g2_o21ai_1 _2460_ (.B1(_0823_),
    .Y(_0287_),
    .A1(_0805_),
    .A2(_0828_));
 sg13g2_a22oi_1 _2461_ (.Y(_0829_),
    .B1(net773),
    .B2(net852),
    .A2(net815),
    .A1(_1133_));
 sg13g2_xnor2_1 _2462_ (.Y(_0288_),
    .A(net782),
    .B(_0829_));
 sg13g2_o21ai_1 _2463_ (.B1(_1373_),
    .Y(_0830_),
    .A1(_1216_),
    .A2(_0793_));
 sg13g2_o21ai_1 _2464_ (.B1(_0830_),
    .Y(_0831_),
    .A1(_1374_),
    .A2(_0792_));
 sg13g2_nor2_1 _2465_ (.A(\uart_0.rx.rx_stop_zeros[1] ),
    .B(net770),
    .Y(_0832_));
 sg13g2_a21oi_1 _2466_ (.A1(_0042_),
    .A2(net782),
    .Y(_0833_),
    .B1(_0832_));
 sg13g2_o21ai_1 _2467_ (.B1(_0833_),
    .Y(_0289_),
    .A1(net782),
    .A2(_0831_));
 sg13g2_or2_1 _2468_ (.X(_0834_),
    .B(_1388_),
    .A(net784));
 sg13g2_xnor2_1 _2469_ (.Y(_0835_),
    .A(\uart_0.rx.rx_marker[2] ),
    .B(_1374_));
 sg13g2_a22oi_1 _2470_ (.Y(_0836_),
    .B1(net773),
    .B2(_1166_),
    .A2(net782),
    .A1(\uart_0.rx.rx_marker[2] ));
 sg13g2_o21ai_1 _2471_ (.B1(_0836_),
    .Y(_0290_),
    .A1(_0834_),
    .A2(_0835_));
 sg13g2_nand3_1 _2472_ (.B(net848),
    .C(_1374_),
    .A(\uart_0.rx.rx_marker[3] ),
    .Y(_0837_));
 sg13g2_a21o_1 _2473_ (.A2(_1374_),
    .A1(net848),
    .B1(\uart_0.rx.rx_marker[3] ),
    .X(_0838_));
 sg13g2_nand2_1 _2474_ (.Y(_0839_),
    .A(_0837_),
    .B(_0838_));
 sg13g2_a21oi_1 _2475_ (.A1(_0830_),
    .A2(_0839_),
    .Y(_0840_),
    .B1(_1389_));
 sg13g2_o21ai_1 _2476_ (.B1(_0840_),
    .Y(_0841_),
    .A1(net850),
    .A2(net770));
 sg13g2_o21ai_1 _2477_ (.B1(_0841_),
    .Y(_0842_),
    .A1(_0043_),
    .A2(_1390_));
 sg13g2_inv_1 _2478_ (.Y(_0291_),
    .A(_0842_));
 sg13g2_nand4_1 _2479_ (.B(net848),
    .C(\uart_0.rx.rx_marker[4] ),
    .A(\uart_0.rx.rx_marker[3] ),
    .Y(_0843_),
    .D(_1374_));
 sg13g2_xor2_1 _2480_ (.B(_0837_),
    .A(\uart_0.rx.rx_marker[4] ),
    .X(_0844_));
 sg13g2_a21oi_1 _2481_ (.A1(_0830_),
    .A2(_0844_),
    .Y(_0845_),
    .B1(net782));
 sg13g2_o21ai_1 _2482_ (.B1(_0845_),
    .Y(_0846_),
    .A1(\uart_0.rx.rx_stop_zeros[4] ),
    .A2(net769));
 sg13g2_o21ai_1 _2483_ (.B1(_0846_),
    .Y(_0847_),
    .A1(_0044_),
    .A2(_1390_));
 sg13g2_inv_1 _2484_ (.Y(_0292_),
    .A(_0847_));
 sg13g2_xor2_1 _2485_ (.B(_0843_),
    .A(_0033_),
    .X(_0848_));
 sg13g2_a221oi_1 _2486_ (.B2(_0848_),
    .C1(net782),
    .B1(_0830_),
    .A1(_1167_),
    .Y(_0849_),
    .A2(net773));
 sg13g2_a21oi_1 _2487_ (.A1(_1135_),
    .A2(_1389_),
    .Y(_0293_),
    .B1(_0849_));
 sg13g2_o21ai_1 _2488_ (.B1(_1134_),
    .Y(_0850_),
    .A1(_1135_),
    .A2(_0843_));
 sg13g2_a22oi_1 _2489_ (.Y(_0851_),
    .B1(net773),
    .B2(_1168_),
    .A2(net782),
    .A1(_0045_));
 sg13g2_o21ai_1 _2490_ (.B1(_0851_),
    .Y(_0294_),
    .A1(net782),
    .A2(_0850_));
 sg13g2_a22oi_1 _2491_ (.Y(_0852_),
    .B1(net774),
    .B2(\tx_data[0] ),
    .A2(net818),
    .A1(\uart_0.tx.tx_data_tmp[2] ));
 sg13g2_inv_1 _2492_ (.Y(_0295_),
    .A(_0852_));
 sg13g2_a22oi_1 _2493_ (.Y(_0853_),
    .B1(_0775_),
    .B2(\tx_data[1] ),
    .A2(_1223_),
    .A1(\uart_0.tx.tx_data_tmp[3] ));
 sg13g2_inv_1 _2494_ (.Y(_0296_),
    .A(_0853_));
 sg13g2_a22oi_1 _2495_ (.Y(_0854_),
    .B1(net774),
    .B2(\tx_data[2] ),
    .A2(_1223_),
    .A1(\uart_0.tx.tx_data_tmp[4] ));
 sg13g2_inv_1 _2496_ (.Y(_0297_),
    .A(_0854_));
 sg13g2_a22oi_1 _2497_ (.Y(_0855_),
    .B1(net774),
    .B2(\tx_data[3] ),
    .A2(net818),
    .A1(\uart_0.tx.tx_data_tmp[5] ));
 sg13g2_inv_1 _2498_ (.Y(_0298_),
    .A(_0855_));
 sg13g2_a22oi_1 _2499_ (.Y(_0856_),
    .B1(net774),
    .B2(\tx_data[4] ),
    .A2(net818),
    .A1(\uart_0.tx.tx_data_tmp[6] ));
 sg13g2_inv_1 _2500_ (.Y(_0299_),
    .A(_0856_));
 sg13g2_a22oi_1 _2501_ (.Y(_0857_),
    .B1(net774),
    .B2(\tx_data[5] ),
    .A2(net818),
    .A1(\uart_0.tx.tx_data_tmp[7] ));
 sg13g2_inv_1 _2502_ (.Y(_0300_),
    .A(_0857_));
 sg13g2_a22oi_1 _2503_ (.Y(_0858_),
    .B1(net774),
    .B2(\tx_data[6] ),
    .A2(net818),
    .A1(\uart_0.tx.tx_data_tmp[8] ));
 sg13g2_inv_1 _2504_ (.Y(_0301_),
    .A(_0858_));
 sg13g2_a22oi_1 _2505_ (.Y(_0859_),
    .B1(net774),
    .B2(\tx_data[7] ),
    .A2(net818),
    .A1(\uart_0.tx.tx_data_tmp[9] ));
 sg13g2_inv_1 _2506_ (.Y(_0302_),
    .A(_0859_));
 sg13g2_nor2_2 _2507_ (.A(net760),
    .B(net785),
    .Y(_0860_));
 sg13g2_or2_2 _2508_ (.X(_0861_),
    .B(net785),
    .A(net765));
 sg13g2_nor2_2 _2509_ (.A(net787),
    .B(net755),
    .Y(_0862_));
 sg13g2_inv_1 _2510_ (.Y(_0863_),
    .A(_0862_));
 sg13g2_nor2_2 _2511_ (.A(net755),
    .B(net785),
    .Y(_0864_));
 sg13g2_inv_1 _2512_ (.Y(_0865_),
    .A(_0864_));
 sg13g2_nor2_2 _2513_ (.A(net755),
    .B(net732),
    .Y(_0866_));
 sg13g2_nor2_2 _2514_ (.A(_0861_),
    .B(_0863_),
    .Y(_0867_));
 sg13g2_and2_2 _2515_ (.A(net849),
    .B(_0807_),
    .X(_0868_));
 sg13g2_nand2_2 _2516_ (.Y(_0869_),
    .A(net849),
    .B(_0807_));
 sg13g2_a21oi_1 _2517_ (.A1(net726),
    .A2(_0868_),
    .Y(_0870_),
    .B1(\uart_0.rx.rx_data_in ));
 sg13g2_mux2_1 _2518_ (.A0(_0046_),
    .A1(_0870_),
    .S(_0786_),
    .X(_0303_));
 sg13g2_a21oi_2 _2519_ (.B1(net748),
    .Y(_0871_),
    .A2(net783),
    .A1(\uart_0.rx.rx_data_in ));
 sg13g2_a21o_1 _2520_ (.A2(net783),
    .A1(\uart_0.rx.rx_data_in ),
    .B1(net740),
    .X(_0872_));
 sg13g2_nand2b_1 _2521_ (.Y(_0873_),
    .B(_0871_),
    .A_N(_0866_));
 sg13g2_nand2b_1 _2522_ (.Y(_0874_),
    .B(\uart_0.rx.rx_stop_zeros[1] ),
    .A_N(net851));
 sg13g2_nand2_2 _2523_ (.Y(_0875_),
    .A(_0809_),
    .B(_0874_));
 sg13g2_and2_1 _2524_ (.A(_0802_),
    .B(_0809_),
    .X(_0876_));
 sg13g2_nand2_2 _2525_ (.Y(_0877_),
    .A(_0802_),
    .B(_0809_));
 sg13g2_nor2_2 _2526_ (.A(net757),
    .B(net786),
    .Y(_0878_));
 sg13g2_nand2_1 _2527_ (.Y(_0879_),
    .A(_0876_),
    .B(_0878_));
 sg13g2_inv_1 _2528_ (.Y(_0880_),
    .A(_0879_));
 sg13g2_a221oi_1 _2529_ (.B2(_0880_),
    .C1(net728),
    .B1(_0866_),
    .A1(\uart_0.rx.rx_samples[0] ),
    .Y(_0881_),
    .A2(net764));
 sg13g2_a21o_1 _2530_ (.A2(net740),
    .A1(_0047_),
    .B1(_0881_),
    .X(_0304_));
 sg13g2_o21ai_1 _2531_ (.B1(_0871_),
    .Y(_0882_),
    .A1(net732),
    .A2(_0863_));
 sg13g2_nor2_2 _2532_ (.A(_0808_),
    .B(net757),
    .Y(_0883_));
 sg13g2_nand2_2 _2533_ (.Y(_0884_),
    .A(_0809_),
    .B(_0814_));
 sg13g2_nor3_2 _2534_ (.A(net756),
    .B(net732),
    .C(_0875_),
    .Y(_0885_));
 sg13g2_a221oi_1 _2535_ (.B2(_0885_),
    .C1(net729),
    .B1(_0862_),
    .A1(\uart_0.rx.rx_samples[1] ),
    .Y(_0886_),
    .A2(net764));
 sg13g2_a21o_1 _2536_ (.A2(net741),
    .A1(_0048_),
    .B1(_0886_),
    .X(_0305_));
 sg13g2_a221oi_1 _2537_ (.B2(_0883_),
    .C1(net729),
    .B1(_0867_),
    .A1(\uart_0.rx.rx_samples[2] ),
    .Y(_0887_),
    .A2(net764));
 sg13g2_a21o_1 _2538_ (.A2(net741),
    .A1(_0049_),
    .B1(_0887_),
    .X(_0306_));
 sg13g2_nor2_1 _2539_ (.A(net849),
    .B(_0809_),
    .Y(_0888_));
 sg13g2_nor3_2 _2540_ (.A(_1166_),
    .B(net849),
    .C(_0801_),
    .Y(_0889_));
 sg13g2_nor2_2 _2541_ (.A(_0883_),
    .B(_0889_),
    .Y(_0890_));
 sg13g2_or2_2 _2542_ (.X(_0891_),
    .B(_0889_),
    .A(_0883_));
 sg13g2_a221oi_1 _2543_ (.B2(_0891_),
    .C1(net729),
    .B1(net726),
    .A1(\uart_0.rx.rx_samples[3] ),
    .Y(_0892_),
    .A2(net764));
 sg13g2_a21o_1 _2544_ (.A2(net740),
    .A1(_0050_),
    .B1(_0892_),
    .X(_0307_));
 sg13g2_nor2_2 _2545_ (.A(_0028_),
    .B(_0802_),
    .Y(_0893_));
 sg13g2_nand2b_2 _2546_ (.Y(_0894_),
    .B(_1166_),
    .A_N(_0802_));
 sg13g2_nand3_1 _2547_ (.B(net726),
    .C(_0894_),
    .A(_0814_),
    .Y(_0895_));
 sg13g2_a21oi_1 _2548_ (.A1(\uart_0.rx.rx_samples[4] ),
    .A2(net765),
    .Y(_0896_),
    .B1(net729));
 sg13g2_a22oi_1 _2549_ (.Y(_0897_),
    .B1(_0895_),
    .B2(_0896_),
    .A2(net740),
    .A1(_0051_));
 sg13g2_inv_1 _2550_ (.Y(_0308_),
    .A(_0897_));
 sg13g2_nor2_2 _2551_ (.A(_0028_),
    .B(_0874_),
    .Y(_0898_));
 sg13g2_nor2_2 _2552_ (.A(net756),
    .B(_0898_),
    .Y(_0899_));
 sg13g2_nor3_2 _2553_ (.A(net763),
    .B(net756),
    .C(_0898_),
    .Y(_0900_));
 sg13g2_nand2_1 _2554_ (.Y(_0901_),
    .A(_0860_),
    .B(_0899_));
 sg13g2_a221oi_1 _2555_ (.B2(_0899_),
    .C1(net727),
    .B1(_0867_),
    .A1(\uart_0.rx.rx_samples[5] ),
    .Y(_0902_),
    .A2(net764));
 sg13g2_a21o_1 _2556_ (.A2(net739),
    .A1(_0052_),
    .B1(_0902_),
    .X(_0309_));
 sg13g2_a221oi_1 _2557_ (.B2(net726),
    .C1(net727),
    .B1(_0814_),
    .A1(\uart_0.rx.rx_samples[6] ),
    .Y(_0903_),
    .A2(net764));
 sg13g2_a21o_1 _2558_ (.A2(net739),
    .A1(_0053_),
    .B1(_0903_),
    .X(_0310_));
 sg13g2_a221oi_1 _2559_ (.B2(net726),
    .C1(net727),
    .B1(_0812_),
    .A1(\uart_0.rx.rx_samples[7] ),
    .Y(_0904_),
    .A2(net766));
 sg13g2_a21o_1 _2560_ (.A2(net739),
    .A1(_0054_),
    .B1(_0904_),
    .X(_0311_));
 sg13g2_a21oi_2 _2561_ (.B1(net786),
    .Y(_0905_),
    .A2(_0877_),
    .A1(net757));
 sg13g2_a221oi_1 _2562_ (.B2(_0905_),
    .C1(net730),
    .B1(_0866_),
    .A1(\uart_0.rx.rx_samples[8] ),
    .Y(_0906_),
    .A2(net762));
 sg13g2_a21o_1 _2563_ (.A2(net738),
    .A1(_0055_),
    .B1(_0906_),
    .X(_0312_));
 sg13g2_a21oi_2 _2564_ (.B1(net732),
    .Y(_0907_),
    .A2(_0875_),
    .A1(net756));
 sg13g2_a221oi_1 _2565_ (.B2(_0907_),
    .C1(net727),
    .B1(_0862_),
    .A1(\uart_0.rx.rx_samples[9] ),
    .Y(_0908_),
    .A2(net762));
 sg13g2_a21o_1 _2566_ (.A2(net738),
    .A1(_0056_),
    .B1(_0908_),
    .X(_0313_));
 sg13g2_and2_2 _2567_ (.A(net850),
    .B(_0808_),
    .X(_0909_));
 sg13g2_nand2_2 _2568_ (.Y(_0910_),
    .A(net849),
    .B(_0808_));
 sg13g2_a221oi_1 _2569_ (.B2(_0910_),
    .C1(net727),
    .B1(net726),
    .A1(\uart_0.rx.rx_samples[10] ),
    .Y(_0911_),
    .A2(net766));
 sg13g2_a21o_1 _2570_ (.A2(net742),
    .A1(_0057_),
    .B1(_0911_),
    .X(_0314_));
 sg13g2_nand2_2 _2571_ (.Y(_0912_),
    .A(_0801_),
    .B(_0909_));
 sg13g2_a221oi_1 _2572_ (.B2(_0912_),
    .C1(net730),
    .B1(net726),
    .A1(\uart_0.rx.rx_samples[11] ),
    .Y(_0913_),
    .A2(net762));
 sg13g2_a21o_1 _2573_ (.A2(net738),
    .A1(_0058_),
    .B1(_0913_),
    .X(_0315_));
 sg13g2_a21oi_2 _2574_ (.B1(net787),
    .Y(_0914_),
    .A2(_0893_),
    .A1(net757));
 sg13g2_a221oi_1 _2575_ (.B2(_0914_),
    .C1(net727),
    .B1(_0866_),
    .A1(\uart_0.rx.rx_samples[12] ),
    .Y(_0915_),
    .A2(net762));
 sg13g2_a21o_1 _2576_ (.A2(net738),
    .A1(_0059_),
    .B1(_0915_),
    .X(_0316_));
 sg13g2_nand2_2 _2577_ (.Y(_0916_),
    .A(net849),
    .B(_0898_));
 sg13g2_a221oi_1 _2578_ (.B2(_0916_),
    .C1(net727),
    .B1(net726),
    .A1(\uart_0.rx.rx_samples[13] ),
    .Y(_0917_),
    .A2(net766));
 sg13g2_a21o_1 _2579_ (.A2(net739),
    .A1(_0060_),
    .B1(_0917_),
    .X(_0317_));
 sg13g2_a21oi_1 _2580_ (.A1(\uart_0.rx.rx_samples[14] ),
    .A2(net762),
    .Y(_0918_),
    .B1(_0882_));
 sg13g2_a21o_1 _2581_ (.A2(net739),
    .A1(_0061_),
    .B1(_0918_),
    .X(_0318_));
 sg13g2_nand2_2 _2582_ (.Y(_0919_),
    .A(_0029_),
    .B(net787));
 sg13g2_nor2_1 _2583_ (.A(net785),
    .B(_0919_),
    .Y(_0920_));
 sg13g2_nor2_2 _2584_ (.A(_0861_),
    .B(_0919_),
    .Y(_0921_));
 sg13g2_a221oi_1 _2585_ (.B2(_0921_),
    .C1(_0882_),
    .B1(_0868_),
    .A1(\uart_0.rx.rx_samples[15] ),
    .Y(_0922_),
    .A2(net762));
 sg13g2_a21o_1 _2586_ (.A2(net739),
    .A1(_0062_),
    .B1(_0922_),
    .X(_0319_));
 sg13g2_nand2_2 _2587_ (.Y(_0923_),
    .A(_0814_),
    .B(net786));
 sg13g2_nor2_1 _2588_ (.A(_0877_),
    .B(_0923_),
    .Y(_0924_));
 sg13g2_o21ai_1 _2589_ (.B1(net786),
    .Y(_0925_),
    .A1(net757),
    .A2(_0877_));
 sg13g2_a21oi_1 _2590_ (.A1(_0864_),
    .A2(_0925_),
    .Y(_0926_),
    .B1(net763));
 sg13g2_nor2_1 _2591_ (.A(\uart_0.rx.rx_samples[16] ),
    .B(net783),
    .Y(_0927_));
 sg13g2_nor3_1 _2592_ (.A(net740),
    .B(_0926_),
    .C(_0927_),
    .Y(_0928_));
 sg13g2_a21oi_1 _2593_ (.A1(_1127_),
    .A2(net741),
    .Y(_0320_),
    .B1(_0928_));
 sg13g2_nand2_1 _2594_ (.Y(_0929_),
    .A(net852),
    .B(_0832_));
 sg13g2_nor2_2 _2595_ (.A(_0884_),
    .B(_0929_),
    .Y(_0930_));
 sg13g2_nand2_1 _2596_ (.Y(_0931_),
    .A(_0920_),
    .B(_0930_));
 sg13g2_a221oi_1 _2597_ (.B2(_0925_),
    .C1(net729),
    .B1(_0866_),
    .A1(\uart_0.rx.rx_samples[17] ),
    .Y(_0932_),
    .A2(net763));
 sg13g2_a22oi_1 _2598_ (.Y(_0933_),
    .B1(_0931_),
    .B2(_0932_),
    .A2(net740),
    .A1(_0064_));
 sg13g2_inv_1 _2599_ (.Y(_0321_),
    .A(_0933_));
 sg13g2_nor2_2 _2600_ (.A(_0860_),
    .B(net728),
    .Y(_0934_));
 sg13g2_nand2_2 _2601_ (.Y(_0935_),
    .A(_0861_),
    .B(_0871_));
 sg13g2_o21ai_1 _2602_ (.B1(_0863_),
    .Y(_0936_),
    .A1(_0884_),
    .A2(_0919_));
 sg13g2_o21ai_1 _2603_ (.B1(net724),
    .Y(_0937_),
    .A1(net728),
    .A2(_0936_));
 sg13g2_a221oi_1 _2604_ (.B2(_0936_),
    .C1(net728),
    .B1(_0860_),
    .A1(\uart_0.rx.rx_samples[18] ),
    .Y(_0938_),
    .A2(net769));
 sg13g2_a21o_1 _2605_ (.A2(net747),
    .A1(_0065_),
    .B1(_0938_),
    .X(_0322_));
 sg13g2_a22oi_1 _2606_ (.Y(_0939_),
    .B1(_0889_),
    .B2(_0921_),
    .A2(net769),
    .A1(\uart_0.rx.rx_samples[19] ));
 sg13g2_a22oi_1 _2607_ (.Y(_0940_),
    .B1(_0937_),
    .B2(_0939_),
    .A2(net747),
    .A1(_0066_));
 sg13g2_inv_1 _2608_ (.Y(_0323_),
    .A(_0940_));
 sg13g2_nand2_1 _2609_ (.Y(_0941_),
    .A(net786),
    .B(_0893_));
 sg13g2_nor2_2 _2610_ (.A(_0814_),
    .B(_0820_),
    .Y(_0942_));
 sg13g2_nor3_1 _2611_ (.A(net755),
    .B(net732),
    .C(_0942_),
    .Y(_0943_));
 sg13g2_a221oi_1 _2612_ (.B2(_0943_),
    .C1(net729),
    .B1(_0941_),
    .A1(\uart_0.rx.rx_samples[20] ),
    .Y(_0944_),
    .A2(net769));
 sg13g2_a21o_1 _2613_ (.A2(net748),
    .A1(_0067_),
    .B1(_0944_),
    .X(_0324_));
 sg13g2_a221oi_1 _2614_ (.B2(_0920_),
    .C1(_0882_),
    .B1(_0900_),
    .A1(\uart_0.rx.rx_samples[21] ),
    .Y(_0945_),
    .A2(net764));
 sg13g2_a21o_1 _2615_ (.A2(net748),
    .A1(_0068_),
    .B1(_0945_),
    .X(_0325_));
 sg13g2_o21ai_1 _2616_ (.B1(net772),
    .Y(_0946_),
    .A1(_0865_),
    .A2(_0942_));
 sg13g2_o21ai_1 _2617_ (.B1(_0946_),
    .Y(_0947_),
    .A1(\uart_0.rx.rx_samples[22] ),
    .A2(net783));
 sg13g2_mux2_1 _2618_ (.A0(_0069_),
    .A1(_0947_),
    .S(_0786_),
    .X(_0326_));
 sg13g2_a22oi_1 _2619_ (.Y(_0948_),
    .B1(_0813_),
    .B2(_0921_),
    .A2(net817),
    .A1(\uart_0.rx.rx_samples[23] ));
 sg13g2_nor2_1 _2620_ (.A(net728),
    .B(_0943_),
    .Y(_0949_));
 sg13g2_a22oi_1 _2621_ (.Y(_0950_),
    .B1(_0948_),
    .B2(_0949_),
    .A2(net748),
    .A1(_0070_));
 sg13g2_inv_1 _2622_ (.Y(_0327_),
    .A(_0950_));
 sg13g2_nand3_1 _2623_ (.B(net787),
    .C(_0877_),
    .A(net756),
    .Y(_0951_));
 sg13g2_a21oi_1 _2624_ (.A1(_0864_),
    .A2(_0951_),
    .Y(_0952_),
    .B1(net769));
 sg13g2_nor2_1 _2625_ (.A(\uart_0.rx.rx_samples[24] ),
    .B(net783),
    .Y(_0953_));
 sg13g2_nor3_1 _2626_ (.A(net747),
    .B(_0952_),
    .C(_0953_),
    .Y(_0954_));
 sg13g2_a21oi_1 _2627_ (.A1(_1126_),
    .A2(net747),
    .Y(_0328_),
    .B1(_0954_));
 sg13g2_nand2_1 _2628_ (.Y(_0955_),
    .A(_0072_),
    .B(net748));
 sg13g2_nor2_2 _2629_ (.A(_0808_),
    .B(_0814_),
    .Y(_0956_));
 sg13g2_nand3_1 _2630_ (.B(_0832_),
    .C(_0956_),
    .A(net852),
    .Y(_0957_));
 sg13g2_nor3_1 _2631_ (.A(net785),
    .B(_0919_),
    .C(_0957_),
    .Y(_0958_));
 sg13g2_nor2_1 _2632_ (.A(\uart_0.rx.rx_samples[25] ),
    .B(net772),
    .Y(_0959_));
 sg13g2_o21ai_1 _2633_ (.B1(_0871_),
    .Y(_0960_),
    .A1(_0952_),
    .A2(_0959_));
 sg13g2_o21ai_1 _2634_ (.B1(_0955_),
    .Y(_0329_),
    .A1(_0958_),
    .A2(_0960_));
 sg13g2_a221oi_1 _2635_ (.B2(_0910_),
    .C1(_0882_),
    .B1(_0866_),
    .A1(\uart_0.rx.rx_samples[26] ),
    .Y(_0961_),
    .A2(net764));
 sg13g2_a21o_1 _2636_ (.A2(net741),
    .A1(_0073_),
    .B1(_0961_),
    .X(_0330_));
 sg13g2_nand2_1 _2637_ (.Y(_0962_),
    .A(_0074_),
    .B(net742));
 sg13g2_nand3_1 _2638_ (.B(_0811_),
    .C(_0921_),
    .A(_0800_),
    .Y(_0963_));
 sg13g2_a22oi_1 _2639_ (.Y(_0964_),
    .B1(_0866_),
    .B2(_0910_),
    .A2(net763),
    .A1(\uart_0.rx.rx_samples[27] ));
 sg13g2_nand2_1 _2640_ (.Y(_0965_),
    .A(_0963_),
    .B(_0964_));
 sg13g2_o21ai_1 _2641_ (.B1(_0962_),
    .Y(_0331_),
    .A1(_0882_),
    .A2(_0965_));
 sg13g2_nand2b_1 _2642_ (.Y(_0966_),
    .B(net756),
    .A_N(_0941_));
 sg13g2_a221oi_1 _2643_ (.B2(_0966_),
    .C1(net727),
    .B1(_0866_),
    .A1(\uart_0.rx.rx_samples[28] ),
    .Y(_0967_),
    .A2(net763));
 sg13g2_a21o_1 _2644_ (.A2(net740),
    .A1(_0075_),
    .B1(_0967_),
    .X(_0332_));
 sg13g2_and2_1 _2645_ (.A(net772),
    .B(_0916_),
    .X(_0968_));
 sg13g2_a221oi_1 _2646_ (.B2(_0968_),
    .C1(_0882_),
    .B1(_0920_),
    .A1(\uart_0.rx.rx_samples[29] ),
    .Y(_0969_),
    .A2(net763));
 sg13g2_a21o_1 _2647_ (.A2(net738),
    .A1(_0076_),
    .B1(_0969_),
    .X(_0333_));
 sg13g2_a21oi_1 _2648_ (.A1(\uart_0.rx.rx_samples[30] ),
    .A2(net762),
    .Y(_0970_),
    .B1(net725));
 sg13g2_a21o_1 _2649_ (.A2(net739),
    .A1(_0077_),
    .B1(_0970_),
    .X(_0334_));
 sg13g2_nor2_2 _2650_ (.A(net786),
    .B(net785),
    .Y(_0971_));
 sg13g2_and2_1 _2651_ (.A(net755),
    .B(_0971_),
    .X(_0972_));
 sg13g2_nand2_1 _2652_ (.Y(_0973_),
    .A(net755),
    .B(_0971_));
 sg13g2_nor2_2 _2653_ (.A(net760),
    .B(_0973_),
    .Y(_0974_));
 sg13g2_a221oi_1 _2654_ (.B2(_0974_),
    .C1(net725),
    .B1(_0868_),
    .A1(\uart_0.rx.rx_samples[31] ),
    .Y(_0975_),
    .A2(net817));
 sg13g2_a21o_1 _2655_ (.A2(net738),
    .A1(_0078_),
    .B1(_0975_),
    .X(_0335_));
 sg13g2_a21o_1 _2656_ (.A2(_0880_),
    .A1(_0860_),
    .B1(_0873_),
    .X(_0976_));
 sg13g2_a21oi_1 _2657_ (.A1(\uart_0.rx.rx_samples[32] ),
    .A2(net762),
    .Y(_0977_),
    .B1(_0976_));
 sg13g2_a21o_1 _2658_ (.A2(net738),
    .A1(_0079_),
    .B1(_0977_),
    .X(_0336_));
 sg13g2_a221oi_1 _2659_ (.B2(_0971_),
    .C1(_0976_),
    .B1(_0930_),
    .A1(\uart_0.rx.rx_samples[33] ),
    .Y(_0978_),
    .A2(net763));
 sg13g2_a21o_1 _2660_ (.A2(net740),
    .A1(_0080_),
    .B1(_0978_),
    .X(_0337_));
 sg13g2_a21oi_2 _2661_ (.B1(net732),
    .Y(_0979_),
    .A2(net786),
    .A1(_1167_));
 sg13g2_nand2_1 _2662_ (.Y(_0980_),
    .A(net755),
    .B(_0884_));
 sg13g2_a221oi_1 _2663_ (.B2(_0980_),
    .C1(net728),
    .B1(_0979_),
    .A1(\uart_0.rx.rx_samples[34] ),
    .Y(_0981_),
    .A2(net763));
 sg13g2_a21o_1 _2664_ (.A2(net736),
    .A1(_0081_),
    .B1(_0981_),
    .X(_0338_));
 sg13g2_a21o_1 _2665_ (.A2(_0974_),
    .A1(_0891_),
    .B1(net725),
    .X(_0982_));
 sg13g2_a21oi_1 _2666_ (.A1(\uart_0.rx.rx_samples[35] ),
    .A2(net817),
    .Y(_0983_),
    .B1(_0982_));
 sg13g2_a21o_1 _2667_ (.A2(net736),
    .A1(_0082_),
    .B1(_0983_),
    .X(_0339_));
 sg13g2_nand2_2 _2668_ (.Y(_0984_),
    .A(_0821_),
    .B(_0828_));
 sg13g2_nor3_1 _2669_ (.A(net756),
    .B(net787),
    .C(_0984_),
    .Y(_0985_));
 sg13g2_nor3_1 _2670_ (.A(net851),
    .B(\uart_0.rx.rx_stop_zeros[1] ),
    .C(_0028_),
    .Y(_0986_));
 sg13g2_nor2_1 _2671_ (.A(net760),
    .B(_0984_),
    .Y(_0987_));
 sg13g2_nand3_1 _2672_ (.B(_0986_),
    .C(_0987_),
    .A(_0878_),
    .Y(_0988_));
 sg13g2_a21oi_1 _2673_ (.A1(\uart_0.rx.rx_samples[36] ),
    .A2(net817),
    .Y(_0989_),
    .B1(_0982_));
 sg13g2_a22oi_1 _2674_ (.Y(_0990_),
    .B1(_0988_),
    .B2(_0989_),
    .A2(net736),
    .A1(_0083_));
 sg13g2_inv_1 _2675_ (.Y(_0340_),
    .A(_0990_));
 sg13g2_a221oi_1 _2676_ (.B2(_0972_),
    .C1(net725),
    .B1(_0900_),
    .A1(\uart_0.rx.rx_samples[37] ),
    .Y(_0991_),
    .A2(net817));
 sg13g2_a21o_1 _2677_ (.A2(net736),
    .A1(_0084_),
    .B1(_0991_),
    .X(_0341_));
 sg13g2_nor2_2 _2678_ (.A(net769),
    .B(_0826_),
    .Y(_0992_));
 sg13g2_o21ai_1 _2679_ (.B1(_0992_),
    .Y(_0993_),
    .A1(_0864_),
    .A2(_0985_));
 sg13g2_nand2_1 _2680_ (.Y(_0994_),
    .A(_0871_),
    .B(_0993_));
 sg13g2_a21oi_1 _2681_ (.A1(\uart_0.rx.rx_samples[38] ),
    .A2(net759),
    .Y(_0995_),
    .B1(_0994_));
 sg13g2_a21o_1 _2682_ (.A2(net735),
    .A1(_0085_),
    .B1(_0995_),
    .X(_0342_));
 sg13g2_a221oi_1 _2683_ (.B2(_0974_),
    .C1(_0994_),
    .B1(_0813_),
    .A1(\uart_0.rx.rx_samples[39] ),
    .Y(_0996_),
    .A2(net760));
 sg13g2_a21o_1 _2684_ (.A2(net735),
    .A1(_0086_),
    .B1(_0996_),
    .X(_0343_));
 sg13g2_nand2_1 _2685_ (.Y(_0997_),
    .A(\uart_0.rx.rx_samples[40] ),
    .B(net759));
 sg13g2_a21oi_1 _2686_ (.A1(_0860_),
    .A2(_0905_),
    .Y(_0998_),
    .B1(net725));
 sg13g2_a22oi_1 _2687_ (.Y(_0999_),
    .B1(_0997_),
    .B2(_0998_),
    .A2(net735),
    .A1(_0087_));
 sg13g2_inv_1 _2688_ (.Y(_0344_),
    .A(_0999_));
 sg13g2_nor2_1 _2689_ (.A(_0957_),
    .B(_0973_),
    .Y(_1000_));
 sg13g2_a21oi_1 _2690_ (.A1(\uart_0.rx.rx_samples[41] ),
    .A2(net759),
    .Y(_1001_),
    .B1(_1000_));
 sg13g2_a22oi_1 _2691_ (.Y(_1002_),
    .B1(_0998_),
    .B2(_1001_),
    .A2(net735),
    .A1(_0088_));
 sg13g2_inv_1 _2692_ (.Y(_0345_),
    .A(_1002_));
 sg13g2_nand2_1 _2693_ (.Y(_1003_),
    .A(net755),
    .B(_0909_));
 sg13g2_a221oi_1 _2694_ (.B2(_1003_),
    .C1(net728),
    .B1(_0979_),
    .A1(\uart_0.rx.rx_samples[42] ),
    .Y(_1004_),
    .A2(net760));
 sg13g2_a21o_1 _2695_ (.A2(net736),
    .A1(_0089_),
    .B1(_1004_),
    .X(_0346_));
 sg13g2_a221oi_1 _2696_ (.B2(_0974_),
    .C1(net725),
    .B1(_0912_),
    .A1(\uart_0.rx.rx_samples[43] ),
    .Y(_1005_),
    .A2(net817));
 sg13g2_a21o_1 _2697_ (.A2(net736),
    .A1(_0090_),
    .B1(_1005_),
    .X(_0347_));
 sg13g2_nor3_2 _2698_ (.A(net851),
    .B(net768),
    .C(_0984_),
    .Y(_1006_));
 sg13g2_and2_1 _2699_ (.A(_0802_),
    .B(_0808_),
    .X(_1007_));
 sg13g2_nand4_1 _2700_ (.B(_0820_),
    .C(_1006_),
    .A(net756),
    .Y(_1008_),
    .D(_1007_));
 sg13g2_a221oi_1 _2701_ (.B2(_0974_),
    .C1(net725),
    .B1(_0912_),
    .A1(\uart_0.rx.rx_samples[44] ),
    .Y(_1009_),
    .A2(net817));
 sg13g2_a22oi_1 _2702_ (.Y(_1010_),
    .B1(_1008_),
    .B2(_1009_),
    .A2(net736),
    .A1(_0091_));
 sg13g2_inv_1 _2703_ (.Y(_0348_),
    .A(_1010_));
 sg13g2_a221oi_1 _2704_ (.B2(_0972_),
    .C1(net725),
    .B1(_0968_),
    .A1(\uart_0.rx.rx_samples[45] ),
    .Y(_1011_),
    .A2(net760));
 sg13g2_a21o_1 _2705_ (.A2(net734),
    .A1(_0092_),
    .B1(_1011_),
    .X(_0349_));
 sg13g2_nand2_1 _2706_ (.Y(_1012_),
    .A(\uart_0.rx.rx_samples[46] ),
    .B(net758));
 sg13g2_nor2_1 _2707_ (.A(net728),
    .B(_0979_),
    .Y(_1013_));
 sg13g2_a22oi_1 _2708_ (.Y(_1014_),
    .B1(_1012_),
    .B2(net721),
    .A2(net733),
    .A1(_0093_));
 sg13g2_inv_1 _2709_ (.Y(_0350_),
    .A(_1014_));
 sg13g2_o21ai_1 _2710_ (.B1(net722),
    .Y(_1015_),
    .A1(_0869_),
    .A2(_0934_));
 sg13g2_a21oi_1 _2711_ (.A1(\uart_0.rx.rx_samples[47] ),
    .A2(net759),
    .Y(_1016_),
    .B1(_1015_));
 sg13g2_a21o_1 _2712_ (.A2(net735),
    .A1(_0094_),
    .B1(_1016_),
    .X(_0351_));
 sg13g2_a221oi_1 _2713_ (.B2(_1006_),
    .C1(_1015_),
    .B1(_0924_),
    .A1(\uart_0.rx.rx_samples[48] ),
    .Y(_1017_),
    .A2(net759));
 sg13g2_a21o_1 _2714_ (.A2(net735),
    .A1(_0095_),
    .B1(_1017_),
    .X(_0352_));
 sg13g2_a21oi_1 _2715_ (.A1(\uart_0.rx.rx_samples[49] ),
    .A2(net759),
    .Y(_1018_),
    .B1(_0885_));
 sg13g2_a22oi_1 _2716_ (.Y(_1019_),
    .B1(net721),
    .B2(_1018_),
    .A2(net733),
    .A1(_0096_));
 sg13g2_inv_1 _2717_ (.Y(_0353_),
    .A(_1019_));
 sg13g2_a22oi_1 _2718_ (.Y(_1020_),
    .B1(_0860_),
    .B2(_0883_),
    .A2(net758),
    .A1(\uart_0.rx.rx_samples[50] ));
 sg13g2_a22oi_1 _2719_ (.Y(_1021_),
    .B1(net722),
    .B2(_1020_),
    .A2(net733),
    .A1(_0097_));
 sg13g2_inv_1 _2720_ (.Y(_0354_),
    .A(_1021_));
 sg13g2_o21ai_1 _2721_ (.B1(net722),
    .Y(_1022_),
    .A1(net732),
    .A2(_0890_));
 sg13g2_a21oi_1 _2722_ (.A1(\uart_0.rx.rx_samples[51] ),
    .A2(net759),
    .Y(_1023_),
    .B1(_1022_));
 sg13g2_a21o_1 _2723_ (.A2(net735),
    .A1(_0098_),
    .B1(_1023_),
    .X(_0355_));
 sg13g2_nor2b_2 _2724_ (.A(_0923_),
    .B_N(_1007_),
    .Y(_1024_));
 sg13g2_a221oi_1 _2725_ (.B2(_1024_),
    .C1(_1022_),
    .B1(_1006_),
    .A1(\uart_0.rx.rx_samples[52] ),
    .Y(_1025_),
    .A2(net759));
 sg13g2_a21o_1 _2726_ (.A2(net733),
    .A1(_0099_),
    .B1(_1025_),
    .X(_0356_));
 sg13g2_nand2_1 _2727_ (.Y(_1026_),
    .A(_0901_),
    .B(net721));
 sg13g2_a21oi_1 _2728_ (.A1(\uart_0.rx.rx_samples[53] ),
    .A2(net758),
    .Y(_1027_),
    .B1(_1026_));
 sg13g2_a21o_1 _2729_ (.A2(net733),
    .A1(_0100_),
    .B1(_1027_),
    .X(_0357_));
 sg13g2_nand4_1 _2730_ (.B(net786),
    .C(_0898_),
    .A(_0814_),
    .Y(_1028_),
    .D(_0987_));
 sg13g2_a21oi_1 _2731_ (.A1(\uart_0.rx.rx_samples[54] ),
    .A2(net817),
    .Y(_1029_),
    .B1(_1026_));
 sg13g2_a22oi_1 _2732_ (.Y(_1030_),
    .B1(_1028_),
    .B2(_1029_),
    .A2(net733),
    .A1(_0101_));
 sg13g2_inv_1 _2733_ (.Y(_0358_),
    .A(_1030_));
 sg13g2_o21ai_1 _2734_ (.B1(net722),
    .Y(_1031_),
    .A1(_0811_),
    .A2(net732));
 sg13g2_a21oi_1 _2735_ (.A1(\uart_0.rx.rx_samples[55] ),
    .A2(net758),
    .Y(_1032_),
    .B1(_1031_));
 sg13g2_a21o_1 _2736_ (.A2(net734),
    .A1(_0102_),
    .B1(_1032_),
    .X(_0359_));
 sg13g2_nand3_1 _2737_ (.B(_0942_),
    .C(_1006_),
    .A(_0876_),
    .Y(_1033_));
 sg13g2_a21oi_1 _2738_ (.A1(\uart_0.rx.rx_samples[56] ),
    .A2(net758),
    .Y(_1034_),
    .B1(_1031_));
 sg13g2_a22oi_1 _2739_ (.Y(_1035_),
    .B1(_1033_),
    .B2(_1034_),
    .A2(net733),
    .A1(_0103_));
 sg13g2_inv_1 _2740_ (.Y(_0360_),
    .A(_1035_));
 sg13g2_a21oi_1 _2741_ (.A1(\uart_0.rx.rx_samples[57] ),
    .A2(net761),
    .Y(_1036_),
    .B1(_0907_));
 sg13g2_a22oi_1 _2742_ (.Y(_1037_),
    .B1(net721),
    .B2(_1036_),
    .A2(net734),
    .A1(_0104_));
 sg13g2_inv_1 _2743_ (.Y(_0361_),
    .A(_1037_));
 sg13g2_a22oi_1 _2744_ (.Y(_1038_),
    .B1(_0860_),
    .B2(_0910_),
    .A2(net761),
    .A1(\uart_0.rx.rx_samples[58] ));
 sg13g2_a22oi_1 _2745_ (.Y(_1039_),
    .B1(net721),
    .B2(_1038_),
    .A2(net734),
    .A1(_0105_));
 sg13g2_inv_1 _2746_ (.Y(_0362_),
    .A(_1039_));
 sg13g2_nand2_1 _2747_ (.Y(_1040_),
    .A(\uart_0.rx.rx_samples[59] ),
    .B(net758));
 sg13g2_nand2_1 _2748_ (.Y(_1041_),
    .A(_0912_),
    .B(_0935_));
 sg13g2_nand3_1 _2749_ (.B(_1040_),
    .C(_1041_),
    .A(net721),
    .Y(_1042_));
 sg13g2_o21ai_1 _2750_ (.B1(_1042_),
    .Y(_0363_),
    .A1(_1125_),
    .A2(_0786_));
 sg13g2_nand3_1 _2751_ (.B(_0986_),
    .C(_0987_),
    .A(_0942_),
    .Y(_1043_));
 sg13g2_nand3_1 _2752_ (.B(_1041_),
    .C(_1043_),
    .A(net721),
    .Y(_1044_));
 sg13g2_a21oi_1 _2753_ (.A1(\uart_0.rx.rx_samples[60] ),
    .A2(net758),
    .Y(_1045_),
    .B1(_1044_));
 sg13g2_a21o_1 _2754_ (.A2(net734),
    .A1(_0107_),
    .B1(_1045_),
    .X(_0364_));
 sg13g2_a22oi_1 _2755_ (.Y(_1046_),
    .B1(_0860_),
    .B2(_0916_),
    .A2(net761),
    .A1(\uart_0.rx.rx_samples[61] ));
 sg13g2_a22oi_1 _2756_ (.Y(_1047_),
    .B1(net721),
    .B2(_1046_),
    .A2(net733),
    .A1(_0108_));
 sg13g2_inv_1 _2757_ (.Y(_0365_),
    .A(_1047_));
 sg13g2_a21oi_1 _2758_ (.A1(\uart_0.rx.rx_samples[62] ),
    .A2(net758),
    .Y(_1048_),
    .B1(_0935_));
 sg13g2_a21o_1 _2759_ (.A2(net735),
    .A1(_0109_),
    .B1(_1048_),
    .X(_0366_));
 sg13g2_and2_1 _2760_ (.A(net772),
    .B(net785),
    .X(_1049_));
 sg13g2_nand2b_2 _2761_ (.Y(_1050_),
    .B(_0862_),
    .A_N(_0828_));
 sg13g2_o21ai_1 _2762_ (.B1(_1049_),
    .Y(_1051_),
    .A1(_0869_),
    .A2(_1050_));
 sg13g2_o21ai_1 _2763_ (.B1(_1051_),
    .Y(_1052_),
    .A1(\uart_0.rx.rx_samples[63] ),
    .A2(net772));
 sg13g2_a22oi_1 _2764_ (.Y(_1053_),
    .B1(_0871_),
    .B2(_1052_),
    .A2(net746),
    .A1(_0110_));
 sg13g2_inv_1 _2765_ (.Y(_0367_),
    .A(_1053_));
 sg13g2_nor3_2 _2766_ (.A(net767),
    .B(_0821_),
    .C(_0826_),
    .Y(_1054_));
 sg13g2_a21oi_2 _2767_ (.B1(net724),
    .Y(_1055_),
    .A2(_1054_),
    .A1(_0878_));
 sg13g2_a21oi_1 _2768_ (.A1(_0877_),
    .A2(_0934_),
    .Y(_1056_),
    .B1(_1055_));
 sg13g2_a21oi_1 _2769_ (.A1(\uart_0.rx.rx_samples[64] ),
    .A2(net767),
    .Y(_1057_),
    .B1(_1056_));
 sg13g2_a21o_1 _2770_ (.A2(net743),
    .A1(_0111_),
    .B1(_1057_),
    .X(_0368_));
 sg13g2_nor2_2 _2771_ (.A(_0929_),
    .B(_1050_),
    .Y(_1058_));
 sg13g2_a221oi_1 _2772_ (.B2(_1058_),
    .C1(_1056_),
    .B1(_0883_),
    .A1(\uart_0.rx.rx_samples[65] ),
    .Y(_1059_),
    .A2(net767));
 sg13g2_a21o_1 _2773_ (.A2(net743),
    .A1(_0112_),
    .B1(_1059_),
    .X(_0369_));
 sg13g2_o21ai_1 _2774_ (.B1(_1049_),
    .Y(_1060_),
    .A1(_0884_),
    .A2(_1050_));
 sg13g2_o21ai_1 _2775_ (.B1(_1060_),
    .Y(_1061_),
    .A1(\uart_0.rx.rx_samples[66] ),
    .A2(net772));
 sg13g2_a22oi_1 _2776_ (.Y(_1062_),
    .B1(_0871_),
    .B2(_1061_),
    .A2(net746),
    .A1(_0113_));
 sg13g2_inv_1 _2777_ (.Y(_0370_),
    .A(_1062_));
 sg13g2_nor2_2 _2778_ (.A(net768),
    .B(_1050_),
    .Y(_1063_));
 sg13g2_a221oi_1 _2779_ (.B2(_1063_),
    .C1(net723),
    .B1(_0891_),
    .A1(\uart_0.rx.rx_samples[67] ),
    .Y(_1064_),
    .A2(net767));
 sg13g2_a21o_1 _2780_ (.A2(net743),
    .A1(_0114_),
    .B1(_1064_),
    .X(_0371_));
 sg13g2_nand2_1 _2781_ (.Y(_1065_),
    .A(\uart_0.rx.rx_samples[68] ),
    .B(net767));
 sg13g2_nand3_1 _2782_ (.B(_0871_),
    .C(_0893_),
    .A(net785),
    .Y(_1066_));
 sg13g2_nand2b_1 _2783_ (.Y(_1067_),
    .B(_1066_),
    .A_N(_1055_));
 sg13g2_a22oi_1 _2784_ (.Y(_1068_),
    .B1(_1065_),
    .B2(_1067_),
    .A2(net743),
    .A1(_0115_));
 sg13g2_inv_1 _2785_ (.Y(_0372_),
    .A(_1068_));
 sg13g2_a22oi_1 _2786_ (.Y(_1069_),
    .B1(_0888_),
    .B2(_1058_),
    .A2(net767),
    .A1(\uart_0.rx.rx_samples[69] ));
 sg13g2_a22oi_1 _2787_ (.Y(_1070_),
    .B1(_1067_),
    .B2(_1069_),
    .A2(net743),
    .A1(_0116_));
 sg13g2_inv_1 _2788_ (.Y(_0373_),
    .A(_1070_));
 sg13g2_nand2_1 _2789_ (.Y(_1071_),
    .A(\uart_0.rx.rx_samples[70] ),
    .B(net767));
 sg13g2_a22oi_1 _2790_ (.Y(_1072_),
    .B1(_1055_),
    .B2(_1071_),
    .A2(net743),
    .A1(_0117_));
 sg13g2_inv_1 _2791_ (.Y(_0374_),
    .A(_1072_));
 sg13g2_a22oi_1 _2792_ (.Y(_1073_),
    .B1(_0813_),
    .B2(_1063_),
    .A2(net767),
    .A1(\uart_0.rx.rx_samples[71] ));
 sg13g2_a22oi_1 _2793_ (.Y(_1074_),
    .B1(_1055_),
    .B2(_1073_),
    .A2(net743),
    .A1(_0118_));
 sg13g2_inv_1 _2794_ (.Y(_0375_),
    .A(_1074_));
 sg13g2_a21o_1 _2795_ (.A2(_1054_),
    .A1(_0905_),
    .B1(net723),
    .X(_1075_));
 sg13g2_a21oi_1 _2796_ (.A1(\uart_0.rx.rx_samples[72] ),
    .A2(net768),
    .Y(_1076_),
    .B1(_1075_));
 sg13g2_a21o_1 _2797_ (.A2(net744),
    .A1(_0119_),
    .B1(_1076_),
    .X(_0376_));
 sg13g2_a221oi_1 _2798_ (.B2(_1058_),
    .C1(_1075_),
    .B1(_0956_),
    .A1(\uart_0.rx.rx_samples[73] ),
    .Y(_1077_),
    .A2(net768));
 sg13g2_a21o_1 _2799_ (.A2(net744),
    .A1(_0120_),
    .B1(_1077_),
    .X(_0377_));
 sg13g2_a221oi_1 _2800_ (.B2(_1063_),
    .C1(net723),
    .B1(_0910_),
    .A1(\uart_0.rx.rx_samples[74] ),
    .Y(_1078_),
    .A2(net815));
 sg13g2_a21o_1 _2801_ (.A2(net744),
    .A1(_0121_),
    .B1(_1078_),
    .X(_0378_));
 sg13g2_a221oi_1 _2802_ (.B2(_1063_),
    .C1(net723),
    .B1(_0912_),
    .A1(\uart_0.rx.rx_samples[75] ),
    .Y(_1079_),
    .A2(net815));
 sg13g2_a21o_1 _2803_ (.A2(net744),
    .A1(_0122_),
    .B1(_1079_),
    .X(_0379_));
 sg13g2_nand2_1 _2804_ (.Y(_1080_),
    .A(\uart_0.rx.rx_samples[76] ),
    .B(net768));
 sg13g2_a21oi_2 _2805_ (.B1(net723),
    .Y(_1081_),
    .A2(_1054_),
    .A1(_0914_));
 sg13g2_a22oi_1 _2806_ (.Y(_1082_),
    .B1(_1080_),
    .B2(_1081_),
    .A2(net744),
    .A1(_0123_));
 sg13g2_inv_1 _2807_ (.Y(_0380_),
    .A(_1082_));
 sg13g2_a22oi_1 _2808_ (.Y(_1083_),
    .B1(_0909_),
    .B2(_1058_),
    .A2(net768),
    .A1(\uart_0.rx.rx_samples[77] ));
 sg13g2_a22oi_1 _2809_ (.Y(_1084_),
    .B1(_1081_),
    .B2(_1083_),
    .A2(net746),
    .A1(_0124_));
 sg13g2_inv_1 _2810_ (.Y(_0381_),
    .A(_1084_));
 sg13g2_o21ai_1 _2811_ (.B1(_0786_),
    .Y(_1085_),
    .A1(\uart_0.rx.rx_samples[78] ),
    .A2(net783));
 sg13g2_a21oi_1 _2812_ (.A1(_1049_),
    .A2(_1050_),
    .Y(_1086_),
    .B1(_1085_));
 sg13g2_a21oi_1 _2813_ (.A1(_1124_),
    .A2(net743),
    .Y(_0382_),
    .B1(_1086_));
 sg13g2_nor2_2 _2814_ (.A(net723),
    .B(_1063_),
    .Y(_1087_));
 sg13g2_nor2_1 _2815_ (.A(_0828_),
    .B(_0919_),
    .Y(_1088_));
 sg13g2_nand2_1 _2816_ (.Y(_1089_),
    .A(net772),
    .B(_1088_));
 sg13g2_nor2_1 _2817_ (.A(_0869_),
    .B(_1089_),
    .Y(_1090_));
 sg13g2_a21oi_1 _2818_ (.A1(\uart_0.rx.rx_samples[79] ),
    .A2(net815),
    .Y(_1091_),
    .B1(_1090_));
 sg13g2_a22oi_1 _2819_ (.Y(_1092_),
    .B1(_1087_),
    .B2(_1091_),
    .A2(net744),
    .A1(_0126_));
 sg13g2_inv_1 _2820_ (.Y(_0383_),
    .A(_1092_));
 sg13g2_a21oi_1 _2821_ (.A1(_0925_),
    .A2(_1054_),
    .Y(_1093_),
    .B1(net723));
 sg13g2_a221oi_1 _2822_ (.B2(_1054_),
    .C1(net723),
    .B1(_0925_),
    .A1(\uart_0.rx.rx_samples[80] ),
    .Y(_1094_),
    .A2(net815));
 sg13g2_a21o_1 _2823_ (.A2(net745),
    .A1(_0127_),
    .B1(_1094_),
    .X(_0384_));
 sg13g2_a22oi_1 _2824_ (.Y(_1095_),
    .B1(_0930_),
    .B2(_1088_),
    .A2(net815),
    .A1(\uart_0.rx.rx_samples[81] ));
 sg13g2_a22oi_1 _2825_ (.Y(_1096_),
    .B1(_1093_),
    .B2(_1095_),
    .A2(net744),
    .A1(_0128_));
 sg13g2_inv_1 _2826_ (.Y(_0385_),
    .A(_1096_));
 sg13g2_a221oi_1 _2827_ (.B2(_0992_),
    .C1(net724),
    .B1(_0936_),
    .A1(\uart_0.rx.rx_samples[82] ),
    .Y(_1097_),
    .A2(net770));
 sg13g2_a21o_1 _2828_ (.A2(net744),
    .A1(_0129_),
    .B1(_1097_),
    .X(_0386_));
 sg13g2_nor2_1 _2829_ (.A(_0890_),
    .B(_1089_),
    .Y(_1098_));
 sg13g2_a21oi_1 _2830_ (.A1(\uart_0.rx.rx_samples[83] ),
    .A2(net815),
    .Y(_1099_),
    .B1(_1098_));
 sg13g2_a22oi_1 _2831_ (.Y(_1100_),
    .B1(_1087_),
    .B2(_1099_),
    .A2(net745),
    .A1(_0130_));
 sg13g2_inv_1 _2832_ (.Y(_0387_),
    .A(_1100_));
 sg13g2_nor3_2 _2833_ (.A(net851),
    .B(_1167_),
    .C(_0031_),
    .Y(_1101_));
 sg13g2_and2_1 _2834_ (.A(net772),
    .B(_1101_),
    .X(_1102_));
 sg13g2_a221oi_1 _2835_ (.B2(_1102_),
    .C1(_1098_),
    .B1(_1024_),
    .A1(\uart_0.rx.rx_samples[84] ),
    .Y(_1103_),
    .A2(net815));
 sg13g2_a22oi_1 _2836_ (.Y(_1104_),
    .B1(_1087_),
    .B2(_1103_),
    .A2(net745),
    .A1(_0131_));
 sg13g2_inv_1 _2837_ (.Y(_0388_),
    .A(_1104_));
 sg13g2_and2_1 _2838_ (.A(_0132_),
    .B(net749),
    .X(_1105_));
 sg13g2_nand2_1 _2839_ (.Y(_1106_),
    .A(\uart_0.rx.rx_samples[85] ),
    .B(net771));
 sg13g2_and2_1 _2840_ (.A(_0900_),
    .B(_1088_),
    .X(_1107_));
 sg13g2_nor3_2 _2841_ (.A(net724),
    .B(_1063_),
    .C(_1107_),
    .Y(_1108_));
 sg13g2_a21o_1 _2842_ (.A2(_1108_),
    .A1(_1106_),
    .B1(_1105_),
    .X(_0389_));
 sg13g2_nor3_2 _2843_ (.A(net769),
    .B(_0894_),
    .C(_0923_),
    .Y(_1109_));
 sg13g2_a22oi_1 _2844_ (.Y(_1110_),
    .B1(_1101_),
    .B2(_1109_),
    .A2(net769),
    .A1(\uart_0.rx.rx_samples[86] ));
 sg13g2_a22oi_1 _2845_ (.Y(_1111_),
    .B1(_1108_),
    .B2(_1110_),
    .A2(net749),
    .A1(_0133_));
 sg13g2_inv_1 _2846_ (.Y(_0390_),
    .A(_1111_));
 sg13g2_o21ai_1 _2847_ (.B1(_1087_),
    .Y(_1112_),
    .A1(_0811_),
    .A2(_1089_));
 sg13g2_a21oi_1 _2848_ (.A1(\uart_0.rx.rx_samples[87] ),
    .A2(net771),
    .Y(_1113_),
    .B1(_1112_));
 sg13g2_a21o_1 _2849_ (.A2(net745),
    .A1(_0134_),
    .B1(_1113_),
    .X(_0391_));
 sg13g2_nor3_1 _2850_ (.A(net852),
    .B(\uart_0.rx.rx_stop_zeros[1] ),
    .C(_1089_),
    .Y(_1114_));
 sg13g2_a221oi_1 _2851_ (.B2(_1114_),
    .C1(_1112_),
    .B1(_0956_),
    .A1(\uart_0.rx.rx_samples[88] ),
    .Y(_1115_),
    .A2(net768));
 sg13g2_a21o_1 _2852_ (.A2(net745),
    .A1(_0135_),
    .B1(_1115_),
    .X(_0392_));
 sg13g2_nor2_1 _2853_ (.A(_1143_),
    .B(_0768_),
    .Y(_1116_));
 sg13g2_a21oi_1 _2854_ (.A1(_1143_),
    .A2(_0771_),
    .Y(_0393_),
    .B1(_1116_));
 sg13g2_nand2_1 _2855_ (.Y(_1117_),
    .A(\uart_0.rx.rx_sample_cnt[1] ),
    .B(_0768_));
 sg13g2_nand2_1 _2856_ (.Y(_1118_),
    .A(\uart_0.rx.rx_sample_cnt[1] ),
    .B(_1116_));
 sg13g2_o21ai_1 _2857_ (.B1(_1118_),
    .Y(_1119_),
    .A1(\uart_0.rx.rx_sample_cnt[0] ),
    .A2(\uart_0.rx.rx_sample_cnt[1] ));
 sg13g2_a21oi_1 _2858_ (.A1(_0771_),
    .A2(_1117_),
    .Y(_0394_),
    .B1(_1119_));
 sg13g2_nor3_1 _2859_ (.A(\uart_0.rx.rx_sample_cnt[3] ),
    .B(net783),
    .C(_0764_),
    .Y(_1120_));
 sg13g2_a21oi_1 _2860_ (.A1(_0770_),
    .A2(_1120_),
    .Y(_1121_),
    .B1(_0768_));
 sg13g2_a21oi_1 _2861_ (.A1(_1142_),
    .A2(_1118_),
    .Y(_0395_),
    .B1(_1121_));
 sg13g2_nand2_1 _2862_ (.Y(_1122_),
    .A(\uart_0.rx.rx_sample_cnt[3] ),
    .B(_0768_));
 sg13g2_nand2_1 _2863_ (.Y(_0396_),
    .A(_0772_),
    .B(_1122_));
 sg13g2_and2_1 _2864_ (.A(\uart_0.rx.rx_sample_cnt[4] ),
    .B(_0768_),
    .X(_0397_));
 sg13g2_and2_1 _2865_ (.A(\uart_0.rx.rx_sample_cnt[5] ),
    .B(net816),
    .X(_0398_));
 sg13g2_and2_1 _2866_ (.A(\uart_0.rx.rx_sample_cnt[6] ),
    .B(_0768_),
    .X(_0399_));
 sg13g2_a21oi_1 _2867_ (.A1(net847),
    .A2(_1389_),
    .Y(_1123_),
    .B1(net773));
 sg13g2_o21ai_1 _2868_ (.B1(_1123_),
    .Y(_0400_),
    .A1(_1169_),
    .A2(_0834_));
 sg13g2_dfrbp_1 _2869_ (.CLK(clknet_1_0__leaf_clk),
    .RESET_B(net927),
    .D(net23),
    .Q_N(_0038_),
    .Q(clk_out));
 sg13g2_dfrbp_1 _2870_ (.CLK(net877),
    .RESET_B(net918),
    .D(net754),
    .Q_N(_1554_),
    .Q(tx_do));
 sg13g2_dfrbp_1 _2871_ (.CLK(net879),
    .RESET_B(net918),
    .D(_0004_),
    .Q_N(_1555_),
    .Q(\tx_data[0] ));
 sg13g2_dfrbp_1 _2872_ (.CLK(net876),
    .RESET_B(net916),
    .D(_0005_),
    .Q_N(_1556_),
    .Q(\tx_data[1] ));
 sg13g2_dfrbp_1 _2873_ (.CLK(net877),
    .RESET_B(net918),
    .D(_0006_),
    .Q_N(_1557_),
    .Q(\tx_data[2] ));
 sg13g2_dfrbp_1 _2874_ (.CLK(net870),
    .RESET_B(net909),
    .D(_0007_),
    .Q_N(_1558_),
    .Q(\tx_data[3] ));
 sg13g2_dfrbp_1 _2875_ (.CLK(net877),
    .RESET_B(net918),
    .D(_0008_),
    .Q_N(_1559_),
    .Q(\tx_data[4] ));
 sg13g2_dfrbp_1 _2876_ (.CLK(net871),
    .RESET_B(net910),
    .D(_0009_),
    .Q_N(_1560_),
    .Q(\tx_data[5] ));
 sg13g2_dfrbp_1 _2877_ (.CLK(net871),
    .RESET_B(net919),
    .D(_0010_),
    .Q_N(_1561_),
    .Q(\tx_data[6] ));
 sg13g2_dfrbp_1 _2878_ (.CLK(net876),
    .RESET_B(net918),
    .D(_0011_),
    .Q_N(_1553_),
    .Q(\tx_data[7] ));
 sg13g2_dfrbp_1 _2879_ (.CLK(net869),
    .RESET_B(net910),
    .D(_0139_),
    .Q_N(_0040_),
    .Q(\fifo_h[0] ));
 sg13g2_dfrbp_1 _2880_ (.CLK(net869),
    .RESET_B(net910),
    .D(_0140_),
    .Q_N(_1552_),
    .Q(\fifo_h[1] ));
 sg13g2_dfrbp_1 _2881_ (.CLK(net869),
    .RESET_B(net910),
    .D(_0141_),
    .Q_N(_1551_),
    .Q(\fifo_h[2] ));
 sg13g2_dfrbp_1 _2882_ (.CLK(net869),
    .RESET_B(net910),
    .D(_0142_),
    .Q_N(_1550_),
    .Q(\fifo_h[3] ));
 sg13g2_dfrbp_1 _2883_ (.CLK(net833),
    .RESET_B(net893),
    .D(_0143_),
    .Q_N(_0039_),
    .Q(\fifo_t[0] ));
 sg13g2_dfrbp_1 _2884_ (.CLK(net833),
    .RESET_B(net892),
    .D(_0144_),
    .Q_N(_1549_),
    .Q(\fifo_t[1] ));
 sg13g2_dfrbp_1 _2885_ (.CLK(net833),
    .RESET_B(net893),
    .D(_0145_),
    .Q_N(_1548_),
    .Q(\fifo_t[2] ));
 sg13g2_dfrbp_1 _2886_ (.CLK(net833),
    .RESET_B(net892),
    .D(_0146_),
    .Q_N(_1547_),
    .Q(\fifo_t[3] ));
 sg13g2_dfrbp_1 _2887_ (.CLK(net844),
    .RESET_B(net917),
    .D(_0147_),
    .Q_N(_1546_),
    .Q(\fifo_d[0][0] ));
 sg13g2_dfrbp_1 _2888_ (.CLK(net844),
    .RESET_B(net916),
    .D(_0148_),
    .Q_N(_1545_),
    .Q(\fifo_d[0][1] ));
 sg13g2_dfrbp_1 _2889_ (.CLK(net844),
    .RESET_B(net917),
    .D(_0149_),
    .Q_N(_1544_),
    .Q(\fifo_d[0][2] ));
 sg13g2_dfrbp_1 _2890_ (.CLK(net840),
    .RESET_B(net910),
    .D(_0150_),
    .Q_N(_1543_),
    .Q(\fifo_d[0][3] ));
 sg13g2_dfrbp_1 _2891_ (.CLK(net844),
    .RESET_B(net917),
    .D(_0151_),
    .Q_N(_1542_),
    .Q(\fifo_d[0][4] ));
 sg13g2_dfrbp_1 _2892_ (.CLK(net839),
    .RESET_B(net909),
    .D(_0152_),
    .Q_N(_1541_),
    .Q(\fifo_d[0][5] ));
 sg13g2_dfrbp_1 _2893_ (.CLK(net839),
    .RESET_B(net910),
    .D(_0153_),
    .Q_N(_1540_),
    .Q(\fifo_d[0][6] ));
 sg13g2_dfrbp_1 _2894_ (.CLK(net840),
    .RESET_B(net918),
    .D(_0154_),
    .Q_N(_1539_),
    .Q(\fifo_d[0][7] ));
 sg13g2_dfrbp_1 _2895_ (.CLK(net826),
    .RESET_B(net888),
    .D(_0155_),
    .Q_N(_1538_),
    .Q(\fifo_d[1][0] ));
 sg13g2_dfrbp_1 _2896_ (.CLK(net827),
    .RESET_B(net886),
    .D(_0156_),
    .Q_N(_1537_),
    .Q(\fifo_d[1][1] ));
 sg13g2_dfrbp_1 _2897_ (.CLK(net827),
    .RESET_B(net885),
    .D(_0157_),
    .Q_N(_1536_),
    .Q(\fifo_d[1][2] ));
 sg13g2_dfrbp_1 _2898_ (.CLK(net832),
    .RESET_B(net907),
    .D(_0158_),
    .Q_N(_1535_),
    .Q(\fifo_d[1][3] ));
 sg13g2_dfrbp_1 _2899_ (.CLK(net839),
    .RESET_B(net909),
    .D(_0159_),
    .Q_N(_1534_),
    .Q(\fifo_d[1][4] ));
 sg13g2_dfrbp_1 _2900_ (.CLK(net839),
    .RESET_B(net907),
    .D(_0160_),
    .Q_N(_1533_),
    .Q(\fifo_d[1][5] ));
 sg13g2_dfrbp_1 _2901_ (.CLK(net824),
    .RESET_B(net885),
    .D(_0161_),
    .Q_N(_1532_),
    .Q(\fifo_d[1][6] ));
 sg13g2_dfrbp_1 _2902_ (.CLK(net830),
    .RESET_B(net890),
    .D(_0162_),
    .Q_N(_1531_),
    .Q(\fifo_d[1][7] ));
 sg13g2_dfrbp_1 _2903_ (.CLK(net826),
    .RESET_B(net888),
    .D(_0163_),
    .Q_N(_1530_),
    .Q(\fifo_d[2][0] ));
 sg13g2_dfrbp_1 _2904_ (.CLK(net841),
    .RESET_B(net912),
    .D(_0164_),
    .Q_N(_1529_),
    .Q(\fifo_d[2][1] ));
 sg13g2_dfrbp_1 _2905_ (.CLK(net837),
    .RESET_B(net911),
    .D(_0165_),
    .Q_N(_1528_),
    .Q(\fifo_d[2][2] ));
 sg13g2_dfrbp_1 _2906_ (.CLK(net831),
    .RESET_B(net905),
    .D(_0166_),
    .Q_N(_1527_),
    .Q(\fifo_d[2][3] ));
 sg13g2_dfrbp_1 _2907_ (.CLK(net826),
    .RESET_B(net888),
    .D(_0167_),
    .Q_N(_1526_),
    .Q(\fifo_d[2][4] ));
 sg13g2_dfrbp_1 _2908_ (.CLK(net829),
    .RESET_B(net889),
    .D(_0168_),
    .Q_N(_1525_),
    .Q(\fifo_d[2][5] ));
 sg13g2_dfrbp_1 _2909_ (.CLK(net835),
    .RESET_B(net906),
    .D(_0169_),
    .Q_N(_1524_),
    .Q(\fifo_d[2][6] ));
 sg13g2_dfrbp_1 _2910_ (.CLK(net841),
    .RESET_B(net912),
    .D(_0170_),
    .Q_N(_1523_),
    .Q(\fifo_d[2][7] ));
 sg13g2_dfrbp_1 _2911_ (.CLK(net843),
    .RESET_B(net914),
    .D(_0171_),
    .Q_N(_1522_),
    .Q(\fifo_d[3][0] ));
 sg13g2_dfrbp_1 _2912_ (.CLK(net827),
    .RESET_B(net886),
    .D(_0172_),
    .Q_N(_1521_),
    .Q(\fifo_d[3][1] ));
 sg13g2_dfrbp_1 _2913_ (.CLK(net827),
    .RESET_B(net885),
    .D(_0173_),
    .Q_N(_1520_),
    .Q(\fifo_d[3][2] ));
 sg13g2_dfrbp_1 _2914_ (.CLK(net837),
    .RESET_B(net908),
    .D(_0174_),
    .Q_N(_1519_),
    .Q(\fifo_d[3][3] ));
 sg13g2_dfrbp_1 _2915_ (.CLK(net825),
    .RESET_B(net884),
    .D(_0175_),
    .Q_N(_1518_),
    .Q(\fifo_d[3][4] ));
 sg13g2_dfrbp_1 _2916_ (.CLK(net829),
    .RESET_B(net888),
    .D(_0176_),
    .Q_N(_1517_),
    .Q(\fifo_d[3][5] ));
 sg13g2_dfrbp_1 _2917_ (.CLK(net824),
    .RESET_B(net884),
    .D(_0177_),
    .Q_N(_1516_),
    .Q(\fifo_d[3][6] ));
 sg13g2_dfrbp_1 _2918_ (.CLK(net844),
    .RESET_B(net915),
    .D(_0178_),
    .Q_N(_1515_),
    .Q(\fifo_d[3][7] ));
 sg13g2_dfrbp_1 _2919_ (.CLK(net824),
    .RESET_B(net887),
    .D(_0179_),
    .Q_N(_1514_),
    .Q(\fifo_d[4][0] ));
 sg13g2_dfrbp_1 _2920_ (.CLK(net824),
    .RESET_B(net885),
    .D(_0180_),
    .Q_N(_1513_),
    .Q(\fifo_d[4][1] ));
 sg13g2_dfrbp_1 _2921_ (.CLK(net824),
    .RESET_B(net885),
    .D(_0181_),
    .Q_N(_1512_),
    .Q(\fifo_d[4][2] ));
 sg13g2_dfrbp_1 _2922_ (.CLK(net831),
    .RESET_B(net905),
    .D(_0182_),
    .Q_N(_1511_),
    .Q(\fifo_d[4][3] ));
 sg13g2_dfrbp_1 _2923_ (.CLK(net825),
    .RESET_B(net885),
    .D(_0183_),
    .Q_N(_1510_),
    .Q(\fifo_d[4][4] ));
 sg13g2_dfrbp_1 _2924_ (.CLK(net831),
    .RESET_B(net905),
    .D(_0184_),
    .Q_N(_1509_),
    .Q(\fifo_d[4][5] ));
 sg13g2_dfrbp_1 _2925_ (.CLK(net825),
    .RESET_B(net884),
    .D(_0185_),
    .Q_N(_1508_),
    .Q(\fifo_d[4][6] ));
 sg13g2_dfrbp_1 _2926_ (.CLK(net825),
    .RESET_B(net884),
    .D(_0186_),
    .Q_N(_1507_),
    .Q(\fifo_d[4][7] ));
 sg13g2_dfrbp_1 _2927_ (.CLK(net826),
    .RESET_B(net891),
    .D(_0187_),
    .Q_N(_1506_),
    .Q(\fifo_d[5][0] ));
 sg13g2_dfrbp_1 _2928_ (.CLK(net837),
    .RESET_B(net908),
    .D(_0188_),
    .Q_N(_1505_),
    .Q(\fifo_d[5][1] ));
 sg13g2_dfrbp_1 _2929_ (.CLK(net837),
    .RESET_B(net911),
    .D(_0189_),
    .Q_N(_1504_),
    .Q(\fifo_d[5][2] ));
 sg13g2_dfrbp_1 _2930_ (.CLK(net829),
    .RESET_B(net890),
    .D(_0190_),
    .Q_N(_1503_),
    .Q(\fifo_d[5][3] ));
 sg13g2_dfrbp_1 _2931_ (.CLK(net826),
    .RESET_B(net888),
    .D(_0191_),
    .Q_N(_1502_),
    .Q(\fifo_d[5][4] ));
 sg13g2_dfrbp_1 _2932_ (.CLK(net835),
    .RESET_B(net906),
    .D(_0192_),
    .Q_N(_1501_),
    .Q(\fifo_d[5][5] ));
 sg13g2_dfrbp_1 _2933_ (.CLK(net829),
    .RESET_B(net889),
    .D(_0193_),
    .Q_N(_1500_),
    .Q(\fifo_d[5][6] ));
 sg13g2_dfrbp_1 _2934_ (.CLK(net830),
    .RESET_B(net889),
    .D(_0194_),
    .Q_N(_1499_),
    .Q(\fifo_d[5][7] ));
 sg13g2_dfrbp_1 _2935_ (.CLK(net843),
    .RESET_B(net913),
    .D(_0195_),
    .Q_N(_1498_),
    .Q(\fifo_d[6][0] ));
 sg13g2_dfrbp_1 _2936_ (.CLK(net841),
    .RESET_B(net911),
    .D(_0196_),
    .Q_N(_1497_),
    .Q(\fifo_d[6][1] ));
 sg13g2_dfrbp_1 _2937_ (.CLK(net842),
    .RESET_B(net913),
    .D(_0197_),
    .Q_N(_1496_),
    .Q(\fifo_d[6][2] ));
 sg13g2_dfrbp_1 _2938_ (.CLK(net837),
    .RESET_B(net911),
    .D(_0198_),
    .Q_N(_1495_),
    .Q(\fifo_d[6][3] ));
 sg13g2_dfrbp_1 _2939_ (.CLK(net835),
    .RESET_B(net905),
    .D(_0199_),
    .Q_N(_1494_),
    .Q(\fifo_d[6][4] ));
 sg13g2_dfrbp_1 _2940_ (.CLK(net835),
    .RESET_B(net906),
    .D(_0200_),
    .Q_N(_1493_),
    .Q(\fifo_d[6][5] ));
 sg13g2_dfrbp_1 _2941_ (.CLK(net835),
    .RESET_B(net905),
    .D(_0201_),
    .Q_N(_1492_),
    .Q(\fifo_d[6][6] ));
 sg13g2_dfrbp_1 _2942_ (.CLK(net841),
    .RESET_B(net912),
    .D(_0202_),
    .Q_N(_1491_),
    .Q(\fifo_d[6][7] ));
 sg13g2_dfrbp_1 _2943_ (.CLK(net842),
    .RESET_B(net914),
    .D(_0203_),
    .Q_N(_1490_),
    .Q(\fifo_d[7][0] ));
 sg13g2_dfrbp_1 _2944_ (.CLK(net841),
    .RESET_B(net912),
    .D(_0204_),
    .Q_N(_1489_),
    .Q(\fifo_d[7][1] ));
 sg13g2_dfrbp_1 _2945_ (.CLK(net842),
    .RESET_B(net913),
    .D(_0205_),
    .Q_N(_1488_),
    .Q(\fifo_d[7][2] ));
 sg13g2_dfrbp_1 _2946_ (.CLK(net837),
    .RESET_B(net911),
    .D(_0206_),
    .Q_N(_1487_),
    .Q(\fifo_d[7][3] ));
 sg13g2_dfrbp_1 _2947_ (.CLK(net845),
    .RESET_B(net917),
    .D(_0207_),
    .Q_N(_1486_),
    .Q(\fifo_d[7][4] ));
 sg13g2_dfrbp_1 _2948_ (.CLK(net840),
    .RESET_B(net916),
    .D(_0208_),
    .Q_N(_1485_),
    .Q(\fifo_d[7][5] ));
 sg13g2_dfrbp_1 _2949_ (.CLK(net835),
    .RESET_B(net905),
    .D(_0209_),
    .Q_N(_1484_),
    .Q(\fifo_d[7][6] ));
 sg13g2_dfrbp_1 _2950_ (.CLK(net831),
    .RESET_B(net889),
    .D(_0210_),
    .Q_N(_1483_),
    .Q(\fifo_d[7][7] ));
 sg13g2_dfrbp_1 _2951_ (.CLK(net844),
    .RESET_B(net917),
    .D(_0211_),
    .Q_N(_1482_),
    .Q(\fifo_d[8][0] ));
 sg13g2_dfrbp_1 _2952_ (.CLK(net827),
    .RESET_B(net886),
    .D(_0212_),
    .Q_N(_1481_),
    .Q(\fifo_d[8][1] ));
 sg13g2_dfrbp_1 _2953_ (.CLK(net827),
    .RESET_B(net886),
    .D(_0213_),
    .Q_N(_1480_),
    .Q(\fifo_d[8][2] ));
 sg13g2_dfrbp_1 _2954_ (.CLK(net839),
    .RESET_B(net909),
    .D(_0214_),
    .Q_N(_1479_),
    .Q(\fifo_d[8][3] ));
 sg13g2_dfrbp_1 _2955_ (.CLK(net845),
    .RESET_B(net917),
    .D(_0215_),
    .Q_N(_1478_),
    .Q(\fifo_d[8][4] ));
 sg13g2_dfrbp_1 _2956_ (.CLK(net840),
    .RESET_B(net909),
    .D(_0216_),
    .Q_N(_1477_),
    .Q(\fifo_d[8][5] ));
 sg13g2_dfrbp_1 _2957_ (.CLK(net839),
    .RESET_B(net909),
    .D(_0217_),
    .Q_N(_1476_),
    .Q(\fifo_d[8][6] ));
 sg13g2_dfrbp_1 _2958_ (.CLK(net844),
    .RESET_B(net916),
    .D(_0218_),
    .Q_N(_1475_),
    .Q(\fifo_d[8][7] ));
 sg13g2_dfrbp_1 _2959_ (.CLK(net828),
    .RESET_B(net886),
    .D(_0219_),
    .Q_N(_1474_),
    .Q(\fifo_d[9][0] ));
 sg13g2_dfrbp_1 _2960_ (.CLK(net837),
    .RESET_B(net912),
    .D(_0220_),
    .Q_N(_1473_),
    .Q(\fifo_d[9][1] ));
 sg13g2_dfrbp_1 _2961_ (.CLK(net828),
    .RESET_B(net886),
    .D(_0221_),
    .Q_N(_1472_),
    .Q(\fifo_d[9][2] ));
 sg13g2_dfrbp_1 _2962_ (.CLK(net836),
    .RESET_B(net908),
    .D(_0222_),
    .Q_N(_1471_),
    .Q(\fifo_d[9][3] ));
 sg13g2_dfrbp_1 _2963_ (.CLK(net840),
    .RESET_B(net909),
    .D(_0223_),
    .Q_N(_1470_),
    .Q(\fifo_d[9][4] ));
 sg13g2_dfrbp_1 _2964_ (.CLK(net840),
    .RESET_B(net909),
    .D(_0224_),
    .Q_N(_1469_),
    .Q(\fifo_d[9][5] ));
 sg13g2_dfrbp_1 _2965_ (.CLK(net836),
    .RESET_B(net907),
    .D(_0225_),
    .Q_N(_1468_),
    .Q(\fifo_d[9][6] ));
 sg13g2_dfrbp_1 _2966_ (.CLK(net838),
    .RESET_B(net912),
    .D(_0226_),
    .Q_N(_1467_),
    .Q(\fifo_d[9][7] ));
 sg13g2_dfrbp_1 _2967_ (.CLK(net842),
    .RESET_B(net913),
    .D(_0227_),
    .Q_N(_1466_),
    .Q(\fifo_d[10][0] ));
 sg13g2_dfrbp_1 _2968_ (.CLK(net837),
    .RESET_B(net911),
    .D(_0228_),
    .Q_N(_1465_),
    .Q(\fifo_d[10][1] ));
 sg13g2_dfrbp_1 _2969_ (.CLK(net842),
    .RESET_B(net913),
    .D(_0229_),
    .Q_N(_1464_),
    .Q(\fifo_d[10][2] ));
 sg13g2_dfrbp_1 _2970_ (.CLK(net835),
    .RESET_B(net908),
    .D(_0230_),
    .Q_N(_1463_),
    .Q(\fifo_d[10][3] ));
 sg13g2_dfrbp_1 _2971_ (.CLK(net845),
    .RESET_B(net914),
    .D(_0231_),
    .Q_N(_1462_),
    .Q(\fifo_d[10][4] ));
 sg13g2_dfrbp_1 _2972_ (.CLK(net839),
    .RESET_B(net907),
    .D(_0232_),
    .Q_N(_1461_),
    .Q(\fifo_d[10][5] ));
 sg13g2_dfrbp_1 _2973_ (.CLK(net839),
    .RESET_B(net908),
    .D(_0233_),
    .Q_N(_1460_),
    .Q(\fifo_d[10][6] ));
 sg13g2_dfrbp_1 _2974_ (.CLK(net831),
    .RESET_B(net890),
    .D(_0234_),
    .Q_N(_1459_),
    .Q(\fifo_d[10][7] ));
 sg13g2_dfrbp_1 _2975_ (.CLK(net843),
    .RESET_B(net914),
    .D(_0235_),
    .Q_N(_1458_),
    .Q(\fifo_d[11][0] ));
 sg13g2_dfrbp_1 _2976_ (.CLK(net841),
    .RESET_B(net911),
    .D(_0236_),
    .Q_N(_1457_),
    .Q(\fifo_d[11][1] ));
 sg13g2_dfrbp_1 _2977_ (.CLK(net842),
    .RESET_B(net913),
    .D(_0237_),
    .Q_N(_1456_),
    .Q(\fifo_d[11][2] ));
 sg13g2_dfrbp_1 _2978_ (.CLK(net831),
    .RESET_B(net906),
    .D(_0238_),
    .Q_N(_1455_),
    .Q(\fifo_d[11][3] ));
 sg13g2_dfrbp_1 _2979_ (.CLK(net835),
    .RESET_B(net908),
    .D(_0239_),
    .Q_N(_1454_),
    .Q(\fifo_d[11][4] ));
 sg13g2_dfrbp_1 _2980_ (.CLK(net831),
    .RESET_B(net905),
    .D(_0240_),
    .Q_N(_1453_),
    .Q(\fifo_d[11][5] ));
 sg13g2_dfrbp_1 _2981_ (.CLK(net832),
    .RESET_B(net907),
    .D(_0241_),
    .Q_N(_1452_),
    .Q(\fifo_d[11][6] ));
 sg13g2_dfrbp_1 _2982_ (.CLK(net841),
    .RESET_B(net911),
    .D(_0242_),
    .Q_N(_1451_),
    .Q(\fifo_d[11][7] ));
 sg13g2_dfrbp_1 _2983_ (.CLK(net825),
    .RESET_B(net884),
    .D(_0243_),
    .Q_N(_1450_),
    .Q(\fifo_d[12][0] ));
 sg13g2_dfrbp_1 _2984_ (.CLK(net824),
    .RESET_B(net884),
    .D(_0244_),
    .Q_N(_1449_),
    .Q(\fifo_d[12][1] ));
 sg13g2_dfrbp_1 _2985_ (.CLK(net824),
    .RESET_B(net885),
    .D(_0245_),
    .Q_N(_1448_),
    .Q(\fifo_d[12][2] ));
 sg13g2_dfrbp_1 _2986_ (.CLK(net829),
    .RESET_B(net889),
    .D(_0246_),
    .Q_N(_1447_),
    .Q(\fifo_d[12][3] ));
 sg13g2_dfrbp_1 _2987_ (.CLK(net826),
    .RESET_B(net888),
    .D(_0247_),
    .Q_N(_1446_),
    .Q(\fifo_d[12][4] ));
 sg13g2_dfrbp_1 _2988_ (.CLK(net829),
    .RESET_B(net889),
    .D(_0248_),
    .Q_N(_1445_),
    .Q(\fifo_d[12][5] ));
 sg13g2_dfrbp_1 _2989_ (.CLK(net829),
    .RESET_B(net889),
    .D(_0249_),
    .Q_N(_1444_),
    .Q(\fifo_d[12][6] ));
 sg13g2_dfrbp_1 _2990_ (.CLK(net825),
    .RESET_B(net884),
    .D(_0250_),
    .Q_N(_1443_),
    .Q(\fifo_d[12][7] ));
 sg13g2_dfrbp_1 _2991_ (.CLK(net828),
    .RESET_B(net893),
    .D(_0251_),
    .Q_N(_1442_),
    .Q(\fifo_d[13][0] ));
 sg13g2_dfrbp_1 _2992_ (.CLK(net828),
    .RESET_B(net893),
    .D(_0252_),
    .Q_N(_1441_),
    .Q(\fifo_d[13][1] ));
 sg13g2_dfrbp_1 _2993_ (.CLK(net828),
    .RESET_B(net888),
    .D(_0253_),
    .Q_N(_1440_),
    .Q(\fifo_d[13][2] ));
 sg13g2_dfrbp_1 _2994_ (.CLK(net833),
    .RESET_B(net890),
    .D(_0254_),
    .Q_N(_1439_),
    .Q(\fifo_d[13][3] ));
 sg13g2_dfrbp_1 _2995_ (.CLK(net833),
    .RESET_B(net892),
    .D(_0255_),
    .Q_N(_1438_),
    .Q(\fifo_d[13][4] ));
 sg13g2_dfrbp_1 _2996_ (.CLK(net830),
    .RESET_B(net891),
    .D(_0256_),
    .Q_N(_1437_),
    .Q(\fifo_d[13][5] ));
 sg13g2_dfrbp_1 _2997_ (.CLK(net831),
    .RESET_B(net890),
    .D(_0257_),
    .Q_N(_1436_),
    .Q(\fifo_d[13][6] ));
 sg13g2_dfrbp_1 _2998_ (.CLK(net830),
    .RESET_B(net890),
    .D(_0258_),
    .Q_N(_1435_),
    .Q(\fifo_d[13][7] ));
 sg13g2_dfrbp_1 _2999_ (.CLK(net824),
    .RESET_B(net887),
    .D(_0259_),
    .Q_N(_1434_),
    .Q(\fifo_d[14][0] ));
 sg13g2_dfrbp_1 _3000_ (.CLK(net827),
    .RESET_B(net886),
    .D(_0260_),
    .Q_N(_1433_),
    .Q(\fifo_d[14][1] ));
 sg13g2_dfrbp_1 _3001_ (.CLK(net827),
    .RESET_B(net886),
    .D(_0261_),
    .Q_N(_1432_),
    .Q(\fifo_d[14][2] ));
 sg13g2_dfrbp_1 _3002_ (.CLK(net830),
    .RESET_B(net890),
    .D(_0262_),
    .Q_N(_1431_),
    .Q(\fifo_d[14][3] ));
 sg13g2_dfrbp_1 _3003_ (.CLK(net826),
    .RESET_B(net888),
    .D(_0263_),
    .Q_N(_1430_),
    .Q(\fifo_d[14][4] ));
 sg13g2_dfrbp_1 _3004_ (.CLK(net833),
    .RESET_B(net892),
    .D(_0264_),
    .Q_N(_1429_),
    .Q(\fifo_d[14][5] ));
 sg13g2_dfrbp_1 _3005_ (.CLK(net825),
    .RESET_B(net884),
    .D(_0265_),
    .Q_N(_1428_),
    .Q(\fifo_d[14][6] ));
 sg13g2_dfrbp_1 _3006_ (.CLK(net829),
    .RESET_B(net889),
    .D(_0266_),
    .Q_N(_1427_),
    .Q(\fifo_d[14][7] ));
 sg13g2_dfrbp_1 _3007_ (.CLK(net842),
    .RESET_B(net914),
    .D(_0267_),
    .Q_N(_1426_),
    .Q(\fifo_d[15][0] ));
 sg13g2_dfrbp_1 _3008_ (.CLK(net828),
    .RESET_B(net893),
    .D(_0268_),
    .Q_N(_1425_),
    .Q(\fifo_d[15][1] ));
 sg13g2_dfrbp_1 _3009_ (.CLK(net842),
    .RESET_B(net913),
    .D(_0269_),
    .Q_N(_1424_),
    .Q(\fifo_d[15][2] ));
 sg13g2_dfrbp_1 _3010_ (.CLK(net836),
    .RESET_B(net908),
    .D(_0270_),
    .Q_N(_1423_),
    .Q(\fifo_d[15][3] ));
 sg13g2_dfrbp_1 _3011_ (.CLK(net844),
    .RESET_B(net913),
    .D(_0271_),
    .Q_N(_1422_),
    .Q(\fifo_d[15][4] ));
 sg13g2_dfrbp_1 _3012_ (.CLK(net840),
    .RESET_B(net916),
    .D(_0272_),
    .Q_N(_1421_),
    .Q(\fifo_d[15][5] ));
 sg13g2_dfrbp_1 _3013_ (.CLK(net836),
    .RESET_B(net905),
    .D(_0273_),
    .Q_N(_1420_),
    .Q(\fifo_d[15][6] ));
 sg13g2_dfrbp_1 _3014_ (.CLK(net841),
    .RESET_B(net912),
    .D(_0274_),
    .Q_N(_1562_),
    .Q(\fifo_d[15][7] ));
 sg13g2_dfrbp_1 _3015_ (.CLK(clknet_1_0__leaf_clk),
    .RESET_B(net928),
    .D(net27),
    .Q_N(_1563_),
    .Q(\clk_out_cnt[0] ));
 sg13g2_dfrbp_1 _3016_ (.CLK(clknet_1_0__leaf_clk),
    .RESET_B(net928),
    .D(_0001_),
    .Q_N(_1564_),
    .Q(\clk_out_cnt[1] ));
 sg13g2_dfrbp_1 _3017_ (.CLK(clknet_1_1__leaf_clk),
    .RESET_B(net928),
    .D(_0002_),
    .Q_N(_1565_),
    .Q(\clk_out_cnt[2] ));
 sg13g2_dfrbp_1 _3018_ (.CLK(clknet_1_1__leaf_clk),
    .RESET_B(net928),
    .D(net25),
    .Q_N(_1419_),
    .Q(\clk_out_cnt[3] ));
 sg13g2_dfrbp_1 _3019_ (.CLK(net882),
    .RESET_B(net927),
    .D(_0275_),
    .Q_N(\uart_0.rx.rx_sample_wrap[0] ),
    .Q(_0041_));
 sg13g2_dfrbp_1 _3020_ (.CLK(net882),
    .RESET_B(net927),
    .D(_0276_),
    .Q_N(_1418_),
    .Q(\uart_0.rx.rx_sample_wrap[3] ));
 sg13g2_dfrbp_1 _3021_ (.CLK(net878),
    .RESET_B(net924),
    .D(_0277_),
    .Q_N(_0037_),
    .Q(\uart_0.tx.tx_bit_cnt[0] ));
 sg13g2_dfrbp_1 _3022_ (.CLK(net878),
    .RESET_B(net924),
    .D(_0278_),
    .Q_N(_1417_),
    .Q(\uart_0.tx.tx_bit_cnt[1] ));
 sg13g2_dfrbp_1 _3023_ (.CLK(net878),
    .RESET_B(net924),
    .D(_0279_),
    .Q_N(_0036_),
    .Q(\uart_0.tx.tx_bit_cnt[2] ));
 sg13g2_dfrbp_1 _3024_ (.CLK(net878),
    .RESET_B(net924),
    .D(_0280_),
    .Q_N(_0035_),
    .Q(\uart_0.tx.tx_bit_cnt[3] ));
 sg13g2_dfrbp_1 _3025_ (.CLK(net874),
    .RESET_B(net923),
    .D(_0281_),
    .Q_N(_1416_),
    .Q(\uart_0.rx.rx_stop_zeros[0] ));
 sg13g2_dfrbp_1 _3026_ (.CLK(net874),
    .RESET_B(net923),
    .D(_0282_),
    .Q_N(_1415_),
    .Q(\uart_0.rx.rx_stop_zeros[1] ));
 sg13g2_dfrbp_1 _3027_ (.CLK(net866),
    .RESET_B(net901),
    .D(_0283_),
    .Q_N(_0028_),
    .Q(\uart_0.rx.rx_stop_zeros[2] ));
 sg13g2_dfrbp_1 _3028_ (.CLK(net874),
    .RESET_B(net923),
    .D(_0284_),
    .Q_N(_1414_),
    .Q(\uart_0.rx.rx_stop_zeros[3] ));
 sg13g2_dfrbp_1 _3029_ (.CLK(net874),
    .RESET_B(net923),
    .D(_0285_),
    .Q_N(_0030_),
    .Q(\uart_0.rx.rx_stop_zeros[4] ));
 sg13g2_dfrbp_1 _3030_ (.CLK(net874),
    .RESET_B(net923),
    .D(_0286_),
    .Q_N(_0029_),
    .Q(\uart_0.rx.rx_stop_zeros[5] ));
 sg13g2_dfrbp_1 _3031_ (.CLK(net874),
    .RESET_B(net923),
    .D(_0287_),
    .Q_N(_0031_),
    .Q(\uart_0.rx.rx_stop_zeros[6] ));
 sg13g2_dfrbp_1 _3032_ (.CLK(net878),
    .RESET_B(net925),
    .D(_0020_),
    .Q_N(_1566_),
    .Q(\uart_0.tx.tx_baudrate_cnt[0] ));
 sg13g2_dfrbp_1 _3033_ (.CLK(net877),
    .RESET_B(net925),
    .D(_0021_),
    .Q_N(_1567_),
    .Q(\uart_0.tx.tx_baudrate_cnt[1] ));
 sg13g2_dfrbp_1 _3034_ (.CLK(net878),
    .RESET_B(net925),
    .D(_0022_),
    .Q_N(_1568_),
    .Q(\uart_0.tx.tx_baudrate_cnt[2] ));
 sg13g2_dfrbp_1 _3035_ (.CLK(net881),
    .RESET_B(net925),
    .D(_0023_),
    .Q_N(_1569_),
    .Q(\uart_0.tx.tx_baudrate_cnt[3] ));
 sg13g2_dfrbp_1 _3036_ (.CLK(net879),
    .RESET_B(net924),
    .D(_0024_),
    .Q_N(_1570_),
    .Q(\uart_0.tx.tx_baudrate_cnt[4] ));
 sg13g2_dfrbp_1 _3037_ (.CLK(net879),
    .RESET_B(net924),
    .D(_0025_),
    .Q_N(_1571_),
    .Q(\uart_0.tx.tx_baudrate_cnt[5] ));
 sg13g2_dfrbp_1 _3038_ (.CLK(net878),
    .RESET_B(net924),
    .D(_0026_),
    .Q_N(_1572_),
    .Q(\uart_0.tx.tx_baudrate_cnt[6] ));
 sg13g2_dfrbp_1 _3039_ (.CLK(net878),
    .RESET_B(net924),
    .D(_0027_),
    .Q_N(_1413_),
    .Q(\uart_0.tx.tx_baudrate_cnt[7] ));
 sg13g2_dfrbp_1 _3040_ (.CLK(net873),
    .RESET_B(net922),
    .D(_0288_),
    .Q_N(_1412_),
    .Q(\uart_0.rx.rx_marker[0] ));
 sg13g2_dfrbp_1 _3041_ (.CLK(net873),
    .RESET_B(net923),
    .D(_0289_),
    .Q_N(\uart_0.rx.rx_marker[1] ),
    .Q(_0042_));
 sg13g2_dfrbp_1 _3042_ (.CLK(net872),
    .RESET_B(net922),
    .D(_0290_),
    .Q_N(_1411_),
    .Q(\uart_0.rx.rx_marker[2] ));
 sg13g2_dfrbp_1 _3043_ (.CLK(net872),
    .RESET_B(net922),
    .D(_0291_),
    .Q_N(\uart_0.rx.rx_marker[3] ),
    .Q(_0043_));
 sg13g2_dfrbp_1 _3044_ (.CLK(net872),
    .RESET_B(net922),
    .D(_0292_),
    .Q_N(\uart_0.rx.rx_marker[4] ),
    .Q(_0044_));
 sg13g2_dfrbp_1 _3045_ (.CLK(net873),
    .RESET_B(net922),
    .D(_0293_),
    .Q_N(_0033_),
    .Q(\uart_0.rx.rx_marker[5] ));
 sg13g2_dfrbp_1 _3046_ (.CLK(net873),
    .RESET_B(net922),
    .D(_0294_),
    .Q_N(\uart_0.rx.rx_marker[6] ),
    .Q(_0045_));
 sg13g2_dfrbp_1 _3047_ (.CLK(net879),
    .RESET_B(net917),
    .D(_0295_),
    .Q_N(_1410_),
    .Q(\uart_0.tx.tx_data_tmp[2] ));
 sg13g2_dfrbp_1 _3048_ (.CLK(net879),
    .RESET_B(net917),
    .D(_0296_),
    .Q_N(_1409_),
    .Q(\uart_0.tx.tx_data_tmp[3] ));
 sg13g2_dfrbp_1 _3049_ (.CLK(net876),
    .RESET_B(net916),
    .D(_0297_),
    .Q_N(_1408_),
    .Q(\uart_0.tx.tx_data_tmp[4] ));
 sg13g2_dfrbp_1 _3050_ (.CLK(net876),
    .RESET_B(net916),
    .D(_0298_),
    .Q_N(_1407_),
    .Q(\uart_0.tx.tx_data_tmp[5] ));
 sg13g2_dfrbp_1 _3051_ (.CLK(net876),
    .RESET_B(net916),
    .D(_0299_),
    .Q_N(_1406_),
    .Q(\uart_0.tx.tx_data_tmp[6] ));
 sg13g2_dfrbp_1 _3052_ (.CLK(net876),
    .RESET_B(net926),
    .D(_0300_),
    .Q_N(_1405_),
    .Q(\uart_0.tx.tx_data_tmp[7] ));
 sg13g2_dfrbp_1 _3053_ (.CLK(net876),
    .RESET_B(net926),
    .D(_0301_),
    .Q_N(_1404_),
    .Q(\uart_0.tx.tx_data_tmp[8] ));
 sg13g2_dfrbp_1 _3054_ (.CLK(net876),
    .RESET_B(net926),
    .D(_0302_),
    .Q_N(_1403_),
    .Q(\uart_0.tx.tx_data_tmp[9] ));
 sg13g2_dfrbp_1 _3055_ (.CLK(net867),
    .RESET_B(net902),
    .D(_0303_),
    .Q_N(\uart_0.rx.rx_samples[0] ),
    .Q(_0046_));
 sg13g2_dfrbp_1 _3056_ (.CLK(net861),
    .RESET_B(net898),
    .D(_0304_),
    .Q_N(\uart_0.rx.rx_samples[1] ),
    .Q(_0047_));
 sg13g2_dfrbp_1 _3057_ (.CLK(net861),
    .RESET_B(net898),
    .D(_0305_),
    .Q_N(\uart_0.rx.rx_samples[2] ),
    .Q(_0048_));
 sg13g2_dfrbp_1 _3058_ (.CLK(net867),
    .RESET_B(net902),
    .D(_0306_),
    .Q_N(\uart_0.rx.rx_samples[3] ),
    .Q(_0049_));
 sg13g2_dfrbp_1 _3059_ (.CLK(net867),
    .RESET_B(net902),
    .D(_0307_),
    .Q_N(\uart_0.rx.rx_samples[4] ),
    .Q(_0050_));
 sg13g2_dfrbp_1 _3060_ (.CLK(net867),
    .RESET_B(net902),
    .D(_0308_),
    .Q_N(\uart_0.rx.rx_samples[5] ),
    .Q(_0051_));
 sg13g2_dfrbp_1 _3061_ (.CLK(net862),
    .RESET_B(net898),
    .D(_0309_),
    .Q_N(\uart_0.rx.rx_samples[6] ),
    .Q(_0052_));
 sg13g2_dfrbp_1 _3062_ (.CLK(net861),
    .RESET_B(net899),
    .D(_0310_),
    .Q_N(\uart_0.rx.rx_samples[7] ),
    .Q(_0053_));
 sg13g2_dfrbp_1 _3063_ (.CLK(net861),
    .RESET_B(net898),
    .D(_0311_),
    .Q_N(\uart_0.rx.rx_samples[8] ),
    .Q(_0054_));
 sg13g2_dfrbp_1 _3064_ (.CLK(net859),
    .RESET_B(net897),
    .D(_0312_),
    .Q_N(\uart_0.rx.rx_samples[9] ),
    .Q(_0055_));
 sg13g2_dfrbp_1 _3065_ (.CLK(net859),
    .RESET_B(net897),
    .D(_0313_),
    .Q_N(\uart_0.rx.rx_samples[10] ),
    .Q(_0056_));
 sg13g2_dfrbp_1 _3066_ (.CLK(net860),
    .RESET_B(net897),
    .D(_0314_),
    .Q_N(\uart_0.rx.rx_samples[11] ),
    .Q(_0057_));
 sg13g2_dfrbp_1 _3067_ (.CLK(net859),
    .RESET_B(net897),
    .D(_0315_),
    .Q_N(\uart_0.rx.rx_samples[12] ),
    .Q(_0058_));
 sg13g2_dfrbp_1 _3068_ (.CLK(net859),
    .RESET_B(net897),
    .D(_0316_),
    .Q_N(\uart_0.rx.rx_samples[13] ),
    .Q(_0059_));
 sg13g2_dfrbp_1 _3069_ (.CLK(net860),
    .RESET_B(net899),
    .D(_0317_),
    .Q_N(\uart_0.rx.rx_samples[14] ),
    .Q(_0060_));
 sg13g2_dfrbp_1 _3070_ (.CLK(net860),
    .RESET_B(net897),
    .D(_0318_),
    .Q_N(\uart_0.rx.rx_samples[15] ),
    .Q(_0061_));
 sg13g2_dfrbp_1 _3071_ (.CLK(net860),
    .RESET_B(net899),
    .D(_0319_),
    .Q_N(\uart_0.rx.rx_samples[16] ),
    .Q(_0062_));
 sg13g2_dfrbp_1 _3072_ (.CLK(net867),
    .RESET_B(net902),
    .D(_0320_),
    .Q_N(\uart_0.rx.rx_samples[17] ),
    .Q(_0063_));
 sg13g2_dfrbp_1 _3073_ (.CLK(net867),
    .RESET_B(net902),
    .D(_0321_),
    .Q_N(\uart_0.rx.rx_samples[18] ),
    .Q(_0064_));
 sg13g2_dfrbp_1 _3074_ (.CLK(net866),
    .RESET_B(net901),
    .D(_0322_),
    .Q_N(\uart_0.rx.rx_samples[19] ),
    .Q(_0065_));
 sg13g2_dfrbp_1 _3075_ (.CLK(net866),
    .RESET_B(net901),
    .D(_0323_),
    .Q_N(\uart_0.rx.rx_samples[20] ),
    .Q(_0066_));
 sg13g2_dfrbp_1 _3076_ (.CLK(net866),
    .RESET_B(net901),
    .D(_0324_),
    .Q_N(\uart_0.rx.rx_samples[21] ),
    .Q(_0067_));
 sg13g2_dfrbp_1 _3077_ (.CLK(net866),
    .RESET_B(net901),
    .D(_0325_),
    .Q_N(\uart_0.rx.rx_samples[22] ),
    .Q(_0068_));
 sg13g2_dfrbp_1 _3078_ (.CLK(net866),
    .RESET_B(net901),
    .D(_0326_),
    .Q_N(\uart_0.rx.rx_samples[23] ),
    .Q(_0069_));
 sg13g2_dfrbp_1 _3079_ (.CLK(net866),
    .RESET_B(net902),
    .D(_0327_),
    .Q_N(\uart_0.rx.rx_samples[24] ),
    .Q(_0070_));
 sg13g2_dfrbp_1 _3080_ (.CLK(net866),
    .RESET_B(net901),
    .D(_0328_),
    .Q_N(\uart_0.rx.rx_samples[25] ),
    .Q(_0071_));
 sg13g2_dfrbp_1 _3081_ (.CLK(net867),
    .RESET_B(net901),
    .D(_0329_),
    .Q_N(\uart_0.rx.rx_samples[26] ),
    .Q(_0072_));
 sg13g2_dfrbp_1 _3082_ (.CLK(net862),
    .RESET_B(net898),
    .D(_0330_),
    .Q_N(\uart_0.rx.rx_samples[27] ),
    .Q(_0073_));
 sg13g2_dfrbp_1 _3083_ (.CLK(net862),
    .RESET_B(net898),
    .D(_0331_),
    .Q_N(\uart_0.rx.rx_samples[28] ),
    .Q(_0074_));
 sg13g2_dfrbp_1 _3084_ (.CLK(net861),
    .RESET_B(net898),
    .D(_0332_),
    .Q_N(\uart_0.rx.rx_samples[29] ),
    .Q(_0075_));
 sg13g2_dfrbp_1 _3085_ (.CLK(net861),
    .RESET_B(net898),
    .D(_0333_),
    .Q_N(\uart_0.rx.rx_samples[30] ),
    .Q(_0076_));
 sg13g2_dfrbp_1 _3086_ (.CLK(net860),
    .RESET_B(net897),
    .D(_0334_),
    .Q_N(\uart_0.rx.rx_samples[31] ),
    .Q(_0077_));
 sg13g2_dfrbp_1 _3087_ (.CLK(net860),
    .RESET_B(net896),
    .D(_0335_),
    .Q_N(\uart_0.rx.rx_samples[32] ),
    .Q(_0078_));
 sg13g2_dfrbp_1 _3088_ (.CLK(net859),
    .RESET_B(net897),
    .D(_0336_),
    .Q_N(\uart_0.rx.rx_samples[33] ),
    .Q(_0079_));
 sg13g2_dfrbp_1 _3089_ (.CLK(net861),
    .RESET_B(net896),
    .D(_0337_),
    .Q_N(\uart_0.rx.rx_samples[34] ),
    .Q(_0080_));
 sg13g2_dfrbp_1 _3090_ (.CLK(net861),
    .RESET_B(net895),
    .D(_0338_),
    .Q_N(\uart_0.rx.rx_samples[35] ),
    .Q(_0081_));
 sg13g2_dfrbp_1 _3091_ (.CLK(net863),
    .RESET_B(net895),
    .D(_0339_),
    .Q_N(\uart_0.rx.rx_samples[36] ),
    .Q(_0082_));
 sg13g2_dfrbp_1 _3092_ (.CLK(net864),
    .RESET_B(net900),
    .D(_0340_),
    .Q_N(\uart_0.rx.rx_samples[37] ),
    .Q(_0083_));
 sg13g2_dfrbp_1 _3093_ (.CLK(net864),
    .RESET_B(net900),
    .D(_0341_),
    .Q_N(\uart_0.rx.rx_samples[38] ),
    .Q(_0084_));
 sg13g2_dfrbp_1 _3094_ (.CLK(net864),
    .RESET_B(net900),
    .D(_0342_),
    .Q_N(\uart_0.rx.rx_samples[39] ),
    .Q(_0085_));
 sg13g2_dfrbp_1 _3095_ (.CLK(net864),
    .RESET_B(net900),
    .D(_0343_),
    .Q_N(\uart_0.rx.rx_samples[40] ),
    .Q(_0086_));
 sg13g2_dfrbp_1 _3096_ (.CLK(net864),
    .RESET_B(net900),
    .D(_0344_),
    .Q_N(\uart_0.rx.rx_samples[41] ),
    .Q(_0087_));
 sg13g2_dfrbp_1 _3097_ (.CLK(net864),
    .RESET_B(net900),
    .D(_0345_),
    .Q_N(\uart_0.rx.rx_samples[42] ),
    .Q(_0088_));
 sg13g2_dfrbp_1 _3098_ (.CLK(net864),
    .RESET_B(net900),
    .D(_0346_),
    .Q_N(\uart_0.rx.rx_samples[43] ),
    .Q(_0089_));
 sg13g2_dfrbp_1 _3099_ (.CLK(net863),
    .RESET_B(net896),
    .D(_0347_),
    .Q_N(\uart_0.rx.rx_samples[44] ),
    .Q(_0090_));
 sg13g2_dfrbp_1 _3100_ (.CLK(net857),
    .RESET_B(net895),
    .D(_0348_),
    .Q_N(\uart_0.rx.rx_samples[45] ),
    .Q(_0091_));
 sg13g2_dfrbp_1 _3101_ (.CLK(net857),
    .RESET_B(net895),
    .D(_0349_),
    .Q_N(\uart_0.rx.rx_samples[46] ),
    .Q(_0092_));
 sg13g2_dfrbp_1 _3102_ (.CLK(net857),
    .RESET_B(net895),
    .D(_0350_),
    .Q_N(\uart_0.rx.rx_samples[47] ),
    .Q(_0093_));
 sg13g2_dfrbp_1 _3103_ (.CLK(net857),
    .RESET_B(net895),
    .D(_0351_),
    .Q_N(\uart_0.rx.rx_samples[48] ),
    .Q(_0094_));
 sg13g2_dfrbp_1 _3104_ (.CLK(net857),
    .RESET_B(net887),
    .D(_0352_),
    .Q_N(\uart_0.rx.rx_samples[49] ),
    .Q(_0095_));
 sg13g2_dfrbp_1 _3105_ (.CLK(net857),
    .RESET_B(net895),
    .D(_0353_),
    .Q_N(\uart_0.rx.rx_samples[50] ),
    .Q(_0096_));
 sg13g2_dfrbp_1 _3106_ (.CLK(net857),
    .RESET_B(net895),
    .D(_0354_),
    .Q_N(\uart_0.rx.rx_samples[51] ),
    .Q(_0097_));
 sg13g2_dfrbp_1 _3107_ (.CLK(net857),
    .RESET_B(net887),
    .D(_0355_),
    .Q_N(\uart_0.rx.rx_samples[52] ),
    .Q(_0098_));
 sg13g2_dfrbp_1 _3108_ (.CLK(net858),
    .RESET_B(net894),
    .D(_0356_),
    .Q_N(\uart_0.rx.rx_samples[53] ),
    .Q(_0099_));
 sg13g2_dfrbp_1 _3109_ (.CLK(net858),
    .RESET_B(net894),
    .D(_0357_),
    .Q_N(\uart_0.rx.rx_samples[54] ),
    .Q(_0100_));
 sg13g2_dfrbp_1 _3110_ (.CLK(net858),
    .RESET_B(net894),
    .D(_0358_),
    .Q_N(\uart_0.rx.rx_samples[55] ),
    .Q(_0101_));
 sg13g2_dfrbp_1 _3111_ (.CLK(net858),
    .RESET_B(net894),
    .D(_0359_),
    .Q_N(\uart_0.rx.rx_samples[56] ),
    .Q(_0102_));
 sg13g2_dfrbp_1 _3112_ (.CLK(net859),
    .RESET_B(net896),
    .D(_0360_),
    .Q_N(\uart_0.rx.rx_samples[57] ),
    .Q(_0103_));
 sg13g2_dfrbp_1 _3113_ (.CLK(net859),
    .RESET_B(net896),
    .D(_0361_),
    .Q_N(\uart_0.rx.rx_samples[58] ),
    .Q(_0104_));
 sg13g2_dfrbp_1 _3114_ (.CLK(net858),
    .RESET_B(net894),
    .D(_0362_),
    .Q_N(\uart_0.rx.rx_samples[59] ),
    .Q(_0105_));
 sg13g2_dfrbp_1 _3115_ (.CLK(net859),
    .RESET_B(net894),
    .D(_0363_),
    .Q_N(\uart_0.rx.rx_samples[60] ),
    .Q(_0106_));
 sg13g2_dfrbp_1 _3116_ (.CLK(net858),
    .RESET_B(net894),
    .D(_0364_),
    .Q_N(\uart_0.rx.rx_samples[61] ),
    .Q(_0107_));
 sg13g2_dfrbp_1 _3117_ (.CLK(net858),
    .RESET_B(net894),
    .D(_0365_),
    .Q_N(\uart_0.rx.rx_samples[62] ),
    .Q(_0108_));
 sg13g2_dfrbp_1 _3118_ (.CLK(net864),
    .RESET_B(net900),
    .D(_0366_),
    .Q_N(\uart_0.rx.rx_samples[63] ),
    .Q(_0109_));
 sg13g2_dfrbp_1 _3119_ (.CLK(net865),
    .RESET_B(net903),
    .D(_0367_),
    .Q_N(\uart_0.rx.rx_samples[64] ),
    .Q(_0110_));
 sg13g2_dfrbp_1 _3120_ (.CLK(net865),
    .RESET_B(net892),
    .D(_0368_),
    .Q_N(\uart_0.rx.rx_samples[65] ),
    .Q(_0111_));
 sg13g2_dfrbp_1 _3121_ (.CLK(net865),
    .RESET_B(net903),
    .D(_0369_),
    .Q_N(\uart_0.rx.rx_samples[66] ),
    .Q(_0112_));
 sg13g2_dfrbp_1 _3122_ (.CLK(net865),
    .RESET_B(net903),
    .D(_0370_),
    .Q_N(\uart_0.rx.rx_samples[67] ),
    .Q(_0113_));
 sg13g2_dfrbp_1 _3123_ (.CLK(net869),
    .RESET_B(net920),
    .D(_0371_),
    .Q_N(\uart_0.rx.rx_samples[68] ),
    .Q(_0114_));
 sg13g2_dfrbp_1 _3124_ (.CLK(net865),
    .RESET_B(net892),
    .D(_0372_),
    .Q_N(\uart_0.rx.rx_samples[69] ),
    .Q(_0115_));
 sg13g2_dfrbp_1 _3125_ (.CLK(net865),
    .RESET_B(net892),
    .D(_0373_),
    .Q_N(\uart_0.rx.rx_samples[70] ),
    .Q(_0116_));
 sg13g2_dfrbp_1 _3126_ (.CLK(net865),
    .RESET_B(net892),
    .D(_0374_),
    .Q_N(\uart_0.rx.rx_samples[71] ),
    .Q(_0117_));
 sg13g2_dfrbp_1 _3127_ (.CLK(net869),
    .RESET_B(net920),
    .D(_0375_),
    .Q_N(\uart_0.rx.rx_samples[72] ),
    .Q(_0118_));
 sg13g2_dfrbp_1 _3128_ (.CLK(net869),
    .RESET_B(net920),
    .D(_0376_),
    .Q_N(\uart_0.rx.rx_samples[73] ),
    .Q(_0119_));
 sg13g2_dfrbp_1 _3129_ (.CLK(net870),
    .RESET_B(net921),
    .D(_0377_),
    .Q_N(\uart_0.rx.rx_samples[74] ),
    .Q(_0120_));
 sg13g2_dfrbp_1 _3130_ (.CLK(net870),
    .RESET_B(net920),
    .D(_0378_),
    .Q_N(\uart_0.rx.rx_samples[75] ),
    .Q(_0121_));
 sg13g2_dfrbp_1 _3131_ (.CLK(net871),
    .RESET_B(net921),
    .D(_0379_),
    .Q_N(\uart_0.rx.rx_samples[76] ),
    .Q(_0122_));
 sg13g2_dfrbp_1 _3132_ (.CLK(net871),
    .RESET_B(net921),
    .D(_0380_),
    .Q_N(\uart_0.rx.rx_samples[77] ),
    .Q(_0123_));
 sg13g2_dfrbp_1 _3133_ (.CLK(net870),
    .RESET_B(net920),
    .D(_0381_),
    .Q_N(\uart_0.rx.rx_samples[78] ),
    .Q(_0124_));
 sg13g2_dfrbp_1 _3134_ (.CLK(net869),
    .RESET_B(net920),
    .D(_0382_),
    .Q_N(\uart_0.rx.rx_samples[79] ),
    .Q(_0125_));
 sg13g2_dfrbp_1 _3135_ (.CLK(net870),
    .RESET_B(net921),
    .D(_0383_),
    .Q_N(\uart_0.rx.rx_samples[80] ),
    .Q(_0126_));
 sg13g2_dfrbp_1 _3136_ (.CLK(net874),
    .RESET_B(net920),
    .D(_0384_),
    .Q_N(\uart_0.rx.rx_samples[81] ),
    .Q(_0127_));
 sg13g2_dfrbp_1 _3137_ (.CLK(net874),
    .RESET_B(net920),
    .D(_0385_),
    .Q_N(\uart_0.rx.rx_samples[82] ),
    .Q(_0128_));
 sg13g2_dfrbp_1 _3138_ (.CLK(net872),
    .RESET_B(net921),
    .D(_0386_),
    .Q_N(\uart_0.rx.rx_samples[83] ),
    .Q(_0129_));
 sg13g2_dfrbp_1 _3139_ (.CLK(net870),
    .RESET_B(net921),
    .D(_0387_),
    .Q_N(\uart_0.rx.rx_samples[84] ),
    .Q(_0130_));
 sg13g2_dfrbp_1 _3140_ (.CLK(net870),
    .RESET_B(net921),
    .D(_0388_),
    .Q_N(\uart_0.rx.rx_samples[85] ),
    .Q(_0131_));
 sg13g2_dfrbp_1 _3141_ (.CLK(net872),
    .RESET_B(net922),
    .D(_0389_),
    .Q_N(\uart_0.rx.rx_samples[86] ),
    .Q(_0132_));
 sg13g2_dfrbp_1 _3142_ (.CLK(net872),
    .RESET_B(net922),
    .D(_0390_),
    .Q_N(\uart_0.rx.rx_samples[87] ),
    .Q(_0133_));
 sg13g2_dfrbp_1 _3143_ (.CLK(net872),
    .RESET_B(net926),
    .D(_0391_),
    .Q_N(\uart_0.rx.rx_samples[88] ),
    .Q(_0134_));
 sg13g2_dfrbp_1 _3144_ (.CLK(net880),
    .RESET_B(net926),
    .D(_0392_),
    .Q_N(\uart_0.rx.rx_samples[89] ),
    .Q(_0135_));
 sg13g2_dfrbp_1 _3145_ (.CLK(net881),
    .RESET_B(net929),
    .D(_0393_),
    .Q_N(_1402_),
    .Q(\uart_0.rx.rx_sample_cnt[0] ));
 sg13g2_dfrbp_1 _3146_ (.CLK(net881),
    .RESET_B(net927),
    .D(_0394_),
    .Q_N(_1401_),
    .Q(\uart_0.rx.rx_sample_cnt[1] ));
 sg13g2_dfrbp_1 _3147_ (.CLK(net881),
    .RESET_B(net927),
    .D(_0395_),
    .Q_N(_1400_),
    .Q(\uart_0.rx.rx_sample_cnt[2] ));
 sg13g2_dfrbp_1 _3148_ (.CLK(net881),
    .RESET_B(net927),
    .D(_0396_),
    .Q_N(_1399_),
    .Q(\uart_0.rx.rx_sample_cnt[3] ));
 sg13g2_dfrbp_1 _3149_ (.CLK(net880),
    .RESET_B(net929),
    .D(_0397_),
    .Q_N(_1398_),
    .Q(\uart_0.rx.rx_sample_cnt[4] ));
 sg13g2_dfrbp_1 _3150_ (.CLK(net882),
    .RESET_B(net929),
    .D(_0398_),
    .Q_N(_1397_),
    .Q(\uart_0.rx.rx_sample_cnt[5] ));
 sg13g2_dfrbp_1 _3151_ (.CLK(net882),
    .RESET_B(net929),
    .D(_0399_),
    .Q_N(_0034_),
    .Q(\uart_0.rx.rx_sample_cnt[6] ));
 sg13g2_dfrbp_1 _3152_ (.CLK(net880),
    .RESET_B(net929),
    .D(_0013_),
    .Q_N(_1573_),
    .Q(\uart_0.rx.rx_sample_clk_cnt[0] ));
 sg13g2_dfrbp_1 _3153_ (.CLK(net880),
    .RESET_B(net927),
    .D(_0014_),
    .Q_N(_1574_),
    .Q(\uart_0.rx.rx_sample_clk_cnt[1] ));
 sg13g2_dfrbp_1 _3154_ (.CLK(net880),
    .RESET_B(net927),
    .D(_0015_),
    .Q_N(_1575_),
    .Q(\uart_0.rx.rx_sample_clk_cnt[2] ));
 sg13g2_dfrbp_1 _3155_ (.CLK(net880),
    .RESET_B(net928),
    .D(_0016_),
    .Q_N(_1576_),
    .Q(\uart_0.rx.rx_sample_clk_cnt[3] ));
 sg13g2_dfrbp_1 _3156_ (.CLK(net880),
    .RESET_B(net928),
    .D(_0017_),
    .Q_N(_1577_),
    .Q(\uart_0.rx.rx_sample_clk_cnt[4] ));
 sg13g2_dfrbp_1 _3157_ (.CLK(net881),
    .RESET_B(net928),
    .D(_0018_),
    .Q_N(_1578_),
    .Q(\uart_0.rx.rx_sample_clk_cnt[5] ));
 sg13g2_dfrbp_1 _3158_ (.CLK(net881),
    .RESET_B(net928),
    .D(_0019_),
    .Q_N(_1396_),
    .Q(\uart_0.rx.rx_sample_clk_cnt[6] ));
 sg13g2_dfrbp_1 _3159_ (.CLK(net872),
    .RESET_B(net929),
    .D(_0400_),
    .Q_N(_0032_),
    .Q(rx_sample_clk));
 sg13g2_dfrbp_1 _3160_ (.CLK(net880),
    .RESET_B(net929),
    .D(_0137_),
    .Q_N(\uart_0.rx.rx_data_in ),
    .Q(_0136_));
 sg13g2_tielo tt_um_uart_bgdtanasa_3 (.L_LO(net3));
 sg13g2_tielo tt_um_uart_bgdtanasa_4 (.L_LO(net4));
 sg13g2_tielo tt_um_uart_bgdtanasa_5 (.L_LO(net5));
 sg13g2_tielo tt_um_uart_bgdtanasa_6 (.L_LO(net6));
 sg13g2_tielo tt_um_uart_bgdtanasa_7 (.L_LO(net7));
 sg13g2_tielo tt_um_uart_bgdtanasa_8 (.L_LO(net8));
 sg13g2_tielo tt_um_uart_bgdtanasa_9 (.L_LO(net9));
 sg13g2_tielo tt_um_uart_bgdtanasa_10 (.L_LO(net10));
 sg13g2_tielo tt_um_uart_bgdtanasa_11 (.L_LO(net11));
 sg13g2_tielo tt_um_uart_bgdtanasa_12 (.L_LO(net12));
 sg13g2_tielo tt_um_uart_bgdtanasa_13 (.L_LO(net13));
 sg13g2_tielo tt_um_uart_bgdtanasa_14 (.L_LO(net14));
 sg13g2_tielo tt_um_uart_bgdtanasa_15 (.L_LO(net15));
 sg13g2_tielo tt_um_uart_bgdtanasa_16 (.L_LO(net16));
 sg13g2_tielo tt_um_uart_bgdtanasa_17 (.L_LO(net17));
 sg13g2_tielo tt_um_uart_bgdtanasa_18 (.L_LO(net18));
 sg13g2_tielo tt_um_uart_bgdtanasa_19 (.L_LO(net19));
 sg13g2_tielo tt_um_uart_bgdtanasa_20 (.L_LO(net20));
 sg13g2_tielo tt_um_uart_bgdtanasa_21 (.L_LO(net21));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_2 _3181_ (.A(rx_data_ready),
    .X(uo_out[0]));
 sg13g2_buf_2 _3182_ (.A(net847),
    .X(uo_out[1]));
 sg13g2_buf_1 _3183_ (.A(tx_data_out),
    .X(uo_out[2]));
 sg13g2_buf_2 _3184_ (.A(tx_data_done),
    .X(uo_out[3]));
 sg13g2_buf_4 fanout701 (.X(net701),
    .A(_0623_));
 sg13g2_buf_4 fanout702 (.X(net702),
    .A(_0623_));
 sg13g2_buf_2 fanout703 (.A(net704),
    .X(net703));
 sg13g2_buf_4 fanout704 (.X(net704),
    .A(net705));
 sg13g2_buf_2 fanout705 (.A(_0600_),
    .X(net705));
 sg13g2_buf_4 fanout706 (.X(net706),
    .A(net707));
 sg13g2_buf_4 fanout707 (.X(net707),
    .A(_0574_));
 sg13g2_buf_4 fanout708 (.X(net708),
    .A(net709));
 sg13g2_buf_4 fanout709 (.X(net709),
    .A(_0550_));
 sg13g2_buf_4 fanout710 (.X(net710),
    .A(net711));
 sg13g2_buf_4 fanout711 (.X(net711),
    .A(_0526_));
 sg13g2_buf_4 fanout712 (.X(net712),
    .A(_0502_));
 sg13g2_buf_4 fanout713 (.X(net713),
    .A(_0502_));
 sg13g2_buf_4 fanout714 (.X(net714),
    .A(_0477_));
 sg13g2_buf_4 fanout715 (.X(net715),
    .A(_0477_));
 sg13g2_buf_4 fanout716 (.X(net716),
    .A(_0451_));
 sg13g2_buf_2 fanout717 (.A(_0451_),
    .X(net717));
 sg13g2_buf_2 fanout718 (.A(_0421_),
    .X(net718));
 sg13g2_buf_2 fanout719 (.A(net720),
    .X(net719));
 sg13g2_buf_4 fanout720 (.X(net720),
    .A(_1191_));
 sg13g2_buf_2 fanout721 (.A(net722),
    .X(net721));
 sg13g2_buf_2 fanout722 (.A(_1013_),
    .X(net722));
 sg13g2_buf_2 fanout723 (.A(net724),
    .X(net723));
 sg13g2_buf_2 fanout724 (.A(_0935_),
    .X(net724));
 sg13g2_buf_2 fanout725 (.A(_0873_),
    .X(net725));
 sg13g2_buf_2 fanout726 (.A(_0867_),
    .X(net726));
 sg13g2_buf_2 fanout727 (.A(net730),
    .X(net727));
 sg13g2_buf_2 fanout728 (.A(net730),
    .X(net728));
 sg13g2_buf_2 fanout729 (.A(net730),
    .X(net729));
 sg13g2_buf_2 fanout730 (.A(_0872_),
    .X(net730));
 sg13g2_buf_2 fanout731 (.A(_0420_),
    .X(net731));
 sg13g2_buf_4 fanout732 (.X(net732),
    .A(_0861_));
 sg13g2_buf_2 fanout733 (.A(net737),
    .X(net733));
 sg13g2_buf_2 fanout734 (.A(net737),
    .X(net734));
 sg13g2_buf_2 fanout735 (.A(net737),
    .X(net735));
 sg13g2_buf_2 fanout736 (.A(net737),
    .X(net736));
 sg13g2_buf_1 fanout737 (.A(net750),
    .X(net737));
 sg13g2_buf_2 fanout738 (.A(net739),
    .X(net738));
 sg13g2_buf_2 fanout739 (.A(net742),
    .X(net739));
 sg13g2_buf_2 fanout740 (.A(net742),
    .X(net740));
 sg13g2_buf_1 fanout741 (.A(net742),
    .X(net741));
 sg13g2_buf_2 fanout742 (.A(net750),
    .X(net742));
 sg13g2_buf_2 fanout743 (.A(net746),
    .X(net743));
 sg13g2_buf_2 fanout744 (.A(net746),
    .X(net744));
 sg13g2_buf_2 fanout745 (.A(net746),
    .X(net745));
 sg13g2_buf_2 fanout746 (.A(net750),
    .X(net746));
 sg13g2_buf_2 fanout747 (.A(net749),
    .X(net747));
 sg13g2_buf_2 fanout748 (.A(net749),
    .X(net748));
 sg13g2_buf_2 fanout749 (.A(net750),
    .X(net749));
 sg13g2_buf_2 fanout750 (.A(_0785_),
    .X(net750));
 sg13g2_buf_4 fanout751 (.X(net751),
    .A(net753));
 sg13g2_buf_1 fanout752 (.A(net753),
    .X(net752));
 sg13g2_buf_4 fanout753 (.X(net753),
    .A(_0754_));
 sg13g2_buf_2 fanout754 (.A(_0012_),
    .X(net754));
 sg13g2_buf_4 fanout755 (.X(net755),
    .A(_0821_));
 sg13g2_buf_4 fanout756 (.X(net756),
    .A(_0815_));
 sg13g2_buf_2 fanout757 (.A(_0815_),
    .X(net757));
 sg13g2_buf_2 fanout758 (.A(net761),
    .X(net758));
 sg13g2_buf_2 fanout759 (.A(net761),
    .X(net759));
 sg13g2_buf_2 fanout760 (.A(net761),
    .X(net760));
 sg13g2_buf_2 fanout761 (.A(_0804_),
    .X(net761));
 sg13g2_buf_2 fanout762 (.A(net766),
    .X(net762));
 sg13g2_buf_2 fanout763 (.A(net765),
    .X(net763));
 sg13g2_buf_2 fanout764 (.A(net765),
    .X(net764));
 sg13g2_buf_1 fanout765 (.A(net766),
    .X(net765));
 sg13g2_buf_2 fanout766 (.A(_0804_),
    .X(net766));
 sg13g2_buf_2 fanout767 (.A(net768),
    .X(net767));
 sg13g2_buf_4 fanout768 (.X(net768),
    .A(net771));
 sg13g2_buf_4 fanout769 (.X(net769),
    .A(net771));
 sg13g2_buf_2 fanout770 (.A(net771),
    .X(net770));
 sg13g2_buf_2 fanout771 (.A(_0804_),
    .X(net771));
 sg13g2_buf_4 fanout772 (.X(net772),
    .A(_0803_));
 sg13g2_buf_2 fanout773 (.A(_0803_),
    .X(net773));
 sg13g2_buf_4 fanout774 (.X(net774),
    .A(_0775_));
 sg13g2_buf_4 fanout775 (.X(net775),
    .A(net777));
 sg13g2_buf_1 fanout776 (.A(net777),
    .X(net776));
 sg13g2_buf_2 fanout777 (.A(_0681_),
    .X(net777));
 sg13g2_buf_4 fanout778 (.X(net778),
    .A(net779));
 sg13g2_buf_2 fanout779 (.A(_0672_),
    .X(net779));
 sg13g2_buf_2 fanout780 (.A(net781),
    .X(net780));
 sg13g2_buf_4 fanout781 (.X(net781),
    .A(_0662_));
 sg13g2_buf_2 fanout782 (.A(_1389_),
    .X(net782));
 sg13g2_buf_4 fanout783 (.X(net783),
    .A(_1380_));
 sg13g2_buf_2 fanout784 (.A(_1380_),
    .X(net784));
 sg13g2_buf_4 fanout785 (.X(net785),
    .A(_0825_));
 sg13g2_buf_4 fanout786 (.X(net786),
    .A(net787));
 sg13g2_buf_2 fanout787 (.A(_0819_),
    .X(net787));
 sg13g2_buf_2 fanout788 (.A(net789),
    .X(net788));
 sg13g2_buf_4 fanout789 (.X(net789),
    .A(_0745_));
 sg13g2_buf_2 fanout790 (.A(net791),
    .X(net790));
 sg13g2_buf_2 fanout791 (.A(_0736_),
    .X(net791));
 sg13g2_buf_2 fanout792 (.A(net793),
    .X(net792));
 sg13g2_buf_4 fanout793 (.X(net793),
    .A(_0727_));
 sg13g2_buf_2 fanout794 (.A(_0718_),
    .X(net794));
 sg13g2_buf_4 fanout795 (.X(net795),
    .A(_0718_));
 sg13g2_buf_2 fanout796 (.A(_0709_),
    .X(net796));
 sg13g2_buf_4 fanout797 (.X(net797),
    .A(_0709_));
 sg13g2_buf_2 fanout798 (.A(net799),
    .X(net798));
 sg13g2_buf_2 fanout799 (.A(net800),
    .X(net799));
 sg13g2_buf_2 fanout800 (.A(_0700_),
    .X(net800));
 sg13g2_buf_2 fanout801 (.A(net803),
    .X(net801));
 sg13g2_buf_1 fanout802 (.A(net803),
    .X(net802));
 sg13g2_buf_4 fanout803 (.X(net803),
    .A(_0691_));
 sg13g2_buf_2 fanout804 (.A(net806),
    .X(net804));
 sg13g2_buf_1 fanout805 (.A(net806),
    .X(net805));
 sg13g2_buf_2 fanout806 (.A(_0652_),
    .X(net806));
 sg13g2_buf_2 fanout807 (.A(net808),
    .X(net807));
 sg13g2_buf_4 fanout808 (.X(net808),
    .A(_0643_));
 sg13g2_buf_4 fanout809 (.X(net809),
    .A(_0634_));
 sg13g2_buf_2 fanout810 (.A(_0634_),
    .X(net810));
 sg13g2_buf_2 fanout811 (.A(net812),
    .X(net811));
 sg13g2_buf_4 fanout812 (.X(net812),
    .A(_0625_));
 sg13g2_buf_2 fanout813 (.A(_0426_),
    .X(net813));
 sg13g2_buf_2 fanout814 (.A(_0426_),
    .X(net814));
 sg13g2_buf_2 fanout815 (.A(net816),
    .X(net815));
 sg13g2_buf_2 fanout816 (.A(_1379_),
    .X(net816));
 sg13g2_buf_4 fanout817 (.X(net817),
    .A(_1379_));
 sg13g2_buf_2 fanout818 (.A(_1223_),
    .X(net818));
 sg13g2_buf_2 fanout819 (.A(\fifo_t[3] ),
    .X(net819));
 sg13g2_buf_2 fanout820 (.A(\fifo_t[3] ),
    .X(net820));
 sg13g2_buf_2 fanout821 (.A(\fifo_t[2] ),
    .X(net821));
 sg13g2_buf_2 fanout822 (.A(net823),
    .X(net822));
 sg13g2_buf_2 fanout823 (.A(_1248_),
    .X(net823));
 sg13g2_buf_2 fanout824 (.A(net825),
    .X(net824));
 sg13g2_buf_2 fanout825 (.A(net826),
    .X(net825));
 sg13g2_buf_2 fanout826 (.A(net834),
    .X(net826));
 sg13g2_buf_2 fanout827 (.A(net834),
    .X(net827));
 sg13g2_buf_2 fanout828 (.A(net834),
    .X(net828));
 sg13g2_buf_2 fanout829 (.A(net832),
    .X(net829));
 sg13g2_buf_1 fanout830 (.A(net832),
    .X(net830));
 sg13g2_buf_2 fanout831 (.A(net832),
    .X(net831));
 sg13g2_buf_1 fanout832 (.A(net833),
    .X(net832));
 sg13g2_buf_2 fanout833 (.A(net834),
    .X(net833));
 sg13g2_buf_2 fanout834 (.A(net847),
    .X(net834));
 sg13g2_buf_2 fanout835 (.A(net838),
    .X(net835));
 sg13g2_buf_1 fanout836 (.A(net838),
    .X(net836));
 sg13g2_buf_2 fanout837 (.A(net838),
    .X(net837));
 sg13g2_buf_1 fanout838 (.A(net846),
    .X(net838));
 sg13g2_buf_2 fanout839 (.A(net846),
    .X(net839));
 sg13g2_buf_2 fanout840 (.A(net846),
    .X(net840));
 sg13g2_buf_2 fanout841 (.A(net843),
    .X(net841));
 sg13g2_buf_2 fanout842 (.A(net843),
    .X(net842));
 sg13g2_buf_2 fanout843 (.A(net845),
    .X(net843));
 sg13g2_buf_2 fanout844 (.A(net845),
    .X(net844));
 sg13g2_buf_2 fanout845 (.A(net846),
    .X(net845));
 sg13g2_buf_1 fanout846 (.A(net847),
    .X(net846));
 sg13g2_buf_2 fanout847 (.A(rx_sample_clk),
    .X(net847));
 sg13g2_buf_2 fanout848 (.A(\uart_0.rx.rx_marker[2] ),
    .X(net848));
 sg13g2_buf_4 fanout849 (.X(net849),
    .A(net850));
 sg13g2_buf_2 fanout850 (.A(\uart_0.rx.rx_stop_zeros[3] ),
    .X(net850));
 sg13g2_buf_4 fanout851 (.X(net851),
    .A(\uart_0.rx.rx_stop_zeros[0] ));
 sg13g2_buf_2 fanout852 (.A(\uart_0.rx.rx_stop_zeros[0] ),
    .X(net852));
 sg13g2_buf_4 fanout853 (.X(net853),
    .A(\fifo_h[3] ));
 sg13g2_buf_4 fanout854 (.X(net854),
    .A(\fifo_h[2] ));
 sg13g2_buf_4 fanout855 (.X(net855),
    .A(\fifo_h[1] ));
 sg13g2_buf_4 fanout856 (.X(net856),
    .A(\fifo_h[0] ));
 sg13g2_buf_2 fanout857 (.A(net858),
    .X(net857));
 sg13g2_buf_2 fanout858 (.A(net863),
    .X(net858));
 sg13g2_buf_2 fanout859 (.A(net860),
    .X(net859));
 sg13g2_buf_2 fanout860 (.A(net862),
    .X(net860));
 sg13g2_buf_2 fanout861 (.A(net862),
    .X(net861));
 sg13g2_buf_2 fanout862 (.A(net863),
    .X(net862));
 sg13g2_buf_1 fanout863 (.A(net868),
    .X(net863));
 sg13g2_buf_2 fanout864 (.A(net868),
    .X(net864));
 sg13g2_buf_2 fanout865 (.A(net868),
    .X(net865));
 sg13g2_buf_2 fanout866 (.A(net867),
    .X(net866));
 sg13g2_buf_2 fanout867 (.A(net868),
    .X(net867));
 sg13g2_buf_4 fanout868 (.X(net868),
    .A(clk_out));
 sg13g2_buf_2 fanout869 (.A(net870),
    .X(net869));
 sg13g2_buf_2 fanout870 (.A(net875),
    .X(net870));
 sg13g2_buf_1 fanout871 (.A(net875),
    .X(net871));
 sg13g2_buf_2 fanout872 (.A(net875),
    .X(net872));
 sg13g2_buf_1 fanout873 (.A(net875),
    .X(net873));
 sg13g2_buf_2 fanout874 (.A(net875),
    .X(net874));
 sg13g2_buf_2 fanout875 (.A(net883),
    .X(net875));
 sg13g2_buf_2 fanout876 (.A(net877),
    .X(net876));
 sg13g2_buf_1 fanout877 (.A(net883),
    .X(net877));
 sg13g2_buf_2 fanout878 (.A(net879),
    .X(net878));
 sg13g2_buf_2 fanout879 (.A(net883),
    .X(net879));
 sg13g2_buf_2 fanout880 (.A(net882),
    .X(net880));
 sg13g2_buf_2 fanout881 (.A(net882),
    .X(net881));
 sg13g2_buf_2 fanout882 (.A(net883),
    .X(net882));
 sg13g2_buf_2 fanout883 (.A(clk_out),
    .X(net883));
 sg13g2_buf_4 fanout884 (.X(net884),
    .A(net885));
 sg13g2_buf_4 fanout885 (.X(net885),
    .A(net887));
 sg13g2_buf_4 fanout886 (.X(net886),
    .A(net887));
 sg13g2_buf_4 fanout887 (.X(net887),
    .A(net904));
 sg13g2_buf_4 fanout888 (.X(net888),
    .A(net891));
 sg13g2_buf_4 fanout889 (.X(net889),
    .A(net890));
 sg13g2_buf_4 fanout890 (.X(net890),
    .A(net891));
 sg13g2_buf_2 fanout891 (.A(net904),
    .X(net891));
 sg13g2_buf_4 fanout892 (.X(net892),
    .A(net893));
 sg13g2_buf_4 fanout893 (.X(net893),
    .A(net904));
 sg13g2_buf_4 fanout894 (.X(net894),
    .A(net896));
 sg13g2_buf_4 fanout895 (.X(net895),
    .A(net896));
 sg13g2_buf_4 fanout896 (.X(net896),
    .A(net904));
 sg13g2_buf_4 fanout897 (.X(net897),
    .A(net899));
 sg13g2_buf_4 fanout898 (.X(net898),
    .A(net899));
 sg13g2_buf_2 fanout899 (.A(net904),
    .X(net899));
 sg13g2_buf_4 fanout900 (.X(net900),
    .A(net903));
 sg13g2_buf_4 fanout901 (.X(net901),
    .A(net902));
 sg13g2_buf_4 fanout902 (.X(net902),
    .A(net903));
 sg13g2_buf_2 fanout903 (.A(net904),
    .X(net903));
 sg13g2_buf_4 fanout904 (.X(net904),
    .A(rst_n));
 sg13g2_buf_4 fanout905 (.X(net905),
    .A(net907));
 sg13g2_buf_2 fanout906 (.A(net907),
    .X(net906));
 sg13g2_buf_4 fanout907 (.X(net907),
    .A(net908));
 sg13g2_buf_4 fanout908 (.X(net908),
    .A(net919));
 sg13g2_buf_4 fanout909 (.X(net909),
    .A(net910));
 sg13g2_buf_4 fanout910 (.X(net910),
    .A(net919));
 sg13g2_buf_4 fanout911 (.X(net911),
    .A(net912));
 sg13g2_buf_4 fanout912 (.X(net912),
    .A(net915));
 sg13g2_buf_4 fanout913 (.X(net913),
    .A(net915));
 sg13g2_buf_2 fanout914 (.A(net915),
    .X(net914));
 sg13g2_buf_2 fanout915 (.A(net919),
    .X(net915));
 sg13g2_buf_4 fanout916 (.X(net916),
    .A(net918));
 sg13g2_buf_4 fanout917 (.X(net917),
    .A(net918));
 sg13g2_buf_4 fanout918 (.X(net918),
    .A(net919));
 sg13g2_buf_2 fanout919 (.A(rst_n),
    .X(net919));
 sg13g2_buf_4 fanout920 (.X(net920),
    .A(net930));
 sg13g2_buf_4 fanout921 (.X(net921),
    .A(net930));
 sg13g2_buf_4 fanout922 (.X(net922),
    .A(net923));
 sg13g2_buf_4 fanout923 (.X(net923),
    .A(net930));
 sg13g2_buf_4 fanout924 (.X(net924),
    .A(net926));
 sg13g2_buf_2 fanout925 (.A(net926),
    .X(net925));
 sg13g2_buf_4 fanout926 (.X(net926),
    .A(net930));
 sg13g2_buf_4 fanout927 (.X(net927),
    .A(net930));
 sg13g2_buf_4 fanout928 (.X(net928),
    .A(net929));
 sg13g2_buf_4 fanout929 (.X(net929),
    .A(net930));
 sg13g2_buf_4 fanout930 (.X(net930),
    .A(rst_n));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_tielo tt_um_uart_bgdtanasa_2 (.L_LO(net2));
 sg13g2_buf_2 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .X(clknet_1_0__leaf_clk));
 sg13g2_buf_2 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .X(clknet_1_1__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_1_1__leaf_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(_0038_),
    .X(net22));
 sg13g2_dlygate4sd3_1 hold2 (.A(_0138_),
    .X(net23));
 sg13g2_dlygate4sd3_1 hold3 (.A(\clk_out_cnt[3] ),
    .X(net24));
 sg13g2_dlygate4sd3_1 hold4 (.A(_0003_),
    .X(net25));
 sg13g2_dlygate4sd3_1 hold5 (.A(\clk_out_cnt[0] ),
    .X(net26));
 sg13g2_dlygate4sd3_1 hold6 (.A(_0000_),
    .X(net27));
 sg13g2_dlygate4sd3_1 hold7 (.A(\clk_out_cnt[1] ),
    .X(net28));
 sg13g2_dlygate4sd3_1 hold8 (.A(\clk_out_cnt[2] ),
    .X(net29));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_4 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_317 ();
 sg13g2_fill_1 FILLER_4_327 ();
 sg13g2_decap_8 FILLER_4_333 ();
 sg13g2_decap_8 FILLER_4_340 ();
 sg13g2_decap_8 FILLER_4_347 ();
 sg13g2_decap_8 FILLER_4_354 ();
 sg13g2_decap_8 FILLER_4_361 ();
 sg13g2_decap_8 FILLER_4_368 ();
 sg13g2_decap_8 FILLER_4_375 ();
 sg13g2_decap_8 FILLER_4_382 ();
 sg13g2_decap_8 FILLER_4_389 ();
 sg13g2_decap_8 FILLER_4_396 ();
 sg13g2_decap_4 FILLER_4_403 ();
 sg13g2_fill_2 FILLER_4_407 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_fill_2 FILLER_5_256 ();
 sg13g2_decap_8 FILLER_5_262 ();
 sg13g2_decap_8 FILLER_5_269 ();
 sg13g2_decap_8 FILLER_5_276 ();
 sg13g2_decap_8 FILLER_5_283 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_4 FILLER_6_238 ();
 sg13g2_fill_2 FILLER_6_242 ();
 sg13g2_decap_4 FILLER_6_279 ();
 sg13g2_fill_2 FILLER_6_283 ();
 sg13g2_fill_1 FILLER_6_311 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_fill_2 FILLER_7_238 ();
 sg13g2_fill_2 FILLER_7_281 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_279 ();
 sg13g2_fill_2 FILLER_8_286 ();
 sg13g2_fill_1 FILLER_8_288 ();
 sg13g2_decap_4 FILLER_8_322 ();
 sg13g2_fill_1 FILLER_8_326 ();
 sg13g2_fill_2 FILLER_8_331 ();
 sg13g2_fill_2 FILLER_8_337 ();
 sg13g2_decap_8 FILLER_8_342 ();
 sg13g2_decap_8 FILLER_8_349 ();
 sg13g2_decap_8 FILLER_8_356 ();
 sg13g2_decap_8 FILLER_8_363 ();
 sg13g2_decap_8 FILLER_8_370 ();
 sg13g2_decap_8 FILLER_8_377 ();
 sg13g2_decap_8 FILLER_8_384 ();
 sg13g2_decap_8 FILLER_8_391 ();
 sg13g2_decap_8 FILLER_8_398 ();
 sg13g2_decap_4 FILLER_8_405 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_4 FILLER_9_245 ();
 sg13g2_fill_2 FILLER_9_249 ();
 sg13g2_fill_2 FILLER_9_256 ();
 sg13g2_fill_1 FILLER_9_258 ();
 sg13g2_decap_8 FILLER_9_263 ();
 sg13g2_decap_8 FILLER_9_270 ();
 sg13g2_decap_4 FILLER_9_277 ();
 sg13g2_fill_1 FILLER_9_281 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_fill_1 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_309 ();
 sg13g2_decap_8 FILLER_9_316 ();
 sg13g2_decap_8 FILLER_9_323 ();
 sg13g2_decap_8 FILLER_9_330 ();
 sg13g2_decap_8 FILLER_9_337 ();
 sg13g2_decap_8 FILLER_9_344 ();
 sg13g2_decap_8 FILLER_9_351 ();
 sg13g2_decap_8 FILLER_9_358 ();
 sg13g2_decap_8 FILLER_9_365 ();
 sg13g2_decap_8 FILLER_9_372 ();
 sg13g2_decap_8 FILLER_9_379 ();
 sg13g2_decap_8 FILLER_9_386 ();
 sg13g2_decap_8 FILLER_9_393 ();
 sg13g2_decap_8 FILLER_9_400 ();
 sg13g2_fill_2 FILLER_9_407 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_4 FILLER_10_224 ();
 sg13g2_fill_2 FILLER_10_228 ();
 sg13g2_fill_2 FILLER_10_256 ();
 sg13g2_fill_1 FILLER_10_258 ();
 sg13g2_fill_1 FILLER_10_288 ();
 sg13g2_decap_4 FILLER_10_297 ();
 sg13g2_fill_1 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_313 ();
 sg13g2_decap_8 FILLER_10_346 ();
 sg13g2_decap_8 FILLER_10_353 ();
 sg13g2_decap_8 FILLER_10_360 ();
 sg13g2_decap_8 FILLER_10_367 ();
 sg13g2_decap_8 FILLER_10_374 ();
 sg13g2_decap_8 FILLER_10_381 ();
 sg13g2_decap_8 FILLER_10_388 ();
 sg13g2_decap_8 FILLER_10_395 ();
 sg13g2_decap_8 FILLER_10_402 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_4 FILLER_11_224 ();
 sg13g2_fill_1 FILLER_11_228 ();
 sg13g2_decap_8 FILLER_11_255 ();
 sg13g2_fill_1 FILLER_11_262 ();
 sg13g2_fill_1 FILLER_11_268 ();
 sg13g2_fill_1 FILLER_11_274 ();
 sg13g2_fill_2 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_353 ();
 sg13g2_decap_8 FILLER_11_360 ();
 sg13g2_decap_8 FILLER_11_367 ();
 sg13g2_decap_8 FILLER_11_374 ();
 sg13g2_decap_8 FILLER_11_381 ();
 sg13g2_decap_8 FILLER_11_388 ();
 sg13g2_decap_8 FILLER_11_395 ();
 sg13g2_decap_8 FILLER_11_402 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_4 FILLER_12_217 ();
 sg13g2_fill_1 FILLER_12_250 ();
 sg13g2_decap_8 FILLER_12_355 ();
 sg13g2_decap_8 FILLER_12_362 ();
 sg13g2_decap_8 FILLER_12_369 ();
 sg13g2_decap_8 FILLER_12_376 ();
 sg13g2_decap_8 FILLER_12_383 ();
 sg13g2_decap_8 FILLER_12_390 ();
 sg13g2_decap_8 FILLER_12_397 ();
 sg13g2_decap_4 FILLER_12_404 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_4 FILLER_13_133 ();
 sg13g2_fill_1 FILLER_13_137 ();
 sg13g2_fill_1 FILLER_13_143 ();
 sg13g2_decap_8 FILLER_13_148 ();
 sg13g2_decap_8 FILLER_13_155 ();
 sg13g2_decap_8 FILLER_13_162 ();
 sg13g2_decap_8 FILLER_13_169 ();
 sg13g2_decap_8 FILLER_13_176 ();
 sg13g2_decap_8 FILLER_13_183 ();
 sg13g2_decap_8 FILLER_13_190 ();
 sg13g2_decap_8 FILLER_13_197 ();
 sg13g2_decap_8 FILLER_13_204 ();
 sg13g2_decap_8 FILLER_13_211 ();
 sg13g2_decap_8 FILLER_13_218 ();
 sg13g2_fill_2 FILLER_13_225 ();
 sg13g2_fill_1 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_351 ();
 sg13g2_decap_8 FILLER_13_358 ();
 sg13g2_decap_8 FILLER_13_365 ();
 sg13g2_decap_8 FILLER_13_372 ();
 sg13g2_decap_8 FILLER_13_379 ();
 sg13g2_decap_8 FILLER_13_386 ();
 sg13g2_decap_8 FILLER_13_393 ();
 sg13g2_decap_8 FILLER_13_400 ();
 sg13g2_fill_2 FILLER_13_407 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_fill_2 FILLER_14_119 ();
 sg13g2_fill_1 FILLER_14_121 ();
 sg13g2_fill_2 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_fill_2 FILLER_14_231 ();
 sg13g2_fill_1 FILLER_14_233 ();
 sg13g2_decap_8 FILLER_14_237 ();
 sg13g2_fill_2 FILLER_14_244 ();
 sg13g2_fill_1 FILLER_14_246 ();
 sg13g2_decap_8 FILLER_14_290 ();
 sg13g2_decap_8 FILLER_14_297 ();
 sg13g2_decap_8 FILLER_14_304 ();
 sg13g2_decap_4 FILLER_14_311 ();
 sg13g2_fill_1 FILLER_14_315 ();
 sg13g2_fill_2 FILLER_14_332 ();
 sg13g2_fill_1 FILLER_14_334 ();
 sg13g2_decap_4 FILLER_14_340 ();
 sg13g2_decap_8 FILLER_14_359 ();
 sg13g2_decap_8 FILLER_14_366 ();
 sg13g2_decap_8 FILLER_14_373 ();
 sg13g2_decap_8 FILLER_14_380 ();
 sg13g2_decap_8 FILLER_14_387 ();
 sg13g2_decap_8 FILLER_14_394 ();
 sg13g2_decap_8 FILLER_14_401 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_fill_2 FILLER_15_105 ();
 sg13g2_fill_2 FILLER_15_133 ();
 sg13g2_fill_1 FILLER_15_166 ();
 sg13g2_decap_8 FILLER_15_193 ();
 sg13g2_decap_8 FILLER_15_200 ();
 sg13g2_decap_8 FILLER_15_207 ();
 sg13g2_decap_8 FILLER_15_214 ();
 sg13g2_decap_8 FILLER_15_221 ();
 sg13g2_decap_8 FILLER_15_228 ();
 sg13g2_decap_4 FILLER_15_235 ();
 sg13g2_fill_1 FILLER_15_239 ();
 sg13g2_decap_8 FILLER_15_247 ();
 sg13g2_decap_8 FILLER_15_254 ();
 sg13g2_fill_1 FILLER_15_261 ();
 sg13g2_decap_8 FILLER_15_281 ();
 sg13g2_fill_2 FILLER_15_288 ();
 sg13g2_fill_1 FILLER_15_290 ();
 sg13g2_fill_1 FILLER_15_298 ();
 sg13g2_fill_1 FILLER_15_309 ();
 sg13g2_fill_2 FILLER_15_318 ();
 sg13g2_decap_8 FILLER_15_332 ();
 sg13g2_fill_1 FILLER_15_339 ();
 sg13g2_decap_8 FILLER_15_366 ();
 sg13g2_decap_8 FILLER_15_373 ();
 sg13g2_decap_8 FILLER_15_380 ();
 sg13g2_decap_8 FILLER_15_387 ();
 sg13g2_decap_8 FILLER_15_394 ();
 sg13g2_decap_8 FILLER_15_401 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_4 FILLER_16_98 ();
 sg13g2_fill_2 FILLER_16_160 ();
 sg13g2_fill_1 FILLER_16_162 ();
 sg13g2_fill_2 FILLER_16_173 ();
 sg13g2_decap_8 FILLER_16_207 ();
 sg13g2_decap_8 FILLER_16_214 ();
 sg13g2_fill_2 FILLER_16_221 ();
 sg13g2_fill_1 FILLER_16_223 ();
 sg13g2_decap_8 FILLER_16_253 ();
 sg13g2_decap_8 FILLER_16_260 ();
 sg13g2_decap_8 FILLER_16_267 ();
 sg13g2_fill_2 FILLER_16_274 ();
 sg13g2_decap_8 FILLER_16_333 ();
 sg13g2_decap_8 FILLER_16_366 ();
 sg13g2_decap_8 FILLER_16_373 ();
 sg13g2_decap_8 FILLER_16_380 ();
 sg13g2_decap_8 FILLER_16_387 ();
 sg13g2_decap_8 FILLER_16_394 ();
 sg13g2_decap_8 FILLER_16_401 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_fill_2 FILLER_17_105 ();
 sg13g2_fill_1 FILLER_17_107 ();
 sg13g2_decap_4 FILLER_17_132 ();
 sg13g2_fill_1 FILLER_17_136 ();
 sg13g2_fill_1 FILLER_17_142 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_4 FILLER_17_161 ();
 sg13g2_decap_4 FILLER_17_177 ();
 sg13g2_fill_1 FILLER_17_181 ();
 sg13g2_decap_4 FILLER_17_191 ();
 sg13g2_decap_8 FILLER_17_203 ();
 sg13g2_decap_8 FILLER_17_210 ();
 sg13g2_decap_4 FILLER_17_217 ();
 sg13g2_decap_8 FILLER_17_272 ();
 sg13g2_fill_2 FILLER_17_279 ();
 sg13g2_fill_1 FILLER_17_291 ();
 sg13g2_decap_8 FILLER_17_300 ();
 sg13g2_fill_1 FILLER_17_307 ();
 sg13g2_decap_8 FILLER_17_315 ();
 sg13g2_decap_8 FILLER_17_322 ();
 sg13g2_decap_4 FILLER_17_329 ();
 sg13g2_fill_1 FILLER_17_333 ();
 sg13g2_fill_2 FILLER_17_337 ();
 sg13g2_fill_1 FILLER_17_339 ();
 sg13g2_fill_1 FILLER_17_362 ();
 sg13g2_decap_8 FILLER_17_378 ();
 sg13g2_decap_8 FILLER_17_385 ();
 sg13g2_decap_8 FILLER_17_392 ();
 sg13g2_decap_8 FILLER_17_399 ();
 sg13g2_fill_2 FILLER_17_406 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_fill_1 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_128 ();
 sg13g2_decap_8 FILLER_18_135 ();
 sg13g2_decap_8 FILLER_18_142 ();
 sg13g2_decap_4 FILLER_18_149 ();
 sg13g2_fill_1 FILLER_18_153 ();
 sg13g2_fill_2 FILLER_18_206 ();
 sg13g2_decap_4 FILLER_18_216 ();
 sg13g2_fill_1 FILLER_18_220 ();
 sg13g2_decap_8 FILLER_18_226 ();
 sg13g2_fill_2 FILLER_18_233 ();
 sg13g2_decap_8 FILLER_18_285 ();
 sg13g2_decap_8 FILLER_18_301 ();
 sg13g2_fill_2 FILLER_18_308 ();
 sg13g2_decap_8 FILLER_18_386 ();
 sg13g2_decap_8 FILLER_18_393 ();
 sg13g2_decap_8 FILLER_18_400 ();
 sg13g2_fill_2 FILLER_18_407 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_fill_2 FILLER_19_105 ();
 sg13g2_fill_1 FILLER_19_107 ();
 sg13g2_fill_2 FILLER_19_160 ();
 sg13g2_fill_2 FILLER_19_172 ();
 sg13g2_fill_1 FILLER_19_174 ();
 sg13g2_decap_4 FILLER_19_209 ();
 sg13g2_fill_1 FILLER_19_213 ();
 sg13g2_decap_4 FILLER_19_240 ();
 sg13g2_fill_2 FILLER_19_244 ();
 sg13g2_decap_8 FILLER_19_251 ();
 sg13g2_decap_4 FILLER_19_258 ();
 sg13g2_decap_4 FILLER_19_266 ();
 sg13g2_fill_1 FILLER_19_270 ();
 sg13g2_fill_2 FILLER_19_279 ();
 sg13g2_decap_4 FILLER_19_340 ();
 sg13g2_decap_8 FILLER_19_352 ();
 sg13g2_decap_4 FILLER_19_359 ();
 sg13g2_decap_8 FILLER_19_386 ();
 sg13g2_decap_8 FILLER_19_393 ();
 sg13g2_decap_8 FILLER_19_400 ();
 sg13g2_fill_2 FILLER_19_407 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_fill_2 FILLER_20_98 ();
 sg13g2_fill_2 FILLER_20_140 ();
 sg13g2_fill_1 FILLER_20_173 ();
 sg13g2_fill_2 FILLER_20_210 ();
 sg13g2_fill_1 FILLER_20_212 ();
 sg13g2_decap_4 FILLER_20_252 ();
 sg13g2_fill_1 FILLER_20_256 ();
 sg13g2_fill_1 FILLER_20_267 ();
 sg13g2_fill_1 FILLER_20_281 ();
 sg13g2_fill_1 FILLER_20_296 ();
 sg13g2_decap_8 FILLER_20_350 ();
 sg13g2_decap_8 FILLER_20_357 ();
 sg13g2_fill_2 FILLER_20_364 ();
 sg13g2_fill_1 FILLER_20_366 ();
 sg13g2_decap_8 FILLER_20_382 ();
 sg13g2_decap_8 FILLER_20_389 ();
 sg13g2_decap_8 FILLER_20_396 ();
 sg13g2_decap_4 FILLER_20_403 ();
 sg13g2_fill_2 FILLER_20_407 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_4 FILLER_21_84 ();
 sg13g2_fill_2 FILLER_21_88 ();
 sg13g2_fill_1 FILLER_21_116 ();
 sg13g2_fill_1 FILLER_21_158 ();
 sg13g2_fill_1 FILLER_21_164 ();
 sg13g2_decap_8 FILLER_21_194 ();
 sg13g2_decap_8 FILLER_21_201 ();
 sg13g2_decap_4 FILLER_21_208 ();
 sg13g2_fill_2 FILLER_21_212 ();
 sg13g2_decap_4 FILLER_21_281 ();
 sg13g2_fill_1 FILLER_21_288 ();
 sg13g2_decap_4 FILLER_21_309 ();
 sg13g2_decap_4 FILLER_21_338 ();
 sg13g2_fill_1 FILLER_21_342 ();
 sg13g2_decap_8 FILLER_21_350 ();
 sg13g2_fill_2 FILLER_21_357 ();
 sg13g2_decap_8 FILLER_21_386 ();
 sg13g2_decap_8 FILLER_21_393 ();
 sg13g2_decap_8 FILLER_21_400 ();
 sg13g2_fill_2 FILLER_21_407 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_4 FILLER_22_91 ();
 sg13g2_fill_1 FILLER_22_95 ();
 sg13g2_fill_2 FILLER_22_106 ();
 sg13g2_fill_1 FILLER_22_108 ();
 sg13g2_decap_8 FILLER_22_118 ();
 sg13g2_decap_4 FILLER_22_125 ();
 sg13g2_decap_8 FILLER_22_139 ();
 sg13g2_fill_2 FILLER_22_146 ();
 sg13g2_fill_1 FILLER_22_148 ();
 sg13g2_fill_2 FILLER_22_154 ();
 sg13g2_decap_8 FILLER_22_160 ();
 sg13g2_decap_8 FILLER_22_167 ();
 sg13g2_decap_8 FILLER_22_174 ();
 sg13g2_decap_4 FILLER_22_181 ();
 sg13g2_fill_2 FILLER_22_185 ();
 sg13g2_decap_8 FILLER_22_191 ();
 sg13g2_decap_8 FILLER_22_198 ();
 sg13g2_decap_8 FILLER_22_205 ();
 sg13g2_decap_8 FILLER_22_212 ();
 sg13g2_fill_2 FILLER_22_219 ();
 sg13g2_fill_1 FILLER_22_221 ();
 sg13g2_decap_8 FILLER_22_225 ();
 sg13g2_decap_4 FILLER_22_232 ();
 sg13g2_fill_2 FILLER_22_236 ();
 sg13g2_fill_2 FILLER_22_244 ();
 sg13g2_fill_1 FILLER_22_246 ();
 sg13g2_fill_2 FILLER_22_253 ();
 sg13g2_decap_4 FILLER_22_261 ();
 sg13g2_decap_4 FILLER_22_270 ();
 sg13g2_decap_8 FILLER_22_279 ();
 sg13g2_decap_8 FILLER_22_286 ();
 sg13g2_decap_4 FILLER_22_293 ();
 sg13g2_decap_4 FILLER_22_306 ();
 sg13g2_fill_2 FILLER_22_310 ();
 sg13g2_decap_4 FILLER_22_319 ();
 sg13g2_decap_4 FILLER_22_328 ();
 sg13g2_fill_2 FILLER_22_336 ();
 sg13g2_fill_1 FILLER_22_338 ();
 sg13g2_decap_8 FILLER_22_378 ();
 sg13g2_decap_8 FILLER_22_385 ();
 sg13g2_decap_8 FILLER_22_392 ();
 sg13g2_decap_8 FILLER_22_399 ();
 sg13g2_fill_2 FILLER_22_406 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_4 FILLER_23_84 ();
 sg13g2_fill_2 FILLER_23_88 ();
 sg13g2_decap_8 FILLER_23_116 ();
 sg13g2_decap_8 FILLER_23_128 ();
 sg13g2_decap_8 FILLER_23_135 ();
 sg13g2_fill_1 FILLER_23_142 ();
 sg13g2_decap_8 FILLER_23_174 ();
 sg13g2_decap_8 FILLER_23_213 ();
 sg13g2_decap_8 FILLER_23_220 ();
 sg13g2_fill_1 FILLER_23_227 ();
 sg13g2_decap_8 FILLER_23_245 ();
 sg13g2_decap_8 FILLER_23_252 ();
 sg13g2_decap_4 FILLER_23_259 ();
 sg13g2_fill_1 FILLER_23_263 ();
 sg13g2_fill_1 FILLER_23_290 ();
 sg13g2_fill_2 FILLER_23_296 ();
 sg13g2_fill_1 FILLER_23_298 ();
 sg13g2_decap_8 FILLER_23_330 ();
 sg13g2_fill_2 FILLER_23_337 ();
 sg13g2_decap_4 FILLER_23_365 ();
 sg13g2_fill_1 FILLER_23_369 ();
 sg13g2_decap_8 FILLER_23_383 ();
 sg13g2_decap_8 FILLER_23_390 ();
 sg13g2_decap_8 FILLER_23_397 ();
 sg13g2_decap_4 FILLER_23_404 ();
 sg13g2_fill_1 FILLER_23_408 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_fill_1 FILLER_24_98 ();
 sg13g2_fill_1 FILLER_24_104 ();
 sg13g2_fill_2 FILLER_24_109 ();
 sg13g2_decap_8 FILLER_24_147 ();
 sg13g2_decap_8 FILLER_24_212 ();
 sg13g2_fill_1 FILLER_24_254 ();
 sg13g2_decap_8 FILLER_24_307 ();
 sg13g2_decap_8 FILLER_24_314 ();
 sg13g2_decap_4 FILLER_24_321 ();
 sg13g2_fill_1 FILLER_24_325 ();
 sg13g2_decap_8 FILLER_24_331 ();
 sg13g2_decap_4 FILLER_24_361 ();
 sg13g2_fill_2 FILLER_24_365 ();
 sg13g2_decap_8 FILLER_24_380 ();
 sg13g2_decap_8 FILLER_24_387 ();
 sg13g2_decap_8 FILLER_24_394 ();
 sg13g2_decap_8 FILLER_24_401 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_4 FILLER_25_84 ();
 sg13g2_fill_2 FILLER_25_88 ();
 sg13g2_fill_2 FILLER_25_120 ();
 sg13g2_fill_1 FILLER_25_122 ();
 sg13g2_decap_4 FILLER_25_164 ();
 sg13g2_fill_1 FILLER_25_168 ();
 sg13g2_fill_2 FILLER_25_179 ();
 sg13g2_fill_1 FILLER_25_181 ();
 sg13g2_fill_2 FILLER_25_198 ();
 sg13g2_fill_1 FILLER_25_200 ();
 sg13g2_fill_2 FILLER_25_209 ();
 sg13g2_fill_1 FILLER_25_211 ();
 sg13g2_fill_1 FILLER_25_224 ();
 sg13g2_decap_8 FILLER_25_263 ();
 sg13g2_fill_1 FILLER_25_270 ();
 sg13g2_fill_2 FILLER_25_278 ();
 sg13g2_fill_1 FILLER_25_291 ();
 sg13g2_decap_4 FILLER_25_307 ();
 sg13g2_decap_4 FILLER_25_342 ();
 sg13g2_decap_8 FILLER_25_379 ();
 sg13g2_decap_8 FILLER_25_386 ();
 sg13g2_decap_8 FILLER_25_393 ();
 sg13g2_decap_8 FILLER_25_400 ();
 sg13g2_fill_2 FILLER_25_407 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_4 FILLER_26_84 ();
 sg13g2_fill_2 FILLER_26_88 ();
 sg13g2_decap_8 FILLER_26_138 ();
 sg13g2_decap_4 FILLER_26_145 ();
 sg13g2_decap_4 FILLER_26_157 ();
 sg13g2_fill_2 FILLER_26_161 ();
 sg13g2_fill_1 FILLER_26_172 ();
 sg13g2_fill_2 FILLER_26_185 ();
 sg13g2_decap_8 FILLER_26_191 ();
 sg13g2_fill_2 FILLER_26_198 ();
 sg13g2_decap_8 FILLER_26_205 ();
 sg13g2_decap_8 FILLER_26_212 ();
 sg13g2_fill_2 FILLER_26_242 ();
 sg13g2_decap_8 FILLER_26_249 ();
 sg13g2_decap_4 FILLER_26_256 ();
 sg13g2_decap_8 FILLER_26_270 ();
 sg13g2_decap_8 FILLER_26_282 ();
 sg13g2_fill_2 FILLER_26_289 ();
 sg13g2_fill_1 FILLER_26_291 ();
 sg13g2_decap_4 FILLER_26_300 ();
 sg13g2_fill_1 FILLER_26_304 ();
 sg13g2_fill_2 FILLER_26_314 ();
 sg13g2_fill_1 FILLER_26_316 ();
 sg13g2_decap_8 FILLER_26_346 ();
 sg13g2_fill_2 FILLER_26_353 ();
 sg13g2_fill_1 FILLER_26_355 ();
 sg13g2_decap_8 FILLER_26_382 ();
 sg13g2_decap_8 FILLER_26_389 ();
 sg13g2_decap_8 FILLER_26_396 ();
 sg13g2_decap_4 FILLER_26_403 ();
 sg13g2_fill_2 FILLER_26_407 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_decap_8 FILLER_27_84 ();
 sg13g2_decap_8 FILLER_27_91 ();
 sg13g2_decap_4 FILLER_27_98 ();
 sg13g2_fill_2 FILLER_27_102 ();
 sg13g2_fill_2 FILLER_27_118 ();
 sg13g2_fill_1 FILLER_27_120 ();
 sg13g2_fill_1 FILLER_27_126 ();
 sg13g2_decap_8 FILLER_27_131 ();
 sg13g2_decap_8 FILLER_27_138 ();
 sg13g2_fill_1 FILLER_27_145 ();
 sg13g2_decap_8 FILLER_27_177 ();
 sg13g2_fill_2 FILLER_27_184 ();
 sg13g2_fill_1 FILLER_27_186 ();
 sg13g2_decap_8 FILLER_27_191 ();
 sg13g2_decap_8 FILLER_27_198 ();
 sg13g2_decap_8 FILLER_27_205 ();
 sg13g2_decap_8 FILLER_27_212 ();
 sg13g2_decap_8 FILLER_27_219 ();
 sg13g2_fill_1 FILLER_27_226 ();
 sg13g2_fill_1 FILLER_27_234 ();
 sg13g2_decap_8 FILLER_27_240 ();
 sg13g2_decap_8 FILLER_27_247 ();
 sg13g2_fill_1 FILLER_27_254 ();
 sg13g2_fill_2 FILLER_27_288 ();
 sg13g2_fill_1 FILLER_27_290 ();
 sg13g2_fill_2 FILLER_27_301 ();
 sg13g2_fill_1 FILLER_27_323 ();
 sg13g2_fill_2 FILLER_27_329 ();
 sg13g2_fill_2 FILLER_27_340 ();
 sg13g2_fill_1 FILLER_27_342 ();
 sg13g2_decap_8 FILLER_27_377 ();
 sg13g2_decap_8 FILLER_27_384 ();
 sg13g2_decap_8 FILLER_27_391 ();
 sg13g2_decap_8 FILLER_27_398 ();
 sg13g2_decap_4 FILLER_27_405 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_decap_8 FILLER_28_84 ();
 sg13g2_decap_8 FILLER_28_91 ();
 sg13g2_decap_8 FILLER_28_98 ();
 sg13g2_decap_4 FILLER_28_105 ();
 sg13g2_fill_1 FILLER_28_109 ();
 sg13g2_fill_2 FILLER_28_142 ();
 sg13g2_decap_4 FILLER_28_153 ();
 sg13g2_fill_2 FILLER_28_157 ();
 sg13g2_decap_8 FILLER_28_169 ();
 sg13g2_fill_2 FILLER_28_176 ();
 sg13g2_fill_2 FILLER_28_242 ();
 sg13g2_fill_1 FILLER_28_244 ();
 sg13g2_decap_4 FILLER_28_271 ();
 sg13g2_fill_2 FILLER_28_275 ();
 sg13g2_decap_8 FILLER_28_315 ();
 sg13g2_fill_2 FILLER_28_322 ();
 sg13g2_fill_1 FILLER_28_329 ();
 sg13g2_decap_8 FILLER_28_372 ();
 sg13g2_decap_8 FILLER_28_379 ();
 sg13g2_decap_8 FILLER_28_386 ();
 sg13g2_decap_8 FILLER_28_393 ();
 sg13g2_decap_8 FILLER_28_400 ();
 sg13g2_fill_2 FILLER_28_407 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_4 FILLER_29_77 ();
 sg13g2_fill_2 FILLER_29_81 ();
 sg13g2_decap_8 FILLER_29_109 ();
 sg13g2_decap_4 FILLER_29_116 ();
 sg13g2_fill_1 FILLER_29_125 ();
 sg13g2_fill_2 FILLER_29_130 ();
 sg13g2_fill_1 FILLER_29_132 ();
 sg13g2_decap_4 FILLER_29_159 ();
 sg13g2_fill_2 FILLER_29_163 ();
 sg13g2_fill_2 FILLER_29_169 ();
 sg13g2_decap_8 FILLER_29_258 ();
 sg13g2_fill_2 FILLER_29_265 ();
 sg13g2_fill_1 FILLER_29_267 ();
 sg13g2_fill_2 FILLER_29_290 ();
 sg13g2_fill_1 FILLER_29_292 ();
 sg13g2_decap_4 FILLER_29_298 ();
 sg13g2_fill_1 FILLER_29_302 ();
 sg13g2_decap_4 FILLER_29_309 ();
 sg13g2_fill_1 FILLER_29_313 ();
 sg13g2_fill_2 FILLER_29_347 ();
 sg13g2_decap_8 FILLER_29_385 ();
 sg13g2_decap_8 FILLER_29_392 ();
 sg13g2_decap_8 FILLER_29_399 ();
 sg13g2_fill_2 FILLER_29_406 ();
 sg13g2_fill_1 FILLER_29_408 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_77 ();
 sg13g2_fill_1 FILLER_30_84 ();
 sg13g2_fill_2 FILLER_30_141 ();
 sg13g2_fill_1 FILLER_30_151 ();
 sg13g2_fill_2 FILLER_30_157 ();
 sg13g2_fill_1 FILLER_30_159 ();
 sg13g2_decap_8 FILLER_30_212 ();
 sg13g2_fill_2 FILLER_30_219 ();
 sg13g2_decap_8 FILLER_30_255 ();
 sg13g2_decap_4 FILLER_30_262 ();
 sg13g2_decap_8 FILLER_30_273 ();
 sg13g2_decap_4 FILLER_30_280 ();
 sg13g2_decap_4 FILLER_30_289 ();
 sg13g2_fill_2 FILLER_30_298 ();
 sg13g2_fill_1 FILLER_30_300 ();
 sg13g2_fill_2 FILLER_30_316 ();
 sg13g2_fill_1 FILLER_30_318 ();
 sg13g2_decap_8 FILLER_30_353 ();
 sg13g2_decap_8 FILLER_30_360 ();
 sg13g2_decap_8 FILLER_30_367 ();
 sg13g2_decap_8 FILLER_30_374 ();
 sg13g2_decap_8 FILLER_30_381 ();
 sg13g2_decap_8 FILLER_30_388 ();
 sg13g2_decap_8 FILLER_30_395 ();
 sg13g2_decap_8 FILLER_30_402 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_decap_4 FILLER_31_84 ();
 sg13g2_fill_2 FILLER_31_88 ();
 sg13g2_fill_2 FILLER_31_104 ();
 sg13g2_fill_1 FILLER_31_106 ();
 sg13g2_decap_8 FILLER_31_113 ();
 sg13g2_decap_8 FILLER_31_120 ();
 sg13g2_decap_4 FILLER_31_127 ();
 sg13g2_fill_2 FILLER_31_131 ();
 sg13g2_decap_8 FILLER_31_200 ();
 sg13g2_decap_8 FILLER_31_207 ();
 sg13g2_decap_8 FILLER_31_214 ();
 sg13g2_decap_8 FILLER_31_221 ();
 sg13g2_decap_8 FILLER_31_228 ();
 sg13g2_decap_8 FILLER_31_235 ();
 sg13g2_decap_8 FILLER_31_242 ();
 sg13g2_fill_2 FILLER_31_249 ();
 sg13g2_fill_1 FILLER_31_289 ();
 sg13g2_fill_2 FILLER_31_299 ();
 sg13g2_fill_1 FILLER_31_301 ();
 sg13g2_fill_1 FILLER_31_331 ();
 sg13g2_decap_8 FILLER_31_340 ();
 sg13g2_decap_8 FILLER_31_352 ();
 sg13g2_decap_8 FILLER_31_359 ();
 sg13g2_decap_8 FILLER_31_374 ();
 sg13g2_decap_8 FILLER_31_381 ();
 sg13g2_decap_8 FILLER_31_388 ();
 sg13g2_decap_8 FILLER_31_395 ();
 sg13g2_decap_8 FILLER_31_402 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_8 FILLER_32_84 ();
 sg13g2_decap_8 FILLER_32_91 ();
 sg13g2_fill_2 FILLER_32_98 ();
 sg13g2_fill_1 FILLER_32_100 ();
 sg13g2_fill_2 FILLER_32_106 ();
 sg13g2_decap_8 FILLER_32_134 ();
 sg13g2_fill_1 FILLER_32_141 ();
 sg13g2_decap_8 FILLER_32_177 ();
 sg13g2_fill_1 FILLER_32_184 ();
 sg13g2_decap_8 FILLER_32_194 ();
 sg13g2_decap_8 FILLER_32_201 ();
 sg13g2_decap_8 FILLER_32_208 ();
 sg13g2_decap_8 FILLER_32_215 ();
 sg13g2_fill_2 FILLER_32_222 ();
 sg13g2_fill_1 FILLER_32_224 ();
 sg13g2_decap_8 FILLER_32_228 ();
 sg13g2_decap_8 FILLER_32_235 ();
 sg13g2_fill_1 FILLER_32_305 ();
 sg13g2_fill_2 FILLER_32_343 ();
 sg13g2_fill_1 FILLER_32_345 ();
 sg13g2_fill_2 FILLER_32_353 ();
 sg13g2_decap_8 FILLER_32_381 ();
 sg13g2_decap_8 FILLER_32_388 ();
 sg13g2_decap_8 FILLER_32_395 ();
 sg13g2_decap_8 FILLER_32_402 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_4 FILLER_33_77 ();
 sg13g2_fill_1 FILLER_33_81 ();
 sg13g2_fill_1 FILLER_33_108 ();
 sg13g2_decap_8 FILLER_33_144 ();
 sg13g2_decap_8 FILLER_33_151 ();
 sg13g2_decap_8 FILLER_33_158 ();
 sg13g2_fill_1 FILLER_33_165 ();
 sg13g2_decap_8 FILLER_33_196 ();
 sg13g2_decap_8 FILLER_33_203 ();
 sg13g2_decap_8 FILLER_33_210 ();
 sg13g2_fill_1 FILLER_33_217 ();
 sg13g2_fill_1 FILLER_33_244 ();
 sg13g2_fill_2 FILLER_33_255 ();
 sg13g2_fill_2 FILLER_33_265 ();
 sg13g2_fill_1 FILLER_33_267 ();
 sg13g2_decap_4 FILLER_33_289 ();
 sg13g2_fill_2 FILLER_33_297 ();
 sg13g2_decap_8 FILLER_33_304 ();
 sg13g2_decap_4 FILLER_33_311 ();
 sg13g2_decap_8 FILLER_33_330 ();
 sg13g2_fill_2 FILLER_33_337 ();
 sg13g2_fill_1 FILLER_33_339 ();
 sg13g2_decap_8 FILLER_33_375 ();
 sg13g2_decap_8 FILLER_33_382 ();
 sg13g2_decap_8 FILLER_33_389 ();
 sg13g2_decap_8 FILLER_33_396 ();
 sg13g2_decap_4 FILLER_33_403 ();
 sg13g2_fill_2 FILLER_33_407 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_fill_1 FILLER_34_77 ();
 sg13g2_decap_4 FILLER_34_115 ();
 sg13g2_decap_8 FILLER_34_142 ();
 sg13g2_decap_4 FILLER_34_158 ();
 sg13g2_fill_1 FILLER_34_167 ();
 sg13g2_decap_8 FILLER_34_194 ();
 sg13g2_decap_8 FILLER_34_201 ();
 sg13g2_decap_8 FILLER_34_208 ();
 sg13g2_fill_2 FILLER_34_215 ();
 sg13g2_decap_4 FILLER_34_261 ();
 sg13g2_decap_8 FILLER_34_278 ();
 sg13g2_fill_1 FILLER_34_295 ();
 sg13g2_fill_2 FILLER_34_302 ();
 sg13g2_fill_2 FILLER_34_308 ();
 sg13g2_fill_1 FILLER_34_310 ();
 sg13g2_fill_1 FILLER_34_316 ();
 sg13g2_decap_4 FILLER_34_322 ();
 sg13g2_decap_4 FILLER_34_334 ();
 sg13g2_decap_4 FILLER_34_346 ();
 sg13g2_fill_2 FILLER_34_350 ();
 sg13g2_decap_8 FILLER_34_384 ();
 sg13g2_decap_8 FILLER_34_391 ();
 sg13g2_decap_8 FILLER_34_398 ();
 sg13g2_decap_4 FILLER_34_405 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_fill_2 FILLER_35_84 ();
 sg13g2_fill_1 FILLER_35_86 ();
 sg13g2_decap_8 FILLER_35_117 ();
 sg13g2_decap_4 FILLER_35_124 ();
 sg13g2_fill_1 FILLER_35_132 ();
 sg13g2_fill_2 FILLER_35_199 ();
 sg13g2_fill_1 FILLER_35_201 ();
 sg13g2_decap_8 FILLER_35_210 ();
 sg13g2_decap_8 FILLER_35_217 ();
 sg13g2_decap_4 FILLER_35_227 ();
 sg13g2_fill_1 FILLER_35_247 ();
 sg13g2_fill_2 FILLER_35_258 ();
 sg13g2_decap_8 FILLER_35_265 ();
 sg13g2_decap_8 FILLER_35_272 ();
 sg13g2_decap_8 FILLER_35_279 ();
 sg13g2_decap_8 FILLER_35_286 ();
 sg13g2_fill_2 FILLER_35_293 ();
 sg13g2_fill_2 FILLER_35_306 ();
 sg13g2_fill_2 FILLER_35_313 ();
 sg13g2_decap_8 FILLER_35_320 ();
 sg13g2_fill_2 FILLER_35_327 ();
 sg13g2_decap_8 FILLER_35_355 ();
 sg13g2_fill_1 FILLER_35_362 ();
 sg13g2_fill_2 FILLER_35_368 ();
 sg13g2_fill_1 FILLER_35_370 ();
 sg13g2_fill_2 FILLER_35_375 ();
 sg13g2_decap_8 FILLER_35_386 ();
 sg13g2_decap_8 FILLER_35_393 ();
 sg13g2_decap_8 FILLER_35_400 ();
 sg13g2_fill_2 FILLER_35_407 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_fill_2 FILLER_36_91 ();
 sg13g2_fill_1 FILLER_36_93 ();
 sg13g2_fill_1 FILLER_36_125 ();
 sg13g2_decap_8 FILLER_36_199 ();
 sg13g2_decap_8 FILLER_36_206 ();
 sg13g2_decap_8 FILLER_36_213 ();
 sg13g2_decap_8 FILLER_36_220 ();
 sg13g2_fill_2 FILLER_36_256 ();
 sg13g2_fill_2 FILLER_36_297 ();
 sg13g2_fill_2 FILLER_36_318 ();
 sg13g2_fill_1 FILLER_36_325 ();
 sg13g2_decap_4 FILLER_36_355 ();
 sg13g2_decap_8 FILLER_36_389 ();
 sg13g2_decap_8 FILLER_36_396 ();
 sg13g2_decap_4 FILLER_36_403 ();
 sg13g2_fill_2 FILLER_36_407 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_fill_1 FILLER_37_112 ();
 sg13g2_fill_2 FILLER_37_118 ();
 sg13g2_fill_1 FILLER_37_152 ();
 sg13g2_decap_8 FILLER_37_163 ();
 sg13g2_decap_8 FILLER_37_170 ();
 sg13g2_fill_2 FILLER_37_177 ();
 sg13g2_fill_1 FILLER_37_179 ();
 sg13g2_decap_4 FILLER_37_184 ();
 sg13g2_fill_1 FILLER_37_188 ();
 sg13g2_decap_4 FILLER_37_197 ();
 sg13g2_fill_2 FILLER_37_295 ();
 sg13g2_decap_4 FILLER_37_314 ();
 sg13g2_fill_1 FILLER_37_330 ();
 sg13g2_decap_8 FILLER_37_398 ();
 sg13g2_decap_4 FILLER_37_405 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_8 FILLER_38_56 ();
 sg13g2_decap_8 FILLER_38_63 ();
 sg13g2_decap_8 FILLER_38_70 ();
 sg13g2_decap_8 FILLER_38_77 ();
 sg13g2_decap_4 FILLER_38_84 ();
 sg13g2_fill_1 FILLER_38_88 ();
 sg13g2_fill_2 FILLER_38_99 ();
 sg13g2_fill_2 FILLER_38_127 ();
 sg13g2_fill_2 FILLER_38_133 ();
 sg13g2_fill_1 FILLER_38_135 ();
 sg13g2_decap_8 FILLER_38_171 ();
 sg13g2_fill_2 FILLER_38_178 ();
 sg13g2_fill_1 FILLER_38_180 ();
 sg13g2_fill_2 FILLER_38_215 ();
 sg13g2_fill_1 FILLER_38_217 ();
 sg13g2_decap_4 FILLER_38_244 ();
 sg13g2_fill_1 FILLER_38_293 ();
 sg13g2_fill_1 FILLER_38_298 ();
 sg13g2_fill_1 FILLER_38_303 ();
 sg13g2_fill_1 FILLER_38_309 ();
 sg13g2_decap_8 FILLER_38_349 ();
 sg13g2_decap_8 FILLER_38_356 ();
 sg13g2_fill_2 FILLER_38_367 ();
 sg13g2_fill_1 FILLER_38_369 ();
 sg13g2_decap_8 FILLER_38_388 ();
 sg13g2_decap_8 FILLER_38_395 ();
 sg13g2_decap_8 FILLER_38_402 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_14 ();
 sg13g2_decap_8 FILLER_39_21 ();
 sg13g2_decap_8 FILLER_39_28 ();
 sg13g2_decap_8 FILLER_39_35 ();
 sg13g2_decap_8 FILLER_39_42 ();
 sg13g2_decap_8 FILLER_39_49 ();
 sg13g2_decap_8 FILLER_39_56 ();
 sg13g2_decap_8 FILLER_39_63 ();
 sg13g2_decap_8 FILLER_39_70 ();
 sg13g2_decap_4 FILLER_39_107 ();
 sg13g2_decap_8 FILLER_39_141 ();
 sg13g2_decap_8 FILLER_39_148 ();
 sg13g2_fill_2 FILLER_39_155 ();
 sg13g2_fill_1 FILLER_39_157 ();
 sg13g2_fill_2 FILLER_39_192 ();
 sg13g2_decap_8 FILLER_39_204 ();
 sg13g2_fill_1 FILLER_39_211 ();
 sg13g2_decap_8 FILLER_39_229 ();
 sg13g2_decap_8 FILLER_39_236 ();
 sg13g2_fill_1 FILLER_39_243 ();
 sg13g2_decap_8 FILLER_39_249 ();
 sg13g2_decap_4 FILLER_39_263 ();
 sg13g2_fill_1 FILLER_39_267 ();
 sg13g2_decap_8 FILLER_39_276 ();
 sg13g2_fill_2 FILLER_39_283 ();
 sg13g2_decap_8 FILLER_39_289 ();
 sg13g2_fill_1 FILLER_39_296 ();
 sg13g2_fill_2 FILLER_39_302 ();
 sg13g2_fill_1 FILLER_39_304 ();
 sg13g2_decap_8 FILLER_39_320 ();
 sg13g2_decap_4 FILLER_39_327 ();
 sg13g2_fill_1 FILLER_39_331 ();
 sg13g2_decap_4 FILLER_39_335 ();
 sg13g2_decap_4 FILLER_39_343 ();
 sg13g2_fill_1 FILLER_39_347 ();
 sg13g2_decap_4 FILLER_39_357 ();
 sg13g2_fill_2 FILLER_39_361 ();
 sg13g2_fill_2 FILLER_39_367 ();
 sg13g2_fill_1 FILLER_39_369 ();
 sg13g2_decap_8 FILLER_39_379 ();
 sg13g2_decap_8 FILLER_39_386 ();
 sg13g2_decap_8 FILLER_39_393 ();
 sg13g2_decap_8 FILLER_39_400 ();
 sg13g2_fill_2 FILLER_39_407 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_14 ();
 sg13g2_decap_8 FILLER_40_21 ();
 sg13g2_decap_8 FILLER_40_28 ();
 sg13g2_decap_8 FILLER_40_35 ();
 sg13g2_decap_8 FILLER_40_42 ();
 sg13g2_decap_8 FILLER_40_49 ();
 sg13g2_decap_8 FILLER_40_56 ();
 sg13g2_decap_8 FILLER_40_63 ();
 sg13g2_decap_8 FILLER_40_70 ();
 sg13g2_fill_1 FILLER_40_77 ();
 sg13g2_decap_4 FILLER_40_114 ();
 sg13g2_decap_4 FILLER_40_128 ();
 sg13g2_decap_8 FILLER_40_137 ();
 sg13g2_fill_2 FILLER_40_144 ();
 sg13g2_fill_1 FILLER_40_159 ();
 sg13g2_fill_2 FILLER_40_191 ();
 sg13g2_decap_8 FILLER_40_224 ();
 sg13g2_decap_8 FILLER_40_231 ();
 sg13g2_decap_8 FILLER_40_238 ();
 sg13g2_decap_8 FILLER_40_245 ();
 sg13g2_decap_8 FILLER_40_252 ();
 sg13g2_decap_8 FILLER_40_259 ();
 sg13g2_decap_8 FILLER_40_266 ();
 sg13g2_decap_8 FILLER_40_273 ();
 sg13g2_decap_8 FILLER_40_280 ();
 sg13g2_fill_1 FILLER_40_287 ();
 sg13g2_fill_2 FILLER_40_292 ();
 sg13g2_fill_1 FILLER_40_314 ();
 sg13g2_fill_1 FILLER_40_334 ();
 sg13g2_decap_8 FILLER_40_374 ();
 sg13g2_decap_8 FILLER_40_381 ();
 sg13g2_decap_8 FILLER_40_388 ();
 sg13g2_decap_8 FILLER_40_395 ();
 sg13g2_decap_8 FILLER_40_402 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_8 FILLER_41_14 ();
 sg13g2_decap_8 FILLER_41_21 ();
 sg13g2_decap_8 FILLER_41_28 ();
 sg13g2_decap_8 FILLER_41_35 ();
 sg13g2_decap_8 FILLER_41_42 ();
 sg13g2_decap_8 FILLER_41_49 ();
 sg13g2_decap_8 FILLER_41_56 ();
 sg13g2_decap_8 FILLER_41_63 ();
 sg13g2_decap_8 FILLER_41_70 ();
 sg13g2_fill_1 FILLER_41_77 ();
 sg13g2_fill_1 FILLER_41_108 ();
 sg13g2_decap_4 FILLER_41_115 ();
 sg13g2_fill_2 FILLER_41_149 ();
 sg13g2_fill_2 FILLER_41_156 ();
 sg13g2_fill_1 FILLER_41_158 ();
 sg13g2_decap_4 FILLER_41_163 ();
 sg13g2_decap_8 FILLER_41_176 ();
 sg13g2_fill_2 FILLER_41_191 ();
 sg13g2_fill_1 FILLER_41_216 ();
 sg13g2_decap_8 FILLER_41_235 ();
 sg13g2_decap_8 FILLER_41_242 ();
 sg13g2_decap_8 FILLER_41_249 ();
 sg13g2_decap_4 FILLER_41_256 ();
 sg13g2_decap_8 FILLER_41_266 ();
 sg13g2_fill_1 FILLER_41_273 ();
 sg13g2_decap_4 FILLER_41_279 ();
 sg13g2_decap_4 FILLER_41_317 ();
 sg13g2_fill_1 FILLER_41_321 ();
 sg13g2_fill_1 FILLER_41_330 ();
 sg13g2_fill_2 FILLER_41_340 ();
 sg13g2_decap_8 FILLER_41_383 ();
 sg13g2_decap_8 FILLER_41_390 ();
 sg13g2_decap_8 FILLER_41_397 ();
 sg13g2_decap_4 FILLER_41_404 ();
 sg13g2_fill_1 FILLER_41_408 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_decap_8 FILLER_42_14 ();
 sg13g2_decap_8 FILLER_42_21 ();
 sg13g2_decap_8 FILLER_42_28 ();
 sg13g2_decap_8 FILLER_42_35 ();
 sg13g2_decap_8 FILLER_42_42 ();
 sg13g2_decap_8 FILLER_42_49 ();
 sg13g2_decap_8 FILLER_42_56 ();
 sg13g2_decap_8 FILLER_42_63 ();
 sg13g2_decap_8 FILLER_42_70 ();
 sg13g2_decap_4 FILLER_42_77 ();
 sg13g2_fill_2 FILLER_42_81 ();
 sg13g2_decap_8 FILLER_42_96 ();
 sg13g2_decap_4 FILLER_42_111 ();
 sg13g2_decap_8 FILLER_42_156 ();
 sg13g2_decap_4 FILLER_42_163 ();
 sg13g2_fill_1 FILLER_42_167 ();
 sg13g2_decap_8 FILLER_42_175 ();
 sg13g2_decap_4 FILLER_42_182 ();
 sg13g2_fill_2 FILLER_42_196 ();
 sg13g2_fill_1 FILLER_42_198 ();
 sg13g2_fill_1 FILLER_42_225 ();
 sg13g2_decap_4 FILLER_42_261 ();
 sg13g2_fill_1 FILLER_42_265 ();
 sg13g2_fill_1 FILLER_42_279 ();
 sg13g2_decap_8 FILLER_42_285 ();
 sg13g2_fill_2 FILLER_42_292 ();
 sg13g2_fill_2 FILLER_42_313 ();
 sg13g2_fill_1 FILLER_42_315 ();
 sg13g2_fill_2 FILLER_42_324 ();
 sg13g2_fill_1 FILLER_42_357 ();
 sg13g2_decap_8 FILLER_42_384 ();
 sg13g2_decap_8 FILLER_42_391 ();
 sg13g2_decap_8 FILLER_42_398 ();
 sg13g2_decap_4 FILLER_42_405 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_decap_8 FILLER_43_14 ();
 sg13g2_decap_8 FILLER_43_21 ();
 sg13g2_decap_8 FILLER_43_28 ();
 sg13g2_decap_8 FILLER_43_35 ();
 sg13g2_decap_8 FILLER_43_42 ();
 sg13g2_decap_8 FILLER_43_49 ();
 sg13g2_decap_8 FILLER_43_56 ();
 sg13g2_decap_8 FILLER_43_63 ();
 sg13g2_decap_8 FILLER_43_70 ();
 sg13g2_fill_2 FILLER_43_77 ();
 sg13g2_fill_2 FILLER_43_95 ();
 sg13g2_fill_1 FILLER_43_97 ();
 sg13g2_fill_1 FILLER_43_159 ();
 sg13g2_decap_8 FILLER_43_172 ();
 sg13g2_fill_2 FILLER_43_179 ();
 sg13g2_fill_1 FILLER_43_181 ();
 sg13g2_fill_1 FILLER_43_223 ();
 sg13g2_fill_1 FILLER_43_291 ();
 sg13g2_fill_1 FILLER_43_297 ();
 sg13g2_fill_2 FILLER_43_315 ();
 sg13g2_fill_1 FILLER_43_317 ();
 sg13g2_fill_2 FILLER_43_329 ();
 sg13g2_decap_8 FILLER_43_348 ();
 sg13g2_decap_8 FILLER_43_355 ();
 sg13g2_fill_2 FILLER_43_362 ();
 sg13g2_decap_8 FILLER_43_374 ();
 sg13g2_decap_8 FILLER_43_381 ();
 sg13g2_decap_8 FILLER_43_388 ();
 sg13g2_decap_8 FILLER_43_395 ();
 sg13g2_decap_8 FILLER_43_402 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_decap_8 FILLER_44_14 ();
 sg13g2_decap_8 FILLER_44_21 ();
 sg13g2_decap_8 FILLER_44_28 ();
 sg13g2_decap_8 FILLER_44_35 ();
 sg13g2_decap_8 FILLER_44_42 ();
 sg13g2_decap_8 FILLER_44_49 ();
 sg13g2_decap_8 FILLER_44_56 ();
 sg13g2_decap_8 FILLER_44_63 ();
 sg13g2_decap_4 FILLER_44_70 ();
 sg13g2_fill_1 FILLER_44_74 ();
 sg13g2_fill_1 FILLER_44_123 ();
 sg13g2_decap_8 FILLER_44_129 ();
 sg13g2_decap_4 FILLER_44_136 ();
 sg13g2_fill_1 FILLER_44_140 ();
 sg13g2_decap_4 FILLER_44_156 ();
 sg13g2_fill_2 FILLER_44_165 ();
 sg13g2_fill_1 FILLER_44_167 ();
 sg13g2_fill_2 FILLER_44_174 ();
 sg13g2_fill_1 FILLER_44_176 ();
 sg13g2_fill_2 FILLER_44_184 ();
 sg13g2_fill_1 FILLER_44_186 ();
 sg13g2_decap_8 FILLER_44_207 ();
 sg13g2_decap_4 FILLER_44_219 ();
 sg13g2_fill_1 FILLER_44_223 ();
 sg13g2_fill_2 FILLER_44_265 ();
 sg13g2_decap_8 FILLER_44_282 ();
 sg13g2_decap_8 FILLER_44_289 ();
 sg13g2_fill_1 FILLER_44_296 ();
 sg13g2_decap_4 FILLER_44_301 ();
 sg13g2_decap_4 FILLER_44_311 ();
 sg13g2_fill_1 FILLER_44_315 ();
 sg13g2_fill_2 FILLER_44_324 ();
 sg13g2_decap_8 FILLER_44_332 ();
 sg13g2_fill_2 FILLER_44_339 ();
 sg13g2_decap_8 FILLER_44_358 ();
 sg13g2_decap_8 FILLER_44_365 ();
 sg13g2_decap_8 FILLER_44_372 ();
 sg13g2_decap_8 FILLER_44_379 ();
 sg13g2_decap_8 FILLER_44_386 ();
 sg13g2_decap_8 FILLER_44_393 ();
 sg13g2_decap_8 FILLER_44_400 ();
 sg13g2_fill_2 FILLER_44_407 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_7 ();
 sg13g2_decap_8 FILLER_45_14 ();
 sg13g2_decap_8 FILLER_45_21 ();
 sg13g2_decap_8 FILLER_45_28 ();
 sg13g2_decap_8 FILLER_45_35 ();
 sg13g2_decap_8 FILLER_45_42 ();
 sg13g2_decap_8 FILLER_45_49 ();
 sg13g2_decap_8 FILLER_45_56 ();
 sg13g2_decap_8 FILLER_45_63 ();
 sg13g2_decap_8 FILLER_45_70 ();
 sg13g2_decap_4 FILLER_45_77 ();
 sg13g2_fill_1 FILLER_45_81 ();
 sg13g2_fill_2 FILLER_45_87 ();
 sg13g2_fill_2 FILLER_45_94 ();
 sg13g2_fill_1 FILLER_45_96 ();
 sg13g2_fill_2 FILLER_45_101 ();
 sg13g2_fill_1 FILLER_45_103 ();
 sg13g2_decap_8 FILLER_45_109 ();
 sg13g2_decap_8 FILLER_45_116 ();
 sg13g2_decap_4 FILLER_45_123 ();
 sg13g2_fill_2 FILLER_45_127 ();
 sg13g2_decap_8 FILLER_45_134 ();
 sg13g2_decap_4 FILLER_45_141 ();
 sg13g2_fill_2 FILLER_45_145 ();
 sg13g2_fill_2 FILLER_45_171 ();
 sg13g2_decap_8 FILLER_45_200 ();
 sg13g2_decap_8 FILLER_45_207 ();
 sg13g2_decap_8 FILLER_45_219 ();
 sg13g2_fill_2 FILLER_45_226 ();
 sg13g2_fill_1 FILLER_45_228 ();
 sg13g2_fill_2 FILLER_45_259 ();
 sg13g2_fill_1 FILLER_45_261 ();
 sg13g2_decap_8 FILLER_45_288 ();
 sg13g2_decap_8 FILLER_45_295 ();
 sg13g2_fill_2 FILLER_45_302 ();
 sg13g2_fill_1 FILLER_45_304 ();
 sg13g2_fill_1 FILLER_45_311 ();
 sg13g2_decap_8 FILLER_45_330 ();
 sg13g2_decap_4 FILLER_45_337 ();
 sg13g2_decap_8 FILLER_45_376 ();
 sg13g2_decap_8 FILLER_45_383 ();
 sg13g2_decap_8 FILLER_45_390 ();
 sg13g2_decap_8 FILLER_45_397 ();
 sg13g2_decap_4 FILLER_45_404 ();
 sg13g2_fill_1 FILLER_45_408 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_7 ();
 sg13g2_decap_8 FILLER_46_14 ();
 sg13g2_decap_8 FILLER_46_21 ();
 sg13g2_decap_8 FILLER_46_28 ();
 sg13g2_decap_8 FILLER_46_35 ();
 sg13g2_decap_8 FILLER_46_42 ();
 sg13g2_decap_8 FILLER_46_49 ();
 sg13g2_decap_8 FILLER_46_56 ();
 sg13g2_decap_8 FILLER_46_63 ();
 sg13g2_fill_2 FILLER_46_70 ();
 sg13g2_fill_2 FILLER_46_98 ();
 sg13g2_fill_1 FILLER_46_108 ();
 sg13g2_fill_2 FILLER_46_135 ();
 sg13g2_fill_2 FILLER_46_142 ();
 sg13g2_fill_2 FILLER_46_153 ();
 sg13g2_decap_8 FILLER_46_180 ();
 sg13g2_fill_1 FILLER_46_187 ();
 sg13g2_decap_4 FILLER_46_196 ();
 sg13g2_fill_1 FILLER_46_200 ();
 sg13g2_decap_8 FILLER_46_225 ();
 sg13g2_decap_8 FILLER_46_232 ();
 sg13g2_fill_1 FILLER_46_239 ();
 sg13g2_fill_2 FILLER_46_248 ();
 sg13g2_fill_1 FILLER_46_250 ();
 sg13g2_fill_1 FILLER_46_323 ();
 sg13g2_fill_1 FILLER_46_339 ();
 sg13g2_decap_4 FILLER_46_371 ();
 sg13g2_decap_8 FILLER_46_383 ();
 sg13g2_decap_8 FILLER_46_390 ();
 sg13g2_decap_8 FILLER_46_397 ();
 sg13g2_decap_4 FILLER_46_404 ();
 sg13g2_fill_1 FILLER_46_408 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_7 ();
 sg13g2_decap_8 FILLER_47_14 ();
 sg13g2_decap_8 FILLER_47_21 ();
 sg13g2_decap_8 FILLER_47_28 ();
 sg13g2_decap_8 FILLER_47_35 ();
 sg13g2_decap_8 FILLER_47_42 ();
 sg13g2_decap_8 FILLER_47_49 ();
 sg13g2_decap_8 FILLER_47_56 ();
 sg13g2_decap_4 FILLER_47_63 ();
 sg13g2_fill_1 FILLER_47_67 ();
 sg13g2_fill_2 FILLER_47_99 ();
 sg13g2_fill_1 FILLER_47_101 ();
 sg13g2_fill_1 FILLER_47_108 ();
 sg13g2_fill_1 FILLER_47_115 ();
 sg13g2_fill_1 FILLER_47_158 ();
 sg13g2_decap_8 FILLER_47_173 ();
 sg13g2_fill_2 FILLER_47_180 ();
 sg13g2_fill_1 FILLER_47_182 ();
 sg13g2_fill_2 FILLER_47_258 ();
 sg13g2_fill_1 FILLER_47_281 ();
 sg13g2_fill_2 FILLER_47_303 ();
 sg13g2_decap_8 FILLER_47_355 ();
 sg13g2_decap_4 FILLER_47_362 ();
 sg13g2_decap_8 FILLER_47_371 ();
 sg13g2_decap_8 FILLER_47_378 ();
 sg13g2_decap_8 FILLER_47_385 ();
 sg13g2_decap_8 FILLER_47_392 ();
 sg13g2_decap_8 FILLER_47_399 ();
 sg13g2_fill_2 FILLER_47_406 ();
 sg13g2_fill_1 FILLER_47_408 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_decap_8 FILLER_48_14 ();
 sg13g2_decap_8 FILLER_48_21 ();
 sg13g2_decap_8 FILLER_48_28 ();
 sg13g2_decap_8 FILLER_48_35 ();
 sg13g2_decap_8 FILLER_48_42 ();
 sg13g2_decap_8 FILLER_48_49 ();
 sg13g2_decap_8 FILLER_48_56 ();
 sg13g2_decap_4 FILLER_48_63 ();
 sg13g2_fill_2 FILLER_48_67 ();
 sg13g2_fill_2 FILLER_48_95 ();
 sg13g2_fill_2 FILLER_48_123 ();
 sg13g2_fill_1 FILLER_48_125 ();
 sg13g2_fill_2 FILLER_48_141 ();
 sg13g2_fill_2 FILLER_48_162 ();
 sg13g2_fill_1 FILLER_48_164 ();
 sg13g2_fill_1 FILLER_48_170 ();
 sg13g2_fill_2 FILLER_48_179 ();
 sg13g2_fill_1 FILLER_48_193 ();
 sg13g2_fill_1 FILLER_48_210 ();
 sg13g2_fill_1 FILLER_48_246 ();
 sg13g2_decap_8 FILLER_48_276 ();
 sg13g2_fill_1 FILLER_48_301 ();
 sg13g2_decap_4 FILLER_48_311 ();
 sg13g2_fill_2 FILLER_48_315 ();
 sg13g2_decap_8 FILLER_48_346 ();
 sg13g2_decap_8 FILLER_48_353 ();
 sg13g2_decap_8 FILLER_48_360 ();
 sg13g2_decap_8 FILLER_48_367 ();
 sg13g2_decap_8 FILLER_48_374 ();
 sg13g2_decap_8 FILLER_48_381 ();
 sg13g2_decap_8 FILLER_48_388 ();
 sg13g2_decap_8 FILLER_48_395 ();
 sg13g2_decap_8 FILLER_48_402 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_7 ();
 sg13g2_decap_8 FILLER_49_14 ();
 sg13g2_decap_8 FILLER_49_21 ();
 sg13g2_decap_8 FILLER_49_28 ();
 sg13g2_decap_8 FILLER_49_35 ();
 sg13g2_decap_8 FILLER_49_42 ();
 sg13g2_decap_8 FILLER_49_49 ();
 sg13g2_decap_8 FILLER_49_56 ();
 sg13g2_decap_8 FILLER_49_63 ();
 sg13g2_decap_8 FILLER_49_70 ();
 sg13g2_decap_4 FILLER_49_77 ();
 sg13g2_fill_1 FILLER_49_81 ();
 sg13g2_fill_1 FILLER_49_100 ();
 sg13g2_fill_1 FILLER_49_106 ();
 sg13g2_decap_4 FILLER_49_111 ();
 sg13g2_fill_1 FILLER_49_115 ();
 sg13g2_decap_4 FILLER_49_122 ();
 sg13g2_fill_1 FILLER_49_126 ();
 sg13g2_fill_1 FILLER_49_131 ();
 sg13g2_fill_2 FILLER_49_137 ();
 sg13g2_fill_1 FILLER_49_139 ();
 sg13g2_decap_8 FILLER_49_144 ();
 sg13g2_decap_4 FILLER_49_164 ();
 sg13g2_fill_1 FILLER_49_168 ();
 sg13g2_decap_4 FILLER_49_181 ();
 sg13g2_fill_1 FILLER_49_193 ();
 sg13g2_decap_8 FILLER_49_203 ();
 sg13g2_fill_2 FILLER_49_210 ();
 sg13g2_fill_1 FILLER_49_212 ();
 sg13g2_decap_8 FILLER_49_223 ();
 sg13g2_decap_8 FILLER_49_230 ();
 sg13g2_fill_1 FILLER_49_264 ();
 sg13g2_fill_2 FILLER_49_271 ();
 sg13g2_decap_8 FILLER_49_281 ();
 sg13g2_decap_8 FILLER_49_288 ();
 sg13g2_fill_1 FILLER_49_295 ();
 sg13g2_fill_2 FILLER_49_349 ();
 sg13g2_decap_4 FILLER_49_354 ();
 sg13g2_fill_2 FILLER_49_358 ();
 sg13g2_decap_8 FILLER_49_368 ();
 sg13g2_decap_8 FILLER_49_375 ();
 sg13g2_decap_8 FILLER_49_382 ();
 sg13g2_decap_8 FILLER_49_389 ();
 sg13g2_decap_8 FILLER_49_396 ();
 sg13g2_decap_4 FILLER_49_403 ();
 sg13g2_fill_2 FILLER_49_407 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_8 FILLER_50_7 ();
 sg13g2_decap_8 FILLER_50_14 ();
 sg13g2_decap_8 FILLER_50_21 ();
 sg13g2_decap_8 FILLER_50_28 ();
 sg13g2_decap_8 FILLER_50_35 ();
 sg13g2_decap_8 FILLER_50_42 ();
 sg13g2_decap_8 FILLER_50_49 ();
 sg13g2_decap_8 FILLER_50_56 ();
 sg13g2_decap_8 FILLER_50_63 ();
 sg13g2_decap_4 FILLER_50_70 ();
 sg13g2_fill_1 FILLER_50_100 ();
 sg13g2_decap_4 FILLER_50_127 ();
 sg13g2_decap_4 FILLER_50_163 ();
 sg13g2_decap_8 FILLER_50_208 ();
 sg13g2_decap_8 FILLER_50_215 ();
 sg13g2_fill_2 FILLER_50_222 ();
 sg13g2_decap_8 FILLER_50_232 ();
 sg13g2_decap_8 FILLER_50_239 ();
 sg13g2_fill_2 FILLER_50_246 ();
 sg13g2_fill_1 FILLER_50_248 ();
 sg13g2_fill_2 FILLER_50_252 ();
 sg13g2_fill_1 FILLER_50_254 ();
 sg13g2_decap_8 FILLER_50_268 ();
 sg13g2_decap_8 FILLER_50_280 ();
 sg13g2_fill_1 FILLER_50_287 ();
 sg13g2_decap_8 FILLER_50_298 ();
 sg13g2_fill_1 FILLER_50_305 ();
 sg13g2_fill_1 FILLER_50_319 ();
 sg13g2_decap_8 FILLER_50_382 ();
 sg13g2_decap_8 FILLER_50_389 ();
 sg13g2_decap_8 FILLER_50_396 ();
 sg13g2_decap_4 FILLER_50_403 ();
 sg13g2_fill_2 FILLER_50_407 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_decap_8 FILLER_51_7 ();
 sg13g2_decap_8 FILLER_51_14 ();
 sg13g2_decap_8 FILLER_51_21 ();
 sg13g2_decap_8 FILLER_51_28 ();
 sg13g2_decap_8 FILLER_51_35 ();
 sg13g2_decap_8 FILLER_51_42 ();
 sg13g2_decap_8 FILLER_51_49 ();
 sg13g2_decap_8 FILLER_51_56 ();
 sg13g2_decap_8 FILLER_51_63 ();
 sg13g2_decap_4 FILLER_51_70 ();
 sg13g2_fill_1 FILLER_51_74 ();
 sg13g2_decap_8 FILLER_51_106 ();
 sg13g2_fill_1 FILLER_51_113 ();
 sg13g2_decap_8 FILLER_51_123 ();
 sg13g2_decap_8 FILLER_51_130 ();
 sg13g2_fill_2 FILLER_51_137 ();
 sg13g2_decap_8 FILLER_51_234 ();
 sg13g2_fill_2 FILLER_51_241 ();
 sg13g2_fill_1 FILLER_51_243 ();
 sg13g2_decap_8 FILLER_51_278 ();
 sg13g2_fill_2 FILLER_51_285 ();
 sg13g2_decap_4 FILLER_51_305 ();
 sg13g2_fill_1 FILLER_51_309 ();
 sg13g2_decap_8 FILLER_51_315 ();
 sg13g2_decap_4 FILLER_51_345 ();
 sg13g2_fill_2 FILLER_51_349 ();
 sg13g2_decap_8 FILLER_51_377 ();
 sg13g2_decap_8 FILLER_51_384 ();
 sg13g2_decap_8 FILLER_51_391 ();
 sg13g2_decap_8 FILLER_51_398 ();
 sg13g2_decap_4 FILLER_51_405 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_decap_8 FILLER_52_7 ();
 sg13g2_decap_8 FILLER_52_14 ();
 sg13g2_decap_8 FILLER_52_21 ();
 sg13g2_decap_8 FILLER_52_28 ();
 sg13g2_decap_8 FILLER_52_35 ();
 sg13g2_decap_8 FILLER_52_42 ();
 sg13g2_decap_8 FILLER_52_49 ();
 sg13g2_decap_8 FILLER_52_56 ();
 sg13g2_decap_8 FILLER_52_63 ();
 sg13g2_decap_8 FILLER_52_70 ();
 sg13g2_decap_8 FILLER_52_77 ();
 sg13g2_fill_1 FILLER_52_84 ();
 sg13g2_fill_1 FILLER_52_94 ();
 sg13g2_decap_4 FILLER_52_99 ();
 sg13g2_decap_4 FILLER_52_111 ();
 sg13g2_fill_2 FILLER_52_115 ();
 sg13g2_decap_4 FILLER_52_126 ();
 sg13g2_fill_1 FILLER_52_130 ();
 sg13g2_fill_2 FILLER_52_169 ();
 sg13g2_decap_8 FILLER_52_177 ();
 sg13g2_fill_1 FILLER_52_184 ();
 sg13g2_fill_1 FILLER_52_194 ();
 sg13g2_fill_2 FILLER_52_233 ();
 sg13g2_decap_8 FILLER_52_264 ();
 sg13g2_decap_4 FILLER_52_271 ();
 sg13g2_fill_1 FILLER_52_275 ();
 sg13g2_decap_4 FILLER_52_279 ();
 sg13g2_decap_8 FILLER_52_296 ();
 sg13g2_decap_8 FILLER_52_303 ();
 sg13g2_fill_1 FILLER_52_327 ();
 sg13g2_fill_1 FILLER_52_354 ();
 sg13g2_decap_4 FILLER_52_364 ();
 sg13g2_decap_8 FILLER_52_400 ();
 sg13g2_fill_2 FILLER_52_407 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_decap_8 FILLER_53_7 ();
 sg13g2_decap_8 FILLER_53_14 ();
 sg13g2_decap_8 FILLER_53_21 ();
 sg13g2_decap_8 FILLER_53_28 ();
 sg13g2_decap_8 FILLER_53_35 ();
 sg13g2_decap_8 FILLER_53_42 ();
 sg13g2_decap_8 FILLER_53_49 ();
 sg13g2_decap_8 FILLER_53_56 ();
 sg13g2_decap_8 FILLER_53_63 ();
 sg13g2_decap_8 FILLER_53_70 ();
 sg13g2_decap_8 FILLER_53_77 ();
 sg13g2_decap_8 FILLER_53_84 ();
 sg13g2_fill_2 FILLER_53_91 ();
 sg13g2_fill_1 FILLER_53_93 ();
 sg13g2_decap_4 FILLER_53_98 ();
 sg13g2_fill_2 FILLER_53_102 ();
 sg13g2_fill_2 FILLER_53_136 ();
 sg13g2_fill_2 FILLER_53_143 ();
 sg13g2_fill_1 FILLER_53_145 ();
 sg13g2_decap_8 FILLER_53_177 ();
 sg13g2_decap_8 FILLER_53_184 ();
 sg13g2_decap_4 FILLER_53_191 ();
 sg13g2_fill_1 FILLER_53_195 ();
 sg13g2_decap_4 FILLER_53_210 ();
 sg13g2_decap_4 FILLER_53_234 ();
 sg13g2_fill_2 FILLER_53_264 ();
 sg13g2_fill_1 FILLER_53_266 ();
 sg13g2_decap_8 FILLER_53_319 ();
 sg13g2_decap_8 FILLER_53_326 ();
 sg13g2_decap_8 FILLER_53_333 ();
 sg13g2_fill_2 FILLER_53_340 ();
 sg13g2_fill_1 FILLER_53_342 ();
 sg13g2_decap_8 FILLER_53_347 ();
 sg13g2_fill_1 FILLER_53_354 ();
 sg13g2_decap_8 FILLER_53_397 ();
 sg13g2_decap_4 FILLER_53_404 ();
 sg13g2_fill_1 FILLER_53_408 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_decap_8 FILLER_54_7 ();
 sg13g2_decap_8 FILLER_54_14 ();
 sg13g2_decap_8 FILLER_54_21 ();
 sg13g2_decap_8 FILLER_54_28 ();
 sg13g2_decap_8 FILLER_54_35 ();
 sg13g2_decap_8 FILLER_54_42 ();
 sg13g2_decap_8 FILLER_54_49 ();
 sg13g2_decap_8 FILLER_54_56 ();
 sg13g2_decap_8 FILLER_54_63 ();
 sg13g2_decap_4 FILLER_54_70 ();
 sg13g2_fill_2 FILLER_54_74 ();
 sg13g2_decap_8 FILLER_54_138 ();
 sg13g2_decap_8 FILLER_54_145 ();
 sg13g2_fill_1 FILLER_54_152 ();
 sg13g2_fill_2 FILLER_54_164 ();
 sg13g2_fill_1 FILLER_54_166 ();
 sg13g2_decap_8 FILLER_54_193 ();
 sg13g2_decap_4 FILLER_54_200 ();
 sg13g2_fill_1 FILLER_54_204 ();
 sg13g2_decap_4 FILLER_54_231 ();
 sg13g2_decap_8 FILLER_54_240 ();
 sg13g2_decap_8 FILLER_54_247 ();
 sg13g2_decap_4 FILLER_54_254 ();
 sg13g2_fill_1 FILLER_54_258 ();
 sg13g2_fill_2 FILLER_54_266 ();
 sg13g2_fill_1 FILLER_54_268 ();
 sg13g2_fill_2 FILLER_54_282 ();
 sg13g2_decap_8 FILLER_54_290 ();
 sg13g2_fill_1 FILLER_54_297 ();
 sg13g2_fill_1 FILLER_54_301 ();
 sg13g2_decap_8 FILLER_54_313 ();
 sg13g2_decap_8 FILLER_54_320 ();
 sg13g2_fill_2 FILLER_54_327 ();
 sg13g2_fill_1 FILLER_54_329 ();
 sg13g2_decap_8 FILLER_54_336 ();
 sg13g2_decap_4 FILLER_54_343 ();
 sg13g2_fill_1 FILLER_54_347 ();
 sg13g2_decap_8 FILLER_54_356 ();
 sg13g2_fill_2 FILLER_54_363 ();
 sg13g2_fill_1 FILLER_54_365 ();
 sg13g2_decap_4 FILLER_54_403 ();
 sg13g2_fill_2 FILLER_54_407 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_decap_8 FILLER_55_7 ();
 sg13g2_decap_8 FILLER_55_14 ();
 sg13g2_decap_8 FILLER_55_21 ();
 sg13g2_decap_8 FILLER_55_28 ();
 sg13g2_decap_8 FILLER_55_35 ();
 sg13g2_decap_8 FILLER_55_42 ();
 sg13g2_decap_8 FILLER_55_49 ();
 sg13g2_decap_8 FILLER_55_56 ();
 sg13g2_decap_8 FILLER_55_63 ();
 sg13g2_decap_4 FILLER_55_70 ();
 sg13g2_fill_2 FILLER_55_74 ();
 sg13g2_fill_2 FILLER_55_112 ();
 sg13g2_fill_1 FILLER_55_114 ();
 sg13g2_decap_8 FILLER_55_134 ();
 sg13g2_fill_2 FILLER_55_141 ();
 sg13g2_decap_8 FILLER_55_149 ();
 sg13g2_fill_2 FILLER_55_156 ();
 sg13g2_fill_1 FILLER_55_158 ();
 sg13g2_fill_2 FILLER_55_195 ();
 sg13g2_fill_1 FILLER_55_197 ();
 sg13g2_decap_4 FILLER_55_203 ();
 sg13g2_fill_1 FILLER_55_207 ();
 sg13g2_decap_4 FILLER_55_234 ();
 sg13g2_fill_2 FILLER_55_238 ();
 sg13g2_decap_8 FILLER_55_279 ();
 sg13g2_fill_1 FILLER_55_286 ();
 sg13g2_fill_2 FILLER_55_292 ();
 sg13g2_fill_2 FILLER_55_317 ();
 sg13g2_fill_1 FILLER_55_319 ();
 sg13g2_fill_1 FILLER_55_360 ();
 sg13g2_decap_8 FILLER_55_366 ();
 sg13g2_fill_2 FILLER_55_373 ();
 sg13g2_fill_2 FILLER_55_385 ();
 sg13g2_decap_8 FILLER_55_400 ();
 sg13g2_fill_2 FILLER_55_407 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_decap_8 FILLER_56_7 ();
 sg13g2_decap_8 FILLER_56_14 ();
 sg13g2_decap_8 FILLER_56_21 ();
 sg13g2_decap_8 FILLER_56_28 ();
 sg13g2_decap_8 FILLER_56_35 ();
 sg13g2_decap_8 FILLER_56_42 ();
 sg13g2_decap_8 FILLER_56_49 ();
 sg13g2_decap_8 FILLER_56_56 ();
 sg13g2_decap_8 FILLER_56_63 ();
 sg13g2_decap_8 FILLER_56_70 ();
 sg13g2_decap_8 FILLER_56_77 ();
 sg13g2_fill_2 FILLER_56_84 ();
 sg13g2_fill_1 FILLER_56_86 ();
 sg13g2_decap_8 FILLER_56_105 ();
 sg13g2_fill_2 FILLER_56_112 ();
 sg13g2_fill_1 FILLER_56_114 ();
 sg13g2_fill_2 FILLER_56_147 ();
 sg13g2_decap_8 FILLER_56_159 ();
 sg13g2_fill_2 FILLER_56_166 ();
 sg13g2_decap_8 FILLER_56_176 ();
 sg13g2_decap_4 FILLER_56_230 ();
 sg13g2_decap_8 FILLER_56_247 ();
 sg13g2_decap_4 FILLER_56_254 ();
 sg13g2_fill_2 FILLER_56_258 ();
 sg13g2_decap_8 FILLER_56_288 ();
 sg13g2_fill_2 FILLER_56_295 ();
 sg13g2_fill_2 FILLER_56_382 ();
 sg13g2_fill_2 FILLER_56_407 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_decap_8 FILLER_57_7 ();
 sg13g2_decap_8 FILLER_57_14 ();
 sg13g2_decap_8 FILLER_57_21 ();
 sg13g2_decap_8 FILLER_57_28 ();
 sg13g2_decap_8 FILLER_57_35 ();
 sg13g2_decap_8 FILLER_57_42 ();
 sg13g2_decap_8 FILLER_57_49 ();
 sg13g2_decap_8 FILLER_57_56 ();
 sg13g2_decap_8 FILLER_57_63 ();
 sg13g2_decap_8 FILLER_57_70 ();
 sg13g2_decap_8 FILLER_57_77 ();
 sg13g2_decap_8 FILLER_57_84 ();
 sg13g2_fill_2 FILLER_57_91 ();
 sg13g2_fill_1 FILLER_57_97 ();
 sg13g2_decap_8 FILLER_57_107 ();
 sg13g2_fill_2 FILLER_57_114 ();
 sg13g2_decap_4 FILLER_57_147 ();
 sg13g2_fill_1 FILLER_57_156 ();
 sg13g2_decap_4 FILLER_57_161 ();
 sg13g2_fill_2 FILLER_57_165 ();
 sg13g2_decap_8 FILLER_57_173 ();
 sg13g2_decap_4 FILLER_57_180 ();
 sg13g2_fill_1 FILLER_57_184 ();
 sg13g2_fill_2 FILLER_57_199 ();
 sg13g2_decap_8 FILLER_57_209 ();
 sg13g2_decap_8 FILLER_57_216 ();
 sg13g2_decap_4 FILLER_57_223 ();
 sg13g2_fill_1 FILLER_57_227 ();
 sg13g2_fill_1 FILLER_57_267 ();
 sg13g2_decap_4 FILLER_57_284 ();
 sg13g2_fill_2 FILLER_57_288 ();
 sg13g2_fill_2 FILLER_57_407 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_decap_8 FILLER_58_7 ();
 sg13g2_decap_8 FILLER_58_14 ();
 sg13g2_decap_8 FILLER_58_21 ();
 sg13g2_decap_8 FILLER_58_28 ();
 sg13g2_decap_8 FILLER_58_35 ();
 sg13g2_decap_8 FILLER_58_42 ();
 sg13g2_decap_8 FILLER_58_49 ();
 sg13g2_decap_8 FILLER_58_56 ();
 sg13g2_decap_8 FILLER_58_63 ();
 sg13g2_decap_8 FILLER_58_70 ();
 sg13g2_decap_8 FILLER_58_77 ();
 sg13g2_decap_4 FILLER_58_84 ();
 sg13g2_fill_1 FILLER_58_88 ();
 sg13g2_decap_8 FILLER_58_120 ();
 sg13g2_fill_2 FILLER_58_140 ();
 sg13g2_decap_8 FILLER_58_176 ();
 sg13g2_fill_2 FILLER_58_183 ();
 sg13g2_decap_4 FILLER_58_211 ();
 sg13g2_fill_2 FILLER_58_215 ();
 sg13g2_decap_8 FILLER_58_225 ();
 sg13g2_decap_8 FILLER_58_232 ();
 sg13g2_decap_4 FILLER_58_239 ();
 sg13g2_fill_2 FILLER_58_243 ();
 sg13g2_decap_8 FILLER_58_253 ();
 sg13g2_fill_2 FILLER_58_260 ();
 sg13g2_fill_1 FILLER_58_262 ();
 sg13g2_decap_4 FILLER_58_300 ();
 sg13g2_decap_8 FILLER_58_336 ();
 sg13g2_decap_8 FILLER_58_343 ();
 sg13g2_decap_8 FILLER_58_350 ();
 sg13g2_fill_2 FILLER_58_357 ();
 sg13g2_fill_1 FILLER_58_362 ();
 sg13g2_fill_1 FILLER_58_368 ();
 sg13g2_fill_2 FILLER_58_377 ();
 sg13g2_fill_1 FILLER_58_384 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_decap_8 FILLER_59_7 ();
 sg13g2_decap_8 FILLER_59_14 ();
 sg13g2_decap_8 FILLER_59_21 ();
 sg13g2_decap_8 FILLER_59_28 ();
 sg13g2_decap_8 FILLER_59_35 ();
 sg13g2_decap_8 FILLER_59_42 ();
 sg13g2_decap_8 FILLER_59_49 ();
 sg13g2_decap_8 FILLER_59_56 ();
 sg13g2_decap_8 FILLER_59_63 ();
 sg13g2_decap_4 FILLER_59_70 ();
 sg13g2_fill_2 FILLER_59_74 ();
 sg13g2_fill_2 FILLER_59_102 ();
 sg13g2_fill_2 FILLER_59_110 ();
 sg13g2_decap_8 FILLER_59_128 ();
 sg13g2_decap_8 FILLER_59_135 ();
 sg13g2_fill_2 FILLER_59_142 ();
 sg13g2_fill_1 FILLER_59_144 ();
 sg13g2_fill_2 FILLER_59_153 ();
 sg13g2_fill_1 FILLER_59_155 ();
 sg13g2_fill_2 FILLER_59_161 ();
 sg13g2_fill_1 FILLER_59_163 ();
 sg13g2_decap_4 FILLER_59_181 ();
 sg13g2_decap_4 FILLER_59_205 ();
 sg13g2_decap_8 FILLER_59_243 ();
 sg13g2_fill_2 FILLER_59_250 ();
 sg13g2_fill_1 FILLER_59_252 ();
 sg13g2_decap_8 FILLER_59_303 ();
 sg13g2_decap_4 FILLER_59_310 ();
 sg13g2_fill_1 FILLER_59_314 ();
 sg13g2_decap_8 FILLER_59_330 ();
 sg13g2_decap_4 FILLER_59_337 ();
 sg13g2_decap_8 FILLER_59_363 ();
 sg13g2_decap_4 FILLER_59_370 ();
 sg13g2_fill_1 FILLER_59_374 ();
 sg13g2_decap_8 FILLER_59_379 ();
 sg13g2_fill_2 FILLER_59_386 ();
 sg13g2_fill_2 FILLER_59_406 ();
 sg13g2_fill_1 FILLER_59_408 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_decap_8 FILLER_60_7 ();
 sg13g2_decap_8 FILLER_60_14 ();
 sg13g2_decap_8 FILLER_60_21 ();
 sg13g2_decap_8 FILLER_60_28 ();
 sg13g2_decap_8 FILLER_60_35 ();
 sg13g2_decap_8 FILLER_60_42 ();
 sg13g2_decap_8 FILLER_60_49 ();
 sg13g2_decap_8 FILLER_60_56 ();
 sg13g2_decap_8 FILLER_60_63 ();
 sg13g2_decap_8 FILLER_60_70 ();
 sg13g2_fill_1 FILLER_60_77 ();
 sg13g2_fill_2 FILLER_60_144 ();
 sg13g2_fill_1 FILLER_60_198 ();
 sg13g2_decap_8 FILLER_60_235 ();
 sg13g2_decap_8 FILLER_60_242 ();
 sg13g2_decap_8 FILLER_60_249 ();
 sg13g2_decap_4 FILLER_60_256 ();
 sg13g2_fill_1 FILLER_60_264 ();
 sg13g2_fill_2 FILLER_60_272 ();
 sg13g2_fill_1 FILLER_60_293 ();
 sg13g2_decap_8 FILLER_60_297 ();
 sg13g2_fill_2 FILLER_60_304 ();
 sg13g2_fill_2 FILLER_60_319 ();
 sg13g2_fill_1 FILLER_60_321 ();
 sg13g2_fill_2 FILLER_60_330 ();
 sg13g2_fill_1 FILLER_60_335 ();
 sg13g2_fill_2 FILLER_60_341 ();
 sg13g2_fill_1 FILLER_60_343 ();
 sg13g2_fill_1 FILLER_60_353 ();
 sg13g2_fill_2 FILLER_60_374 ();
 sg13g2_fill_1 FILLER_60_376 ();
 sg13g2_fill_2 FILLER_60_385 ();
 sg13g2_decap_4 FILLER_60_405 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_decap_8 FILLER_61_7 ();
 sg13g2_decap_8 FILLER_61_14 ();
 sg13g2_decap_8 FILLER_61_21 ();
 sg13g2_decap_8 FILLER_61_28 ();
 sg13g2_decap_8 FILLER_61_35 ();
 sg13g2_decap_8 FILLER_61_42 ();
 sg13g2_decap_8 FILLER_61_49 ();
 sg13g2_decap_8 FILLER_61_56 ();
 sg13g2_decap_8 FILLER_61_63 ();
 sg13g2_decap_4 FILLER_61_70 ();
 sg13g2_fill_1 FILLER_61_74 ();
 sg13g2_fill_2 FILLER_61_110 ();
 sg13g2_fill_2 FILLER_61_142 ();
 sg13g2_fill_2 FILLER_61_149 ();
 sg13g2_fill_1 FILLER_61_151 ();
 sg13g2_decap_8 FILLER_61_161 ();
 sg13g2_fill_2 FILLER_61_177 ();
 sg13g2_fill_1 FILLER_61_213 ();
 sg13g2_decap_8 FILLER_61_240 ();
 sg13g2_fill_2 FILLER_61_247 ();
 sg13g2_fill_1 FILLER_61_249 ();
 sg13g2_fill_1 FILLER_61_276 ();
 sg13g2_decap_4 FILLER_61_283 ();
 sg13g2_fill_2 FILLER_61_326 ();
 sg13g2_fill_1 FILLER_61_353 ();
 sg13g2_fill_1 FILLER_61_373 ();
 sg13g2_fill_2 FILLER_61_407 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_decap_8 FILLER_62_7 ();
 sg13g2_decap_8 FILLER_62_14 ();
 sg13g2_decap_8 FILLER_62_21 ();
 sg13g2_decap_8 FILLER_62_28 ();
 sg13g2_decap_8 FILLER_62_35 ();
 sg13g2_decap_8 FILLER_62_42 ();
 sg13g2_decap_8 FILLER_62_49 ();
 sg13g2_decap_8 FILLER_62_56 ();
 sg13g2_decap_8 FILLER_62_63 ();
 sg13g2_decap_8 FILLER_62_70 ();
 sg13g2_decap_8 FILLER_62_77 ();
 sg13g2_decap_8 FILLER_62_84 ();
 sg13g2_fill_2 FILLER_62_91 ();
 sg13g2_fill_1 FILLER_62_93 ();
 sg13g2_decap_8 FILLER_62_98 ();
 sg13g2_decap_8 FILLER_62_105 ();
 sg13g2_decap_8 FILLER_62_112 ();
 sg13g2_fill_2 FILLER_62_119 ();
 sg13g2_fill_1 FILLER_62_121 ();
 sg13g2_fill_2 FILLER_62_127 ();
 sg13g2_decap_4 FILLER_62_133 ();
 sg13g2_fill_1 FILLER_62_162 ();
 sg13g2_decap_8 FILLER_62_169 ();
 sg13g2_decap_8 FILLER_62_176 ();
 sg13g2_decap_8 FILLER_62_183 ();
 sg13g2_fill_2 FILLER_62_190 ();
 sg13g2_fill_1 FILLER_62_192 ();
 sg13g2_decap_8 FILLER_62_197 ();
 sg13g2_decap_8 FILLER_62_204 ();
 sg13g2_decap_8 FILLER_62_211 ();
 sg13g2_decap_8 FILLER_62_218 ();
 sg13g2_decap_8 FILLER_62_225 ();
 sg13g2_decap_8 FILLER_62_232 ();
 sg13g2_decap_8 FILLER_62_239 ();
 sg13g2_decap_8 FILLER_62_246 ();
 sg13g2_fill_2 FILLER_62_253 ();
 sg13g2_fill_1 FILLER_62_255 ();
 sg13g2_fill_2 FILLER_62_282 ();
 sg13g2_decap_4 FILLER_62_287 ();
 sg13g2_fill_2 FILLER_62_291 ();
 sg13g2_fill_2 FILLER_62_319 ();
 sg13g2_fill_2 FILLER_62_350 ();
 sg13g2_fill_1 FILLER_62_352 ();
 sg13g2_decap_4 FILLER_62_388 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_decap_8 FILLER_63_7 ();
 sg13g2_decap_8 FILLER_63_14 ();
 sg13g2_decap_8 FILLER_63_21 ();
 sg13g2_decap_8 FILLER_63_28 ();
 sg13g2_decap_8 FILLER_63_35 ();
 sg13g2_decap_8 FILLER_63_42 ();
 sg13g2_decap_8 FILLER_63_49 ();
 sg13g2_decap_8 FILLER_63_56 ();
 sg13g2_decap_8 FILLER_63_63 ();
 sg13g2_decap_8 FILLER_63_70 ();
 sg13g2_fill_2 FILLER_63_77 ();
 sg13g2_decap_4 FILLER_63_111 ();
 sg13g2_fill_1 FILLER_63_121 ();
 sg13g2_decap_4 FILLER_63_128 ();
 sg13g2_fill_2 FILLER_63_138 ();
 sg13g2_fill_1 FILLER_63_140 ();
 sg13g2_fill_1 FILLER_63_181 ();
 sg13g2_fill_1 FILLER_63_192 ();
 sg13g2_decap_8 FILLER_63_202 ();
 sg13g2_fill_1 FILLER_63_209 ();
 sg13g2_fill_2 FILLER_63_218 ();
 sg13g2_fill_1 FILLER_63_220 ();
 sg13g2_decap_4 FILLER_63_224 ();
 sg13g2_fill_1 FILLER_63_234 ();
 sg13g2_fill_1 FILLER_63_261 ();
 sg13g2_decap_8 FILLER_63_265 ();
 sg13g2_fill_2 FILLER_63_272 ();
 sg13g2_decap_8 FILLER_63_300 ();
 sg13g2_decap_4 FILLER_63_307 ();
 sg13g2_fill_2 FILLER_63_324 ();
 sg13g2_decap_8 FILLER_63_349 ();
 sg13g2_fill_2 FILLER_63_356 ();
 sg13g2_fill_1 FILLER_63_358 ();
 sg13g2_fill_1 FILLER_63_369 ();
 sg13g2_decap_8 FILLER_63_378 ();
 sg13g2_decap_8 FILLER_63_385 ();
 sg13g2_fill_2 FILLER_63_392 ();
 sg13g2_decap_8 FILLER_63_399 ();
 sg13g2_fill_2 FILLER_63_406 ();
 sg13g2_fill_1 FILLER_63_408 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_8 FILLER_64_7 ();
 sg13g2_decap_8 FILLER_64_14 ();
 sg13g2_decap_8 FILLER_64_21 ();
 sg13g2_decap_8 FILLER_64_28 ();
 sg13g2_decap_8 FILLER_64_35 ();
 sg13g2_decap_8 FILLER_64_42 ();
 sg13g2_decap_8 FILLER_64_49 ();
 sg13g2_decap_8 FILLER_64_56 ();
 sg13g2_decap_8 FILLER_64_63 ();
 sg13g2_decap_8 FILLER_64_70 ();
 sg13g2_fill_1 FILLER_64_77 ();
 sg13g2_fill_1 FILLER_64_134 ();
 sg13g2_fill_2 FILLER_64_150 ();
 sg13g2_fill_1 FILLER_64_152 ();
 sg13g2_fill_1 FILLER_64_179 ();
 sg13g2_decap_4 FILLER_64_211 ();
 sg13g2_fill_2 FILLER_64_299 ();
 sg13g2_decap_8 FILLER_64_307 ();
 sg13g2_fill_2 FILLER_64_314 ();
 sg13g2_fill_1 FILLER_64_316 ();
 sg13g2_fill_2 FILLER_64_322 ();
 sg13g2_fill_1 FILLER_64_324 ();
 sg13g2_decap_8 FILLER_64_338 ();
 sg13g2_decap_8 FILLER_64_345 ();
 sg13g2_fill_2 FILLER_64_352 ();
 sg13g2_fill_1 FILLER_64_354 ();
 sg13g2_fill_2 FILLER_64_378 ();
 sg13g2_fill_1 FILLER_64_380 ();
 sg13g2_decap_8 FILLER_64_394 ();
 sg13g2_decap_8 FILLER_64_401 ();
 sg13g2_fill_1 FILLER_64_408 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_8 FILLER_65_7 ();
 sg13g2_decap_8 FILLER_65_14 ();
 sg13g2_decap_8 FILLER_65_21 ();
 sg13g2_decap_8 FILLER_65_28 ();
 sg13g2_decap_8 FILLER_65_35 ();
 sg13g2_decap_8 FILLER_65_42 ();
 sg13g2_decap_8 FILLER_65_49 ();
 sg13g2_decap_8 FILLER_65_56 ();
 sg13g2_decap_8 FILLER_65_63 ();
 sg13g2_decap_8 FILLER_65_70 ();
 sg13g2_decap_8 FILLER_65_77 ();
 sg13g2_decap_4 FILLER_65_84 ();
 sg13g2_decap_8 FILLER_65_121 ();
 sg13g2_fill_2 FILLER_65_128 ();
 sg13g2_fill_2 FILLER_65_149 ();
 sg13g2_fill_1 FILLER_65_151 ();
 sg13g2_decap_8 FILLER_65_156 ();
 sg13g2_decap_8 FILLER_65_163 ();
 sg13g2_decap_8 FILLER_65_170 ();
 sg13g2_decap_4 FILLER_65_177 ();
 sg13g2_fill_1 FILLER_65_181 ();
 sg13g2_decap_8 FILLER_65_187 ();
 sg13g2_fill_1 FILLER_65_194 ();
 sg13g2_fill_2 FILLER_65_229 ();
 sg13g2_fill_1 FILLER_65_231 ();
 sg13g2_decap_8 FILLER_65_250 ();
 sg13g2_decap_4 FILLER_65_257 ();
 sg13g2_fill_2 FILLER_65_261 ();
 sg13g2_fill_2 FILLER_65_283 ();
 sg13g2_decap_4 FILLER_65_311 ();
 sg13g2_fill_1 FILLER_65_315 ();
 sg13g2_fill_2 FILLER_65_337 ();
 sg13g2_fill_1 FILLER_65_339 ();
 sg13g2_decap_8 FILLER_65_366 ();
 sg13g2_decap_8 FILLER_65_373 ();
 sg13g2_decap_8 FILLER_65_380 ();
 sg13g2_fill_2 FILLER_65_387 ();
 sg13g2_decap_8 FILLER_65_393 ();
 sg13g2_decap_8 FILLER_65_400 ();
 sg13g2_fill_2 FILLER_65_407 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_8 FILLER_66_7 ();
 sg13g2_decap_8 FILLER_66_14 ();
 sg13g2_decap_8 FILLER_66_21 ();
 sg13g2_decap_8 FILLER_66_28 ();
 sg13g2_decap_8 FILLER_66_35 ();
 sg13g2_decap_8 FILLER_66_42 ();
 sg13g2_decap_8 FILLER_66_49 ();
 sg13g2_decap_8 FILLER_66_56 ();
 sg13g2_decap_8 FILLER_66_63 ();
 sg13g2_decap_4 FILLER_66_70 ();
 sg13g2_fill_1 FILLER_66_74 ();
 sg13g2_decap_8 FILLER_66_105 ();
 sg13g2_fill_2 FILLER_66_112 ();
 sg13g2_fill_1 FILLER_66_144 ();
 sg13g2_fill_2 FILLER_66_153 ();
 sg13g2_fill_1 FILLER_66_155 ();
 sg13g2_decap_4 FILLER_66_162 ();
 sg13g2_fill_1 FILLER_66_166 ();
 sg13g2_decap_4 FILLER_66_183 ();
 sg13g2_fill_2 FILLER_66_187 ();
 sg13g2_fill_1 FILLER_66_193 ();
 sg13g2_decap_8 FILLER_66_197 ();
 sg13g2_decap_4 FILLER_66_204 ();
 sg13g2_decap_4 FILLER_66_216 ();
 sg13g2_fill_2 FILLER_66_220 ();
 sg13g2_decap_8 FILLER_66_225 ();
 sg13g2_fill_2 FILLER_66_232 ();
 sg13g2_decap_4 FILLER_66_243 ();
 sg13g2_fill_2 FILLER_66_247 ();
 sg13g2_decap_8 FILLER_66_259 ();
 sg13g2_decap_8 FILLER_66_266 ();
 sg13g2_decap_8 FILLER_66_273 ();
 sg13g2_decap_8 FILLER_66_280 ();
 sg13g2_decap_4 FILLER_66_287 ();
 sg13g2_fill_2 FILLER_66_291 ();
 sg13g2_fill_1 FILLER_66_296 ();
 sg13g2_fill_2 FILLER_66_338 ();
 sg13g2_decap_8 FILLER_66_366 ();
 sg13g2_decap_4 FILLER_66_373 ();
 sg13g2_fill_1 FILLER_66_377 ();
 sg13g2_decap_8 FILLER_66_402 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_8 FILLER_67_7 ();
 sg13g2_decap_8 FILLER_67_14 ();
 sg13g2_decap_8 FILLER_67_21 ();
 sg13g2_decap_8 FILLER_67_28 ();
 sg13g2_decap_8 FILLER_67_35 ();
 sg13g2_decap_8 FILLER_67_42 ();
 sg13g2_decap_8 FILLER_67_49 ();
 sg13g2_decap_8 FILLER_67_56 ();
 sg13g2_decap_8 FILLER_67_63 ();
 sg13g2_decap_8 FILLER_67_70 ();
 sg13g2_decap_8 FILLER_67_77 ();
 sg13g2_decap_4 FILLER_67_84 ();
 sg13g2_fill_2 FILLER_67_88 ();
 sg13g2_decap_4 FILLER_67_95 ();
 sg13g2_fill_1 FILLER_67_99 ();
 sg13g2_decap_4 FILLER_67_104 ();
 sg13g2_fill_2 FILLER_67_113 ();
 sg13g2_fill_1 FILLER_67_115 ();
 sg13g2_fill_2 FILLER_67_124 ();
 sg13g2_fill_1 FILLER_67_131 ();
 sg13g2_decap_4 FILLER_67_178 ();
 sg13g2_fill_1 FILLER_67_182 ();
 sg13g2_fill_1 FILLER_67_192 ();
 sg13g2_fill_2 FILLER_67_233 ();
 sg13g2_fill_2 FILLER_67_261 ();
 sg13g2_fill_1 FILLER_67_263 ();
 sg13g2_decap_4 FILLER_67_272 ();
 sg13g2_decap_8 FILLER_67_280 ();
 sg13g2_decap_8 FILLER_67_287 ();
 sg13g2_decap_4 FILLER_67_294 ();
 sg13g2_decap_4 FILLER_67_327 ();
 sg13g2_decap_8 FILLER_67_343 ();
 sg13g2_decap_8 FILLER_67_350 ();
 sg13g2_decap_8 FILLER_67_357 ();
 sg13g2_fill_2 FILLER_67_364 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_8 FILLER_68_7 ();
 sg13g2_decap_8 FILLER_68_14 ();
 sg13g2_decap_8 FILLER_68_21 ();
 sg13g2_decap_8 FILLER_68_28 ();
 sg13g2_decap_8 FILLER_68_35 ();
 sg13g2_decap_8 FILLER_68_42 ();
 sg13g2_decap_8 FILLER_68_49 ();
 sg13g2_decap_8 FILLER_68_56 ();
 sg13g2_decap_8 FILLER_68_63 ();
 sg13g2_decap_8 FILLER_68_70 ();
 sg13g2_decap_8 FILLER_68_77 ();
 sg13g2_fill_1 FILLER_68_84 ();
 sg13g2_fill_2 FILLER_68_93 ();
 sg13g2_fill_1 FILLER_68_100 ();
 sg13g2_fill_1 FILLER_68_127 ();
 sg13g2_fill_2 FILLER_68_267 ();
 sg13g2_fill_2 FILLER_68_278 ();
 sg13g2_fill_1 FILLER_68_280 ();
 sg13g2_decap_8 FILLER_68_289 ();
 sg13g2_decap_8 FILLER_68_296 ();
 sg13g2_decap_4 FILLER_68_303 ();
 sg13g2_fill_2 FILLER_68_307 ();
 sg13g2_decap_8 FILLER_68_316 ();
 sg13g2_decap_8 FILLER_68_323 ();
 sg13g2_fill_1 FILLER_68_369 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_8 FILLER_69_7 ();
 sg13g2_decap_8 FILLER_69_14 ();
 sg13g2_decap_8 FILLER_69_21 ();
 sg13g2_decap_8 FILLER_69_28 ();
 sg13g2_decap_8 FILLER_69_35 ();
 sg13g2_decap_8 FILLER_69_42 ();
 sg13g2_decap_8 FILLER_69_49 ();
 sg13g2_decap_8 FILLER_69_56 ();
 sg13g2_decap_8 FILLER_69_63 ();
 sg13g2_decap_8 FILLER_69_70 ();
 sg13g2_decap_8 FILLER_69_77 ();
 sg13g2_fill_2 FILLER_69_84 ();
 sg13g2_decap_8 FILLER_69_130 ();
 sg13g2_fill_2 FILLER_69_137 ();
 sg13g2_fill_2 FILLER_69_149 ();
 sg13g2_fill_1 FILLER_69_151 ();
 sg13g2_decap_4 FILLER_69_204 ();
 sg13g2_decap_8 FILLER_69_239 ();
 sg13g2_decap_4 FILLER_69_246 ();
 sg13g2_fill_2 FILLER_69_250 ();
 sg13g2_fill_1 FILLER_69_257 ();
 sg13g2_fill_1 FILLER_69_263 ();
 sg13g2_decap_8 FILLER_69_303 ();
 sg13g2_decap_8 FILLER_69_310 ();
 sg13g2_decap_8 FILLER_69_317 ();
 sg13g2_fill_2 FILLER_69_324 ();
 sg13g2_decap_8 FILLER_69_339 ();
 sg13g2_fill_2 FILLER_69_346 ();
 sg13g2_fill_1 FILLER_69_348 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_decap_8 FILLER_70_14 ();
 sg13g2_decap_8 FILLER_70_21 ();
 sg13g2_decap_8 FILLER_70_28 ();
 sg13g2_decap_8 FILLER_70_35 ();
 sg13g2_decap_8 FILLER_70_42 ();
 sg13g2_decap_8 FILLER_70_49 ();
 sg13g2_decap_8 FILLER_70_56 ();
 sg13g2_decap_8 FILLER_70_63 ();
 sg13g2_decap_8 FILLER_70_70 ();
 sg13g2_decap_4 FILLER_70_77 ();
 sg13g2_fill_2 FILLER_70_81 ();
 sg13g2_decap_4 FILLER_70_113 ();
 sg13g2_fill_2 FILLER_70_117 ();
 sg13g2_decap_8 FILLER_70_124 ();
 sg13g2_fill_2 FILLER_70_131 ();
 sg13g2_fill_1 FILLER_70_141 ();
 sg13g2_decap_8 FILLER_70_147 ();
 sg13g2_fill_2 FILLER_70_154 ();
 sg13g2_fill_2 FILLER_70_165 ();
 sg13g2_decap_8 FILLER_70_171 ();
 sg13g2_fill_2 FILLER_70_178 ();
 sg13g2_decap_8 FILLER_70_206 ();
 sg13g2_decap_4 FILLER_70_213 ();
 sg13g2_fill_2 FILLER_70_217 ();
 sg13g2_decap_8 FILLER_70_222 ();
 sg13g2_decap_8 FILLER_70_229 ();
 sg13g2_decap_8 FILLER_70_236 ();
 sg13g2_decap_4 FILLER_70_243 ();
 sg13g2_fill_2 FILLER_70_247 ();
 sg13g2_fill_2 FILLER_70_275 ();
 sg13g2_fill_1 FILLER_70_277 ();
 sg13g2_decap_8 FILLER_70_304 ();
 sg13g2_decap_4 FILLER_70_311 ();
 sg13g2_fill_1 FILLER_70_315 ();
 sg13g2_decap_4 FILLER_70_321 ();
 sg13g2_fill_1 FILLER_70_325 ();
 sg13g2_decap_8 FILLER_70_370 ();
 sg13g2_fill_2 FILLER_70_377 ();
 sg13g2_decap_4 FILLER_70_404 ();
 sg13g2_fill_1 FILLER_70_408 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_decap_8 FILLER_71_7 ();
 sg13g2_decap_8 FILLER_71_14 ();
 sg13g2_decap_8 FILLER_71_21 ();
 sg13g2_decap_8 FILLER_71_28 ();
 sg13g2_decap_8 FILLER_71_35 ();
 sg13g2_decap_8 FILLER_71_42 ();
 sg13g2_decap_8 FILLER_71_49 ();
 sg13g2_decap_8 FILLER_71_56 ();
 sg13g2_decap_8 FILLER_71_63 ();
 sg13g2_decap_8 FILLER_71_70 ();
 sg13g2_decap_8 FILLER_71_77 ();
 sg13g2_decap_8 FILLER_71_84 ();
 sg13g2_decap_8 FILLER_71_91 ();
 sg13g2_decap_8 FILLER_71_98 ();
 sg13g2_decap_8 FILLER_71_105 ();
 sg13g2_fill_2 FILLER_71_112 ();
 sg13g2_fill_1 FILLER_71_114 ();
 sg13g2_decap_4 FILLER_71_119 ();
 sg13g2_decap_4 FILLER_71_162 ();
 sg13g2_fill_2 FILLER_71_180 ();
 sg13g2_fill_1 FILLER_71_182 ();
 sg13g2_decap_4 FILLER_71_219 ();
 sg13g2_fill_2 FILLER_71_223 ();
 sg13g2_decap_4 FILLER_71_231 ();
 sg13g2_fill_2 FILLER_71_240 ();
 sg13g2_decap_4 FILLER_71_260 ();
 sg13g2_fill_2 FILLER_71_268 ();
 sg13g2_fill_1 FILLER_71_270 ();
 sg13g2_fill_1 FILLER_71_309 ();
 sg13g2_fill_2 FILLER_71_341 ();
 sg13g2_fill_2 FILLER_71_385 ();
 sg13g2_decap_8 FILLER_71_395 ();
 sg13g2_decap_8 FILLER_71_402 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_decap_8 FILLER_72_14 ();
 sg13g2_decap_8 FILLER_72_21 ();
 sg13g2_decap_8 FILLER_72_28 ();
 sg13g2_decap_8 FILLER_72_35 ();
 sg13g2_decap_8 FILLER_72_42 ();
 sg13g2_decap_8 FILLER_72_49 ();
 sg13g2_decap_8 FILLER_72_56 ();
 sg13g2_decap_8 FILLER_72_63 ();
 sg13g2_decap_8 FILLER_72_70 ();
 sg13g2_decap_8 FILLER_72_77 ();
 sg13g2_decap_8 FILLER_72_84 ();
 sg13g2_decap_4 FILLER_72_91 ();
 sg13g2_fill_1 FILLER_72_132 ();
 sg13g2_fill_1 FILLER_72_165 ();
 sg13g2_decap_4 FILLER_72_192 ();
 sg13g2_fill_2 FILLER_72_222 ();
 sg13g2_fill_1 FILLER_72_224 ();
 sg13g2_decap_4 FILLER_72_266 ();
 sg13g2_decap_8 FILLER_72_275 ();
 sg13g2_fill_1 FILLER_72_352 ();
 sg13g2_decap_4 FILLER_72_405 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_decap_8 FILLER_73_14 ();
 sg13g2_decap_8 FILLER_73_21 ();
 sg13g2_decap_8 FILLER_73_28 ();
 sg13g2_decap_8 FILLER_73_35 ();
 sg13g2_decap_8 FILLER_73_42 ();
 sg13g2_decap_8 FILLER_73_49 ();
 sg13g2_decap_8 FILLER_73_56 ();
 sg13g2_decap_8 FILLER_73_63 ();
 sg13g2_decap_8 FILLER_73_70 ();
 sg13g2_decap_8 FILLER_73_77 ();
 sg13g2_decap_8 FILLER_73_84 ();
 sg13g2_decap_8 FILLER_73_91 ();
 sg13g2_fill_1 FILLER_73_135 ();
 sg13g2_fill_1 FILLER_73_141 ();
 sg13g2_fill_1 FILLER_73_151 ();
 sg13g2_fill_1 FILLER_73_163 ();
 sg13g2_fill_2 FILLER_73_176 ();
 sg13g2_fill_1 FILLER_73_178 ();
 sg13g2_fill_1 FILLER_73_184 ();
 sg13g2_fill_1 FILLER_73_190 ();
 sg13g2_decap_8 FILLER_73_196 ();
 sg13g2_decap_4 FILLER_73_203 ();
 sg13g2_fill_1 FILLER_73_207 ();
 sg13g2_fill_1 FILLER_73_237 ();
 sg13g2_decap_8 FILLER_73_272 ();
 sg13g2_decap_8 FILLER_73_279 ();
 sg13g2_fill_2 FILLER_73_306 ();
 sg13g2_fill_1 FILLER_73_308 ();
 sg13g2_fill_2 FILLER_73_313 ();
 sg13g2_fill_1 FILLER_73_315 ();
 sg13g2_decap_8 FILLER_73_335 ();
 sg13g2_decap_4 FILLER_73_345 ();
 sg13g2_fill_2 FILLER_73_349 ();
 sg13g2_decap_8 FILLER_73_355 ();
 sg13g2_decap_8 FILLER_73_362 ();
 sg13g2_decap_8 FILLER_73_372 ();
 sg13g2_decap_8 FILLER_73_379 ();
 sg13g2_decap_8 FILLER_73_386 ();
 sg13g2_decap_8 FILLER_73_393 ();
 sg13g2_decap_8 FILLER_73_400 ();
 sg13g2_fill_2 FILLER_73_407 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_decap_8 FILLER_74_14 ();
 sg13g2_decap_8 FILLER_74_21 ();
 sg13g2_decap_8 FILLER_74_28 ();
 sg13g2_decap_8 FILLER_74_35 ();
 sg13g2_decap_8 FILLER_74_42 ();
 sg13g2_decap_8 FILLER_74_49 ();
 sg13g2_decap_8 FILLER_74_56 ();
 sg13g2_decap_8 FILLER_74_63 ();
 sg13g2_decap_8 FILLER_74_70 ();
 sg13g2_decap_8 FILLER_74_77 ();
 sg13g2_decap_8 FILLER_74_84 ();
 sg13g2_decap_8 FILLER_74_91 ();
 sg13g2_decap_4 FILLER_74_98 ();
 sg13g2_decap_8 FILLER_74_122 ();
 sg13g2_decap_4 FILLER_74_129 ();
 sg13g2_fill_2 FILLER_74_133 ();
 sg13g2_decap_4 FILLER_74_187 ();
 sg13g2_fill_1 FILLER_74_191 ();
 sg13g2_fill_1 FILLER_74_200 ();
 sg13g2_fill_2 FILLER_74_232 ();
 sg13g2_fill_2 FILLER_74_298 ();
 sg13g2_fill_2 FILLER_74_319 ();
 sg13g2_fill_2 FILLER_74_330 ();
 sg13g2_fill_1 FILLER_74_332 ();
 sg13g2_fill_1 FILLER_74_374 ();
 sg13g2_decap_8 FILLER_74_385 ();
 sg13g2_decap_8 FILLER_74_392 ();
 sg13g2_decap_8 FILLER_74_399 ();
 sg13g2_fill_2 FILLER_74_406 ();
 sg13g2_fill_1 FILLER_74_408 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_14 ();
 sg13g2_decap_8 FILLER_75_21 ();
 sg13g2_decap_8 FILLER_75_28 ();
 sg13g2_decap_8 FILLER_75_35 ();
 sg13g2_decap_8 FILLER_75_42 ();
 sg13g2_decap_8 FILLER_75_49 ();
 sg13g2_decap_8 FILLER_75_56 ();
 sg13g2_decap_8 FILLER_75_63 ();
 sg13g2_decap_8 FILLER_75_70 ();
 sg13g2_decap_8 FILLER_75_77 ();
 sg13g2_decap_8 FILLER_75_84 ();
 sg13g2_decap_8 FILLER_75_91 ();
 sg13g2_decap_8 FILLER_75_98 ();
 sg13g2_decap_4 FILLER_75_105 ();
 sg13g2_decap_8 FILLER_75_113 ();
 sg13g2_decap_4 FILLER_75_120 ();
 sg13g2_fill_1 FILLER_75_124 ();
 sg13g2_decap_8 FILLER_75_134 ();
 sg13g2_fill_1 FILLER_75_141 ();
 sg13g2_decap_8 FILLER_75_146 ();
 sg13g2_fill_1 FILLER_75_153 ();
 sg13g2_decap_8 FILLER_75_160 ();
 sg13g2_fill_1 FILLER_75_167 ();
 sg13g2_fill_1 FILLER_75_172 ();
 sg13g2_fill_1 FILLER_75_202 ();
 sg13g2_fill_2 FILLER_75_237 ();
 sg13g2_fill_1 FILLER_75_263 ();
 sg13g2_fill_2 FILLER_75_305 ();
 sg13g2_fill_1 FILLER_75_333 ();
 sg13g2_fill_1 FILLER_75_365 ();
 sg13g2_fill_1 FILLER_75_372 ();
 sg13g2_decap_8 FILLER_75_399 ();
 sg13g2_fill_2 FILLER_75_406 ();
 sg13g2_fill_1 FILLER_75_408 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_8 FILLER_76_21 ();
 sg13g2_decap_8 FILLER_76_28 ();
 sg13g2_decap_8 FILLER_76_35 ();
 sg13g2_decap_8 FILLER_76_42 ();
 sg13g2_decap_8 FILLER_76_49 ();
 sg13g2_decap_8 FILLER_76_56 ();
 sg13g2_decap_8 FILLER_76_63 ();
 sg13g2_decap_8 FILLER_76_70 ();
 sg13g2_decap_8 FILLER_76_77 ();
 sg13g2_decap_8 FILLER_76_84 ();
 sg13g2_decap_4 FILLER_76_91 ();
 sg13g2_fill_2 FILLER_76_95 ();
 sg13g2_decap_8 FILLER_76_158 ();
 sg13g2_decap_4 FILLER_76_165 ();
 sg13g2_fill_2 FILLER_76_169 ();
 sg13g2_decap_8 FILLER_76_202 ();
 sg13g2_decap_8 FILLER_76_209 ();
 sg13g2_fill_2 FILLER_76_216 ();
 sg13g2_fill_1 FILLER_76_218 ();
 sg13g2_decap_4 FILLER_76_222 ();
 sg13g2_decap_8 FILLER_76_232 ();
 sg13g2_decap_8 FILLER_76_239 ();
 sg13g2_decap_8 FILLER_76_259 ();
 sg13g2_decap_8 FILLER_76_266 ();
 sg13g2_fill_2 FILLER_76_283 ();
 sg13g2_fill_2 FILLER_76_353 ();
 sg13g2_decap_8 FILLER_76_402 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_decap_8 FILLER_77_28 ();
 sg13g2_decap_8 FILLER_77_35 ();
 sg13g2_decap_8 FILLER_77_42 ();
 sg13g2_decap_8 FILLER_77_49 ();
 sg13g2_decap_8 FILLER_77_56 ();
 sg13g2_decap_8 FILLER_77_63 ();
 sg13g2_decap_8 FILLER_77_70 ();
 sg13g2_decap_8 FILLER_77_77 ();
 sg13g2_decap_8 FILLER_77_84 ();
 sg13g2_fill_2 FILLER_77_91 ();
 sg13g2_decap_8 FILLER_77_163 ();
 sg13g2_decap_8 FILLER_77_170 ();
 sg13g2_decap_4 FILLER_77_177 ();
 sg13g2_fill_1 FILLER_77_181 ();
 sg13g2_decap_8 FILLER_77_195 ();
 sg13g2_decap_8 FILLER_77_202 ();
 sg13g2_decap_8 FILLER_77_209 ();
 sg13g2_decap_8 FILLER_77_216 ();
 sg13g2_decap_8 FILLER_77_223 ();
 sg13g2_decap_8 FILLER_77_230 ();
 sg13g2_decap_8 FILLER_77_263 ();
 sg13g2_fill_2 FILLER_77_369 ();
 sg13g2_decap_8 FILLER_77_394 ();
 sg13g2_decap_8 FILLER_77_401 ();
 sg13g2_fill_1 FILLER_77_408 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_decap_8 FILLER_78_28 ();
 sg13g2_decap_8 FILLER_78_35 ();
 sg13g2_decap_8 FILLER_78_42 ();
 sg13g2_decap_8 FILLER_78_49 ();
 sg13g2_decap_8 FILLER_78_56 ();
 sg13g2_decap_8 FILLER_78_63 ();
 sg13g2_decap_8 FILLER_78_70 ();
 sg13g2_decap_8 FILLER_78_77 ();
 sg13g2_decap_8 FILLER_78_84 ();
 sg13g2_decap_8 FILLER_78_91 ();
 sg13g2_decap_4 FILLER_78_98 ();
 sg13g2_fill_1 FILLER_78_102 ();
 sg13g2_fill_2 FILLER_78_134 ();
 sg13g2_fill_1 FILLER_78_136 ();
 sg13g2_fill_2 FILLER_78_142 ();
 sg13g2_decap_8 FILLER_78_170 ();
 sg13g2_decap_8 FILLER_78_177 ();
 sg13g2_decap_8 FILLER_78_184 ();
 sg13g2_decap_8 FILLER_78_191 ();
 sg13g2_decap_8 FILLER_78_198 ();
 sg13g2_decap_8 FILLER_78_205 ();
 sg13g2_decap_8 FILLER_78_212 ();
 sg13g2_decap_8 FILLER_78_219 ();
 sg13g2_decap_8 FILLER_78_226 ();
 sg13g2_fill_2 FILLER_78_233 ();
 sg13g2_fill_1 FILLER_78_261 ();
 sg13g2_fill_1 FILLER_78_332 ();
 sg13g2_decap_8 FILLER_78_387 ();
 sg13g2_decap_8 FILLER_78_394 ();
 sg13g2_decap_8 FILLER_78_401 ();
 sg13g2_fill_1 FILLER_78_408 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_decap_8 FILLER_79_35 ();
 sg13g2_decap_8 FILLER_79_42 ();
 sg13g2_decap_8 FILLER_79_49 ();
 sg13g2_decap_8 FILLER_79_56 ();
 sg13g2_decap_8 FILLER_79_63 ();
 sg13g2_decap_8 FILLER_79_70 ();
 sg13g2_decap_8 FILLER_79_77 ();
 sg13g2_decap_8 FILLER_79_84 ();
 sg13g2_decap_8 FILLER_79_91 ();
 sg13g2_decap_8 FILLER_79_98 ();
 sg13g2_decap_4 FILLER_79_105 ();
 sg13g2_fill_1 FILLER_79_109 ();
 sg13g2_decap_4 FILLER_79_114 ();
 sg13g2_fill_1 FILLER_79_118 ();
 sg13g2_decap_8 FILLER_79_155 ();
 sg13g2_decap_8 FILLER_79_162 ();
 sg13g2_decap_8 FILLER_79_169 ();
 sg13g2_decap_8 FILLER_79_176 ();
 sg13g2_decap_8 FILLER_79_183 ();
 sg13g2_decap_8 FILLER_79_190 ();
 sg13g2_decap_8 FILLER_79_197 ();
 sg13g2_decap_8 FILLER_79_204 ();
 sg13g2_decap_8 FILLER_79_211 ();
 sg13g2_decap_8 FILLER_79_218 ();
 sg13g2_decap_8 FILLER_79_225 ();
 sg13g2_decap_8 FILLER_79_232 ();
 sg13g2_fill_2 FILLER_79_239 ();
 sg13g2_fill_1 FILLER_79_241 ();
 sg13g2_decap_4 FILLER_79_263 ();
 sg13g2_fill_1 FILLER_79_267 ();
 sg13g2_decap_4 FILLER_79_272 ();
 sg13g2_decap_8 FILLER_79_288 ();
 sg13g2_decap_8 FILLER_79_295 ();
 sg13g2_decap_8 FILLER_79_302 ();
 sg13g2_decap_8 FILLER_79_309 ();
 sg13g2_fill_2 FILLER_79_316 ();
 sg13g2_decap_8 FILLER_79_327 ();
 sg13g2_decap_4 FILLER_79_334 ();
 sg13g2_fill_2 FILLER_79_346 ();
 sg13g2_fill_1 FILLER_79_353 ();
 sg13g2_fill_2 FILLER_79_363 ();
 sg13g2_fill_1 FILLER_79_365 ();
 sg13g2_decap_8 FILLER_79_392 ();
 sg13g2_decap_8 FILLER_79_399 ();
 sg13g2_fill_2 FILLER_79_406 ();
 sg13g2_fill_1 FILLER_79_408 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_42 ();
 sg13g2_decap_8 FILLER_80_49 ();
 sg13g2_decap_4 FILLER_80_60 ();
 sg13g2_decap_4 FILLER_80_68 ();
 sg13g2_decap_4 FILLER_80_76 ();
 sg13g2_decap_4 FILLER_80_84 ();
 sg13g2_decap_4 FILLER_80_92 ();
 sg13g2_decap_4 FILLER_80_100 ();
 sg13g2_decap_4 FILLER_80_108 ();
 sg13g2_decap_4 FILLER_80_116 ();
 sg13g2_decap_4 FILLER_80_124 ();
 sg13g2_decap_4 FILLER_80_132 ();
 sg13g2_decap_4 FILLER_80_140 ();
 sg13g2_decap_4 FILLER_80_148 ();
 sg13g2_decap_4 FILLER_80_156 ();
 sg13g2_decap_4 FILLER_80_164 ();
 sg13g2_decap_4 FILLER_80_172 ();
 sg13g2_decap_4 FILLER_80_180 ();
 sg13g2_decap_4 FILLER_80_188 ();
 sg13g2_decap_4 FILLER_80_196 ();
 sg13g2_decap_4 FILLER_80_204 ();
 sg13g2_decap_8 FILLER_80_212 ();
 sg13g2_decap_8 FILLER_80_219 ();
 sg13g2_decap_8 FILLER_80_226 ();
 sg13g2_decap_8 FILLER_80_233 ();
 sg13g2_decap_8 FILLER_80_240 ();
 sg13g2_decap_4 FILLER_80_247 ();
 sg13g2_decap_8 FILLER_80_255 ();
 sg13g2_decap_8 FILLER_80_262 ();
 sg13g2_decap_8 FILLER_80_269 ();
 sg13g2_decap_8 FILLER_80_276 ();
 sg13g2_decap_8 FILLER_80_283 ();
 sg13g2_decap_8 FILLER_80_290 ();
 sg13g2_decap_8 FILLER_80_297 ();
 sg13g2_decap_8 FILLER_80_304 ();
 sg13g2_decap_8 FILLER_80_319 ();
 sg13g2_decap_8 FILLER_80_326 ();
 sg13g2_decap_8 FILLER_80_333 ();
 sg13g2_decap_8 FILLER_80_340 ();
 sg13g2_decap_8 FILLER_80_347 ();
 sg13g2_decap_8 FILLER_80_354 ();
 sg13g2_decap_8 FILLER_80_361 ();
 sg13g2_decap_8 FILLER_80_372 ();
 sg13g2_decap_8 FILLER_80_379 ();
 sg13g2_decap_8 FILLER_80_386 ();
 sg13g2_decap_8 FILLER_80_393 ();
 sg13g2_decap_8 FILLER_80_400 ();
 sg13g2_fill_2 FILLER_80_407 ();
 assign uio_oe[0] = net2;
 assign uio_oe[1] = net3;
 assign uio_oe[2] = net4;
 assign uio_oe[3] = net5;
 assign uio_oe[4] = net6;
 assign uio_oe[5] = net7;
 assign uio_oe[6] = net8;
 assign uio_oe[7] = net9;
 assign uio_out[0] = net10;
 assign uio_out[1] = net11;
 assign uio_out[2] = net12;
 assign uio_out[3] = net13;
 assign uio_out[4] = net14;
 assign uio_out[5] = net15;
 assign uio_out[6] = net16;
 assign uio_out[7] = net17;
 assign uo_out[4] = net18;
 assign uo_out[5] = net19;
 assign uo_out[6] = net20;
 assign uo_out[7] = net21;
endmodule

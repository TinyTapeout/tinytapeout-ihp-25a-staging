module tt_um_led_cipher (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire \bitserial_cipher.bcount[0] ;
 wire \bitserial_cipher.bcount[1] ;
 wire \bitserial_cipher.bcount[2] ;
 wire \bitserial_cipher.bcount[3] ;
 wire \bitserial_cipher.ctlstate[0] ;
 wire \bitserial_cipher.ctlstate[1] ;
 wire \bitserial_cipher.ctlstate[2] ;
 wire \bitserial_cipher.ctlstate[3] ;
 wire \bitserial_cipher.ctlstate_next[0] ;
 wire \bitserial_cipher.ctlstate_next[1] ;
 wire \bitserial_cipher.ctlstate_next[2] ;
 wire \bitserial_cipher.ctlstate_next[3] ;
 wire \bitserial_cipher.dataq ;
 wire \bitserial_cipher.done ;
 wire \bitserial_cipher.key[0] ;
 wire \bitserial_cipher.key[100] ;
 wire \bitserial_cipher.key[101] ;
 wire \bitserial_cipher.key[102] ;
 wire \bitserial_cipher.key[103] ;
 wire \bitserial_cipher.key[104] ;
 wire \bitserial_cipher.key[105] ;
 wire \bitserial_cipher.key[106] ;
 wire \bitserial_cipher.key[107] ;
 wire \bitserial_cipher.key[108] ;
 wire \bitserial_cipher.key[109] ;
 wire \bitserial_cipher.key[10] ;
 wire \bitserial_cipher.key[110] ;
 wire \bitserial_cipher.key[111] ;
 wire \bitserial_cipher.key[112] ;
 wire \bitserial_cipher.key[113] ;
 wire \bitserial_cipher.key[114] ;
 wire \bitserial_cipher.key[115] ;
 wire \bitserial_cipher.key[116] ;
 wire \bitserial_cipher.key[117] ;
 wire \bitserial_cipher.key[118] ;
 wire \bitserial_cipher.key[119] ;
 wire \bitserial_cipher.key[11] ;
 wire \bitserial_cipher.key[120] ;
 wire \bitserial_cipher.key[121] ;
 wire \bitserial_cipher.key[122] ;
 wire \bitserial_cipher.key[123] ;
 wire \bitserial_cipher.key[124] ;
 wire \bitserial_cipher.key[125] ;
 wire \bitserial_cipher.key[126] ;
 wire \bitserial_cipher.key[127] ;
 wire \bitserial_cipher.key[12] ;
 wire \bitserial_cipher.key[13] ;
 wire \bitserial_cipher.key[14] ;
 wire \bitserial_cipher.key[15] ;
 wire \bitserial_cipher.key[16] ;
 wire \bitserial_cipher.key[17] ;
 wire \bitserial_cipher.key[18] ;
 wire \bitserial_cipher.key[19] ;
 wire \bitserial_cipher.key[1] ;
 wire \bitserial_cipher.key[20] ;
 wire \bitserial_cipher.key[21] ;
 wire \bitserial_cipher.key[22] ;
 wire \bitserial_cipher.key[23] ;
 wire \bitserial_cipher.key[24] ;
 wire \bitserial_cipher.key[25] ;
 wire \bitserial_cipher.key[26] ;
 wire \bitserial_cipher.key[27] ;
 wire \bitserial_cipher.key[28] ;
 wire \bitserial_cipher.key[29] ;
 wire \bitserial_cipher.key[2] ;
 wire \bitserial_cipher.key[30] ;
 wire \bitserial_cipher.key[31] ;
 wire \bitserial_cipher.key[32] ;
 wire \bitserial_cipher.key[33] ;
 wire \bitserial_cipher.key[34] ;
 wire \bitserial_cipher.key[35] ;
 wire \bitserial_cipher.key[36] ;
 wire \bitserial_cipher.key[37] ;
 wire \bitserial_cipher.key[38] ;
 wire \bitserial_cipher.key[39] ;
 wire \bitserial_cipher.key[3] ;
 wire \bitserial_cipher.key[40] ;
 wire \bitserial_cipher.key[41] ;
 wire \bitserial_cipher.key[42] ;
 wire \bitserial_cipher.key[43] ;
 wire \bitserial_cipher.key[44] ;
 wire \bitserial_cipher.key[45] ;
 wire \bitserial_cipher.key[46] ;
 wire \bitserial_cipher.key[47] ;
 wire \bitserial_cipher.key[48] ;
 wire \bitserial_cipher.key[49] ;
 wire \bitserial_cipher.key[4] ;
 wire \bitserial_cipher.key[50] ;
 wire \bitserial_cipher.key[51] ;
 wire \bitserial_cipher.key[52] ;
 wire \bitserial_cipher.key[53] ;
 wire \bitserial_cipher.key[54] ;
 wire \bitserial_cipher.key[55] ;
 wire \bitserial_cipher.key[56] ;
 wire \bitserial_cipher.key[57] ;
 wire \bitserial_cipher.key[58] ;
 wire \bitserial_cipher.key[59] ;
 wire \bitserial_cipher.key[5] ;
 wire \bitserial_cipher.key[60] ;
 wire \bitserial_cipher.key[61] ;
 wire \bitserial_cipher.key[62] ;
 wire \bitserial_cipher.key[63] ;
 wire \bitserial_cipher.key[64] ;
 wire \bitserial_cipher.key[65] ;
 wire \bitserial_cipher.key[66] ;
 wire \bitserial_cipher.key[67] ;
 wire \bitserial_cipher.key[68] ;
 wire \bitserial_cipher.key[69] ;
 wire \bitserial_cipher.key[6] ;
 wire \bitserial_cipher.key[70] ;
 wire \bitserial_cipher.key[71] ;
 wire \bitserial_cipher.key[72] ;
 wire \bitserial_cipher.key[73] ;
 wire \bitserial_cipher.key[74] ;
 wire \bitserial_cipher.key[75] ;
 wire \bitserial_cipher.key[76] ;
 wire \bitserial_cipher.key[77] ;
 wire \bitserial_cipher.key[78] ;
 wire \bitserial_cipher.key[79] ;
 wire \bitserial_cipher.key[7] ;
 wire \bitserial_cipher.key[80] ;
 wire \bitserial_cipher.key[81] ;
 wire \bitserial_cipher.key[82] ;
 wire \bitserial_cipher.key[83] ;
 wire \bitserial_cipher.key[84] ;
 wire \bitserial_cipher.key[85] ;
 wire \bitserial_cipher.key[86] ;
 wire \bitserial_cipher.key[87] ;
 wire \bitserial_cipher.key[88] ;
 wire \bitserial_cipher.key[89] ;
 wire \bitserial_cipher.key[8] ;
 wire \bitserial_cipher.key[90] ;
 wire \bitserial_cipher.key[91] ;
 wire \bitserial_cipher.key[92] ;
 wire \bitserial_cipher.key[93] ;
 wire \bitserial_cipher.key[94] ;
 wire \bitserial_cipher.key[95] ;
 wire \bitserial_cipher.key[96] ;
 wire \bitserial_cipher.key[97] ;
 wire \bitserial_cipher.key[98] ;
 wire \bitserial_cipher.key[99] ;
 wire \bitserial_cipher.key[9] ;
 wire \bitserial_cipher.rc[0] ;
 wire \bitserial_cipher.rc[1] ;
 wire \bitserial_cipher.rc[2] ;
 wire \bitserial_cipher.rc[3] ;
 wire \bitserial_cipher.rc[4] ;
 wire \bitserial_cipher.rc[5] ;
 wire \bitserial_cipher.rcount[0] ;
 wire \bitserial_cipher.rcount[1] ;
 wire \bitserial_cipher.rcount[2] ;
 wire \bitserial_cipher.rcount[3] ;
 wire \bitserial_cipher.scount[0] ;
 wire \bitserial_cipher.scount[1] ;
 wire \bitserial_cipher.scount[2] ;
 wire \bitserial_cipher.scount[3] ;
 wire \bitserial_cipher.state[0] ;
 wire \bitserial_cipher.state[10] ;
 wire \bitserial_cipher.state[11] ;
 wire \bitserial_cipher.state[12] ;
 wire \bitserial_cipher.state[13] ;
 wire \bitserial_cipher.state[14] ;
 wire \bitserial_cipher.state[15] ;
 wire \bitserial_cipher.state[16] ;
 wire \bitserial_cipher.state[17] ;
 wire \bitserial_cipher.state[18] ;
 wire \bitserial_cipher.state[19] ;
 wire \bitserial_cipher.state[1] ;
 wire \bitserial_cipher.state[20] ;
 wire \bitserial_cipher.state[21] ;
 wire \bitserial_cipher.state[22] ;
 wire \bitserial_cipher.state[23] ;
 wire \bitserial_cipher.state[24] ;
 wire \bitserial_cipher.state[25] ;
 wire \bitserial_cipher.state[26] ;
 wire \bitserial_cipher.state[27] ;
 wire \bitserial_cipher.state[28] ;
 wire \bitserial_cipher.state[29] ;
 wire \bitserial_cipher.state[2] ;
 wire \bitserial_cipher.state[30] ;
 wire \bitserial_cipher.state[31] ;
 wire \bitserial_cipher.state[32] ;
 wire \bitserial_cipher.state[33] ;
 wire \bitserial_cipher.state[34] ;
 wire \bitserial_cipher.state[35] ;
 wire \bitserial_cipher.state[36] ;
 wire \bitserial_cipher.state[37] ;
 wire \bitserial_cipher.state[38] ;
 wire \bitserial_cipher.state[39] ;
 wire \bitserial_cipher.state[3] ;
 wire \bitserial_cipher.state[40] ;
 wire \bitserial_cipher.state[41] ;
 wire \bitserial_cipher.state[42] ;
 wire \bitserial_cipher.state[43] ;
 wire \bitserial_cipher.state[44] ;
 wire \bitserial_cipher.state[45] ;
 wire \bitserial_cipher.state[46] ;
 wire \bitserial_cipher.state[47] ;
 wire \bitserial_cipher.state[48] ;
 wire \bitserial_cipher.state[49] ;
 wire \bitserial_cipher.state[4] ;
 wire \bitserial_cipher.state[50] ;
 wire \bitserial_cipher.state[51] ;
 wire \bitserial_cipher.state[52] ;
 wire \bitserial_cipher.state[53] ;
 wire \bitserial_cipher.state[54] ;
 wire \bitserial_cipher.state[55] ;
 wire \bitserial_cipher.state[56] ;
 wire \bitserial_cipher.state[57] ;
 wire \bitserial_cipher.state[58] ;
 wire \bitserial_cipher.state[59] ;
 wire \bitserial_cipher.state[5] ;
 wire \bitserial_cipher.state[60] ;
 wire \bitserial_cipher.state[61] ;
 wire \bitserial_cipher.state[62] ;
 wire \bitserial_cipher.state[6] ;
 wire \bitserial_cipher.state[7] ;
 wire \bitserial_cipher.state[8] ;
 wire \bitserial_cipher.state[9] ;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire clknet_leaf_0_clk;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;

 sg13g2_inv_1 _1119_ (.Y(_0452_),
    .A(\bitserial_cipher.ctlstate[0] ));
 sg13g2_inv_1 _1120_ (.Y(_0453_),
    .A(\bitserial_cipher.ctlstate[2] ));
 sg13g2_inv_1 _1121_ (.Y(_0454_),
    .A(net4));
 sg13g2_inv_1 _1122_ (.Y(_0455_),
    .A(\bitserial_cipher.scount[1] ));
 sg13g2_inv_1 _1123_ (.Y(_0456_),
    .A(net327));
 sg13g2_inv_1 _1124_ (.Y(_0457_),
    .A(\bitserial_cipher.rc[4] ));
 sg13g2_inv_1 _1125_ (.Y(_0458_),
    .A(net87));
 sg13g2_inv_1 _1126_ (.Y(_0459_),
    .A(net89));
 sg13g2_inv_1 _1127_ (.Y(_0460_),
    .A(\bitserial_cipher.key[113] ));
 sg13g2_inv_1 _1128_ (.Y(_0461_),
    .A(net75));
 sg13g2_inv_1 _1129_ (.Y(_0462_),
    .A(net181));
 sg13g2_inv_1 _1130_ (.Y(_0463_),
    .A(net221));
 sg13g2_inv_1 _1131_ (.Y(_0464_),
    .A(net130));
 sg13g2_inv_1 _1132_ (.Y(_0465_),
    .A(net224));
 sg13g2_inv_1 _1133_ (.Y(_0466_),
    .A(net36));
 sg13g2_inv_1 _1134_ (.Y(_0467_),
    .A(net141));
 sg13g2_inv_1 _1135_ (.Y(_0468_),
    .A(\bitserial_cipher.state[33] ));
 sg13g2_inv_1 _1136_ (.Y(_0469_),
    .A(net105));
 sg13g2_inv_1 _1137_ (.Y(_0470_),
    .A(net71));
 sg13g2_inv_1 _1138_ (.Y(_0471_),
    .A(net63));
 sg13g2_inv_1 _1139_ (.Y(_0472_),
    .A(net91));
 sg13g2_inv_1 _1140_ (.Y(_0473_),
    .A(net57));
 sg13g2_inv_1 _1141_ (.Y(_0474_),
    .A(net170));
 sg13g2_inv_1 _1142_ (.Y(_0475_),
    .A(net111));
 sg13g2_inv_1 _1143_ (.Y(_0476_),
    .A(net55));
 sg13g2_inv_1 _1144_ (.Y(_0477_),
    .A(net101));
 sg13g2_inv_1 _1145_ (.Y(_0478_),
    .A(net85));
 sg13g2_inv_1 _1146_ (.Y(_0479_),
    .A(net118));
 sg13g2_inv_1 _1147_ (.Y(_0480_),
    .A(net69));
 sg13g2_inv_1 _1148_ (.Y(_0481_),
    .A(net107));
 sg13g2_inv_1 _1149_ (.Y(_0482_),
    .A(net147));
 sg13g2_inv_1 _1150_ (.Y(_0483_),
    .A(net126));
 sg13g2_inv_1 _1151_ (.Y(_0484_),
    .A(net128));
 sg13g2_inv_1 _1152_ (.Y(_0485_),
    .A(net67));
 sg13g2_inv_1 _1153_ (.Y(_0486_),
    .A(net121));
 sg13g2_inv_1 _1154_ (.Y(_0487_),
    .A(net172));
 sg13g2_inv_1 _1155_ (.Y(_0488_),
    .A(net93));
 sg13g2_inv_1 _1156_ (.Y(_0489_),
    .A(\bitserial_cipher.key[29] ));
 sg13g2_inv_1 _1157_ (.Y(_0490_),
    .A(net230));
 sg13g2_inv_1 _1158_ (.Y(_0491_),
    .A(net133));
 sg13g2_inv_1 _1159_ (.Y(_0492_),
    .A(net59));
 sg13g2_inv_1 _1160_ (.Y(_0493_),
    .A(net83));
 sg13g2_inv_1 _1161_ (.Y(_0494_),
    .A(net203));
 sg13g2_inv_1 _1162_ (.Y(_0495_),
    .A(net38));
 sg13g2_inv_1 _1163_ (.Y(_0496_),
    .A(net132));
 sg13g2_inv_1 _1164_ (.Y(_0497_),
    .A(net283));
 sg13g2_inv_1 _1165_ (.Y(_0498_),
    .A(net243));
 sg13g2_inv_1 _1166_ (.Y(_0499_),
    .A(\bitserial_cipher.state[49] ));
 sg13g2_inv_1 _1167_ (.Y(_0500_),
    .A(net326));
 sg13g2_inv_1 _1168_ (.Y(_0501_),
    .A(\bitserial_cipher.state[13] ));
 sg13g2_inv_1 _1169_ (.Y(_0502_),
    .A(net304));
 sg13g2_inv_1 _1170_ (.Y(_0503_),
    .A(net329));
 sg13g2_inv_1 _1171_ (.Y(_0504_),
    .A(net340));
 sg13g2_inv_1 _1172_ (.Y(_0505_),
    .A(net331));
 sg13g2_inv_1 _1173_ (.Y(_0506_),
    .A(net324));
 sg13g2_inv_1 _1174_ (.Y(_0507_),
    .A(net361));
 sg13g2_inv_1 _1175_ (.Y(_0508_),
    .A(net346));
 sg13g2_nor2_2 _1176_ (.A(\bitserial_cipher.ctlstate[3] ),
    .B(\bitserial_cipher.ctlstate[2] ),
    .Y(_0509_));
 sg13g2_nor2_2 _1177_ (.A(\bitserial_cipher.ctlstate[1] ),
    .B(\bitserial_cipher.ctlstate[0] ),
    .Y(_0510_));
 sg13g2_nand2_1 _1178_ (.Y(_0511_),
    .A(_0509_),
    .B(_0510_));
 sg13g2_inv_2 _1179_ (.Y(\bitserial_cipher.done ),
    .A(_0511_));
 sg13g2_and2_1 _1180_ (.A(\bitserial_cipher.bcount[0] ),
    .B(\bitserial_cipher.bcount[1] ),
    .X(_0512_));
 sg13g2_nand2_1 _1181_ (.Y(_0513_),
    .A(\bitserial_cipher.bcount[0] ),
    .B(\bitserial_cipher.bcount[1] ));
 sg13g2_nand3_1 _1182_ (.B(net362),
    .C(_0512_),
    .A(\bitserial_cipher.bcount[2] ),
    .Y(_0514_));
 sg13g2_nand2b_1 _1183_ (.Y(_0515_),
    .B(\bitserial_cipher.ctlstate[0] ),
    .A_N(\bitserial_cipher.ctlstate[1] ));
 sg13g2_nor3_1 _1184_ (.A(\bitserial_cipher.ctlstate[1] ),
    .B(net617),
    .C(\bitserial_cipher.ctlstate[2] ),
    .Y(_0516_));
 sg13g2_and2_1 _1185_ (.A(\bitserial_cipher.ctlstate[0] ),
    .B(_0516_),
    .X(_0517_));
 sg13g2_nor2b_1 _1186_ (.A(\bitserial_cipher.ctlstate[2] ),
    .B_N(\bitserial_cipher.ctlstate[1] ),
    .Y(_0518_));
 sg13g2_and2_1 _1187_ (.A(_0452_),
    .B(_0518_),
    .X(_0519_));
 sg13g2_nor2b_1 _1188_ (.A(_0514_),
    .B_N(_0519_),
    .Y(_0520_));
 sg13g2_a21oi_1 _1189_ (.A1(net363),
    .A2(_0517_),
    .Y(_0521_),
    .B1(_0520_));
 sg13g2_nor2_1 _1190_ (.A(net617),
    .B(_0453_),
    .Y(_0522_));
 sg13g2_nor2b_1 _1191_ (.A(\bitserial_cipher.ctlstate[2] ),
    .B_N(net617),
    .Y(_0523_));
 sg13g2_nand2_1 _1192_ (.Y(_0524_),
    .A(net617),
    .B(_0453_));
 sg13g2_and2_2 _1193_ (.A(_0510_),
    .B(_0523_),
    .X(_0525_));
 sg13g2_inv_1 _1194_ (.Y(_0526_),
    .A(net611));
 sg13g2_nor3_2 _1195_ (.A(net354),
    .B(net346),
    .C(_0513_),
    .Y(_0527_));
 sg13g2_nand2_1 _1196_ (.Y(_0528_),
    .A(net611),
    .B(_0527_));
 sg13g2_a22oi_1 _1197_ (.Y(_0529_),
    .B1(net615),
    .B2(_0452_),
    .A2(\bitserial_cipher.done ),
    .A1(net5));
 sg13g2_nand3_1 _1198_ (.B(_0528_),
    .C(_0529_),
    .A(net364),
    .Y(\bitserial_cipher.ctlstate_next[0] ));
 sg13g2_nand2_1 _1199_ (.Y(_0530_),
    .A(\bitserial_cipher.ctlstate[1] ),
    .B(\bitserial_cipher.ctlstate[0] ));
 sg13g2_nand3_1 _1200_ (.B(\bitserial_cipher.ctlstate[0] ),
    .C(_0523_),
    .A(\bitserial_cipher.ctlstate[1] ),
    .Y(_0531_));
 sg13g2_nor3_1 _1201_ (.A(_0455_),
    .B(_0456_),
    .C(net360),
    .Y(_0532_));
 sg13g2_a21oi_1 _1202_ (.A1(net30),
    .A2(_0532_),
    .Y(_0533_),
    .B1(_0531_));
 sg13g2_nor2_2 _1203_ (.A(_0515_),
    .B(_0524_),
    .Y(_0534_));
 sg13g2_nand2b_1 _1204_ (.Y(_0535_),
    .B(_0523_),
    .A_N(_0515_));
 sg13g2_nand2_1 _1205_ (.Y(_0536_),
    .A(net615),
    .B(_0530_));
 sg13g2_nand2b_1 _1206_ (.Y(_0537_),
    .B(_0517_),
    .A_N(_0514_));
 sg13g2_o21ai_1 _1207_ (.B1(_0537_),
    .Y(_0538_),
    .A1(_0510_),
    .A2(_0536_));
 sg13g2_or4_1 _1208_ (.A(_0519_),
    .B(_0533_),
    .C(_0534_),
    .D(_0538_),
    .X(\bitserial_cipher.ctlstate_next[1] ));
 sg13g2_nor3_1 _1209_ (.A(net617),
    .B(\bitserial_cipher.ctlstate[2] ),
    .C(_0530_),
    .Y(_0539_));
 sg13g2_nor2_1 _1210_ (.A(_0526_),
    .B(_0527_),
    .Y(_0540_));
 sg13g2_a21oi_1 _1211_ (.A1(net615),
    .A2(_0530_),
    .Y(_0541_),
    .B1(net608));
 sg13g2_o21ai_1 _1212_ (.B1(_0541_),
    .Y(\bitserial_cipher.ctlstate_next[2] ),
    .A1(_0526_),
    .A2(_0527_));
 sg13g2_nand3_1 _1213_ (.B(\bitserial_cipher.ctlstate[0] ),
    .C(net615),
    .A(\bitserial_cipher.ctlstate[1] ),
    .Y(_0542_));
 sg13g2_nand2_1 _1214_ (.Y(_0543_),
    .A(net343),
    .B(net239));
 sg13g2_nor4_2 _1215_ (.A(net61),
    .B(net318),
    .C(_0535_),
    .Y(_0544_),
    .D(_0543_));
 sg13g2_nand2_1 _1216_ (.Y(_0545_),
    .A(net617),
    .B(_0519_));
 sg13g2_nand3_1 _1217_ (.B(_0542_),
    .C(_0545_),
    .A(_0528_),
    .Y(_0546_));
 sg13g2_or2_1 _1218_ (.X(\bitserial_cipher.ctlstate_next[3] ),
    .B(_0546_),
    .A(_0544_));
 sg13g2_mux2_1 _1219_ (.A0(_0516_),
    .A1(_0518_),
    .S(_0452_),
    .X(_0547_));
 sg13g2_nor2_1 _1220_ (.A(net611),
    .B(net601),
    .Y(_0548_));
 sg13g2_or2_1 _1221_ (.X(_0549_),
    .B(net601),
    .A(net611));
 sg13g2_nand3b_1 _1222_ (.B(net2),
    .C(\bitserial_cipher.done ),
    .Y(_0550_),
    .A_N(net3));
 sg13g2_or2_1 _1223_ (.X(_0551_),
    .B(net2),
    .A(net3));
 sg13g2_o21ai_1 _1224_ (.B1(_0510_),
    .Y(_0552_),
    .A1(_0454_),
    .A2(_0551_));
 sg13g2_nand2_1 _1225_ (.Y(_0553_),
    .A(_0509_),
    .B(_0552_));
 sg13g2_a22oi_1 _1226_ (.Y(_0554_),
    .B1(_0552_),
    .B2(_0509_),
    .A2(_0519_),
    .A1(net617));
 sg13g2_nand2_2 _1227_ (.Y(_0555_),
    .A(_0545_),
    .B(_0553_));
 sg13g2_a21oi_1 _1228_ (.A1(\bitserial_cipher.ctlstate[0] ),
    .A2(_0453_),
    .Y(_0556_),
    .B1(net617));
 sg13g2_nand2_2 _1229_ (.Y(_0557_),
    .A(_0550_),
    .B(_0556_));
 sg13g2_a22oi_1 _1230_ (.Y(_0558_),
    .B1(\bitserial_cipher.done ),
    .B2(_0551_),
    .A2(_0509_),
    .A1(\bitserial_cipher.ctlstate[1] ));
 sg13g2_nor2b_1 _1231_ (.A(_0557_),
    .B_N(_0558_),
    .Y(_0559_));
 sg13g2_nand3_1 _1232_ (.B(_0556_),
    .C(_0558_),
    .A(_0550_),
    .Y(_0560_));
 sg13g2_nand2_1 _1233_ (.Y(_0561_),
    .A(_0555_),
    .B(_0559_));
 sg13g2_o21ai_1 _1234_ (.B1(_0550_),
    .Y(_0562_),
    .A1(_0554_),
    .A2(_0560_));
 sg13g2_nor2_1 _1235_ (.A(net593),
    .B(net581),
    .Y(_0563_));
 sg13g2_nor2_2 _1236_ (.A(net613),
    .B(net595),
    .Y(_0564_));
 sg13g2_or2_1 _1237_ (.X(_0565_),
    .B(net604),
    .A(net610));
 sg13g2_nor2_2 _1238_ (.A(net608),
    .B(net596),
    .Y(_0566_));
 sg13g2_nand2b_1 _1239_ (.Y(_0567_),
    .B(net597),
    .A_N(net604));
 sg13g2_nor2_1 _1240_ (.A(net612),
    .B(net585),
    .Y(_0568_));
 sg13g2_nor2b_2 _1241_ (.A(net580),
    .B_N(_0564_),
    .Y(_0569_));
 sg13g2_nand2_1 _1242_ (.Y(_0570_),
    .A(net553),
    .B(net583));
 sg13g2_a22oi_1 _1243_ (.Y(_0571_),
    .B1(net582),
    .B2(\bitserial_cipher.state[44] ),
    .A2(net614),
    .A1(\bitserial_cipher.state[29] ));
 sg13g2_o21ai_1 _1244_ (.B1(_0571_),
    .Y(_0572_),
    .A1(_0465_),
    .A2(net588));
 sg13g2_mux2_1 _1245_ (.A0(net337),
    .A1(_0572_),
    .S(net512),
    .X(_0001_));
 sg13g2_nor2_1 _1246_ (.A(net307),
    .B(net512),
    .Y(_0573_));
 sg13g2_and2_1 _1247_ (.A(\bitserial_cipher.state[30] ),
    .B(net612),
    .X(_0574_));
 sg13g2_a221oi_1 _1248_ (.B2(net337),
    .C1(_0574_),
    .B1(net582),
    .A1(net79),
    .Y(_0575_),
    .A2(net584));
 sg13g2_a21oi_1 _1249_ (.A1(net512),
    .A2(_0575_),
    .Y(_0002_),
    .B1(_0573_));
 sg13g2_and2_1 _1250_ (.A(\bitserial_cipher.state[31] ),
    .B(net612),
    .X(_0576_));
 sg13g2_a221oi_1 _1251_ (.B2(net307),
    .C1(_0576_),
    .B1(net582),
    .A1(net341),
    .Y(_0577_),
    .A2(net584));
 sg13g2_nor2_1 _1252_ (.A(net162),
    .B(net512),
    .Y(_0578_));
 sg13g2_a21oi_1 _1253_ (.A1(net512),
    .A2(_0577_),
    .Y(_0003_),
    .B1(_0578_));
 sg13g2_nand2_1 _1254_ (.Y(_0579_),
    .A(net162),
    .B(net597));
 sg13g2_a22oi_1 _1255_ (.Y(_0580_),
    .B1(net600),
    .B2(net366),
    .A2(net611),
    .A1(\bitserial_cipher.state[60] ));
 sg13g2_a21oi_1 _1256_ (.A1(_0579_),
    .A2(_0580_),
    .Y(_0581_),
    .B1(net553));
 sg13g2_a21o_1 _1257_ (.A2(net554),
    .A1(net109),
    .B1(_0581_),
    .X(_0004_));
 sg13g2_nand2_1 _1258_ (.Y(_0582_),
    .A(net109),
    .B(net597));
 sg13g2_a221oi_1 _1259_ (.B2(\bitserial_cipher.state[45] ),
    .C1(net553),
    .B1(net600),
    .A1(\bitserial_cipher.state[61] ),
    .Y(_0583_),
    .A2(net611));
 sg13g2_a22oi_1 _1260_ (.Y(_0005_),
    .B1(_0582_),
    .B2(_0583_),
    .A2(net553),
    .A1(_0499_));
 sg13g2_nand2_1 _1261_ (.Y(_0584_),
    .A(net228),
    .B(net597));
 sg13g2_a221oi_1 _1262_ (.B2(\bitserial_cipher.state[46] ),
    .C1(net553),
    .B1(net600),
    .A1(\bitserial_cipher.state[62] ),
    .Y(_0585_),
    .A2(net610));
 sg13g2_a22oi_1 _1263_ (.Y(_0006_),
    .B1(_0584_),
    .B2(_0585_),
    .A2(net553),
    .A1(_0500_));
 sg13g2_a22oi_1 _1264_ (.Y(_0586_),
    .B1(net600),
    .B2(net162),
    .A2(net610),
    .A1(\bitserial_cipher.dataq ));
 sg13g2_o21ai_1 _1265_ (.B1(_0586_),
    .Y(_0587_),
    .A1(_0500_),
    .A2(net593));
 sg13g2_mux2_1 _1266_ (.A0(_0587_),
    .A1(net95),
    .S(net553),
    .X(_0007_));
 sg13g2_xnor2_1 _1267_ (.Y(_0588_),
    .A(\bitserial_cipher.state[44] ),
    .B(\bitserial_cipher.state[31] ));
 sg13g2_xor2_1 _1268_ (.B(\bitserial_cipher.state[62] ),
    .A(\bitserial_cipher.state[15] ),
    .X(_0589_));
 sg13g2_xnor2_1 _1269_ (.Y(_0590_),
    .A(_0588_),
    .B(_0589_));
 sg13g2_a22oi_1 _1270_ (.Y(_0591_),
    .B1(net594),
    .B2(\bitserial_cipher.state[8] ),
    .A2(net606),
    .A1(\bitserial_cipher.state[0] ));
 sg13g2_inv_1 _1271_ (.Y(_0592_),
    .A(_0591_));
 sg13g2_a221oi_1 _1272_ (.B2(net613),
    .C1(_0592_),
    .B1(_0590_),
    .A1(net310),
    .Y(_0593_),
    .A2(net583));
 sg13g2_nor2_1 _1273_ (.A(net349),
    .B(_0570_),
    .Y(_0594_));
 sg13g2_a21oi_1 _1274_ (.A1(net513),
    .A2(_0593_),
    .Y(_0008_),
    .B1(_0594_));
 sg13g2_nor2_1 _1275_ (.A(net344),
    .B(net513),
    .Y(_0595_));
 sg13g2_xor2_1 _1276_ (.B(\bitserial_cipher.dataq ),
    .A(\bitserial_cipher.state[62] ),
    .X(_0596_));
 sg13g2_xor2_1 _1277_ (.B(\bitserial_cipher.state[15] ),
    .A(\bitserial_cipher.state[12] ),
    .X(_0597_));
 sg13g2_xnor2_1 _1278_ (.Y(_0598_),
    .A(_0596_),
    .B(_0597_));
 sg13g2_xnor2_1 _1279_ (.Y(_0599_),
    .A(\bitserial_cipher.state[31] ),
    .B(\bitserial_cipher.state[45] ));
 sg13g2_xnor2_1 _1280_ (.Y(_0600_),
    .A(\bitserial_cipher.state[28] ),
    .B(_0599_));
 sg13g2_xnor2_1 _1281_ (.Y(_0601_),
    .A(_0598_),
    .B(_0600_));
 sg13g2_a22oi_1 _1282_ (.Y(_0602_),
    .B1(net594),
    .B2(\bitserial_cipher.state[9] ),
    .A2(net605),
    .A1(\bitserial_cipher.state[1] ));
 sg13g2_inv_1 _1283_ (.Y(_0603_),
    .A(_0602_));
 sg13g2_a221oi_1 _1284_ (.B2(net613),
    .C1(_0603_),
    .B1(_0601_),
    .A1(net367),
    .Y(_0604_),
    .A2(net583));
 sg13g2_a21oi_1 _1285_ (.A1(net513),
    .A2(_0604_),
    .Y(_0009_),
    .B1(_0595_));
 sg13g2_xnor2_1 _1286_ (.Y(_0605_),
    .A(\bitserial_cipher.dataq ),
    .B(\bitserial_cipher.state[60] ));
 sg13g2_xor2_1 _1287_ (.B(\bitserial_cipher.state[46] ),
    .A(\bitserial_cipher.state[29] ),
    .X(_0606_));
 sg13g2_xnor2_1 _1288_ (.Y(_0607_),
    .A(_0605_),
    .B(_0606_));
 sg13g2_nand3_1 _1289_ (.B(net613),
    .C(_0607_),
    .A(\bitserial_cipher.state[13] ),
    .Y(_0608_));
 sg13g2_o21ai_1 _1290_ (.B1(net590),
    .Y(_0609_),
    .A1(\bitserial_cipher.state[13] ),
    .A2(_0607_));
 sg13g2_nand2b_1 _1291_ (.Y(_0610_),
    .B(_0608_),
    .A_N(_0609_));
 sg13g2_a22oi_1 _1292_ (.Y(_0611_),
    .B1(net594),
    .B2(net355),
    .A2(net605),
    .A1(\bitserial_cipher.state[2] ));
 sg13g2_a22oi_1 _1293_ (.Y(_0612_),
    .B1(_0610_),
    .B2(_0611_),
    .A2(net583),
    .A1(_0501_));
 sg13g2_mux2_1 _1294_ (.A0(net352),
    .A1(_0612_),
    .S(net513),
    .X(_0010_));
 sg13g2_nor2_1 _1295_ (.A(net321),
    .B(net513),
    .Y(_0613_));
 sg13g2_xnor2_1 _1296_ (.Y(_0614_),
    .A(\bitserial_cipher.state[30] ),
    .B(\bitserial_cipher.state[47] ));
 sg13g2_xor2_1 _1297_ (.B(\bitserial_cipher.state[61] ),
    .A(\bitserial_cipher.state[14] ),
    .X(_0615_));
 sg13g2_xnor2_1 _1298_ (.Y(_0616_),
    .A(_0614_),
    .B(_0615_));
 sg13g2_a22oi_1 _1299_ (.Y(_0617_),
    .B1(net593),
    .B2(net310),
    .A2(net609),
    .A1(\bitserial_cipher.state[3] ));
 sg13g2_inv_1 _1300_ (.Y(_0618_),
    .A(_0617_));
 sg13g2_a221oi_1 _1301_ (.B2(net613),
    .C1(_0618_),
    .B1(_0616_),
    .A1(net352),
    .Y(_0619_),
    .A2(net583));
 sg13g2_a21oi_1 _1302_ (.A1(net513),
    .A2(net353),
    .Y(_0011_),
    .B1(_0613_));
 sg13g2_a22oi_1 _1303_ (.Y(_0620_),
    .B1(net592),
    .B2(\bitserial_cipher.state[24] ),
    .A2(net612),
    .A1(\bitserial_cipher.state[12] ));
 sg13g2_a22oi_1 _1304_ (.Y(_0621_),
    .B1(net582),
    .B2(net303),
    .A2(net604),
    .A1(net215));
 sg13g2_nand3_1 _1305_ (.B(_0620_),
    .C(_0621_),
    .A(net511),
    .Y(_0622_));
 sg13g2_o21ai_1 _1306_ (.B1(_0622_),
    .Y(_0623_),
    .A1(net358),
    .A2(net511));
 sg13g2_inv_1 _1307_ (.Y(_0012_),
    .A(net359));
 sg13g2_nor2_1 _1308_ (.A(net356),
    .B(net511),
    .Y(_0624_));
 sg13g2_a22oi_1 _1309_ (.Y(_0625_),
    .B1(net591),
    .B2(net293),
    .A2(net612),
    .A1(\bitserial_cipher.state[13] ));
 sg13g2_inv_1 _1310_ (.Y(_0626_),
    .A(_0625_));
 sg13g2_a221oi_1 _1311_ (.B2(\bitserial_cipher.state[28] ),
    .C1(_0626_),
    .B1(net582),
    .A1(net301),
    .Y(_0627_),
    .A2(net603));
 sg13g2_a21oi_1 _1312_ (.A1(net511),
    .A2(_0627_),
    .Y(_0013_),
    .B1(_0624_));
 sg13g2_a22oi_1 _1313_ (.Y(_0628_),
    .B1(net591),
    .B2(net295),
    .A2(net612),
    .A1(\bitserial_cipher.state[14] ));
 sg13g2_a22oi_1 _1314_ (.Y(_0629_),
    .B1(net582),
    .B2(\bitserial_cipher.state[29] ),
    .A2(net602),
    .A1(net335));
 sg13g2_nand3_1 _1315_ (.B(_0628_),
    .C(_0629_),
    .A(net511),
    .Y(_0630_));
 sg13g2_o21ai_1 _1316_ (.B1(_0630_),
    .Y(_0631_),
    .A1(net342),
    .A2(net511));
 sg13g2_inv_1 _1317_ (.Y(_0014_),
    .A(_0631_));
 sg13g2_and2_1 _1318_ (.A(\bitserial_cipher.state[15] ),
    .B(net612),
    .X(_0632_));
 sg13g2_a221oi_1 _1319_ (.B2(net303),
    .C1(_0632_),
    .B1(net592),
    .A1(net285),
    .Y(_0633_),
    .A2(net603));
 sg13g2_nor2_1 _1320_ (.A(net291),
    .B(net512),
    .Y(_0634_));
 sg13g2_o21ai_1 _1321_ (.B1(net582),
    .Y(_0635_),
    .A1(net342),
    .A2(net553));
 sg13g2_a21oi_1 _1322_ (.A1(_0633_),
    .A2(_0635_),
    .Y(_0015_),
    .B1(_0634_));
 sg13g2_nor3_2 _1323_ (.A(net615),
    .B(net611),
    .C(_0555_),
    .Y(_0636_));
 sg13g2_a21oi_2 _1324_ (.B1(net607),
    .Y(_0637_),
    .A2(_0636_),
    .A1(_0559_));
 sg13g2_xor2_1 _1325_ (.B(\bitserial_cipher.rc[4] ),
    .A(\bitserial_cipher.rc[5] ),
    .X(_0638_));
 sg13g2_a22oi_1 _1326_ (.Y(_0639_),
    .B1(_0638_),
    .B2(net607),
    .A2(_0637_),
    .A1(net32));
 sg13g2_inv_1 _1327_ (.Y(_0016_),
    .A(net33));
 sg13g2_a22oi_1 _1328_ (.Y(_0640_),
    .B1(_0637_),
    .B2(\bitserial_cipher.rc[1] ),
    .A2(net607),
    .A1(net28));
 sg13g2_inv_1 _1329_ (.Y(_0017_),
    .A(net29));
 sg13g2_a22oi_1 _1330_ (.Y(_0641_),
    .B1(_0637_),
    .B2(net45),
    .A2(net607),
    .A1(\bitserial_cipher.rc[1] ));
 sg13g2_inv_1 _1331_ (.Y(_0018_),
    .A(net46));
 sg13g2_a22oi_1 _1332_ (.Y(_0642_),
    .B1(_0637_),
    .B2(net43),
    .A2(net607),
    .A1(\bitserial_cipher.rc[2] ));
 sg13g2_inv_1 _1333_ (.Y(_0019_),
    .A(net44));
 sg13g2_a22oi_1 _1334_ (.Y(_0643_),
    .B1(_0637_),
    .B2(net174),
    .A2(net607),
    .A1(net43));
 sg13g2_inv_1 _1335_ (.Y(_0020_),
    .A(_0643_));
 sg13g2_a22oi_1 _1336_ (.Y(_0644_),
    .B1(_0637_),
    .B2(net65),
    .A2(net607),
    .A1(\bitserial_cipher.rc[4] ));
 sg13g2_inv_1 _1337_ (.Y(_0021_),
    .A(net66));
 sg13g2_a22oi_1 _1338_ (.Y(_0645_),
    .B1(_0564_),
    .B2(net277),
    .A2(net595),
    .A1(net47));
 sg13g2_a22oi_1 _1339_ (.Y(_0646_),
    .B1(_0569_),
    .B2(\bitserial_cipher.state[60] ),
    .A2(net613),
    .A1(\bitserial_cipher.state[44] ));
 sg13g2_o21ai_1 _1340_ (.B1(_0646_),
    .Y(_0022_),
    .A1(_0569_),
    .A2(_0645_));
 sg13g2_a22oi_1 _1341_ (.Y(_0647_),
    .B1(_0564_),
    .B2(\bitserial_cipher.state[60] ),
    .A2(net595),
    .A1(net34));
 sg13g2_a22oi_1 _1342_ (.Y(_0648_),
    .B1(_0569_),
    .B2(\bitserial_cipher.state[61] ),
    .A2(net614),
    .A1(net337));
 sg13g2_o21ai_1 _1343_ (.B1(net338),
    .Y(_0023_),
    .A1(_0569_),
    .A2(_0647_));
 sg13g2_a22oi_1 _1344_ (.Y(_0649_),
    .B1(_0564_),
    .B2(\bitserial_cipher.state[61] ),
    .A2(net595),
    .A1(net81));
 sg13g2_a22oi_1 _1345_ (.Y(_0650_),
    .B1(_0569_),
    .B2(\bitserial_cipher.state[62] ),
    .A2(net613),
    .A1(net307));
 sg13g2_o21ai_1 _1346_ (.B1(net308),
    .Y(_0024_),
    .A1(_0569_),
    .A2(_0649_));
 sg13g2_nand2_1 _1347_ (.Y(_0651_),
    .A(net162),
    .B(net613));
 sg13g2_a221oi_1 _1348_ (.B2(\bitserial_cipher.state[62] ),
    .C1(_0569_),
    .B1(_0564_),
    .A1(net277),
    .Y(_0652_),
    .A2(net595));
 sg13g2_a22oi_1 _1349_ (.Y(_0025_),
    .B1(_0651_),
    .B2(_0652_),
    .A2(_0569_),
    .A1(_0504_));
 sg13g2_nand2_1 _1350_ (.Y(_0653_),
    .A(_0561_),
    .B(net589));
 sg13g2_nor2_1 _1351_ (.A(net579),
    .B(net584),
    .Y(_0654_));
 sg13g2_nand2b_2 _1352_ (.Y(_0655_),
    .B(net590),
    .A_N(net581));
 sg13g2_a22oi_1 _1353_ (.Y(_0656_),
    .B1(net589),
    .B2(\bitserial_cipher.state[3] ),
    .A2(net594),
    .A1(net117));
 sg13g2_a22oi_1 _1354_ (.Y(_0657_),
    .B1(net551),
    .B2(net263),
    .A2(net606),
    .A1(\bitserial_cipher.state[8] ));
 sg13g2_o21ai_1 _1355_ (.B1(net264),
    .Y(_0026_),
    .A1(net550),
    .A2(_0656_));
 sg13g2_nor2_1 _1356_ (.A(net316),
    .B(_0655_),
    .Y(_0658_));
 sg13g2_nor2_1 _1357_ (.A(_0505_),
    .B(net598),
    .Y(_0659_));
 sg13g2_a221oi_1 _1358_ (.B2(net263),
    .C1(_0659_),
    .B1(net589),
    .A1(\bitserial_cipher.state[9] ),
    .Y(_0660_),
    .A2(net606));
 sg13g2_a21oi_1 _1359_ (.A1(_0655_),
    .A2(_0660_),
    .Y(_0027_),
    .B1(_0658_));
 sg13g2_a22oi_1 _1360_ (.Y(_0661_),
    .B1(net590),
    .B2(\bitserial_cipher.state[5] ),
    .A2(net594),
    .A1(\bitserial_cipher.state[2] ));
 sg13g2_a22oi_1 _1361_ (.Y(_0662_),
    .B1(net549),
    .B2(net298),
    .A2(net605),
    .A1(net280));
 sg13g2_o21ai_1 _1362_ (.B1(_0662_),
    .Y(_0028_),
    .A1(net549),
    .A2(_0661_));
 sg13g2_a22oi_1 _1363_ (.Y(_0663_),
    .B1(net590),
    .B2(net298),
    .A2(net594),
    .A1(net313));
 sg13g2_a22oi_1 _1364_ (.Y(_0664_),
    .B1(net549),
    .B2(net334),
    .A2(net605),
    .A1(net310));
 sg13g2_o21ai_1 _1365_ (.B1(_0664_),
    .Y(_0029_),
    .A1(net549),
    .A2(_0663_));
 sg13g2_nand2_1 _1366_ (.Y(_0665_),
    .A(net266),
    .B(net589));
 sg13g2_a22oi_1 _1367_ (.Y(_0666_),
    .B1(net589),
    .B2(\bitserial_cipher.state[7] ),
    .A2(net596),
    .A1(net263));
 sg13g2_a22oi_1 _1368_ (.Y(_0667_),
    .B1(net550),
    .B2(net266),
    .A2(net606),
    .A1(\bitserial_cipher.state[12] ));
 sg13g2_o21ai_1 _1369_ (.B1(net267),
    .Y(_0030_),
    .A1(net550),
    .A2(_0666_));
 sg13g2_a22oi_1 _1370_ (.Y(_0668_),
    .B1(net594),
    .B2(net316),
    .A2(net605),
    .A1(\bitserial_cipher.state[13] ));
 sg13g2_a21oi_1 _1371_ (.A1(_0665_),
    .A2(_0668_),
    .Y(_0669_),
    .B1(net550));
 sg13g2_a21o_1 _1372_ (.A2(net550),
    .A1(net333),
    .B1(_0669_),
    .X(_0031_));
 sg13g2_a22oi_1 _1373_ (.Y(_0670_),
    .B1(net590),
    .B2(\bitserial_cipher.state[9] ),
    .A2(net594),
    .A1(\bitserial_cipher.state[6] ));
 sg13g2_a22oi_1 _1374_ (.Y(_0671_),
    .B1(net549),
    .B2(net280),
    .A2(net605),
    .A1(\bitserial_cipher.state[14] ));
 sg13g2_o21ai_1 _1375_ (.B1(net281),
    .Y(_0032_),
    .A1(net549),
    .A2(_0670_));
 sg13g2_a22oi_1 _1376_ (.Y(_0672_),
    .B1(net590),
    .B2(net280),
    .A2(net593),
    .A1(\bitserial_cipher.state[7] ));
 sg13g2_a22oi_1 _1377_ (.Y(_0673_),
    .B1(net549),
    .B2(net310),
    .A2(net609),
    .A1(\bitserial_cipher.state[15] ));
 sg13g2_o21ai_1 _1378_ (.B1(net311),
    .Y(_0033_),
    .A1(net549),
    .A2(_0672_));
 sg13g2_nor2_1 _1379_ (.A(_0502_),
    .B(net597),
    .Y(_0674_));
 sg13g2_a221oi_1 _1380_ (.B2(\bitserial_cipher.state[19] ),
    .C1(_0674_),
    .B1(net586),
    .A1(\bitserial_cipher.state[28] ),
    .Y(_0675_),
    .A2(net602));
 sg13g2_nor2_1 _1381_ (.A(net215),
    .B(_0655_),
    .Y(_0676_));
 sg13g2_a21oi_1 _1382_ (.A1(_0655_),
    .A2(_0675_),
    .Y(_0034_),
    .B1(_0676_));
 sg13g2_a22oi_1 _1383_ (.Y(_0677_),
    .B1(net588),
    .B2(net215),
    .A2(net592),
    .A1(net300));
 sg13g2_a22oi_1 _1384_ (.Y(_0678_),
    .B1(net545),
    .B2(net301),
    .A2(net602),
    .A1(\bitserial_cipher.state[29] ));
 sg13g2_o21ai_1 _1385_ (.B1(net302),
    .Y(_0035_),
    .A1(net545),
    .A2(_0677_));
 sg13g2_a22oi_1 _1386_ (.Y(_0679_),
    .B1(net586),
    .B2(net301),
    .A2(net591),
    .A1(net329));
 sg13g2_a22oi_1 _1387_ (.Y(_0680_),
    .B1(net543),
    .B2(net335),
    .A2(net602),
    .A1(\bitserial_cipher.state[30] ));
 sg13g2_o21ai_1 _1388_ (.B1(net336),
    .Y(_0036_),
    .A1(net543),
    .A2(_0679_));
 sg13g2_a22oi_1 _1389_ (.Y(_0681_),
    .B1(net586),
    .B2(\bitserial_cipher.state[22] ),
    .A2(net591),
    .A1(net274));
 sg13g2_a22oi_1 _1390_ (.Y(_0682_),
    .B1(net544),
    .B2(net285),
    .A2(net603),
    .A1(\bitserial_cipher.state[31] ));
 sg13g2_o21ai_1 _1391_ (.B1(net286),
    .Y(_0037_),
    .A1(net544),
    .A2(_0681_));
 sg13g2_nand2_1 _1392_ (.Y(_0683_),
    .A(\bitserial_cipher.state[24] ),
    .B(net586));
 sg13g2_a22oi_1 _1393_ (.Y(_0684_),
    .B1(net588),
    .B2(net285),
    .A2(net591),
    .A1(net215));
 sg13g2_a22oi_1 _1394_ (.Y(_0685_),
    .B1(net548),
    .B2(\bitserial_cipher.state[24] ),
    .A2(net603),
    .A1(net304));
 sg13g2_o21ai_1 _1395_ (.B1(net305),
    .Y(_0038_),
    .A1(net545),
    .A2(_0684_));
 sg13g2_a22oi_1 _1396_ (.Y(_0686_),
    .B1(net591),
    .B2(\bitserial_cipher.state[21] ),
    .A2(net602),
    .A1(\bitserial_cipher.state[17] ));
 sg13g2_a21oi_1 _1397_ (.A1(_0683_),
    .A2(_0686_),
    .Y(_0687_),
    .B1(net545));
 sg13g2_a21o_1 _1398_ (.A2(net543),
    .A1(net293),
    .B1(_0687_),
    .X(_0039_));
 sg13g2_a22oi_1 _1399_ (.Y(_0688_),
    .B1(net586),
    .B2(net293),
    .A2(net591),
    .A1(\bitserial_cipher.state[22] ));
 sg13g2_a22oi_1 _1400_ (.Y(_0689_),
    .B1(net543),
    .B2(net295),
    .A2(net602),
    .A1(\bitserial_cipher.state[18] ));
 sg13g2_o21ai_1 _1401_ (.B1(net296),
    .Y(_0040_),
    .A1(net543),
    .A2(_0688_));
 sg13g2_a22oi_1 _1402_ (.Y(_0690_),
    .B1(net586),
    .B2(net295),
    .A2(net591),
    .A1(net285));
 sg13g2_a22oi_1 _1403_ (.Y(_0691_),
    .B1(net543),
    .B2(net303),
    .A2(net603),
    .A1(net274));
 sg13g2_o21ai_1 _1404_ (.B1(_0691_),
    .Y(_0041_),
    .A1(net544),
    .A2(_0690_));
 sg13g2_nor2_1 _1405_ (.A(_0502_),
    .B(net585),
    .Y(_0692_));
 sg13g2_a221oi_1 _1406_ (.B2(\bitserial_cipher.state[12] ),
    .C1(net548),
    .B1(net599),
    .A1(\bitserial_cipher.state[24] ),
    .Y(_0693_),
    .A2(net603));
 sg13g2_a22oi_1 _1407_ (.Y(_0694_),
    .B1(_0566_),
    .B2(net321),
    .A2(net610),
    .A1(\bitserial_cipher.state[28] ));
 sg13g2_a22oi_1 _1408_ (.Y(_0042_),
    .B1(_0693_),
    .B2(net322),
    .A2(net548),
    .A1(_0502_));
 sg13g2_a221oi_1 _1409_ (.B2(\bitserial_cipher.state[13] ),
    .C1(_0692_),
    .B1(net599),
    .A1(\bitserial_cipher.state[29] ),
    .Y(_0695_),
    .A2(net610));
 sg13g2_a22oi_1 _1410_ (.Y(_0696_),
    .B1(net545),
    .B2(net300),
    .A2(net602),
    .A1(net293));
 sg13g2_o21ai_1 _1411_ (.B1(_0696_),
    .Y(_0043_),
    .A1(net543),
    .A2(_0695_));
 sg13g2_and2_1 _1412_ (.A(net295),
    .B(net602),
    .X(_0697_));
 sg13g2_a21oi_1 _1413_ (.A1(\bitserial_cipher.state[14] ),
    .A2(net599),
    .Y(_0698_),
    .B1(net545));
 sg13g2_a221oi_1 _1414_ (.B2(net300),
    .C1(_0697_),
    .B1(net586),
    .A1(\bitserial_cipher.state[30] ),
    .Y(_0699_),
    .A2(net610));
 sg13g2_a22oi_1 _1415_ (.Y(_0044_),
    .B1(_0698_),
    .B2(_0699_),
    .A2(net543),
    .A1(_0503_));
 sg13g2_a22oi_1 _1416_ (.Y(_0700_),
    .B1(net599),
    .B2(\bitserial_cipher.state[15] ),
    .A2(net603),
    .A1(\bitserial_cipher.state[27] ));
 sg13g2_a22oi_1 _1417_ (.Y(_0701_),
    .B1(net586),
    .B2(\bitserial_cipher.state[18] ),
    .A2(net610),
    .A1(\bitserial_cipher.state[31] ));
 sg13g2_a21oi_1 _1418_ (.A1(_0700_),
    .A2(_0701_),
    .Y(_0702_),
    .B1(net544));
 sg13g2_a21o_1 _1419_ (.A2(net544),
    .A1(net274),
    .B1(_0702_),
    .X(_0045_));
 sg13g2_nand2_1 _1420_ (.Y(_0703_),
    .A(net117),
    .B(net551));
 sg13g2_nor3_1 _1421_ (.A(_0507_),
    .B(\bitserial_cipher.bcount[1] ),
    .C(\bitserial_cipher.bcount[2] ),
    .Y(_0704_));
 sg13g2_nor2b_1 _1422_ (.A(\bitserial_cipher.bcount[1] ),
    .B_N(\bitserial_cipher.bcount[2] ),
    .Y(_0705_));
 sg13g2_nand2b_1 _1423_ (.Y(_0706_),
    .B(\bitserial_cipher.bcount[0] ),
    .A_N(\bitserial_cipher.rc[0] ));
 sg13g2_nor2_1 _1424_ (.A(\bitserial_cipher.bcount[0] ),
    .B(\bitserial_cipher.bcount[1] ),
    .Y(_0707_));
 sg13g2_and2_1 _1425_ (.A(\bitserial_cipher.bcount[0] ),
    .B(_0705_),
    .X(_0708_));
 sg13g2_a22oi_1 _1426_ (.Y(_0709_),
    .B1(_0705_),
    .B2(_0706_),
    .A2(_0704_),
    .A1(\bitserial_cipher.rc[3] ));
 sg13g2_xnor2_1 _1427_ (.Y(_0710_),
    .A(\bitserial_cipher.state[60] ),
    .B(_0709_));
 sg13g2_xor2_1 _1428_ (.B(_0709_),
    .A(\bitserial_cipher.state[60] ),
    .X(_0711_));
 sg13g2_or4_1 _1429_ (.A(_0457_),
    .B(_0507_),
    .C(\bitserial_cipher.bcount[1] ),
    .D(\bitserial_cipher.bcount[2] ),
    .X(_0712_));
 sg13g2_nand2_1 _1430_ (.Y(_0713_),
    .A(\bitserial_cipher.bcount[3] ),
    .B(_0707_));
 sg13g2_nand3_1 _1431_ (.B(\bitserial_cipher.bcount[0] ),
    .C(_0705_),
    .A(\bitserial_cipher.rc[1] ),
    .Y(_0714_));
 sg13g2_nand3_1 _1432_ (.B(_0713_),
    .C(_0714_),
    .A(_0712_),
    .Y(_0715_));
 sg13g2_xor2_1 _1433_ (.B(_0715_),
    .A(\bitserial_cipher.state[61] ),
    .X(_0716_));
 sg13g2_xnor2_1 _1434_ (.Y(_0717_),
    .A(\bitserial_cipher.state[61] ),
    .B(_0715_));
 sg13g2_nand2_1 _1435_ (.Y(_0718_),
    .A(_0711_),
    .B(_0717_));
 sg13g2_a22oi_1 _1436_ (.Y(_0719_),
    .B1(_0708_),
    .B2(\bitserial_cipher.rc[2] ),
    .A2(_0704_),
    .A1(\bitserial_cipher.rc[5] ));
 sg13g2_xor2_1 _1437_ (.B(_0719_),
    .A(\bitserial_cipher.state[62] ),
    .X(_0720_));
 sg13g2_nor2_1 _1438_ (.A(_0711_),
    .B(_0717_),
    .Y(_0721_));
 sg13g2_nand2b_1 _1439_ (.Y(_0722_),
    .B(_0711_),
    .A_N(_0720_));
 sg13g2_nor2_1 _1440_ (.A(_0716_),
    .B(_0720_),
    .Y(_0723_));
 sg13g2_a21oi_1 _1441_ (.A1(_0710_),
    .A2(_0716_),
    .Y(_0724_),
    .B1(_0720_));
 sg13g2_a22oi_1 _1442_ (.Y(_0725_),
    .B1(_0724_),
    .B2(_0718_),
    .A2(_0720_),
    .A1(_0711_));
 sg13g2_nor3_2 _1443_ (.A(\bitserial_cipher.bcount[0] ),
    .B(\bitserial_cipher.bcount[1] ),
    .C(\bitserial_cipher.bcount[3] ),
    .Y(_0726_));
 sg13g2_xnor2_1 _1444_ (.Y(_0727_),
    .A(\bitserial_cipher.dataq ),
    .B(_0726_));
 sg13g2_xnor2_1 _1445_ (.Y(_0728_),
    .A(_0504_),
    .B(_0726_));
 sg13g2_nor2_2 _1446_ (.A(_0557_),
    .B(_0558_),
    .Y(_0729_));
 sg13g2_nand2_1 _1447_ (.Y(_0730_),
    .A(_0555_),
    .B(_0729_));
 sg13g2_inv_1 _1448_ (.Y(_0731_),
    .A(_0730_));
 sg13g2_and3_1 _1449_ (.X(_0732_),
    .A(_0555_),
    .B(_0557_),
    .C(_0558_));
 sg13g2_nand3_1 _1450_ (.B(_0557_),
    .C(_0558_),
    .A(_0555_),
    .Y(_0733_));
 sg13g2_xnor2_1 _1451_ (.Y(_0734_),
    .A(\bitserial_cipher.key[124] ),
    .B(\bitserial_cipher.state[60] ));
 sg13g2_a22oi_1 _1452_ (.Y(_0735_),
    .B1(net606),
    .B2(net365),
    .A2(_0525_),
    .A1(\bitserial_cipher.state[12] ));
 sg13g2_xnor2_1 _1453_ (.Y(_0736_),
    .A(_0725_),
    .B(_0727_));
 sg13g2_o21ai_1 _1454_ (.B1(_0735_),
    .Y(_0737_),
    .A1(net569),
    .A2(_0734_));
 sg13g2_a221oi_1 _1455_ (.B2(_0736_),
    .C1(_0737_),
    .B1(_0731_),
    .A1(_0561_),
    .Y(_0738_),
    .A2(net589));
 sg13g2_o21ai_1 _1456_ (.B1(_0655_),
    .Y(_0739_),
    .A1(net1),
    .A2(_0653_));
 sg13g2_o21ai_1 _1457_ (.B1(_0703_),
    .Y(_0046_),
    .A1(_0738_),
    .A2(_0739_));
 sg13g2_a21oi_1 _1458_ (.A1(_0720_),
    .A2(_0721_),
    .Y(_0740_),
    .B1(_0730_));
 sg13g2_nand3_1 _1459_ (.B(_0728_),
    .C(_0740_),
    .A(_0722_),
    .Y(_0741_));
 sg13g2_o21ai_1 _1460_ (.B1(_0716_),
    .Y(_0742_),
    .A1(_0711_),
    .A2(_0720_));
 sg13g2_nor3_1 _1461_ (.A(_0728_),
    .B(_0730_),
    .C(_0742_),
    .Y(_0743_));
 sg13g2_xnor2_1 _1462_ (.Y(_0744_),
    .A(\bitserial_cipher.key[125] ),
    .B(\bitserial_cipher.state[61] ));
 sg13g2_nor2_1 _1463_ (.A(_0501_),
    .B(_0526_),
    .Y(_0745_));
 sg13g2_a221oi_1 _1464_ (.B2(\bitserial_cipher.state[0] ),
    .C1(_0745_),
    .B1(net589),
    .A1(\bitserial_cipher.state[5] ),
    .Y(_0746_),
    .A2(net607));
 sg13g2_o21ai_1 _1465_ (.B1(_0746_),
    .Y(_0747_),
    .A1(net569),
    .A2(_0744_));
 sg13g2_nor3_1 _1466_ (.A(net551),
    .B(_0743_),
    .C(_0747_),
    .Y(_0748_));
 sg13g2_a22oi_1 _1467_ (.Y(_0047_),
    .B1(_0741_),
    .B2(_0748_),
    .A2(net550),
    .A1(_0505_));
 sg13g2_nand2_1 _1468_ (.Y(_0749_),
    .A(_0718_),
    .B(_0720_));
 sg13g2_nor2_1 _1469_ (.A(_0723_),
    .B(_0727_),
    .Y(_0750_));
 sg13g2_a22oi_1 _1470_ (.Y(_0751_),
    .B1(_0749_),
    .B2(_0750_),
    .A2(_0727_),
    .A1(_0724_));
 sg13g2_xor2_1 _1471_ (.B(\bitserial_cipher.state[62] ),
    .A(\bitserial_cipher.key[126] ),
    .X(_0752_));
 sg13g2_a22oi_1 _1472_ (.Y(_0753_),
    .B1(net605),
    .B2(\bitserial_cipher.state[6] ),
    .A2(_0525_),
    .A1(\bitserial_cipher.state[14] ));
 sg13g2_inv_1 _1473_ (.Y(_0754_),
    .A(_0753_));
 sg13g2_a221oi_1 _1474_ (.B2(net576),
    .C1(_0754_),
    .B1(_0752_),
    .A1(_0740_),
    .Y(_0755_),
    .A2(_0751_));
 sg13g2_a21oi_1 _1475_ (.A1(\bitserial_cipher.state[1] ),
    .A2(net589),
    .Y(_0756_),
    .B1(net550));
 sg13g2_a22oi_1 _1476_ (.Y(_0048_),
    .B1(_0755_),
    .B2(_0756_),
    .A2(net550),
    .A1(_0506_));
 sg13g2_a21o_1 _1477_ (.A2(_0720_),
    .A1(_0711_),
    .B1(_0717_),
    .X(_0757_));
 sg13g2_xnor2_1 _1478_ (.Y(_0758_),
    .A(\bitserial_cipher.key[127] ),
    .B(\bitserial_cipher.dataq ));
 sg13g2_a22oi_1 _1479_ (.Y(_0759_),
    .B1(net605),
    .B2(\bitserial_cipher.state[7] ),
    .A2(net610),
    .A1(\bitserial_cipher.state[15] ));
 sg13g2_o21ai_1 _1480_ (.B1(_0759_),
    .Y(_0760_),
    .A1(net560),
    .A2(_0758_));
 sg13g2_a21oi_1 _1481_ (.A1(_0711_),
    .A2(_0717_),
    .Y(_0761_),
    .B1(_0728_));
 sg13g2_a221oi_1 _1482_ (.B2(_0761_),
    .C1(_0730_),
    .B1(_0757_),
    .A1(_0728_),
    .Y(_0762_),
    .A2(_0749_));
 sg13g2_nor2_1 _1483_ (.A(_0760_),
    .B(_0762_),
    .Y(_0763_));
 sg13g2_a22oi_1 _1484_ (.Y(_0764_),
    .B1(net552),
    .B2(net313),
    .A2(net581),
    .A1(\bitserial_cipher.state[2] ));
 sg13g2_nand2_1 _1485_ (.Y(_0049_),
    .A(_0763_),
    .B(net314));
 sg13g2_and2_1 _1486_ (.A(net616),
    .B(_0531_),
    .X(_0765_));
 sg13g2_nor2_2 _1487_ (.A(_0456_),
    .B(_0765_),
    .Y(_0766_));
 sg13g2_a21oi_1 _1488_ (.A1(_0456_),
    .A2(_0531_),
    .Y(_0050_),
    .B1(_0766_));
 sg13g2_o21ai_1 _1489_ (.B1(net616),
    .Y(_0767_),
    .A1(net232),
    .A2(_0766_));
 sg13g2_a21oi_1 _1490_ (.A1(net232),
    .A2(_0766_),
    .Y(_0051_),
    .B1(_0767_));
 sg13g2_nand3_1 _1491_ (.B(\bitserial_cipher.scount[0] ),
    .C(net40),
    .A(\bitserial_cipher.scount[1] ),
    .Y(_0768_));
 sg13g2_a21oi_1 _1492_ (.A1(_0533_),
    .A2(_0768_),
    .Y(_0769_),
    .B1(_0765_));
 sg13g2_a21oi_1 _1493_ (.A1(\bitserial_cipher.scount[1] ),
    .A2(_0766_),
    .Y(_0770_),
    .B1(net40));
 sg13g2_nor2_1 _1494_ (.A(_0769_),
    .B(net41),
    .Y(_0052_));
 sg13g2_nor2_1 _1495_ (.A(_0531_),
    .B(_0768_),
    .Y(_0771_));
 sg13g2_nor2_1 _1496_ (.A(net30),
    .B(_0771_),
    .Y(_0772_));
 sg13g2_a21oi_1 _1497_ (.A1(net30),
    .A2(_0769_),
    .Y(_0053_),
    .B1(_0772_));
 sg13g2_o21ai_1 _1498_ (.B1(net616),
    .Y(_0773_),
    .A1(_0507_),
    .A2(net598));
 sg13g2_a21oi_1 _1499_ (.A1(_0507_),
    .A2(net598),
    .Y(_0054_),
    .B1(_0773_));
 sg13g2_nand2_1 _1500_ (.Y(_0774_),
    .A(net616),
    .B(net598));
 sg13g2_nand3_1 _1501_ (.B(net616),
    .C(net598),
    .A(net348),
    .Y(_0775_));
 sg13g2_or2_1 _1502_ (.X(_0776_),
    .B(_0707_),
    .A(net597));
 sg13g2_o21ai_1 _1503_ (.B1(_0775_),
    .Y(_0055_),
    .A1(_0512_),
    .A2(_0776_));
 sg13g2_a21oi_1 _1504_ (.A1(net616),
    .A2(net597),
    .Y(_0777_),
    .B1(_0513_));
 sg13g2_nand2_1 _1505_ (.Y(_0778_),
    .A(\bitserial_cipher.bcount[2] ),
    .B(_0777_));
 sg13g2_nor2_1 _1506_ (.A(_0540_),
    .B(net601),
    .Y(_0779_));
 sg13g2_xnor2_1 _1507_ (.Y(_0780_),
    .A(net354),
    .B(_0777_));
 sg13g2_a21oi_1 _1508_ (.A1(_0774_),
    .A2(_0779_),
    .Y(_0056_),
    .B1(_0780_));
 sg13g2_nand2_1 _1509_ (.Y(_0781_),
    .A(_0514_),
    .B(_0549_));
 sg13g2_a22oi_1 _1510_ (.Y(_0057_),
    .B1(_0781_),
    .B2(_0774_),
    .A2(_0778_),
    .A1(_0508_));
 sg13g2_nand2_2 _1511_ (.Y(_0782_),
    .A(_0636_),
    .B(_0729_));
 sg13g2_a21oi_1 _1512_ (.A1(_0636_),
    .A2(_0729_),
    .Y(_0783_),
    .B1(net577));
 sg13g2_nand2_1 _1513_ (.Y(_0784_),
    .A(net556),
    .B(net522));
 sg13g2_a22oi_1 _1514_ (.Y(_0785_),
    .B1(net519),
    .B2(net77),
    .A2(net576),
    .A1(\bitserial_cipher.key[124] ));
 sg13g2_inv_1 _1515_ (.Y(_0058_),
    .A(net78));
 sg13g2_nor3_1 _1516_ (.A(net77),
    .B(net573),
    .C(net536),
    .Y(_0786_));
 sg13g2_nor2_1 _1517_ (.A(net132),
    .B(net574),
    .Y(_0787_));
 sg13g2_a221oi_1 _1518_ (.B2(_0787_),
    .C1(_0786_),
    .B1(net536),
    .A1(_0497_),
    .Y(_0059_),
    .A2(net576));
 sg13g2_nor2_1 _1519_ (.A(net160),
    .B(net501),
    .Y(_0788_));
 sg13g2_nor3_1 _1520_ (.A(net132),
    .B(net572),
    .C(net536),
    .Y(_0789_));
 sg13g2_nor2_1 _1521_ (.A(net276),
    .B(net569),
    .Y(_0790_));
 sg13g2_nor3_1 _1522_ (.A(_0788_),
    .B(_0789_),
    .C(_0790_),
    .Y(_0060_));
 sg13g2_nor2_1 _1523_ (.A(net160),
    .B(net529),
    .Y(_0791_));
 sg13g2_nor2_1 _1524_ (.A(net113),
    .B(net573),
    .Y(_0792_));
 sg13g2_a221oi_1 _1525_ (.B2(_0792_),
    .C1(_0791_),
    .B1(net528),
    .A1(_0498_),
    .Y(_0061_),
    .A2(net573));
 sg13g2_nor2_1 _1526_ (.A(net103),
    .B(net501),
    .Y(_0793_));
 sg13g2_nor2b_1 _1527_ (.A(net529),
    .B_N(_0792_),
    .Y(_0794_));
 sg13g2_nor2_1 _1528_ (.A(net77),
    .B(net561),
    .Y(_0795_));
 sg13g2_nor3_1 _1529_ (.A(_0793_),
    .B(_0794_),
    .C(_0795_),
    .Y(_0062_));
 sg13g2_nor2_1 _1530_ (.A(net103),
    .B(net529),
    .Y(_0796_));
 sg13g2_a221oi_1 _1531_ (.B2(_0495_),
    .C1(_0796_),
    .B1(net515),
    .A1(_0496_),
    .Y(_0063_),
    .A2(net572));
 sg13g2_nor2_1 _1532_ (.A(\bitserial_cipher.key[6] ),
    .B(net501),
    .Y(_0797_));
 sg13g2_nor2_1 _1533_ (.A(\bitserial_cipher.key[2] ),
    .B(net559),
    .Y(_0798_));
 sg13g2_nor2_1 _1534_ (.A(net38),
    .B(net529),
    .Y(_0799_));
 sg13g2_nor3_1 _1535_ (.A(_0797_),
    .B(_0798_),
    .C(_0799_),
    .Y(_0064_));
 sg13g2_nor2_1 _1536_ (.A(\bitserial_cipher.key[7] ),
    .B(net501),
    .Y(_0800_));
 sg13g2_nor2_1 _1537_ (.A(\bitserial_cipher.key[6] ),
    .B(net528),
    .Y(_0801_));
 sg13g2_nor2_1 _1538_ (.A(net113),
    .B(net561),
    .Y(_0802_));
 sg13g2_nor3_1 _1539_ (.A(_0800_),
    .B(_0801_),
    .C(_0802_),
    .Y(_0065_));
 sg13g2_nor2_1 _1540_ (.A(\bitserial_cipher.key[8] ),
    .B(net501),
    .Y(_0803_));
 sg13g2_nor2_1 _1541_ (.A(\bitserial_cipher.key[7] ),
    .B(net528),
    .Y(_0804_));
 sg13g2_nor2_1 _1542_ (.A(net103),
    .B(net561),
    .Y(_0805_));
 sg13g2_nor3_1 _1543_ (.A(_0803_),
    .B(_0804_),
    .C(_0805_),
    .Y(_0066_));
 sg13g2_nor2_1 _1544_ (.A(net191),
    .B(net528),
    .Y(_0806_));
 sg13g2_a221oi_1 _1545_ (.B2(_0494_),
    .C1(_0806_),
    .B1(net515),
    .A1(_0495_),
    .Y(_0067_),
    .A2(net572));
 sg13g2_nor2_1 _1546_ (.A(\bitserial_cipher.key[10] ),
    .B(net500),
    .Y(_0807_));
 sg13g2_nor2_1 _1547_ (.A(net203),
    .B(net524),
    .Y(_0808_));
 sg13g2_nor2_1 _1548_ (.A(\bitserial_cipher.key[6] ),
    .B(net559),
    .Y(_0809_));
 sg13g2_nor3_1 _1549_ (.A(_0807_),
    .B(_0808_),
    .C(_0809_),
    .Y(_0068_));
 sg13g2_nor2_1 _1550_ (.A(\bitserial_cipher.key[11] ),
    .B(net502),
    .Y(_0810_));
 sg13g2_nor2_1 _1551_ (.A(\bitserial_cipher.key[10] ),
    .B(net528),
    .Y(_0811_));
 sg13g2_nor2_1 _1552_ (.A(net245),
    .B(net561),
    .Y(_0812_));
 sg13g2_nor3_1 _1553_ (.A(_0810_),
    .B(_0811_),
    .C(_0812_),
    .Y(_0069_));
 sg13g2_nor2_1 _1554_ (.A(net195),
    .B(net502),
    .Y(_0813_));
 sg13g2_nor2_1 _1555_ (.A(net191),
    .B(net559),
    .Y(_0814_));
 sg13g2_nor2_1 _1556_ (.A(net273),
    .B(net528),
    .Y(_0815_));
 sg13g2_nor3_1 _1557_ (.A(_0813_),
    .B(_0814_),
    .C(_0815_),
    .Y(_0070_));
 sg13g2_nor2_1 _1558_ (.A(net195),
    .B(net527),
    .Y(_0816_));
 sg13g2_a221oi_1 _1559_ (.B2(_0493_),
    .C1(_0816_),
    .B1(net514),
    .A1(_0494_),
    .Y(_0071_),
    .A2(net571));
 sg13g2_nor2_1 _1560_ (.A(\bitserial_cipher.key[14] ),
    .B(net502),
    .Y(_0817_));
 sg13g2_nor2_1 _1561_ (.A(\bitserial_cipher.key[10] ),
    .B(net559),
    .Y(_0818_));
 sg13g2_nor2_1 _1562_ (.A(net83),
    .B(net528),
    .Y(_0819_));
 sg13g2_nor3_1 _1563_ (.A(_0817_),
    .B(_0818_),
    .C(_0819_),
    .Y(_0072_));
 sg13g2_nor2_1 _1564_ (.A(\bitserial_cipher.key[15] ),
    .B(net499),
    .Y(_0820_));
 sg13g2_nor2_1 _1565_ (.A(\bitserial_cipher.key[11] ),
    .B(net561),
    .Y(_0821_));
 sg13g2_nor2_1 _1566_ (.A(net158),
    .B(net528),
    .Y(_0822_));
 sg13g2_nor3_1 _1567_ (.A(_0820_),
    .B(_0821_),
    .C(_0822_),
    .Y(_0073_));
 sg13g2_nor2_1 _1568_ (.A(\bitserial_cipher.key[16] ),
    .B(net498),
    .Y(_0823_));
 sg13g2_nor2_1 _1569_ (.A(\bitserial_cipher.key[15] ),
    .B(net527),
    .Y(_0824_));
 sg13g2_nor2_1 _1570_ (.A(net195),
    .B(net560),
    .Y(_0825_));
 sg13g2_nor3_1 _1571_ (.A(_0823_),
    .B(_0824_),
    .C(_0825_),
    .Y(_0074_));
 sg13g2_nor2_1 _1572_ (.A(net254),
    .B(net527),
    .Y(_0826_));
 sg13g2_a221oi_1 _1573_ (.B2(_0492_),
    .C1(_0826_),
    .B1(net515),
    .A1(_0493_),
    .Y(_0075_),
    .A2(net571));
 sg13g2_nor2_1 _1574_ (.A(\bitserial_cipher.key[18] ),
    .B(net499),
    .Y(_0827_));
 sg13g2_nor2_1 _1575_ (.A(\bitserial_cipher.key[14] ),
    .B(net560),
    .Y(_0828_));
 sg13g2_nor2_1 _1576_ (.A(net59),
    .B(net527),
    .Y(_0829_));
 sg13g2_nor3_1 _1577_ (.A(_0827_),
    .B(_0828_),
    .C(_0829_),
    .Y(_0076_));
 sg13g2_nor2_1 _1578_ (.A(net258),
    .B(net498),
    .Y(_0830_));
 sg13g2_nor2_1 _1579_ (.A(\bitserial_cipher.key[18] ),
    .B(net530),
    .Y(_0831_));
 sg13g2_nor2_1 _1580_ (.A(net261),
    .B(net560),
    .Y(_0832_));
 sg13g2_nor3_1 _1581_ (.A(_0830_),
    .B(_0831_),
    .C(_0832_),
    .Y(_0077_));
 sg13g2_nor2_1 _1582_ (.A(net149),
    .B(net498),
    .Y(_0833_));
 sg13g2_nor2_1 _1583_ (.A(net258),
    .B(net526),
    .Y(_0834_));
 sg13g2_nor2_1 _1584_ (.A(net254),
    .B(net560),
    .Y(_0835_));
 sg13g2_nor3_1 _1585_ (.A(_0833_),
    .B(_0834_),
    .C(_0835_),
    .Y(_0078_));
 sg13g2_nor2_1 _1586_ (.A(net149),
    .B(net526),
    .Y(_0836_));
 sg13g2_a221oi_1 _1587_ (.B2(_0491_),
    .C1(_0836_),
    .B1(net515),
    .A1(_0492_),
    .Y(_0079_),
    .A2(net572));
 sg13g2_nor2_1 _1588_ (.A(\bitserial_cipher.key[22] ),
    .B(net498),
    .Y(_0837_));
 sg13g2_nor2_1 _1589_ (.A(\bitserial_cipher.key[18] ),
    .B(net560),
    .Y(_0838_));
 sg13g2_nor2_1 _1590_ (.A(net133),
    .B(net526),
    .Y(_0839_));
 sg13g2_nor3_1 _1591_ (.A(_0837_),
    .B(_0838_),
    .C(_0839_),
    .Y(_0080_));
 sg13g2_nor2_1 _1592_ (.A(net209),
    .B(net498),
    .Y(_0840_));
 sg13g2_nor2_1 _1593_ (.A(net258),
    .B(net560),
    .Y(_0841_));
 sg13g2_nor2_1 _1594_ (.A(net163),
    .B(net526),
    .Y(_0842_));
 sg13g2_nor3_1 _1595_ (.A(_0840_),
    .B(_0841_),
    .C(_0842_),
    .Y(_0081_));
 sg13g2_nor2_1 _1596_ (.A(net208),
    .B(net498),
    .Y(_0843_));
 sg13g2_nor2_1 _1597_ (.A(net209),
    .B(net526),
    .Y(_0844_));
 sg13g2_nor2_1 _1598_ (.A(net149),
    .B(net560),
    .Y(_0845_));
 sg13g2_nor3_1 _1599_ (.A(_0843_),
    .B(_0844_),
    .C(_0845_),
    .Y(_0082_));
 sg13g2_nor2_1 _1600_ (.A(net208),
    .B(net526),
    .Y(_0846_));
 sg13g2_a221oi_1 _1601_ (.B2(_0490_),
    .C1(_0846_),
    .B1(net514),
    .A1(_0491_),
    .Y(_0083_),
    .A2(net572));
 sg13g2_nor2_1 _1602_ (.A(\bitserial_cipher.key[26] ),
    .B(net498),
    .Y(_0847_));
 sg13g2_nor2_1 _1603_ (.A(\bitserial_cipher.key[25] ),
    .B(net526),
    .Y(_0848_));
 sg13g2_nor2_1 _1604_ (.A(net163),
    .B(net557),
    .Y(_0849_));
 sg13g2_nor3_1 _1605_ (.A(_0847_),
    .B(_0848_),
    .C(_0849_),
    .Y(_0084_));
 sg13g2_nor2_1 _1606_ (.A(net139),
    .B(net498),
    .Y(_0850_));
 sg13g2_nor2_1 _1607_ (.A(\bitserial_cipher.key[26] ),
    .B(net526),
    .Y(_0851_));
 sg13g2_nor2_1 _1608_ (.A(net209),
    .B(net557),
    .Y(_0852_));
 sg13g2_nor3_1 _1609_ (.A(_0850_),
    .B(_0851_),
    .C(_0852_),
    .Y(_0085_));
 sg13g2_nor2_1 _1610_ (.A(net145),
    .B(net497),
    .Y(_0853_));
 sg13g2_nor2_1 _1611_ (.A(net139),
    .B(net522),
    .Y(_0854_));
 sg13g2_nor2_1 _1612_ (.A(net208),
    .B(net557),
    .Y(_0855_));
 sg13g2_nor3_1 _1613_ (.A(_0853_),
    .B(_0854_),
    .C(_0855_),
    .Y(_0086_));
 sg13g2_nor2_1 _1614_ (.A(net145),
    .B(net525),
    .Y(_0856_));
 sg13g2_a221oi_1 _1615_ (.B2(_0489_),
    .C1(_0856_),
    .B1(net514),
    .A1(_0490_),
    .Y(_0087_),
    .A2(net571));
 sg13g2_nor2_1 _1616_ (.A(\bitserial_cipher.key[30] ),
    .B(net497),
    .Y(_0857_));
 sg13g2_nor2_1 _1617_ (.A(net219),
    .B(net556),
    .Y(_0858_));
 sg13g2_nor2_1 _1618_ (.A(\bitserial_cipher.key[29] ),
    .B(net525),
    .Y(_0859_));
 sg13g2_nor3_1 _1619_ (.A(_0857_),
    .B(_0858_),
    .C(_0859_),
    .Y(_0088_));
 sg13g2_nor2_1 _1620_ (.A(\bitserial_cipher.key[31] ),
    .B(net496),
    .Y(_0860_));
 sg13g2_nor2_1 _1621_ (.A(\bitserial_cipher.key[30] ),
    .B(net522),
    .Y(_0861_));
 sg13g2_nor2_1 _1622_ (.A(net139),
    .B(net556),
    .Y(_0862_));
 sg13g2_nor3_1 _1623_ (.A(_0860_),
    .B(_0861_),
    .C(_0862_),
    .Y(_0089_));
 sg13g2_nor2_1 _1624_ (.A(net123),
    .B(net496),
    .Y(_0863_));
 sg13g2_nor2_1 _1625_ (.A(net214),
    .B(net522),
    .Y(_0864_));
 sg13g2_nor2_1 _1626_ (.A(net145),
    .B(net556),
    .Y(_0865_));
 sg13g2_nor3_1 _1627_ (.A(_0863_),
    .B(_0864_),
    .C(_0865_),
    .Y(_0090_));
 sg13g2_nor2_1 _1628_ (.A(net123),
    .B(net522),
    .Y(_0866_));
 sg13g2_a221oi_1 _1629_ (.B2(_0488_),
    .C1(_0866_),
    .B1(net514),
    .A1(_0489_),
    .Y(_0091_),
    .A2(net571));
 sg13g2_nor2_1 _1630_ (.A(\bitserial_cipher.key[34] ),
    .B(net496),
    .Y(_0867_));
 sg13g2_nor2_1 _1631_ (.A(\bitserial_cipher.key[30] ),
    .B(net557),
    .Y(_0868_));
 sg13g2_nor2_1 _1632_ (.A(net93),
    .B(net522),
    .Y(_0869_));
 sg13g2_nor3_1 _1633_ (.A(_0867_),
    .B(_0868_),
    .C(_0869_),
    .Y(_0092_));
 sg13g2_nor2_1 _1634_ (.A(net73),
    .B(net496),
    .Y(_0870_));
 sg13g2_nor2_1 _1635_ (.A(net255),
    .B(net520),
    .Y(_0871_));
 sg13g2_nor2_1 _1636_ (.A(net214),
    .B(net555),
    .Y(_0872_));
 sg13g2_nor3_1 _1637_ (.A(_0870_),
    .B(_0871_),
    .C(_0872_),
    .Y(_0093_));
 sg13g2_nor2_1 _1638_ (.A(\bitserial_cipher.key[36] ),
    .B(net496),
    .Y(_0873_));
 sg13g2_nor2_1 _1639_ (.A(\bitserial_cipher.key[32] ),
    .B(net555),
    .Y(_0874_));
 sg13g2_nor2_1 _1640_ (.A(net73),
    .B(net520),
    .Y(_0875_));
 sg13g2_nor3_1 _1641_ (.A(_0873_),
    .B(_0874_),
    .C(_0875_),
    .Y(_0094_));
 sg13g2_nor2_1 _1642_ (.A(net207),
    .B(net520),
    .Y(_0876_));
 sg13g2_a221oi_1 _1643_ (.B2(_0487_),
    .C1(_0876_),
    .B1(net514),
    .A1(_0488_),
    .Y(_0095_),
    .A2(net571));
 sg13g2_nor2_1 _1644_ (.A(net166),
    .B(net496),
    .Y(_0877_));
 sg13g2_nor2_1 _1645_ (.A(net255),
    .B(net555),
    .Y(_0878_));
 sg13g2_nor2_1 _1646_ (.A(net172),
    .B(net520),
    .Y(_0879_));
 sg13g2_nor3_1 _1647_ (.A(_0877_),
    .B(_0878_),
    .C(_0879_),
    .Y(_0096_));
 sg13g2_nor2_1 _1648_ (.A(net49),
    .B(net496),
    .Y(_0880_));
 sg13g2_nor2_1 _1649_ (.A(net166),
    .B(net520),
    .Y(_0881_));
 sg13g2_nor2_1 _1650_ (.A(net73),
    .B(net555),
    .Y(_0882_));
 sg13g2_nor3_1 _1651_ (.A(_0880_),
    .B(_0881_),
    .C(_0882_),
    .Y(_0097_));
 sg13g2_nor2_1 _1652_ (.A(\bitserial_cipher.key[40] ),
    .B(net496),
    .Y(_0883_));
 sg13g2_nor2_1 _1653_ (.A(net49),
    .B(net520),
    .Y(_0884_));
 sg13g2_nor2_1 _1654_ (.A(\bitserial_cipher.key[36] ),
    .B(net555),
    .Y(_0885_));
 sg13g2_nor3_1 _1655_ (.A(_0883_),
    .B(_0884_),
    .C(_0885_),
    .Y(_0098_));
 sg13g2_nor2_1 _1656_ (.A(\bitserial_cipher.key[40] ),
    .B(net520),
    .Y(_0886_));
 sg13g2_a221oi_1 _1657_ (.B2(_0486_),
    .C1(_0886_),
    .B1(net514),
    .A1(_0487_),
    .Y(_0099_),
    .A2(net571));
 sg13g2_nor2_1 _1658_ (.A(net99),
    .B(net497),
    .Y(_0887_));
 sg13g2_nor2_1 _1659_ (.A(net121),
    .B(net521),
    .Y(_0888_));
 sg13g2_nor2_1 _1660_ (.A(\bitserial_cipher.key[38] ),
    .B(net555),
    .Y(_0889_));
 sg13g2_nor3_1 _1661_ (.A(_0887_),
    .B(_0888_),
    .C(_0889_),
    .Y(_0100_));
 sg13g2_nor2_1 _1662_ (.A(\bitserial_cipher.key[43] ),
    .B(net497),
    .Y(_0890_));
 sg13g2_nor2_1 _1663_ (.A(net99),
    .B(net521),
    .Y(_0891_));
 sg13g2_nor2_1 _1664_ (.A(net49),
    .B(net555),
    .Y(_0892_));
 sg13g2_nor3_1 _1665_ (.A(_0890_),
    .B(_0891_),
    .C(_0892_),
    .Y(_0101_));
 sg13g2_nor2_1 _1666_ (.A(net152),
    .B(net497),
    .Y(_0893_));
 sg13g2_nor2_1 _1667_ (.A(net237),
    .B(net555),
    .Y(_0894_));
 sg13g2_nor2_1 _1668_ (.A(\bitserial_cipher.key[43] ),
    .B(net520),
    .Y(_0895_));
 sg13g2_nor3_1 _1669_ (.A(_0893_),
    .B(_0894_),
    .C(_0895_),
    .Y(_0102_));
 sg13g2_nor2_1 _1670_ (.A(net152),
    .B(net521),
    .Y(_0896_));
 sg13g2_a221oi_1 _1671_ (.B2(_0485_),
    .C1(_0896_),
    .B1(net514),
    .A1(_0486_),
    .Y(_0103_),
    .A2(net571));
 sg13g2_nor2_1 _1672_ (.A(\bitserial_cipher.key[46] ),
    .B(net497),
    .Y(_0897_));
 sg13g2_nor2_1 _1673_ (.A(\bitserial_cipher.key[42] ),
    .B(net556),
    .Y(_0898_));
 sg13g2_nor2_1 _1674_ (.A(net67),
    .B(net521),
    .Y(_0899_));
 sg13g2_nor3_1 _1675_ (.A(_0897_),
    .B(_0898_),
    .C(_0899_),
    .Y(_0104_));
 sg13g2_nor2_1 _1676_ (.A(\bitserial_cipher.key[47] ),
    .B(net500),
    .Y(_0900_));
 sg13g2_nor2_1 _1677_ (.A(\bitserial_cipher.key[43] ),
    .B(net556),
    .Y(_0901_));
 sg13g2_nor2_1 _1678_ (.A(net175),
    .B(net521),
    .Y(_0902_));
 sg13g2_nor3_1 _1679_ (.A(_0900_),
    .B(_0901_),
    .C(_0902_),
    .Y(_0105_));
 sg13g2_nor2_1 _1680_ (.A(\bitserial_cipher.key[48] ),
    .B(net500),
    .Y(_0903_));
 sg13g2_nor2_1 _1681_ (.A(\bitserial_cipher.key[47] ),
    .B(net523),
    .Y(_0904_));
 sg13g2_nor2_1 _1682_ (.A(net152),
    .B(net556),
    .Y(_0905_));
 sg13g2_nor3_1 _1683_ (.A(_0903_),
    .B(_0904_),
    .C(_0905_),
    .Y(_0106_));
 sg13g2_nor2_1 _1684_ (.A(net187),
    .B(net523),
    .Y(_0211_));
 sg13g2_a221oi_1 _1685_ (.B2(_0484_),
    .C1(_0211_),
    .B1(net514),
    .A1(_0485_),
    .Y(_0107_),
    .A2(net571));
 sg13g2_nor2_1 _1686_ (.A(\bitserial_cipher.key[50] ),
    .B(net500),
    .Y(_0212_));
 sg13g2_nor2_1 _1687_ (.A(\bitserial_cipher.key[46] ),
    .B(net558),
    .Y(_0213_));
 sg13g2_nor2_1 _1688_ (.A(net128),
    .B(net523),
    .Y(_0214_));
 sg13g2_nor3_1 _1689_ (.A(_0212_),
    .B(_0213_),
    .C(_0214_),
    .Y(_0108_));
 sg13g2_nor2_1 _1690_ (.A(net188),
    .B(net500),
    .Y(_0215_));
 sg13g2_nor2_1 _1691_ (.A(\bitserial_cipher.key[50] ),
    .B(net523),
    .Y(_0216_));
 sg13g2_nor2_1 _1692_ (.A(net251),
    .B(net558),
    .Y(_0217_));
 sg13g2_nor3_1 _1693_ (.A(_0215_),
    .B(_0216_),
    .C(_0217_),
    .Y(_0109_));
 sg13g2_nor2_1 _1694_ (.A(\bitserial_cipher.key[52] ),
    .B(net500),
    .Y(_0218_));
 sg13g2_nor2_1 _1695_ (.A(net188),
    .B(net523),
    .Y(_0219_));
 sg13g2_nor2_1 _1696_ (.A(net187),
    .B(net558),
    .Y(_0220_));
 sg13g2_nor3_1 _1697_ (.A(_0218_),
    .B(_0219_),
    .C(_0220_),
    .Y(_0110_));
 sg13g2_nor2_1 _1698_ (.A(net213),
    .B(net523),
    .Y(_0221_));
 sg13g2_a221oi_1 _1699_ (.B2(_0483_),
    .C1(_0221_),
    .B1(net515),
    .A1(_0484_),
    .Y(_0111_),
    .A2(net572));
 sg13g2_nor2_1 _1700_ (.A(\bitserial_cipher.key[54] ),
    .B(net501),
    .Y(_0222_));
 sg13g2_nor2_1 _1701_ (.A(\bitserial_cipher.key[50] ),
    .B(net558),
    .Y(_0223_));
 sg13g2_nor2_1 _1702_ (.A(net126),
    .B(net524),
    .Y(_0224_));
 sg13g2_nor3_1 _1703_ (.A(_0222_),
    .B(_0223_),
    .C(_0224_),
    .Y(_0112_));
 sg13g2_nor2_1 _1704_ (.A(\bitserial_cipher.key[55] ),
    .B(net500),
    .Y(_0225_));
 sg13g2_nor2_1 _1705_ (.A(\bitserial_cipher.key[51] ),
    .B(net558),
    .Y(_0226_));
 sg13g2_nor2_1 _1706_ (.A(net183),
    .B(net523),
    .Y(_0227_));
 sg13g2_nor3_1 _1707_ (.A(_0225_),
    .B(_0226_),
    .C(_0227_),
    .Y(_0113_));
 sg13g2_nor2_1 _1708_ (.A(net165),
    .B(net500),
    .Y(_0228_));
 sg13g2_nor2_1 _1709_ (.A(net217),
    .B(net524),
    .Y(_0229_));
 sg13g2_nor2_1 _1710_ (.A(net213),
    .B(net559),
    .Y(_0230_));
 sg13g2_nor3_1 _1711_ (.A(_0228_),
    .B(_0229_),
    .C(_0230_),
    .Y(_0114_));
 sg13g2_nor2_1 _1712_ (.A(net165),
    .B(net524),
    .Y(_0231_));
 sg13g2_a221oi_1 _1713_ (.B2(_0482_),
    .C1(_0231_),
    .B1(net515),
    .A1(_0483_),
    .Y(_0115_),
    .A2(net572));
 sg13g2_nor2_1 _1714_ (.A(\bitserial_cipher.key[58] ),
    .B(net501),
    .Y(_0232_));
 sg13g2_nor2_1 _1715_ (.A(net147),
    .B(net524),
    .Y(_0233_));
 sg13g2_nor2_1 _1716_ (.A(\bitserial_cipher.key[54] ),
    .B(net558),
    .Y(_0234_));
 sg13g2_nor3_1 _1717_ (.A(_0232_),
    .B(_0233_),
    .C(_0234_),
    .Y(_0116_));
 sg13g2_nor2_1 _1718_ (.A(net135),
    .B(net503),
    .Y(_0235_));
 sg13g2_nor2_1 _1719_ (.A(net253),
    .B(net524),
    .Y(_0236_));
 sg13g2_nor2_1 _1720_ (.A(net217),
    .B(net558),
    .Y(_0237_));
 sg13g2_nor3_1 _1721_ (.A(_0235_),
    .B(_0236_),
    .C(_0237_),
    .Y(_0117_));
 sg13g2_nor2_1 _1722_ (.A(\bitserial_cipher.key[60] ),
    .B(net503),
    .Y(_0238_));
 sg13g2_nor2_1 _1723_ (.A(net135),
    .B(net523),
    .Y(_0239_));
 sg13g2_nor2_1 _1724_ (.A(\bitserial_cipher.key[56] ),
    .B(net558),
    .Y(_0240_));
 sg13g2_nor3_1 _1725_ (.A(_0238_),
    .B(_0239_),
    .C(_0240_),
    .Y(_0118_));
 sg13g2_nor2_1 _1726_ (.A(net198),
    .B(net532),
    .Y(_0241_));
 sg13g2_a221oi_1 _1727_ (.B2(_0481_),
    .C1(_0241_),
    .B1(net516),
    .A1(_0482_),
    .Y(_0119_),
    .A2(net574));
 sg13g2_nor2_1 _1728_ (.A(\bitserial_cipher.key[62] ),
    .B(net503),
    .Y(_0242_));
 sg13g2_nor2_1 _1729_ (.A(\bitserial_cipher.key[58] ),
    .B(net563),
    .Y(_0243_));
 sg13g2_nor2_1 _1730_ (.A(net107),
    .B(net532),
    .Y(_0244_));
 sg13g2_nor3_1 _1731_ (.A(_0242_),
    .B(_0243_),
    .C(_0244_),
    .Y(_0120_));
 sg13g2_nor2_1 _1732_ (.A(net177),
    .B(net503),
    .Y(_0245_));
 sg13g2_nor2_1 _1733_ (.A(\bitserial_cipher.key[62] ),
    .B(net531),
    .Y(_0246_));
 sg13g2_nor2_1 _1734_ (.A(net135),
    .B(net563),
    .Y(_0247_));
 sg13g2_nor3_1 _1735_ (.A(_0245_),
    .B(_0246_),
    .C(_0247_),
    .Y(_0121_));
 sg13g2_nor2_1 _1736_ (.A(net212),
    .B(net503),
    .Y(_0248_));
 sg13g2_nor2_1 _1737_ (.A(net177),
    .B(net531),
    .Y(_0249_));
 sg13g2_nor2_1 _1738_ (.A(net198),
    .B(net563),
    .Y(_0250_));
 sg13g2_nor3_1 _1739_ (.A(_0248_),
    .B(_0249_),
    .C(_0250_),
    .Y(_0122_));
 sg13g2_nor2_1 _1740_ (.A(net212),
    .B(net532),
    .Y(_0251_));
 sg13g2_a221oi_1 _1741_ (.B2(_0480_),
    .C1(_0251_),
    .B1(net516),
    .A1(_0481_),
    .Y(_0123_),
    .A2(net574));
 sg13g2_nor2_1 _1742_ (.A(\bitserial_cipher.key[66] ),
    .B(net504),
    .Y(_0252_));
 sg13g2_nor2_1 _1743_ (.A(\bitserial_cipher.key[62] ),
    .B(net564),
    .Y(_0253_));
 sg13g2_nor2_1 _1744_ (.A(net69),
    .B(net532),
    .Y(_0254_));
 sg13g2_nor3_1 _1745_ (.A(_0252_),
    .B(_0253_),
    .C(_0254_),
    .Y(_0124_));
 sg13g2_nor2_1 _1746_ (.A(net199),
    .B(net504),
    .Y(_0255_));
 sg13g2_nor2_1 _1747_ (.A(net202),
    .B(net531),
    .Y(_0256_));
 sg13g2_nor2_1 _1748_ (.A(net177),
    .B(net563),
    .Y(_0257_));
 sg13g2_nor3_1 _1749_ (.A(_0255_),
    .B(_0256_),
    .C(_0257_),
    .Y(_0125_));
 sg13g2_nor2_1 _1750_ (.A(net120),
    .B(net504),
    .Y(_0258_));
 sg13g2_nor2_1 _1751_ (.A(\bitserial_cipher.key[64] ),
    .B(net563),
    .Y(_0259_));
 sg13g2_nor2_1 _1752_ (.A(net199),
    .B(net531),
    .Y(_0260_));
 sg13g2_nor3_1 _1753_ (.A(_0258_),
    .B(_0259_),
    .C(_0260_),
    .Y(_0126_));
 sg13g2_nor2_1 _1754_ (.A(net120),
    .B(net531),
    .Y(_0261_));
 sg13g2_a221oi_1 _1755_ (.B2(_0479_),
    .C1(_0261_),
    .B1(net516),
    .A1(_0480_),
    .Y(_0127_),
    .A2(net574));
 sg13g2_nor2_1 _1756_ (.A(\bitserial_cipher.key[70] ),
    .B(net503),
    .Y(_0262_));
 sg13g2_nor2_1 _1757_ (.A(\bitserial_cipher.key[66] ),
    .B(net564),
    .Y(_0263_));
 sg13g2_nor2_1 _1758_ (.A(net118),
    .B(net532),
    .Y(_0264_));
 sg13g2_nor3_1 _1759_ (.A(_0262_),
    .B(_0263_),
    .C(_0264_),
    .Y(_0128_));
 sg13g2_nor2_1 _1760_ (.A(net201),
    .B(net503),
    .Y(_0265_));
 sg13g2_nor2_1 _1761_ (.A(net223),
    .B(net531),
    .Y(_0266_));
 sg13g2_nor2_1 _1762_ (.A(net199),
    .B(net564),
    .Y(_0267_));
 sg13g2_nor3_1 _1763_ (.A(_0265_),
    .B(_0266_),
    .C(_0267_),
    .Y(_0129_));
 sg13g2_nor2_1 _1764_ (.A(net150),
    .B(net503),
    .Y(_0268_));
 sg13g2_nor2_1 _1765_ (.A(net201),
    .B(net531),
    .Y(_0269_));
 sg13g2_nor2_1 _1766_ (.A(net120),
    .B(net563),
    .Y(_0270_));
 sg13g2_nor3_1 _1767_ (.A(_0268_),
    .B(_0269_),
    .C(_0270_),
    .Y(_0130_));
 sg13g2_nor2_1 _1768_ (.A(net150),
    .B(net531),
    .Y(_0271_));
 sg13g2_a221oi_1 _1769_ (.B2(_0478_),
    .C1(_0271_),
    .B1(net517),
    .A1(_0479_),
    .Y(_0131_),
    .A2(net575));
 sg13g2_nor2_1 _1770_ (.A(\bitserial_cipher.key[74] ),
    .B(net506),
    .Y(_0272_));
 sg13g2_nor2_1 _1771_ (.A(net85),
    .B(net533),
    .Y(_0273_));
 sg13g2_nor2_1 _1772_ (.A(\bitserial_cipher.key[70] ),
    .B(net564),
    .Y(_0274_));
 sg13g2_nor3_1 _1773_ (.A(_0272_),
    .B(_0273_),
    .C(_0274_),
    .Y(_0132_));
 sg13g2_nor2_1 _1774_ (.A(net256),
    .B(net506),
    .Y(_0275_));
 sg13g2_nor2_1 _1775_ (.A(\bitserial_cipher.key[74] ),
    .B(net533),
    .Y(_0276_));
 sg13g2_nor2_1 _1776_ (.A(net201),
    .B(net563),
    .Y(_0277_));
 sg13g2_nor3_1 _1777_ (.A(_0275_),
    .B(_0276_),
    .C(_0277_),
    .Y(_0133_));
 sg13g2_nor2_1 _1778_ (.A(\bitserial_cipher.key[76] ),
    .B(net506),
    .Y(_0278_));
 sg13g2_nor2_1 _1779_ (.A(net150),
    .B(net563),
    .Y(_0279_));
 sg13g2_nor2_1 _1780_ (.A(\bitserial_cipher.key[75] ),
    .B(net533),
    .Y(_0280_));
 sg13g2_nor3_1 _1781_ (.A(_0278_),
    .B(_0279_),
    .C(_0280_),
    .Y(_0134_));
 sg13g2_nor2_1 _1782_ (.A(net226),
    .B(net533),
    .Y(_0281_));
 sg13g2_a221oi_1 _1783_ (.B2(_0477_),
    .C1(_0281_),
    .B1(net517),
    .A1(_0478_),
    .Y(_0135_),
    .A2(net575));
 sg13g2_nor2_1 _1784_ (.A(\bitserial_cipher.key[78] ),
    .B(net506),
    .Y(_0282_));
 sg13g2_nor2_1 _1785_ (.A(\bitserial_cipher.key[74] ),
    .B(net565),
    .Y(_0283_));
 sg13g2_nor2_1 _1786_ (.A(net101),
    .B(net533),
    .Y(_0284_));
 sg13g2_nor3_1 _1787_ (.A(_0282_),
    .B(_0283_),
    .C(_0284_),
    .Y(_0136_));
 sg13g2_nor2_1 _1788_ (.A(\bitserial_cipher.key[79] ),
    .B(net505),
    .Y(_0285_));
 sg13g2_nor2_1 _1789_ (.A(\bitserial_cipher.key[75] ),
    .B(net565),
    .Y(_0286_));
 sg13g2_nor2_1 _1790_ (.A(net205),
    .B(net535),
    .Y(_0287_));
 sg13g2_nor3_1 _1791_ (.A(_0285_),
    .B(_0286_),
    .C(_0287_),
    .Y(_0137_));
 sg13g2_nor2_1 _1792_ (.A(net242),
    .B(net505),
    .Y(_0288_));
 sg13g2_nor2_1 _1793_ (.A(net269),
    .B(net533),
    .Y(_0289_));
 sg13g2_nor2_1 _1794_ (.A(net226),
    .B(net565),
    .Y(_0290_));
 sg13g2_nor3_1 _1795_ (.A(_0288_),
    .B(_0289_),
    .C(_0290_),
    .Y(_0138_));
 sg13g2_nor2_1 _1796_ (.A(net242),
    .B(net533),
    .Y(_0291_));
 sg13g2_a221oi_1 _1797_ (.B2(_0476_),
    .C1(_0291_),
    .B1(net517),
    .A1(_0477_),
    .Y(_0139_),
    .A2(net575));
 sg13g2_nor2_1 _1798_ (.A(\bitserial_cipher.key[82] ),
    .B(net505),
    .Y(_0292_));
 sg13g2_nor2_1 _1799_ (.A(\bitserial_cipher.key[78] ),
    .B(net565),
    .Y(_0293_));
 sg13g2_nor2_1 _1800_ (.A(net55),
    .B(net533),
    .Y(_0294_));
 sg13g2_nor3_1 _1801_ (.A(_0292_),
    .B(_0293_),
    .C(_0294_),
    .Y(_0140_));
 sg13g2_nor2_1 _1802_ (.A(net270),
    .B(net505),
    .Y(_0295_));
 sg13g2_nor2_1 _1803_ (.A(\bitserial_cipher.key[82] ),
    .B(net535),
    .Y(_0296_));
 sg13g2_nor2_1 _1804_ (.A(net269),
    .B(net565),
    .Y(_0297_));
 sg13g2_nor3_1 _1805_ (.A(_0295_),
    .B(_0296_),
    .C(_0297_),
    .Y(_0141_));
 sg13g2_nor2_1 _1806_ (.A(net125),
    .B(net505),
    .Y(_0298_));
 sg13g2_nor2_1 _1807_ (.A(net270),
    .B(net535),
    .Y(_0299_));
 sg13g2_nor2_1 _1808_ (.A(net242),
    .B(net565),
    .Y(_0300_));
 sg13g2_nor3_1 _1809_ (.A(_0298_),
    .B(_0299_),
    .C(_0300_),
    .Y(_0142_));
 sg13g2_nor2_1 _1810_ (.A(net125),
    .B(net534),
    .Y(_0301_));
 sg13g2_a221oi_1 _1811_ (.B2(_0475_),
    .C1(_0301_),
    .B1(net517),
    .A1(_0476_),
    .Y(_0143_),
    .A2(net575));
 sg13g2_nor2_1 _1812_ (.A(\bitserial_cipher.key[86] ),
    .B(net505),
    .Y(_0302_));
 sg13g2_nor2_1 _1813_ (.A(\bitserial_cipher.key[82] ),
    .B(net565),
    .Y(_0303_));
 sg13g2_nor2_1 _1814_ (.A(net111),
    .B(net534),
    .Y(_0304_));
 sg13g2_nor3_1 _1815_ (.A(_0302_),
    .B(_0303_),
    .C(_0304_),
    .Y(_0144_));
 sg13g2_nor2_1 _1816_ (.A(\bitserial_cipher.key[87] ),
    .B(net505),
    .Y(_0305_));
 sg13g2_nor2_1 _1817_ (.A(\bitserial_cipher.key[83] ),
    .B(net565),
    .Y(_0306_));
 sg13g2_nor2_1 _1818_ (.A(net156),
    .B(net534),
    .Y(_0307_));
 sg13g2_nor3_1 _1819_ (.A(_0305_),
    .B(_0306_),
    .C(_0307_),
    .Y(_0145_));
 sg13g2_nor2_1 _1820_ (.A(net211),
    .B(net506),
    .Y(_0308_));
 sg13g2_nor2_1 _1821_ (.A(net248),
    .B(net534),
    .Y(_0309_));
 sg13g2_nor2_1 _1822_ (.A(net125),
    .B(net566),
    .Y(_0310_));
 sg13g2_nor3_1 _1823_ (.A(_0308_),
    .B(_0309_),
    .C(_0310_),
    .Y(_0146_));
 sg13g2_nor2_1 _1824_ (.A(net211),
    .B(net534),
    .Y(_0311_));
 sg13g2_a221oi_1 _1825_ (.B2(_0474_),
    .C1(_0311_),
    .B1(net517),
    .A1(_0475_),
    .Y(_0147_),
    .A2(net575));
 sg13g2_nor2_1 _1826_ (.A(\bitserial_cipher.key[90] ),
    .B(net506),
    .Y(_0312_));
 sg13g2_nor2_1 _1827_ (.A(net170),
    .B(net534),
    .Y(_0313_));
 sg13g2_nor2_1 _1828_ (.A(net156),
    .B(net566),
    .Y(_0314_));
 sg13g2_nor3_1 _1829_ (.A(_0312_),
    .B(_0313_),
    .C(_0314_),
    .Y(_0148_));
 sg13g2_nor2_1 _1830_ (.A(net179),
    .B(net506),
    .Y(_0315_));
 sg13g2_nor2_1 _1831_ (.A(net235),
    .B(net534),
    .Y(_0316_));
 sg13g2_nor2_1 _1832_ (.A(\bitserial_cipher.key[87] ),
    .B(net566),
    .Y(_0317_));
 sg13g2_nor3_1 _1833_ (.A(_0315_),
    .B(_0316_),
    .C(_0317_),
    .Y(_0149_));
 sg13g2_nor2_1 _1834_ (.A(net143),
    .B(net505),
    .Y(_0318_));
 sg13g2_nor2_1 _1835_ (.A(net179),
    .B(net534),
    .Y(_0319_));
 sg13g2_nor2_1 _1836_ (.A(net211),
    .B(net566),
    .Y(_0320_));
 sg13g2_nor3_1 _1837_ (.A(_0318_),
    .B(_0319_),
    .C(_0320_),
    .Y(_0150_));
 sg13g2_nor2_1 _1838_ (.A(net143),
    .B(net535),
    .Y(_0321_));
 sg13g2_a221oi_1 _1839_ (.B2(_0473_),
    .C1(_0321_),
    .B1(net517),
    .A1(_0474_),
    .Y(_0151_),
    .A2(net574));
 sg13g2_nor2_1 _1840_ (.A(\bitserial_cipher.key[94] ),
    .B(net507),
    .Y(_0322_));
 sg13g2_nor2_1 _1841_ (.A(\bitserial_cipher.key[90] ),
    .B(net566),
    .Y(_0323_));
 sg13g2_nor2_1 _1842_ (.A(net57),
    .B(net540),
    .Y(_0324_));
 sg13g2_nor3_1 _1843_ (.A(_0322_),
    .B(_0323_),
    .C(_0324_),
    .Y(_0152_));
 sg13g2_nor2_1 _1844_ (.A(\bitserial_cipher.key[95] ),
    .B(net507),
    .Y(_0325_));
 sg13g2_nor2_1 _1845_ (.A(\bitserial_cipher.key[94] ),
    .B(net540),
    .Y(_0326_));
 sg13g2_nor2_1 _1846_ (.A(net179),
    .B(net566),
    .Y(_0327_));
 sg13g2_nor3_1 _1847_ (.A(_0325_),
    .B(_0326_),
    .C(_0327_),
    .Y(_0153_));
 sg13g2_nor2_1 _1848_ (.A(net218),
    .B(net507),
    .Y(_0328_));
 sg13g2_nor2_1 _1849_ (.A(net193),
    .B(net540),
    .Y(_0329_));
 sg13g2_nor2_1 _1850_ (.A(net143),
    .B(net566),
    .Y(_0330_));
 sg13g2_nor3_1 _1851_ (.A(_0328_),
    .B(_0329_),
    .C(_0330_),
    .Y(_0154_));
 sg13g2_nor2_1 _1852_ (.A(net218),
    .B(net540),
    .Y(_0331_));
 sg13g2_a221oi_1 _1853_ (.B2(_0472_),
    .C1(_0331_),
    .B1(net517),
    .A1(_0473_),
    .Y(_0155_),
    .A2(net575));
 sg13g2_nor2_1 _1854_ (.A(\bitserial_cipher.key[98] ),
    .B(net507),
    .Y(_0332_));
 sg13g2_nor2_1 _1855_ (.A(\bitserial_cipher.key[94] ),
    .B(net568),
    .Y(_0333_));
 sg13g2_nor2_1 _1856_ (.A(net91),
    .B(net540),
    .Y(_0334_));
 sg13g2_nor3_1 _1857_ (.A(_0332_),
    .B(_0333_),
    .C(_0334_),
    .Y(_0156_));
 sg13g2_nor2_1 _1858_ (.A(\bitserial_cipher.key[99] ),
    .B(net509),
    .Y(_0335_));
 sg13g2_nor2_1 _1859_ (.A(\bitserial_cipher.key[98] ),
    .B(net540),
    .Y(_0336_));
 sg13g2_nor2_1 _1860_ (.A(net193),
    .B(net567),
    .Y(_0337_));
 sg13g2_nor3_1 _1861_ (.A(_0335_),
    .B(_0336_),
    .C(_0337_),
    .Y(_0157_));
 sg13g2_nor2_1 _1862_ (.A(net231),
    .B(net507),
    .Y(_0338_));
 sg13g2_nor2_1 _1863_ (.A(net218),
    .B(net567),
    .Y(_0339_));
 sg13g2_nor2_1 _1864_ (.A(net247),
    .B(net539),
    .Y(_0340_));
 sg13g2_nor3_1 _1865_ (.A(_0338_),
    .B(_0339_),
    .C(_0340_),
    .Y(_0158_));
 sg13g2_nor2_1 _1866_ (.A(net231),
    .B(net539),
    .Y(_0341_));
 sg13g2_a221oi_1 _1867_ (.B2(_0470_),
    .C1(_0341_),
    .B1(net518),
    .A1(_0472_),
    .Y(_0159_),
    .A2(net577));
 sg13g2_nor2_1 _1868_ (.A(\bitserial_cipher.key[102] ),
    .B(net509),
    .Y(_0342_));
 sg13g2_nor2_1 _1869_ (.A(\bitserial_cipher.key[98] ),
    .B(net567),
    .Y(_0343_));
 sg13g2_nor2_1 _1870_ (.A(net71),
    .B(net538),
    .Y(_0344_));
 sg13g2_nor3_1 _1871_ (.A(_0342_),
    .B(_0343_),
    .C(_0344_),
    .Y(_0160_));
 sg13g2_nor2_1 _1872_ (.A(net259),
    .B(net507),
    .Y(_0345_));
 sg13g2_nor2_1 _1873_ (.A(net279),
    .B(net539),
    .Y(_0346_));
 sg13g2_nor2_1 _1874_ (.A(net247),
    .B(net567),
    .Y(_0347_));
 sg13g2_nor3_1 _1875_ (.A(_0345_),
    .B(_0346_),
    .C(_0347_),
    .Y(_0161_));
 sg13g2_nor2_1 _1876_ (.A(net234),
    .B(net507),
    .Y(_0348_));
 sg13g2_nor2_1 _1877_ (.A(net259),
    .B(net539),
    .Y(_0349_));
 sg13g2_nor2_1 _1878_ (.A(net231),
    .B(net567),
    .Y(_0350_));
 sg13g2_nor3_1 _1879_ (.A(_0348_),
    .B(_0349_),
    .C(_0350_),
    .Y(_0162_));
 sg13g2_nor2_1 _1880_ (.A(net234),
    .B(net539),
    .Y(_0351_));
 sg13g2_a221oi_1 _1881_ (.B2(_0471_),
    .C1(_0351_),
    .B1(net518),
    .A1(_0470_),
    .Y(_0163_),
    .A2(net576));
 sg13g2_nor2_1 _1882_ (.A(\bitserial_cipher.key[106] ),
    .B(net509),
    .Y(_0352_));
 sg13g2_nor2_1 _1883_ (.A(net63),
    .B(net539),
    .Y(_0353_));
 sg13g2_nor2_1 _1884_ (.A(\bitserial_cipher.key[102] ),
    .B(net568),
    .Y(_0354_));
 sg13g2_nor3_1 _1885_ (.A(_0352_),
    .B(_0353_),
    .C(_0354_),
    .Y(_0164_));
 sg13g2_nor2_1 _1886_ (.A(\bitserial_cipher.key[107] ),
    .B(net507),
    .Y(_0355_));
 sg13g2_nor2_1 _1887_ (.A(\bitserial_cipher.key[106] ),
    .B(net539),
    .Y(_0356_));
 sg13g2_nor2_1 _1888_ (.A(net259),
    .B(net568),
    .Y(_0357_));
 sg13g2_nor3_1 _1889_ (.A(_0355_),
    .B(_0356_),
    .C(_0357_),
    .Y(_0165_));
 sg13g2_nor2_1 _1890_ (.A(net185),
    .B(net508),
    .Y(_0358_));
 sg13g2_nor2_1 _1891_ (.A(net272),
    .B(net538),
    .Y(_0359_));
 sg13g2_nor2_1 _1892_ (.A(net234),
    .B(net568),
    .Y(_0360_));
 sg13g2_nor3_1 _1893_ (.A(_0358_),
    .B(_0359_),
    .C(_0360_),
    .Y(_0166_));
 sg13g2_nor2_1 _1894_ (.A(net185),
    .B(net538),
    .Y(_0361_));
 sg13g2_a221oi_1 _1895_ (.B2(_0459_),
    .C1(_0361_),
    .B1(net518),
    .A1(_0471_),
    .Y(_0167_),
    .A2(net577));
 sg13g2_nor2_1 _1896_ (.A(\bitserial_cipher.key[110] ),
    .B(net508),
    .Y(_0362_));
 sg13g2_nor2_1 _1897_ (.A(\bitserial_cipher.key[106] ),
    .B(net568),
    .Y(_0363_));
 sg13g2_nor2_1 _1898_ (.A(net89),
    .B(net538),
    .Y(_0364_));
 sg13g2_nor3_1 _1899_ (.A(_0362_),
    .B(_0363_),
    .C(_0364_),
    .Y(_0168_));
 sg13g2_nor2_1 _1900_ (.A(\bitserial_cipher.key[111] ),
    .B(net508),
    .Y(_0365_));
 sg13g2_nor2_1 _1901_ (.A(\bitserial_cipher.key[107] ),
    .B(net568),
    .Y(_0366_));
 sg13g2_nor2_1 _1902_ (.A(net167),
    .B(net538),
    .Y(_0367_));
 sg13g2_nor3_1 _1903_ (.A(_0365_),
    .B(_0366_),
    .C(_0367_),
    .Y(_0169_));
 sg13g2_nor2_1 _1904_ (.A(net137),
    .B(net508),
    .Y(_0368_));
 sg13g2_nor2_1 _1905_ (.A(net185),
    .B(net568),
    .Y(_0369_));
 sg13g2_nor2_1 _1906_ (.A(\bitserial_cipher.key[111] ),
    .B(net538),
    .Y(_0370_));
 sg13g2_nor3_1 _1907_ (.A(_0368_),
    .B(_0369_),
    .C(_0370_),
    .Y(_0170_));
 sg13g2_nor2_1 _1908_ (.A(net137),
    .B(net538),
    .Y(_0371_));
 sg13g2_a221oi_1 _1909_ (.B2(_0460_),
    .C1(_0371_),
    .B1(net517),
    .A1(_0459_),
    .Y(_0171_),
    .A2(net577));
 sg13g2_nor2_1 _1910_ (.A(net154),
    .B(net508),
    .Y(_0372_));
 sg13g2_nor2_1 _1911_ (.A(net169),
    .B(net538),
    .Y(_0373_));
 sg13g2_nor2_1 _1912_ (.A(net167),
    .B(net567),
    .Y(_0374_));
 sg13g2_nor3_1 _1913_ (.A(_0372_),
    .B(_0373_),
    .C(_0374_),
    .Y(_0172_));
 sg13g2_nor2_1 _1914_ (.A(\bitserial_cipher.key[115] ),
    .B(net508),
    .Y(_0375_));
 sg13g2_nor2_1 _1915_ (.A(\bitserial_cipher.key[111] ),
    .B(net567),
    .Y(_0376_));
 sg13g2_nor2_1 _1916_ (.A(net154),
    .B(net540),
    .Y(_0377_));
 sg13g2_nor3_1 _1917_ (.A(_0375_),
    .B(_0376_),
    .C(_0377_),
    .Y(_0173_));
 sg13g2_nor2_1 _1918_ (.A(net115),
    .B(net504),
    .Y(_0378_));
 sg13g2_nor2_1 _1919_ (.A(net227),
    .B(net536),
    .Y(_0379_));
 sg13g2_nor2_1 _1920_ (.A(net137),
    .B(net569),
    .Y(_0380_));
 sg13g2_nor3_1 _1921_ (.A(_0378_),
    .B(_0379_),
    .C(_0380_),
    .Y(_0174_));
 sg13g2_nor2_1 _1922_ (.A(net115),
    .B(net536),
    .Y(_0381_));
 sg13g2_a221oi_1 _1923_ (.B2(_0461_),
    .C1(_0381_),
    .B1(net518),
    .A1(_0460_),
    .Y(_0175_),
    .A2(net577));
 sg13g2_nor2_1 _1924_ (.A(\bitserial_cipher.key[118] ),
    .B(net508),
    .Y(_0382_));
 sg13g2_nor2_1 _1925_ (.A(\bitserial_cipher.key[114] ),
    .B(net567),
    .Y(_0383_));
 sg13g2_nor2_1 _1926_ (.A(net75),
    .B(net540),
    .Y(_0384_));
 sg13g2_nor3_1 _1927_ (.A(_0382_),
    .B(_0383_),
    .C(_0384_),
    .Y(_0176_));
 sg13g2_nor2_1 _1928_ (.A(net249),
    .B(net504),
    .Y(_0385_));
 sg13g2_nor2_1 _1929_ (.A(net227),
    .B(net564),
    .Y(_0386_));
 sg13g2_nor2_1 _1930_ (.A(\bitserial_cipher.key[118] ),
    .B(net536),
    .Y(_0387_));
 sg13g2_nor3_1 _1931_ (.A(_0385_),
    .B(_0386_),
    .C(_0387_),
    .Y(_0177_));
 sg13g2_nor2_1 _1932_ (.A(net190),
    .B(net504),
    .Y(_0388_));
 sg13g2_nor2_1 _1933_ (.A(net249),
    .B(net537),
    .Y(_0389_));
 sg13g2_nor2_1 _1934_ (.A(net115),
    .B(net569),
    .Y(_0390_));
 sg13g2_nor3_1 _1935_ (.A(_0388_),
    .B(_0389_),
    .C(_0390_),
    .Y(_0178_));
 sg13g2_nor2_1 _1936_ (.A(net190),
    .B(net537),
    .Y(_0391_));
 sg13g2_a221oi_1 _1937_ (.B2(_0462_),
    .C1(_0391_),
    .B1(net519),
    .A1(_0461_),
    .Y(_0179_),
    .A2(net576));
 sg13g2_nor2_1 _1938_ (.A(\bitserial_cipher.key[122] ),
    .B(net510),
    .Y(_0392_));
 sg13g2_nor2_1 _1939_ (.A(net181),
    .B(net537),
    .Y(_0393_));
 sg13g2_nor2_1 _1940_ (.A(\bitserial_cipher.key[118] ),
    .B(net564),
    .Y(_0394_));
 sg13g2_nor3_1 _1941_ (.A(_0392_),
    .B(_0393_),
    .C(_0394_),
    .Y(_0180_));
 sg13g2_nand2b_1 _1942_ (.Y(_0395_),
    .B(net574),
    .A_N(\bitserial_cipher.key[119] ));
 sg13g2_o21ai_1 _1943_ (.B1(_0395_),
    .Y(_0396_),
    .A1(\bitserial_cipher.key[122] ),
    .A2(net574));
 sg13g2_nand2_1 _1944_ (.Y(_0397_),
    .A(net97),
    .B(net516));
 sg13g2_o21ai_1 _1945_ (.B1(_0397_),
    .Y(_0181_),
    .A1(net516),
    .A2(_0396_));
 sg13g2_nor2_1 _1946_ (.A(net288),
    .B(net504),
    .Y(_0398_));
 sg13g2_nor2_1 _1947_ (.A(net97),
    .B(net536),
    .Y(_0399_));
 sg13g2_nor2_1 _1948_ (.A(net190),
    .B(net569),
    .Y(_0400_));
 sg13g2_nor3_1 _1949_ (.A(_0398_),
    .B(_0399_),
    .C(_0400_),
    .Y(_0182_));
 sg13g2_nor3_1 _1950_ (.A(\bitserial_cipher.key[124] ),
    .B(net576),
    .C(net537),
    .Y(_0401_));
 sg13g2_a221oi_1 _1951_ (.B2(_0497_),
    .C1(_0401_),
    .B1(net516),
    .A1(_0462_),
    .Y(_0183_),
    .A2(net576));
 sg13g2_a22oi_1 _1952_ (.Y(_0402_),
    .B1(net516),
    .B2(net276),
    .A2(net574),
    .A1(net306));
 sg13g2_o21ai_1 _1953_ (.B1(_0402_),
    .Y(_0184_),
    .A1(_0497_),
    .A2(net536));
 sg13g2_nand2_1 _1954_ (.Y(_0403_),
    .A(net97),
    .B(net576));
 sg13g2_a21oi_1 _1955_ (.A1(\bitserial_cipher.key[126] ),
    .A2(net569),
    .Y(_0404_),
    .B1(net516));
 sg13g2_a22oi_1 _1956_ (.Y(_0185_),
    .B1(_0403_),
    .B2(_0404_),
    .A2(net515),
    .A1(_0498_));
 sg13g2_o21ai_1 _1957_ (.B1(net343),
    .Y(_0405_),
    .A1(\bitserial_cipher.done ),
    .A2(_0534_));
 sg13g2_o21ai_1 _1958_ (.B1(_0405_),
    .Y(_0406_),
    .A1(net343),
    .A2(_0534_));
 sg13g2_inv_1 _1959_ (.Y(_0186_),
    .A(_0406_));
 sg13g2_nor2b_1 _1960_ (.A(net239),
    .B_N(_0405_),
    .Y(_0407_));
 sg13g2_a21oi_1 _1961_ (.A1(_0511_),
    .A2(_0535_),
    .Y(_0408_),
    .B1(_0543_));
 sg13g2_nor3_1 _1962_ (.A(\bitserial_cipher.done ),
    .B(net240),
    .C(_0408_),
    .Y(_0187_));
 sg13g2_nor2_1 _1963_ (.A(net318),
    .B(_0408_),
    .Y(_0409_));
 sg13g2_nand4_1 _1964_ (.B(\bitserial_cipher.rcount[1] ),
    .C(\bitserial_cipher.rcount[2] ),
    .A(\bitserial_cipher.rcount[0] ),
    .Y(_0410_),
    .D(_0534_));
 sg13g2_nand2_1 _1965_ (.Y(_0411_),
    .A(net616),
    .B(_0410_));
 sg13g2_nor3_1 _1966_ (.A(_0544_),
    .B(net319),
    .C(_0411_),
    .Y(_0188_));
 sg13g2_nand3_1 _1967_ (.B(net616),
    .C(_0410_),
    .A(net61),
    .Y(_0412_));
 sg13g2_o21ai_1 _1968_ (.B1(_0412_),
    .Y(_0189_),
    .A1(net61),
    .A2(_0410_));
 sg13g2_and3_1 _1969_ (.X(_0413_),
    .A(_0467_),
    .B(net579),
    .C(net587));
 sg13g2_a221oi_1 _1970_ (.B2(_0463_),
    .C1(_0413_),
    .B1(net547),
    .A1(_0466_),
    .Y(_0190_),
    .A2(net584));
 sg13g2_a22oi_1 _1971_ (.Y(_0414_),
    .B1(net584),
    .B2(\bitserial_cipher.state[33] ),
    .A2(net579),
    .A1(\bitserial_cipher.state[36] ));
 sg13g2_o21ai_1 _1972_ (.B1(_0414_),
    .Y(_0191_),
    .A1(_0464_),
    .A2(_0655_));
 sg13g2_a22oi_1 _1973_ (.Y(_0415_),
    .B1(net546),
    .B2(net197),
    .A2(net579),
    .A1(net130));
 sg13g2_o21ai_1 _1974_ (.B1(_0415_),
    .Y(_0192_),
    .A1(_0469_),
    .A2(net587));
 sg13g2_a22oi_1 _1975_ (.Y(_0416_),
    .B1(net546),
    .B2(\bitserial_cipher.state[39] ),
    .A2(net579),
    .A1(\bitserial_cipher.state[38] ));
 sg13g2_o21ai_1 _1976_ (.B1(_0416_),
    .Y(_0193_),
    .A1(_0467_),
    .A2(net587));
 sg13g2_a22oi_1 _1977_ (.Y(_0417_),
    .B1(net546),
    .B2(\bitserial_cipher.state[40] ),
    .A2(net579),
    .A1(\bitserial_cipher.state[39] ));
 sg13g2_o21ai_1 _1978_ (.B1(_0417_),
    .Y(_0194_),
    .A1(_0463_),
    .A2(net587));
 sg13g2_a22oi_1 _1979_ (.Y(_0418_),
    .B1(net584),
    .B2(net130),
    .A2(net581),
    .A1(\bitserial_cipher.state[40] ));
 sg13g2_o21ai_1 _1980_ (.B1(_0418_),
    .Y(_0195_),
    .A1(_0465_),
    .A2(_0655_));
 sg13g2_nand2_1 _1981_ (.Y(_0419_),
    .A(net79),
    .B(net547));
 sg13g2_nand2_1 _1982_ (.Y(_0420_),
    .A(net197),
    .B(net584));
 sg13g2_nand3_1 _1983_ (.B(net579),
    .C(net588),
    .A(net224),
    .Y(_0421_));
 sg13g2_nand3_1 _1984_ (.B(_0420_),
    .C(_0421_),
    .A(_0419_),
    .Y(_0196_));
 sg13g2_nand3_1 _1985_ (.B(net579),
    .C(net588),
    .A(net79),
    .Y(_0422_));
 sg13g2_a22oi_1 _1986_ (.Y(_0423_),
    .B1(net547),
    .B2(\bitserial_cipher.state[43] ),
    .A2(net585),
    .A1(\bitserial_cipher.state[39] ));
 sg13g2_nand2_1 _1987_ (.Y(_0197_),
    .A(_0422_),
    .B(_0423_));
 sg13g2_nand2_1 _1988_ (.Y(_0424_),
    .A(net291),
    .B(net587));
 sg13g2_nand2_1 _1989_ (.Y(_0425_),
    .A(net36),
    .B(net587));
 sg13g2_a221oi_1 _1990_ (.B2(\bitserial_cipher.state[44] ),
    .C1(net547),
    .B1(_0565_),
    .A1(\bitserial_cipher.state[28] ),
    .Y(_0426_),
    .A2(net599));
 sg13g2_a22oi_1 _1991_ (.Y(_0198_),
    .B1(_0424_),
    .B2(_0426_),
    .A2(net546),
    .A1(_0466_));
 sg13g2_a221oi_1 _1992_ (.B2(\bitserial_cipher.state[45] ),
    .C1(net547),
    .B1(_0565_),
    .A1(\bitserial_cipher.state[29] ),
    .Y(_0427_),
    .A2(net599));
 sg13g2_a22oi_1 _1993_ (.Y(_0199_),
    .B1(_0425_),
    .B2(_0427_),
    .A2(net546),
    .A1(_0468_));
 sg13g2_a22oi_1 _1994_ (.Y(_0428_),
    .B1(_0565_),
    .B2(\bitserial_cipher.state[46] ),
    .A2(net599),
    .A1(\bitserial_cipher.state[30] ));
 sg13g2_nand2_1 _1995_ (.Y(_0429_),
    .A(net105),
    .B(net587));
 sg13g2_a21oi_1 _1996_ (.A1(net289),
    .A2(net587),
    .Y(_0430_),
    .B1(net546));
 sg13g2_a22oi_1 _1997_ (.Y(_0200_),
    .B1(_0428_),
    .B2(_0430_),
    .A2(net546),
    .A1(_0469_));
 sg13g2_a221oi_1 _1998_ (.B2(\bitserial_cipher.state[47] ),
    .C1(net547),
    .B1(_0565_),
    .A1(\bitserial_cipher.state[31] ),
    .Y(_0431_),
    .A2(net599));
 sg13g2_a22oi_1 _1999_ (.Y(_0201_),
    .B1(_0429_),
    .B2(_0431_),
    .A2(net546),
    .A1(_0467_));
 sg13g2_nand2_1 _2000_ (.Y(_0432_),
    .A(net95),
    .B(net580));
 sg13g2_a22oi_1 _2001_ (.Y(_0433_),
    .B1(net554),
    .B2(net53),
    .A2(net593),
    .A1(\bitserial_cipher.state[48] ));
 sg13g2_nand2_1 _2002_ (.Y(_0202_),
    .A(_0432_),
    .B(_0433_));
 sg13g2_nand2_1 _2003_ (.Y(_0434_),
    .A(net53),
    .B(net580));
 sg13g2_a22oi_1 _2004_ (.Y(_0435_),
    .B1(net554),
    .B2(\bitserial_cipher.state[53] ),
    .A2(net593),
    .A1(\bitserial_cipher.state[49] ));
 sg13g2_nand2_1 _2005_ (.Y(_0203_),
    .A(_0434_),
    .B(_0435_));
 sg13g2_nand2_1 _2006_ (.Y(_0436_),
    .A(net51),
    .B(_0563_));
 sg13g2_a22oi_1 _2007_ (.Y(_0437_),
    .B1(net580),
    .B2(\bitserial_cipher.state[53] ),
    .A2(net593),
    .A1(\bitserial_cipher.state[50] ));
 sg13g2_nand2_1 _2008_ (.Y(_0204_),
    .A(_0436_),
    .B(_0437_));
 sg13g2_nand2_1 _2009_ (.Y(_0438_),
    .A(net51),
    .B(net581));
 sg13g2_a22oi_1 _2010_ (.Y(_0439_),
    .B1(_0563_),
    .B2(net87),
    .A2(net596),
    .A1(\bitserial_cipher.state[51] ));
 sg13g2_nand2_1 _2011_ (.Y(_0205_),
    .A(_0438_),
    .B(net88));
 sg13g2_nand2b_1 _2012_ (.Y(_0440_),
    .B(net554),
    .A_N(net47));
 sg13g2_o21ai_1 _2013_ (.B1(_0440_),
    .Y(_0441_),
    .A1(net53),
    .A2(net597));
 sg13g2_a21oi_1 _2014_ (.A1(_0458_),
    .A2(net580),
    .Y(_0206_),
    .B1(_0441_));
 sg13g2_nand2_1 _2015_ (.Y(_0442_),
    .A(net47),
    .B(net580));
 sg13g2_a22oi_1 _2016_ (.Y(_0443_),
    .B1(net554),
    .B2(net34),
    .A2(net595),
    .A1(\bitserial_cipher.state[53] ));
 sg13g2_nand2_1 _2017_ (.Y(_0207_),
    .A(_0442_),
    .B(_0443_));
 sg13g2_nand2_1 _2018_ (.Y(_0444_),
    .A(net34),
    .B(net580));
 sg13g2_a22oi_1 _2019_ (.Y(_0445_),
    .B1(net554),
    .B2(\bitserial_cipher.state[58] ),
    .A2(net595),
    .A1(\bitserial_cipher.state[54] ));
 sg13g2_nand2_1 _2020_ (.Y(_0208_),
    .A(_0444_),
    .B(_0445_));
 sg13g2_nand2_1 _2021_ (.Y(_0446_),
    .A(net81),
    .B(net580));
 sg13g2_a22oi_1 _2022_ (.Y(_0447_),
    .B1(net554),
    .B2(\bitserial_cipher.state[59] ),
    .A2(net595),
    .A1(\bitserial_cipher.state[55] ));
 sg13g2_nand2_1 _2023_ (.Y(_0209_),
    .A(_0446_),
    .B(_0447_));
 sg13g2_nand2_1 _2024_ (.Y(_0448_),
    .A(net341),
    .B(net582));
 sg13g2_a22oi_1 _2025_ (.Y(_0449_),
    .B1(net584),
    .B2(net351),
    .A2(net612),
    .A1(\bitserial_cipher.state[28] ));
 sg13g2_nand3_1 _2026_ (.B(_0448_),
    .C(_0449_),
    .A(net511),
    .Y(_0450_));
 sg13g2_o21ai_1 _2027_ (.B1(_0450_),
    .Y(_0451_),
    .A1(net345),
    .A2(net511));
 sg13g2_inv_1 _2028_ (.Y(_0210_),
    .A(_0451_));
 sg13g2_dfrbp_1 _2029_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net631),
    .D(_0001_),
    .Q_N(_1114_),
    .Q(\bitserial_cipher.state[45] ));
 sg13g2_dfrbp_1 _2030_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net634),
    .D(_0002_),
    .Q_N(_1113_),
    .Q(\bitserial_cipher.state[46] ));
 sg13g2_dfrbp_1 _2031_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net631),
    .D(_0003_),
    .Q_N(_1112_),
    .Q(\bitserial_cipher.state[47] ));
 sg13g2_dfrbp_1 _2032_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net634),
    .D(_0004_),
    .Q_N(_1111_),
    .Q(\bitserial_cipher.state[48] ));
 sg13g2_dfrbp_1 _2033_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net634),
    .D(net110),
    .Q_N(_1110_),
    .Q(\bitserial_cipher.state[49] ));
 sg13g2_dfrbp_1 _2034_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net634),
    .D(net229),
    .Q_N(_1109_),
    .Q(\bitserial_cipher.state[50] ));
 sg13g2_dfrbp_1 _2035_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net635),
    .D(_0007_),
    .Q_N(_1108_),
    .Q(\bitserial_cipher.state[51] ));
 sg13g2_dfrbp_1 _2036_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net632),
    .D(net350),
    .Q_N(_1107_),
    .Q(\bitserial_cipher.state[12] ));
 sg13g2_dfrbp_1 _2037_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net632),
    .D(_0009_),
    .Q_N(_1106_),
    .Q(\bitserial_cipher.state[13] ));
 sg13g2_dfrbp_1 _2038_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net632),
    .D(_0010_),
    .Q_N(_1105_),
    .Q(\bitserial_cipher.state[14] ));
 sg13g2_dfrbp_1 _2039_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net632),
    .D(_0011_),
    .Q_N(_1104_),
    .Q(\bitserial_cipher.state[15] ));
 sg13g2_dfrbp_1 _2040_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net632),
    .D(_0012_),
    .Q_N(_1103_),
    .Q(\bitserial_cipher.state[28] ));
 sg13g2_dfrbp_1 _2041_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net632),
    .D(net357),
    .Q_N(_1102_),
    .Q(\bitserial_cipher.state[29] ));
 sg13g2_dfrbp_1 _2042_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net628),
    .D(_0014_),
    .Q_N(_1101_),
    .Q(\bitserial_cipher.state[30] ));
 sg13g2_dfrbp_1 _2043_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net632),
    .D(_0015_),
    .Q_N(_1115_),
    .Q(\bitserial_cipher.state[31] ));
 sg13g2_dfrbp_1 _2044_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net654),
    .D(\bitserial_cipher.ctlstate_next[0] ),
    .Q_N(_1116_),
    .Q(\bitserial_cipher.ctlstate[0] ));
 sg13g2_dfrbp_1 _2045_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net653),
    .D(\bitserial_cipher.ctlstate_next[1] ),
    .Q_N(_1117_),
    .Q(\bitserial_cipher.ctlstate[1] ));
 sg13g2_dfrbp_1 _2046_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net654),
    .D(\bitserial_cipher.ctlstate_next[2] ),
    .Q_N(_1118_),
    .Q(\bitserial_cipher.ctlstate[2] ));
 sg13g2_dfrbp_1 _2047_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net654),
    .D(\bitserial_cipher.ctlstate_next[3] ),
    .Q_N(_1100_),
    .Q(\bitserial_cipher.ctlstate[3] ));
 sg13g2_dfrbp_1 _2048_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net649),
    .D(_0016_),
    .Q_N(\bitserial_cipher.rc[0] ),
    .Q(_0000_));
 sg13g2_dfrbp_1 _2049_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net649),
    .D(_0017_),
    .Q_N(_1099_),
    .Q(\bitserial_cipher.rc[1] ));
 sg13g2_dfrbp_1 _2050_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net649),
    .D(_0018_),
    .Q_N(_1098_),
    .Q(\bitserial_cipher.rc[2] ));
 sg13g2_dfrbp_1 _2051_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net649),
    .D(_0019_),
    .Q_N(_1097_),
    .Q(\bitserial_cipher.rc[3] ));
 sg13g2_dfrbp_1 _2052_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net648),
    .D(_0020_),
    .Q_N(_1096_),
    .Q(\bitserial_cipher.rc[4] ));
 sg13g2_dfrbp_1 _2053_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net649),
    .D(_0021_),
    .Q_N(_1095_),
    .Q(\bitserial_cipher.rc[5] ));
 sg13g2_dfrbp_1 _2054_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net648),
    .D(net278),
    .Q_N(_1094_),
    .Q(\bitserial_cipher.state[60] ));
 sg13g2_dfrbp_1 _2055_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net634),
    .D(net339),
    .Q_N(_1093_),
    .Q(\bitserial_cipher.state[61] ));
 sg13g2_dfrbp_1 _2056_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net648),
    .D(net309),
    .Q_N(_1092_),
    .Q(\bitserial_cipher.state[62] ));
 sg13g2_dfrbp_1 _2057_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net648),
    .D(_0025_),
    .Q_N(_1091_),
    .Q(\bitserial_cipher.dataq ));
 sg13g2_dfrbp_1 _2058_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net647),
    .D(net265),
    .Q_N(_1090_),
    .Q(\bitserial_cipher.state[4] ));
 sg13g2_dfrbp_1 _2059_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net647),
    .D(net317),
    .Q_N(_1089_),
    .Q(\bitserial_cipher.state[5] ));
 sg13g2_dfrbp_1 _2060_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net633),
    .D(net299),
    .Q_N(_1088_),
    .Q(\bitserial_cipher.state[6] ));
 sg13g2_dfrbp_1 _2061_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net633),
    .D(_0029_),
    .Q_N(_1087_),
    .Q(\bitserial_cipher.state[7] ));
 sg13g2_dfrbp_1 _2062_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net647),
    .D(net268),
    .Q_N(_1086_),
    .Q(\bitserial_cipher.state[8] ));
 sg13g2_dfrbp_1 _2063_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net647),
    .D(_0031_),
    .Q_N(_1085_),
    .Q(\bitserial_cipher.state[9] ));
 sg13g2_dfrbp_1 _2064_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net633),
    .D(net282),
    .Q_N(_1084_),
    .Q(\bitserial_cipher.state[10] ));
 sg13g2_dfrbp_1 _2065_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net632),
    .D(net312),
    .Q_N(_1083_),
    .Q(\bitserial_cipher.state[11] ));
 sg13g2_dfrbp_1 _2066_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net629),
    .D(net216),
    .Q_N(_1082_),
    .Q(\bitserial_cipher.state[20] ));
 sg13g2_dfrbp_1 _2067_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net629),
    .D(_0035_),
    .Q_N(_1081_),
    .Q(\bitserial_cipher.state[21] ));
 sg13g2_dfrbp_1 _2068_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net628),
    .D(_0036_),
    .Q_N(_1080_),
    .Q(\bitserial_cipher.state[22] ));
 sg13g2_dfrbp_1 _2069_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net629),
    .D(net287),
    .Q_N(_1079_),
    .Q(\bitserial_cipher.state[23] ));
 sg13g2_dfrbp_1 _2070_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net629),
    .D(_0038_),
    .Q_N(_1078_),
    .Q(\bitserial_cipher.state[24] ));
 sg13g2_dfrbp_1 _2071_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net628),
    .D(net294),
    .Q_N(_1077_),
    .Q(\bitserial_cipher.state[25] ));
 sg13g2_dfrbp_1 _2072_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net628),
    .D(net297),
    .Q_N(_1076_),
    .Q(\bitserial_cipher.state[26] ));
 sg13g2_dfrbp_1 _2073_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net628),
    .D(_0041_),
    .Q_N(_1075_),
    .Q(\bitserial_cipher.state[27] ));
 sg13g2_dfrbp_1 _2074_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net629),
    .D(net323),
    .Q_N(_1074_),
    .Q(\bitserial_cipher.state[16] ));
 sg13g2_dfrbp_1 _2075_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net628),
    .D(_0043_),
    .Q_N(_1073_),
    .Q(\bitserial_cipher.state[17] ));
 sg13g2_dfrbp_1 _2076_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net628),
    .D(net330),
    .Q_N(_1072_),
    .Q(\bitserial_cipher.state[18] ));
 sg13g2_dfrbp_1 _2077_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net628),
    .D(net275),
    .Q_N(_1071_),
    .Q(\bitserial_cipher.state[19] ));
 sg13g2_dfrbp_1 _2078_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net647),
    .D(_0046_),
    .Q_N(_1070_),
    .Q(\bitserial_cipher.state[0] ));
 sg13g2_dfrbp_1 _2079_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net647),
    .D(net332),
    .Q_N(_1069_),
    .Q(\bitserial_cipher.state[1] ));
 sg13g2_dfrbp_1 _2080_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net647),
    .D(net325),
    .Q_N(_1068_),
    .Q(\bitserial_cipher.state[2] ));
 sg13g2_dfrbp_1 _2081_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net647),
    .D(net315),
    .Q_N(_1067_),
    .Q(\bitserial_cipher.state[3] ));
 sg13g2_dfrbp_1 _2082_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net653),
    .D(net328),
    .Q_N(_1066_),
    .Q(\bitserial_cipher.scount[0] ));
 sg13g2_dfrbp_1 _2083_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net653),
    .D(net233),
    .Q_N(_1065_),
    .Q(\bitserial_cipher.scount[1] ));
 sg13g2_dfrbp_1 _2084_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net653),
    .D(net42),
    .Q_N(_1064_),
    .Q(\bitserial_cipher.scount[2] ));
 sg13g2_dfrbp_1 _2085_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net653),
    .D(net31),
    .Q_N(_1063_),
    .Q(\bitserial_cipher.scount[3] ));
 sg13g2_dfrbp_1 _2086_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net654),
    .D(_0054_),
    .Q_N(_1062_),
    .Q(\bitserial_cipher.bcount[0] ));
 sg13g2_dfrbp_1 _2087_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net652),
    .D(_0055_),
    .Q_N(_1061_),
    .Q(\bitserial_cipher.bcount[1] ));
 sg13g2_dfrbp_1 _2088_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net651),
    .D(_0056_),
    .Q_N(_1060_),
    .Q(\bitserial_cipher.bcount[2] ));
 sg13g2_dfrbp_1 _2089_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net651),
    .D(net347),
    .Q_N(_1059_),
    .Q(\bitserial_cipher.bcount[3] ));
 sg13g2_dfrbp_1 _2090_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net639),
    .D(_0058_),
    .Q_N(_1058_),
    .Q(\bitserial_cipher.key[0] ));
 sg13g2_dfrbp_1 _2091_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net639),
    .D(_0059_),
    .Q_N(_1057_),
    .Q(\bitserial_cipher.key[1] ));
 sg13g2_dfrbp_1 _2092_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net639),
    .D(_0060_),
    .Q_N(_1056_),
    .Q(\bitserial_cipher.key[2] ));
 sg13g2_dfrbp_1 _2093_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net626),
    .D(net161),
    .Q_N(_1055_),
    .Q(\bitserial_cipher.key[3] ));
 sg13g2_dfrbp_1 _2094_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net625),
    .D(_0062_),
    .Q_N(_1054_),
    .Q(\bitserial_cipher.key[4] ));
 sg13g2_dfrbp_1 _2095_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net625),
    .D(_0063_),
    .Q_N(_1053_),
    .Q(\bitserial_cipher.key[5] ));
 sg13g2_dfrbp_1 _2096_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net626),
    .D(net39),
    .Q_N(_1052_),
    .Q(\bitserial_cipher.key[6] ));
 sg13g2_dfrbp_1 _2097_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net626),
    .D(net114),
    .Q_N(_1051_),
    .Q(\bitserial_cipher.key[7] ));
 sg13g2_dfrbp_1 _2098_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net626),
    .D(net104),
    .Q_N(_1050_),
    .Q(\bitserial_cipher.key[8] ));
 sg13g2_dfrbp_1 _2099_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net626),
    .D(net192),
    .Q_N(_1049_),
    .Q(\bitserial_cipher.key[9] ));
 sg13g2_dfrbp_1 _2100_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net625),
    .D(net204),
    .Q_N(_1048_),
    .Q(\bitserial_cipher.key[10] ));
 sg13g2_dfrbp_1 _2101_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net625),
    .D(net246),
    .Q_N(_1047_),
    .Q(\bitserial_cipher.key[11] ));
 sg13g2_dfrbp_1 _2102_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net625),
    .D(_0070_),
    .Q_N(_1046_),
    .Q(\bitserial_cipher.key[12] ));
 sg13g2_dfrbp_1 _2103_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net625),
    .D(_0071_),
    .Q_N(_1045_),
    .Q(\bitserial_cipher.key[13] ));
 sg13g2_dfrbp_1 _2104_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net625),
    .D(net84),
    .Q_N(_1044_),
    .Q(\bitserial_cipher.key[14] ));
 sg13g2_dfrbp_1 _2105_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net625),
    .D(net159),
    .Q_N(_1043_),
    .Q(\bitserial_cipher.key[15] ));
 sg13g2_dfrbp_1 _2106_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net621),
    .D(net196),
    .Q_N(_1042_),
    .Q(\bitserial_cipher.key[16] ));
 sg13g2_dfrbp_1 _2107_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net620),
    .D(_0075_),
    .Q_N(_1041_),
    .Q(\bitserial_cipher.key[17] ));
 sg13g2_dfrbp_1 _2108_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net621),
    .D(net60),
    .Q_N(_1040_),
    .Q(\bitserial_cipher.key[18] ));
 sg13g2_dfrbp_1 _2109_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net621),
    .D(net262),
    .Q_N(_1039_),
    .Q(\bitserial_cipher.key[19] ));
 sg13g2_dfrbp_1 _2110_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net620),
    .D(_0078_),
    .Q_N(_1038_),
    .Q(\bitserial_cipher.key[20] ));
 sg13g2_dfrbp_1 _2111_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net621),
    .D(_0079_),
    .Q_N(_1037_),
    .Q(\bitserial_cipher.key[21] ));
 sg13g2_dfrbp_1 _2112_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net620),
    .D(net134),
    .Q_N(_1036_),
    .Q(\bitserial_cipher.key[22] ));
 sg13g2_dfrbp_1 _2113_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net620),
    .D(_0081_),
    .Q_N(_1035_),
    .Q(\bitserial_cipher.key[23] ));
 sg13g2_dfrbp_1 _2114_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net620),
    .D(_0082_),
    .Q_N(_1034_),
    .Q(\bitserial_cipher.key[24] ));
 sg13g2_dfrbp_1 _2115_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net621),
    .D(_0083_),
    .Q_N(_1033_),
    .Q(\bitserial_cipher.key[25] ));
 sg13g2_dfrbp_1 _2116_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net620),
    .D(net164),
    .Q_N(_1032_),
    .Q(\bitserial_cipher.key[26] ));
 sg13g2_dfrbp_1 _2117_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net620),
    .D(net210),
    .Q_N(_1031_),
    .Q(\bitserial_cipher.key[27] ));
 sg13g2_dfrbp_1 _2118_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net620),
    .D(_0086_),
    .Q_N(_1030_),
    .Q(\bitserial_cipher.key[28] ));
 sg13g2_dfrbp_1 _2119_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net618),
    .D(net146),
    .Q_N(_1029_),
    .Q(\bitserial_cipher.key[29] ));
 sg13g2_dfrbp_1 _2120_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net619),
    .D(net220),
    .Q_N(_1028_),
    .Q(\bitserial_cipher.key[30] ));
 sg13g2_dfrbp_1 _2121_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net619),
    .D(net140),
    .Q_N(_1027_),
    .Q(\bitserial_cipher.key[31] ));
 sg13g2_dfrbp_1 _2122_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net619),
    .D(_0090_),
    .Q_N(_1026_),
    .Q(\bitserial_cipher.key[32] ));
 sg13g2_dfrbp_1 _2123_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net618),
    .D(net124),
    .Q_N(_1025_),
    .Q(\bitserial_cipher.key[33] ));
 sg13g2_dfrbp_1 _2124_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net619),
    .D(net94),
    .Q_N(_1024_),
    .Q(\bitserial_cipher.key[34] ));
 sg13g2_dfrbp_1 _2125_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net619),
    .D(_0093_),
    .Q_N(_1023_),
    .Q(\bitserial_cipher.key[35] ));
 sg13g2_dfrbp_1 _2126_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net619),
    .D(net74),
    .Q_N(_1022_),
    .Q(\bitserial_cipher.key[36] ));
 sg13g2_dfrbp_1 _2127_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net618),
    .D(_0095_),
    .Q_N(_1021_),
    .Q(\bitserial_cipher.key[37] ));
 sg13g2_dfrbp_1 _2128_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net619),
    .D(_0096_),
    .Q_N(_1020_),
    .Q(\bitserial_cipher.key[38] ));
 sg13g2_dfrbp_1 _2129_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net619),
    .D(_0097_),
    .Q_N(_1019_),
    .Q(\bitserial_cipher.key[39] ));
 sg13g2_dfrbp_1 _2130_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net618),
    .D(net50),
    .Q_N(_1018_),
    .Q(\bitserial_cipher.key[40] ));
 sg13g2_dfrbp_1 _2131_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net618),
    .D(net173),
    .Q_N(_1017_),
    .Q(\bitserial_cipher.key[41] ));
 sg13g2_dfrbp_1 _2132_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net618),
    .D(net122),
    .Q_N(_1016_),
    .Q(\bitserial_cipher.key[42] ));
 sg13g2_dfrbp_1 _2133_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net618),
    .D(net100),
    .Q_N(_1015_),
    .Q(\bitserial_cipher.key[43] ));
 sg13g2_dfrbp_1 _2134_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net618),
    .D(net238),
    .Q_N(_1014_),
    .Q(\bitserial_cipher.key[44] ));
 sg13g2_dfrbp_1 _2135_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net622),
    .D(_0103_),
    .Q_N(_1013_),
    .Q(\bitserial_cipher.key[45] ));
 sg13g2_dfrbp_1 _2136_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net623),
    .D(net68),
    .Q_N(_1012_),
    .Q(\bitserial_cipher.key[46] ));
 sg13g2_dfrbp_1 _2137_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net623),
    .D(net176),
    .Q_N(_1011_),
    .Q(\bitserial_cipher.key[47] ));
 sg13g2_dfrbp_1 _2138_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net623),
    .D(net153),
    .Q_N(_1010_),
    .Q(\bitserial_cipher.key[48] ));
 sg13g2_dfrbp_1 _2139_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net623),
    .D(_0107_),
    .Q_N(_1009_),
    .Q(\bitserial_cipher.key[49] ));
 sg13g2_dfrbp_1 _2140_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net623),
    .D(net129),
    .Q_N(_1008_),
    .Q(\bitserial_cipher.key[50] ));
 sg13g2_dfrbp_1 _2141_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net624),
    .D(net252),
    .Q_N(_1007_),
    .Q(\bitserial_cipher.key[51] ));
 sg13g2_dfrbp_1 _2142_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net623),
    .D(net189),
    .Q_N(_1006_),
    .Q(\bitserial_cipher.key[52] ));
 sg13g2_dfrbp_1 _2143_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net624),
    .D(_0111_),
    .Q_N(_1005_),
    .Q(\bitserial_cipher.key[53] ));
 sg13g2_dfrbp_1 _2144_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net624),
    .D(net127),
    .Q_N(_1004_),
    .Q(\bitserial_cipher.key[54] ));
 sg13g2_dfrbp_1 _2145_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net623),
    .D(net184),
    .Q_N(_1003_),
    .Q(\bitserial_cipher.key[55] ));
 sg13g2_dfrbp_1 _2146_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net623),
    .D(_0114_),
    .Q_N(_1002_),
    .Q(\bitserial_cipher.key[56] ));
 sg13g2_dfrbp_1 _2147_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net624),
    .D(_0115_),
    .Q_N(_1001_),
    .Q(\bitserial_cipher.key[57] ));
 sg13g2_dfrbp_1 _2148_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net624),
    .D(net148),
    .Q_N(_1000_),
    .Q(\bitserial_cipher.key[58] ));
 sg13g2_dfrbp_1 _2149_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net637),
    .D(_0117_),
    .Q_N(_0999_),
    .Q(\bitserial_cipher.key[59] ));
 sg13g2_dfrbp_1 _2150_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net637),
    .D(net136),
    .Q_N(_0998_),
    .Q(\bitserial_cipher.key[60] ));
 sg13g2_dfrbp_1 _2151_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net637),
    .D(_0119_),
    .Q_N(_0997_),
    .Q(\bitserial_cipher.key[61] ));
 sg13g2_dfrbp_1 _2152_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net637),
    .D(net108),
    .Q_N(_0996_),
    .Q(\bitserial_cipher.key[62] ));
 sg13g2_dfrbp_1 _2153_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net637),
    .D(net178),
    .Q_N(_0995_),
    .Q(\bitserial_cipher.key[63] ));
 sg13g2_dfrbp_1 _2154_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net637),
    .D(_0122_),
    .Q_N(_0994_),
    .Q(\bitserial_cipher.key[64] ));
 sg13g2_dfrbp_1 _2155_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net638),
    .D(_0123_),
    .Q_N(_0993_),
    .Q(\bitserial_cipher.key[65] ));
 sg13g2_dfrbp_1 _2156_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net638),
    .D(net70),
    .Q_N(_0992_),
    .Q(\bitserial_cipher.key[66] ));
 sg13g2_dfrbp_1 _2157_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net638),
    .D(_0125_),
    .Q_N(_0991_),
    .Q(\bitserial_cipher.key[67] ));
 sg13g2_dfrbp_1 _2158_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net638),
    .D(net200),
    .Q_N(_0990_),
    .Q(\bitserial_cipher.key[68] ));
 sg13g2_dfrbp_1 _2159_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net637),
    .D(_0127_),
    .Q_N(_0989_),
    .Q(\bitserial_cipher.key[69] ));
 sg13g2_dfrbp_1 _2160_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net638),
    .D(net119),
    .Q_N(_0988_),
    .Q(\bitserial_cipher.key[70] ));
 sg13g2_dfrbp_1 _2161_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net637),
    .D(_0129_),
    .Q_N(_0987_),
    .Q(\bitserial_cipher.key[71] ));
 sg13g2_dfrbp_1 _2162_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net638),
    .D(_0130_),
    .Q_N(_0986_),
    .Q(\bitserial_cipher.key[72] ));
 sg13g2_dfrbp_1 _2163_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net643),
    .D(_0131_),
    .Q_N(_0985_),
    .Q(\bitserial_cipher.key[73] ));
 sg13g2_dfrbp_1 _2164_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net643),
    .D(net86),
    .Q_N(_0984_),
    .Q(\bitserial_cipher.key[74] ));
 sg13g2_dfrbp_1 _2165_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net643),
    .D(net257),
    .Q_N(_0983_),
    .Q(\bitserial_cipher.key[75] ));
 sg13g2_dfrbp_1 _2166_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net643),
    .D(net151),
    .Q_N(_0982_),
    .Q(\bitserial_cipher.key[76] ));
 sg13g2_dfrbp_1 _2167_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net643),
    .D(_0135_),
    .Q_N(_0981_),
    .Q(\bitserial_cipher.key[77] ));
 sg13g2_dfrbp_1 _2168_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net643),
    .D(net102),
    .Q_N(_0980_),
    .Q(\bitserial_cipher.key[78] ));
 sg13g2_dfrbp_1 _2169_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net642),
    .D(net206),
    .Q_N(_0979_),
    .Q(\bitserial_cipher.key[79] ));
 sg13g2_dfrbp_1 _2170_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net642),
    .D(_0138_),
    .Q_N(_0978_),
    .Q(\bitserial_cipher.key[80] ));
 sg13g2_dfrbp_1 _2171_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net642),
    .D(_0139_),
    .Q_N(_0977_),
    .Q(\bitserial_cipher.key[81] ));
 sg13g2_dfrbp_1 _2172_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net642),
    .D(net56),
    .Q_N(_0976_),
    .Q(\bitserial_cipher.key[82] ));
 sg13g2_dfrbp_1 _2173_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net642),
    .D(net271),
    .Q_N(_0975_),
    .Q(\bitserial_cipher.key[83] ));
 sg13g2_dfrbp_1 _2174_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net646),
    .D(_0142_),
    .Q_N(_0974_),
    .Q(\bitserial_cipher.key[84] ));
 sg13g2_dfrbp_1 _2175_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net646),
    .D(_0143_),
    .Q_N(_0973_),
    .Q(\bitserial_cipher.key[85] ));
 sg13g2_dfrbp_1 _2176_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net642),
    .D(net112),
    .Q_N(_0972_),
    .Q(\bitserial_cipher.key[86] ));
 sg13g2_dfrbp_1 _2177_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net642),
    .D(net157),
    .Q_N(_0971_),
    .Q(\bitserial_cipher.key[87] ));
 sg13g2_dfrbp_1 _2178_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net646),
    .D(_0146_),
    .Q_N(_0970_),
    .Q(\bitserial_cipher.key[88] ));
 sg13g2_dfrbp_1 _2179_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net643),
    .D(_0147_),
    .Q_N(_0969_),
    .Q(\bitserial_cipher.key[89] ));
 sg13g2_dfrbp_1 _2180_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net642),
    .D(net171),
    .Q_N(_0968_),
    .Q(\bitserial_cipher.key[90] ));
 sg13g2_dfrbp_1 _2181_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net644),
    .D(net236),
    .Q_N(_0967_),
    .Q(\bitserial_cipher.key[91] ));
 sg13g2_dfrbp_1 _2182_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net644),
    .D(_0150_),
    .Q_N(_0966_),
    .Q(\bitserial_cipher.key[92] ));
 sg13g2_dfrbp_1 _2183_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net644),
    .D(net144),
    .Q_N(_0965_),
    .Q(\bitserial_cipher.key[93] ));
 sg13g2_dfrbp_1 _2184_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net644),
    .D(net58),
    .Q_N(_0964_),
    .Q(\bitserial_cipher.key[94] ));
 sg13g2_dfrbp_1 _2185_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net644),
    .D(net180),
    .Q_N(_0963_),
    .Q(\bitserial_cipher.key[95] ));
 sg13g2_dfrbp_1 _2186_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net644),
    .D(_0154_),
    .Q_N(_0962_),
    .Q(\bitserial_cipher.key[96] ));
 sg13g2_dfrbp_1 _2187_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net645),
    .D(_0155_),
    .Q_N(_0961_),
    .Q(\bitserial_cipher.key[97] ));
 sg13g2_dfrbp_1 _2188_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net645),
    .D(net92),
    .Q_N(_0960_),
    .Q(\bitserial_cipher.key[98] ));
 sg13g2_dfrbp_1 _2189_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net646),
    .D(net194),
    .Q_N(_0959_),
    .Q(\bitserial_cipher.key[99] ));
 sg13g2_dfrbp_1 _2190_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net644),
    .D(_0158_),
    .Q_N(_0958_),
    .Q(\bitserial_cipher.key[100] ));
 sg13g2_dfrbp_1 _2191_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net644),
    .D(_0159_),
    .Q_N(_0957_),
    .Q(\bitserial_cipher.key[101] ));
 sg13g2_dfrbp_1 _2192_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net652),
    .D(net72),
    .Q_N(_0956_),
    .Q(\bitserial_cipher.key[102] ));
 sg13g2_dfrbp_1 _2193_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net651),
    .D(_0161_),
    .Q_N(_0955_),
    .Q(\bitserial_cipher.key[103] ));
 sg13g2_dfrbp_1 _2194_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net652),
    .D(_0162_),
    .Q_N(_0954_),
    .Q(\bitserial_cipher.key[104] ));
 sg13g2_dfrbp_1 _2195_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net652),
    .D(_0163_),
    .Q_N(_0953_),
    .Q(\bitserial_cipher.key[105] ));
 sg13g2_dfrbp_1 _2196_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net651),
    .D(net64),
    .Q_N(_0952_),
    .Q(\bitserial_cipher.key[106] ));
 sg13g2_dfrbp_1 _2197_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net651),
    .D(net260),
    .Q_N(_0951_),
    .Q(\bitserial_cipher.key[107] ));
 sg13g2_dfrbp_1 _2198_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net651),
    .D(_0166_),
    .Q_N(_0950_),
    .Q(\bitserial_cipher.key[108] ));
 sg13g2_dfrbp_1 _2199_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net651),
    .D(_0167_),
    .Q_N(_0949_),
    .Q(\bitserial_cipher.key[109] ));
 sg13g2_dfrbp_1 _2200_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net651),
    .D(net90),
    .Q_N(_0948_),
    .Q(\bitserial_cipher.key[110] ));
 sg13g2_dfrbp_1 _2201_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net645),
    .D(net168),
    .Q_N(_0947_),
    .Q(\bitserial_cipher.key[111] ));
 sg13g2_dfrbp_1 _2202_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net650),
    .D(net186),
    .Q_N(_0946_),
    .Q(\bitserial_cipher.key[112] ));
 sg13g2_dfrbp_1 _2203_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net645),
    .D(net138),
    .Q_N(_0945_),
    .Q(\bitserial_cipher.key[113] ));
 sg13g2_dfrbp_1 _2204_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net645),
    .D(_0172_),
    .Q_N(_0944_),
    .Q(\bitserial_cipher.key[114] ));
 sg13g2_dfrbp_1 _2205_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net645),
    .D(net155),
    .Q_N(_0943_),
    .Q(\bitserial_cipher.key[115] ));
 sg13g2_dfrbp_1 _2206_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net639),
    .D(_0174_),
    .Q_N(_0942_),
    .Q(\bitserial_cipher.key[116] ));
 sg13g2_dfrbp_1 _2207_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net640),
    .D(net116),
    .Q_N(_0941_),
    .Q(\bitserial_cipher.key[117] ));
 sg13g2_dfrbp_1 _2208_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net645),
    .D(net76),
    .Q_N(_0940_),
    .Q(\bitserial_cipher.key[118] ));
 sg13g2_dfrbp_1 _2209_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net640),
    .D(net250),
    .Q_N(_0939_),
    .Q(\bitserial_cipher.key[119] ));
 sg13g2_dfrbp_1 _2210_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net640),
    .D(_0178_),
    .Q_N(_0938_),
    .Q(\bitserial_cipher.key[120] ));
 sg13g2_dfrbp_1 _2211_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net640),
    .D(_0179_),
    .Q_N(_0937_),
    .Q(\bitserial_cipher.key[121] ));
 sg13g2_dfrbp_1 _2212_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net639),
    .D(net182),
    .Q_N(_0936_),
    .Q(\bitserial_cipher.key[122] ));
 sg13g2_dfrbp_1 _2213_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net639),
    .D(net98),
    .Q_N(_0935_),
    .Q(\bitserial_cipher.key[123] ));
 sg13g2_dfrbp_1 _2214_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net639),
    .D(_0182_),
    .Q_N(_0934_),
    .Q(\bitserial_cipher.key[124] ));
 sg13g2_dfrbp_1 _2215_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net650),
    .D(net284),
    .Q_N(_0933_),
    .Q(\bitserial_cipher.key[125] ));
 sg13g2_dfrbp_1 _2216_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net639),
    .D(_0184_),
    .Q_N(_0932_),
    .Q(\bitserial_cipher.key[126] ));
 sg13g2_dfrbp_1 _2217_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net633),
    .D(net244),
    .Q_N(_0931_),
    .Q(\bitserial_cipher.key[127] ));
 sg13g2_dfrbp_1 _2218_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net654),
    .D(_0186_),
    .Q_N(_0930_),
    .Q(\bitserial_cipher.rcount[0] ));
 sg13g2_dfrbp_1 _2219_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net653),
    .D(net241),
    .Q_N(_0929_),
    .Q(\bitserial_cipher.rcount[1] ));
 sg13g2_dfrbp_1 _2220_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net653),
    .D(net320),
    .Q_N(_0928_),
    .Q(\bitserial_cipher.rcount[2] ));
 sg13g2_dfrbp_1 _2221_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net653),
    .D(net62),
    .Q_N(_0927_),
    .Q(\bitserial_cipher.rcount[3] ));
 sg13g2_dfrbp_1 _2222_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net630),
    .D(_0190_),
    .Q_N(_0926_),
    .Q(\bitserial_cipher.state[36] ));
 sg13g2_dfrbp_1 _2223_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net630),
    .D(net131),
    .Q_N(_0925_),
    .Q(\bitserial_cipher.state[37] ));
 sg13g2_dfrbp_1 _2224_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net630),
    .D(_0192_),
    .Q_N(_0924_),
    .Q(\bitserial_cipher.state[38] ));
 sg13g2_dfrbp_1 _2225_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net630),
    .D(net142),
    .Q_N(_0923_),
    .Q(\bitserial_cipher.state[39] ));
 sg13g2_dfrbp_1 _2226_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net630),
    .D(net222),
    .Q_N(_0922_),
    .Q(\bitserial_cipher.state[40] ));
 sg13g2_dfrbp_1 _2227_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net631),
    .D(net225),
    .Q_N(_0921_),
    .Q(\bitserial_cipher.state[41] ));
 sg13g2_dfrbp_1 _2228_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net631),
    .D(_0196_),
    .Q_N(_0920_),
    .Q(\bitserial_cipher.state[42] ));
 sg13g2_dfrbp_1 _2229_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net631),
    .D(net80),
    .Q_N(_0919_),
    .Q(\bitserial_cipher.state[43] ));
 sg13g2_dfrbp_1 _2230_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net630),
    .D(net292),
    .Q_N(_0918_),
    .Q(\bitserial_cipher.state[32] ));
 sg13g2_dfrbp_1 _2231_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net630),
    .D(net37),
    .Q_N(_0917_),
    .Q(\bitserial_cipher.state[33] ));
 sg13g2_dfrbp_1 _2232_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net630),
    .D(net290),
    .Q_N(_0916_),
    .Q(\bitserial_cipher.state[34] ));
 sg13g2_dfrbp_1 _2233_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net631),
    .D(net106),
    .Q_N(_0915_),
    .Q(\bitserial_cipher.state[35] ));
 sg13g2_dfrbp_1 _2234_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net634),
    .D(net96),
    .Q_N(_0914_),
    .Q(\bitserial_cipher.state[52] ));
 sg13g2_dfrbp_1 _2235_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net635),
    .D(net54),
    .Q_N(_0913_),
    .Q(\bitserial_cipher.state[53] ));
 sg13g2_dfrbp_1 _2236_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net648),
    .D(net52),
    .Q_N(_0912_),
    .Q(\bitserial_cipher.state[54] ));
 sg13g2_dfrbp_1 _2237_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net648),
    .D(_0205_),
    .Q_N(_0911_),
    .Q(\bitserial_cipher.state[55] ));
 sg13g2_dfrbp_1 _2238_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net635),
    .D(_0206_),
    .Q_N(_0910_),
    .Q(\bitserial_cipher.state[56] ));
 sg13g2_dfrbp_1 _2239_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net634),
    .D(net48),
    .Q_N(_0909_),
    .Q(\bitserial_cipher.state[57] ));
 sg13g2_dfrbp_1 _2240_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net648),
    .D(net35),
    .Q_N(_0908_),
    .Q(\bitserial_cipher.state[58] ));
 sg13g2_dfrbp_1 _2241_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net648),
    .D(net82),
    .Q_N(_0907_),
    .Q(\bitserial_cipher.state[59] ));
 sg13g2_dfrbp_1 _2242_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net634),
    .D(_0210_),
    .Q_N(_0906_),
    .Q(\bitserial_cipher.state[44] ));
 sg13g2_tielo tt_um_led_cipher_7 (.L_LO(net7));
 sg13g2_tielo tt_um_led_cipher_8 (.L_LO(net8));
 sg13g2_tielo tt_um_led_cipher_9 (.L_LO(net9));
 sg13g2_tielo tt_um_led_cipher_10 (.L_LO(net10));
 sg13g2_tielo tt_um_led_cipher_11 (.L_LO(net11));
 sg13g2_tielo tt_um_led_cipher_12 (.L_LO(net12));
 sg13g2_tielo tt_um_led_cipher_13 (.L_LO(net13));
 sg13g2_tielo tt_um_led_cipher_14 (.L_LO(net14));
 sg13g2_tielo tt_um_led_cipher_15 (.L_LO(net15));
 sg13g2_tielo tt_um_led_cipher_16 (.L_LO(net16));
 sg13g2_tielo tt_um_led_cipher_17 (.L_LO(net17));
 sg13g2_tielo tt_um_led_cipher_18 (.L_LO(net18));
 sg13g2_tielo tt_um_led_cipher_19 (.L_LO(net19));
 sg13g2_tielo tt_um_led_cipher_20 (.L_LO(net20));
 sg13g2_tielo tt_um_led_cipher_21 (.L_LO(net21));
 sg13g2_tielo tt_um_led_cipher_22 (.L_LO(net22));
 sg13g2_tielo tt_um_led_cipher_23 (.L_LO(net23));
 sg13g2_tielo tt_um_led_cipher_24 (.L_LO(net24));
 sg13g2_tielo tt_um_led_cipher_25 (.L_LO(net25));
 sg13g2_tielo tt_um_led_cipher_26 (.L_LO(net26));
 sg13g2_tielo tt_um_led_cipher_27 (.L_LO(net27));
 sg13g2_buf_2 clkbuf_leaf_0_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_buf_1 _2265_ (.A(\bitserial_cipher.dataq ),
    .X(uo_out[0]));
 sg13g2_buf_1 _2266_ (.A(\bitserial_cipher.done ),
    .X(uo_out[1]));
 sg13g2_buf_2 fanout496 (.A(net497),
    .X(net496));
 sg13g2_buf_2 fanout497 (.A(net499),
    .X(net497));
 sg13g2_buf_2 fanout498 (.A(net499),
    .X(net498));
 sg13g2_buf_1 fanout499 (.A(net502),
    .X(net499));
 sg13g2_buf_2 fanout500 (.A(net501),
    .X(net500));
 sg13g2_buf_2 fanout501 (.A(net502),
    .X(net501));
 sg13g2_buf_2 fanout502 (.A(net510),
    .X(net502));
 sg13g2_buf_2 fanout503 (.A(net504),
    .X(net503));
 sg13g2_buf_2 fanout504 (.A(net510),
    .X(net504));
 sg13g2_buf_2 fanout505 (.A(net506),
    .X(net505));
 sg13g2_buf_2 fanout506 (.A(net509),
    .X(net506));
 sg13g2_buf_2 fanout507 (.A(net508),
    .X(net507));
 sg13g2_buf_2 fanout508 (.A(net509),
    .X(net508));
 sg13g2_buf_2 fanout509 (.A(net510),
    .X(net509));
 sg13g2_buf_2 fanout510 (.A(_0784_),
    .X(net510));
 sg13g2_buf_2 fanout511 (.A(net513),
    .X(net511));
 sg13g2_buf_2 fanout512 (.A(net513),
    .X(net512));
 sg13g2_buf_2 fanout513 (.A(_0570_),
    .X(net513));
 sg13g2_buf_2 fanout514 (.A(net515),
    .X(net514));
 sg13g2_buf_2 fanout515 (.A(_0783_),
    .X(net515));
 sg13g2_buf_2 fanout516 (.A(net519),
    .X(net516));
 sg13g2_buf_2 fanout517 (.A(net519),
    .X(net517));
 sg13g2_buf_1 fanout518 (.A(net519),
    .X(net518));
 sg13g2_buf_2 fanout519 (.A(_0783_),
    .X(net519));
 sg13g2_buf_2 fanout520 (.A(net522),
    .X(net520));
 sg13g2_buf_1 fanout521 (.A(net522),
    .X(net521));
 sg13g2_buf_2 fanout522 (.A(net525),
    .X(net522));
 sg13g2_buf_2 fanout523 (.A(net524),
    .X(net523));
 sg13g2_buf_2 fanout524 (.A(net525),
    .X(net524));
 sg13g2_buf_1 fanout525 (.A(_0782_),
    .X(net525));
 sg13g2_buf_2 fanout526 (.A(net530),
    .X(net526));
 sg13g2_buf_1 fanout527 (.A(net530),
    .X(net527));
 sg13g2_buf_2 fanout528 (.A(net530),
    .X(net528));
 sg13g2_buf_1 fanout529 (.A(net530),
    .X(net529));
 sg13g2_buf_1 fanout530 (.A(_0782_),
    .X(net530));
 sg13g2_buf_2 fanout531 (.A(net542),
    .X(net531));
 sg13g2_buf_1 fanout532 (.A(net542),
    .X(net532));
 sg13g2_buf_2 fanout533 (.A(net535),
    .X(net533));
 sg13g2_buf_2 fanout534 (.A(net535),
    .X(net534));
 sg13g2_buf_2 fanout535 (.A(net542),
    .X(net535));
 sg13g2_buf_2 fanout536 (.A(net537),
    .X(net536));
 sg13g2_buf_1 fanout537 (.A(net541),
    .X(net537));
 sg13g2_buf_2 fanout538 (.A(net541),
    .X(net538));
 sg13g2_buf_2 fanout539 (.A(net541),
    .X(net539));
 sg13g2_buf_2 fanout540 (.A(net541),
    .X(net540));
 sg13g2_buf_1 fanout541 (.A(net542),
    .X(net541));
 sg13g2_buf_1 fanout542 (.A(_0782_),
    .X(net542));
 sg13g2_buf_2 fanout543 (.A(net545),
    .X(net543));
 sg13g2_buf_1 fanout544 (.A(net545),
    .X(net544));
 sg13g2_buf_2 fanout545 (.A(net548),
    .X(net545));
 sg13g2_buf_2 fanout546 (.A(net547),
    .X(net546));
 sg13g2_buf_2 fanout547 (.A(net548),
    .X(net547));
 sg13g2_buf_2 fanout548 (.A(net552),
    .X(net548));
 sg13g2_buf_2 fanout549 (.A(net552),
    .X(net549));
 sg13g2_buf_2 fanout550 (.A(net551),
    .X(net550));
 sg13g2_buf_1 fanout551 (.A(net552),
    .X(net551));
 sg13g2_buf_2 fanout552 (.A(_0654_),
    .X(net552));
 sg13g2_buf_2 fanout553 (.A(net554),
    .X(net553));
 sg13g2_buf_2 fanout554 (.A(_0563_),
    .X(net554));
 sg13g2_buf_2 fanout555 (.A(net556),
    .X(net555));
 sg13g2_buf_2 fanout556 (.A(net562),
    .X(net556));
 sg13g2_buf_1 fanout557 (.A(net562),
    .X(net557));
 sg13g2_buf_2 fanout558 (.A(net559),
    .X(net558));
 sg13g2_buf_2 fanout559 (.A(net562),
    .X(net559));
 sg13g2_buf_4 fanout560 (.X(net560),
    .A(net562));
 sg13g2_buf_1 fanout561 (.A(net562),
    .X(net561));
 sg13g2_buf_2 fanout562 (.A(_0733_),
    .X(net562));
 sg13g2_buf_2 fanout563 (.A(net564),
    .X(net563));
 sg13g2_buf_2 fanout564 (.A(net570),
    .X(net564));
 sg13g2_buf_2 fanout565 (.A(net570),
    .X(net565));
 sg13g2_buf_2 fanout566 (.A(net570),
    .X(net566));
 sg13g2_buf_2 fanout567 (.A(net568),
    .X(net567));
 sg13g2_buf_2 fanout568 (.A(net569),
    .X(net568));
 sg13g2_buf_4 fanout569 (.X(net569),
    .A(net570));
 sg13g2_buf_2 fanout570 (.A(_0733_),
    .X(net570));
 sg13g2_buf_2 fanout571 (.A(net572),
    .X(net571));
 sg13g2_buf_2 fanout572 (.A(net573),
    .X(net572));
 sg13g2_buf_1 fanout573 (.A(_0732_),
    .X(net573));
 sg13g2_buf_2 fanout574 (.A(net578),
    .X(net574));
 sg13g2_buf_2 fanout575 (.A(net578),
    .X(net575));
 sg13g2_buf_2 fanout576 (.A(net578),
    .X(net576));
 sg13g2_buf_2 fanout577 (.A(net578),
    .X(net577));
 sg13g2_buf_1 fanout578 (.A(_0732_),
    .X(net578));
 sg13g2_buf_2 fanout579 (.A(net581),
    .X(net579));
 sg13g2_buf_2 fanout580 (.A(net581),
    .X(net580));
 sg13g2_buf_2 fanout581 (.A(_0562_),
    .X(net581));
 sg13g2_buf_2 fanout582 (.A(_0568_),
    .X(net582));
 sg13g2_buf_2 fanout583 (.A(_0568_),
    .X(net583));
 sg13g2_buf_2 fanout584 (.A(net585),
    .X(net584));
 sg13g2_buf_1 fanout585 (.A(_0567_),
    .X(net585));
 sg13g2_buf_2 fanout586 (.A(net588),
    .X(net586));
 sg13g2_buf_2 fanout587 (.A(net588),
    .X(net587));
 sg13g2_buf_2 fanout588 (.A(_0566_),
    .X(net588));
 sg13g2_buf_2 fanout589 (.A(net590),
    .X(net589));
 sg13g2_buf_2 fanout590 (.A(_0566_),
    .X(net590));
 sg13g2_buf_2 fanout591 (.A(net592),
    .X(net591));
 sg13g2_buf_1 fanout592 (.A(net593),
    .X(net592));
 sg13g2_buf_4 fanout593 (.X(net593),
    .A(_0549_));
 sg13g2_buf_2 fanout594 (.A(net596),
    .X(net594));
 sg13g2_buf_2 fanout595 (.A(net596),
    .X(net595));
 sg13g2_buf_2 fanout596 (.A(_0549_),
    .X(net596));
 sg13g2_buf_4 fanout597 (.X(net597),
    .A(_0548_));
 sg13g2_buf_2 fanout598 (.A(_0548_),
    .X(net598));
 sg13g2_buf_2 fanout599 (.A(net601),
    .X(net599));
 sg13g2_buf_1 fanout600 (.A(net601),
    .X(net600));
 sg13g2_buf_2 fanout601 (.A(_0547_),
    .X(net601));
 sg13g2_buf_2 fanout602 (.A(net603),
    .X(net602));
 sg13g2_buf_2 fanout603 (.A(net604),
    .X(net603));
 sg13g2_buf_1 fanout604 (.A(net609),
    .X(net604));
 sg13g2_buf_2 fanout605 (.A(net608),
    .X(net605));
 sg13g2_buf_1 fanout606 (.A(net608),
    .X(net606));
 sg13g2_buf_2 fanout607 (.A(net608),
    .X(net607));
 sg13g2_buf_2 fanout608 (.A(net609),
    .X(net608));
 sg13g2_buf_2 fanout609 (.A(_0539_),
    .X(net609));
 sg13g2_buf_4 fanout610 (.X(net610),
    .A(net611));
 sg13g2_buf_2 fanout611 (.A(_0525_),
    .X(net611));
 sg13g2_buf_2 fanout612 (.A(net614),
    .X(net612));
 sg13g2_buf_2 fanout613 (.A(net614),
    .X(net613));
 sg13g2_buf_1 fanout614 (.A(net615),
    .X(net614));
 sg13g2_buf_2 fanout615 (.A(_0522_),
    .X(net615));
 sg13g2_buf_2 fanout616 (.A(_0511_),
    .X(net616));
 sg13g2_buf_2 fanout617 (.A(\bitserial_cipher.ctlstate[3] ),
    .X(net617));
 sg13g2_buf_4 fanout618 (.X(net618),
    .A(net622));
 sg13g2_buf_4 fanout619 (.X(net619),
    .A(net622));
 sg13g2_buf_4 fanout620 (.X(net620),
    .A(net622));
 sg13g2_buf_2 fanout621 (.A(net622),
    .X(net621));
 sg13g2_buf_2 fanout622 (.A(net636),
    .X(net622));
 sg13g2_buf_4 fanout623 (.X(net623),
    .A(net627));
 sg13g2_buf_2 fanout624 (.A(net627),
    .X(net624));
 sg13g2_buf_4 fanout625 (.X(net625),
    .A(net627));
 sg13g2_buf_4 fanout626 (.X(net626),
    .A(net627));
 sg13g2_buf_2 fanout627 (.A(net636),
    .X(net627));
 sg13g2_buf_4 fanout628 (.X(net628),
    .A(net629));
 sg13g2_buf_4 fanout629 (.X(net629),
    .A(net636));
 sg13g2_buf_4 fanout630 (.X(net630),
    .A(net631));
 sg13g2_buf_4 fanout631 (.X(net631),
    .A(net636));
 sg13g2_buf_4 fanout632 (.X(net632),
    .A(net635));
 sg13g2_buf_2 fanout633 (.A(net635),
    .X(net633));
 sg13g2_buf_4 fanout634 (.X(net634),
    .A(net635));
 sg13g2_buf_4 fanout635 (.X(net635),
    .A(net636));
 sg13g2_buf_2 fanout636 (.A(net656),
    .X(net636));
 sg13g2_buf_4 fanout637 (.X(net637),
    .A(net641));
 sg13g2_buf_4 fanout638 (.X(net638),
    .A(net641));
 sg13g2_buf_4 fanout639 (.X(net639),
    .A(net641));
 sg13g2_buf_2 fanout640 (.A(net641),
    .X(net640));
 sg13g2_buf_1 fanout641 (.A(net656),
    .X(net641));
 sg13g2_buf_4 fanout642 (.X(net642),
    .A(net643));
 sg13g2_buf_4 fanout643 (.X(net643),
    .A(net646));
 sg13g2_buf_4 fanout644 (.X(net644),
    .A(net645));
 sg13g2_buf_4 fanout645 (.X(net645),
    .A(net646));
 sg13g2_buf_4 fanout646 (.X(net646),
    .A(net656));
 sg13g2_buf_4 fanout647 (.X(net647),
    .A(net650));
 sg13g2_buf_4 fanout648 (.X(net648),
    .A(net650));
 sg13g2_buf_2 fanout649 (.A(net650),
    .X(net649));
 sg13g2_buf_2 fanout650 (.A(net655),
    .X(net650));
 sg13g2_buf_4 fanout651 (.X(net651),
    .A(net655));
 sg13g2_buf_2 fanout652 (.A(net655),
    .X(net652));
 sg13g2_buf_4 fanout653 (.X(net653),
    .A(net654));
 sg13g2_buf_4 fanout654 (.X(net654),
    .A(net655));
 sg13g2_buf_2 fanout655 (.A(net656),
    .X(net655));
 sg13g2_buf_1 fanout656 (.A(rst_n),
    .X(net656));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[2]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[3]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[4]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[5]),
    .X(net5));
 sg13g2_tielo tt_um_led_cipher_6 (.L_LO(net6));
 sg13g2_buf_2 clkbuf_leaf_1_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_2 clkbuf_leaf_2_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_2 clkbuf_leaf_3_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_2 clkbuf_leaf_4_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_2 clkbuf_leaf_5_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_2 clkbuf_leaf_6_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_2 clkbuf_leaf_7_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_2 clkbuf_leaf_8_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_2 clkbuf_leaf_9_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_2 clkbuf_leaf_10_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_2 clkbuf_leaf_11_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_2 clkbuf_leaf_12_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_2 clkbuf_leaf_13_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_2 clkbuf_leaf_14_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_2 clkbuf_leaf_15_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_2 clkbuf_leaf_16_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_2 clkbuf_leaf_17_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_2 clkbuf_leaf_18_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_2 clkbuf_leaf_19_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_2 clkbuf_leaf_20_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_2 clkbuf_leaf_21_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_2 clkbuf_leaf_22_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_2 clkbuf_leaf_23_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_2 clkbuf_leaf_24_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_2 clkbuf_leaf_25_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_2 clkbuf_leaf_26_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_2 clkbuf_leaf_27_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_2 clkbuf_leaf_28_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_2 clkbuf_leaf_29_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_2 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sg13g2_buf_2 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sg13g2_buf_2 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sg13g2_buf_2 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sg13g2_buf_2 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sg13g2_buf_2 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sg13g2_buf_2 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sg13g2_buf_2 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sg13g2_buf_2 clkload0 (.A(clknet_3_3__leaf_clk));
 sg13g2_buf_2 clkload1 (.A(clknet_3_7__leaf_clk));
 sg13g2_inv_2 clkload2 (.A(clknet_leaf_1_clk));
 sg13g2_inv_4 clkload3 (.A(clknet_leaf_29_clk));
 sg13g2_inv_4 clkload4 (.A(clknet_leaf_25_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_leaf_26_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_leaf_5_clk));
 sg13g2_inv_1 clkload7 (.A(clknet_leaf_7_clk));
 sg13g2_inv_4 clkload8 (.A(clknet_leaf_9_clk));
 sg13g2_inv_8 clkload9 (.A(clknet_leaf_10_clk));
 sg13g2_inv_2 clkload10 (.A(clknet_leaf_22_clk));
 sg13g2_inv_1 clkload11 (.A(clknet_leaf_11_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\bitserial_cipher.rc[0] ),
    .X(net28));
 sg13g2_dlygate4sd3_1 hold2 (.A(_0640_),
    .X(net29));
 sg13g2_dlygate4sd3_1 hold3 (.A(\bitserial_cipher.scount[3] ),
    .X(net30));
 sg13g2_dlygate4sd3_1 hold4 (.A(_0053_),
    .X(net31));
 sg13g2_dlygate4sd3_1 hold5 (.A(_0000_),
    .X(net32));
 sg13g2_dlygate4sd3_1 hold6 (.A(_0639_),
    .X(net33));
 sg13g2_dlygate4sd3_1 hold7 (.A(\bitserial_cipher.state[57] ),
    .X(net34));
 sg13g2_dlygate4sd3_1 hold8 (.A(_0208_),
    .X(net35));
 sg13g2_dlygate4sd3_1 hold9 (.A(\bitserial_cipher.state[32] ),
    .X(net36));
 sg13g2_dlygate4sd3_1 hold10 (.A(_0199_),
    .X(net37));
 sg13g2_dlygate4sd3_1 hold11 (.A(\bitserial_cipher.key[5] ),
    .X(net38));
 sg13g2_dlygate4sd3_1 hold12 (.A(_0064_),
    .X(net39));
 sg13g2_dlygate4sd3_1 hold13 (.A(\bitserial_cipher.scount[2] ),
    .X(net40));
 sg13g2_dlygate4sd3_1 hold14 (.A(_0770_),
    .X(net41));
 sg13g2_dlygate4sd3_1 hold15 (.A(_0052_),
    .X(net42));
 sg13g2_dlygate4sd3_1 hold16 (.A(\bitserial_cipher.rc[3] ),
    .X(net43));
 sg13g2_dlygate4sd3_1 hold17 (.A(_0642_),
    .X(net44));
 sg13g2_dlygate4sd3_1 hold18 (.A(\bitserial_cipher.rc[2] ),
    .X(net45));
 sg13g2_dlygate4sd3_1 hold19 (.A(_0641_),
    .X(net46));
 sg13g2_dlygate4sd3_1 hold20 (.A(\bitserial_cipher.state[56] ),
    .X(net47));
 sg13g2_dlygate4sd3_1 hold21 (.A(_0207_),
    .X(net48));
 sg13g2_dlygate4sd3_1 hold22 (.A(\bitserial_cipher.key[39] ),
    .X(net49));
 sg13g2_dlygate4sd3_1 hold23 (.A(_0098_),
    .X(net50));
 sg13g2_dlygate4sd3_1 hold24 (.A(\bitserial_cipher.state[54] ),
    .X(net51));
 sg13g2_dlygate4sd3_1 hold25 (.A(_0204_),
    .X(net52));
 sg13g2_dlygate4sd3_1 hold26 (.A(\bitserial_cipher.state[52] ),
    .X(net53));
 sg13g2_dlygate4sd3_1 hold27 (.A(_0203_),
    .X(net54));
 sg13g2_dlygate4sd3_1 hold28 (.A(\bitserial_cipher.key[81] ),
    .X(net55));
 sg13g2_dlygate4sd3_1 hold29 (.A(_0140_),
    .X(net56));
 sg13g2_dlygate4sd3_1 hold30 (.A(\bitserial_cipher.key[93] ),
    .X(net57));
 sg13g2_dlygate4sd3_1 hold31 (.A(_0152_),
    .X(net58));
 sg13g2_dlygate4sd3_1 hold32 (.A(\bitserial_cipher.key[17] ),
    .X(net59));
 sg13g2_dlygate4sd3_1 hold33 (.A(_0076_),
    .X(net60));
 sg13g2_dlygate4sd3_1 hold34 (.A(\bitserial_cipher.rcount[3] ),
    .X(net61));
 sg13g2_dlygate4sd3_1 hold35 (.A(_0189_),
    .X(net62));
 sg13g2_dlygate4sd3_1 hold36 (.A(\bitserial_cipher.key[105] ),
    .X(net63));
 sg13g2_dlygate4sd3_1 hold37 (.A(_0164_),
    .X(net64));
 sg13g2_dlygate4sd3_1 hold38 (.A(\bitserial_cipher.rc[5] ),
    .X(net65));
 sg13g2_dlygate4sd3_1 hold39 (.A(_0644_),
    .X(net66));
 sg13g2_dlygate4sd3_1 hold40 (.A(\bitserial_cipher.key[45] ),
    .X(net67));
 sg13g2_dlygate4sd3_1 hold41 (.A(_0104_),
    .X(net68));
 sg13g2_dlygate4sd3_1 hold42 (.A(\bitserial_cipher.key[65] ),
    .X(net69));
 sg13g2_dlygate4sd3_1 hold43 (.A(_0124_),
    .X(net70));
 sg13g2_dlygate4sd3_1 hold44 (.A(\bitserial_cipher.key[101] ),
    .X(net71));
 sg13g2_dlygate4sd3_1 hold45 (.A(_0160_),
    .X(net72));
 sg13g2_dlygate4sd3_1 hold46 (.A(\bitserial_cipher.key[35] ),
    .X(net73));
 sg13g2_dlygate4sd3_1 hold47 (.A(_0094_),
    .X(net74));
 sg13g2_dlygate4sd3_1 hold48 (.A(\bitserial_cipher.key[117] ),
    .X(net75));
 sg13g2_dlygate4sd3_1 hold49 (.A(_0176_),
    .X(net76));
 sg13g2_dlygate4sd3_1 hold50 (.A(\bitserial_cipher.key[0] ),
    .X(net77));
 sg13g2_dlygate4sd3_1 hold51 (.A(_0785_),
    .X(net78));
 sg13g2_dlygate4sd3_1 hold52 (.A(\bitserial_cipher.state[42] ),
    .X(net79));
 sg13g2_dlygate4sd3_1 hold53 (.A(_0197_),
    .X(net80));
 sg13g2_dlygate4sd3_1 hold54 (.A(\bitserial_cipher.state[58] ),
    .X(net81));
 sg13g2_dlygate4sd3_1 hold55 (.A(_0209_),
    .X(net82));
 sg13g2_dlygate4sd3_1 hold56 (.A(\bitserial_cipher.key[13] ),
    .X(net83));
 sg13g2_dlygate4sd3_1 hold57 (.A(_0072_),
    .X(net84));
 sg13g2_dlygate4sd3_1 hold58 (.A(\bitserial_cipher.key[73] ),
    .X(net85));
 sg13g2_dlygate4sd3_1 hold59 (.A(_0132_),
    .X(net86));
 sg13g2_dlygate4sd3_1 hold60 (.A(\bitserial_cipher.state[55] ),
    .X(net87));
 sg13g2_dlygate4sd3_1 hold61 (.A(_0439_),
    .X(net88));
 sg13g2_dlygate4sd3_1 hold62 (.A(\bitserial_cipher.key[109] ),
    .X(net89));
 sg13g2_dlygate4sd3_1 hold63 (.A(_0168_),
    .X(net90));
 sg13g2_dlygate4sd3_1 hold64 (.A(\bitserial_cipher.key[97] ),
    .X(net91));
 sg13g2_dlygate4sd3_1 hold65 (.A(_0156_),
    .X(net92));
 sg13g2_dlygate4sd3_1 hold66 (.A(\bitserial_cipher.key[33] ),
    .X(net93));
 sg13g2_dlygate4sd3_1 hold67 (.A(_0092_),
    .X(net94));
 sg13g2_dlygate4sd3_1 hold68 (.A(\bitserial_cipher.state[51] ),
    .X(net95));
 sg13g2_dlygate4sd3_1 hold69 (.A(_0202_),
    .X(net96));
 sg13g2_dlygate4sd3_1 hold70 (.A(\bitserial_cipher.key[123] ),
    .X(net97));
 sg13g2_dlygate4sd3_1 hold71 (.A(_0181_),
    .X(net98));
 sg13g2_dlygate4sd3_1 hold72 (.A(\bitserial_cipher.key[42] ),
    .X(net99));
 sg13g2_dlygate4sd3_1 hold73 (.A(_0101_),
    .X(net100));
 sg13g2_dlygate4sd3_1 hold74 (.A(\bitserial_cipher.key[77] ),
    .X(net101));
 sg13g2_dlygate4sd3_1 hold75 (.A(_0136_),
    .X(net102));
 sg13g2_dlygate4sd3_1 hold76 (.A(\bitserial_cipher.key[4] ),
    .X(net103));
 sg13g2_dlygate4sd3_1 hold77 (.A(_0066_),
    .X(net104));
 sg13g2_dlygate4sd3_1 hold78 (.A(\bitserial_cipher.state[34] ),
    .X(net105));
 sg13g2_dlygate4sd3_1 hold79 (.A(_0201_),
    .X(net106));
 sg13g2_dlygate4sd3_1 hold80 (.A(\bitserial_cipher.key[61] ),
    .X(net107));
 sg13g2_dlygate4sd3_1 hold81 (.A(_0120_),
    .X(net108));
 sg13g2_dlygate4sd3_1 hold82 (.A(\bitserial_cipher.state[48] ),
    .X(net109));
 sg13g2_dlygate4sd3_1 hold83 (.A(_0005_),
    .X(net110));
 sg13g2_dlygate4sd3_1 hold84 (.A(\bitserial_cipher.key[85] ),
    .X(net111));
 sg13g2_dlygate4sd3_1 hold85 (.A(_0144_),
    .X(net112));
 sg13g2_dlygate4sd3_1 hold86 (.A(\bitserial_cipher.key[3] ),
    .X(net113));
 sg13g2_dlygate4sd3_1 hold87 (.A(_0065_),
    .X(net114));
 sg13g2_dlygate4sd3_1 hold88 (.A(\bitserial_cipher.key[116] ),
    .X(net115));
 sg13g2_dlygate4sd3_1 hold89 (.A(_0175_),
    .X(net116));
 sg13g2_dlygate4sd3_1 hold90 (.A(\bitserial_cipher.state[0] ),
    .X(net117));
 sg13g2_dlygate4sd3_1 hold91 (.A(\bitserial_cipher.key[69] ),
    .X(net118));
 sg13g2_dlygate4sd3_1 hold92 (.A(_0128_),
    .X(net119));
 sg13g2_dlygate4sd3_1 hold93 (.A(\bitserial_cipher.key[68] ),
    .X(net120));
 sg13g2_dlygate4sd3_1 hold94 (.A(\bitserial_cipher.key[41] ),
    .X(net121));
 sg13g2_dlygate4sd3_1 hold95 (.A(_0100_),
    .X(net122));
 sg13g2_dlygate4sd3_1 hold96 (.A(\bitserial_cipher.key[32] ),
    .X(net123));
 sg13g2_dlygate4sd3_1 hold97 (.A(_0091_),
    .X(net124));
 sg13g2_dlygate4sd3_1 hold98 (.A(\bitserial_cipher.key[84] ),
    .X(net125));
 sg13g2_dlygate4sd3_1 hold99 (.A(\bitserial_cipher.key[53] ),
    .X(net126));
 sg13g2_dlygate4sd3_1 hold100 (.A(_0112_),
    .X(net127));
 sg13g2_dlygate4sd3_1 hold101 (.A(\bitserial_cipher.key[49] ),
    .X(net128));
 sg13g2_dlygate4sd3_1 hold102 (.A(_0108_),
    .X(net129));
 sg13g2_dlygate4sd3_1 hold103 (.A(\bitserial_cipher.state[37] ),
    .X(net130));
 sg13g2_dlygate4sd3_1 hold104 (.A(_0191_),
    .X(net131));
 sg13g2_dlygate4sd3_1 hold105 (.A(\bitserial_cipher.key[1] ),
    .X(net132));
 sg13g2_dlygate4sd3_1 hold106 (.A(\bitserial_cipher.key[21] ),
    .X(net133));
 sg13g2_dlygate4sd3_1 hold107 (.A(_0080_),
    .X(net134));
 sg13g2_dlygate4sd3_1 hold108 (.A(\bitserial_cipher.key[59] ),
    .X(net135));
 sg13g2_dlygate4sd3_1 hold109 (.A(_0118_),
    .X(net136));
 sg13g2_dlygate4sd3_1 hold110 (.A(\bitserial_cipher.key[112] ),
    .X(net137));
 sg13g2_dlygate4sd3_1 hold111 (.A(_0171_),
    .X(net138));
 sg13g2_dlygate4sd3_1 hold112 (.A(\bitserial_cipher.key[27] ),
    .X(net139));
 sg13g2_dlygate4sd3_1 hold113 (.A(_0089_),
    .X(net140));
 sg13g2_dlygate4sd3_1 hold114 (.A(\bitserial_cipher.state[35] ),
    .X(net141));
 sg13g2_dlygate4sd3_1 hold115 (.A(_0193_),
    .X(net142));
 sg13g2_dlygate4sd3_1 hold116 (.A(\bitserial_cipher.key[92] ),
    .X(net143));
 sg13g2_dlygate4sd3_1 hold117 (.A(_0151_),
    .X(net144));
 sg13g2_dlygate4sd3_1 hold118 (.A(\bitserial_cipher.key[28] ),
    .X(net145));
 sg13g2_dlygate4sd3_1 hold119 (.A(_0087_),
    .X(net146));
 sg13g2_dlygate4sd3_1 hold120 (.A(\bitserial_cipher.key[57] ),
    .X(net147));
 sg13g2_dlygate4sd3_1 hold121 (.A(_0116_),
    .X(net148));
 sg13g2_dlygate4sd3_1 hold122 (.A(\bitserial_cipher.key[20] ),
    .X(net149));
 sg13g2_dlygate4sd3_1 hold123 (.A(\bitserial_cipher.key[72] ),
    .X(net150));
 sg13g2_dlygate4sd3_1 hold124 (.A(_0134_),
    .X(net151));
 sg13g2_dlygate4sd3_1 hold125 (.A(\bitserial_cipher.key[44] ),
    .X(net152));
 sg13g2_dlygate4sd3_1 hold126 (.A(_0106_),
    .X(net153));
 sg13g2_dlygate4sd3_1 hold127 (.A(\bitserial_cipher.key[114] ),
    .X(net154));
 sg13g2_dlygate4sd3_1 hold128 (.A(_0173_),
    .X(net155));
 sg13g2_dlygate4sd3_1 hold129 (.A(\bitserial_cipher.key[86] ),
    .X(net156));
 sg13g2_dlygate4sd3_1 hold130 (.A(_0145_),
    .X(net157));
 sg13g2_dlygate4sd3_1 hold131 (.A(\bitserial_cipher.key[14] ),
    .X(net158));
 sg13g2_dlygate4sd3_1 hold132 (.A(_0073_),
    .X(net159));
 sg13g2_dlygate4sd3_1 hold133 (.A(\bitserial_cipher.key[2] ),
    .X(net160));
 sg13g2_dlygate4sd3_1 hold134 (.A(_0061_),
    .X(net161));
 sg13g2_dlygate4sd3_1 hold135 (.A(\bitserial_cipher.state[47] ),
    .X(net162));
 sg13g2_dlygate4sd3_1 hold136 (.A(\bitserial_cipher.key[22] ),
    .X(net163));
 sg13g2_dlygate4sd3_1 hold137 (.A(_0084_),
    .X(net164));
 sg13g2_dlygate4sd3_1 hold138 (.A(\bitserial_cipher.key[56] ),
    .X(net165));
 sg13g2_dlygate4sd3_1 hold139 (.A(\bitserial_cipher.key[38] ),
    .X(net166));
 sg13g2_dlygate4sd3_1 hold140 (.A(\bitserial_cipher.key[110] ),
    .X(net167));
 sg13g2_dlygate4sd3_1 hold141 (.A(_0169_),
    .X(net168));
 sg13g2_dlygate4sd3_1 hold142 (.A(\bitserial_cipher.key[113] ),
    .X(net169));
 sg13g2_dlygate4sd3_1 hold143 (.A(\bitserial_cipher.key[89] ),
    .X(net170));
 sg13g2_dlygate4sd3_1 hold144 (.A(_0148_),
    .X(net171));
 sg13g2_dlygate4sd3_1 hold145 (.A(\bitserial_cipher.key[37] ),
    .X(net172));
 sg13g2_dlygate4sd3_1 hold146 (.A(_0099_),
    .X(net173));
 sg13g2_dlygate4sd3_1 hold147 (.A(\bitserial_cipher.rc[4] ),
    .X(net174));
 sg13g2_dlygate4sd3_1 hold148 (.A(\bitserial_cipher.key[46] ),
    .X(net175));
 sg13g2_dlygate4sd3_1 hold149 (.A(_0105_),
    .X(net176));
 sg13g2_dlygate4sd3_1 hold150 (.A(\bitserial_cipher.key[63] ),
    .X(net177));
 sg13g2_dlygate4sd3_1 hold151 (.A(_0121_),
    .X(net178));
 sg13g2_dlygate4sd3_1 hold152 (.A(\bitserial_cipher.key[91] ),
    .X(net179));
 sg13g2_dlygate4sd3_1 hold153 (.A(_0153_),
    .X(net180));
 sg13g2_dlygate4sd3_1 hold154 (.A(\bitserial_cipher.key[121] ),
    .X(net181));
 sg13g2_dlygate4sd3_1 hold155 (.A(_0180_),
    .X(net182));
 sg13g2_dlygate4sd3_1 hold156 (.A(\bitserial_cipher.key[54] ),
    .X(net183));
 sg13g2_dlygate4sd3_1 hold157 (.A(_0113_),
    .X(net184));
 sg13g2_dlygate4sd3_1 hold158 (.A(\bitserial_cipher.key[108] ),
    .X(net185));
 sg13g2_dlygate4sd3_1 hold159 (.A(_0170_),
    .X(net186));
 sg13g2_dlygate4sd3_1 hold160 (.A(\bitserial_cipher.key[48] ),
    .X(net187));
 sg13g2_dlygate4sd3_1 hold161 (.A(\bitserial_cipher.key[51] ),
    .X(net188));
 sg13g2_dlygate4sd3_1 hold162 (.A(_0110_),
    .X(net189));
 sg13g2_dlygate4sd3_1 hold163 (.A(\bitserial_cipher.key[120] ),
    .X(net190));
 sg13g2_dlygate4sd3_1 hold164 (.A(\bitserial_cipher.key[8] ),
    .X(net191));
 sg13g2_dlygate4sd3_1 hold165 (.A(_0067_),
    .X(net192));
 sg13g2_dlygate4sd3_1 hold166 (.A(\bitserial_cipher.key[95] ),
    .X(net193));
 sg13g2_dlygate4sd3_1 hold167 (.A(_0157_),
    .X(net194));
 sg13g2_dlygate4sd3_1 hold168 (.A(\bitserial_cipher.key[12] ),
    .X(net195));
 sg13g2_dlygate4sd3_1 hold169 (.A(_0074_),
    .X(net196));
 sg13g2_dlygate4sd3_1 hold170 (.A(\bitserial_cipher.state[38] ),
    .X(net197));
 sg13g2_dlygate4sd3_1 hold171 (.A(\bitserial_cipher.key[60] ),
    .X(net198));
 sg13g2_dlygate4sd3_1 hold172 (.A(\bitserial_cipher.key[67] ),
    .X(net199));
 sg13g2_dlygate4sd3_1 hold173 (.A(_0126_),
    .X(net200));
 sg13g2_dlygate4sd3_1 hold174 (.A(\bitserial_cipher.key[71] ),
    .X(net201));
 sg13g2_dlygate4sd3_1 hold175 (.A(\bitserial_cipher.key[66] ),
    .X(net202));
 sg13g2_dlygate4sd3_1 hold176 (.A(\bitserial_cipher.key[9] ),
    .X(net203));
 sg13g2_dlygate4sd3_1 hold177 (.A(_0068_),
    .X(net204));
 sg13g2_dlygate4sd3_1 hold178 (.A(\bitserial_cipher.key[78] ),
    .X(net205));
 sg13g2_dlygate4sd3_1 hold179 (.A(_0137_),
    .X(net206));
 sg13g2_dlygate4sd3_1 hold180 (.A(\bitserial_cipher.key[36] ),
    .X(net207));
 sg13g2_dlygate4sd3_1 hold181 (.A(\bitserial_cipher.key[24] ),
    .X(net208));
 sg13g2_dlygate4sd3_1 hold182 (.A(\bitserial_cipher.key[23] ),
    .X(net209));
 sg13g2_dlygate4sd3_1 hold183 (.A(_0085_),
    .X(net210));
 sg13g2_dlygate4sd3_1 hold184 (.A(\bitserial_cipher.key[88] ),
    .X(net211));
 sg13g2_dlygate4sd3_1 hold185 (.A(\bitserial_cipher.key[64] ),
    .X(net212));
 sg13g2_dlygate4sd3_1 hold186 (.A(\bitserial_cipher.key[52] ),
    .X(net213));
 sg13g2_dlygate4sd3_1 hold187 (.A(\bitserial_cipher.key[31] ),
    .X(net214));
 sg13g2_dlygate4sd3_1 hold188 (.A(\bitserial_cipher.state[20] ),
    .X(net215));
 sg13g2_dlygate4sd3_1 hold189 (.A(_0034_),
    .X(net216));
 sg13g2_dlygate4sd3_1 hold190 (.A(\bitserial_cipher.key[55] ),
    .X(net217));
 sg13g2_dlygate4sd3_1 hold191 (.A(\bitserial_cipher.key[96] ),
    .X(net218));
 sg13g2_dlygate4sd3_1 hold192 (.A(\bitserial_cipher.key[26] ),
    .X(net219));
 sg13g2_dlygate4sd3_1 hold193 (.A(_0088_),
    .X(net220));
 sg13g2_dlygate4sd3_1 hold194 (.A(\bitserial_cipher.state[36] ),
    .X(net221));
 sg13g2_dlygate4sd3_1 hold195 (.A(_0194_),
    .X(net222));
 sg13g2_dlygate4sd3_1 hold196 (.A(\bitserial_cipher.key[70] ),
    .X(net223));
 sg13g2_dlygate4sd3_1 hold197 (.A(\bitserial_cipher.state[41] ),
    .X(net224));
 sg13g2_dlygate4sd3_1 hold198 (.A(_0195_),
    .X(net225));
 sg13g2_dlygate4sd3_1 hold199 (.A(\bitserial_cipher.key[76] ),
    .X(net226));
 sg13g2_dlygate4sd3_1 hold200 (.A(\bitserial_cipher.key[115] ),
    .X(net227));
 sg13g2_dlygate4sd3_1 hold201 (.A(\bitserial_cipher.state[49] ),
    .X(net228));
 sg13g2_dlygate4sd3_1 hold202 (.A(_0006_),
    .X(net229));
 sg13g2_dlygate4sd3_1 hold203 (.A(\bitserial_cipher.key[25] ),
    .X(net230));
 sg13g2_dlygate4sd3_1 hold204 (.A(\bitserial_cipher.key[100] ),
    .X(net231));
 sg13g2_dlygate4sd3_1 hold205 (.A(\bitserial_cipher.scount[1] ),
    .X(net232));
 sg13g2_dlygate4sd3_1 hold206 (.A(_0051_),
    .X(net233));
 sg13g2_dlygate4sd3_1 hold207 (.A(\bitserial_cipher.key[104] ),
    .X(net234));
 sg13g2_dlygate4sd3_1 hold208 (.A(\bitserial_cipher.key[90] ),
    .X(net235));
 sg13g2_dlygate4sd3_1 hold209 (.A(_0149_),
    .X(net236));
 sg13g2_dlygate4sd3_1 hold210 (.A(\bitserial_cipher.key[40] ),
    .X(net237));
 sg13g2_dlygate4sd3_1 hold211 (.A(_0102_),
    .X(net238));
 sg13g2_dlygate4sd3_1 hold212 (.A(\bitserial_cipher.rcount[1] ),
    .X(net239));
 sg13g2_dlygate4sd3_1 hold213 (.A(_0407_),
    .X(net240));
 sg13g2_dlygate4sd3_1 hold214 (.A(_0187_),
    .X(net241));
 sg13g2_dlygate4sd3_1 hold215 (.A(\bitserial_cipher.key[80] ),
    .X(net242));
 sg13g2_dlygate4sd3_1 hold216 (.A(\bitserial_cipher.key[127] ),
    .X(net243));
 sg13g2_dlygate4sd3_1 hold217 (.A(_0185_),
    .X(net244));
 sg13g2_dlygate4sd3_1 hold218 (.A(\bitserial_cipher.key[7] ),
    .X(net245));
 sg13g2_dlygate4sd3_1 hold219 (.A(_0069_),
    .X(net246));
 sg13g2_dlygate4sd3_1 hold220 (.A(\bitserial_cipher.key[99] ),
    .X(net247));
 sg13g2_dlygate4sd3_1 hold221 (.A(\bitserial_cipher.key[87] ),
    .X(net248));
 sg13g2_dlygate4sd3_1 hold222 (.A(\bitserial_cipher.key[119] ),
    .X(net249));
 sg13g2_dlygate4sd3_1 hold223 (.A(_0177_),
    .X(net250));
 sg13g2_dlygate4sd3_1 hold224 (.A(\bitserial_cipher.key[47] ),
    .X(net251));
 sg13g2_dlygate4sd3_1 hold225 (.A(_0109_),
    .X(net252));
 sg13g2_dlygate4sd3_1 hold226 (.A(\bitserial_cipher.key[58] ),
    .X(net253));
 sg13g2_dlygate4sd3_1 hold227 (.A(\bitserial_cipher.key[16] ),
    .X(net254));
 sg13g2_dlygate4sd3_1 hold228 (.A(\bitserial_cipher.key[34] ),
    .X(net255));
 sg13g2_dlygate4sd3_1 hold229 (.A(\bitserial_cipher.key[75] ),
    .X(net256));
 sg13g2_dlygate4sd3_1 hold230 (.A(_0133_),
    .X(net257));
 sg13g2_dlygate4sd3_1 hold231 (.A(\bitserial_cipher.key[19] ),
    .X(net258));
 sg13g2_dlygate4sd3_1 hold232 (.A(\bitserial_cipher.key[103] ),
    .X(net259));
 sg13g2_dlygate4sd3_1 hold233 (.A(_0165_),
    .X(net260));
 sg13g2_dlygate4sd3_1 hold234 (.A(\bitserial_cipher.key[15] ),
    .X(net261));
 sg13g2_dlygate4sd3_1 hold235 (.A(_0077_),
    .X(net262));
 sg13g2_dlygate4sd3_1 hold236 (.A(\bitserial_cipher.state[4] ),
    .X(net263));
 sg13g2_dlygate4sd3_1 hold237 (.A(_0657_),
    .X(net264));
 sg13g2_dlygate4sd3_1 hold238 (.A(_0026_),
    .X(net265));
 sg13g2_dlygate4sd3_1 hold239 (.A(\bitserial_cipher.state[8] ),
    .X(net266));
 sg13g2_dlygate4sd3_1 hold240 (.A(_0667_),
    .X(net267));
 sg13g2_dlygate4sd3_1 hold241 (.A(_0030_),
    .X(net268));
 sg13g2_dlygate4sd3_1 hold242 (.A(\bitserial_cipher.key[79] ),
    .X(net269));
 sg13g2_dlygate4sd3_1 hold243 (.A(\bitserial_cipher.key[83] ),
    .X(net270));
 sg13g2_dlygate4sd3_1 hold244 (.A(_0141_),
    .X(net271));
 sg13g2_dlygate4sd3_1 hold245 (.A(\bitserial_cipher.key[107] ),
    .X(net272));
 sg13g2_dlygate4sd3_1 hold246 (.A(\bitserial_cipher.key[11] ),
    .X(net273));
 sg13g2_dlygate4sd3_1 hold247 (.A(\bitserial_cipher.state[19] ),
    .X(net274));
 sg13g2_dlygate4sd3_1 hold248 (.A(_0045_),
    .X(net275));
 sg13g2_dlygate4sd3_1 hold249 (.A(\bitserial_cipher.key[126] ),
    .X(net276));
 sg13g2_dlygate4sd3_1 hold250 (.A(\bitserial_cipher.state[59] ),
    .X(net277));
 sg13g2_dlygate4sd3_1 hold251 (.A(_0022_),
    .X(net278));
 sg13g2_dlygate4sd3_1 hold252 (.A(\bitserial_cipher.key[102] ),
    .X(net279));
 sg13g2_dlygate4sd3_1 hold253 (.A(\bitserial_cipher.state[10] ),
    .X(net280));
 sg13g2_dlygate4sd3_1 hold254 (.A(_0671_),
    .X(net281));
 sg13g2_dlygate4sd3_1 hold255 (.A(_0032_),
    .X(net282));
 sg13g2_dlygate4sd3_1 hold256 (.A(\bitserial_cipher.key[125] ),
    .X(net283));
 sg13g2_dlygate4sd3_1 hold257 (.A(_0183_),
    .X(net284));
 sg13g2_dlygate4sd3_1 hold258 (.A(\bitserial_cipher.state[23] ),
    .X(net285));
 sg13g2_dlygate4sd3_1 hold259 (.A(_0682_),
    .X(net286));
 sg13g2_dlygate4sd3_1 hold260 (.A(_0037_),
    .X(net287));
 sg13g2_dlygate4sd3_1 hold261 (.A(\bitserial_cipher.key[124] ),
    .X(net288));
 sg13g2_dlygate4sd3_1 hold262 (.A(\bitserial_cipher.state[33] ),
    .X(net289));
 sg13g2_dlygate4sd3_1 hold263 (.A(_0200_),
    .X(net290));
 sg13g2_dlygate4sd3_1 hold264 (.A(\bitserial_cipher.state[31] ),
    .X(net291));
 sg13g2_dlygate4sd3_1 hold265 (.A(_0198_),
    .X(net292));
 sg13g2_dlygate4sd3_1 hold266 (.A(\bitserial_cipher.state[25] ),
    .X(net293));
 sg13g2_dlygate4sd3_1 hold267 (.A(_0039_),
    .X(net294));
 sg13g2_dlygate4sd3_1 hold268 (.A(\bitserial_cipher.state[26] ),
    .X(net295));
 sg13g2_dlygate4sd3_1 hold269 (.A(_0689_),
    .X(net296));
 sg13g2_dlygate4sd3_1 hold270 (.A(_0040_),
    .X(net297));
 sg13g2_dlygate4sd3_1 hold271 (.A(\bitserial_cipher.state[6] ),
    .X(net298));
 sg13g2_dlygate4sd3_1 hold272 (.A(_0028_),
    .X(net299));
 sg13g2_dlygate4sd3_1 hold273 (.A(\bitserial_cipher.state[17] ),
    .X(net300));
 sg13g2_dlygate4sd3_1 hold274 (.A(\bitserial_cipher.state[21] ),
    .X(net301));
 sg13g2_dlygate4sd3_1 hold275 (.A(_0678_),
    .X(net302));
 sg13g2_dlygate4sd3_1 hold276 (.A(\bitserial_cipher.state[27] ),
    .X(net303));
 sg13g2_dlygate4sd3_1 hold277 (.A(\bitserial_cipher.state[16] ),
    .X(net304));
 sg13g2_dlygate4sd3_1 hold278 (.A(_0685_),
    .X(net305));
 sg13g2_dlygate4sd3_1 hold279 (.A(\bitserial_cipher.key[122] ),
    .X(net306));
 sg13g2_dlygate4sd3_1 hold280 (.A(\bitserial_cipher.state[46] ),
    .X(net307));
 sg13g2_dlygate4sd3_1 hold281 (.A(_0650_),
    .X(net308));
 sg13g2_dlygate4sd3_1 hold282 (.A(_0024_),
    .X(net309));
 sg13g2_dlygate4sd3_1 hold283 (.A(\bitserial_cipher.state[11] ),
    .X(net310));
 sg13g2_dlygate4sd3_1 hold284 (.A(_0673_),
    .X(net311));
 sg13g2_dlygate4sd3_1 hold285 (.A(_0033_),
    .X(net312));
 sg13g2_dlygate4sd3_1 hold286 (.A(\bitserial_cipher.state[3] ),
    .X(net313));
 sg13g2_dlygate4sd3_1 hold287 (.A(_0764_),
    .X(net314));
 sg13g2_dlygate4sd3_1 hold288 (.A(_0049_),
    .X(net315));
 sg13g2_dlygate4sd3_1 hold289 (.A(\bitserial_cipher.state[5] ),
    .X(net316));
 sg13g2_dlygate4sd3_1 hold290 (.A(_0027_),
    .X(net317));
 sg13g2_dlygate4sd3_1 hold291 (.A(\bitserial_cipher.rcount[2] ),
    .X(net318));
 sg13g2_dlygate4sd3_1 hold292 (.A(_0409_),
    .X(net319));
 sg13g2_dlygate4sd3_1 hold293 (.A(_0188_),
    .X(net320));
 sg13g2_dlygate4sd3_1 hold294 (.A(\bitserial_cipher.state[15] ),
    .X(net321));
 sg13g2_dlygate4sd3_1 hold295 (.A(_0694_),
    .X(net322));
 sg13g2_dlygate4sd3_1 hold296 (.A(_0042_),
    .X(net323));
 sg13g2_dlygate4sd3_1 hold297 (.A(\bitserial_cipher.state[2] ),
    .X(net324));
 sg13g2_dlygate4sd3_1 hold298 (.A(_0048_),
    .X(net325));
 sg13g2_dlygate4sd3_1 hold299 (.A(\bitserial_cipher.state[50] ),
    .X(net326));
 sg13g2_dlygate4sd3_1 hold300 (.A(\bitserial_cipher.scount[0] ),
    .X(net327));
 sg13g2_dlygate4sd3_1 hold301 (.A(_0050_),
    .X(net328));
 sg13g2_dlygate4sd3_1 hold302 (.A(\bitserial_cipher.state[18] ),
    .X(net329));
 sg13g2_dlygate4sd3_1 hold303 (.A(_0044_),
    .X(net330));
 sg13g2_dlygate4sd3_1 hold304 (.A(\bitserial_cipher.state[1] ),
    .X(net331));
 sg13g2_dlygate4sd3_1 hold305 (.A(_0047_),
    .X(net332));
 sg13g2_dlygate4sd3_1 hold306 (.A(\bitserial_cipher.state[9] ),
    .X(net333));
 sg13g2_dlygate4sd3_1 hold307 (.A(\bitserial_cipher.state[7] ),
    .X(net334));
 sg13g2_dlygate4sd3_1 hold308 (.A(\bitserial_cipher.state[22] ),
    .X(net335));
 sg13g2_dlygate4sd3_1 hold309 (.A(_0680_),
    .X(net336));
 sg13g2_dlygate4sd3_1 hold310 (.A(\bitserial_cipher.state[45] ),
    .X(net337));
 sg13g2_dlygate4sd3_1 hold311 (.A(_0648_),
    .X(net338));
 sg13g2_dlygate4sd3_1 hold312 (.A(_0023_),
    .X(net339));
 sg13g2_dlygate4sd3_1 hold313 (.A(\bitserial_cipher.dataq ),
    .X(net340));
 sg13g2_dlygate4sd3_1 hold314 (.A(\bitserial_cipher.state[43] ),
    .X(net341));
 sg13g2_dlygate4sd3_1 hold315 (.A(\bitserial_cipher.state[30] ),
    .X(net342));
 sg13g2_dlygate4sd3_1 hold316 (.A(\bitserial_cipher.rcount[0] ),
    .X(net343));
 sg13g2_dlygate4sd3_1 hold317 (.A(\bitserial_cipher.state[13] ),
    .X(net344));
 sg13g2_dlygate4sd3_1 hold318 (.A(\bitserial_cipher.state[44] ),
    .X(net345));
 sg13g2_dlygate4sd3_1 hold319 (.A(\bitserial_cipher.bcount[3] ),
    .X(net346));
 sg13g2_dlygate4sd3_1 hold320 (.A(_0057_),
    .X(net347));
 sg13g2_dlygate4sd3_1 hold321 (.A(\bitserial_cipher.bcount[1] ),
    .X(net348));
 sg13g2_dlygate4sd3_1 hold322 (.A(\bitserial_cipher.state[12] ),
    .X(net349));
 sg13g2_dlygate4sd3_1 hold323 (.A(_0008_),
    .X(net350));
 sg13g2_dlygate4sd3_1 hold324 (.A(\bitserial_cipher.state[40] ),
    .X(net351));
 sg13g2_dlygate4sd3_1 hold325 (.A(\bitserial_cipher.state[14] ),
    .X(net352));
 sg13g2_dlygate4sd3_1 hold326 (.A(_0619_),
    .X(net353));
 sg13g2_dlygate4sd3_1 hold327 (.A(\bitserial_cipher.bcount[2] ),
    .X(net354));
 sg13g2_dlygate4sd3_1 hold328 (.A(\bitserial_cipher.state[10] ),
    .X(net355));
 sg13g2_dlygate4sd3_1 hold329 (.A(\bitserial_cipher.state[29] ),
    .X(net356));
 sg13g2_dlygate4sd3_1 hold330 (.A(_0013_),
    .X(net357));
 sg13g2_dlygate4sd3_1 hold331 (.A(\bitserial_cipher.state[28] ),
    .X(net358));
 sg13g2_dlygate4sd3_1 hold332 (.A(_0623_),
    .X(net359));
 sg13g2_dlygate4sd3_1 hold333 (.A(\bitserial_cipher.scount[2] ),
    .X(net360));
 sg13g2_dlygate4sd3_1 hold334 (.A(\bitserial_cipher.bcount[0] ),
    .X(net361));
 sg13g2_dlygate4sd3_1 hold335 (.A(\bitserial_cipher.bcount[3] ),
    .X(net362));
 sg13g2_dlygate4sd3_1 hold336 (.A(_0514_),
    .X(net363));
 sg13g2_dlygate4sd3_1 hold337 (.A(_0521_),
    .X(net364));
 sg13g2_dlygate4sd3_1 hold338 (.A(\bitserial_cipher.state[4] ),
    .X(net365));
 sg13g2_dlygate4sd3_1 hold339 (.A(\bitserial_cipher.state[44] ),
    .X(net366));
 sg13g2_dlygate4sd3_1 hold340 (.A(\bitserial_cipher.state[12] ),
    .X(net367));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_4 FILLER_0_21 ();
 sg13g2_fill_1 FILLER_0_25 ();
 sg13g2_fill_1 FILLER_0_30 ();
 sg13g2_fill_1 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_40 ();
 sg13g2_decap_8 FILLER_0_47 ();
 sg13g2_fill_1 FILLER_0_54 ();
 sg13g2_decap_8 FILLER_0_59 ();
 sg13g2_decap_8 FILLER_0_66 ();
 sg13g2_fill_2 FILLER_0_73 ();
 sg13g2_fill_1 FILLER_0_75 ();
 sg13g2_fill_1 FILLER_0_84 ();
 sg13g2_fill_1 FILLER_0_92 ();
 sg13g2_decap_8 FILLER_0_97 ();
 sg13g2_decap_8 FILLER_0_108 ();
 sg13g2_fill_1 FILLER_0_115 ();
 sg13g2_decap_8 FILLER_0_124 ();
 sg13g2_decap_8 FILLER_0_131 ();
 sg13g2_decap_8 FILLER_0_138 ();
 sg13g2_decap_8 FILLER_0_145 ();
 sg13g2_decap_8 FILLER_0_152 ();
 sg13g2_decap_8 FILLER_0_159 ();
 sg13g2_decap_8 FILLER_0_166 ();
 sg13g2_decap_8 FILLER_0_173 ();
 sg13g2_decap_8 FILLER_0_180 ();
 sg13g2_decap_8 FILLER_0_187 ();
 sg13g2_decap_8 FILLER_0_194 ();
 sg13g2_decap_8 FILLER_0_201 ();
 sg13g2_decap_8 FILLER_0_208 ();
 sg13g2_decap_8 FILLER_0_215 ();
 sg13g2_decap_8 FILLER_0_222 ();
 sg13g2_decap_8 FILLER_0_229 ();
 sg13g2_decap_8 FILLER_0_236 ();
 sg13g2_decap_8 FILLER_0_243 ();
 sg13g2_decap_8 FILLER_0_250 ();
 sg13g2_decap_8 FILLER_0_257 ();
 sg13g2_decap_8 FILLER_0_264 ();
 sg13g2_decap_8 FILLER_0_271 ();
 sg13g2_decap_8 FILLER_0_278 ();
 sg13g2_decap_8 FILLER_0_285 ();
 sg13g2_decap_8 FILLER_0_292 ();
 sg13g2_decap_8 FILLER_0_299 ();
 sg13g2_decap_8 FILLER_0_306 ();
 sg13g2_decap_8 FILLER_0_313 ();
 sg13g2_decap_8 FILLER_0_320 ();
 sg13g2_decap_8 FILLER_0_327 ();
 sg13g2_decap_8 FILLER_0_334 ();
 sg13g2_decap_8 FILLER_0_341 ();
 sg13g2_decap_8 FILLER_0_348 ();
 sg13g2_fill_2 FILLER_0_355 ();
 sg13g2_fill_1 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_366 ();
 sg13g2_decap_8 FILLER_0_373 ();
 sg13g2_decap_8 FILLER_0_380 ();
 sg13g2_decap_8 FILLER_0_387 ();
 sg13g2_decap_8 FILLER_0_394 ();
 sg13g2_decap_8 FILLER_0_401 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_fill_1 FILLER_1_21 ();
 sg13g2_fill_1 FILLER_1_30 ();
 sg13g2_fill_2 FILLER_1_43 ();
 sg13g2_fill_1 FILLER_1_49 ();
 sg13g2_fill_2 FILLER_1_55 ();
 sg13g2_fill_2 FILLER_1_110 ();
 sg13g2_fill_2 FILLER_1_117 ();
 sg13g2_fill_1 FILLER_1_119 ();
 sg13g2_fill_2 FILLER_1_132 ();
 sg13g2_fill_1 FILLER_1_134 ();
 sg13g2_fill_1 FILLER_1_139 ();
 sg13g2_fill_1 FILLER_1_144 ();
 sg13g2_fill_2 FILLER_1_170 ();
 sg13g2_fill_1 FILLER_1_172 ();
 sg13g2_fill_2 FILLER_1_177 ();
 sg13g2_fill_1 FILLER_1_179 ();
 sg13g2_decap_8 FILLER_1_184 ();
 sg13g2_decap_8 FILLER_1_191 ();
 sg13g2_decap_8 FILLER_1_198 ();
 sg13g2_decap_8 FILLER_1_205 ();
 sg13g2_decap_8 FILLER_1_212 ();
 sg13g2_decap_8 FILLER_1_219 ();
 sg13g2_decap_8 FILLER_1_226 ();
 sg13g2_decap_8 FILLER_1_233 ();
 sg13g2_decap_4 FILLER_1_240 ();
 sg13g2_fill_2 FILLER_1_244 ();
 sg13g2_decap_8 FILLER_1_250 ();
 sg13g2_decap_8 FILLER_1_257 ();
 sg13g2_decap_8 FILLER_1_264 ();
 sg13g2_decap_8 FILLER_1_271 ();
 sg13g2_decap_8 FILLER_1_278 ();
 sg13g2_decap_8 FILLER_1_285 ();
 sg13g2_decap_8 FILLER_1_292 ();
 sg13g2_decap_8 FILLER_1_299 ();
 sg13g2_fill_2 FILLER_1_310 ();
 sg13g2_decap_8 FILLER_1_320 ();
 sg13g2_decap_8 FILLER_1_327 ();
 sg13g2_decap_8 FILLER_1_334 ();
 sg13g2_decap_4 FILLER_1_341 ();
 sg13g2_fill_1 FILLER_1_345 ();
 sg13g2_fill_2 FILLER_1_354 ();
 sg13g2_fill_1 FILLER_1_356 ();
 sg13g2_fill_1 FILLER_1_365 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_fill_2 FILLER_2_7 ();
 sg13g2_decap_4 FILLER_2_13 ();
 sg13g2_fill_1 FILLER_2_17 ();
 sg13g2_fill_1 FILLER_2_44 ();
 sg13g2_fill_2 FILLER_2_50 ();
 sg13g2_fill_2 FILLER_2_87 ();
 sg13g2_fill_1 FILLER_2_115 ();
 sg13g2_fill_2 FILLER_2_186 ();
 sg13g2_fill_2 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_207 ();
 sg13g2_decap_4 FILLER_2_214 ();
 sg13g2_fill_2 FILLER_2_218 ();
 sg13g2_fill_2 FILLER_2_234 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_4 FILLER_2_273 ();
 sg13g2_decap_4 FILLER_2_281 ();
 sg13g2_fill_2 FILLER_2_293 ();
 sg13g2_fill_2 FILLER_2_308 ();
 sg13g2_fill_1 FILLER_2_310 ();
 sg13g2_fill_2 FILLER_2_329 ();
 sg13g2_fill_2 FILLER_2_335 ();
 sg13g2_fill_1 FILLER_2_337 ();
 sg13g2_fill_2 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_387 ();
 sg13g2_decap_8 FILLER_2_394 ();
 sg13g2_decap_8 FILLER_2_401 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_fill_1 FILLER_3_49 ();
 sg13g2_fill_2 FILLER_3_99 ();
 sg13g2_fill_2 FILLER_3_148 ();
 sg13g2_fill_1 FILLER_3_150 ();
 sg13g2_fill_2 FILLER_3_259 ();
 sg13g2_fill_1 FILLER_3_361 ();
 sg13g2_decap_8 FILLER_3_398 ();
 sg13g2_decap_4 FILLER_3_405 ();
 sg13g2_fill_2 FILLER_4_0 ();
 sg13g2_fill_2 FILLER_4_15 ();
 sg13g2_fill_1 FILLER_4_33 ();
 sg13g2_fill_1 FILLER_4_121 ();
 sg13g2_fill_2 FILLER_4_184 ();
 sg13g2_fill_1 FILLER_4_213 ();
 sg13g2_fill_2 FILLER_4_231 ();
 sg13g2_fill_2 FILLER_4_263 ();
 sg13g2_fill_2 FILLER_4_270 ();
 sg13g2_fill_1 FILLER_4_298 ();
 sg13g2_fill_2 FILLER_4_317 ();
 sg13g2_fill_1 FILLER_4_319 ();
 sg13g2_fill_1 FILLER_4_329 ();
 sg13g2_fill_2 FILLER_4_357 ();
 sg13g2_fill_2 FILLER_4_368 ();
 sg13g2_decap_4 FILLER_4_404 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_fill_1 FILLER_5_39 ();
 sg13g2_fill_1 FILLER_5_82 ();
 sg13g2_fill_1 FILLER_5_118 ();
 sg13g2_fill_1 FILLER_5_160 ();
 sg13g2_fill_2 FILLER_5_201 ();
 sg13g2_fill_2 FILLER_5_229 ();
 sg13g2_fill_1 FILLER_5_235 ();
 sg13g2_fill_2 FILLER_5_301 ();
 sg13g2_fill_1 FILLER_5_303 ();
 sg13g2_fill_1 FILLER_5_330 ();
 sg13g2_fill_2 FILLER_5_344 ();
 sg13g2_fill_2 FILLER_5_407 ();
 sg13g2_decap_4 FILLER_6_0 ();
 sg13g2_fill_1 FILLER_6_39 ();
 sg13g2_fill_1 FILLER_6_54 ();
 sg13g2_fill_2 FILLER_6_64 ();
 sg13g2_fill_2 FILLER_6_105 ();
 sg13g2_fill_2 FILLER_6_130 ();
 sg13g2_fill_1 FILLER_6_159 ();
 sg13g2_fill_2 FILLER_6_173 ();
 sg13g2_fill_2 FILLER_6_184 ();
 sg13g2_fill_1 FILLER_6_186 ();
 sg13g2_fill_2 FILLER_6_196 ();
 sg13g2_fill_1 FILLER_6_198 ();
 sg13g2_fill_2 FILLER_6_221 ();
 sg13g2_fill_2 FILLER_6_231 ();
 sg13g2_fill_1 FILLER_6_233 ();
 sg13g2_fill_1 FILLER_6_340 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_fill_2 FILLER_7_0 ();
 sg13g2_fill_2 FILLER_7_37 ();
 sg13g2_fill_1 FILLER_7_124 ();
 sg13g2_fill_1 FILLER_7_168 ();
 sg13g2_fill_2 FILLER_7_195 ();
 sg13g2_fill_1 FILLER_7_246 ();
 sg13g2_fill_2 FILLER_7_270 ();
 sg13g2_fill_1 FILLER_7_272 ();
 sg13g2_fill_1 FILLER_7_309 ();
 sg13g2_fill_1 FILLER_8_145 ();
 sg13g2_fill_1 FILLER_8_187 ();
 sg13g2_fill_2 FILLER_8_206 ();
 sg13g2_fill_1 FILLER_8_217 ();
 sg13g2_fill_1 FILLER_8_249 ();
 sg13g2_fill_2 FILLER_8_328 ();
 sg13g2_fill_1 FILLER_8_335 ();
 sg13g2_fill_1 FILLER_8_344 ();
 sg13g2_fill_2 FILLER_8_353 ();
 sg13g2_fill_1 FILLER_8_382 ();
 sg13g2_decap_4 FILLER_9_0 ();
 sg13g2_fill_2 FILLER_9_4 ();
 sg13g2_fill_1 FILLER_9_58 ();
 sg13g2_fill_2 FILLER_9_63 ();
 sg13g2_fill_2 FILLER_9_82 ();
 sg13g2_fill_2 FILLER_9_110 ();
 sg13g2_fill_1 FILLER_9_121 ();
 sg13g2_fill_1 FILLER_9_173 ();
 sg13g2_fill_1 FILLER_9_217 ();
 sg13g2_fill_1 FILLER_9_252 ();
 sg13g2_fill_2 FILLER_9_301 ();
 sg13g2_fill_2 FILLER_9_311 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_4 FILLER_10_7 ();
 sg13g2_fill_1 FILLER_10_11 ();
 sg13g2_fill_1 FILLER_10_47 ();
 sg13g2_decap_8 FILLER_10_199 ();
 sg13g2_fill_2 FILLER_10_248 ();
 sg13g2_fill_1 FILLER_10_372 ();
 sg13g2_fill_1 FILLER_10_382 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_4 FILLER_11_7 ();
 sg13g2_fill_1 FILLER_11_11 ();
 sg13g2_fill_2 FILLER_11_43 ();
 sg13g2_fill_1 FILLER_11_61 ();
 sg13g2_fill_2 FILLER_11_120 ();
 sg13g2_fill_1 FILLER_11_174 ();
 sg13g2_decap_8 FILLER_11_205 ();
 sg13g2_fill_1 FILLER_11_212 ();
 sg13g2_decap_8 FILLER_11_216 ();
 sg13g2_fill_2 FILLER_11_223 ();
 sg13g2_fill_1 FILLER_11_225 ();
 sg13g2_fill_1 FILLER_11_232 ();
 sg13g2_fill_2 FILLER_11_306 ();
 sg13g2_fill_1 FILLER_11_313 ();
 sg13g2_fill_1 FILLER_11_335 ();
 sg13g2_fill_2 FILLER_11_341 ();
 sg13g2_fill_2 FILLER_11_348 ();
 sg13g2_fill_1 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_4 FILLER_12_14 ();
 sg13g2_fill_2 FILLER_12_35 ();
 sg13g2_fill_1 FILLER_12_37 ();
 sg13g2_fill_2 FILLER_12_102 ();
 sg13g2_fill_1 FILLER_12_109 ();
 sg13g2_fill_2 FILLER_12_261 ();
 sg13g2_fill_2 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_4 FILLER_13_7 ();
 sg13g2_fill_2 FILLER_13_11 ();
 sg13g2_fill_1 FILLER_13_39 ();
 sg13g2_fill_2 FILLER_13_112 ();
 sg13g2_fill_1 FILLER_13_145 ();
 sg13g2_fill_2 FILLER_13_163 ();
 sg13g2_fill_1 FILLER_13_207 ();
 sg13g2_fill_2 FILLER_13_234 ();
 sg13g2_fill_2 FILLER_13_281 ();
 sg13g2_fill_2 FILLER_13_292 ();
 sg13g2_fill_1 FILLER_13_294 ();
 sg13g2_fill_2 FILLER_13_300 ();
 sg13g2_fill_1 FILLER_13_302 ();
 sg13g2_fill_1 FILLER_13_313 ();
 sg13g2_fill_2 FILLER_13_352 ();
 sg13g2_fill_2 FILLER_13_367 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_4 FILLER_14_7 ();
 sg13g2_fill_2 FILLER_14_37 ();
 sg13g2_fill_1 FILLER_14_39 ();
 sg13g2_fill_1 FILLER_14_79 ();
 sg13g2_fill_1 FILLER_14_167 ();
 sg13g2_fill_1 FILLER_14_244 ();
 sg13g2_fill_2 FILLER_14_269 ();
 sg13g2_fill_1 FILLER_14_271 ();
 sg13g2_fill_2 FILLER_14_298 ();
 sg13g2_fill_1 FILLER_14_300 ();
 sg13g2_fill_2 FILLER_14_306 ();
 sg13g2_fill_1 FILLER_14_330 ();
 sg13g2_fill_2 FILLER_14_339 ();
 sg13g2_fill_2 FILLER_14_381 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_4 FILLER_15_14 ();
 sg13g2_fill_1 FILLER_15_18 ();
 sg13g2_fill_2 FILLER_15_74 ();
 sg13g2_fill_1 FILLER_15_84 ();
 sg13g2_fill_1 FILLER_15_118 ();
 sg13g2_fill_1 FILLER_15_128 ();
 sg13g2_fill_2 FILLER_15_147 ();
 sg13g2_fill_1 FILLER_15_176 ();
 sg13g2_fill_1 FILLER_15_201 ();
 sg13g2_fill_2 FILLER_15_220 ();
 sg13g2_fill_2 FILLER_15_226 ();
 sg13g2_fill_1 FILLER_15_233 ();
 sg13g2_fill_2 FILLER_15_240 ();
 sg13g2_fill_1 FILLER_15_242 ();
 sg13g2_fill_1 FILLER_15_248 ();
 sg13g2_fill_2 FILLER_15_268 ();
 sg13g2_fill_1 FILLER_15_270 ();
 sg13g2_fill_2 FILLER_15_288 ();
 sg13g2_fill_1 FILLER_15_290 ();
 sg13g2_fill_1 FILLER_15_296 ();
 sg13g2_fill_1 FILLER_15_305 ();
 sg13g2_fill_1 FILLER_15_390 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_fill_2 FILLER_16_14 ();
 sg13g2_fill_2 FILLER_16_75 ();
 sg13g2_fill_2 FILLER_16_134 ();
 sg13g2_fill_1 FILLER_16_136 ();
 sg13g2_fill_1 FILLER_16_172 ();
 sg13g2_fill_1 FILLER_16_190 ();
 sg13g2_fill_2 FILLER_16_222 ();
 sg13g2_fill_2 FILLER_16_259 ();
 sg13g2_fill_1 FILLER_16_261 ();
 sg13g2_fill_2 FILLER_16_292 ();
 sg13g2_fill_1 FILLER_16_294 ();
 sg13g2_fill_1 FILLER_16_300 ();
 sg13g2_fill_2 FILLER_16_306 ();
 sg13g2_fill_2 FILLER_16_381 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_fill_2 FILLER_17_28 ();
 sg13g2_fill_2 FILLER_17_56 ();
 sg13g2_fill_1 FILLER_17_58 ();
 sg13g2_fill_1 FILLER_17_115 ();
 sg13g2_fill_1 FILLER_17_130 ();
 sg13g2_fill_2 FILLER_17_162 ();
 sg13g2_fill_1 FILLER_17_164 ();
 sg13g2_fill_2 FILLER_17_234 ();
 sg13g2_fill_1 FILLER_17_295 ();
 sg13g2_fill_2 FILLER_17_383 ();
 sg13g2_fill_2 FILLER_17_407 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_4 FILLER_18_42 ();
 sg13g2_fill_2 FILLER_18_46 ();
 sg13g2_fill_2 FILLER_18_61 ();
 sg13g2_fill_1 FILLER_18_68 ();
 sg13g2_fill_2 FILLER_18_108 ();
 sg13g2_fill_2 FILLER_18_136 ();
 sg13g2_fill_1 FILLER_18_138 ();
 sg13g2_fill_1 FILLER_18_174 ();
 sg13g2_fill_1 FILLER_18_193 ();
 sg13g2_fill_2 FILLER_18_214 ();
 sg13g2_fill_2 FILLER_18_277 ();
 sg13g2_fill_2 FILLER_18_328 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_fill_2 FILLER_19_28 ();
 sg13g2_fill_1 FILLER_19_30 ();
 sg13g2_fill_1 FILLER_19_76 ();
 sg13g2_fill_2 FILLER_19_113 ();
 sg13g2_fill_2 FILLER_19_123 ();
 sg13g2_fill_1 FILLER_19_129 ();
 sg13g2_fill_1 FILLER_19_195 ();
 sg13g2_fill_2 FILLER_19_247 ();
 sg13g2_fill_2 FILLER_19_262 ();
 sg13g2_fill_2 FILLER_19_273 ();
 sg13g2_fill_1 FILLER_19_275 ();
 sg13g2_fill_2 FILLER_19_298 ();
 sg13g2_fill_2 FILLER_19_375 ();
 sg13g2_fill_1 FILLER_19_385 ();
 sg13g2_fill_2 FILLER_19_407 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_fill_1 FILLER_20_21 ();
 sg13g2_fill_2 FILLER_20_41 ();
 sg13g2_fill_1 FILLER_20_80 ();
 sg13g2_fill_1 FILLER_20_107 ();
 sg13g2_fill_2 FILLER_20_141 ();
 sg13g2_fill_2 FILLER_20_188 ();
 sg13g2_fill_1 FILLER_20_221 ();
 sg13g2_fill_2 FILLER_20_248 ();
 sg13g2_fill_1 FILLER_20_333 ();
 sg13g2_fill_1 FILLER_20_338 ();
 sg13g2_fill_2 FILLER_20_352 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_fill_1 FILLER_21_14 ();
 sg13g2_fill_2 FILLER_21_136 ();
 sg13g2_fill_2 FILLER_21_148 ();
 sg13g2_fill_1 FILLER_21_150 ();
 sg13g2_fill_1 FILLER_21_160 ();
 sg13g2_fill_2 FILLER_21_300 ();
 sg13g2_fill_2 FILLER_21_316 ();
 sg13g2_fill_1 FILLER_21_366 ();
 sg13g2_fill_1 FILLER_21_394 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_fill_2 FILLER_22_0 ();
 sg13g2_fill_1 FILLER_22_2 ();
 sg13g2_fill_1 FILLER_22_38 ();
 sg13g2_fill_1 FILLER_22_57 ();
 sg13g2_fill_2 FILLER_22_64 ();
 sg13g2_fill_1 FILLER_22_90 ();
 sg13g2_fill_1 FILLER_22_132 ();
 sg13g2_fill_2 FILLER_22_168 ();
 sg13g2_fill_1 FILLER_22_170 ();
 sg13g2_fill_2 FILLER_22_180 ();
 sg13g2_fill_2 FILLER_22_200 ();
 sg13g2_fill_1 FILLER_22_202 ();
 sg13g2_fill_2 FILLER_22_238 ();
 sg13g2_fill_1 FILLER_22_263 ();
 sg13g2_fill_1 FILLER_22_281 ();
 sg13g2_fill_1 FILLER_22_351 ();
 sg13g2_fill_2 FILLER_22_366 ();
 sg13g2_fill_1 FILLER_22_382 ();
 sg13g2_fill_2 FILLER_23_0 ();
 sg13g2_fill_1 FILLER_23_2 ();
 sg13g2_fill_1 FILLER_23_62 ();
 sg13g2_fill_1 FILLER_23_79 ();
 sg13g2_fill_2 FILLER_23_91 ();
 sg13g2_fill_2 FILLER_23_116 ();
 sg13g2_fill_2 FILLER_23_149 ();
 sg13g2_fill_1 FILLER_23_151 ();
 sg13g2_fill_2 FILLER_23_211 ();
 sg13g2_fill_1 FILLER_23_213 ();
 sg13g2_fill_1 FILLER_23_235 ();
 sg13g2_fill_1 FILLER_23_284 ();
 sg13g2_fill_2 FILLER_23_303 ();
 sg13g2_fill_1 FILLER_23_318 ();
 sg13g2_fill_1 FILLER_23_335 ();
 sg13g2_fill_2 FILLER_23_380 ();
 sg13g2_fill_1 FILLER_23_408 ();
 sg13g2_fill_2 FILLER_24_0 ();
 sg13g2_fill_1 FILLER_24_28 ();
 sg13g2_fill_2 FILLER_24_64 ();
 sg13g2_fill_2 FILLER_24_140 ();
 sg13g2_fill_1 FILLER_24_142 ();
 sg13g2_fill_2 FILLER_24_192 ();
 sg13g2_fill_1 FILLER_24_194 ();
 sg13g2_fill_2 FILLER_24_227 ();
 sg13g2_fill_1 FILLER_24_238 ();
 sg13g2_fill_2 FILLER_24_329 ();
 sg13g2_fill_1 FILLER_24_363 ();
 sg13g2_fill_1 FILLER_24_378 ();
 sg13g2_fill_2 FILLER_25_69 ();
 sg13g2_fill_1 FILLER_25_71 ();
 sg13g2_fill_2 FILLER_25_143 ();
 sg13g2_fill_1 FILLER_25_145 ();
 sg13g2_fill_2 FILLER_25_160 ();
 sg13g2_fill_2 FILLER_25_196 ();
 sg13g2_fill_1 FILLER_25_244 ();
 sg13g2_fill_1 FILLER_25_303 ();
 sg13g2_fill_2 FILLER_25_407 ();
 sg13g2_fill_2 FILLER_26_0 ();
 sg13g2_fill_1 FILLER_26_42 ();
 sg13g2_fill_1 FILLER_26_125 ();
 sg13g2_fill_2 FILLER_26_164 ();
 sg13g2_fill_2 FILLER_26_301 ();
 sg13g2_fill_2 FILLER_26_329 ();
 sg13g2_fill_1 FILLER_26_340 ();
 sg13g2_fill_2 FILLER_26_380 ();
 sg13g2_fill_2 FILLER_26_407 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_fill_2 FILLER_27_7 ();
 sg13g2_fill_1 FILLER_27_26 ();
 sg13g2_fill_1 FILLER_27_36 ();
 sg13g2_fill_2 FILLER_27_72 ();
 sg13g2_fill_1 FILLER_27_74 ();
 sg13g2_fill_2 FILLER_27_140 ();
 sg13g2_fill_1 FILLER_27_292 ();
 sg13g2_fill_1 FILLER_27_298 ();
 sg13g2_fill_1 FILLER_27_307 ();
 sg13g2_fill_1 FILLER_27_373 ();
 sg13g2_fill_2 FILLER_28_0 ();
 sg13g2_fill_1 FILLER_28_2 ();
 sg13g2_fill_1 FILLER_28_51 ();
 sg13g2_fill_1 FILLER_28_66 ();
 sg13g2_fill_1 FILLER_28_92 ();
 sg13g2_fill_1 FILLER_28_102 ();
 sg13g2_fill_1 FILLER_28_117 ();
 sg13g2_fill_1 FILLER_28_142 ();
 sg13g2_fill_1 FILLER_28_151 ();
 sg13g2_fill_2 FILLER_28_168 ();
 sg13g2_fill_1 FILLER_28_170 ();
 sg13g2_fill_2 FILLER_28_192 ();
 sg13g2_fill_1 FILLER_28_248 ();
 sg13g2_fill_2 FILLER_28_300 ();
 sg13g2_fill_2 FILLER_28_313 ();
 sg13g2_fill_2 FILLER_28_407 ();
 sg13g2_fill_1 FILLER_29_92 ();
 sg13g2_fill_2 FILLER_29_133 ();
 sg13g2_fill_2 FILLER_29_143 ();
 sg13g2_fill_2 FILLER_29_166 ();
 sg13g2_fill_2 FILLER_29_207 ();
 sg13g2_fill_1 FILLER_29_261 ();
 sg13g2_fill_1 FILLER_29_267 ();
 sg13g2_fill_1 FILLER_29_290 ();
 sg13g2_fill_1 FILLER_29_296 ();
 sg13g2_fill_1 FILLER_29_305 ();
 sg13g2_fill_2 FILLER_29_330 ();
 sg13g2_fill_2 FILLER_29_407 ();
 sg13g2_fill_2 FILLER_30_0 ();
 sg13g2_fill_1 FILLER_30_28 ();
 sg13g2_fill_1 FILLER_30_50 ();
 sg13g2_fill_1 FILLER_30_94 ();
 sg13g2_fill_1 FILLER_30_137 ();
 sg13g2_fill_2 FILLER_30_193 ();
 sg13g2_fill_1 FILLER_30_195 ();
 sg13g2_fill_2 FILLER_30_273 ();
 sg13g2_fill_2 FILLER_30_279 ();
 sg13g2_fill_2 FILLER_30_289 ();
 sg13g2_fill_1 FILLER_30_296 ();
 sg13g2_fill_1 FILLER_30_315 ();
 sg13g2_fill_2 FILLER_31_30 ();
 sg13g2_fill_1 FILLER_31_71 ();
 sg13g2_fill_2 FILLER_31_92 ();
 sg13g2_fill_1 FILLER_31_94 ();
 sg13g2_fill_2 FILLER_31_117 ();
 sg13g2_fill_2 FILLER_31_165 ();
 sg13g2_fill_1 FILLER_31_167 ();
 sg13g2_fill_1 FILLER_31_200 ();
 sg13g2_fill_2 FILLER_31_240 ();
 sg13g2_fill_1 FILLER_31_266 ();
 sg13g2_fill_1 FILLER_31_292 ();
 sg13g2_fill_2 FILLER_31_314 ();
 sg13g2_fill_2 FILLER_31_342 ();
 sg13g2_fill_1 FILLER_32_0 ();
 sg13g2_fill_2 FILLER_32_35 ();
 sg13g2_fill_2 FILLER_32_65 ();
 sg13g2_fill_2 FILLER_32_102 ();
 sg13g2_fill_1 FILLER_32_140 ();
 sg13g2_fill_1 FILLER_32_312 ();
 sg13g2_fill_1 FILLER_32_319 ();
 sg13g2_fill_1 FILLER_33_26 ();
 sg13g2_fill_2 FILLER_33_36 ();
 sg13g2_fill_2 FILLER_33_95 ();
 sg13g2_fill_1 FILLER_33_133 ();
 sg13g2_fill_2 FILLER_33_242 ();
 sg13g2_fill_2 FILLER_33_264 ();
 sg13g2_fill_2 FILLER_33_318 ();
 sg13g2_fill_2 FILLER_33_325 ();
 sg13g2_fill_1 FILLER_33_376 ();
 sg13g2_fill_1 FILLER_33_408 ();
 sg13g2_fill_2 FILLER_34_0 ();
 sg13g2_fill_1 FILLER_34_2 ();
 sg13g2_fill_1 FILLER_34_29 ();
 sg13g2_fill_2 FILLER_34_72 ();
 sg13g2_fill_1 FILLER_34_84 ();
 sg13g2_fill_2 FILLER_34_130 ();
 sg13g2_fill_1 FILLER_34_164 ();
 sg13g2_fill_2 FILLER_34_265 ();
 sg13g2_fill_1 FILLER_34_313 ();
 sg13g2_fill_1 FILLER_34_399 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_fill_2 FILLER_35_7 ();
 sg13g2_fill_1 FILLER_35_9 ();
 sg13g2_fill_1 FILLER_35_28 ();
 sg13g2_fill_1 FILLER_35_73 ();
 sg13g2_fill_2 FILLER_35_159 ();
 sg13g2_fill_1 FILLER_35_337 ();
 sg13g2_fill_1 FILLER_35_373 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_4 FILLER_36_14 ();
 sg13g2_fill_1 FILLER_36_135 ();
 sg13g2_fill_2 FILLER_36_152 ();
 sg13g2_fill_1 FILLER_36_197 ();
 sg13g2_fill_1 FILLER_36_253 ();
 sg13g2_fill_1 FILLER_36_322 ();
 sg13g2_fill_1 FILLER_36_328 ();
 sg13g2_fill_1 FILLER_36_338 ();
 sg13g2_fill_2 FILLER_36_347 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_4 FILLER_37_21 ();
 sg13g2_fill_1 FILLER_37_25 ();
 sg13g2_fill_1 FILLER_37_29 ();
 sg13g2_fill_2 FILLER_37_40 ();
 sg13g2_fill_2 FILLER_37_69 ();
 sg13g2_fill_2 FILLER_37_81 ();
 sg13g2_fill_2 FILLER_37_172 ();
 sg13g2_fill_2 FILLER_37_237 ();
 sg13g2_fill_2 FILLER_37_319 ();
 sg13g2_fill_1 FILLER_37_408 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_4 FILLER_38_28 ();
 sg13g2_fill_1 FILLER_38_32 ();
 sg13g2_fill_2 FILLER_38_220 ();
 sg13g2_fill_2 FILLER_38_252 ();
 sg13g2_fill_2 FILLER_38_287 ();
 sg13g2_fill_1 FILLER_38_328 ();
 assign uio_oe[0] = net6;
 assign uio_oe[1] = net7;
 assign uio_oe[2] = net8;
 assign uio_oe[3] = net9;
 assign uio_oe[4] = net10;
 assign uio_oe[5] = net11;
 assign uio_oe[6] = net12;
 assign uio_oe[7] = net13;
 assign uio_out[0] = net14;
 assign uio_out[1] = net15;
 assign uio_out[2] = net16;
 assign uio_out[3] = net17;
 assign uio_out[4] = net18;
 assign uio_out[5] = net19;
 assign uio_out[6] = net20;
 assign uio_out[7] = net21;
 assign uo_out[2] = net22;
 assign uo_out[3] = net23;
 assign uo_out[4] = net24;
 assign uo_out[5] = net25;
 assign uo_out[6] = net26;
 assign uo_out[7] = net27;
endmodule

module tt_um_cejmu (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire \bav0._02_ ;
 wire \bav0.state_q[0] ;
 wire \bav0.state_q[1] ;
 wire \bav0.state_q[2] ;
 wire \bav1._02_ ;
 wire \bav1.state_q[0] ;
 wire \bav1.state_q[1] ;
 wire \bav1.state_q[2] ;
 wire \bav1.x[0] ;
 wire \bav1.x[1] ;
 wire \ca._07_[0] ;
 wire \ca._08_[0] ;
 wire \ca._11_ ;
 wire \ca._13_ ;
 wire \ca._15_ ;
 wire \ca.coin_out[2] ;
 wire \ca.coin_out[3] ;
 wire \ca.coin_out[4] ;
 wire \ca.coin_out[5] ;
 wire \ca.commit_count[0] ;
 wire \ca.commit_count[10] ;
 wire \ca.commit_count[11] ;
 wire \ca.commit_count[12] ;
 wire \ca.commit_count[13] ;
 wire \ca.commit_count[14] ;
 wire \ca.commit_count[15] ;
 wire \ca.commit_count[16] ;
 wire \ca.commit_count[17] ;
 wire \ca.commit_count[18] ;
 wire \ca.commit_count[19] ;
 wire \ca.commit_count[1] ;
 wire \ca.commit_count[20] ;
 wire \ca.commit_count[21] ;
 wire \ca.commit_count[2] ;
 wire \ca.commit_count[3] ;
 wire \ca.commit_count[4] ;
 wire \ca.commit_count[5] ;
 wire \ca.commit_count[6] ;
 wire \ca.commit_count[7] ;
 wire \ca.commit_count[8] ;
 wire \ca.commit_count[9] ;
 wire \ca.pulse0 ;
 wire \ca.pulse_count[0] ;
 wire \ca.pulse_count[1] ;
 wire \ca.pulse_count[2] ;
 wire \ca.pulse_count[3] ;
 wire \ca.pulse_count[4] ;
 wire \ca.pulse_count[5] ;
 wire \cla_z[0] ;
 wire \cla_z[10] ;
 wire \cla_z[11] ;
 wire \cla_z[12] ;
 wire \cla_z[13] ;
 wire \cla_z[14] ;
 wire \cla_z[15] ;
 wire \cla_z[16] ;
 wire \cla_z[17] ;
 wire \cla_z[18] ;
 wire \cla_z[19] ;
 wire \cla_z[1] ;
 wire \cla_z[20] ;
 wire \cla_z[21] ;
 wire \cla_z[22] ;
 wire \cla_z[23] ;
 wire \cla_z[2] ;
 wire \cla_z[3] ;
 wire \cla_z[4] ;
 wire \cla_z[5] ;
 wire \cla_z[6] ;
 wire \cla_z[7] ;
 wire \cla_z[8] ;
 wire \cla_z[9] ;
 wire \io_sd._052_[0] ;
 wire \io_sd._052_[10] ;
 wire \io_sd._052_[11] ;
 wire \io_sd._052_[12] ;
 wire \io_sd._052_[13] ;
 wire \io_sd._052_[14] ;
 wire \io_sd._052_[15] ;
 wire \io_sd._052_[16] ;
 wire \io_sd._052_[17] ;
 wire \io_sd._052_[18] ;
 wire \io_sd._052_[19] ;
 wire \io_sd._052_[1] ;
 wire \io_sd._052_[20] ;
 wire \io_sd._052_[21] ;
 wire \io_sd._052_[22] ;
 wire \io_sd._052_[23] ;
 wire \io_sd._052_[2] ;
 wire \io_sd._052_[3] ;
 wire \io_sd._052_[4] ;
 wire \io_sd._052_[5] ;
 wire \io_sd._052_[6] ;
 wire \io_sd._052_[7] ;
 wire \io_sd._052_[8] ;
 wire \io_sd._052_[9] ;
 wire \io_sd._053_[0] ;
 wire \io_sd._053_[10] ;
 wire \io_sd._053_[11] ;
 wire \io_sd._053_[12] ;
 wire \io_sd._053_[13] ;
 wire \io_sd._053_[14] ;
 wire \io_sd._053_[15] ;
 wire \io_sd._053_[16] ;
 wire \io_sd._053_[17] ;
 wire \io_sd._053_[18] ;
 wire \io_sd._053_[19] ;
 wire \io_sd._053_[1] ;
 wire \io_sd._053_[20] ;
 wire \io_sd._053_[21] ;
 wire \io_sd._053_[22] ;
 wire \io_sd._053_[23] ;
 wire \io_sd._053_[2] ;
 wire \io_sd._053_[3] ;
 wire \io_sd._053_[4] ;
 wire \io_sd._053_[5] ;
 wire \io_sd._053_[6] ;
 wire \io_sd._053_[7] ;
 wire \io_sd._053_[8] ;
 wire \io_sd._053_[9] ;
 wire \io_sd._080_ ;
 wire \io_sd._083_ ;
 wire \io_sd._209_[0] ;
 wire \io_sd._210_[0] ;
 wire \io_sd.input_index[3] ;
 wire \io_sd.input_index[4] ;
 wire \io_sd.input_index[5] ;
 wire \io_sd.output_index[3] ;
 wire \io_sd.output_index[4] ;
 wire \io_sd.output_index[5] ;
 wire \io_sd.outputs[0] ;
 wire \io_sd.outputs[1] ;
 wire \io_sd.outputs[2] ;
 wire \io_sd.outputs[3] ;
 wire \io_sd.outputs[4] ;
 wire \io_sd.outputs[5] ;
 wire \io_sd.outputs[6] ;
 wire \io_sd.outputs[7] ;
 wire \rca.generate_adder_modules[0].fa.a ;
 wire \rca.generate_adder_modules[0].fa.b ;
 wire \rca.generate_adder_modules[10].fa.a ;
 wire \rca.generate_adder_modules[10].fa.b ;
 wire \rca.generate_adder_modules[11].fa.a ;
 wire \rca.generate_adder_modules[11].fa.b ;
 wire \rca.generate_adder_modules[12].fa.a ;
 wire \rca.generate_adder_modules[12].fa.b ;
 wire \rca.generate_adder_modules[13].fa.a ;
 wire \rca.generate_adder_modules[13].fa.b ;
 wire \rca.generate_adder_modules[14].fa.a ;
 wire \rca.generate_adder_modules[14].fa.b ;
 wire \rca.generate_adder_modules[15].fa.a ;
 wire \rca.generate_adder_modules[15].fa.b ;
 wire \rca.generate_adder_modules[16].fa.a ;
 wire \rca.generate_adder_modules[16].fa.b ;
 wire \rca.generate_adder_modules[17].fa.a ;
 wire \rca.generate_adder_modules[17].fa.b ;
 wire \rca.generate_adder_modules[18].fa.a ;
 wire \rca.generate_adder_modules[18].fa.b ;
 wire \rca.generate_adder_modules[19].fa.a ;
 wire \rca.generate_adder_modules[19].fa.b ;
 wire \rca.generate_adder_modules[1].fa.a ;
 wire \rca.generate_adder_modules[1].fa.b ;
 wire \rca.generate_adder_modules[20].fa.a ;
 wire \rca.generate_adder_modules[20].fa.b ;
 wire \rca.generate_adder_modules[21].fa.a ;
 wire \rca.generate_adder_modules[21].fa.b ;
 wire \rca.generate_adder_modules[22].fa.a ;
 wire \rca.generate_adder_modules[22].fa.b ;
 wire \rca.generate_adder_modules[23].fa._02_ ;
 wire \rca.generate_adder_modules[23].fa.a ;
 wire \rca.generate_adder_modules[23].fa.b ;
 wire \rca.generate_adder_modules[2].fa.a ;
 wire \rca.generate_adder_modules[2].fa.b ;
 wire \rca.generate_adder_modules[3].fa.a ;
 wire \rca.generate_adder_modules[3].fa.b ;
 wire \rca.generate_adder_modules[4].fa.a ;
 wire \rca.generate_adder_modules[4].fa.b ;
 wire \rca.generate_adder_modules[5].fa.a ;
 wire \rca.generate_adder_modules[5].fa.b ;
 wire \rca.generate_adder_modules[6].fa.a ;
 wire \rca.generate_adder_modules[6].fa.b ;
 wire \rca.generate_adder_modules[7].fa.a ;
 wire \rca.generate_adder_modules[7].fa.b ;
 wire \rca.generate_adder_modules[8].fa.a ;
 wire \rca.generate_adder_modules[8].fa.b ;
 wire \rca.generate_adder_modules[9].fa.a ;
 wire \rca.generate_adder_modules[9].fa.b ;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net138;
 wire clknet_0_clk;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire \cla/_0341_ ;
 wire \cla/_342_ ;
 wire \cla/_343_ ;
 wire \cla/_344_ ;
 wire \cla/_345_ ;
 wire \cla/_346_ ;
 wire \cla/_347_ ;
 wire \cla/_348_ ;
 wire \cla/_349_ ;
 wire \cla/_350_ ;
 wire \cla/_351_ ;
 wire \cla/_352_ ;
 wire \cla/_353_ ;
 wire \cla/_354_ ;
 wire \cla/_355_ ;
 wire \cla/_356_ ;
 wire \cla/_357_ ;
 wire \cla/_358_ ;
 wire \cla/_359_ ;
 wire \cla/_360_ ;
 wire \cla/_361_ ;
 wire \cla/_362_ ;
 wire \cla/_363_ ;
 wire \cla/_364_ ;
 wire \cla/_365_ ;
 wire \cla/_366_ ;
 wire \cla/_367_ ;
 wire \cla/_368_ ;
 wire \cla/_369_ ;
 wire \cla/_370_ ;
 wire \cla/_371_ ;
 wire \cla/_372_ ;
 wire \cla/_373_ ;
 wire \cla/_374_ ;
 wire \cla/_375_ ;
 wire \cla/_376_ ;
 wire \cla/_377_ ;
 wire \cla/_378_ ;
 wire \cla/_379_ ;
 wire \cla/_380_ ;
 wire \cla/_381_ ;
 wire \cla/_382_ ;
 wire \cla/_383_ ;
 wire \cla/_384_ ;
 wire \cla/_385_ ;
 wire \cla/_386_ ;
 wire \cla/_387_ ;
 wire \cla/_388_ ;
 wire \cla/_389_ ;
 wire \cla/_390_ ;
 wire \cla/_391_ ;
 wire \cla/_392_ ;
 wire \cla/_393_ ;
 wire \cla/_394_ ;
 wire \cla/_395_ ;
 wire \cla/_396_ ;
 wire \cla/_397_ ;
 wire \cla/_398_ ;
 wire \cla/_399_ ;
 wire \cla/_400_ ;
 wire \cla/_401_ ;
 wire \cla/_402_ ;
 wire \cla/_403_ ;
 wire \cla/_404_ ;
 wire \cla/_405_ ;
 wire \cla/_406_ ;
 wire \cla/_407_ ;
 wire \cla/_408_ ;
 wire \cla/_409_ ;
 wire \cla/_410_ ;
 wire \cla/_411_ ;
 wire \cla/_412_ ;
 wire \cla/_413_ ;
 wire \cla/_414_ ;
 wire \cla/_415_ ;
 wire \cla/_416_ ;
 wire \cla/_417_ ;
 wire \cla/_418_ ;
 wire \cla/_419_ ;
 wire \cla/_420_ ;
 wire \cla/_421_ ;
 wire \cla/_422_ ;
 wire \cla/_423_ ;
 wire \cla/_424_ ;
 wire \cla/_425_ ;
 wire \cla/_426_ ;
 wire \cla/_427_ ;
 wire \cla/_428_ ;
 wire \cla/_429_ ;
 wire \cla/_430_ ;
 wire \cla/_431_ ;
 wire \cla/_432_ ;
 wire \cla/_433_ ;
 wire \cla/_434_ ;
 wire \cla/_435_ ;
 wire \cla/_436_ ;
 wire \cla/_437_ ;
 wire \cla/_438_ ;
 wire \cla/_439_ ;
 wire \cla/_440_ ;
 wire \cla/_441_ ;
 wire \cla/_442_ ;
 wire \cla/_443_ ;
 wire \cla/_444_ ;
 wire \cla/_445_ ;
 wire \cla/_446_ ;
 wire \cla/_447_ ;
 wire \cla/_448_ ;
 wire \cla/_449_ ;
 wire \cla/_450_ ;
 wire \cla/_451_ ;
 wire \cla/_452_ ;
 wire \cla/_453_ ;
 wire \cla/_454_ ;
 wire \cla/_455_ ;
 wire \cla/_456_ ;
 wire \cla/_457_ ;
 wire \cla/_458_ ;
 wire \cla/_459_ ;
 wire \cla/_460_ ;
 wire \cla/_461_ ;
 wire \cla/_462_ ;
 wire \cla/_463_ ;
 wire \cla/_464_ ;
 wire \cla/_465_ ;
 wire \cla/_466_ ;
 wire \cla/_467_ ;
 wire \cla/_468_ ;
 wire \cla/_469_ ;
 wire \cla/_470_ ;
 wire \cla/_471_ ;
 wire \cla/_472_ ;
 wire \cla/_473_ ;
 wire \cla/_474_ ;
 wire \cla/_475_ ;
 wire \cla/_476_ ;
 wire \cla/_477_ ;
 wire \cla/_478_ ;
 wire \cla/_479_ ;
 wire \cla/_480_ ;
 wire \cla/_481_ ;
 wire \cla/_482_ ;
 wire \cla/_483_ ;
 wire \cla/_484_ ;
 wire \cla/_485_ ;
 wire \cla/_486_ ;
 wire \cla/_487_ ;
 wire \cla/_488_ ;
 wire \cla/_489_ ;
 wire \cla/_490_ ;
 wire \cla/_491_ ;
 wire \cla/_492_ ;
 wire \cla/_493_ ;
 wire \cla/_494_ ;
 wire \cla/_495_ ;
 wire \cla/_496_ ;
 wire \cla/_497_ ;
 wire \cla/_498_ ;
 wire \cla/_499_ ;
 wire \cla/_500_ ;
 wire \cla/_501_ ;
 wire \cla/_502_ ;
 wire \cla/_503_ ;
 wire \cla/_504_ ;
 wire \cla/_505_ ;
 wire \cla/_506_ ;
 wire \cla/_507_ ;
 wire \cla/_508_ ;
 wire \cla/_509_ ;
 wire \cla/_510_ ;
 wire \cla/_511_ ;
 wire \cla/_512_ ;
 wire \cla/_513_ ;
 wire \cla/_514_ ;
 wire \cla/_515_ ;
 wire \cla/_516_ ;
 wire \cla/_517_ ;
 wire \cla/_518_ ;
 wire \cla/_519_ ;
 wire \cla/_520_ ;
 wire \cla/_521_ ;
 wire \cla/_522_ ;
 wire \cla/_523_ ;
 wire \cla/_524_ ;
 wire \cla/_525_ ;
 wire \cla/_526_ ;
 wire \cla/_527_ ;
 wire \cla/_528_ ;
 wire \cla/_529_ ;
 wire \cla/_530_ ;
 wire \cla/_531_ ;
 wire \cla/_532_ ;
 wire \cla/_533_ ;
 wire \cla/_534_ ;
 wire \cla/_535_ ;
 wire \cla/_536_ ;
 wire \cla/_537_ ;
 wire \cla/_538_ ;
 wire \cla/_539_ ;
 wire \cla/_540_ ;
 wire \cla/_541_ ;
 wire \cla/_542_ ;
 wire \cla/_543_ ;
 wire \cla/_544_ ;
 wire \cla/_545_ ;
 wire \cla/_546_ ;
 wire \cla/_547_ ;
 wire \cla/_548_ ;
 wire \cla/_549_ ;
 wire \cla/_550_ ;
 wire \cla/_551_ ;
 wire \cla/_552_ ;
 wire \cla/_553_ ;
 wire \cla/_554_ ;
 wire \cla/_555_ ;
 wire \cla/_556_ ;
 wire \cla/_557_ ;
 wire \cla/_558_ ;
 wire \cla/_559_ ;
 wire \cla/_560_ ;
 wire \cla/_561_ ;
 wire \cla/_562_ ;
 wire \cla/_563_ ;
 wire \cla/_564_ ;
 wire \cla/_565_ ;
 wire \cla/_566_ ;
 wire \cla/_567_ ;
 wire \cla/_568_ ;
 wire \cla/_569_ ;
 wire \cla/_570_ ;
 wire \cla/_571_ ;
 wire \cla/_572_ ;
 wire \cla/_573_ ;
 wire \cla/_574_ ;
 wire \cla/_575_ ;
 wire \cla/_576_ ;
 wire \cla/_577_ ;
 wire \cla/_578_ ;
 wire \cla/_579_ ;
 wire \cla/_580_ ;
 wire \cla/_581_ ;
 wire \cla/_582_ ;
 wire \cla/_583_ ;
 wire \cla/_584_ ;
 wire \cla/_585_ ;
 wire \cla/_586_ ;
 wire \cla/_587_ ;
 wire \cla/_588_ ;
 wire \cla/_589_ ;
 wire \cla/_590_ ;
 wire \cla/generate_adder_modules[0].fa_i._2_ ;
 wire \cla/generate_adder_modules[10].fa_i._3_ ;
 wire \cla/generate_adder_modules[11].fa_i._3_ ;
 wire \cla/generate_adder_modules[12].fa_i._3_ ;
 wire \cla/generate_adder_modules[13].fa_i._3_ ;
 wire \cla/generate_adder_modules[14].fa_i._3_ ;
 wire \cla/generate_adder_modules[15].fa_i._3_ ;
 wire \cla/generate_adder_modules[16].fa_i._3_ ;
 wire \cla/generate_adder_modules[17].fa_i._3_ ;
 wire \cla/generate_adder_modules[18].fa_i._3_ ;
 wire \cla/generate_adder_modules[19].fa_i._3_ ;
 wire \cla/generate_adder_modules[1].fa_i._3_ ;
 wire \cla/generate_adder_modules[20].fa_i._3_ ;
 wire \cla/generate_adder_modules[21].fa_i._3_ ;
 wire \cla/generate_adder_modules[22].fa_i._3_ ;
 wire \cla/generate_adder_modules[23].fa_i._3_ ;
 wire \cla/generate_adder_modules[2].fa_i._3_ ;
 wire \cla/generate_adder_modules[3].fa_i._3_ ;
 wire \cla/generate_adder_modules[4].fa_i._3_ ;
 wire \cla/generate_adder_modules[5].fa_i._3_ ;
 wire \cla/generate_adder_modules[6].fa_i._3_ ;
 wire \cla/generate_adder_modules[7].fa_i._3_ ;
 wire \cla/generate_adder_modules[8].fa_i._3_ ;
 wire \cla/generate_adder_modules[9].fa_i._3_ ;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;

 sg13g2_inv_1 _0863_ (.Y(_0131_),
    .A(net12));
 sg13g2_inv_1 _0864_ (.Y(_0132_),
    .A(\ca.commit_count[19] ));
 sg13g2_inv_1 _0865_ (.Y(_0133_),
    .A(net218));
 sg13g2_inv_2 _0866_ (.Y(_0134_),
    .A(net219));
 sg13g2_inv_2 _0867_ (.Y(_0135_),
    .A(net249));
 sg13g2_inv_1 _0868_ (.Y(_0136_),
    .A(net334));
 sg13g2_inv_1 _0869_ (.Y(_0137_),
    .A(net9));
 sg13g2_nand2_1 _0870_ (.Y(_0138_),
    .A(net12),
    .B(net247));
 sg13g2_nor2_1 _0871_ (.A(net331),
    .B(net220),
    .Y(_0139_));
 sg13g2_nor2_1 _0872_ (.A(net214),
    .B(\io_sd.output_index[5] ),
    .Y(_0140_));
 sg13g2_o21ai_1 _0873_ (.B1(_0139_),
    .Y(_0141_),
    .A1(_0010_),
    .A2(_0140_));
 sg13g2_nor2b_1 _0874_ (.A(_0138_),
    .B_N(_0141_),
    .Y(_0142_));
 sg13g2_nor2_1 _0875_ (.A(net12),
    .B(net235),
    .Y(_0143_));
 sg13g2_nor2b_1 _0876_ (.A(\io_sd.input_index[5] ),
    .B_N(net216),
    .Y(_0144_));
 sg13g2_nor2_1 _0877_ (.A(net328),
    .B(net217),
    .Y(_0145_));
 sg13g2_o21ai_1 _0878_ (.B1(_0145_),
    .Y(_0146_),
    .A1(_0011_),
    .A2(_0144_));
 sg13g2_a21oi_1 _0879_ (.A1(net211),
    .A2(_0146_),
    .Y(_0147_),
    .B1(_0142_));
 sg13g2_o21ai_1 _0880_ (.B1(net1),
    .Y(_0004_),
    .A1(_0136_),
    .A2(_0147_));
 sg13g2_nor2b_2 _0881_ (.A(\bav1.x[0] ),
    .B_N(\bav1.x[1] ),
    .Y(_0148_));
 sg13g2_nor2b_2 _0882_ (.A(net325),
    .B_N(\bav1.x[0] ),
    .Y(_0149_));
 sg13g2_nor2_1 _0883_ (.A(_0148_),
    .B(_0149_),
    .Y(_0150_));
 sg13g2_nand3_1 _0884_ (.B(net251),
    .C(_0150_),
    .A(net248),
    .Y(_0151_));
 sg13g2_nand3_1 _0885_ (.B(net279),
    .C(_0148_),
    .A(net248),
    .Y(_0152_));
 sg13g2_nand3_1 _0886_ (.B(net184),
    .C(_0149_),
    .A(net248),
    .Y(_0153_));
 sg13g2_nand3_1 _0887_ (.B(_0152_),
    .C(_0153_),
    .A(_0151_),
    .Y(_0001_));
 sg13g2_nor2b_1 _0888_ (.A(net3),
    .B_N(net2),
    .Y(_0154_));
 sg13g2_nor2b_2 _0889_ (.A(net2),
    .B_N(net3),
    .Y(_0155_));
 sg13g2_nor2_1 _0890_ (.A(_0154_),
    .B(_0155_),
    .Y(_0156_));
 sg13g2_nor3_1 _0891_ (.A(net237),
    .B(_0154_),
    .C(_0155_),
    .Y(_0157_));
 sg13g2_a21o_1 _0892_ (.A2(_0156_),
    .A1(net182),
    .B1(net237),
    .X(_0006_));
 sg13g2_and2_1 _0893_ (.A(net249),
    .B(_0154_),
    .X(_0158_));
 sg13g2_a22oi_1 _0894_ (.Y(_0159_),
    .B1(_0158_),
    .B2(net182),
    .A2(_0157_),
    .A1(net175));
 sg13g2_inv_1 _0895_ (.Y(_0008_),
    .A(_0159_));
 sg13g2_a21o_1 _0896_ (.A2(_0150_),
    .A1(net279),
    .B1(net231),
    .X(_0000_));
 sg13g2_nand2b_1 _0897_ (.Y(_0160_),
    .B(net262),
    .A_N(_0147_));
 sg13g2_nand2_1 _0898_ (.Y(_0161_),
    .A(\io_sd._083_ ),
    .B(net211));
 sg13g2_o21ai_1 _0899_ (.B1(_0160_),
    .Y(_0005_),
    .A1(_0146_),
    .A2(_0161_));
 sg13g2_nand2b_1 _0900_ (.Y(_0056_),
    .B(net1),
    .A_N(net2));
 sg13g2_nand3_1 _0901_ (.B(\bav0.state_q[0] ),
    .C(_0155_),
    .A(net249),
    .Y(_0162_));
 sg13g2_a22oi_1 _0902_ (.Y(_0163_),
    .B1(_0158_),
    .B2(net175),
    .A2(_0157_),
    .A1(net167));
 sg13g2_nand2_1 _0903_ (.Y(_0007_),
    .A(_0162_),
    .B(_0163_));
 sg13g2_nand3_1 _0904_ (.B(net184),
    .C(_0150_),
    .A(net248),
    .Y(_0164_));
 sg13g2_nand3_1 _0905_ (.B(\bav1.state_q[0] ),
    .C(_0149_),
    .A(net248),
    .Y(_0165_));
 sg13g2_nand2_1 _0906_ (.Y(_0002_),
    .A(_0164_),
    .B(_0165_));
 sg13g2_o21ai_1 _0907_ (.B1(net249),
    .Y(_0166_),
    .A1(_0154_),
    .A2(_0155_));
 sg13g2_nand2b_1 _0908_ (.Y(_0167_),
    .B(net167),
    .A_N(_0166_));
 sg13g2_a21oi_1 _0909_ (.A1(\bav0.state_q[2] ),
    .A2(_0155_),
    .Y(_0168_),
    .B1(\bav0._02_ ));
 sg13g2_o21ai_1 _0910_ (.B1(_0167_),
    .Y(_0009_),
    .A1(net236),
    .A2(_0168_));
 sg13g2_o21ai_1 _0911_ (.B1(net251),
    .Y(_0169_),
    .A1(_0148_),
    .A2(_0149_));
 sg13g2_a21oi_1 _0912_ (.A1(net184),
    .A2(_0148_),
    .Y(_0170_),
    .B1(\bav1._02_ ));
 sg13g2_a21oi_1 _0913_ (.A1(net252),
    .A2(_0170_),
    .Y(_0003_),
    .B1(net231));
 sg13g2_and2_1 _0914_ (.A(\io_sd._053_[0] ),
    .B(net243),
    .X(\rca.generate_adder_modules[0].fa.b ));
 sg13g2_and2_1 _0915_ (.A(\io_sd._053_[1] ),
    .B(net242),
    .X(\rca.generate_adder_modules[1].fa.b ));
 sg13g2_and2_1 _0916_ (.A(\io_sd._053_[2] ),
    .B(net242),
    .X(\rca.generate_adder_modules[2].fa.b ));
 sg13g2_and2_1 _0917_ (.A(\io_sd._053_[3] ),
    .B(net242),
    .X(\rca.generate_adder_modules[3].fa.b ));
 sg13g2_and2_1 _0918_ (.A(\io_sd._053_[4] ),
    .B(net244),
    .X(\rca.generate_adder_modules[4].fa.b ));
 sg13g2_and2_1 _0919_ (.A(\io_sd._053_[5] ),
    .B(net244),
    .X(\rca.generate_adder_modules[5].fa.b ));
 sg13g2_and2_1 _0920_ (.A(\io_sd._053_[6] ),
    .B(net244),
    .X(\rca.generate_adder_modules[6].fa.b ));
 sg13g2_and2_1 _0921_ (.A(\io_sd._053_[7] ),
    .B(net244),
    .X(\rca.generate_adder_modules[7].fa.b ));
 sg13g2_and2_1 _0922_ (.A(\io_sd._053_[8] ),
    .B(net240),
    .X(\rca.generate_adder_modules[8].fa.b ));
 sg13g2_and2_1 _0923_ (.A(\io_sd._053_[9] ),
    .B(net241),
    .X(\rca.generate_adder_modules[9].fa.b ));
 sg13g2_and2_2 _0924_ (.A(\io_sd._053_[10] ),
    .B(net240),
    .X(\rca.generate_adder_modules[10].fa.b ));
 sg13g2_and2_2 _0925_ (.A(\io_sd._053_[11] ),
    .B(net240),
    .X(\rca.generate_adder_modules[11].fa.b ));
 sg13g2_and2_1 _0926_ (.A(\io_sd._053_[12] ),
    .B(net240),
    .X(\rca.generate_adder_modules[12].fa.b ));
 sg13g2_and2_1 _0927_ (.A(\io_sd._053_[13] ),
    .B(net241),
    .X(\rca.generate_adder_modules[13].fa.b ));
 sg13g2_and2_2 _0928_ (.A(\io_sd._053_[14] ),
    .B(net241),
    .X(\rca.generate_adder_modules[14].fa.b ));
 sg13g2_and2_2 _0929_ (.A(\io_sd._053_[15] ),
    .B(net239),
    .X(\rca.generate_adder_modules[15].fa.b ));
 sg13g2_and2_1 _0930_ (.A(\io_sd._053_[16] ),
    .B(net239),
    .X(\rca.generate_adder_modules[16].fa.b ));
 sg13g2_and2_1 _0931_ (.A(\io_sd._053_[17] ),
    .B(net238),
    .X(\rca.generate_adder_modules[17].fa.b ));
 sg13g2_and2_2 _0932_ (.A(\io_sd._053_[18] ),
    .B(net238),
    .X(\rca.generate_adder_modules[18].fa.b ));
 sg13g2_and2_2 _0933_ (.A(\io_sd._053_[19] ),
    .B(net238),
    .X(\rca.generate_adder_modules[19].fa.b ));
 sg13g2_and2_2 _0934_ (.A(\io_sd._053_[20] ),
    .B(net238),
    .X(\rca.generate_adder_modules[20].fa.b ));
 sg13g2_and2_1 _0935_ (.A(\io_sd._053_[21] ),
    .B(net245),
    .X(\rca.generate_adder_modules[21].fa.b ));
 sg13g2_and2_2 _0936_ (.A(\io_sd._053_[22] ),
    .B(net239),
    .X(\rca.generate_adder_modules[22].fa.b ));
 sg13g2_and2_1 _0937_ (.A(\io_sd._053_[23] ),
    .B(net239),
    .X(\rca.generate_adder_modules[23].fa.b ));
 sg13g2_and2_1 _0938_ (.A(\io_sd._052_[0] ),
    .B(net243),
    .X(\rca.generate_adder_modules[0].fa.a ));
 sg13g2_and2_1 _0939_ (.A(\io_sd._052_[1] ),
    .B(net243),
    .X(\rca.generate_adder_modules[1].fa.a ));
 sg13g2_and2_1 _0940_ (.A(\io_sd._052_[2] ),
    .B(net242),
    .X(\rca.generate_adder_modules[2].fa.a ));
 sg13g2_and2_1 _0941_ (.A(\io_sd._052_[3] ),
    .B(net242),
    .X(\rca.generate_adder_modules[3].fa.a ));
 sg13g2_and2_2 _0942_ (.A(\io_sd._052_[4] ),
    .B(net242),
    .X(\rca.generate_adder_modules[4].fa.a ));
 sg13g2_and2_2 _0943_ (.A(\io_sd._052_[5] ),
    .B(net244),
    .X(\rca.generate_adder_modules[5].fa.a ));
 sg13g2_and2_2 _0944_ (.A(\io_sd._052_[6] ),
    .B(net244),
    .X(\rca.generate_adder_modules[6].fa.a ));
 sg13g2_and2_2 _0945_ (.A(\io_sd._052_[7] ),
    .B(net244),
    .X(\rca.generate_adder_modules[7].fa.a ));
 sg13g2_and2_2 _0946_ (.A(\io_sd._052_[8] ),
    .B(net242),
    .X(\rca.generate_adder_modules[8].fa.a ));
 sg13g2_and2_2 _0947_ (.A(\io_sd._052_[9] ),
    .B(net241),
    .X(\rca.generate_adder_modules[9].fa.a ));
 sg13g2_and2_2 _0948_ (.A(\io_sd._052_[10] ),
    .B(net240),
    .X(\rca.generate_adder_modules[10].fa.a ));
 sg13g2_and2_2 _0949_ (.A(\io_sd._052_[11] ),
    .B(net240),
    .X(\rca.generate_adder_modules[11].fa.a ));
 sg13g2_and2_2 _0950_ (.A(\io_sd._052_[12] ),
    .B(net240),
    .X(\rca.generate_adder_modules[12].fa.a ));
 sg13g2_and2_2 _0951_ (.A(\io_sd._052_[13] ),
    .B(net240),
    .X(\rca.generate_adder_modules[13].fa.a ));
 sg13g2_and2_2 _0952_ (.A(\io_sd._052_[14] ),
    .B(net241),
    .X(\rca.generate_adder_modules[14].fa.a ));
 sg13g2_and2_2 _0953_ (.A(\io_sd._052_[15] ),
    .B(net241),
    .X(\rca.generate_adder_modules[15].fa.a ));
 sg13g2_and2_2 _0954_ (.A(\io_sd._052_[16] ),
    .B(net241),
    .X(\rca.generate_adder_modules[16].fa.a ));
 sg13g2_and2_2 _0955_ (.A(\io_sd._052_[17] ),
    .B(net238),
    .X(\rca.generate_adder_modules[17].fa.a ));
 sg13g2_and2_2 _0956_ (.A(\io_sd._052_[18] ),
    .B(net238),
    .X(\rca.generate_adder_modules[18].fa.a ));
 sg13g2_and2_2 _0957_ (.A(\io_sd._052_[19] ),
    .B(net238),
    .X(\rca.generate_adder_modules[19].fa.a ));
 sg13g2_and2_2 _0958_ (.A(\io_sd._052_[20] ),
    .B(net238),
    .X(\rca.generate_adder_modules[20].fa.a ));
 sg13g2_and2_2 _0959_ (.A(\io_sd._052_[21] ),
    .B(net239),
    .X(\rca.generate_adder_modules[21].fa.a ));
 sg13g2_and2_2 _0960_ (.A(\io_sd._052_[22] ),
    .B(net239),
    .X(\rca.generate_adder_modules[22].fa.a ));
 sg13g2_and2_1 _0961_ (.A(\io_sd._052_[23] ),
    .B(net239),
    .X(\rca.generate_adder_modules[23].fa.a ));
 sg13g2_nand2_1 _0962_ (.Y(_0171_),
    .A(\io_sd.outputs[0] ),
    .B(net11));
 sg13g2_nand2b_1 _0963_ (.Y(_0172_),
    .B(net10),
    .A_N(\bav1._02_ ));
 sg13g2_o21ai_1 _0964_ (.B1(_0172_),
    .Y(_0173_),
    .A1(\bav0._02_ ),
    .A2(net10));
 sg13g2_o21ai_1 _0965_ (.B1(_0171_),
    .Y(uo_out[0]),
    .A1(net11),
    .A2(_0173_));
 sg13g2_nor2b_2 _0966_ (.A(net11),
    .B_N(net10),
    .Y(_0174_));
 sg13g2_a22oi_1 _0967_ (.Y(_0175_),
    .B1(_0174_),
    .B2(\ca._13_ ),
    .A2(net246),
    .A1(\io_sd.outputs[1] ));
 sg13g2_inv_1 _0968_ (.Y(uo_out[1]),
    .A(_0175_));
 sg13g2_a22oi_1 _0969_ (.Y(_0176_),
    .B1(_0174_),
    .B2(\bav1.x[0] ),
    .A2(net246),
    .A1(\io_sd.outputs[2] ));
 sg13g2_inv_1 _0970_ (.Y(uo_out[2]),
    .A(_0176_));
 sg13g2_a22oi_1 _0971_ (.Y(_0177_),
    .B1(_0174_),
    .B2(\bav1.x[1] ),
    .A2(net246),
    .A1(\io_sd.outputs[3] ));
 sg13g2_inv_1 _0972_ (.Y(uo_out[3]),
    .A(_0177_));
 sg13g2_a22oi_1 _0973_ (.Y(_0178_),
    .B1(\ca.coin_out[2] ),
    .B2(_0174_),
    .A2(net246),
    .A1(\io_sd.outputs[4] ));
 sg13g2_inv_1 _0974_ (.Y(uo_out[4]),
    .A(_0178_));
 sg13g2_a22oi_1 _0975_ (.Y(_0179_),
    .B1(\ca.coin_out[3] ),
    .B2(_0174_),
    .A2(net246),
    .A1(\io_sd.outputs[5] ));
 sg13g2_inv_1 _0976_ (.Y(uo_out[5]),
    .A(_0179_));
 sg13g2_a22oi_1 _0977_ (.Y(_0180_),
    .B1(\ca.coin_out[4] ),
    .B2(_0174_),
    .A2(net246),
    .A1(\io_sd.outputs[6] ));
 sg13g2_inv_1 _0978_ (.Y(uo_out[6]),
    .A(_0180_));
 sg13g2_a22oi_1 _0979_ (.Y(_0181_),
    .B1(\ca.coin_out[5] ),
    .B2(_0174_),
    .A2(net246),
    .A1(\io_sd.outputs[7] ));
 sg13g2_inv_1 _0980_ (.Y(uo_out[7]),
    .A(_0181_));
 sg13g2_nand2_1 _0981_ (.Y(_0182_),
    .A(\io_sd._053_[23] ),
    .B(\rca.generate_adder_modules[23].fa.a ));
 sg13g2_nand2_1 _0982_ (.Y(_0183_),
    .A(\io_sd._053_[21] ),
    .B(\rca.generate_adder_modules[21].fa.a ));
 sg13g2_nand2_1 _0983_ (.Y(_0184_),
    .A(\io_sd._053_[19] ),
    .B(\rca.generate_adder_modules[19].fa.a ));
 sg13g2_nand2_1 _0984_ (.Y(_0185_),
    .A(\io_sd._053_[17] ),
    .B(\rca.generate_adder_modules[17].fa.a ));
 sg13g2_nand2_1 _0985_ (.Y(_0186_),
    .A(\io_sd._053_[15] ),
    .B(\rca.generate_adder_modules[15].fa.a ));
 sg13g2_nand2_1 _0986_ (.Y(_0187_),
    .A(\io_sd._053_[13] ),
    .B(\rca.generate_adder_modules[13].fa.a ));
 sg13g2_nand2_1 _0987_ (.Y(_0188_),
    .A(\io_sd._053_[11] ),
    .B(\rca.generate_adder_modules[11].fa.a ));
 sg13g2_nand2_1 _0988_ (.Y(_0189_),
    .A(\io_sd._053_[9] ),
    .B(\rca.generate_adder_modules[9].fa.a ));
 sg13g2_nor2_1 _0989_ (.A(\rca.generate_adder_modules[9].fa.b ),
    .B(\rca.generate_adder_modules[9].fa.a ),
    .Y(_0190_));
 sg13g2_a21oi_1 _0990_ (.A1(\io_sd._053_[9] ),
    .A2(\rca.generate_adder_modules[9].fa.a ),
    .Y(_0191_),
    .B1(_0190_));
 sg13g2_nand2_1 _0991_ (.Y(_0192_),
    .A(\io_sd._053_[7] ),
    .B(\rca.generate_adder_modules[7].fa.a ));
 sg13g2_nand2_1 _0992_ (.Y(_0193_),
    .A(\io_sd._053_[5] ),
    .B(\rca.generate_adder_modules[5].fa.a ));
 sg13g2_nand2_1 _0993_ (.Y(_0194_),
    .A(\io_sd._053_[3] ),
    .B(\rca.generate_adder_modules[3].fa.a ));
 sg13g2_nand3_1 _0994_ (.B(\io_sd._052_[1] ),
    .C(net243),
    .A(\io_sd._053_[1] ),
    .Y(_0195_));
 sg13g2_nand3_1 _0995_ (.B(\io_sd._052_[0] ),
    .C(net243),
    .A(\io_sd._053_[0] ),
    .Y(_0196_));
 sg13g2_inv_1 _0996_ (.Y(_0197_),
    .A(_0196_));
 sg13g2_o21ai_1 _0997_ (.B1(net243),
    .Y(_0198_),
    .A1(\io_sd._053_[1] ),
    .A2(\io_sd._052_[1] ));
 sg13g2_a21oi_1 _0998_ (.A1(\io_sd._053_[1] ),
    .A2(\rca.generate_adder_modules[1].fa.a ),
    .Y(_0199_),
    .B1(_0198_));
 sg13g2_o21ai_1 _0999_ (.B1(_0195_),
    .Y(_0200_),
    .A1(_0196_),
    .A2(_0198_));
 sg13g2_o21ai_1 _1000_ (.B1(net242),
    .Y(_0201_),
    .A1(\io_sd._053_[2] ),
    .A2(\io_sd._052_[2] ));
 sg13g2_a21oi_1 _1001_ (.A1(\io_sd._053_[2] ),
    .A2(\rca.generate_adder_modules[2].fa.a ),
    .Y(_0202_),
    .B1(_0201_));
 sg13g2_a22oi_1 _1002_ (.Y(_0203_),
    .B1(_0200_),
    .B2(_0202_),
    .A2(\rca.generate_adder_modules[2].fa.a ),
    .A1(\io_sd._053_[2] ));
 sg13g2_nor2_1 _1003_ (.A(\rca.generate_adder_modules[3].fa.b ),
    .B(\rca.generate_adder_modules[3].fa.a ),
    .Y(_0204_));
 sg13g2_a21oi_1 _1004_ (.A1(\io_sd._053_[3] ),
    .A2(\rca.generate_adder_modules[3].fa.a ),
    .Y(_0205_),
    .B1(_0204_));
 sg13g2_o21ai_1 _1005_ (.B1(_0194_),
    .Y(_0206_),
    .A1(_0203_),
    .A2(_0204_));
 sg13g2_nor2_1 _1006_ (.A(\rca.generate_adder_modules[4].fa.b ),
    .B(\rca.generate_adder_modules[4].fa.a ),
    .Y(_0207_));
 sg13g2_a21oi_1 _1007_ (.A1(\io_sd._053_[4] ),
    .A2(\rca.generate_adder_modules[4].fa.a ),
    .Y(_0208_),
    .B1(_0207_));
 sg13g2_a22oi_1 _1008_ (.Y(_0209_),
    .B1(_0206_),
    .B2(_0208_),
    .A2(\rca.generate_adder_modules[4].fa.a ),
    .A1(\io_sd._053_[4] ));
 sg13g2_nor2_1 _1009_ (.A(\rca.generate_adder_modules[5].fa.b ),
    .B(\rca.generate_adder_modules[5].fa.a ),
    .Y(_0210_));
 sg13g2_a21oi_1 _1010_ (.A1(\io_sd._053_[5] ),
    .A2(\rca.generate_adder_modules[5].fa.a ),
    .Y(_0211_),
    .B1(_0210_));
 sg13g2_o21ai_1 _1011_ (.B1(_0193_),
    .Y(_0212_),
    .A1(_0209_),
    .A2(_0210_));
 sg13g2_nor2_1 _1012_ (.A(\rca.generate_adder_modules[6].fa.b ),
    .B(\rca.generate_adder_modules[6].fa.a ),
    .Y(_0213_));
 sg13g2_a21oi_1 _1013_ (.A1(\io_sd._053_[6] ),
    .A2(\rca.generate_adder_modules[6].fa.a ),
    .Y(_0214_),
    .B1(_0213_));
 sg13g2_a22oi_1 _1014_ (.Y(_0215_),
    .B1(_0212_),
    .B2(_0214_),
    .A2(\rca.generate_adder_modules[6].fa.a ),
    .A1(\io_sd._053_[6] ));
 sg13g2_nor2_1 _1015_ (.A(\rca.generate_adder_modules[7].fa.b ),
    .B(\rca.generate_adder_modules[7].fa.a ),
    .Y(_0216_));
 sg13g2_a21oi_1 _1016_ (.A1(\io_sd._053_[7] ),
    .A2(\rca.generate_adder_modules[7].fa.a ),
    .Y(_0217_),
    .B1(_0216_));
 sg13g2_o21ai_1 _1017_ (.B1(_0192_),
    .Y(_0218_),
    .A1(_0215_),
    .A2(_0216_));
 sg13g2_nor2_1 _1018_ (.A(\rca.generate_adder_modules[8].fa.b ),
    .B(\rca.generate_adder_modules[8].fa.a ),
    .Y(_0219_));
 sg13g2_a21oi_1 _1019_ (.A1(\io_sd._053_[8] ),
    .A2(\rca.generate_adder_modules[8].fa.a ),
    .Y(_0220_),
    .B1(_0219_));
 sg13g2_a22oi_1 _1020_ (.Y(_0221_),
    .B1(_0218_),
    .B2(_0220_),
    .A2(\rca.generate_adder_modules[8].fa.a ),
    .A1(\io_sd._053_[8] ));
 sg13g2_o21ai_1 _1021_ (.B1(_0189_),
    .Y(_0222_),
    .A1(_0190_),
    .A2(_0221_));
 sg13g2_nor2_1 _1022_ (.A(\rca.generate_adder_modules[10].fa.b ),
    .B(\rca.generate_adder_modules[10].fa.a ),
    .Y(_0223_));
 sg13g2_a21oi_1 _1023_ (.A1(\io_sd._053_[10] ),
    .A2(\rca.generate_adder_modules[10].fa.a ),
    .Y(_0224_),
    .B1(_0223_));
 sg13g2_a22oi_1 _1024_ (.Y(_0225_),
    .B1(_0222_),
    .B2(_0224_),
    .A2(\rca.generate_adder_modules[10].fa.a ),
    .A1(\io_sd._053_[10] ));
 sg13g2_nor2_1 _1025_ (.A(\rca.generate_adder_modules[11].fa.b ),
    .B(\rca.generate_adder_modules[11].fa.a ),
    .Y(_0226_));
 sg13g2_a21oi_1 _1026_ (.A1(\io_sd._053_[11] ),
    .A2(\rca.generate_adder_modules[11].fa.a ),
    .Y(_0227_),
    .B1(_0226_));
 sg13g2_o21ai_1 _1027_ (.B1(_0188_),
    .Y(_0228_),
    .A1(_0225_),
    .A2(_0226_));
 sg13g2_nor2_1 _1028_ (.A(\rca.generate_adder_modules[12].fa.b ),
    .B(\rca.generate_adder_modules[12].fa.a ),
    .Y(_0229_));
 sg13g2_a21oi_1 _1029_ (.A1(\io_sd._053_[12] ),
    .A2(\rca.generate_adder_modules[12].fa.a ),
    .Y(_0230_),
    .B1(_0229_));
 sg13g2_a22oi_1 _1030_ (.Y(_0231_),
    .B1(_0228_),
    .B2(_0230_),
    .A2(\rca.generate_adder_modules[12].fa.a ),
    .A1(\io_sd._053_[12] ));
 sg13g2_nor2_1 _1031_ (.A(\rca.generate_adder_modules[13].fa.b ),
    .B(\rca.generate_adder_modules[13].fa.a ),
    .Y(_0232_));
 sg13g2_a21oi_1 _1032_ (.A1(\io_sd._053_[13] ),
    .A2(\rca.generate_adder_modules[13].fa.a ),
    .Y(_0233_),
    .B1(_0232_));
 sg13g2_o21ai_1 _1033_ (.B1(_0187_),
    .Y(_0234_),
    .A1(_0231_),
    .A2(_0232_));
 sg13g2_nor2_1 _1034_ (.A(\rca.generate_adder_modules[14].fa.b ),
    .B(\rca.generate_adder_modules[14].fa.a ),
    .Y(_0235_));
 sg13g2_a21oi_1 _1035_ (.A1(\io_sd._053_[14] ),
    .A2(\rca.generate_adder_modules[14].fa.a ),
    .Y(_0236_),
    .B1(_0235_));
 sg13g2_a22oi_1 _1036_ (.Y(_0237_),
    .B1(_0234_),
    .B2(_0236_),
    .A2(\rca.generate_adder_modules[14].fa.a ),
    .A1(\io_sd._053_[14] ));
 sg13g2_nor2_1 _1037_ (.A(\rca.generate_adder_modules[15].fa.b ),
    .B(\rca.generate_adder_modules[15].fa.a ),
    .Y(_0238_));
 sg13g2_a21oi_1 _1038_ (.A1(\io_sd._053_[15] ),
    .A2(\rca.generate_adder_modules[15].fa.a ),
    .Y(_0239_),
    .B1(_0238_));
 sg13g2_o21ai_1 _1039_ (.B1(_0186_),
    .Y(_0240_),
    .A1(_0237_),
    .A2(_0238_));
 sg13g2_nor2_1 _1040_ (.A(\rca.generate_adder_modules[16].fa.b ),
    .B(\rca.generate_adder_modules[16].fa.a ),
    .Y(_0241_));
 sg13g2_a21oi_1 _1041_ (.A1(\io_sd._053_[16] ),
    .A2(\rca.generate_adder_modules[16].fa.a ),
    .Y(_0242_),
    .B1(_0241_));
 sg13g2_a22oi_1 _1042_ (.Y(_0243_),
    .B1(_0240_),
    .B2(_0242_),
    .A2(\rca.generate_adder_modules[16].fa.a ),
    .A1(\io_sd._053_[16] ));
 sg13g2_nor2_1 _1043_ (.A(\rca.generate_adder_modules[17].fa.b ),
    .B(\rca.generate_adder_modules[17].fa.a ),
    .Y(_0244_));
 sg13g2_a21oi_1 _1044_ (.A1(\io_sd._053_[17] ),
    .A2(\rca.generate_adder_modules[17].fa.a ),
    .Y(_0245_),
    .B1(_0244_));
 sg13g2_o21ai_1 _1045_ (.B1(_0185_),
    .Y(_0246_),
    .A1(_0243_),
    .A2(_0244_));
 sg13g2_nor2_1 _1046_ (.A(\rca.generate_adder_modules[18].fa.b ),
    .B(\rca.generate_adder_modules[18].fa.a ),
    .Y(_0247_));
 sg13g2_a21oi_1 _1047_ (.A1(\io_sd._053_[18] ),
    .A2(\rca.generate_adder_modules[18].fa.a ),
    .Y(_0248_),
    .B1(_0247_));
 sg13g2_a22oi_1 _1048_ (.Y(_0249_),
    .B1(_0246_),
    .B2(_0248_),
    .A2(\rca.generate_adder_modules[18].fa.a ),
    .A1(\io_sd._053_[18] ));
 sg13g2_nor2_1 _1049_ (.A(\rca.generate_adder_modules[19].fa.b ),
    .B(\rca.generate_adder_modules[19].fa.a ),
    .Y(_0250_));
 sg13g2_a21oi_1 _1050_ (.A1(\io_sd._053_[19] ),
    .A2(\rca.generate_adder_modules[19].fa.a ),
    .Y(_0251_),
    .B1(_0250_));
 sg13g2_o21ai_1 _1051_ (.B1(_0184_),
    .Y(_0252_),
    .A1(_0249_),
    .A2(_0250_));
 sg13g2_nor2_1 _1052_ (.A(\rca.generate_adder_modules[20].fa.b ),
    .B(\rca.generate_adder_modules[20].fa.a ),
    .Y(_0253_));
 sg13g2_a21oi_1 _1053_ (.A1(\io_sd._053_[20] ),
    .A2(\rca.generate_adder_modules[20].fa.a ),
    .Y(_0254_),
    .B1(_0253_));
 sg13g2_a22oi_1 _1054_ (.Y(_0255_),
    .B1(_0252_),
    .B2(_0254_),
    .A2(\rca.generate_adder_modules[20].fa.a ),
    .A1(\io_sd._053_[20] ));
 sg13g2_nor2_1 _1055_ (.A(\rca.generate_adder_modules[21].fa.b ),
    .B(\rca.generate_adder_modules[21].fa.a ),
    .Y(_0256_));
 sg13g2_a21oi_1 _1056_ (.A1(\io_sd._053_[21] ),
    .A2(\rca.generate_adder_modules[21].fa.a ),
    .Y(_0257_),
    .B1(_0256_));
 sg13g2_o21ai_1 _1057_ (.B1(_0183_),
    .Y(_0258_),
    .A1(_0255_),
    .A2(_0256_));
 sg13g2_nor2_1 _1058_ (.A(\rca.generate_adder_modules[22].fa.b ),
    .B(\rca.generate_adder_modules[22].fa.a ),
    .Y(_0259_));
 sg13g2_a21oi_1 _1059_ (.A1(\io_sd._053_[22] ),
    .A2(\rca.generate_adder_modules[22].fa.a ),
    .Y(_0260_),
    .B1(_0259_));
 sg13g2_a22oi_1 _1060_ (.Y(_0261_),
    .B1(_0258_),
    .B2(_0260_),
    .A2(\rca.generate_adder_modules[22].fa.a ),
    .A1(\io_sd._053_[22] ));
 sg13g2_o21ai_1 _1061_ (.B1(_0182_),
    .Y(_0262_),
    .A1(\rca.generate_adder_modules[23].fa.b ),
    .A2(\rca.generate_adder_modules[23].fa.a ));
 sg13g2_o21ai_1 _1062_ (.B1(_0182_),
    .Y(\rca.generate_adder_modules[23].fa._02_ ),
    .A1(_0261_),
    .A2(_0262_));
 sg13g2_mux2_1 _1063_ (.A0(_0142_),
    .A1(net211),
    .S(net220),
    .X(_0016_));
 sg13g2_nand2_1 _1064_ (.Y(_0263_),
    .A(net12),
    .B(_0139_));
 sg13g2_o21ai_1 _1065_ (.B1(net331),
    .Y(_0264_),
    .A1(_0131_),
    .A2(net220));
 sg13g2_nand3_1 _1066_ (.B(_0263_),
    .C(net332),
    .A(net247),
    .Y(_0017_));
 sg13g2_nor3_1 _1067_ (.A(_0010_),
    .B(_0138_),
    .C(_0139_),
    .Y(_0265_));
 sg13g2_a21o_1 _1068_ (.A2(net210),
    .A1(net292),
    .B1(_0265_),
    .X(_0018_));
 sg13g2_nor2b_1 _1069_ (.A(\ca.commit_count[16] ),
    .B_N(\ca.commit_count[17] ),
    .Y(_0266_));
 sg13g2_nand3b_1 _1070_ (.B(\ca.commit_count[11] ),
    .C(_0266_),
    .Y(_0267_),
    .A_N(\ca.commit_count[12] ));
 sg13g2_nand4_1 _1071_ (.B(\ca.commit_count[20] ),
    .C(_0132_),
    .A(\ca.commit_count[21] ),
    .Y(_0268_),
    .D(\ca.commit_count[18] ));
 sg13g2_nor4_1 _1072_ (.A(\ca.commit_count[6] ),
    .B(\ca.commit_count[5] ),
    .C(\ca.commit_count[4] ),
    .D(\ca.commit_count[3] ),
    .Y(_0269_));
 sg13g2_nor2b_1 _1073_ (.A(\ca.commit_count[8] ),
    .B_N(\ca.commit_count[7] ),
    .Y(_0270_));
 sg13g2_nand4_1 _1074_ (.B(\ca.commit_count[9] ),
    .C(_0269_),
    .A(\ca.commit_count[10] ),
    .Y(_0271_),
    .D(_0270_));
 sg13g2_nand3_1 _1075_ (.B(\ca.commit_count[14] ),
    .C(\ca.commit_count[13] ),
    .A(\ca.commit_count[15] ),
    .Y(_0272_));
 sg13g2_inv_1 _1076_ (.Y(_0273_),
    .A(_0272_));
 sg13g2_or4_1 _1077_ (.A(\ca.commit_count[2] ),
    .B(\ca.commit_count[1] ),
    .C(\ca.commit_count[0] ),
    .D(_0272_),
    .X(_0274_));
 sg13g2_nor4_2 _1078_ (.A(_0267_),
    .B(_0268_),
    .C(_0271_),
    .Y(_0275_),
    .D(_0274_));
 sg13g2_and2_2 _1079_ (.A(net247),
    .B(_0275_),
    .X(_0276_));
 sg13g2_and2_1 _1080_ (.A(net160),
    .B(_0276_),
    .X(_0019_));
 sg13g2_and2_1 _1081_ (.A(net152),
    .B(_0276_),
    .X(_0020_));
 sg13g2_and2_1 _1082_ (.A(net144),
    .B(_0276_),
    .X(_0021_));
 sg13g2_and2_1 _1083_ (.A(net143),
    .B(_0276_),
    .X(_0022_));
 sg13g2_and2_1 _1084_ (.A(net159),
    .B(_0276_),
    .X(_0023_));
 sg13g2_and2_1 _1085_ (.A(net161),
    .B(_0276_),
    .X(_0024_));
 sg13g2_nand3_1 _1086_ (.B(net344),
    .C(_0139_),
    .A(net12),
    .Y(_0277_));
 sg13g2_nand3_1 _1087_ (.B(net247),
    .C(_0277_),
    .A(net214),
    .Y(_0025_));
 sg13g2_nand2b_1 _1088_ (.Y(_0026_),
    .B(net247),
    .A_N(net163));
 sg13g2_and2_1 _1089_ (.A(\ca.commit_count[11] ),
    .B(\ca.commit_count[10] ),
    .X(_0278_));
 sg13g2_nand2b_2 _1090_ (.Y(_0279_),
    .B(net247),
    .A_N(_0275_));
 sg13g2_inv_1 _1091_ (.Y(_0280_),
    .A(_0279_));
 sg13g2_nor2b_1 _1092_ (.A(net162),
    .B_N(net169),
    .Y(_0281_));
 sg13g2_or2_1 _1093_ (.X(_0282_),
    .B(_0281_),
    .A(_0279_));
 sg13g2_inv_1 _1094_ (.Y(_0283_),
    .A(net194));
 sg13g2_nor2b_1 _1095_ (.A(\ca._15_ ),
    .B_N(\ca.commit_count[0] ),
    .Y(_0284_));
 sg13g2_a21oi_1 _1096_ (.A1(\ca._15_ ),
    .A2(net141),
    .Y(_0285_),
    .B1(_0284_));
 sg13g2_nor2_1 _1097_ (.A(net195),
    .B(net142),
    .Y(_0027_));
 sg13g2_and3_1 _1098_ (.X(_0286_),
    .A(\ca._15_ ),
    .B(net164),
    .C(\ca.commit_count[0] ));
 sg13g2_a21oi_1 _1099_ (.A1(\ca._15_ ),
    .A2(\ca.commit_count[0] ),
    .Y(_0287_),
    .B1(net164));
 sg13g2_nor3_1 _1100_ (.A(net195),
    .B(_0286_),
    .C(net165),
    .Y(_0028_));
 sg13g2_and2_1 _1101_ (.A(net260),
    .B(_0286_),
    .X(_0288_));
 sg13g2_nor2_1 _1102_ (.A(net260),
    .B(_0286_),
    .Y(_0289_));
 sg13g2_nor3_1 _1103_ (.A(net193),
    .B(_0288_),
    .C(net261),
    .Y(_0029_));
 sg13g2_and2_1 _1104_ (.A(net277),
    .B(_0288_),
    .X(_0290_));
 sg13g2_nor2_1 _1105_ (.A(net277),
    .B(_0288_),
    .Y(_0291_));
 sg13g2_nor3_1 _1106_ (.A(net195),
    .B(_0290_),
    .C(_0291_),
    .Y(_0030_));
 sg13g2_and2_1 _1107_ (.A(net269),
    .B(_0290_),
    .X(_0292_));
 sg13g2_nor2_1 _1108_ (.A(net269),
    .B(_0290_),
    .Y(_0293_));
 sg13g2_nor3_1 _1109_ (.A(net193),
    .B(_0292_),
    .C(net270),
    .Y(_0031_));
 sg13g2_and2_1 _1110_ (.A(net271),
    .B(_0292_),
    .X(_0294_));
 sg13g2_nor2_1 _1111_ (.A(net271),
    .B(_0292_),
    .Y(_0295_));
 sg13g2_nor3_1 _1112_ (.A(net193),
    .B(_0294_),
    .C(_0295_),
    .Y(_0032_));
 sg13g2_nor2_1 _1113_ (.A(net303),
    .B(_0294_),
    .Y(_0296_));
 sg13g2_and2_1 _1114_ (.A(net303),
    .B(_0294_),
    .X(_0297_));
 sg13g2_nor3_1 _1115_ (.A(net193),
    .B(_0296_),
    .C(_0297_),
    .Y(_0033_));
 sg13g2_nor2_1 _1116_ (.A(net280),
    .B(_0297_),
    .Y(_0298_));
 sg13g2_and2_1 _1117_ (.A(net280),
    .B(_0297_),
    .X(_0299_));
 sg13g2_nor3_1 _1118_ (.A(net193),
    .B(net281),
    .C(_0299_),
    .Y(_0034_));
 sg13g2_xnor2_1 _1119_ (.Y(_0300_),
    .A(net318),
    .B(_0299_));
 sg13g2_nor2_1 _1120_ (.A(net193),
    .B(_0300_),
    .Y(_0035_));
 sg13g2_a21oi_1 _1121_ (.A1(\ca.commit_count[8] ),
    .A2(_0299_),
    .Y(_0301_),
    .B1(net172));
 sg13g2_and3_1 _1122_ (.X(_0302_),
    .A(net172),
    .B(net318),
    .C(_0299_));
 sg13g2_nor3_1 _1123_ (.A(net193),
    .B(net173),
    .C(_0302_),
    .Y(_0036_));
 sg13g2_and2_1 _1124_ (.A(net337),
    .B(_0302_),
    .X(_0303_));
 sg13g2_o21ai_1 _1125_ (.B1(_0283_),
    .Y(_0304_),
    .A1(net337),
    .A2(_0302_));
 sg13g2_nor2_1 _1126_ (.A(_0303_),
    .B(_0304_),
    .Y(_0037_));
 sg13g2_and2_1 _1127_ (.A(net335),
    .B(_0303_),
    .X(_0305_));
 sg13g2_o21ai_1 _1128_ (.B1(_0283_),
    .Y(_0306_),
    .A1(net335),
    .A2(_0303_));
 sg13g2_nor2_1 _1129_ (.A(_0305_),
    .B(net336),
    .Y(_0038_));
 sg13g2_nor2_1 _1130_ (.A(net316),
    .B(_0305_),
    .Y(_0307_));
 sg13g2_and2_1 _1131_ (.A(net316),
    .B(_0305_),
    .X(_0308_));
 sg13g2_nor3_1 _1132_ (.A(net193),
    .B(net317),
    .C(_0308_),
    .Y(_0039_));
 sg13g2_nor2_1 _1133_ (.A(net312),
    .B(_0308_),
    .Y(_0309_));
 sg13g2_and2_1 _1134_ (.A(net312),
    .B(_0308_),
    .X(_0310_));
 sg13g2_and4_1 _1135_ (.A(net312),
    .B(net316),
    .C(_0278_),
    .D(_0302_),
    .X(_0311_));
 sg13g2_nor3_1 _1136_ (.A(net194),
    .B(net313),
    .C(_0310_),
    .Y(_0040_));
 sg13g2_and2_1 _1137_ (.A(net330),
    .B(_0310_),
    .X(_0312_));
 sg13g2_o21ai_1 _1138_ (.B1(_0283_),
    .Y(_0313_),
    .A1(net330),
    .A2(_0311_));
 sg13g2_nor2_1 _1139_ (.A(_0312_),
    .B(_0313_),
    .Y(_0041_));
 sg13g2_nor2_1 _1140_ (.A(net306),
    .B(_0312_),
    .Y(_0314_));
 sg13g2_and2_1 _1141_ (.A(net306),
    .B(_0312_),
    .X(_0315_));
 sg13g2_nor3_1 _1142_ (.A(net194),
    .B(net307),
    .C(_0315_),
    .Y(_0042_));
 sg13g2_a21oi_1 _1143_ (.A1(net338),
    .A2(_0315_),
    .Y(_0316_),
    .B1(net194));
 sg13g2_and4_1 _1144_ (.A(\ca.commit_count[16] ),
    .B(net306),
    .C(\ca.commit_count[14] ),
    .D(_0311_),
    .X(_0317_));
 sg13g2_o21ai_1 _1145_ (.B1(_0316_),
    .Y(_0318_),
    .A1(net338),
    .A2(_0315_));
 sg13g2_inv_1 _1146_ (.Y(_0043_),
    .A(_0318_));
 sg13g2_nor2_1 _1147_ (.A(net309),
    .B(_0317_),
    .Y(_0319_));
 sg13g2_and4_2 _1148_ (.A(net309),
    .B(\ca.commit_count[16] ),
    .C(_0273_),
    .D(_0308_),
    .X(_0320_));
 sg13g2_nor3_1 _1149_ (.A(net194),
    .B(net310),
    .C(_0320_),
    .Y(_0044_));
 sg13g2_o21ai_1 _1150_ (.B1(_0283_),
    .Y(_0321_),
    .A1(net297),
    .A2(_0320_));
 sg13g2_a21oi_1 _1151_ (.A1(net297),
    .A2(_0320_),
    .Y(_0045_),
    .B1(_0321_));
 sg13g2_a21oi_1 _1152_ (.A1(\ca.commit_count[18] ),
    .A2(_0320_),
    .Y(_0322_),
    .B1(net257));
 sg13g2_and4_1 _1153_ (.A(net257),
    .B(\ca.commit_count[18] ),
    .C(\ca.commit_count[17] ),
    .D(_0317_),
    .X(_0323_));
 sg13g2_nor3_1 _1154_ (.A(net194),
    .B(net258),
    .C(_0323_),
    .Y(_0046_));
 sg13g2_nor2_1 _1155_ (.A(net295),
    .B(_0323_),
    .Y(_0324_));
 sg13g2_and4_1 _1156_ (.A(net295),
    .B(net257),
    .C(net297),
    .D(_0320_),
    .X(_0325_));
 sg13g2_nor3_1 _1157_ (.A(net194),
    .B(net296),
    .C(_0325_),
    .Y(_0047_));
 sg13g2_a21oi_1 _1158_ (.A1(net327),
    .A2(_0325_),
    .Y(_0326_),
    .B1(net194));
 sg13g2_o21ai_1 _1159_ (.B1(_0326_),
    .Y(_0327_),
    .A1(net327),
    .A2(_0325_));
 sg13g2_inv_1 _1160_ (.Y(_0048_),
    .A(_0327_));
 sg13g2_a22oi_1 _1161_ (.Y(_0328_),
    .B1(_0281_),
    .B2(net247),
    .A2(_0280_),
    .A1(net323));
 sg13g2_inv_1 _1162_ (.Y(_0049_),
    .A(_0328_));
 sg13g2_nor2b_2 _1163_ (.A(net169),
    .B_N(net162),
    .Y(_0329_));
 sg13g2_nor2b_1 _1164_ (.A(_0329_),
    .B_N(\ca.pulse_count[0] ),
    .Y(_0330_));
 sg13g2_a21oi_1 _1165_ (.A1(net139),
    .A2(_0329_),
    .Y(_0331_),
    .B1(_0330_));
 sg13g2_nor2_1 _1166_ (.A(_0279_),
    .B(net140),
    .Y(_0050_));
 sg13g2_and3_1 _1167_ (.X(_0332_),
    .A(net152),
    .B(net160),
    .C(_0329_));
 sg13g2_a21oi_1 _1168_ (.A1(net160),
    .A2(_0329_),
    .Y(_0333_),
    .B1(net152));
 sg13g2_nor3_1 _1169_ (.A(_0279_),
    .B(_0332_),
    .C(_0333_),
    .Y(_0051_));
 sg13g2_and2_1 _1170_ (.A(net144),
    .B(_0332_),
    .X(_0334_));
 sg13g2_nor2_1 _1171_ (.A(net144),
    .B(_0332_),
    .Y(_0335_));
 sg13g2_nor3_1 _1172_ (.A(_0279_),
    .B(_0334_),
    .C(_0335_),
    .Y(_0052_));
 sg13g2_and2_1 _1173_ (.A(net143),
    .B(_0334_),
    .X(_0336_));
 sg13g2_nor2_1 _1174_ (.A(net143),
    .B(_0334_),
    .Y(_0337_));
 sg13g2_nor3_1 _1175_ (.A(_0279_),
    .B(_0336_),
    .C(_0337_),
    .Y(_0053_));
 sg13g2_nor2_1 _1176_ (.A(net159),
    .B(_0336_),
    .Y(_0338_));
 sg13g2_and2_1 _1177_ (.A(net159),
    .B(_0336_),
    .X(_0339_));
 sg13g2_nor3_1 _1178_ (.A(_0279_),
    .B(_0338_),
    .C(_0339_),
    .Y(_0054_));
 sg13g2_a21oi_1 _1179_ (.A1(net161),
    .A2(_0339_),
    .Y(_0340_),
    .B1(_0279_));
 sg13g2_o21ai_1 _1180_ (.B1(_0340_),
    .Y(_0341_),
    .A1(net161),
    .A2(_0339_));
 sg13g2_inv_1 _1181_ (.Y(_0055_),
    .A(_0341_));
 sg13g2_nand2b_1 _1182_ (.Y(_0057_),
    .B(net247),
    .A_N(net162));
 sg13g2_nor2_2 _1183_ (.A(net12),
    .B(_0136_),
    .Y(_0342_));
 sg13g2_nand2_1 _1184_ (.Y(_0343_),
    .A(_0131_),
    .B(\io_sd._083_ ));
 sg13g2_nor2b_2 _1185_ (.A(net12),
    .B_N(\io_sd._080_ ),
    .Y(_0344_));
 sg13g2_nand2_1 _1186_ (.Y(_0345_),
    .A(_0131_),
    .B(net262));
 sg13g2_nor2_2 _1187_ (.A(net202),
    .B(net206),
    .Y(_0346_));
 sg13g2_xnor2_1 _1188_ (.Y(_0347_),
    .A(net343),
    .B(_0346_));
 sg13g2_and3_1 _1189_ (.X(_0058_),
    .A(net249),
    .B(_0146_),
    .C(_0347_));
 sg13g2_o21ai_1 _1190_ (.B1(net328),
    .Y(_0348_),
    .A1(\io_sd.input_index[3] ),
    .A2(_0346_));
 sg13g2_o21ai_1 _1191_ (.B1(_0145_),
    .Y(_0349_),
    .A1(net202),
    .A2(net206));
 sg13g2_nand3_1 _1192_ (.B(net329),
    .C(_0349_),
    .A(net249),
    .Y(_0059_));
 sg13g2_nor2_1 _1193_ (.A(_0011_),
    .B(_0145_),
    .Y(_0350_));
 sg13g2_nor2_1 _1194_ (.A(_0346_),
    .B(_0350_),
    .Y(_0351_));
 sg13g2_nor3_1 _1195_ (.A(net339),
    .B(net202),
    .C(net206),
    .Y(_0352_));
 sg13g2_nor3_1 _1196_ (.A(net236),
    .B(_0351_),
    .C(_0352_),
    .Y(_0060_));
 sg13g2_nand2_1 _1197_ (.Y(_0353_),
    .A(net153),
    .B(net211));
 sg13g2_nor2_2 _1198_ (.A(net218),
    .B(net219),
    .Y(_0354_));
 sg13g2_nand2_2 _1199_ (.Y(_0355_),
    .A(net212),
    .B(_0134_));
 sg13g2_nand2_1 _1200_ (.Y(_0356_),
    .A(_0013_),
    .B(_0354_));
 sg13g2_nand2_1 _1201_ (.Y(_0357_),
    .A(_0010_),
    .B(_0356_));
 sg13g2_or2_1 _1202_ (.X(_0358_),
    .B(_0356_),
    .A(_0010_));
 sg13g2_nor2_2 _1203_ (.A(net212),
    .B(_0134_),
    .Y(_0359_));
 sg13g2_nand2_2 _1204_ (.Y(_0360_),
    .A(\io_sd._209_[0] ),
    .B(net219));
 sg13g2_nor2_1 _1205_ (.A(_0013_),
    .B(_0360_),
    .Y(_0361_));
 sg13g2_a21oi_1 _1206_ (.A1(_0013_),
    .A2(_0354_),
    .Y(_0362_),
    .B1(_0361_));
 sg13g2_o21ai_1 _1207_ (.B1(_0357_),
    .Y(_0363_),
    .A1(_0010_),
    .A2(_0361_));
 sg13g2_a21o_2 _1208_ (.A2(_0358_),
    .A1(_0357_),
    .B1(_0138_),
    .X(_0364_));
 sg13g2_nand2_2 _1209_ (.Y(_0365_),
    .A(_0355_),
    .B(_0360_));
 sg13g2_nor2_2 _1210_ (.A(_0013_),
    .B(_0365_),
    .Y(_0366_));
 sg13g2_or2_1 _1211_ (.X(_0367_),
    .B(_0365_),
    .A(_0013_));
 sg13g2_nand2_2 _1212_ (.Y(_0368_),
    .A(_0362_),
    .B(_0367_));
 sg13g2_nor2b_1 _1213_ (.A(net10),
    .B_N(net246),
    .Y(_0369_));
 sg13g2_xor2_1 _1214_ (.B(_0221_),
    .A(_0191_),
    .X(_0370_));
 sg13g2_nand3_1 _1215_ (.B(\io_sd.output_index[4] ),
    .C(_0359_),
    .A(\io_sd.output_index[5] ),
    .Y(_0371_));
 sg13g2_xor2_1 _1216_ (.B(_0371_),
    .A(_0363_),
    .X(_0372_));
 sg13g2_xnor2_1 _1217_ (.Y(_0373_),
    .A(_0363_),
    .B(_0371_));
 sg13g2_a21oi_1 _1218_ (.A1(net224),
    .A2(_0370_),
    .Y(_0374_),
    .B1(_0372_));
 sg13g2_o21ai_1 _1219_ (.B1(_0374_),
    .Y(_0375_),
    .A1(\cla_z[9] ),
    .A2(net224));
 sg13g2_nor2_1 _1220_ (.A(_0355_),
    .B(_0375_),
    .Y(_0376_));
 sg13g2_nor2_1 _1221_ (.A(\cla_z[1] ),
    .B(net228),
    .Y(_0377_));
 sg13g2_xnor2_1 _1222_ (.Y(_0378_),
    .A(_0197_),
    .B(_0199_));
 sg13g2_a21oi_1 _1223_ (.A1(net226),
    .A2(_0378_),
    .Y(_0379_),
    .B1(_0377_));
 sg13g2_nor2_1 _1224_ (.A(\rca.generate_adder_modules[0].fa.b ),
    .B(\rca.generate_adder_modules[0].fa.a ),
    .Y(_0380_));
 sg13g2_o21ai_1 _1225_ (.B1(net226),
    .Y(_0381_),
    .A1(_0197_),
    .A2(_0380_));
 sg13g2_o21ai_1 _1226_ (.B1(_0381_),
    .Y(_0382_),
    .A1(\cla_z[0] ),
    .A2(net226));
 sg13g2_a21oi_1 _1227_ (.A1(_0134_),
    .A2(_0382_),
    .Y(_0383_),
    .B1(_0365_));
 sg13g2_o21ai_1 _1228_ (.B1(_0383_),
    .Y(_0384_),
    .A1(net218),
    .A2(_0379_));
 sg13g2_xnor2_1 _1229_ (.Y(_0385_),
    .A(_0218_),
    .B(_0220_));
 sg13g2_o21ai_1 _1230_ (.B1(net191),
    .Y(_0386_),
    .A1(\cla_z[8] ),
    .A2(net225));
 sg13g2_a21oi_2 _1231_ (.B1(_0386_),
    .Y(_0387_),
    .A2(_0385_),
    .A1(net226));
 sg13g2_a21oi_1 _1232_ (.A1(_0359_),
    .A2(_0387_),
    .Y(_0388_),
    .B1(_0376_));
 sg13g2_a21oi_1 _1233_ (.A1(_0384_),
    .A2(_0388_),
    .Y(_0389_),
    .B1(_0368_));
 sg13g2_xor2_1 _1234_ (.B(_0245_),
    .A(_0243_),
    .X(_0390_));
 sg13g2_a21oi_1 _1235_ (.A1(net221),
    .A2(_0390_),
    .Y(_0391_),
    .B1(net192));
 sg13g2_o21ai_1 _1236_ (.B1(_0391_),
    .Y(_0392_),
    .A1(\cla_z[17] ),
    .A2(net221));
 sg13g2_nand2_1 _1237_ (.Y(_0393_),
    .A(net212),
    .B(_0392_));
 sg13g2_xnor2_1 _1238_ (.Y(_0394_),
    .A(_0240_),
    .B(_0242_));
 sg13g2_a21oi_1 _1239_ (.A1(net222),
    .A2(_0394_),
    .Y(_0395_),
    .B1(net192));
 sg13g2_o21ai_1 _1240_ (.B1(_0395_),
    .Y(_0396_),
    .A1(\cla_z[16] ),
    .A2(net222));
 sg13g2_a21oi_1 _1241_ (.A1(\io_sd._209_[0] ),
    .A2(_0396_),
    .Y(_0397_),
    .B1(_0367_));
 sg13g2_a21oi_1 _1242_ (.A1(_0393_),
    .A2(_0397_),
    .Y(_0398_),
    .B1(_0389_));
 sg13g2_o21ai_1 _1243_ (.B1(_0353_),
    .Y(_0061_),
    .A1(_0364_),
    .A2(_0398_));
 sg13g2_nand2_1 _1244_ (.Y(_0399_),
    .A(net150),
    .B(net210));
 sg13g2_xnor2_1 _1245_ (.Y(_0400_),
    .A(_0222_),
    .B(_0224_));
 sg13g2_o21ai_1 _1246_ (.B1(net191),
    .Y(_0401_),
    .A1(\cla_z[10] ),
    .A2(net224));
 sg13g2_a21oi_1 _1247_ (.A1(net224),
    .A2(_0400_),
    .Y(_0402_),
    .B1(_0401_));
 sg13g2_inv_1 _1248_ (.Y(_0403_),
    .A(_0402_));
 sg13g2_xnor2_1 _1249_ (.Y(_0404_),
    .A(_0200_),
    .B(_0202_));
 sg13g2_o21ai_1 _1250_ (.B1(net191),
    .Y(_0405_),
    .A1(\cla_z[2] ),
    .A2(net226));
 sg13g2_a21oi_1 _1251_ (.A1(net226),
    .A2(_0404_),
    .Y(_0406_),
    .B1(_0405_));
 sg13g2_nor2_1 _1252_ (.A(net213),
    .B(net192),
    .Y(_0407_));
 sg13g2_a221oi_1 _1253_ (.B2(_0379_),
    .C1(_0365_),
    .B1(_0407_),
    .A1(net212),
    .Y(_0408_),
    .A2(_0406_));
 sg13g2_nor2_1 _1254_ (.A(_0368_),
    .B(_0408_),
    .Y(_0409_));
 sg13g2_a22oi_1 _1255_ (.Y(_0410_),
    .B1(_0403_),
    .B2(_0354_),
    .A2(_0375_),
    .A1(_0359_));
 sg13g2_xnor2_1 _1256_ (.Y(_0411_),
    .A(_0246_),
    .B(_0248_));
 sg13g2_o21ai_1 _1257_ (.B1(net190),
    .Y(_0412_),
    .A1(\cla_z[18] ),
    .A2(net221));
 sg13g2_a21oi_2 _1258_ (.B1(_0412_),
    .Y(_0413_),
    .A2(_0411_),
    .A1(net221));
 sg13g2_nor2_1 _1259_ (.A(net218),
    .B(_0413_),
    .Y(_0414_));
 sg13g2_a21oi_1 _1260_ (.A1(_0134_),
    .A2(_0392_),
    .Y(_0415_),
    .B1(_0414_));
 sg13g2_a22oi_1 _1261_ (.Y(_0416_),
    .B1(_0415_),
    .B2(_0366_),
    .A2(_0410_),
    .A1(_0409_));
 sg13g2_o21ai_1 _1262_ (.B1(_0399_),
    .Y(_0062_),
    .A1(_0364_),
    .A2(_0416_));
 sg13g2_nand2_1 _1263_ (.Y(_0417_),
    .A(net148),
    .B(net210));
 sg13g2_xor2_1 _1264_ (.B(_0227_),
    .A(_0225_),
    .X(_0418_));
 sg13g2_a21oi_1 _1265_ (.A1(net224),
    .A2(_0418_),
    .Y(_0419_),
    .B1(_0372_));
 sg13g2_o21ai_1 _1266_ (.B1(_0419_),
    .Y(_0420_),
    .A1(\cla_z[11] ),
    .A2(net224));
 sg13g2_xor2_1 _1267_ (.B(_0205_),
    .A(_0203_),
    .X(_0421_));
 sg13g2_a21oi_1 _1268_ (.A1(net226),
    .A2(_0421_),
    .Y(_0422_),
    .B1(net192));
 sg13g2_o21ai_1 _1269_ (.B1(_0422_),
    .Y(_0423_),
    .A1(\cla_z[3] ),
    .A2(net226));
 sg13g2_nand2_1 _1270_ (.Y(_0424_),
    .A(net212),
    .B(_0423_));
 sg13g2_o21ai_1 _1271_ (.B1(_0424_),
    .Y(_0425_),
    .A1(net220),
    .A2(_0406_));
 sg13g2_a21oi_1 _1272_ (.A1(_0355_),
    .A2(_0425_),
    .Y(_0426_),
    .B1(_0368_));
 sg13g2_a22oi_1 _1273_ (.Y(_0427_),
    .B1(_0420_),
    .B2(_0354_),
    .A2(_0403_),
    .A1(_0359_));
 sg13g2_xor2_1 _1274_ (.B(_0251_),
    .A(_0249_),
    .X(_0428_));
 sg13g2_a21oi_1 _1275_ (.A1(net221),
    .A2(_0428_),
    .Y(_0429_),
    .B1(net192));
 sg13g2_o21ai_1 _1276_ (.B1(_0429_),
    .Y(_0430_),
    .A1(\cla_z[19] ),
    .A2(net221));
 sg13g2_nor2_1 _1277_ (.A(net219),
    .B(_0413_),
    .Y(_0431_));
 sg13g2_a21oi_1 _1278_ (.A1(net212),
    .A2(_0430_),
    .Y(_0432_),
    .B1(_0431_));
 sg13g2_a22oi_1 _1279_ (.Y(_0433_),
    .B1(_0432_),
    .B2(_0366_),
    .A2(_0427_),
    .A1(_0426_));
 sg13g2_o21ai_1 _1280_ (.B1(_0417_),
    .Y(_0063_),
    .A1(_0364_),
    .A2(_0433_));
 sg13g2_nand2_1 _1281_ (.Y(_0434_),
    .A(net157),
    .B(net210));
 sg13g2_xnor2_1 _1282_ (.Y(_0435_),
    .A(_0228_),
    .B(_0230_));
 sg13g2_o21ai_1 _1283_ (.B1(net191),
    .Y(_0436_),
    .A1(\cla_z[12] ),
    .A2(net224));
 sg13g2_a21oi_1 _1284_ (.A1(net224),
    .A2(_0435_),
    .Y(_0437_),
    .B1(_0436_));
 sg13g2_inv_1 _1285_ (.Y(_0438_),
    .A(_0437_));
 sg13g2_xnor2_1 _1286_ (.Y(_0439_),
    .A(_0206_),
    .B(_0208_));
 sg13g2_o21ai_1 _1287_ (.B1(net190),
    .Y(_0440_),
    .A1(\cla_z[4] ),
    .A2(net227));
 sg13g2_a21oi_1 _1288_ (.A1(net227),
    .A2(_0439_),
    .Y(_0441_),
    .B1(_0440_));
 sg13g2_and2_1 _1289_ (.A(net213),
    .B(_0441_),
    .X(_0442_));
 sg13g2_nor2_1 _1290_ (.A(net220),
    .B(_0423_),
    .Y(_0443_));
 sg13g2_nor3_1 _1291_ (.A(_0365_),
    .B(_0442_),
    .C(_0443_),
    .Y(_0444_));
 sg13g2_nor2_1 _1292_ (.A(_0368_),
    .B(_0444_),
    .Y(_0445_));
 sg13g2_a22oi_1 _1293_ (.Y(_0446_),
    .B1(_0438_),
    .B2(_0354_),
    .A2(_0420_),
    .A1(_0359_));
 sg13g2_xnor2_1 _1294_ (.Y(_0447_),
    .A(_0252_),
    .B(_0254_));
 sg13g2_o21ai_1 _1295_ (.B1(net190),
    .Y(_0448_),
    .A1(\cla_z[20] ),
    .A2(net221));
 sg13g2_a21oi_1 _1296_ (.A1(net221),
    .A2(_0447_),
    .Y(_0449_),
    .B1(_0448_));
 sg13g2_nor2_1 _1297_ (.A(net218),
    .B(_0449_),
    .Y(_0450_));
 sg13g2_a21oi_1 _1298_ (.A1(_0134_),
    .A2(_0430_),
    .Y(_0451_),
    .B1(_0450_));
 sg13g2_a22oi_1 _1299_ (.Y(_0452_),
    .B1(_0451_),
    .B2(_0366_),
    .A2(_0446_),
    .A1(_0445_));
 sg13g2_o21ai_1 _1300_ (.B1(_0434_),
    .Y(_0064_),
    .A1(_0364_),
    .A2(_0452_));
 sg13g2_nand2_1 _1301_ (.Y(_0453_),
    .A(net146),
    .B(net210));
 sg13g2_xor2_1 _1302_ (.B(_0233_),
    .A(_0231_),
    .X(_0454_));
 sg13g2_a21oi_1 _1303_ (.A1(net225),
    .A2(_0454_),
    .Y(_0455_),
    .B1(net192));
 sg13g2_o21ai_1 _1304_ (.B1(_0455_),
    .Y(_0456_),
    .A1(\cla_z[13] ),
    .A2(net225));
 sg13g2_xor2_1 _1305_ (.B(_0211_),
    .A(_0209_),
    .X(_0457_));
 sg13g2_a21oi_1 _1306_ (.A1(net227),
    .A2(_0457_),
    .Y(_0458_),
    .B1(net192));
 sg13g2_o21ai_1 _1307_ (.B1(_0458_),
    .Y(_0459_),
    .A1(\cla_z[5] ),
    .A2(net223));
 sg13g2_nand2_1 _1308_ (.Y(_0460_),
    .A(net212),
    .B(_0459_));
 sg13g2_o21ai_1 _1309_ (.B1(_0460_),
    .Y(_0461_),
    .A1(net220),
    .A2(_0441_));
 sg13g2_a21oi_1 _1310_ (.A1(_0355_),
    .A2(_0461_),
    .Y(_0462_),
    .B1(_0368_));
 sg13g2_a22oi_1 _1311_ (.Y(_0463_),
    .B1(_0456_),
    .B2(_0354_),
    .A2(_0438_),
    .A1(_0359_));
 sg13g2_xor2_1 _1312_ (.B(_0257_),
    .A(_0255_),
    .X(_0464_));
 sg13g2_a21oi_1 _1313_ (.A1(net223),
    .A2(_0464_),
    .Y(_0465_),
    .B1(net192));
 sg13g2_o21ai_1 _1314_ (.B1(_0465_),
    .Y(_0466_),
    .A1(\cla_z[21] ),
    .A2(net228));
 sg13g2_nor2_1 _1315_ (.A(net219),
    .B(_0449_),
    .Y(_0467_));
 sg13g2_a21oi_1 _1316_ (.A1(net212),
    .A2(_0466_),
    .Y(_0468_),
    .B1(_0467_));
 sg13g2_a22oi_1 _1317_ (.Y(_0469_),
    .B1(_0468_),
    .B2(_0366_),
    .A2(_0463_),
    .A1(_0462_));
 sg13g2_o21ai_1 _1318_ (.B1(_0453_),
    .Y(_0065_),
    .A1(_0364_),
    .A2(_0469_));
 sg13g2_nand2_1 _1319_ (.Y(_0470_),
    .A(net155),
    .B(net210));
 sg13g2_xnor2_1 _1320_ (.Y(_0471_),
    .A(_0234_),
    .B(_0236_));
 sg13g2_o21ai_1 _1321_ (.B1(net191),
    .Y(_0472_),
    .A1(\cla_z[14] ),
    .A2(net225));
 sg13g2_a21oi_2 _1322_ (.B1(_0472_),
    .Y(_0473_),
    .A2(_0471_),
    .A1(net225));
 sg13g2_nand2b_1 _1323_ (.Y(_0474_),
    .B(_0354_),
    .A_N(_0473_));
 sg13g2_xnor2_1 _1324_ (.Y(_0475_),
    .A(_0212_),
    .B(_0214_));
 sg13g2_o21ai_1 _1325_ (.B1(net190),
    .Y(_0476_),
    .A1(\cla_z[6] ),
    .A2(net227));
 sg13g2_a21oi_1 _1326_ (.A1(net227),
    .A2(_0475_),
    .Y(_0477_),
    .B1(_0476_));
 sg13g2_nand2_1 _1327_ (.Y(_0478_),
    .A(net213),
    .B(_0477_));
 sg13g2_nor2_1 _1328_ (.A(net219),
    .B(_0459_),
    .Y(_0479_));
 sg13g2_nor2_1 _1329_ (.A(_0365_),
    .B(_0479_),
    .Y(_0480_));
 sg13g2_a221oi_1 _1330_ (.B2(_0480_),
    .C1(_0368_),
    .B1(_0478_),
    .A1(_0359_),
    .Y(_0481_),
    .A2(_0456_));
 sg13g2_xnor2_1 _1331_ (.Y(_0482_),
    .A(_0258_),
    .B(_0260_));
 sg13g2_o21ai_1 _1332_ (.B1(net190),
    .Y(_0483_),
    .A1(\cla_z[22] ),
    .A2(net223));
 sg13g2_a21oi_1 _1333_ (.A1(net223),
    .A2(_0482_),
    .Y(_0484_),
    .B1(_0483_));
 sg13g2_nor2_1 _1334_ (.A(net218),
    .B(_0484_),
    .Y(_0485_));
 sg13g2_a21oi_1 _1335_ (.A1(_0134_),
    .A2(_0466_),
    .Y(_0486_),
    .B1(_0485_));
 sg13g2_a22oi_1 _1336_ (.Y(_0487_),
    .B1(_0486_),
    .B2(_0366_),
    .A2(_0481_),
    .A1(_0474_));
 sg13g2_o21ai_1 _1337_ (.B1(_0470_),
    .Y(_0066_),
    .A1(_0364_),
    .A2(_0487_));
 sg13g2_nand2_1 _1338_ (.Y(_0488_),
    .A(net145),
    .B(net210));
 sg13g2_xnor2_1 _1339_ (.Y(_0489_),
    .A(_0261_),
    .B(_0262_));
 sg13g2_o21ai_1 _1340_ (.B1(net190),
    .Y(_0490_),
    .A1(\cla_z[23] ),
    .A2(net223));
 sg13g2_a21oi_1 _1341_ (.A1(net223),
    .A2(_0489_),
    .Y(_0491_),
    .B1(_0490_));
 sg13g2_or2_1 _1342_ (.X(_0492_),
    .B(_0491_),
    .A(\io_sd._209_[0] ));
 sg13g2_o21ai_1 _1343_ (.B1(_0366_),
    .Y(_0493_),
    .A1(net219),
    .A2(_0484_));
 sg13g2_inv_1 _1344_ (.Y(_0494_),
    .A(_0493_));
 sg13g2_xor2_1 _1345_ (.B(_0239_),
    .A(_0237_),
    .X(_0495_));
 sg13g2_o21ai_1 _1346_ (.B1(net190),
    .Y(_0496_),
    .A1(\cla_z[15] ),
    .A2(net222));
 sg13g2_a21oi_2 _1347_ (.B1(_0496_),
    .Y(_0497_),
    .A2(_0495_),
    .A1(net222));
 sg13g2_nor2_1 _1348_ (.A(_0355_),
    .B(_0497_),
    .Y(_0498_));
 sg13g2_xor2_1 _1349_ (.B(_0217_),
    .A(_0215_),
    .X(_0499_));
 sg13g2_o21ai_1 _1350_ (.B1(net190),
    .Y(_0500_),
    .A1(\cla_z[7] ),
    .A2(net227));
 sg13g2_a21oi_1 _1351_ (.A1(net227),
    .A2(_0499_),
    .Y(_0501_),
    .B1(_0500_));
 sg13g2_nor2_1 _1352_ (.A(_0134_),
    .B(_0501_),
    .Y(_0502_));
 sg13g2_nor2_1 _1353_ (.A(net213),
    .B(_0477_),
    .Y(_0503_));
 sg13g2_o21ai_1 _1354_ (.B1(_0360_),
    .Y(_0504_),
    .A1(_0502_),
    .A2(_0503_));
 sg13g2_nor2_1 _1355_ (.A(_0360_),
    .B(_0473_),
    .Y(_0505_));
 sg13g2_nor3_1 _1356_ (.A(_0368_),
    .B(_0498_),
    .C(_0505_),
    .Y(_0506_));
 sg13g2_a22oi_1 _1357_ (.Y(_0507_),
    .B1(_0504_),
    .B2(_0506_),
    .A2(_0494_),
    .A1(_0492_));
 sg13g2_o21ai_1 _1358_ (.B1(_0488_),
    .Y(_0067_),
    .A1(_0364_),
    .A2(_0507_));
 sg13g2_or2_1 _1359_ (.X(_0508_),
    .B(_0396_),
    .A(_0355_));
 sg13g2_or2_1 _1360_ (.X(_0509_),
    .B(_0387_),
    .A(net218));
 sg13g2_nor2_1 _1361_ (.A(net219),
    .B(_0501_),
    .Y(_0510_));
 sg13g2_nor2_1 _1362_ (.A(_0365_),
    .B(_0510_),
    .Y(_0511_));
 sg13g2_a22oi_1 _1363_ (.Y(_0512_),
    .B1(_0509_),
    .B2(_0511_),
    .A2(_0497_),
    .A1(_0359_));
 sg13g2_a21oi_1 _1364_ (.A1(_0508_),
    .A2(_0512_),
    .Y(_0513_),
    .B1(_0368_));
 sg13g2_nor2_1 _1365_ (.A(net287),
    .B(_0367_),
    .Y(_0514_));
 sg13g2_a21oi_1 _1366_ (.A1(_0491_),
    .A2(_0514_),
    .Y(_0515_),
    .B1(_0513_));
 sg13g2_nor4_1 _1367_ (.A(net218),
    .B(_0138_),
    .C(_0363_),
    .D(_0382_),
    .Y(_0516_));
 sg13g2_a21oi_1 _1368_ (.A1(\io_sd.outputs[7] ),
    .A2(net210),
    .Y(_0517_),
    .B1(_0516_));
 sg13g2_o21ai_1 _1369_ (.B1(_0517_),
    .Y(_0068_),
    .A1(_0364_),
    .A2(_0515_));
 sg13g2_nand2b_2 _1370_ (.Y(_0518_),
    .B(net215),
    .A_N(net217));
 sg13g2_nand2_2 _1371_ (.Y(_0519_),
    .A(_0011_),
    .B(_0014_));
 sg13g2_nor2_2 _1372_ (.A(_0518_),
    .B(_0519_),
    .Y(_0520_));
 sg13g2_nand2_1 _1373_ (.Y(_0521_),
    .A(net202),
    .B(_0520_));
 sg13g2_nand2_1 _1374_ (.Y(_0522_),
    .A(net2),
    .B(_0520_));
 sg13g2_nor2_2 _1375_ (.A(net215),
    .B(net217),
    .Y(_0523_));
 sg13g2_nand2_1 _1376_ (.Y(_0524_),
    .A(_0011_),
    .B(_0523_));
 sg13g2_o21ai_1 _1377_ (.B1(_0011_),
    .Y(_0525_),
    .A1(_0014_),
    .A2(_0523_));
 sg13g2_a21oi_1 _1378_ (.A1(_0014_),
    .A2(_0523_),
    .Y(_0526_),
    .B1(_0525_));
 sg13g2_nand2_1 _1379_ (.Y(_0527_),
    .A(_0518_),
    .B(_0526_));
 sg13g2_inv_1 _1380_ (.Y(_0528_),
    .A(net196));
 sg13g2_nand2_1 _1381_ (.Y(_0529_),
    .A(net215),
    .B(net217));
 sg13g2_nor2b_2 _1382_ (.A(_0523_),
    .B_N(_0529_),
    .Y(_0530_));
 sg13g2_inv_1 _1383_ (.Y(_0531_),
    .A(net199));
 sg13g2_nand4_1 _1384_ (.B(\io_sd.input_index[5] ),
    .C(\io_sd.input_index[4] ),
    .A(net215),
    .Y(_0532_),
    .D(net217));
 sg13g2_nand2b_1 _1385_ (.Y(_0533_),
    .B(_0011_),
    .A_N(_0014_));
 sg13g2_o21ai_1 _1386_ (.B1(_0524_),
    .Y(_0534_),
    .A1(_0014_),
    .A2(_0529_));
 sg13g2_and2_1 _1387_ (.A(_0533_),
    .B(_0534_),
    .X(_0535_));
 sg13g2_xor2_1 _1388_ (.B(_0535_),
    .A(_0532_),
    .X(_0536_));
 sg13g2_nor2b_1 _1389_ (.A(_0015_),
    .B_N(_0536_),
    .Y(_0537_));
 sg13g2_nand2_1 _1390_ (.Y(_0538_),
    .A(net2),
    .B(_0537_));
 sg13g2_nand3_1 _1391_ (.B(_0530_),
    .C(_0537_),
    .A(net2),
    .Y(_0539_));
 sg13g2_o21ai_1 _1392_ (.B1(_0522_),
    .Y(_0540_),
    .A1(_0527_),
    .A2(_0539_));
 sg13g2_a22oi_1 _1393_ (.Y(_0541_),
    .B1(_0540_),
    .B2(net202),
    .A2(_0521_),
    .A1(net302));
 sg13g2_nor2_1 _1394_ (.A(net236),
    .B(_0541_),
    .Y(_0069_));
 sg13g2_nor2b_1 _1395_ (.A(net217),
    .B_N(_0015_),
    .Y(_0542_));
 sg13g2_nor3_2 _1396_ (.A(_0519_),
    .B(_0531_),
    .C(_0542_),
    .Y(_0543_));
 sg13g2_nand2_2 _1397_ (.Y(_0544_),
    .A(net203),
    .B(_0543_));
 sg13g2_nand2_1 _1398_ (.Y(_0545_),
    .A(net3),
    .B(_0520_));
 sg13g2_mux2_1 _1399_ (.A0(net2),
    .A1(net3),
    .S(net216),
    .X(_0546_));
 sg13g2_nand2_1 _1400_ (.Y(_0547_),
    .A(net199),
    .B(_0546_));
 sg13g2_o21ai_1 _1401_ (.B1(_0545_),
    .Y(_0548_),
    .A1(net196),
    .A2(_0547_));
 sg13g2_a22oi_1 _1402_ (.Y(_0549_),
    .B1(_0548_),
    .B2(net202),
    .A2(_0544_),
    .A1(net322));
 sg13g2_nor2_1 _1403_ (.A(net236),
    .B(_0549_),
    .Y(_0070_));
 sg13g2_nand2_1 _1404_ (.Y(_0550_),
    .A(net4),
    .B(_0520_));
 sg13g2_mux2_1 _1405_ (.A0(net3),
    .A1(net4),
    .S(net216),
    .X(_0551_));
 sg13g2_nand2_1 _1406_ (.Y(_0552_),
    .A(net199),
    .B(_0551_));
 sg13g2_o21ai_1 _1407_ (.B1(_0550_),
    .Y(_0553_),
    .A1(net196),
    .A2(_0552_));
 sg13g2_a22oi_1 _1408_ (.Y(_0554_),
    .B1(_0553_),
    .B2(net202),
    .A2(_0544_),
    .A1(net304));
 sg13g2_nor2_1 _1409_ (.A(net236),
    .B(_0554_),
    .Y(_0071_));
 sg13g2_nand2_1 _1410_ (.Y(_0555_),
    .A(net5),
    .B(_0520_));
 sg13g2_mux2_1 _1411_ (.A0(net4),
    .A1(net5),
    .S(net216),
    .X(_0556_));
 sg13g2_nand2_1 _1412_ (.Y(_0557_),
    .A(net199),
    .B(_0556_));
 sg13g2_o21ai_1 _1413_ (.B1(_0555_),
    .Y(_0558_),
    .A1(net196),
    .A2(_0557_));
 sg13g2_a22oi_1 _1414_ (.Y(_0559_),
    .B1(_0558_),
    .B2(net200),
    .A2(_0544_),
    .A1(net268));
 sg13g2_nor2_1 _1415_ (.A(net233),
    .B(_0559_),
    .Y(_0072_));
 sg13g2_mux2_1 _1416_ (.A0(net5),
    .A1(net6),
    .S(net216),
    .X(_0560_));
 sg13g2_nand2_1 _1417_ (.Y(_0561_),
    .A(net199),
    .B(_0560_));
 sg13g2_nor3_2 _1418_ (.A(_0015_),
    .B(_0518_),
    .C(_0519_),
    .Y(_0562_));
 sg13g2_nand2_1 _1419_ (.Y(_0563_),
    .A(net6),
    .B(_0562_));
 sg13g2_o21ai_1 _1420_ (.B1(_0563_),
    .Y(_0564_),
    .A1(net196),
    .A2(_0561_));
 sg13g2_a22oi_1 _1421_ (.Y(_0565_),
    .B1(_0564_),
    .B2(net201),
    .A2(_0544_),
    .A1(net272));
 sg13g2_nor2_1 _1422_ (.A(net233),
    .B(net273),
    .Y(_0073_));
 sg13g2_nand2_1 _1423_ (.Y(_0566_),
    .A(net7),
    .B(_0562_));
 sg13g2_mux2_1 _1424_ (.A0(net6),
    .A1(net7),
    .S(net216),
    .X(_0567_));
 sg13g2_nand2_1 _1425_ (.Y(_0568_),
    .A(net199),
    .B(_0567_));
 sg13g2_o21ai_1 _1426_ (.B1(_0566_),
    .Y(_0569_),
    .A1(net196),
    .A2(_0568_));
 sg13g2_a22oi_1 _1427_ (.Y(_0570_),
    .B1(_0569_),
    .B2(net200),
    .A2(_0544_),
    .A1(net314));
 sg13g2_nor2_1 _1428_ (.A(net233),
    .B(net315),
    .Y(_0074_));
 sg13g2_nand2_1 _1429_ (.Y(_0571_),
    .A(net8),
    .B(_0562_));
 sg13g2_mux2_1 _1430_ (.A0(net7),
    .A1(net8),
    .S(net216),
    .X(_0572_));
 sg13g2_nand2_1 _1431_ (.Y(_0573_),
    .A(net199),
    .B(_0572_));
 sg13g2_o21ai_1 _1432_ (.B1(_0571_),
    .Y(_0574_),
    .A1(net196),
    .A2(_0573_));
 sg13g2_a22oi_1 _1433_ (.Y(_0575_),
    .B1(_0574_),
    .B2(net203),
    .A2(_0544_),
    .A1(net291));
 sg13g2_nor2_1 _1434_ (.A(net235),
    .B(_0575_),
    .Y(_0075_));
 sg13g2_nand2_1 _1435_ (.Y(_0576_),
    .A(net9),
    .B(_0562_));
 sg13g2_nor2_1 _1436_ (.A(net215),
    .B(net8),
    .Y(_0577_));
 sg13g2_a21oi_2 _1437_ (.B1(_0577_),
    .Y(_0578_),
    .A2(_0137_),
    .A1(net215));
 sg13g2_nand2_1 _1438_ (.Y(_0579_),
    .A(_0530_),
    .B(_0578_));
 sg13g2_o21ai_1 _1439_ (.B1(_0576_),
    .Y(_0580_),
    .A1(net196),
    .A2(_0579_));
 sg13g2_a22oi_1 _1440_ (.Y(_0581_),
    .B1(_0580_),
    .B2(net203),
    .A2(_0544_),
    .A1(net250));
 sg13g2_nor2_1 _1441_ (.A(net235),
    .B(_0581_),
    .Y(_0076_));
 sg13g2_o21ai_1 _1442_ (.B1(_0528_),
    .Y(_0582_),
    .A1(net199),
    .A2(_0537_));
 sg13g2_o21ai_1 _1443_ (.B1(net299),
    .Y(_0583_),
    .A1(_0343_),
    .A2(_0582_));
 sg13g2_nor3_1 _1444_ (.A(net215),
    .B(_0137_),
    .C(_0535_),
    .Y(_0584_));
 sg13g2_nand2_1 _1445_ (.Y(_0585_),
    .A(net217),
    .B(_0584_));
 sg13g2_o21ai_1 _1446_ (.B1(_0585_),
    .Y(_0586_),
    .A1(_0530_),
    .A2(_0538_));
 sg13g2_nand3_1 _1447_ (.B(_0528_),
    .C(_0586_),
    .A(net202),
    .Y(_0587_));
 sg13g2_a21oi_1 _1448_ (.A1(net300),
    .A2(_0587_),
    .Y(_0077_),
    .B1(net235));
 sg13g2_and2_2 _1449_ (.A(_0526_),
    .B(_0531_),
    .X(_0588_));
 sg13g2_nand2_2 _1450_ (.Y(_0589_),
    .A(_0536_),
    .B(_0588_));
 sg13g2_nand3_1 _1451_ (.B(_0536_),
    .C(_0588_),
    .A(net200),
    .Y(_0590_));
 sg13g2_nor2b_1 _1452_ (.A(_0589_),
    .B_N(_0546_),
    .Y(_0591_));
 sg13g2_a22oi_1 _1453_ (.Y(_0592_),
    .B1(_0591_),
    .B2(net200),
    .A2(_0590_),
    .A1(net264));
 sg13g2_nor2_1 _1454_ (.A(net232),
    .B(_0592_),
    .Y(_0078_));
 sg13g2_nor2b_1 _1455_ (.A(_0589_),
    .B_N(_0551_),
    .Y(_0593_));
 sg13g2_a22oi_1 _1456_ (.Y(_0594_),
    .B1(_0593_),
    .B2(net200),
    .A2(_0590_),
    .A1(net178));
 sg13g2_nor2_1 _1457_ (.A(net232),
    .B(_0594_),
    .Y(_0079_));
 sg13g2_nor2b_1 _1458_ (.A(_0589_),
    .B_N(_0556_),
    .Y(_0595_));
 sg13g2_a22oi_1 _1459_ (.Y(_0596_),
    .B1(_0595_),
    .B2(net200),
    .A2(_0590_),
    .A1(net179));
 sg13g2_nor2_1 _1460_ (.A(net232),
    .B(_0596_),
    .Y(_0080_));
 sg13g2_nor2b_1 _1461_ (.A(_0589_),
    .B_N(_0560_),
    .Y(_0597_));
 sg13g2_a22oi_1 _1462_ (.Y(_0598_),
    .B1(_0597_),
    .B2(net200),
    .A2(_0590_),
    .A1(net254));
 sg13g2_nor2_1 _1463_ (.A(net232),
    .B(_0598_),
    .Y(_0081_));
 sg13g2_nor2b_1 _1464_ (.A(_0589_),
    .B_N(_0567_),
    .Y(_0599_));
 sg13g2_a22oi_1 _1465_ (.Y(_0600_),
    .B1(_0599_),
    .B2(net200),
    .A2(_0590_),
    .A1(net266));
 sg13g2_nor2_1 _1466_ (.A(net234),
    .B(_0600_),
    .Y(_0082_));
 sg13g2_nor2b_1 _1467_ (.A(_0589_),
    .B_N(_0572_),
    .Y(_0601_));
 sg13g2_a22oi_1 _1468_ (.Y(_0602_),
    .B1(_0601_),
    .B2(net201),
    .A2(_0590_),
    .A1(net267));
 sg13g2_nor2_1 _1469_ (.A(net234),
    .B(_0602_),
    .Y(_0083_));
 sg13g2_nor2b_1 _1470_ (.A(_0589_),
    .B_N(_0578_),
    .Y(_0603_));
 sg13g2_a22oi_1 _1471_ (.Y(_0604_),
    .B1(_0603_),
    .B2(net201),
    .A2(_0590_),
    .A1(net181));
 sg13g2_nor2_1 _1472_ (.A(net234),
    .B(_0604_),
    .Y(_0084_));
 sg13g2_nor2_1 _1473_ (.A(net217),
    .B(_0533_),
    .Y(_0605_));
 sg13g2_nand2_1 _1474_ (.Y(_0606_),
    .A(net203),
    .B(_0605_));
 sg13g2_a21oi_1 _1475_ (.A1(_0014_),
    .A2(_0523_),
    .Y(_0607_),
    .B1(_0011_));
 sg13g2_nor2b_1 _1476_ (.A(_0607_),
    .B_N(_0525_),
    .Y(_0608_));
 sg13g2_inv_4 _1477_ (.A(_0608_),
    .Y(_0609_));
 sg13g2_nand2_1 _1478_ (.Y(_0610_),
    .A(_0584_),
    .B(_0588_));
 sg13g2_o21ai_1 _1479_ (.B1(_0610_),
    .Y(_0611_),
    .A1(_0539_),
    .A2(_0609_));
 sg13g2_a22oi_1 _1480_ (.Y(_0612_),
    .B1(_0611_),
    .B2(net203),
    .A2(_0606_),
    .A1(net324));
 sg13g2_nor2_1 _1481_ (.A(net235),
    .B(_0612_),
    .Y(_0085_));
 sg13g2_nor2_2 _1482_ (.A(_0531_),
    .B(_0533_),
    .Y(_0613_));
 sg13g2_nand2_2 _1483_ (.Y(_0614_),
    .A(net204),
    .B(_0613_));
 sg13g2_nor2_2 _1484_ (.A(_0547_),
    .B(_0609_),
    .Y(_0615_));
 sg13g2_a22oi_1 _1485_ (.Y(_0616_),
    .B1(_0615_),
    .B2(net204),
    .A2(_0614_),
    .A1(net278));
 sg13g2_nor2_1 _1486_ (.A(net229),
    .B(_0616_),
    .Y(_0086_));
 sg13g2_nor2_2 _1487_ (.A(_0552_),
    .B(_0609_),
    .Y(_0617_));
 sg13g2_a22oi_1 _1488_ (.Y(_0618_),
    .B1(_0617_),
    .B2(net204),
    .A2(_0614_),
    .A1(net186));
 sg13g2_nor2_1 _1489_ (.A(net229),
    .B(_0618_),
    .Y(_0087_));
 sg13g2_nor2_2 _1490_ (.A(_0557_),
    .B(_0609_),
    .Y(_0619_));
 sg13g2_a22oi_1 _1491_ (.Y(_0620_),
    .B1(_0619_),
    .B2(net204),
    .A2(_0614_),
    .A1(net180));
 sg13g2_nor2_1 _1492_ (.A(net229),
    .B(_0620_),
    .Y(_0088_));
 sg13g2_nor2_2 _1493_ (.A(_0561_),
    .B(_0609_),
    .Y(_0621_));
 sg13g2_a22oi_1 _1494_ (.Y(_0622_),
    .B1(_0621_),
    .B2(net204),
    .A2(_0614_),
    .A1(net177));
 sg13g2_nor2_1 _1495_ (.A(net230),
    .B(_0622_),
    .Y(_0089_));
 sg13g2_nor2_2 _1496_ (.A(_0568_),
    .B(_0609_),
    .Y(_0623_));
 sg13g2_a22oi_1 _1497_ (.Y(_0624_),
    .B1(_0623_),
    .B2(net204),
    .A2(_0614_),
    .A1(net183));
 sg13g2_nor2_1 _1498_ (.A(net229),
    .B(_0624_),
    .Y(_0090_));
 sg13g2_nor2_2 _1499_ (.A(_0573_),
    .B(_0609_),
    .Y(_0625_));
 sg13g2_a22oi_1 _1500_ (.Y(_0626_),
    .B1(_0625_),
    .B2(net204),
    .A2(_0614_),
    .A1(net170));
 sg13g2_nor2_1 _1501_ (.A(net231),
    .B(_0626_),
    .Y(_0091_));
 sg13g2_nor2_2 _1502_ (.A(_0579_),
    .B(_0609_),
    .Y(_0627_));
 sg13g2_a22oi_1 _1503_ (.Y(_0628_),
    .B1(_0627_),
    .B2(net204),
    .A2(_0614_),
    .A1(net189));
 sg13g2_nor2_1 _1504_ (.A(net231),
    .B(_0628_),
    .Y(_0092_));
 sg13g2_nand2_1 _1505_ (.Y(_0629_),
    .A(net206),
    .B(_0520_));
 sg13g2_a22oi_1 _1506_ (.Y(_0630_),
    .B1(_0629_),
    .B2(net187),
    .A2(_0540_),
    .A1(net206));
 sg13g2_nor2_1 _1507_ (.A(net237),
    .B(_0630_),
    .Y(_0093_));
 sg13g2_nand2_2 _1508_ (.Y(_0631_),
    .A(net206),
    .B(_0543_));
 sg13g2_a22oi_1 _1509_ (.Y(_0632_),
    .B1(_0631_),
    .B2(net308),
    .A2(_0548_),
    .A1(net206));
 sg13g2_nor2_1 _1510_ (.A(net236),
    .B(_0632_),
    .Y(_0094_));
 sg13g2_a22oi_1 _1511_ (.Y(_0633_),
    .B1(_0631_),
    .B2(net319),
    .A2(_0553_),
    .A1(net206));
 sg13g2_nor2_1 _1512_ (.A(net236),
    .B(_0633_),
    .Y(_0095_));
 sg13g2_a22oi_1 _1513_ (.Y(_0634_),
    .B1(_0631_),
    .B2(net286),
    .A2(_0558_),
    .A1(net205));
 sg13g2_nor2_1 _1514_ (.A(net233),
    .B(_0634_),
    .Y(_0096_));
 sg13g2_a22oi_1 _1515_ (.Y(_0635_),
    .B1(_0631_),
    .B2(net289),
    .A2(_0564_),
    .A1(net205));
 sg13g2_nor2_1 _1516_ (.A(net233),
    .B(_0635_),
    .Y(_0097_));
 sg13g2_a22oi_1 _1517_ (.Y(_0636_),
    .B1(_0631_),
    .B2(net320),
    .A2(_0569_),
    .A1(net205));
 sg13g2_nor2_1 _1518_ (.A(net233),
    .B(net321),
    .Y(_0098_));
 sg13g2_a22oi_1 _1519_ (.Y(_0637_),
    .B1(_0631_),
    .B2(net283),
    .A2(_0574_),
    .A1(net207));
 sg13g2_nor2_1 _1520_ (.A(net235),
    .B(_0637_),
    .Y(_0099_));
 sg13g2_a22oi_1 _1521_ (.Y(_0638_),
    .B1(_0631_),
    .B2(net290),
    .A2(_0580_),
    .A1(net207));
 sg13g2_nor2_1 _1522_ (.A(net235),
    .B(_0638_),
    .Y(_0100_));
 sg13g2_o21ai_1 _1523_ (.B1(net333),
    .Y(_0639_),
    .A1(_0345_),
    .A2(_0582_));
 sg13g2_nand3_1 _1524_ (.B(_0528_),
    .C(_0586_),
    .A(net207),
    .Y(_0640_));
 sg13g2_a21oi_1 _1525_ (.A1(_0639_),
    .A2(_0640_),
    .Y(_0101_),
    .B1(net235));
 sg13g2_nand3_1 _1526_ (.B(_0536_),
    .C(_0588_),
    .A(net205),
    .Y(_0641_));
 sg13g2_a22oi_1 _1527_ (.Y(_0642_),
    .B1(_0641_),
    .B2(net274),
    .A2(_0591_),
    .A1(net208));
 sg13g2_nor2_1 _1528_ (.A(net232),
    .B(_0642_),
    .Y(_0102_));
 sg13g2_a22oi_1 _1529_ (.Y(_0643_),
    .B1(_0641_),
    .B2(net188),
    .A2(_0593_),
    .A1(net208));
 sg13g2_nor2_1 _1530_ (.A(net232),
    .B(_0643_),
    .Y(_0103_));
 sg13g2_a22oi_1 _1531_ (.Y(_0644_),
    .B1(_0641_),
    .B2(net276),
    .A2(_0595_),
    .A1(net208));
 sg13g2_nor2_1 _1532_ (.A(net232),
    .B(_0644_),
    .Y(_0104_));
 sg13g2_a22oi_1 _1533_ (.Y(_0645_),
    .B1(_0641_),
    .B2(net282),
    .A2(_0597_),
    .A1(net205));
 sg13g2_nor2_1 _1534_ (.A(net232),
    .B(_0645_),
    .Y(_0105_));
 sg13g2_a22oi_1 _1535_ (.Y(_0646_),
    .B1(_0641_),
    .B2(net305),
    .A2(_0599_),
    .A1(net205));
 sg13g2_nor2_1 _1536_ (.A(net234),
    .B(_0646_),
    .Y(_0106_));
 sg13g2_a22oi_1 _1537_ (.Y(_0118_),
    .B1(_0641_),
    .B2(net284),
    .A2(_0601_),
    .A1(net205));
 sg13g2_nor2_1 _1538_ (.A(net234),
    .B(_0118_),
    .Y(_0107_));
 sg13g2_a22oi_1 _1539_ (.Y(_0119_),
    .B1(_0641_),
    .B2(net342),
    .A2(_0603_),
    .A1(net205));
 sg13g2_nor2_1 _1540_ (.A(net230),
    .B(_0119_),
    .Y(_0108_));
 sg13g2_nand2_1 _1541_ (.Y(_0120_),
    .A(net207),
    .B(_0605_));
 sg13g2_a22oi_1 _1542_ (.Y(_0121_),
    .B1(_0120_),
    .B2(net341),
    .A2(_0611_),
    .A1(net207));
 sg13g2_nor2_1 _1543_ (.A(net237),
    .B(_0121_),
    .Y(_0109_));
 sg13g2_nand2_2 _1544_ (.Y(_0122_),
    .A(net209),
    .B(_0613_));
 sg13g2_a22oi_1 _1545_ (.Y(_0123_),
    .B1(_0122_),
    .B2(net285),
    .A2(_0615_),
    .A1(net209));
 sg13g2_nor2_1 _1546_ (.A(net229),
    .B(_0123_),
    .Y(_0110_));
 sg13g2_a22oi_1 _1547_ (.Y(_0124_),
    .B1(_0122_),
    .B2(net275),
    .A2(_0617_),
    .A1(net209));
 sg13g2_nor2_1 _1548_ (.A(net229),
    .B(_0124_),
    .Y(_0111_));
 sg13g2_a22oi_1 _1549_ (.Y(_0125_),
    .B1(_0122_),
    .B2(net255),
    .A2(_0619_),
    .A1(net209));
 sg13g2_nor2_1 _1550_ (.A(net229),
    .B(_0125_),
    .Y(_0112_));
 sg13g2_a22oi_1 _1551_ (.Y(_0126_),
    .B1(_0122_),
    .B2(net256),
    .A2(_0621_),
    .A1(net209));
 sg13g2_nor2_1 _1552_ (.A(net230),
    .B(_0126_),
    .Y(_0113_));
 sg13g2_a22oi_1 _1553_ (.Y(_0127_),
    .B1(_0122_),
    .B2(net294),
    .A2(_0623_),
    .A1(net209));
 sg13g2_nor2_1 _1554_ (.A(net229),
    .B(_0127_),
    .Y(_0114_));
 sg13g2_a22oi_1 _1555_ (.Y(_0128_),
    .B1(_0122_),
    .B2(net265),
    .A2(_0625_),
    .A1(net209));
 sg13g2_nor2_1 _1556_ (.A(net231),
    .B(_0128_),
    .Y(_0115_));
 sg13g2_a22oi_1 _1557_ (.Y(_0129_),
    .B1(_0122_),
    .B2(net171),
    .A2(_0627_),
    .A1(net209));
 sg13g2_nor2_1 _1558_ (.A(net231),
    .B(_0129_),
    .Y(_0116_));
 sg13g2_nor2_1 _1559_ (.A(net215),
    .B(net236),
    .Y(_0130_));
 sg13g2_o21ai_1 _1560_ (.B1(_0130_),
    .Y(_0117_),
    .A1(_0146_),
    .A2(_0346_));
 sg13g2_dfrbp_1 _1561_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net34),
    .D(_0016_),
    .Q_N(_0741_),
    .Q(\io_sd.output_index[3] ));
 sg13g2_dfrbp_1 _1562_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net28),
    .D(_0017_),
    .Q_N(_0013_),
    .Q(\io_sd.output_index[4] ));
 sg13g2_dfrbp_1 _1563_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net26),
    .D(net293),
    .Q_N(_0010_),
    .Q(\io_sd.output_index[5] ));
 sg13g2_dfrbp_1 _1564_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net130),
    .D(_0019_),
    .Q_N(_0740_),
    .Q(\bav1.x[0] ));
 sg13g2_dfrbp_1 _1565_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net129),
    .D(_0020_),
    .Q_N(_0739_),
    .Q(\bav1.x[1] ));
 sg13g2_dfrbp_1 _1566_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net128),
    .D(_0021_),
    .Q_N(_0738_),
    .Q(\ca.coin_out[2] ));
 sg13g2_dfrbp_1 _1567_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net127),
    .D(_0022_),
    .Q_N(_0737_),
    .Q(\ca.coin_out[3] ));
 sg13g2_dfrbp_1 _1568_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net126),
    .D(_0023_),
    .Q_N(_0736_),
    .Q(\ca.coin_out[4] ));
 sg13g2_dfrbp_1 _1569_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net35),
    .D(_0024_),
    .Q_N(_0742_),
    .Q(\ca.coin_out[5] ));
 sg13g2_dfrbp_1 _1570_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net36),
    .D(_0006_),
    .Q_N(_0743_),
    .Q(\bav0.state_q[0] ));
 sg13g2_dfrbp_1 _1571_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net37),
    .D(net176),
    .Q_N(_0744_),
    .Q(\bav0.state_q[1] ));
 sg13g2_dfrbp_1 _1572_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net131),
    .D(_0008_),
    .Q_N(_0745_),
    .Q(\bav0.state_q[2] ));
 sg13g2_dfrbp_1 _1573_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net125),
    .D(net168),
    .Q_N(_0735_),
    .Q(\bav0._02_ ));
 sg13g2_dfrbp_1 _1574_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net124),
    .D(_0025_),
    .Q_N(_0012_),
    .Q(\io_sd._209_[0] ));
 sg13g2_dfrbp_1 _1575_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net122),
    .D(_0026_),
    .Q_N(_0734_),
    .Q(\ca._11_ ));
 sg13g2_dfrbp_1 _1576_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net121),
    .D(_0027_),
    .Q_N(\ca._08_[0] ),
    .Q(\ca.commit_count[0] ));
 sg13g2_dfrbp_1 _1577_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net119),
    .D(net166),
    .Q_N(_0733_),
    .Q(\ca.commit_count[1] ));
 sg13g2_dfrbp_1 _1578_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net117),
    .D(_0029_),
    .Q_N(_0732_),
    .Q(\ca.commit_count[2] ));
 sg13g2_dfrbp_1 _1579_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net115),
    .D(_0030_),
    .Q_N(_0731_),
    .Q(\ca.commit_count[3] ));
 sg13g2_dfrbp_1 _1580_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net113),
    .D(_0031_),
    .Q_N(_0730_),
    .Q(\ca.commit_count[4] ));
 sg13g2_dfrbp_1 _1581_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net111),
    .D(_0032_),
    .Q_N(_0729_),
    .Q(\ca.commit_count[5] ));
 sg13g2_dfrbp_1 _1582_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net109),
    .D(_0033_),
    .Q_N(_0728_),
    .Q(\ca.commit_count[6] ));
 sg13g2_dfrbp_1 _1583_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net107),
    .D(_0034_),
    .Q_N(_0727_),
    .Q(\ca.commit_count[7] ));
 sg13g2_dfrbp_1 _1584_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net105),
    .D(_0035_),
    .Q_N(_0726_),
    .Q(\ca.commit_count[8] ));
 sg13g2_dfrbp_1 _1585_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net103),
    .D(net174),
    .Q_N(_0725_),
    .Q(\ca.commit_count[9] ));
 sg13g2_dfrbp_1 _1586_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net101),
    .D(_0037_),
    .Q_N(_0724_),
    .Q(\ca.commit_count[10] ));
 sg13g2_dfrbp_1 _1587_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net99),
    .D(_0038_),
    .Q_N(_0723_),
    .Q(\ca.commit_count[11] ));
 sg13g2_dfrbp_1 _1588_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net97),
    .D(_0039_),
    .Q_N(_0722_),
    .Q(\ca.commit_count[12] ));
 sg13g2_dfrbp_1 _1589_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net95),
    .D(_0040_),
    .Q_N(_0721_),
    .Q(\ca.commit_count[13] ));
 sg13g2_dfrbp_1 _1590_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net93),
    .D(_0041_),
    .Q_N(_0720_),
    .Q(\ca.commit_count[14] ));
 sg13g2_dfrbp_1 _1591_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net91),
    .D(_0042_),
    .Q_N(_0719_),
    .Q(\ca.commit_count[15] ));
 sg13g2_dfrbp_1 _1592_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net89),
    .D(_0043_),
    .Q_N(_0718_),
    .Q(\ca.commit_count[16] ));
 sg13g2_dfrbp_1 _1593_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net87),
    .D(net311),
    .Q_N(_0717_),
    .Q(\ca.commit_count[17] ));
 sg13g2_dfrbp_1 _1594_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net85),
    .D(net298),
    .Q_N(_0716_),
    .Q(\ca.commit_count[18] ));
 sg13g2_dfrbp_1 _1595_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net83),
    .D(net259),
    .Q_N(_0715_),
    .Q(\ca.commit_count[19] ));
 sg13g2_dfrbp_1 _1596_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net81),
    .D(_0047_),
    .Q_N(_0714_),
    .Q(\ca.commit_count[20] ));
 sg13g2_dfrbp_1 _1597_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net79),
    .D(_0048_),
    .Q_N(_0713_),
    .Q(\ca.commit_count[21] ));
 sg13g2_dfrbp_1 _1598_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net77),
    .D(_0049_),
    .Q_N(_0712_),
    .Q(\ca._15_ ));
 sg13g2_dfrbp_1 _1599_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net75),
    .D(_0050_),
    .Q_N(\ca._07_[0] ),
    .Q(\ca.pulse_count[0] ));
 sg13g2_dfrbp_1 _1600_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net73),
    .D(_0051_),
    .Q_N(_0711_),
    .Q(\ca.pulse_count[1] ));
 sg13g2_dfrbp_1 _1601_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net71),
    .D(_0052_),
    .Q_N(_0710_),
    .Q(\ca.pulse_count[2] ));
 sg13g2_dfrbp_1 _1602_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net69),
    .D(_0053_),
    .Q_N(_0709_),
    .Q(\ca.pulse_count[3] ));
 sg13g2_dfrbp_1 _1603_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net67),
    .D(_0054_),
    .Q_N(_0708_),
    .Q(\ca.pulse_count[4] ));
 sg13g2_dfrbp_1 _1604_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net65),
    .D(_0055_),
    .Q_N(_0707_),
    .Q(\ca.pulse_count[5] ));
 sg13g2_dfrbp_1 _1605_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net63),
    .D(_0056_),
    .Q_N(_0706_),
    .Q(\ca.pulse0 ));
 sg13g2_dfrbp_1 _1606_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net62),
    .D(_0057_),
    .Q_N(_0705_),
    .Q(\ca._13_ ));
 sg13g2_dfrbp_1 _1607_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net61),
    .D(_0058_),
    .Q_N(_0704_),
    .Q(\io_sd.input_index[3] ));
 sg13g2_dfrbp_1 _1608_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net59),
    .D(_0059_),
    .Q_N(_0014_),
    .Q(\io_sd.input_index[4] ));
 sg13g2_dfrbp_1 _1609_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net57),
    .D(net340),
    .Q_N(_0011_),
    .Q(\io_sd.input_index[5] ));
 sg13g2_dfrbp_1 _1610_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net55),
    .D(net154),
    .Q_N(_0703_),
    .Q(\io_sd.outputs[0] ));
 sg13g2_dfrbp_1 _1611_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net53),
    .D(net151),
    .Q_N(_0702_),
    .Q(\io_sd.outputs[1] ));
 sg13g2_dfrbp_1 _1612_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net51),
    .D(net149),
    .Q_N(_0701_),
    .Q(\io_sd.outputs[2] ));
 sg13g2_dfrbp_1 _1613_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net49),
    .D(net158),
    .Q_N(_0700_),
    .Q(\io_sd.outputs[3] ));
 sg13g2_dfrbp_1 _1614_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net47),
    .D(net147),
    .Q_N(_0699_),
    .Q(\io_sd.outputs[4] ));
 sg13g2_dfrbp_1 _1615_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net45),
    .D(net156),
    .Q_N(_0698_),
    .Q(\io_sd.outputs[5] ));
 sg13g2_dfrbp_1 _1616_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net43),
    .D(_0067_),
    .Q_N(_0697_),
    .Q(\io_sd.outputs[6] ));
 sg13g2_dfrbp_1 _1617_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net41),
    .D(net288),
    .Q_N(_0696_),
    .Q(\io_sd.outputs[7] ));
 sg13g2_dfrbp_1 _1618_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net39),
    .D(_0069_),
    .Q_N(_0695_),
    .Q(\io_sd._052_[0] ));
 sg13g2_dfrbp_1 _1619_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net33),
    .D(_0070_),
    .Q_N(_0694_),
    .Q(\io_sd._052_[1] ));
 sg13g2_dfrbp_1 _1620_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net31),
    .D(_0071_),
    .Q_N(_0693_),
    .Q(\io_sd._052_[2] ));
 sg13g2_dfrbp_1 _1621_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net29),
    .D(_0072_),
    .Q_N(_0692_),
    .Q(\io_sd._052_[3] ));
 sg13g2_dfrbp_1 _1622_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net25),
    .D(_0073_),
    .Q_N(_0691_),
    .Q(\io_sd._052_[4] ));
 sg13g2_dfrbp_1 _1623_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net120),
    .D(_0074_),
    .Q_N(_0690_),
    .Q(\io_sd._052_[5] ));
 sg13g2_dfrbp_1 _1624_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net116),
    .D(_0075_),
    .Q_N(_0689_),
    .Q(\io_sd._052_[6] ));
 sg13g2_dfrbp_1 _1625_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net112),
    .D(_0076_),
    .Q_N(_0688_),
    .Q(\io_sd._052_[7] ));
 sg13g2_dfrbp_1 _1626_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net108),
    .D(net301),
    .Q_N(_0687_),
    .Q(\io_sd._052_[8] ));
 sg13g2_dfrbp_1 _1627_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net104),
    .D(_0078_),
    .Q_N(_0686_),
    .Q(\io_sd._052_[9] ));
 sg13g2_dfrbp_1 _1628_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net100),
    .D(_0079_),
    .Q_N(_0685_),
    .Q(\io_sd._052_[10] ));
 sg13g2_dfrbp_1 _1629_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net96),
    .D(_0080_),
    .Q_N(_0684_),
    .Q(\io_sd._052_[11] ));
 sg13g2_dfrbp_1 _1630_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net92),
    .D(_0081_),
    .Q_N(_0683_),
    .Q(\io_sd._052_[12] ));
 sg13g2_dfrbp_1 _1631_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net88),
    .D(_0082_),
    .Q_N(_0682_),
    .Q(\io_sd._052_[13] ));
 sg13g2_dfrbp_1 _1632_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net84),
    .D(_0083_),
    .Q_N(_0681_),
    .Q(\io_sd._052_[14] ));
 sg13g2_dfrbp_1 _1633_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net80),
    .D(_0084_),
    .Q_N(_0680_),
    .Q(\io_sd._052_[15] ));
 sg13g2_dfrbp_1 _1634_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net76),
    .D(_0085_),
    .Q_N(_0679_),
    .Q(\io_sd._052_[16] ));
 sg13g2_dfrbp_1 _1635_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net72),
    .D(_0086_),
    .Q_N(_0678_),
    .Q(\io_sd._052_[17] ));
 sg13g2_dfrbp_1 _1636_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net68),
    .D(_0087_),
    .Q_N(_0677_),
    .Q(\io_sd._052_[18] ));
 sg13g2_dfrbp_1 _1637_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net64),
    .D(_0088_),
    .Q_N(_0676_),
    .Q(\io_sd._052_[19] ));
 sg13g2_dfrbp_1 _1638_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net58),
    .D(_0089_),
    .Q_N(_0675_),
    .Q(\io_sd._052_[20] ));
 sg13g2_dfrbp_1 _1639_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net54),
    .D(_0090_),
    .Q_N(_0674_),
    .Q(\io_sd._052_[21] ));
 sg13g2_dfrbp_1 _1640_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net50),
    .D(_0091_),
    .Q_N(_0673_),
    .Q(\io_sd._052_[22] ));
 sg13g2_dfrbp_1 _1641_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net46),
    .D(_0092_),
    .Q_N(_0672_),
    .Q(\io_sd._052_[23] ));
 sg13g2_dfrbp_1 _1642_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net42),
    .D(_0093_),
    .Q_N(_0671_),
    .Q(\io_sd._053_[0] ));
 sg13g2_dfrbp_1 _1643_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net38),
    .D(_0094_),
    .Q_N(_0670_),
    .Q(\io_sd._053_[1] ));
 sg13g2_dfrbp_1 _1644_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net30),
    .D(_0095_),
    .Q_N(_0669_),
    .Q(\io_sd._053_[2] ));
 sg13g2_dfrbp_1 _1645_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net123),
    .D(_0096_),
    .Q_N(_0668_),
    .Q(\io_sd._053_[3] ));
 sg13g2_dfrbp_1 _1646_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net114),
    .D(_0097_),
    .Q_N(_0667_),
    .Q(\io_sd._053_[4] ));
 sg13g2_dfrbp_1 _1647_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net106),
    .D(_0098_),
    .Q_N(_0666_),
    .Q(\io_sd._053_[5] ));
 sg13g2_dfrbp_1 _1648_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net98),
    .D(_0099_),
    .Q_N(_0665_),
    .Q(\io_sd._053_[6] ));
 sg13g2_dfrbp_1 _1649_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net90),
    .D(_0100_),
    .Q_N(_0664_),
    .Q(\io_sd._053_[7] ));
 sg13g2_dfrbp_1 _1650_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net82),
    .D(_0101_),
    .Q_N(_0663_),
    .Q(\io_sd._053_[8] ));
 sg13g2_dfrbp_1 _1651_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net74),
    .D(_0102_),
    .Q_N(_0662_),
    .Q(\io_sd._053_[9] ));
 sg13g2_dfrbp_1 _1652_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net66),
    .D(_0103_),
    .Q_N(_0661_),
    .Q(\io_sd._053_[10] ));
 sg13g2_dfrbp_1 _1653_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net56),
    .D(_0104_),
    .Q_N(_0660_),
    .Q(\io_sd._053_[11] ));
 sg13g2_dfrbp_1 _1654_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net48),
    .D(_0105_),
    .Q_N(_0659_),
    .Q(\io_sd._053_[12] ));
 sg13g2_dfrbp_1 _1655_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net40),
    .D(_0106_),
    .Q_N(_0658_),
    .Q(\io_sd._053_[13] ));
 sg13g2_dfrbp_1 _1656_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net27),
    .D(_0107_),
    .Q_N(_0657_),
    .Q(\io_sd._053_[14] ));
 sg13g2_dfrbp_1 _1657_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net110),
    .D(_0108_),
    .Q_N(_0656_),
    .Q(\io_sd._053_[15] ));
 sg13g2_dfrbp_1 _1658_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net94),
    .D(_0109_),
    .Q_N(_0655_),
    .Q(\io_sd._053_[16] ));
 sg13g2_dfrbp_1 _1659_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net78),
    .D(_0110_),
    .Q_N(_0654_),
    .Q(\io_sd._053_[17] ));
 sg13g2_dfrbp_1 _1660_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net60),
    .D(_0111_),
    .Q_N(_0653_),
    .Q(\io_sd._053_[18] ));
 sg13g2_dfrbp_1 _1661_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net44),
    .D(_0112_),
    .Q_N(_0652_),
    .Q(\io_sd._053_[19] ));
 sg13g2_dfrbp_1 _1662_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net118),
    .D(_0113_),
    .Q_N(_0651_),
    .Q(\io_sd._053_[20] ));
 sg13g2_dfrbp_1 _1663_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net86),
    .D(_0114_),
    .Q_N(_0650_),
    .Q(\io_sd._053_[21] ));
 sg13g2_dfrbp_1 _1664_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net52),
    .D(_0115_),
    .Q_N(_0649_),
    .Q(\io_sd._053_[22] ));
 sg13g2_dfrbp_1 _1665_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net102),
    .D(_0116_),
    .Q_N(_0648_),
    .Q(\io_sd._053_[23] ));
 sg13g2_dfrbp_1 _1666_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net132),
    .D(_0117_),
    .Q_N(_0015_),
    .Q(\io_sd._210_[0] ));
 sg13g2_dfrbp_1 _1667_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net133),
    .D(_0000_),
    .Q_N(_0746_),
    .Q(\bav1.state_q[0] ));
 sg13g2_dfrbp_1 _1668_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net134),
    .D(net326),
    .Q_N(_0747_),
    .Q(\bav1.state_q[1] ));
 sg13g2_dfrbp_1 _1669_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net135),
    .D(net185),
    .Q_N(_0748_),
    .Q(\bav1.state_q[2] ));
 sg13g2_dfrbp_1 _1670_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net136),
    .D(net253),
    .Q_N(_0749_),
    .Q(\bav1._02_ ));
 sg13g2_dfrbp_1 _1671_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net70),
    .D(_0004_),
    .Q_N(_0750_),
    .Q(\io_sd._083_ ));
 sg13g2_dfrbp_1 _1672_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net32),
    .D(net263),
    .Q_N(_0647_),
    .Q(\io_sd._080_ ));
 sg13g2_tiehi _1563__26 (.L_HI(net26));
 sg13g2_tiehi _1656__27 (.L_HI(net27));
 sg13g2_tiehi _1562__28 (.L_HI(net28));
 sg13g2_tiehi _1621__29 (.L_HI(net29));
 sg13g2_tiehi _1644__30 (.L_HI(net30));
 sg13g2_tiehi _1620__31 (.L_HI(net31));
 sg13g2_tiehi _1672__32 (.L_HI(net32));
 sg13g2_tiehi _1619__33 (.L_HI(net33));
 sg13g2_tiehi _1561__34 (.L_HI(net34));
 sg13g2_tiehi _1569__35 (.L_HI(net35));
 sg13g2_tiehi _1570__36 (.L_HI(net36));
 sg13g2_tiehi _1571__37 (.L_HI(net37));
 sg13g2_tiehi _1643__38 (.L_HI(net38));
 sg13g2_tiehi _1618__39 (.L_HI(net39));
 sg13g2_tiehi _1655__40 (.L_HI(net40));
 sg13g2_tiehi _1617__41 (.L_HI(net41));
 sg13g2_tiehi _1642__42 (.L_HI(net42));
 sg13g2_tiehi _1616__43 (.L_HI(net43));
 sg13g2_tiehi _1661__44 (.L_HI(net44));
 sg13g2_tiehi _1615__45 (.L_HI(net45));
 sg13g2_tiehi _1641__46 (.L_HI(net46));
 sg13g2_tiehi _1614__47 (.L_HI(net47));
 sg13g2_tiehi _1654__48 (.L_HI(net48));
 sg13g2_tiehi _1613__49 (.L_HI(net49));
 sg13g2_tiehi _1640__50 (.L_HI(net50));
 sg13g2_tiehi _1612__51 (.L_HI(net51));
 sg13g2_tiehi _1664__52 (.L_HI(net52));
 sg13g2_tiehi _1611__53 (.L_HI(net53));
 sg13g2_tiehi _1639__54 (.L_HI(net54));
 sg13g2_tiehi _1610__55 (.L_HI(net55));
 sg13g2_tiehi _1653__56 (.L_HI(net56));
 sg13g2_tiehi _1609__57 (.L_HI(net57));
 sg13g2_tiehi _1638__58 (.L_HI(net58));
 sg13g2_tiehi _1608__59 (.L_HI(net59));
 sg13g2_tiehi _1660__60 (.L_HI(net60));
 sg13g2_tiehi _1607__61 (.L_HI(net61));
 sg13g2_tiehi _1606__62 (.L_HI(net62));
 sg13g2_tiehi _1605__63 (.L_HI(net63));
 sg13g2_tiehi _1637__64 (.L_HI(net64));
 sg13g2_tiehi _1604__65 (.L_HI(net65));
 sg13g2_tiehi _1652__66 (.L_HI(net66));
 sg13g2_tiehi _1603__67 (.L_HI(net67));
 sg13g2_tiehi _1636__68 (.L_HI(net68));
 sg13g2_tiehi _1602__69 (.L_HI(net69));
 sg13g2_tiehi _1671__70 (.L_HI(net70));
 sg13g2_tiehi _1601__71 (.L_HI(net71));
 sg13g2_tiehi _1635__72 (.L_HI(net72));
 sg13g2_tiehi _1600__73 (.L_HI(net73));
 sg13g2_tiehi _1651__74 (.L_HI(net74));
 sg13g2_tiehi _1599__75 (.L_HI(net75));
 sg13g2_tiehi _1634__76 (.L_HI(net76));
 sg13g2_tiehi _1598__77 (.L_HI(net77));
 sg13g2_tiehi _1659__78 (.L_HI(net78));
 sg13g2_tiehi _1597__79 (.L_HI(net79));
 sg13g2_tiehi _1633__80 (.L_HI(net80));
 sg13g2_tiehi _1596__81 (.L_HI(net81));
 sg13g2_tiehi _1650__82 (.L_HI(net82));
 sg13g2_tiehi _1595__83 (.L_HI(net83));
 sg13g2_tiehi _1632__84 (.L_HI(net84));
 sg13g2_tiehi _1594__85 (.L_HI(net85));
 sg13g2_tiehi _1663__86 (.L_HI(net86));
 sg13g2_tiehi _1593__87 (.L_HI(net87));
 sg13g2_tiehi _1631__88 (.L_HI(net88));
 sg13g2_tiehi _1592__89 (.L_HI(net89));
 sg13g2_tiehi _1649__90 (.L_HI(net90));
 sg13g2_tiehi _1591__91 (.L_HI(net91));
 sg13g2_tiehi _1630__92 (.L_HI(net92));
 sg13g2_tiehi _1590__93 (.L_HI(net93));
 sg13g2_tiehi _1658__94 (.L_HI(net94));
 sg13g2_tiehi _1589__95 (.L_HI(net95));
 sg13g2_tiehi _1629__96 (.L_HI(net96));
 sg13g2_tiehi _1588__97 (.L_HI(net97));
 sg13g2_tiehi _1648__98 (.L_HI(net98));
 sg13g2_tiehi _1587__99 (.L_HI(net99));
 sg13g2_tiehi _1628__100 (.L_HI(net100));
 sg13g2_tiehi _1586__101 (.L_HI(net101));
 sg13g2_tiehi _1665__102 (.L_HI(net102));
 sg13g2_tiehi _1585__103 (.L_HI(net103));
 sg13g2_tiehi _1627__104 (.L_HI(net104));
 sg13g2_tiehi _1584__105 (.L_HI(net105));
 sg13g2_tiehi _1647__106 (.L_HI(net106));
 sg13g2_tiehi _1583__107 (.L_HI(net107));
 sg13g2_tiehi _1626__108 (.L_HI(net108));
 sg13g2_tiehi _1582__109 (.L_HI(net109));
 sg13g2_tiehi _1657__110 (.L_HI(net110));
 sg13g2_tiehi _1581__111 (.L_HI(net111));
 sg13g2_tiehi _1625__112 (.L_HI(net112));
 sg13g2_tiehi _1580__113 (.L_HI(net113));
 sg13g2_tiehi _1646__114 (.L_HI(net114));
 sg13g2_tiehi _1579__115 (.L_HI(net115));
 sg13g2_tiehi _1624__116 (.L_HI(net116));
 sg13g2_tiehi _1578__117 (.L_HI(net117));
 sg13g2_tiehi _1662__118 (.L_HI(net118));
 sg13g2_tiehi _1577__119 (.L_HI(net119));
 sg13g2_tiehi _1623__120 (.L_HI(net120));
 sg13g2_tiehi _1576__121 (.L_HI(net121));
 sg13g2_tiehi _1575__122 (.L_HI(net122));
 sg13g2_tiehi _1645__123 (.L_HI(net123));
 sg13g2_tiehi _1574__124 (.L_HI(net124));
 sg13g2_tiehi _1573__125 (.L_HI(net125));
 sg13g2_tiehi _1568__126 (.L_HI(net126));
 sg13g2_tiehi _1567__127 (.L_HI(net127));
 sg13g2_tiehi _1566__128 (.L_HI(net128));
 sg13g2_tiehi _1565__129 (.L_HI(net129));
 sg13g2_tiehi _1564__130 (.L_HI(net130));
 sg13g2_tiehi _1572__131 (.L_HI(net131));
 sg13g2_tiehi _1666__132 (.L_HI(net132));
 sg13g2_tiehi _1667__133 (.L_HI(net133));
 sg13g2_tiehi _1668__134 (.L_HI(net134));
 sg13g2_tiehi _1669__135 (.L_HI(net135));
 sg13g2_tiehi _1670__136 (.L_HI(net136));
 sg13g2_tiehi tt_um_cejmu_137 (.L_HI(net137));
 sg13g2_tiehi tt_um_cejmu_138 (.L_HI(net138));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_cejmu_14 (.L_LO(net14));
 sg13g2_tielo tt_um_cejmu_15 (.L_LO(net15));
 sg13g2_tielo tt_um_cejmu_16 (.L_LO(net16));
 sg13g2_tielo tt_um_cejmu_17 (.L_LO(net17));
 sg13g2_tielo tt_um_cejmu_18 (.L_LO(net18));
 sg13g2_tielo tt_um_cejmu_19 (.L_LO(net19));
 sg13g2_tielo tt_um_cejmu_20 (.L_LO(net20));
 sg13g2_tielo tt_um_cejmu_21 (.L_LO(net21));
 sg13g2_tielo tt_um_cejmu_22 (.L_LO(net22));
 sg13g2_tielo tt_um_cejmu_23 (.L_LO(net23));
 sg13g2_tielo tt_um_cejmu_24 (.L_LO(net24));
 sg13g2_tiehi _1622__25 (.L_HI(net25));
 sg13g2_buf_1 _1799_ (.A(\rca.generate_adder_modules[23].fa._02_ ),
    .X(uio_out[6]));
 sg13g2_and2_1 \cla/_591_  (.A(\rca.generate_adder_modules[21].fa.b ),
    .B(\rca.generate_adder_modules[21].fa.a ),
    .X(\cla/_565_ ));
 sg13g2_nor2_1 \cla/_592_  (.A(\rca.generate_adder_modules[21].fa.b ),
    .B(\rca.generate_adder_modules[21].fa.a ),
    .Y(\cla/_566_ ));
 sg13g2_nor2_2 \cla/_593_  (.A(\cla/_565_ ),
    .B(\cla/_566_ ),
    .Y(\cla/_567_ ));
 sg13g2_or2_2 \cla/_594_  (.X(\cla/_568_ ),
    .B(\cla/_566_ ),
    .A(\cla/_565_ ));
 sg13g2_nand2_1 \cla/_595_  (.Y(\cla/_569_ ),
    .A(\rca.generate_adder_modules[19].fa.b ),
    .B(\rca.generate_adder_modules[19].fa.a ));
 sg13g2_nor2_1 \cla/_596_  (.A(\rca.generate_adder_modules[19].fa.b ),
    .B(\rca.generate_adder_modules[19].fa.a ),
    .Y(\cla/_570_ ));
 sg13g2_xor2_1 \cla/_597_  (.B(\rca.generate_adder_modules[19].fa.a ),
    .A(\rca.generate_adder_modules[19].fa.b ),
    .X(\cla/_571_ ));
 sg13g2_xnor2_1 \cla/_598_  (.Y(\cla/_572_ ),
    .A(\rca.generate_adder_modules[19].fa.b ),
    .B(\rca.generate_adder_modules[19].fa.a ));
 sg13g2_nor2_1 \cla/_599_  (.A(\rca.generate_adder_modules[20].fa.b ),
    .B(\rca.generate_adder_modules[20].fa.a ),
    .Y(\cla/_573_ ));
 sg13g2_xor2_1 \cla/_600_  (.B(\rca.generate_adder_modules[20].fa.a ),
    .A(\rca.generate_adder_modules[20].fa.b ),
    .X(\cla/_574_ ));
 sg13g2_xnor2_1 \cla/_601_  (.Y(\cla/_575_ ),
    .A(\rca.generate_adder_modules[20].fa.b ),
    .B(\rca.generate_adder_modules[20].fa.a ));
 sg13g2_nor2_1 \cla/_602_  (.A(\cla/_572_ ),
    .B(\cla/_575_ ),
    .Y(\cla/_576_ ));
 sg13g2_nand2_1 \cla/_603_  (.Y(\cla/_577_ ),
    .A(\rca.generate_adder_modules[18].fa.b ),
    .B(\rca.generate_adder_modules[18].fa.a ));
 sg13g2_and2_1 \cla/_604_  (.A(\rca.generate_adder_modules[15].fa.b ),
    .B(\rca.generate_adder_modules[15].fa.a ),
    .X(\cla/_578_ ));
 sg13g2_or2_1 \cla/_605_  (.X(\cla/_579_ ),
    .B(\rca.generate_adder_modules[15].fa.a ),
    .A(\rca.generate_adder_modules[15].fa.b ));
 sg13g2_xor2_1 \cla/_606_  (.B(\rca.generate_adder_modules[15].fa.a ),
    .A(\rca.generate_adder_modules[15].fa.b ),
    .X(\cla/_580_ ));
 sg13g2_xnor2_1 \cla/_607_  (.Y(\cla/_581_ ),
    .A(\rca.generate_adder_modules[15].fa.b ),
    .B(\rca.generate_adder_modules[15].fa.a ));
 sg13g2_xor2_1 \cla/_608_  (.B(\rca.generate_adder_modules[18].fa.a ),
    .A(\rca.generate_adder_modules[18].fa.b ),
    .X(\cla/_582_ ));
 sg13g2_xnor2_1 \cla/_609_  (.Y(\cla/_583_ ),
    .A(\rca.generate_adder_modules[18].fa.b ),
    .B(\rca.generate_adder_modules[18].fa.a ));
 sg13g2_nand2_1 \cla/_610_  (.Y(\cla/_584_ ),
    .A(\rca.generate_adder_modules[16].fa.b ),
    .B(\rca.generate_adder_modules[16].fa.a ));
 sg13g2_xor2_1 \cla/_611_  (.B(\rca.generate_adder_modules[16].fa.a ),
    .A(\rca.generate_adder_modules[16].fa.b ),
    .X(\cla/_585_ ));
 sg13g2_nand2_2 \cla/_612_  (.Y(\cla/_586_ ),
    .A(\rca.generate_adder_modules[17].fa.b ),
    .B(\rca.generate_adder_modules[17].fa.a ));
 sg13g2_xor2_1 \cla/_613_  (.B(\rca.generate_adder_modules[17].fa.a ),
    .A(\rca.generate_adder_modules[17].fa.b ),
    .X(\cla/_587_ ));
 sg13g2_and2_1 \cla/_614_  (.A(\cla/_585_ ),
    .B(net197),
    .X(\cla/_588_ ));
 sg13g2_nand2_1 \cla/_615_  (.Y(\cla/_589_ ),
    .A(net198),
    .B(net197));
 sg13g2_nand2_1 \cla/_616_  (.Y(\cla/_590_ ),
    .A(\cla/_582_ ),
    .B(net197));
 sg13g2_nand3_1 \cla/_617_  (.B(net198),
    .C(net197),
    .A(\cla/_582_ ),
    .Y(\cla/_342_ ));
 sg13g2_nor2_1 \cla/_618_  (.A(\cla/_581_ ),
    .B(\cla/_342_ ),
    .Y(\cla/_343_ ));
 sg13g2_nand2_1 \cla/_619_  (.Y(\cla/_344_ ),
    .A(\rca.generate_adder_modules[14].fa.b ),
    .B(\rca.generate_adder_modules[14].fa.a ));
 sg13g2_xor2_1 \cla/_620_  (.B(\rca.generate_adder_modules[14].fa.a ),
    .A(\rca.generate_adder_modules[14].fa.b ),
    .X(\cla/_345_ ));
 sg13g2_xnor2_1 \cla/_621_  (.Y(\cla/_346_ ),
    .A(\rca.generate_adder_modules[14].fa.b ),
    .B(\rca.generate_adder_modules[14].fa.a ));
 sg13g2_nand2_2 \cla/_622_  (.Y(\cla/_347_ ),
    .A(\rca.generate_adder_modules[13].fa.b ),
    .B(\rca.generate_adder_modules[13].fa.a ));
 sg13g2_xor2_1 \cla/_623_  (.B(\rca.generate_adder_modules[13].fa.a ),
    .A(\rca.generate_adder_modules[13].fa.b ),
    .X(\cla/_348_ ));
 sg13g2_nand2_2 \cla/_624_  (.Y(\cla/_349_ ),
    .A(\cla/_345_ ),
    .B(\cla/_348_ ));
 sg13g2_inv_1 \cla/_625_  (.Y(\cla/_350_ ),
    .A(\cla/_349_ ));
 sg13g2_nand2_1 \cla/_626_  (.Y(\cla/_351_ ),
    .A(\rca.generate_adder_modules[10].fa.b ),
    .B(\rca.generate_adder_modules[10].fa.a ));
 sg13g2_nor2_1 \cla/_627_  (.A(\rca.generate_adder_modules[11].fa.b ),
    .B(\rca.generate_adder_modules[11].fa.a ),
    .Y(\cla/_352_ ));
 sg13g2_xor2_1 \cla/_628_  (.B(\rca.generate_adder_modules[11].fa.a ),
    .A(\rca.generate_adder_modules[11].fa.b ),
    .X(\cla/_353_ ));
 sg13g2_xnor2_1 \cla/_629_  (.Y(\cla/_354_ ),
    .A(\rca.generate_adder_modules[11].fa.b ),
    .B(\rca.generate_adder_modules[11].fa.a ));
 sg13g2_nand2_1 \cla/_630_  (.Y(\cla/_355_ ),
    .A(\rca.generate_adder_modules[12].fa.b ),
    .B(\rca.generate_adder_modules[12].fa.a ));
 sg13g2_xor2_1 \cla/_631_  (.B(\rca.generate_adder_modules[12].fa.a ),
    .A(\rca.generate_adder_modules[12].fa.b ),
    .X(\cla/_356_ ));
 sg13g2_nand2_1 \cla/_632_  (.Y(\cla/_357_ ),
    .A(\cla/_353_ ),
    .B(\cla/_356_ ));
 sg13g2_nand4_1 \cla/_633_  (.B(\rca.generate_adder_modules[10].fa.a ),
    .C(\cla/_353_ ),
    .A(\rca.generate_adder_modules[10].fa.b ),
    .Y(\cla/_358_ ),
    .D(\cla/_356_ ));
 sg13g2_o21ai_1 \cla/_634_  (.B1(\cla/_344_ ),
    .Y(\cla/_359_ ),
    .A1(\cla/_349_ ),
    .A2(\cla/_358_ ));
 sg13g2_nor4_2 \cla/_635_  (.A(\cla/_581_ ),
    .B(\cla/_342_ ),
    .C(\cla/_349_ ),
    .Y(\cla/_360_ ),
    .D(\cla/_358_ ));
 sg13g2_nand4_1 \cla/_636_  (.B(\rca.generate_adder_modules[14].fa.a ),
    .C(\cla/_580_ ),
    .A(\rca.generate_adder_modules[14].fa.b ),
    .Y(\cla/_361_ ),
    .D(net198));
 sg13g2_o21ai_1 \cla/_637_  (.B1(\cla/_577_ ),
    .Y(\cla/_362_ ),
    .A1(\cla/_590_ ),
    .A2(\cla/_361_ ));
 sg13g2_o21ai_1 \cla/_638_  (.B1(\cla/_576_ ),
    .Y(\cla/_363_ ),
    .A1(\cla/_360_ ),
    .A2(\cla/_362_ ));
 sg13g2_nor2_1 \cla/_639_  (.A(\cla/_568_ ),
    .B(\cla/_363_ ),
    .Y(\cla/_364_ ));
 sg13g2_nand2_1 \cla/_640_  (.Y(\cla/_365_ ),
    .A(\cla/_571_ ),
    .B(\cla/_582_ ));
 sg13g2_nor3_2 \cla/_641_  (.A(\cla/_572_ ),
    .B(\cla/_575_ ),
    .C(\cla/_583_ ),
    .Y(\cla/_366_ ));
 sg13g2_nand3_1 \cla/_642_  (.B(\cla/_574_ ),
    .C(\cla/_582_ ),
    .A(\cla/_571_ ),
    .Y(\cla/_367_ ));
 sg13g2_nand2_2 \cla/_643_  (.Y(\cla/_368_ ),
    .A(\cla/_567_ ),
    .B(\cla/_366_ ));
 sg13g2_nor2_2 \cla/_644_  (.A(\cla/_581_ ),
    .B(\cla/_346_ ),
    .Y(\cla/_369_ ));
 sg13g2_nand2_1 \cla/_645_  (.Y(\cla/_370_ ),
    .A(\cla/_580_ ),
    .B(\cla/_345_ ));
 sg13g2_nor2_1 \cla/_646_  (.A(\cla/_581_ ),
    .B(\cla/_589_ ),
    .Y(\cla/_371_ ));
 sg13g2_nand4_1 \cla/_647_  (.B(net198),
    .C(net197),
    .A(\cla/_580_ ),
    .Y(\cla/_372_ ),
    .D(\cla/_345_ ));
 sg13g2_o21ai_1 \cla/_648_  (.B1(\cla/_586_ ),
    .Y(\cla/_373_ ),
    .A1(\cla/_347_ ),
    .A2(\cla/_372_ ));
 sg13g2_and2_1 \cla/_649_  (.A(\cla/_348_ ),
    .B(\cla/_356_ ),
    .X(\cla/_374_ ));
 sg13g2_nand2_1 \cla/_650_  (.Y(\cla/_375_ ),
    .A(\cla/_348_ ),
    .B(\cla/_356_ ));
 sg13g2_xor2_1 \cla/_651_  (.B(\rca.generate_adder_modules[10].fa.a ),
    .A(\rca.generate_adder_modules[10].fa.b ),
    .X(\cla/_376_ ));
 sg13g2_xnor2_1 \cla/_652_  (.Y(\cla/_377_ ),
    .A(\rca.generate_adder_modules[10].fa.b ),
    .B(\rca.generate_adder_modules[10].fa.a ));
 sg13g2_and4_1 \cla/_653_  (.A(\rca.generate_adder_modules[9].fa.b ),
    .B(\rca.generate_adder_modules[9].fa.a ),
    .C(\cla/_353_ ),
    .D(\cla/_376_ ),
    .X(\cla/_378_ ));
 sg13g2_nand4_1 \cla/_654_  (.B(\rca.generate_adder_modules[9].fa.a ),
    .C(\cla/_353_ ),
    .A(\rca.generate_adder_modules[9].fa.b ),
    .Y(\cla/_379_ ),
    .D(\cla/_376_ ));
 sg13g2_nand4_1 \cla/_655_  (.B(\cla/_369_ ),
    .C(\cla/_374_ ),
    .A(\cla/_588_ ),
    .Y(\cla/_380_ ),
    .D(\cla/_378_ ));
 sg13g2_nor2b_1 \cla/_656_  (.A(\cla/_373_ ),
    .B_N(\cla/_380_ ),
    .Y(\cla/_381_ ));
 sg13g2_nor2_1 \cla/_657_  (.A(\cla/_368_ ),
    .B(\cla/_381_ ),
    .Y(\cla/_382_ ));
 sg13g2_and2_1 \cla/_658_  (.A(net197),
    .B(\cla/_366_ ),
    .X(\cla/_383_ ));
 sg13g2_nand2_1 \cla/_659_  (.Y(\cla/_384_ ),
    .A(\cla/_588_ ),
    .B(\cla/_366_ ));
 sg13g2_nor2_1 \cla/_660_  (.A(\cla/_568_ ),
    .B(\cla/_384_ ),
    .Y(\cla/_385_ ));
 sg13g2_nand2_1 \cla/_661_  (.Y(\cla/_386_ ),
    .A(\rca.generate_adder_modules[8].fa.b ),
    .B(\rca.generate_adder_modules[8].fa.a ));
 sg13g2_xnor2_1 \cla/_662_  (.Y(\cla/_387_ ),
    .A(\rca.generate_adder_modules[8].fa.b ),
    .B(\rca.generate_adder_modules[8].fa.a ));
 sg13g2_xnor2_1 \cla/_663_  (.Y(\cla/_388_ ),
    .A(\rca.generate_adder_modules[9].fa.b ),
    .B(\rca.generate_adder_modules[9].fa.a ));
 sg13g2_nor2_1 \cla/_664_  (.A(\cla/_387_ ),
    .B(\cla/_388_ ),
    .Y(\cla/_389_ ));
 sg13g2_nor4_2 \cla/_665_  (.A(\cla/_354_ ),
    .B(\cla/_377_ ),
    .C(\cla/_387_ ),
    .Y(\cla/_390_ ),
    .D(\cla/_388_ ));
 sg13g2_or4_2 \cla/_666_  (.A(\cla/_354_ ),
    .B(\cla/_377_ ),
    .C(\cla/_387_ ),
    .D(\cla/_388_ ),
    .X(\cla/_391_ ));
 sg13g2_nand2_1 \cla/_667_  (.Y(\cla/_392_ ),
    .A(\cla/_374_ ),
    .B(\cla/_390_ ));
 sg13g2_nor3_1 \cla/_668_  (.A(\cla/_370_ ),
    .B(\cla/_375_ ),
    .C(\cla/_391_ ),
    .Y(\cla/_393_ ));
 sg13g2_nand3_1 \cla/_669_  (.B(\cla/_374_ ),
    .C(\cla/_390_ ),
    .A(\cla/_369_ ),
    .Y(\cla/_394_ ));
 sg13g2_nand2_2 \cla/_670_  (.Y(\cla/_395_ ),
    .A(\rca.generate_adder_modules[4].fa.b ),
    .B(\rca.generate_adder_modules[4].fa.a ));
 sg13g2_nand2_1 \cla/_671_  (.Y(\cla/_396_ ),
    .A(\rca.generate_adder_modules[5].fa.b ),
    .B(\rca.generate_adder_modules[5].fa.a ));
 sg13g2_xnor2_1 \cla/_672_  (.Y(\cla/_397_ ),
    .A(\rca.generate_adder_modules[5].fa.b ),
    .B(\rca.generate_adder_modules[5].fa.a ));
 sg13g2_nor2_1 \cla/_673_  (.A(\rca.generate_adder_modules[7].fa.b ),
    .B(\rca.generate_adder_modules[7].fa.a ),
    .Y(\cla/_398_ ));
 sg13g2_nand2_1 \cla/_674_  (.Y(\cla/_399_ ),
    .A(\rca.generate_adder_modules[7].fa.b ),
    .B(\rca.generate_adder_modules[7].fa.a ));
 sg13g2_xnor2_1 \cla/_675_  (.Y(\cla/_400_ ),
    .A(\rca.generate_adder_modules[7].fa.b ),
    .B(\rca.generate_adder_modules[7].fa.a ));
 sg13g2_nand2_1 \cla/_676_  (.Y(\cla/_401_ ),
    .A(\rca.generate_adder_modules[6].fa.b ),
    .B(\rca.generate_adder_modules[6].fa.a ));
 sg13g2_nor2_1 \cla/_677_  (.A(\rca.generate_adder_modules[6].fa.b ),
    .B(\rca.generate_adder_modules[6].fa.a ),
    .Y(\cla/_402_ ));
 sg13g2_xnor2_1 \cla/_678_  (.Y(\cla/_403_ ),
    .A(\rca.generate_adder_modules[6].fa.b ),
    .B(\rca.generate_adder_modules[6].fa.a ));
 sg13g2_nor2_2 \cla/_679_  (.A(\cla/_400_ ),
    .B(\cla/_403_ ),
    .Y(\cla/_404_ ));
 sg13g2_nor3_2 \cla/_680_  (.A(\cla/_397_ ),
    .B(\cla/_400_ ),
    .C(\cla/_403_ ),
    .Y(\cla/_405_ ));
 sg13g2_nand2b_1 \cla/_681_  (.Y(\cla/_406_ ),
    .B(\cla/_404_ ),
    .A_N(\cla/_397_ ));
 sg13g2_nor2_1 \cla/_682_  (.A(\rca.generate_adder_modules[22].fa.b ),
    .B(\rca.generate_adder_modules[22].fa.a ),
    .Y(\cla/_407_ ));
 sg13g2_xnor2_1 \cla/_683_  (.Y(\cla/_408_ ),
    .A(\rca.generate_adder_modules[22].fa.b ),
    .B(\rca.generate_adder_modules[22].fa.a ));
 sg13g2_nor2_1 \cla/_684_  (.A(\cla/_406_ ),
    .B(\cla/_408_ ),
    .Y(\cla/_409_ ));
 sg13g2_nor4_1 \cla/_685_  (.A(\cla/_394_ ),
    .B(\cla/_395_ ),
    .C(\cla/_406_ ),
    .D(\cla/_408_ ),
    .Y(\cla/_410_ ));
 sg13g2_and2_1 \cla/_686_  (.A(\cla/_385_ ),
    .B(\cla/_410_ ),
    .X(\cla/_411_ ));
 sg13g2_xnor2_1 \cla/_687_  (.Y(\cla/_412_ ),
    .A(\rca.generate_adder_modules[4].fa.b ),
    .B(\rca.generate_adder_modules[4].fa.a ));
 sg13g2_and2_1 \cla/_688_  (.A(\rca.generate_adder_modules[2].fa.b ),
    .B(\rca.generate_adder_modules[2].fa.a ),
    .X(\cla/_413_ ));
 sg13g2_nand2_1 \cla/_689_  (.Y(\cla/_414_ ),
    .A(\rca.generate_adder_modules[2].fa.b ),
    .B(\rca.generate_adder_modules[2].fa.a ));
 sg13g2_nand2_1 \cla/_690_  (.Y(\cla/_415_ ),
    .A(\rca.generate_adder_modules[3].fa.b ),
    .B(\rca.generate_adder_modules[3].fa.a ));
 sg13g2_xnor2_1 \cla/_691_  (.Y(\cla/_416_ ),
    .A(\rca.generate_adder_modules[3].fa.b ),
    .B(\rca.generate_adder_modules[3].fa.a ));
 sg13g2_or2_1 \cla/_692_  (.X(\cla/_417_ ),
    .B(\cla/_416_ ),
    .A(\cla/_414_ ));
 sg13g2_nor2_2 \cla/_693_  (.A(\cla/_412_ ),
    .B(\cla/_416_ ),
    .Y(\cla/_418_ ));
 sg13g2_nand2_2 \cla/_694_  (.Y(\cla/_419_ ),
    .A(\cla/_413_ ),
    .B(\cla/_418_ ));
 sg13g2_nor4_1 \cla/_695_  (.A(\cla/_368_ ),
    .B(\cla/_372_ ),
    .C(\cla/_392_ ),
    .D(\cla/_419_ ),
    .Y(\cla/_420_ ));
 sg13g2_and2_1 \cla/_696_  (.A(\cla/_405_ ),
    .B(\cla/_420_ ),
    .X(\cla/_421_ ));
 sg13g2_nor2_1 \cla/_697_  (.A(\cla/_412_ ),
    .B(\cla/_415_ ),
    .Y(\cla/_422_ ));
 sg13g2_or4_1 \cla/_698_  (.A(\cla/_565_ ),
    .B(\cla/_382_ ),
    .C(\cla/_411_ ),
    .D(\cla/_421_ ),
    .X(\cla/_423_ ));
 sg13g2_nand4_1 \cla/_699_  (.B(\cla/_366_ ),
    .C(\cla/_393_ ),
    .A(\cla/_588_ ),
    .Y(\cla/_424_ ),
    .D(\cla/_422_ ));
 sg13g2_nor3_1 \cla/_700_  (.A(\cla/_568_ ),
    .B(\cla/_397_ ),
    .C(\cla/_424_ ),
    .Y(\cla/_425_ ));
 sg13g2_a21o_1 \cla/_701_  (.A2(\cla/_425_ ),
    .A1(\cla/_404_ ),
    .B1(\cla/_364_ ),
    .X(\cla/_426_ ));
 sg13g2_nor3_1 \cla/_702_  (.A(\cla/_372_ ),
    .B(\cla/_392_ ),
    .C(\cla/_419_ ),
    .Y(\cla/_427_ ));
 sg13g2_nand2_1 \cla/_703_  (.Y(\cla/_428_ ),
    .A(\cla/_405_ ),
    .B(\cla/_427_ ));
 sg13g2_xnor2_1 \cla/_704_  (.Y(\cla/_429_ ),
    .A(\rca.generate_adder_modules[23].fa.b ),
    .B(\rca.generate_adder_modules[23].fa.a ));
 sg13g2_nor2_1 \cla/_705_  (.A(\cla/_408_ ),
    .B(\cla/_429_ ),
    .Y(\cla/_430_ ));
 sg13g2_o21ai_1 \cla/_706_  (.B1(\cla/_430_ ),
    .Y(\cla/_431_ ),
    .A1(\cla/_423_ ),
    .A2(\cla/_426_ ));
 sg13g2_a22oi_1 \cla/_707_  (.Y(\cla/_432_ ),
    .B1(\rca.generate_adder_modules[22].fa.b ),
    .B2(\rca.generate_adder_modules[22].fa.a ),
    .A2(\rca.generate_adder_modules[23].fa.a ),
    .A1(\rca.generate_adder_modules[23].fa.b ));
 sg13g2_inv_1 \cla/_708_  (.Y(\cla/_433_ ),
    .A(\cla/_432_ ));
 sg13g2_o21ai_1 \cla/_709_  (.B1(\cla/_433_ ),
    .Y(\cla/_434_ ),
    .A1(\rca.generate_adder_modules[23].fa.b ),
    .A2(\rca.generate_adder_modules[23].fa.a ));
 sg13g2_and4_1 \cla/_710_  (.A(\cla/_580_ ),
    .B(net198),
    .C(\cla/_345_ ),
    .D(\cla/_348_ ),
    .X(\cla/_435_ ));
 sg13g2_nand4_1 \cla/_711_  (.B(net198),
    .C(\cla/_345_ ),
    .A(\cla/_580_ ),
    .Y(\cla/_436_ ),
    .D(\cla/_348_ ));
 sg13g2_nor2_1 \cla/_712_  (.A(\cla/_386_ ),
    .B(\cla/_388_ ),
    .Y(\cla/_437_ ));
 sg13g2_or3_1 \cla/_713_  (.A(\cla/_377_ ),
    .B(\cla/_386_ ),
    .C(\cla/_388_ ),
    .X(\cla/_438_ ));
 sg13g2_nor2_1 \cla/_714_  (.A(\cla/_357_ ),
    .B(\cla/_438_ ),
    .Y(\cla/_439_ ));
 sg13g2_nand3_1 \cla/_715_  (.B(\cla/_435_ ),
    .C(\cla/_439_ ),
    .A(\cla/_383_ ),
    .Y(\cla/_440_ ));
 sg13g2_nor2_1 \cla/_716_  (.A(\cla/_569_ ),
    .B(\cla/_573_ ),
    .Y(\cla/_441_ ));
 sg13g2_o21ai_1 \cla/_717_  (.B1(\cla/_584_ ),
    .Y(\cla/_442_ ),
    .A1(\cla/_355_ ),
    .A2(\cla/_436_ ));
 sg13g2_a221oi_1 \cla/_718_  (.B2(\cla/_442_ ),
    .C1(\cla/_441_ ),
    .B1(\cla/_383_ ),
    .A1(\rca.generate_adder_modules[20].fa.b ),
    .Y(\cla/_443_ ),
    .A2(\rca.generate_adder_modules[20].fa.a ));
 sg13g2_nand2_1 \cla/_719_  (.Y(\cla/_444_ ),
    .A(\cla/_440_ ),
    .B(\cla/_443_ ));
 sg13g2_and4_1 \cla/_720_  (.A(\rca.generate_adder_modules[11].fa.b ),
    .B(\rca.generate_adder_modules[11].fa.a ),
    .C(\cla/_348_ ),
    .D(\cla/_356_ ),
    .X(\cla/_445_ ));
 sg13g2_a21oi_1 \cla/_721_  (.A1(\cla/_369_ ),
    .A2(\cla/_445_ ),
    .Y(\cla/_446_ ),
    .B1(\cla/_578_ ));
 sg13g2_a21o_1 \cla/_722_  (.A2(\cla/_445_ ),
    .A1(\cla/_369_ ),
    .B1(\cla/_578_ ),
    .X(\cla/_447_ ));
 sg13g2_nor3_1 \cla/_723_  (.A(\cla/_396_ ),
    .B(\cla/_400_ ),
    .C(\cla/_403_ ),
    .Y(\cla/_448_ ));
 sg13g2_a21oi_2 \cla/_724_  (.B1(\cla/_398_ ),
    .Y(\cla/_449_ ),
    .A2(\cla/_401_ ),
    .A1(\cla/_399_ ));
 sg13g2_or2_1 \cla/_725_  (.X(\cla/_450_ ),
    .B(\cla/_449_ ),
    .A(\cla/_448_ ));
 sg13g2_a21oi_1 \cla/_726_  (.A1(\cla/_393_ ),
    .A2(\cla/_450_ ),
    .Y(\cla/_451_ ),
    .B1(\cla/_447_ ));
 sg13g2_nor3_1 \cla/_727_  (.A(\cla/_581_ ),
    .B(\cla/_589_ ),
    .C(\cla/_367_ ),
    .Y(\cla/_452_ ));
 sg13g2_nor2_1 \cla/_728_  (.A(\cla/_397_ ),
    .B(\cla/_412_ ),
    .Y(\cla/_453_ ));
 sg13g2_and2_1 \cla/_729_  (.A(\cla/_405_ ),
    .B(\cla/_418_ ),
    .X(\cla/_454_ ));
 sg13g2_nand2_2 \cla/_730_  (.Y(\cla/_455_ ),
    .A(\cla/_405_ ),
    .B(\cla/_418_ ));
 sg13g2_and2_1 \cla/_731_  (.A(\rca.generate_adder_modules[1].fa.b ),
    .B(\rca.generate_adder_modules[1].fa.a ),
    .X(\cla/_456_ ));
 sg13g2_and2_1 \cla/_732_  (.A(\rca.generate_adder_modules[0].fa.b ),
    .B(\rca.generate_adder_modules[0].fa.a ),
    .X(\cla/_457_ ));
 sg13g2_xor2_1 \cla/_733_  (.B(\rca.generate_adder_modules[1].fa.a ),
    .A(\rca.generate_adder_modules[1].fa.b ),
    .X(\cla/_458_ ));
 sg13g2_a21oi_2 \cla/_734_  (.B1(\cla/_456_ ),
    .Y(\cla/_459_ ),
    .A2(\cla/_458_ ),
    .A1(\cla/_457_ ));
 sg13g2_a21o_1 \cla/_735_  (.A2(\cla/_458_ ),
    .A1(\cla/_457_ ),
    .B1(\cla/_456_ ),
    .X(\cla/_460_ ));
 sg13g2_xor2_1 \cla/_736_  (.B(\rca.generate_adder_modules[2].fa.a ),
    .A(\rca.generate_adder_modules[2].fa.b ),
    .X(\cla/_461_ ));
 sg13g2_nand2_1 \cla/_737_  (.Y(\cla/_462_ ),
    .A(\cla/_460_ ),
    .B(\cla/_461_ ));
 sg13g2_nand2_1 \cla/_738_  (.Y(\cla/_463_ ),
    .A(\cla/_356_ ),
    .B(\cla/_461_ ));
 sg13g2_nor4_1 \cla/_739_  (.A(\cla/_391_ ),
    .B(\cla/_455_ ),
    .C(\cla/_459_ ),
    .D(\cla/_463_ ),
    .Y(\cla/_464_ ));
 sg13g2_nor4_2 \cla/_740_  (.A(\cla/_349_ ),
    .B(\cla/_391_ ),
    .C(\cla/_459_ ),
    .Y(\cla/_465_ ),
    .D(\cla/_463_ ));
 sg13g2_nand3_1 \cla/_741_  (.B(\cla/_454_ ),
    .C(\cla/_465_ ),
    .A(\cla/_452_ ),
    .Y(\cla/_466_ ));
 sg13g2_o21ai_1 \cla/_742_  (.B1(\cla/_466_ ),
    .Y(\cla/_467_ ),
    .A1(\cla/_384_ ),
    .A2(\cla/_451_ ));
 sg13g2_nor2_1 \cla/_743_  (.A(\cla/_568_ ),
    .B(\cla/_408_ ),
    .Y(\cla/_468_ ));
 sg13g2_nor3_1 \cla/_744_  (.A(\cla/_568_ ),
    .B(\cla/_408_ ),
    .C(\cla/_429_ ),
    .Y(\cla/_469_ ));
 sg13g2_o21ai_1 \cla/_745_  (.B1(\cla/_469_ ),
    .Y(\cla/_470_ ),
    .A1(\cla/_444_ ),
    .A2(\cla/_467_ ));
 sg13g2_nand3_1 \cla/_746_  (.B(\cla/_434_ ),
    .C(\cla/_470_ ),
    .A(\cla/_431_ ),
    .Y(\cla/_0341_ ));
 sg13g2_xor2_1 \cla/_747_  (.B(\rca.generate_adder_modules[0].fa.a ),
    .A(\rca.generate_adder_modules[0].fa.b ),
    .X(\cla/generate_adder_modules[0].fa_i._2_ ));
 sg13g2_o21ai_1 \cla/_748_  (.B1(\cla/_396_ ),
    .Y(\cla/_471_ ),
    .A1(\cla/_395_ ),
    .A2(\cla/_397_ ));
 sg13g2_a21oi_1 \cla/_749_  (.A1(\cla/_404_ ),
    .A2(\cla/_471_ ),
    .Y(\cla/_472_ ),
    .B1(\cla/_449_ ));
 sg13g2_a221oi_1 \cla/_750_  (.B2(\cla/_404_ ),
    .C1(\cla/_449_ ),
    .B1(\cla/_471_ ),
    .A1(\cla/_405_ ),
    .Y(\cla/_473_ ),
    .A2(\cla/_422_ ));
 sg13g2_a21oi_1 \cla/_751_  (.A1(\cla/_460_ ),
    .A2(\cla/_461_ ),
    .Y(\cla/_474_ ),
    .B1(\cla/_413_ ));
 sg13g2_nand2_1 \cla/_752_  (.Y(\cla/_475_ ),
    .A(\cla/_413_ ),
    .B(\cla/_454_ ));
 sg13g2_o21ai_1 \cla/_753_  (.B1(\cla/_473_ ),
    .Y(\cla/_476_ ),
    .A1(\cla/_455_ ),
    .A2(\cla/_474_ ));
 sg13g2_a221oi_1 \cla/_754_  (.B2(\cla/_476_ ),
    .C1(\cla/_437_ ),
    .B1(\cla/_389_ ),
    .A1(\rca.generate_adder_modules[9].fa.b ),
    .Y(\cla/_477_ ),
    .A2(\rca.generate_adder_modules[9].fa.a ));
 sg13g2_xnor2_1 \cla/_755_  (.Y(\cla/generate_adder_modules[10].fa_i._3_ ),
    .A(\cla/_376_ ),
    .B(\cla/_477_ ));
 sg13g2_o21ai_1 \cla/_756_  (.B1(\cla/_351_ ),
    .Y(\cla/_478_ ),
    .A1(\cla/_377_ ),
    .A2(\cla/_477_ ));
 sg13g2_xnor2_1 \cla/_757_  (.Y(\cla/generate_adder_modules[11].fa_i._3_ ),
    .A(\cla/_354_ ),
    .B(\cla/_478_ ));
 sg13g2_a21oi_1 \cla/_758_  (.A1(\cla/_351_ ),
    .A2(\cla/_438_ ),
    .Y(\cla/_479_ ),
    .B1(\cla/_352_ ));
 sg13g2_nand2_1 \cla/_759_  (.Y(\cla/_480_ ),
    .A(\cla/_390_ ),
    .B(\cla/_476_ ));
 sg13g2_a21oi_1 \cla/_760_  (.A1(\rca.generate_adder_modules[11].fa.b ),
    .A2(\rca.generate_adder_modules[11].fa.a ),
    .Y(\cla/_481_ ),
    .B1(\cla/_378_ ));
 sg13g2_nand2_1 \cla/_761_  (.Y(\cla/_482_ ),
    .A(\cla/_480_ ),
    .B(\cla/_481_ ));
 sg13g2_nor2_1 \cla/_762_  (.A(\cla/_479_ ),
    .B(\cla/_482_ ),
    .Y(\cla/_483_ ));
 sg13g2_xnor2_1 \cla/_763_  (.Y(\cla/generate_adder_modules[12].fa_i._3_ ),
    .A(\cla/_356_ ),
    .B(\cla/_483_ ));
 sg13g2_a21oi_2 \cla/_764_  (.B1(\cla/_439_ ),
    .Y(\cla/_484_ ),
    .A2(\rca.generate_adder_modules[12].fa.a ),
    .A1(\rca.generate_adder_modules[12].fa.b ));
 sg13g2_o21ai_1 \cla/_765_  (.B1(\cla/_355_ ),
    .Y(\cla/_485_ ),
    .A1(\cla/_357_ ),
    .A2(\cla/_438_ ));
 sg13g2_nand2_1 \cla/_766_  (.Y(\cla/_486_ ),
    .A(\cla/_358_ ),
    .B(\cla/_484_ ));
 sg13g2_a21oi_1 \cla/_767_  (.A1(\cla/_356_ ),
    .A2(\cla/_482_ ),
    .Y(\cla/_487_ ),
    .B1(\cla/_486_ ));
 sg13g2_xnor2_1 \cla/_768_  (.Y(\cla/generate_adder_modules[13].fa_i._3_ ),
    .A(\cla/_348_ ),
    .B(\cla/_487_ ));
 sg13g2_a21oi_1 \cla/_769_  (.A1(\cla/_473_ ),
    .A2(\cla/_475_ ),
    .Y(\cla/_488_ ),
    .B1(\cla/_392_ ));
 sg13g2_o21ai_1 \cla/_770_  (.B1(\cla/_347_ ),
    .Y(\cla/_489_ ),
    .A1(\cla/_375_ ),
    .A2(\cla/_379_ ));
 sg13g2_nor3_1 \cla/_771_  (.A(\cla/_445_ ),
    .B(\cla/_488_ ),
    .C(\cla/_489_ ),
    .Y(\cla/_490_ ));
 sg13g2_o21ai_1 \cla/_772_  (.B1(\cla/_348_ ),
    .Y(\cla/_491_ ),
    .A1(\cla/_464_ ),
    .A2(\cla/_486_ ));
 sg13g2_nand2_1 \cla/_773_  (.Y(\cla/_492_ ),
    .A(\cla/_490_ ),
    .B(\cla/_491_ ));
 sg13g2_xnor2_1 \cla/_774_  (.Y(\cla/generate_adder_modules[14].fa_i._3_ ),
    .A(\cla/_346_ ),
    .B(\cla/_492_ ));
 sg13g2_a22oi_1 \cla/_775_  (.Y(\cla/_493_ ),
    .B1(\cla/_485_ ),
    .B2(\cla/_350_ ),
    .A2(\cla/_465_ ),
    .A1(\cla/_454_ ));
 sg13g2_a21o_1 \cla/_776_  (.A2(\cla/_485_ ),
    .A1(\cla/_350_ ),
    .B1(\cla/_359_ ),
    .X(\cla/_494_ ));
 sg13g2_nor2b_1 \cla/_777_  (.A(\cla/_359_ ),
    .B_N(\cla/_493_ ),
    .Y(\cla/_495_ ));
 sg13g2_nand2b_1 \cla/_778_  (.Y(\cla/_496_ ),
    .B(\cla/_493_ ),
    .A_N(\cla/_359_ ));
 sg13g2_o21ai_1 \cla/_779_  (.B1(\cla/_495_ ),
    .Y(\cla/_497_ ),
    .A1(\cla/_346_ ),
    .A2(\cla/_490_ ));
 sg13g2_xnor2_1 \cla/_780_  (.Y(\cla/generate_adder_modules[15].fa_i._3_ ),
    .A(\cla/_581_ ),
    .B(\cla/_497_ ));
 sg13g2_and2_1 \cla/_781_  (.A(\cla/_369_ ),
    .B(\cla/_489_ ),
    .X(\cla/_498_ ));
 sg13g2_nor2_1 \cla/_782_  (.A(\cla/_394_ ),
    .B(\cla/_473_ ),
    .Y(\cla/_499_ ));
 sg13g2_o21ai_1 \cla/_783_  (.B1(\cla/_446_ ),
    .Y(\cla/_500_ ),
    .A1(\cla/_394_ ),
    .A2(\cla/_473_ ));
 sg13g2_nor4_1 \cla/_784_  (.A(\cla/_346_ ),
    .B(\cla/_375_ ),
    .C(\cla/_391_ ),
    .D(\cla/_417_ ),
    .Y(\cla/_501_ ));
 sg13g2_o21ai_1 \cla/_785_  (.B1(\cla/_580_ ),
    .Y(\cla/_502_ ),
    .A1(\cla/_465_ ),
    .A2(\cla/_501_ ));
 sg13g2_nor2_1 \cla/_786_  (.A(\cla/_455_ ),
    .B(\cla/_502_ ),
    .Y(\cla/_503_ ));
 sg13g2_or3_1 \cla/_787_  (.A(\cla/_498_ ),
    .B(\cla/_500_ ),
    .C(\cla/_503_ ),
    .X(\cla/_504_ ));
 sg13g2_a21o_1 \cla/_788_  (.A2(\cla/_494_ ),
    .A1(\cla/_579_ ),
    .B1(\cla/_504_ ),
    .X(\cla/_505_ ));
 sg13g2_xor2_1 \cla/_789_  (.B(\cla/_505_ ),
    .A(net198),
    .X(\cla/generate_adder_modules[16].fa_i._3_ ));
 sg13g2_nand2_1 \cla/_790_  (.Y(\cla/_506_ ),
    .A(\cla/_584_ ),
    .B(\cla/_361_ ));
 sg13g2_a221oi_1 \cla/_791_  (.B2(net198),
    .C1(\cla/_506_ ),
    .B1(\cla/_504_ ),
    .A1(\cla/_435_ ),
    .Y(\cla/_507_ ),
    .A2(\cla/_486_ ));
 sg13g2_xnor2_1 \cla/_792_  (.Y(\cla/generate_adder_modules[17].fa_i._3_ ),
    .A(net197),
    .B(\cla/_507_ ));
 sg13g2_a21o_1 \cla/_793_  (.A2(\cla/_371_ ),
    .A1(\cla/_359_ ),
    .B1(\cla/_500_ ),
    .X(\cla/_508_ ));
 sg13g2_o21ai_1 \cla/_794_  (.B1(\cla/_588_ ),
    .Y(\cla/_509_ ),
    .A1(\cla/_503_ ),
    .A2(\cla/_508_ ));
 sg13g2_o21ai_1 \cla/_795_  (.B1(\cla/_584_ ),
    .Y(\cla/_510_ ),
    .A1(\cla/_436_ ),
    .A2(\cla/_484_ ));
 sg13g2_nand2_1 \cla/_796_  (.Y(\cla/_511_ ),
    .A(net197),
    .B(\cla/_510_ ));
 sg13g2_nand3_1 \cla/_797_  (.B(\cla/_509_ ),
    .C(\cla/_511_ ),
    .A(\cla/_381_ ),
    .Y(\cla/_512_ ));
 sg13g2_xnor2_1 \cla/_798_  (.Y(\cla/generate_adder_modules[18].fa_i._3_ ),
    .A(\cla/_583_ ),
    .B(\cla/_512_ ));
 sg13g2_o21ai_1 \cla/_799_  (.B1(\cla/_373_ ),
    .Y(\cla/_513_ ),
    .A1(\rca.generate_adder_modules[18].fa.b ),
    .A2(\rca.generate_adder_modules[18].fa.a ));
 sg13g2_or2_1 \cla/_800_  (.X(\cla/_514_ ),
    .B(\cla/_380_ ),
    .A(\cla/_583_ ));
 sg13g2_or2_1 \cla/_801_  (.X(\cla/_515_ ),
    .B(\cla/_590_ ),
    .A(\cla/_584_ ));
 sg13g2_nand4_1 \cla/_802_  (.B(\cla/_513_ ),
    .C(\cla/_514_ ),
    .A(\cla/_577_ ),
    .Y(\cla/_516_ ),
    .D(\cla/_515_ ));
 sg13g2_a21oi_1 \cla/_803_  (.A1(\cla/_405_ ),
    .A2(\cla/_427_ ),
    .Y(\cla/_517_ ),
    .B1(\cla/_500_ ));
 sg13g2_a21oi_1 \cla/_804_  (.A1(\cla/_343_ ),
    .A2(\cla/_496_ ),
    .Y(\cla/_518_ ),
    .B1(\cla/_516_ ));
 sg13g2_o21ai_1 \cla/_805_  (.B1(\cla/_518_ ),
    .Y(\cla/_519_ ),
    .A1(\cla/_342_ ),
    .A2(\cla/_517_ ));
 sg13g2_xnor2_1 \cla/_806_  (.Y(\cla/generate_adder_modules[19].fa_i._3_ ),
    .A(\cla/_572_ ),
    .B(\cla/_519_ ));
 sg13g2_xor2_1 \cla/_807_  (.B(\cla/_458_ ),
    .A(\cla/_457_ ),
    .X(\cla/generate_adder_modules[1].fa_i._3_ ));
 sg13g2_nand2b_1 \cla/_808_  (.Y(\cla/_520_ ),
    .B(\cla/_343_ ),
    .A_N(\cla/_493_ ));
 sg13g2_nor2b_1 \cla/_809_  (.A(\cla/_360_ ),
    .B_N(\cla/_514_ ),
    .Y(\cla/_521_ ));
 sg13g2_a21oi_1 \cla/_810_  (.A1(\cla/_520_ ),
    .A2(\cla/_521_ ),
    .Y(\cla/_522_ ),
    .B1(\cla/_572_ ));
 sg13g2_o21ai_1 \cla/_811_  (.B1(\cla/_446_ ),
    .Y(\cla/_523_ ),
    .A1(\cla/_347_ ),
    .A2(\cla/_370_ ));
 sg13g2_nor2_1 \cla/_812_  (.A(\cla/_589_ ),
    .B(\cla/_365_ ),
    .Y(\cla/_524_ ));
 sg13g2_o21ai_1 \cla/_813_  (.B1(\cla/_524_ ),
    .Y(\cla/_525_ ),
    .A1(\cla/_499_ ),
    .A2(\cla/_523_ ));
 sg13g2_o21ai_1 \cla/_814_  (.B1(\cla/_569_ ),
    .Y(\cla/_526_ ),
    .A1(\cla/_586_ ),
    .A2(\cla/_365_ ));
 sg13g2_or2_1 \cla/_815_  (.X(\cla/_527_ ),
    .B(\cla/_577_ ),
    .A(\cla/_570_ ));
 sg13g2_nand2_1 \cla/_816_  (.Y(\cla/_528_ ),
    .A(\cla/_587_ ),
    .B(\cla/_506_ ));
 sg13g2_a21oi_1 \cla/_817_  (.A1(\cla/_428_ ),
    .A2(\cla/_528_ ),
    .Y(\cla/_529_ ),
    .B1(\cla/_365_ ));
 sg13g2_nand3b_1 \cla/_818_  (.B(\cla/_527_ ),
    .C(\cla/_525_ ),
    .Y(\cla/_530_ ),
    .A_N(\cla/_526_ ));
 sg13g2_nor3_1 \cla/_819_  (.A(\cla/_522_ ),
    .B(\cla/_529_ ),
    .C(\cla/_530_ ),
    .Y(\cla/_531_ ));
 sg13g2_xnor2_1 \cla/_820_  (.Y(\cla/generate_adder_modules[20].fa_i._3_ ),
    .A(\cla/_574_ ),
    .B(\cla/_531_ ));
 sg13g2_a21oi_1 \cla/_821_  (.A1(\cla/_586_ ),
    .A2(\cla/_428_ ),
    .Y(\cla/_532_ ),
    .B1(\cla/_367_ ));
 sg13g2_nor2_1 \cla/_822_  (.A(\cla/_394_ ),
    .B(\cla/_472_ ),
    .Y(\cla/_533_ ));
 sg13g2_nor3_1 \cla/_823_  (.A(\cla/_447_ ),
    .B(\cla/_498_ ),
    .C(\cla/_533_ ),
    .Y(\cla/_534_ ));
 sg13g2_nor2_1 \cla/_824_  (.A(\cla/_384_ ),
    .B(\cla/_534_ ),
    .Y(\cla/_535_ ));
 sg13g2_nand3_1 \cla/_825_  (.B(\cla/_440_ ),
    .C(\cla/_443_ ),
    .A(\cla/_363_ ),
    .Y(\cla/_536_ ));
 sg13g2_nand3_1 \cla/_826_  (.B(\cla/_452_ ),
    .C(\cla/_465_ ),
    .A(\cla/_418_ ),
    .Y(\cla/_537_ ));
 sg13g2_a21oi_1 \cla/_827_  (.A1(\cla/_424_ ),
    .A2(\cla/_537_ ),
    .Y(\cla/_538_ ),
    .B1(\cla/_406_ ));
 sg13g2_nor4_1 \cla/_828_  (.A(\cla/_532_ ),
    .B(\cla/_535_ ),
    .C(\cla/_536_ ),
    .D(\cla/_538_ ),
    .Y(\cla/_539_ ));
 sg13g2_xnor2_1 \cla/_829_  (.Y(\cla/generate_adder_modules[21].fa_i._3_ ),
    .A(\cla/_567_ ),
    .B(\cla/_539_ ));
 sg13g2_o21ai_1 \cla/_830_  (.B1(\cla/_385_ ),
    .Y(\cla/_540_ ),
    .A1(\cla/_523_ ),
    .A2(\cla/_533_ ));
 sg13g2_nand3_1 \cla/_831_  (.B(\cla/_574_ ),
    .C(\cla/_526_ ),
    .A(\cla/_567_ ),
    .Y(\cla/_541_ ));
 sg13g2_a22oi_1 \cla/_832_  (.Y(\cla/_542_ ),
    .B1(\rca.generate_adder_modules[21].fa.b ),
    .B2(\rca.generate_adder_modules[21].fa.a ),
    .A2(\rca.generate_adder_modules[20].fa.a ),
    .A1(\rca.generate_adder_modules[20].fa.b ));
 sg13g2_nor2_1 \cla/_833_  (.A(\cla/_566_ ),
    .B(\cla/_542_ ),
    .Y(\cla/_543_ ));
 sg13g2_nand2_1 \cla/_834_  (.Y(\cla/_544_ ),
    .A(\cla/_567_ ),
    .B(\cla/_538_ ));
 sg13g2_o21ai_1 \cla/_835_  (.B1(\cla/_541_ ),
    .Y(\cla/_545_ ),
    .A1(\cla/_368_ ),
    .A2(\cla/_380_ ));
 sg13g2_nor4_1 \cla/_836_  (.A(\cla/_364_ ),
    .B(\cla/_421_ ),
    .C(\cla/_543_ ),
    .D(\cla/_545_ ),
    .Y(\cla/_546_ ));
 sg13g2_nand3_1 \cla/_837_  (.B(\cla/_383_ ),
    .C(\cla/_510_ ),
    .A(\cla/_567_ ),
    .Y(\cla/_547_ ));
 sg13g2_nand4_1 \cla/_838_  (.B(\cla/_544_ ),
    .C(\cla/_546_ ),
    .A(\cla/_540_ ),
    .Y(\cla/_548_ ),
    .D(\cla/_547_ ));
 sg13g2_xnor2_1 \cla/_839_  (.Y(\cla/generate_adder_modules[22].fa_i._3_ ),
    .A(\cla/_408_ ),
    .B(\cla/_548_ ));
 sg13g2_o21ai_1 \cla/_840_  (.B1(\cla/_468_ ),
    .Y(\cla/_549_ ),
    .A1(\cla/_467_ ),
    .A2(\cla/_536_ ));
 sg13g2_nor3_1 \cla/_841_  (.A(\cla/_368_ ),
    .B(\cla/_381_ ),
    .C(\cla/_408_ ),
    .Y(\cla/_550_ ));
 sg13g2_a22oi_1 \cla/_842_  (.Y(\cla/_551_ ),
    .B1(\rca.generate_adder_modules[22].fa.b ),
    .B2(\rca.generate_adder_modules[22].fa.a ),
    .A2(\rca.generate_adder_modules[21].fa.a ),
    .A1(\rca.generate_adder_modules[21].fa.b ));
 sg13g2_nor2_1 \cla/_843_  (.A(\cla/_407_ ),
    .B(\cla/_551_ ),
    .Y(\cla/_552_ ));
 sg13g2_nor3_1 \cla/_844_  (.A(\cla/_411_ ),
    .B(\cla/_550_ ),
    .C(\cla/_552_ ),
    .Y(\cla/_553_ ));
 sg13g2_o21ai_1 \cla/_845_  (.B1(\cla/_409_ ),
    .Y(\cla/_554_ ),
    .A1(\cla/_420_ ),
    .A2(\cla/_425_ ));
 sg13g2_nand3_1 \cla/_846_  (.B(\cla/_553_ ),
    .C(\cla/_554_ ),
    .A(\cla/_549_ ),
    .Y(\cla/_555_ ));
 sg13g2_xnor2_1 \cla/_847_  (.Y(\cla/generate_adder_modules[23].fa_i._3_ ),
    .A(\cla/_429_ ),
    .B(\cla/_555_ ));
 sg13g2_xnor2_1 \cla/_848_  (.Y(\cla/generate_adder_modules[2].fa_i._3_ ),
    .A(\cla/_459_ ),
    .B(\cla/_461_ ));
 sg13g2_xor2_1 \cla/_849_  (.B(\cla/_474_ ),
    .A(\cla/_416_ ),
    .X(\cla/generate_adder_modules[3].fa_i._3_ ));
 sg13g2_o21ai_1 \cla/_850_  (.B1(\cla/_415_ ),
    .Y(\cla/_556_ ),
    .A1(\cla/_416_ ),
    .A2(\cla/_462_ ));
 sg13g2_nand2b_1 \cla/_851_  (.Y(\cla/_557_ ),
    .B(\cla/_417_ ),
    .A_N(\cla/_556_ ));
 sg13g2_xnor2_1 \cla/_852_  (.Y(\cla/generate_adder_modules[4].fa_i._3_ ),
    .A(\cla/_412_ ),
    .B(\cla/_557_ ));
 sg13g2_o21ai_1 \cla/_853_  (.B1(\cla/_556_ ),
    .Y(\cla/_558_ ),
    .A1(\rca.generate_adder_modules[4].fa.b ),
    .A2(\rca.generate_adder_modules[4].fa.a ));
 sg13g2_nand3_1 \cla/_854_  (.B(\cla/_419_ ),
    .C(\cla/_558_ ),
    .A(\cla/_395_ ),
    .Y(\cla/_559_ ));
 sg13g2_xnor2_1 \cla/_855_  (.Y(\cla/generate_adder_modules[5].fa_i._3_ ),
    .A(\cla/_397_ ),
    .B(\cla/_559_ ));
 sg13g2_a21oi_1 \cla/_856_  (.A1(\cla/_395_ ),
    .A2(\cla/_419_ ),
    .Y(\cla/_560_ ),
    .B1(\cla/_397_ ));
 sg13g2_a221oi_1 \cla/_857_  (.B2(\cla/_556_ ),
    .C1(\cla/_560_ ),
    .B1(\cla/_453_ ),
    .A1(\rca.generate_adder_modules[5].fa.b ),
    .Y(\cla/_561_ ),
    .A2(\rca.generate_adder_modules[5].fa.a ));
 sg13g2_xor2_1 \cla/_858_  (.B(\cla/_561_ ),
    .A(\cla/_403_ ),
    .X(\cla/generate_adder_modules[6].fa_i._3_ ));
 sg13g2_o21ai_1 \cla/_859_  (.B1(\cla/_401_ ),
    .Y(\cla/_562_ ),
    .A1(\cla/_402_ ),
    .A2(\cla/_561_ ));
 sg13g2_xnor2_1 \cla/_860_  (.Y(\cla/generate_adder_modules[7].fa_i._3_ ),
    .A(\cla/_400_ ),
    .B(\cla/_562_ ));
 sg13g2_xnor2_1 \cla/_861_  (.Y(\cla/generate_adder_modules[8].fa_i._3_ ),
    .A(\cla/_387_ ),
    .B(\cla/_476_ ));
 sg13g2_o21ai_1 \cla/_862_  (.B1(\cla/_476_ ),
    .Y(\cla/_563_ ),
    .A1(\rca.generate_adder_modules[8].fa.b ),
    .A2(\rca.generate_adder_modules[8].fa.a ));
 sg13g2_nand2_1 \cla/_863_  (.Y(\cla/_564_ ),
    .A(\cla/_386_ ),
    .B(\cla/_563_ ));
 sg13g2_xnor2_1 \cla/_864_  (.Y(\cla/generate_adder_modules[9].fa_i._3_ ),
    .A(\cla/_388_ ),
    .B(\cla/_564_ ));
 sg13g2_buf_1 \cla/_865_  (.A(\cla/generate_adder_modules[0].fa_i._2_ ),
    .X(\cla_z[0] ));
 sg13g2_buf_1 \cla/_866_  (.A(\cla/generate_adder_modules[1].fa_i._3_ ),
    .X(\cla_z[1] ));
 sg13g2_buf_1 \cla/_867_  (.A(\cla/generate_adder_modules[2].fa_i._3_ ),
    .X(\cla_z[2] ));
 sg13g2_buf_1 \cla/_868_  (.A(\cla/generate_adder_modules[3].fa_i._3_ ),
    .X(\cla_z[3] ));
 sg13g2_buf_1 \cla/_869_  (.A(\cla/generate_adder_modules[4].fa_i._3_ ),
    .X(\cla_z[4] ));
 sg13g2_buf_1 \cla/_870_  (.A(\cla/generate_adder_modules[5].fa_i._3_ ),
    .X(\cla_z[5] ));
 sg13g2_buf_1 \cla/_871_  (.A(\cla/generate_adder_modules[6].fa_i._3_ ),
    .X(\cla_z[6] ));
 sg13g2_buf_1 \cla/_872_  (.A(\cla/generate_adder_modules[7].fa_i._3_ ),
    .X(\cla_z[7] ));
 sg13g2_buf_1 \cla/_873_  (.A(\cla/generate_adder_modules[8].fa_i._3_ ),
    .X(\cla_z[8] ));
 sg13g2_buf_1 \cla/_874_  (.A(\cla/generate_adder_modules[9].fa_i._3_ ),
    .X(\cla_z[9] ));
 sg13g2_buf_1 \cla/_875_  (.A(\cla/generate_adder_modules[10].fa_i._3_ ),
    .X(\cla_z[10] ));
 sg13g2_buf_1 \cla/_876_  (.A(\cla/generate_adder_modules[11].fa_i._3_ ),
    .X(\cla_z[11] ));
 sg13g2_buf_1 \cla/_877_  (.A(\cla/generate_adder_modules[12].fa_i._3_ ),
    .X(\cla_z[12] ));
 sg13g2_buf_1 \cla/_878_  (.A(\cla/generate_adder_modules[13].fa_i._3_ ),
    .X(\cla_z[13] ));
 sg13g2_buf_1 \cla/_879_  (.A(\cla/generate_adder_modules[14].fa_i._3_ ),
    .X(\cla_z[14] ));
 sg13g2_buf_1 \cla/_880_  (.A(\cla/generate_adder_modules[15].fa_i._3_ ),
    .X(\cla_z[15] ));
 sg13g2_buf_1 \cla/_881_  (.A(\cla/generate_adder_modules[16].fa_i._3_ ),
    .X(\cla_z[16] ));
 sg13g2_buf_1 \cla/_882_  (.A(\cla/generate_adder_modules[17].fa_i._3_ ),
    .X(\cla_z[17] ));
 sg13g2_buf_1 \cla/_883_  (.A(\cla/generate_adder_modules[18].fa_i._3_ ),
    .X(\cla_z[18] ));
 sg13g2_buf_1 \cla/_884_  (.A(\cla/generate_adder_modules[19].fa_i._3_ ),
    .X(\cla_z[19] ));
 sg13g2_buf_1 \cla/_885_  (.A(\cla/generate_adder_modules[20].fa_i._3_ ),
    .X(\cla_z[20] ));
 sg13g2_buf_1 \cla/_886_  (.A(\cla/generate_adder_modules[21].fa_i._3_ ),
    .X(\cla_z[21] ));
 sg13g2_buf_1 \cla/_887_  (.A(\cla/generate_adder_modules[22].fa_i._3_ ),
    .X(\cla_z[22] ));
 sg13g2_buf_1 \cla/_888_  (.A(\cla/generate_adder_modules[23].fa_i._3_ ),
    .X(\cla_z[23] ));
 sg13g2_buf_2 \cla/_889_  (.A(\cla/_0341_ ),
    .X(uio_out[7]));
 sg13g2_buf_4 fanout190 (.X(net190),
    .A(_0373_));
 sg13g2_buf_2 fanout191 (.A(_0373_),
    .X(net191));
 sg13g2_buf_4 fanout192 (.X(net192),
    .A(_0372_));
 sg13g2_buf_2 fanout193 (.A(net195),
    .X(net193));
 sg13g2_buf_2 fanout194 (.A(net195),
    .X(net194));
 sg13g2_buf_2 fanout195 (.A(_0282_),
    .X(net195));
 sg13g2_buf_2 fanout196 (.A(_0527_),
    .X(net196));
 sg13g2_buf_2 fanout197 (.A(\cla/_587_ ),
    .X(net197));
 sg13g2_buf_2 fanout198 (.A(\cla/_585_ ),
    .X(net198));
 sg13g2_buf_2 fanout199 (.A(_0530_),
    .X(net199));
 sg13g2_buf_4 fanout200 (.X(net200),
    .A(net201));
 sg13g2_buf_2 fanout201 (.A(_0342_),
    .X(net201));
 sg13g2_buf_4 fanout202 (.X(net202),
    .A(net203));
 sg13g2_buf_2 fanout203 (.A(_0342_),
    .X(net203));
 sg13g2_buf_4 fanout204 (.X(net204),
    .A(_0342_));
 sg13g2_buf_2 fanout205 (.A(net208),
    .X(net205));
 sg13g2_buf_4 fanout206 (.X(net206),
    .A(net207));
 sg13g2_buf_2 fanout207 (.A(net208),
    .X(net207));
 sg13g2_buf_2 fanout208 (.A(_0344_),
    .X(net208));
 sg13g2_buf_4 fanout209 (.X(net209),
    .A(_0344_));
 sg13g2_buf_2 fanout210 (.A(_0143_),
    .X(net210));
 sg13g2_buf_1 fanout211 (.A(_0143_),
    .X(net211));
 sg13g2_buf_2 fanout212 (.A(net214),
    .X(net212));
 sg13g2_buf_1 fanout213 (.A(net214),
    .X(net213));
 sg13g2_buf_1 fanout214 (.A(_0133_),
    .X(net214));
 sg13g2_buf_4 fanout215 (.X(net215),
    .A(net216));
 sg13g2_buf_4 fanout216 (.X(net216),
    .A(\io_sd._210_[0] ));
 sg13g2_buf_2 fanout217 (.A(\io_sd.input_index[3] ),
    .X(net217));
 sg13g2_buf_2 fanout218 (.A(\io_sd._209_[0] ),
    .X(net218));
 sg13g2_buf_2 fanout219 (.A(net220),
    .X(net219));
 sg13g2_buf_2 fanout220 (.A(net345),
    .X(net220));
 sg13g2_buf_2 fanout221 (.A(net223),
    .X(net221));
 sg13g2_buf_1 fanout222 (.A(net223),
    .X(net222));
 sg13g2_buf_2 fanout223 (.A(net228),
    .X(net223));
 sg13g2_buf_2 fanout224 (.A(net225),
    .X(net224));
 sg13g2_buf_2 fanout225 (.A(net228),
    .X(net225));
 sg13g2_buf_2 fanout226 (.A(net227),
    .X(net226));
 sg13g2_buf_2 fanout227 (.A(net228),
    .X(net227));
 sg13g2_buf_2 fanout228 (.A(_0369_),
    .X(net228));
 sg13g2_buf_2 fanout229 (.A(net230),
    .X(net229));
 sg13g2_buf_2 fanout230 (.A(net231),
    .X(net230));
 sg13g2_buf_4 fanout231 (.X(net231),
    .A(_0135_));
 sg13g2_buf_2 fanout232 (.A(net234),
    .X(net232));
 sg13g2_buf_2 fanout233 (.A(net234),
    .X(net233));
 sg13g2_buf_2 fanout234 (.A(_0135_),
    .X(net234));
 sg13g2_buf_2 fanout235 (.A(net237),
    .X(net235));
 sg13g2_buf_2 fanout236 (.A(net237),
    .X(net236));
 sg13g2_buf_2 fanout237 (.A(_0135_),
    .X(net237));
 sg13g2_buf_2 fanout238 (.A(net239),
    .X(net238));
 sg13g2_buf_2 fanout239 (.A(net245),
    .X(net239));
 sg13g2_buf_2 fanout240 (.A(net241),
    .X(net240));
 sg13g2_buf_2 fanout241 (.A(net245),
    .X(net241));
 sg13g2_buf_2 fanout242 (.A(net245),
    .X(net242));
 sg13g2_buf_1 fanout243 (.A(net244),
    .X(net243));
 sg13g2_buf_2 fanout244 (.A(net245),
    .X(net244));
 sg13g2_buf_2 fanout245 (.A(uio_in[2]),
    .X(net245));
 sg13g2_buf_2 fanout246 (.A(net11),
    .X(net246));
 sg13g2_buf_4 fanout247 (.X(net247),
    .A(net249));
 sg13g2_buf_1 fanout248 (.A(net249),
    .X(net248));
 sg13g2_buf_2 fanout249 (.A(net1),
    .X(net249));
 sg13g2_buf_1 input1 (.A(rst_n),
    .X(net1));
 sg13g2_buf_2 input2 (.A(ui_in[0]),
    .X(net2));
 sg13g2_buf_2 input3 (.A(ui_in[1]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[2]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[3]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[4]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[5]),
    .X(net7));
 sg13g2_buf_2 input8 (.A(ui_in[6]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(ui_in[7]),
    .X(net9));
 sg13g2_buf_1 input10 (.A(uio_in[0]),
    .X(net10));
 sg13g2_buf_1 input11 (.A(uio_in[1]),
    .X(net11));
 sg13g2_buf_2 input12 (.A(uio_in[3]),
    .X(net12));
 sg13g2_tielo tt_um_cejmu_13 (.L_LO(net13));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\ca._07_[0] ),
    .X(net139));
 sg13g2_dlygate4sd3_1 hold2 (.A(_0331_),
    .X(net140));
 sg13g2_dlygate4sd3_1 hold3 (.A(\ca._08_[0] ),
    .X(net141));
 sg13g2_dlygate4sd3_1 hold4 (.A(_0285_),
    .X(net142));
 sg13g2_dlygate4sd3_1 hold5 (.A(\ca.pulse_count[3] ),
    .X(net143));
 sg13g2_dlygate4sd3_1 hold6 (.A(\ca.pulse_count[2] ),
    .X(net144));
 sg13g2_dlygate4sd3_1 hold7 (.A(\io_sd.outputs[6] ),
    .X(net145));
 sg13g2_dlygate4sd3_1 hold8 (.A(\io_sd.outputs[4] ),
    .X(net146));
 sg13g2_dlygate4sd3_1 hold9 (.A(_0065_),
    .X(net147));
 sg13g2_dlygate4sd3_1 hold10 (.A(\io_sd.outputs[2] ),
    .X(net148));
 sg13g2_dlygate4sd3_1 hold11 (.A(_0063_),
    .X(net149));
 sg13g2_dlygate4sd3_1 hold12 (.A(\io_sd.outputs[1] ),
    .X(net150));
 sg13g2_dlygate4sd3_1 hold13 (.A(_0062_),
    .X(net151));
 sg13g2_dlygate4sd3_1 hold14 (.A(\ca.pulse_count[1] ),
    .X(net152));
 sg13g2_dlygate4sd3_1 hold15 (.A(\io_sd.outputs[0] ),
    .X(net153));
 sg13g2_dlygate4sd3_1 hold16 (.A(_0061_),
    .X(net154));
 sg13g2_dlygate4sd3_1 hold17 (.A(\io_sd.outputs[5] ),
    .X(net155));
 sg13g2_dlygate4sd3_1 hold18 (.A(_0066_),
    .X(net156));
 sg13g2_dlygate4sd3_1 hold19 (.A(\io_sd.outputs[3] ),
    .X(net157));
 sg13g2_dlygate4sd3_1 hold20 (.A(_0064_),
    .X(net158));
 sg13g2_dlygate4sd3_1 hold21 (.A(\ca.pulse_count[4] ),
    .X(net159));
 sg13g2_dlygate4sd3_1 hold22 (.A(\ca.pulse_count[0] ),
    .X(net160));
 sg13g2_dlygate4sd3_1 hold23 (.A(\ca.pulse_count[5] ),
    .X(net161));
 sg13g2_dlygate4sd3_1 hold24 (.A(\ca._11_ ),
    .X(net162));
 sg13g2_dlygate4sd3_1 hold25 (.A(\ca.pulse0 ),
    .X(net163));
 sg13g2_dlygate4sd3_1 hold26 (.A(\ca.commit_count[1] ),
    .X(net164));
 sg13g2_dlygate4sd3_1 hold27 (.A(_0287_),
    .X(net165));
 sg13g2_dlygate4sd3_1 hold28 (.A(_0028_),
    .X(net166));
 sg13g2_dlygate4sd3_1 hold29 (.A(\bav0.state_q[1] ),
    .X(net167));
 sg13g2_dlygate4sd3_1 hold30 (.A(_0009_),
    .X(net168));
 sg13g2_dlygate4sd3_1 hold31 (.A(\ca._13_ ),
    .X(net169));
 sg13g2_dlygate4sd3_1 hold32 (.A(\io_sd._052_[22] ),
    .X(net170));
 sg13g2_dlygate4sd3_1 hold33 (.A(\io_sd._053_[23] ),
    .X(net171));
 sg13g2_dlygate4sd3_1 hold34 (.A(\ca.commit_count[9] ),
    .X(net172));
 sg13g2_dlygate4sd3_1 hold35 (.A(_0301_),
    .X(net173));
 sg13g2_dlygate4sd3_1 hold36 (.A(_0036_),
    .X(net174));
 sg13g2_dlygate4sd3_1 hold37 (.A(\bav0.state_q[2] ),
    .X(net175));
 sg13g2_dlygate4sd3_1 hold38 (.A(_0007_),
    .X(net176));
 sg13g2_dlygate4sd3_1 hold39 (.A(\io_sd._052_[20] ),
    .X(net177));
 sg13g2_dlygate4sd3_1 hold40 (.A(\io_sd._052_[10] ),
    .X(net178));
 sg13g2_dlygate4sd3_1 hold41 (.A(\io_sd._052_[11] ),
    .X(net179));
 sg13g2_dlygate4sd3_1 hold42 (.A(\io_sd._052_[19] ),
    .X(net180));
 sg13g2_dlygate4sd3_1 hold43 (.A(\io_sd._052_[15] ),
    .X(net181));
 sg13g2_dlygate4sd3_1 hold44 (.A(\bav0.state_q[0] ),
    .X(net182));
 sg13g2_dlygate4sd3_1 hold45 (.A(\io_sd._052_[21] ),
    .X(net183));
 sg13g2_dlygate4sd3_1 hold46 (.A(\bav1.state_q[2] ),
    .X(net184));
 sg13g2_dlygate4sd3_1 hold47 (.A(_0002_),
    .X(net185));
 sg13g2_dlygate4sd3_1 hold48 (.A(\io_sd._052_[18] ),
    .X(net186));
 sg13g2_dlygate4sd3_1 hold49 (.A(\io_sd._053_[0] ),
    .X(net187));
 sg13g2_dlygate4sd3_1 hold50 (.A(\io_sd._053_[10] ),
    .X(net188));
 sg13g2_dlygate4sd3_1 hold51 (.A(\io_sd._052_[23] ),
    .X(net189));
 sg13g2_dlygate4sd3_1 hold52 (.A(\io_sd._052_[7] ),
    .X(net250));
 sg13g2_dlygate4sd3_1 hold53 (.A(\bav1.state_q[1] ),
    .X(net251));
 sg13g2_dlygate4sd3_1 hold54 (.A(_0169_),
    .X(net252));
 sg13g2_dlygate4sd3_1 hold55 (.A(_0003_),
    .X(net253));
 sg13g2_dlygate4sd3_1 hold56 (.A(\io_sd._052_[12] ),
    .X(net254));
 sg13g2_dlygate4sd3_1 hold57 (.A(\io_sd._053_[19] ),
    .X(net255));
 sg13g2_dlygate4sd3_1 hold58 (.A(\io_sd._053_[20] ),
    .X(net256));
 sg13g2_dlygate4sd3_1 hold59 (.A(\ca.commit_count[19] ),
    .X(net257));
 sg13g2_dlygate4sd3_1 hold60 (.A(_0322_),
    .X(net258));
 sg13g2_dlygate4sd3_1 hold61 (.A(_0046_),
    .X(net259));
 sg13g2_dlygate4sd3_1 hold62 (.A(\ca.commit_count[2] ),
    .X(net260));
 sg13g2_dlygate4sd3_1 hold63 (.A(_0289_),
    .X(net261));
 sg13g2_dlygate4sd3_1 hold64 (.A(\io_sd._080_ ),
    .X(net262));
 sg13g2_dlygate4sd3_1 hold65 (.A(_0005_),
    .X(net263));
 sg13g2_dlygate4sd3_1 hold66 (.A(\io_sd._052_[9] ),
    .X(net264));
 sg13g2_dlygate4sd3_1 hold67 (.A(\io_sd._053_[22] ),
    .X(net265));
 sg13g2_dlygate4sd3_1 hold68 (.A(\io_sd._052_[13] ),
    .X(net266));
 sg13g2_dlygate4sd3_1 hold69 (.A(\io_sd._052_[14] ),
    .X(net267));
 sg13g2_dlygate4sd3_1 hold70 (.A(\io_sd._052_[3] ),
    .X(net268));
 sg13g2_dlygate4sd3_1 hold71 (.A(\ca.commit_count[4] ),
    .X(net269));
 sg13g2_dlygate4sd3_1 hold72 (.A(_0293_),
    .X(net270));
 sg13g2_dlygate4sd3_1 hold73 (.A(\ca.commit_count[5] ),
    .X(net271));
 sg13g2_dlygate4sd3_1 hold74 (.A(\io_sd._052_[4] ),
    .X(net272));
 sg13g2_dlygate4sd3_1 hold75 (.A(_0565_),
    .X(net273));
 sg13g2_dlygate4sd3_1 hold76 (.A(\io_sd._053_[9] ),
    .X(net274));
 sg13g2_dlygate4sd3_1 hold77 (.A(\io_sd._053_[18] ),
    .X(net275));
 sg13g2_dlygate4sd3_1 hold78 (.A(\io_sd._053_[11] ),
    .X(net276));
 sg13g2_dlygate4sd3_1 hold79 (.A(\ca.commit_count[3] ),
    .X(net277));
 sg13g2_dlygate4sd3_1 hold80 (.A(\io_sd._052_[17] ),
    .X(net278));
 sg13g2_dlygate4sd3_1 hold81 (.A(\bav1.state_q[0] ),
    .X(net279));
 sg13g2_dlygate4sd3_1 hold82 (.A(\ca.commit_count[7] ),
    .X(net280));
 sg13g2_dlygate4sd3_1 hold83 (.A(_0298_),
    .X(net281));
 sg13g2_dlygate4sd3_1 hold84 (.A(\io_sd._053_[12] ),
    .X(net282));
 sg13g2_dlygate4sd3_1 hold85 (.A(\io_sd._053_[6] ),
    .X(net283));
 sg13g2_dlygate4sd3_1 hold86 (.A(\io_sd._053_[14] ),
    .X(net284));
 sg13g2_dlygate4sd3_1 hold87 (.A(\io_sd._053_[17] ),
    .X(net285));
 sg13g2_dlygate4sd3_1 hold88 (.A(\io_sd._053_[3] ),
    .X(net286));
 sg13g2_dlygate4sd3_1 hold89 (.A(_0012_),
    .X(net287));
 sg13g2_dlygate4sd3_1 hold90 (.A(_0068_),
    .X(net288));
 sg13g2_dlygate4sd3_1 hold91 (.A(\io_sd._053_[4] ),
    .X(net289));
 sg13g2_dlygate4sd3_1 hold92 (.A(\io_sd._053_[7] ),
    .X(net290));
 sg13g2_dlygate4sd3_1 hold93 (.A(\io_sd._052_[6] ),
    .X(net291));
 sg13g2_dlygate4sd3_1 hold94 (.A(\io_sd.output_index[5] ),
    .X(net292));
 sg13g2_dlygate4sd3_1 hold95 (.A(_0018_),
    .X(net293));
 sg13g2_dlygate4sd3_1 hold96 (.A(\io_sd._053_[21] ),
    .X(net294));
 sg13g2_dlygate4sd3_1 hold97 (.A(\ca.commit_count[20] ),
    .X(net295));
 sg13g2_dlygate4sd3_1 hold98 (.A(_0324_),
    .X(net296));
 sg13g2_dlygate4sd3_1 hold99 (.A(\ca.commit_count[18] ),
    .X(net297));
 sg13g2_dlygate4sd3_1 hold100 (.A(_0045_),
    .X(net298));
 sg13g2_dlygate4sd3_1 hold101 (.A(\io_sd._052_[8] ),
    .X(net299));
 sg13g2_dlygate4sd3_1 hold102 (.A(_0583_),
    .X(net300));
 sg13g2_dlygate4sd3_1 hold103 (.A(_0077_),
    .X(net301));
 sg13g2_dlygate4sd3_1 hold104 (.A(\io_sd._052_[0] ),
    .X(net302));
 sg13g2_dlygate4sd3_1 hold105 (.A(\ca.commit_count[6] ),
    .X(net303));
 sg13g2_dlygate4sd3_1 hold106 (.A(\io_sd._052_[2] ),
    .X(net304));
 sg13g2_dlygate4sd3_1 hold107 (.A(\io_sd._053_[13] ),
    .X(net305));
 sg13g2_dlygate4sd3_1 hold108 (.A(\ca.commit_count[15] ),
    .X(net306));
 sg13g2_dlygate4sd3_1 hold109 (.A(_0314_),
    .X(net307));
 sg13g2_dlygate4sd3_1 hold110 (.A(\io_sd._053_[1] ),
    .X(net308));
 sg13g2_dlygate4sd3_1 hold111 (.A(\ca.commit_count[17] ),
    .X(net309));
 sg13g2_dlygate4sd3_1 hold112 (.A(_0319_),
    .X(net310));
 sg13g2_dlygate4sd3_1 hold113 (.A(_0044_),
    .X(net311));
 sg13g2_dlygate4sd3_1 hold114 (.A(\ca.commit_count[13] ),
    .X(net312));
 sg13g2_dlygate4sd3_1 hold115 (.A(_0309_),
    .X(net313));
 sg13g2_dlygate4sd3_1 hold116 (.A(\io_sd._052_[5] ),
    .X(net314));
 sg13g2_dlygate4sd3_1 hold117 (.A(_0570_),
    .X(net315));
 sg13g2_dlygate4sd3_1 hold118 (.A(\ca.commit_count[12] ),
    .X(net316));
 sg13g2_dlygate4sd3_1 hold119 (.A(_0307_),
    .X(net317));
 sg13g2_dlygate4sd3_1 hold120 (.A(\ca.commit_count[8] ),
    .X(net318));
 sg13g2_dlygate4sd3_1 hold121 (.A(\io_sd._053_[2] ),
    .X(net319));
 sg13g2_dlygate4sd3_1 hold122 (.A(\io_sd._053_[5] ),
    .X(net320));
 sg13g2_dlygate4sd3_1 hold123 (.A(_0636_),
    .X(net321));
 sg13g2_dlygate4sd3_1 hold124 (.A(\io_sd._052_[1] ),
    .X(net322));
 sg13g2_dlygate4sd3_1 hold125 (.A(\ca._15_ ),
    .X(net323));
 sg13g2_dlygate4sd3_1 hold126 (.A(\io_sd._052_[16] ),
    .X(net324));
 sg13g2_dlygate4sd3_1 hold127 (.A(\bav1.x[1] ),
    .X(net325));
 sg13g2_dlygate4sd3_1 hold128 (.A(_0001_),
    .X(net326));
 sg13g2_dlygate4sd3_1 hold129 (.A(\ca.commit_count[21] ),
    .X(net327));
 sg13g2_dlygate4sd3_1 hold130 (.A(\io_sd.input_index[4] ),
    .X(net328));
 sg13g2_dlygate4sd3_1 hold131 (.A(_0348_),
    .X(net329));
 sg13g2_dlygate4sd3_1 hold132 (.A(\ca.commit_count[14] ),
    .X(net330));
 sg13g2_dlygate4sd3_1 hold133 (.A(\io_sd.output_index[4] ),
    .X(net331));
 sg13g2_dlygate4sd3_1 hold134 (.A(_0264_),
    .X(net332));
 sg13g2_dlygate4sd3_1 hold135 (.A(\io_sd._053_[8] ),
    .X(net333));
 sg13g2_dlygate4sd3_1 hold136 (.A(\io_sd._083_ ),
    .X(net334));
 sg13g2_dlygate4sd3_1 hold137 (.A(\ca.commit_count[11] ),
    .X(net335));
 sg13g2_dlygate4sd3_1 hold138 (.A(_0306_),
    .X(net336));
 sg13g2_dlygate4sd3_1 hold139 (.A(\ca.commit_count[10] ),
    .X(net337));
 sg13g2_dlygate4sd3_1 hold140 (.A(\ca.commit_count[16] ),
    .X(net338));
 sg13g2_dlygate4sd3_1 hold141 (.A(\io_sd.input_index[5] ),
    .X(net339));
 sg13g2_dlygate4sd3_1 hold142 (.A(_0060_),
    .X(net340));
 sg13g2_dlygate4sd3_1 hold143 (.A(\io_sd._053_[16] ),
    .X(net341));
 sg13g2_dlygate4sd3_1 hold144 (.A(\io_sd._053_[15] ),
    .X(net342));
 sg13g2_dlygate4sd3_1 hold145 (.A(\io_sd.input_index[3] ),
    .X(net343));
 sg13g2_dlygate4sd3_1 hold146 (.A(_0010_),
    .X(net344));
 sg13g2_dlygate4sd3_1 hold147 (.A(\io_sd.output_index[3] ),
    .X(net345));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_fill_1 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_348 ();
 sg13g2_decap_8 FILLER_5_355 ();
 sg13g2_decap_8 FILLER_5_362 ();
 sg13g2_decap_8 FILLER_5_369 ();
 sg13g2_decap_8 FILLER_5_376 ();
 sg13g2_decap_8 FILLER_5_383 ();
 sg13g2_decap_8 FILLER_5_390 ();
 sg13g2_decap_8 FILLER_5_397 ();
 sg13g2_decap_4 FILLER_5_404 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_4 FILLER_6_168 ();
 sg13g2_fill_1 FILLER_6_172 ();
 sg13g2_decap_8 FILLER_6_177 ();
 sg13g2_decap_8 FILLER_6_184 ();
 sg13g2_fill_1 FILLER_6_191 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_291 ();
 sg13g2_decap_8 FILLER_6_324 ();
 sg13g2_fill_2 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_363 ();
 sg13g2_decap_8 FILLER_6_370 ();
 sg13g2_decap_8 FILLER_6_377 ();
 sg13g2_decap_8 FILLER_6_384 ();
 sg13g2_decap_8 FILLER_6_391 ();
 sg13g2_decap_8 FILLER_6_398 ();
 sg13g2_decap_4 FILLER_6_405 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_4 FILLER_7_140 ();
 sg13g2_decap_4 FILLER_7_153 ();
 sg13g2_fill_1 FILLER_7_157 ();
 sg13g2_decap_8 FILLER_7_204 ();
 sg13g2_decap_8 FILLER_7_211 ();
 sg13g2_decap_8 FILLER_7_218 ();
 sg13g2_decap_8 FILLER_7_225 ();
 sg13g2_decap_4 FILLER_7_232 ();
 sg13g2_fill_1 FILLER_7_236 ();
 sg13g2_fill_1 FILLER_7_241 ();
 sg13g2_fill_1 FILLER_7_248 ();
 sg13g2_decap_4 FILLER_7_254 ();
 sg13g2_fill_2 FILLER_7_258 ();
 sg13g2_decap_4 FILLER_7_271 ();
 sg13g2_fill_2 FILLER_7_275 ();
 sg13g2_decap_4 FILLER_7_303 ();
 sg13g2_fill_1 FILLER_7_320 ();
 sg13g2_decap_8 FILLER_7_382 ();
 sg13g2_decap_8 FILLER_7_389 ();
 sg13g2_decap_8 FILLER_7_396 ();
 sg13g2_decap_4 FILLER_7_403 ();
 sg13g2_fill_2 FILLER_7_407 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_fill_2 FILLER_8_42 ();
 sg13g2_fill_1 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_75 ();
 sg13g2_decap_8 FILLER_8_82 ();
 sg13g2_decap_4 FILLER_8_89 ();
 sg13g2_fill_2 FILLER_8_97 ();
 sg13g2_fill_1 FILLER_8_99 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_4 FILLER_8_112 ();
 sg13g2_fill_1 FILLER_8_116 ();
 sg13g2_fill_1 FILLER_8_122 ();
 sg13g2_decap_8 FILLER_8_127 ();
 sg13g2_fill_1 FILLER_8_134 ();
 sg13g2_decap_4 FILLER_8_157 ();
 sg13g2_fill_1 FILLER_8_161 ();
 sg13g2_decap_4 FILLER_8_166 ();
 sg13g2_fill_2 FILLER_8_170 ();
 sg13g2_decap_8 FILLER_8_177 ();
 sg13g2_fill_2 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_223 ();
 sg13g2_fill_2 FILLER_8_230 ();
 sg13g2_fill_2 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_277 ();
 sg13g2_decap_4 FILLER_8_290 ();
 sg13g2_fill_2 FILLER_8_294 ();
 sg13g2_fill_2 FILLER_8_301 ();
 sg13g2_fill_2 FILLER_8_316 ();
 sg13g2_fill_1 FILLER_8_318 ();
 sg13g2_fill_2 FILLER_8_331 ();
 sg13g2_fill_1 FILLER_8_333 ();
 sg13g2_fill_1 FILLER_8_361 ();
 sg13g2_fill_2 FILLER_8_388 ();
 sg13g2_decap_8 FILLER_8_398 ();
 sg13g2_decap_4 FILLER_8_405 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_4 FILLER_9_56 ();
 sg13g2_fill_2 FILLER_9_86 ();
 sg13g2_fill_1 FILLER_9_114 ();
 sg13g2_decap_4 FILLER_9_133 ();
 sg13g2_fill_1 FILLER_9_137 ();
 sg13g2_fill_2 FILLER_9_147 ();
 sg13g2_decap_4 FILLER_9_185 ();
 sg13g2_fill_1 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_202 ();
 sg13g2_fill_2 FILLER_9_237 ();
 sg13g2_decap_8 FILLER_9_244 ();
 sg13g2_fill_2 FILLER_9_251 ();
 sg13g2_fill_1 FILLER_9_253 ();
 sg13g2_fill_2 FILLER_9_276 ();
 sg13g2_fill_2 FILLER_9_294 ();
 sg13g2_fill_1 FILLER_9_296 ();
 sg13g2_fill_2 FILLER_9_349 ();
 sg13g2_fill_2 FILLER_9_381 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_fill_2 FILLER_10_50 ();
 sg13g2_fill_1 FILLER_10_52 ();
 sg13g2_fill_2 FILLER_10_82 ();
 sg13g2_fill_1 FILLER_10_84 ();
 sg13g2_fill_2 FILLER_10_90 ();
 sg13g2_fill_2 FILLER_10_96 ();
 sg13g2_decap_8 FILLER_10_104 ();
 sg13g2_decap_8 FILLER_10_111 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_fill_1 FILLER_10_140 ();
 sg13g2_fill_2 FILLER_10_145 ();
 sg13g2_fill_1 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_162 ();
 sg13g2_decap_8 FILLER_10_169 ();
 sg13g2_decap_8 FILLER_10_176 ();
 sg13g2_fill_1 FILLER_10_183 ();
 sg13g2_decap_8 FILLER_10_200 ();
 sg13g2_fill_1 FILLER_10_207 ();
 sg13g2_decap_8 FILLER_10_225 ();
 sg13g2_decap_8 FILLER_10_232 ();
 sg13g2_decap_4 FILLER_10_259 ();
 sg13g2_fill_1 FILLER_10_263 ();
 sg13g2_fill_2 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_293 ();
 sg13g2_decap_4 FILLER_10_300 ();
 sg13g2_fill_1 FILLER_10_304 ();
 sg13g2_decap_4 FILLER_10_314 ();
 sg13g2_decap_4 FILLER_10_322 ();
 sg13g2_fill_1 FILLER_10_326 ();
 sg13g2_fill_1 FILLER_10_337 ();
 sg13g2_fill_2 FILLER_10_364 ();
 sg13g2_fill_1 FILLER_10_366 ();
 sg13g2_fill_1 FILLER_10_404 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_fill_2 FILLER_11_28 ();
 sg13g2_fill_1 FILLER_11_30 ();
 sg13g2_decap_4 FILLER_11_35 ();
 sg13g2_fill_2 FILLER_11_65 ();
 sg13g2_fill_1 FILLER_11_67 ();
 sg13g2_fill_1 FILLER_11_100 ();
 sg13g2_decap_4 FILLER_11_109 ();
 sg13g2_fill_1 FILLER_11_113 ();
 sg13g2_fill_1 FILLER_11_153 ();
 sg13g2_fill_2 FILLER_11_159 ();
 sg13g2_fill_1 FILLER_11_161 ();
 sg13g2_fill_2 FILLER_11_167 ();
 sg13g2_fill_1 FILLER_11_178 ();
 sg13g2_fill_1 FILLER_11_185 ();
 sg13g2_decap_4 FILLER_11_192 ();
 sg13g2_fill_2 FILLER_11_196 ();
 sg13g2_decap_4 FILLER_11_231 ();
 sg13g2_fill_1 FILLER_11_235 ();
 sg13g2_fill_2 FILLER_11_253 ();
 sg13g2_fill_1 FILLER_11_255 ();
 sg13g2_decap_8 FILLER_11_282 ();
 sg13g2_fill_1 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_327 ();
 sg13g2_decap_8 FILLER_11_334 ();
 sg13g2_fill_2 FILLER_11_364 ();
 sg13g2_fill_2 FILLER_11_377 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_4 FILLER_12_14 ();
 sg13g2_fill_2 FILLER_12_18 ();
 sg13g2_fill_1 FILLER_12_46 ();
 sg13g2_fill_2 FILLER_12_81 ();
 sg13g2_fill_1 FILLER_12_83 ();
 sg13g2_fill_2 FILLER_12_101 ();
 sg13g2_decap_8 FILLER_12_120 ();
 sg13g2_decap_4 FILLER_12_127 ();
 sg13g2_fill_1 FILLER_12_131 ();
 sg13g2_fill_1 FILLER_12_148 ();
 sg13g2_fill_2 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_198 ();
 sg13g2_decap_4 FILLER_12_205 ();
 sg13g2_decap_4 FILLER_12_228 ();
 sg13g2_decap_4 FILLER_12_244 ();
 sg13g2_decap_8 FILLER_12_253 ();
 sg13g2_fill_2 FILLER_12_265 ();
 sg13g2_fill_1 FILLER_12_267 ();
 sg13g2_decap_4 FILLER_12_273 ();
 sg13g2_fill_2 FILLER_12_289 ();
 sg13g2_decap_8 FILLER_12_299 ();
 sg13g2_fill_2 FILLER_12_306 ();
 sg13g2_fill_2 FILLER_12_313 ();
 sg13g2_fill_1 FILLER_12_315 ();
 sg13g2_fill_2 FILLER_12_338 ();
 sg13g2_fill_1 FILLER_12_340 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_fill_1 FILLER_13_28 ();
 sg13g2_decap_4 FILLER_13_33 ();
 sg13g2_fill_2 FILLER_13_37 ();
 sg13g2_decap_4 FILLER_13_75 ();
 sg13g2_fill_2 FILLER_13_104 ();
 sg13g2_fill_1 FILLER_13_106 ();
 sg13g2_fill_1 FILLER_13_116 ();
 sg13g2_decap_4 FILLER_13_122 ();
 sg13g2_fill_1 FILLER_13_126 ();
 sg13g2_decap_4 FILLER_13_159 ();
 sg13g2_fill_2 FILLER_13_163 ();
 sg13g2_fill_2 FILLER_13_170 ();
 sg13g2_fill_1 FILLER_13_180 ();
 sg13g2_fill_2 FILLER_13_185 ();
 sg13g2_decap_8 FILLER_13_198 ();
 sg13g2_fill_2 FILLER_13_216 ();
 sg13g2_fill_1 FILLER_13_244 ();
 sg13g2_fill_2 FILLER_13_269 ();
 sg13g2_fill_1 FILLER_13_271 ();
 sg13g2_decap_8 FILLER_13_288 ();
 sg13g2_fill_2 FILLER_13_295 ();
 sg13g2_decap_4 FILLER_13_311 ();
 sg13g2_fill_2 FILLER_13_315 ();
 sg13g2_decap_4 FILLER_13_329 ();
 sg13g2_fill_2 FILLER_13_333 ();
 sg13g2_fill_1 FILLER_13_366 ();
 sg13g2_fill_1 FILLER_13_382 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_4 FILLER_14_35 ();
 sg13g2_fill_1 FILLER_14_39 ();
 sg13g2_fill_2 FILLER_14_48 ();
 sg13g2_decap_4 FILLER_14_54 ();
 sg13g2_fill_1 FILLER_14_58 ();
 sg13g2_fill_1 FILLER_14_74 ();
 sg13g2_fill_2 FILLER_14_89 ();
 sg13g2_fill_2 FILLER_14_99 ();
 sg13g2_decap_4 FILLER_14_123 ();
 sg13g2_fill_2 FILLER_14_127 ();
 sg13g2_fill_2 FILLER_14_133 ();
 sg13g2_fill_1 FILLER_14_144 ();
 sg13g2_decap_4 FILLER_14_150 ();
 sg13g2_fill_2 FILLER_14_159 ();
 sg13g2_fill_2 FILLER_14_180 ();
 sg13g2_fill_2 FILLER_14_208 ();
 sg13g2_decap_4 FILLER_14_224 ();
 sg13g2_decap_4 FILLER_14_236 ();
 sg13g2_decap_8 FILLER_14_244 ();
 sg13g2_decap_4 FILLER_14_251 ();
 sg13g2_fill_1 FILLER_14_255 ();
 sg13g2_decap_8 FILLER_14_260 ();
 sg13g2_decap_4 FILLER_14_267 ();
 sg13g2_fill_1 FILLER_14_271 ();
 sg13g2_fill_1 FILLER_14_289 ();
 sg13g2_fill_1 FILLER_14_298 ();
 sg13g2_fill_1 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_337 ();
 sg13g2_decap_4 FILLER_14_344 ();
 sg13g2_fill_2 FILLER_14_348 ();
 sg13g2_fill_1 FILLER_14_367 ();
 sg13g2_fill_2 FILLER_14_407 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_fill_1 FILLER_15_28 ();
 sg13g2_decap_4 FILLER_15_59 ();
 sg13g2_fill_1 FILLER_15_69 ();
 sg13g2_fill_2 FILLER_15_91 ();
 sg13g2_fill_1 FILLER_15_139 ();
 sg13g2_fill_1 FILLER_15_148 ();
 sg13g2_decap_4 FILLER_15_160 ();
 sg13g2_fill_2 FILLER_15_164 ();
 sg13g2_decap_4 FILLER_15_177 ();
 sg13g2_fill_2 FILLER_15_181 ();
 sg13g2_fill_2 FILLER_15_187 ();
 sg13g2_decap_8 FILLER_15_194 ();
 sg13g2_fill_2 FILLER_15_201 ();
 sg13g2_fill_1 FILLER_15_203 ();
 sg13g2_fill_2 FILLER_15_209 ();
 sg13g2_fill_1 FILLER_15_211 ();
 sg13g2_decap_8 FILLER_15_221 ();
 sg13g2_decap_4 FILLER_15_228 ();
 sg13g2_fill_2 FILLER_15_246 ();
 sg13g2_fill_2 FILLER_15_257 ();
 sg13g2_fill_1 FILLER_15_259 ();
 sg13g2_decap_4 FILLER_15_269 ();
 sg13g2_fill_1 FILLER_15_273 ();
 sg13g2_fill_2 FILLER_15_282 ();
 sg13g2_fill_1 FILLER_15_297 ();
 sg13g2_fill_2 FILLER_15_306 ();
 sg13g2_fill_2 FILLER_15_317 ();
 sg13g2_decap_8 FILLER_15_331 ();
 sg13g2_fill_1 FILLER_15_338 ();
 sg13g2_decap_4 FILLER_15_344 ();
 sg13g2_fill_2 FILLER_15_353 ();
 sg13g2_fill_1 FILLER_15_355 ();
 sg13g2_fill_1 FILLER_15_365 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_4 FILLER_16_35 ();
 sg13g2_fill_2 FILLER_16_39 ();
 sg13g2_decap_8 FILLER_16_95 ();
 sg13g2_decap_8 FILLER_16_102 ();
 sg13g2_fill_1 FILLER_16_109 ();
 sg13g2_fill_1 FILLER_16_119 ();
 sg13g2_decap_4 FILLER_16_135 ();
 sg13g2_decap_8 FILLER_16_164 ();
 sg13g2_fill_2 FILLER_16_171 ();
 sg13g2_fill_1 FILLER_16_173 ();
 sg13g2_fill_2 FILLER_16_183 ();
 sg13g2_fill_1 FILLER_16_191 ();
 sg13g2_decap_4 FILLER_16_197 ();
 sg13g2_decap_8 FILLER_16_223 ();
 sg13g2_fill_1 FILLER_16_230 ();
 sg13g2_fill_1 FILLER_16_239 ();
 sg13g2_decap_8 FILLER_16_253 ();
 sg13g2_fill_2 FILLER_16_260 ();
 sg13g2_fill_2 FILLER_16_280 ();
 sg13g2_fill_1 FILLER_16_282 ();
 sg13g2_fill_2 FILLER_16_297 ();
 sg13g2_fill_1 FILLER_16_299 ();
 sg13g2_decap_8 FILLER_16_322 ();
 sg13g2_decap_8 FILLER_16_329 ();
 sg13g2_fill_2 FILLER_16_336 ();
 sg13g2_fill_2 FILLER_16_342 ();
 sg13g2_fill_1 FILLER_16_344 ();
 sg13g2_fill_2 FILLER_16_371 ();
 sg13g2_fill_2 FILLER_16_407 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_fill_1 FILLER_17_21 ();
 sg13g2_decap_4 FILLER_17_48 ();
 sg13g2_decap_8 FILLER_17_96 ();
 sg13g2_fill_2 FILLER_17_103 ();
 sg13g2_fill_1 FILLER_17_111 ();
 sg13g2_decap_8 FILLER_17_132 ();
 sg13g2_fill_2 FILLER_17_139 ();
 sg13g2_fill_1 FILLER_17_141 ();
 sg13g2_fill_1 FILLER_17_152 ();
 sg13g2_decap_4 FILLER_17_161 ();
 sg13g2_fill_1 FILLER_17_165 ();
 sg13g2_fill_2 FILLER_17_171 ();
 sg13g2_fill_1 FILLER_17_187 ();
 sg13g2_decap_8 FILLER_17_202 ();
 sg13g2_decap_8 FILLER_17_209 ();
 sg13g2_fill_1 FILLER_17_235 ();
 sg13g2_fill_1 FILLER_17_258 ();
 sg13g2_fill_2 FILLER_17_264 ();
 sg13g2_fill_1 FILLER_17_266 ();
 sg13g2_decap_4 FILLER_17_272 ();
 sg13g2_fill_2 FILLER_17_276 ();
 sg13g2_decap_8 FILLER_17_287 ();
 sg13g2_decap_4 FILLER_17_316 ();
 sg13g2_fill_2 FILLER_17_320 ();
 sg13g2_fill_1 FILLER_17_369 ();
 sg13g2_fill_2 FILLER_17_388 ();
 sg13g2_fill_2 FILLER_17_407 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_fill_1 FILLER_18_28 ();
 sg13g2_decap_4 FILLER_18_45 ();
 sg13g2_fill_1 FILLER_18_49 ();
 sg13g2_fill_2 FILLER_18_68 ();
 sg13g2_fill_2 FILLER_18_80 ();
 sg13g2_fill_1 FILLER_18_95 ();
 sg13g2_fill_2 FILLER_18_105 ();
 sg13g2_fill_1 FILLER_18_107 ();
 sg13g2_decap_8 FILLER_18_117 ();
 sg13g2_fill_2 FILLER_18_124 ();
 sg13g2_fill_1 FILLER_18_140 ();
 sg13g2_decap_4 FILLER_18_164 ();
 sg13g2_decap_4 FILLER_18_189 ();
 sg13g2_fill_2 FILLER_18_211 ();
 sg13g2_fill_1 FILLER_18_213 ();
 sg13g2_fill_2 FILLER_18_219 ();
 sg13g2_decap_8 FILLER_18_225 ();
 sg13g2_decap_4 FILLER_18_242 ();
 sg13g2_decap_4 FILLER_18_258 ();
 sg13g2_fill_1 FILLER_18_262 ();
 sg13g2_fill_2 FILLER_18_297 ();
 sg13g2_fill_2 FILLER_18_314 ();
 sg13g2_fill_1 FILLER_18_316 ();
 sg13g2_fill_2 FILLER_18_322 ();
 sg13g2_fill_1 FILLER_18_373 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_fill_2 FILLER_19_28 ();
 sg13g2_fill_1 FILLER_19_56 ();
 sg13g2_decap_4 FILLER_19_93 ();
 sg13g2_fill_2 FILLER_19_97 ();
 sg13g2_decap_4 FILLER_19_121 ();
 sg13g2_fill_2 FILLER_19_125 ();
 sg13g2_decap_4 FILLER_19_135 ();
 sg13g2_fill_1 FILLER_19_153 ();
 sg13g2_fill_1 FILLER_19_164 ();
 sg13g2_fill_2 FILLER_19_172 ();
 sg13g2_fill_1 FILLER_19_174 ();
 sg13g2_decap_8 FILLER_19_179 ();
 sg13g2_decap_4 FILLER_19_191 ();
 sg13g2_fill_2 FILLER_19_215 ();
 sg13g2_decap_4 FILLER_19_242 ();
 sg13g2_fill_2 FILLER_19_246 ();
 sg13g2_decap_8 FILLER_19_269 ();
 sg13g2_fill_1 FILLER_19_281 ();
 sg13g2_decap_4 FILLER_19_295 ();
 sg13g2_fill_2 FILLER_19_313 ();
 sg13g2_fill_1 FILLER_19_337 ();
 sg13g2_fill_1 FILLER_19_357 ();
 sg13g2_fill_1 FILLER_19_373 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_fill_2 FILLER_20_49 ();
 sg13g2_fill_2 FILLER_20_86 ();
 sg13g2_fill_1 FILLER_20_102 ();
 sg13g2_fill_2 FILLER_20_112 ();
 sg13g2_fill_1 FILLER_20_114 ();
 sg13g2_decap_8 FILLER_20_123 ();
 sg13g2_fill_1 FILLER_20_130 ();
 sg13g2_decap_4 FILLER_20_140 ();
 sg13g2_fill_2 FILLER_20_144 ();
 sg13g2_decap_8 FILLER_20_164 ();
 sg13g2_decap_4 FILLER_20_171 ();
 sg13g2_fill_1 FILLER_20_175 ();
 sg13g2_decap_8 FILLER_20_194 ();
 sg13g2_decap_8 FILLER_20_201 ();
 sg13g2_decap_8 FILLER_20_208 ();
 sg13g2_fill_2 FILLER_20_215 ();
 sg13g2_fill_1 FILLER_20_217 ();
 sg13g2_fill_1 FILLER_20_222 ();
 sg13g2_decap_8 FILLER_20_244 ();
 sg13g2_fill_2 FILLER_20_251 ();
 sg13g2_fill_1 FILLER_20_267 ();
 sg13g2_fill_1 FILLER_20_277 ();
 sg13g2_decap_8 FILLER_20_294 ();
 sg13g2_decap_8 FILLER_20_301 ();
 sg13g2_decap_4 FILLER_20_316 ();
 sg13g2_decap_4 FILLER_20_326 ();
 sg13g2_fill_2 FILLER_20_354 ();
 sg13g2_fill_2 FILLER_20_374 ();
 sg13g2_fill_1 FILLER_20_376 ();
 sg13g2_fill_2 FILLER_20_407 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_4 FILLER_21_35 ();
 sg13g2_fill_1 FILLER_21_39 ();
 sg13g2_fill_2 FILLER_21_66 ();
 sg13g2_fill_1 FILLER_21_73 ();
 sg13g2_fill_2 FILLER_21_94 ();
 sg13g2_fill_1 FILLER_21_96 ();
 sg13g2_fill_1 FILLER_21_116 ();
 sg13g2_decap_4 FILLER_21_125 ();
 sg13g2_fill_2 FILLER_21_129 ();
 sg13g2_decap_8 FILLER_21_141 ();
 sg13g2_decap_4 FILLER_21_162 ();
 sg13g2_fill_2 FILLER_21_190 ();
 sg13g2_fill_2 FILLER_21_197 ();
 sg13g2_fill_1 FILLER_21_204 ();
 sg13g2_fill_2 FILLER_21_209 ();
 sg13g2_fill_1 FILLER_21_211 ();
 sg13g2_fill_2 FILLER_21_217 ();
 sg13g2_fill_1 FILLER_21_229 ();
 sg13g2_fill_2 FILLER_21_235 ();
 sg13g2_fill_1 FILLER_21_237 ();
 sg13g2_decap_4 FILLER_21_260 ();
 sg13g2_fill_1 FILLER_21_264 ();
 sg13g2_fill_1 FILLER_21_278 ();
 sg13g2_fill_2 FILLER_21_290 ();
 sg13g2_fill_1 FILLER_21_292 ();
 sg13g2_decap_4 FILLER_21_321 ();
 sg13g2_fill_2 FILLER_21_325 ();
 sg13g2_fill_1 FILLER_21_343 ();
 sg13g2_fill_2 FILLER_21_354 ();
 sg13g2_fill_1 FILLER_21_356 ();
 sg13g2_fill_1 FILLER_21_380 ();
 sg13g2_fill_2 FILLER_21_407 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_fill_2 FILLER_22_42 ();
 sg13g2_fill_1 FILLER_22_44 ();
 sg13g2_fill_2 FILLER_22_66 ();
 sg13g2_fill_2 FILLER_22_97 ();
 sg13g2_fill_1 FILLER_22_105 ();
 sg13g2_decap_8 FILLER_22_116 ();
 sg13g2_fill_2 FILLER_22_123 ();
 sg13g2_decap_8 FILLER_22_143 ();
 sg13g2_decap_8 FILLER_22_150 ();
 sg13g2_fill_1 FILLER_22_161 ();
 sg13g2_fill_2 FILLER_22_221 ();
 sg13g2_fill_1 FILLER_22_223 ();
 sg13g2_fill_1 FILLER_22_232 ();
 sg13g2_decap_8 FILLER_22_238 ();
 sg13g2_decap_4 FILLER_22_245 ();
 sg13g2_fill_2 FILLER_22_249 ();
 sg13g2_decap_4 FILLER_22_269 ();
 sg13g2_fill_1 FILLER_22_273 ();
 sg13g2_decap_8 FILLER_22_292 ();
 sg13g2_decap_8 FILLER_22_318 ();
 sg13g2_fill_1 FILLER_22_325 ();
 sg13g2_fill_2 FILLER_22_341 ();
 sg13g2_fill_1 FILLER_22_343 ();
 sg13g2_fill_2 FILLER_22_362 ();
 sg13g2_fill_1 FILLER_22_364 ();
 sg13g2_fill_2 FILLER_22_377 ();
 sg13g2_fill_1 FILLER_22_379 ();
 sg13g2_fill_2 FILLER_22_406 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_fill_1 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_34 ();
 sg13g2_decap_4 FILLER_23_41 ();
 sg13g2_fill_2 FILLER_23_45 ();
 sg13g2_fill_2 FILLER_23_73 ();
 sg13g2_decap_4 FILLER_23_118 ();
 sg13g2_fill_1 FILLER_23_122 ();
 sg13g2_fill_1 FILLER_23_153 ();
 sg13g2_fill_2 FILLER_23_166 ();
 sg13g2_fill_1 FILLER_23_168 ();
 sg13g2_decap_8 FILLER_23_193 ();
 sg13g2_decap_8 FILLER_23_209 ();
 sg13g2_decap_4 FILLER_23_216 ();
 sg13g2_fill_1 FILLER_23_220 ();
 sg13g2_fill_2 FILLER_23_243 ();
 sg13g2_decap_8 FILLER_23_255 ();
 sg13g2_decap_4 FILLER_23_262 ();
 sg13g2_fill_1 FILLER_23_266 ();
 sg13g2_decap_4 FILLER_23_272 ();
 sg13g2_fill_1 FILLER_23_276 ();
 sg13g2_decap_8 FILLER_23_281 ();
 sg13g2_decap_8 FILLER_23_314 ();
 sg13g2_decap_8 FILLER_23_321 ();
 sg13g2_fill_2 FILLER_23_360 ();
 sg13g2_fill_1 FILLER_23_362 ();
 sg13g2_fill_2 FILLER_23_377 ();
 sg13g2_decap_4 FILLER_23_405 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_fill_2 FILLER_24_14 ();
 sg13g2_fill_1 FILLER_24_16 ();
 sg13g2_fill_1 FILLER_24_21 ();
 sg13g2_fill_2 FILLER_24_31 ();
 sg13g2_fill_1 FILLER_24_33 ();
 sg13g2_decap_4 FILLER_24_47 ();
 sg13g2_fill_2 FILLER_24_60 ();
 sg13g2_fill_1 FILLER_24_62 ();
 sg13g2_fill_2 FILLER_24_110 ();
 sg13g2_decap_4 FILLER_24_118 ();
 sg13g2_fill_2 FILLER_24_122 ();
 sg13g2_decap_8 FILLER_24_144 ();
 sg13g2_fill_2 FILLER_24_151 ();
 sg13g2_fill_2 FILLER_24_157 ();
 sg13g2_fill_1 FILLER_24_159 ();
 sg13g2_fill_1 FILLER_24_165 ();
 sg13g2_decap_8 FILLER_24_182 ();
 sg13g2_decap_4 FILLER_24_207 ();
 sg13g2_fill_2 FILLER_24_211 ();
 sg13g2_decap_8 FILLER_24_227 ();
 sg13g2_fill_1 FILLER_24_234 ();
 sg13g2_decap_4 FILLER_24_249 ();
 sg13g2_fill_2 FILLER_24_253 ();
 sg13g2_fill_1 FILLER_24_281 ();
 sg13g2_fill_2 FILLER_24_315 ();
 sg13g2_fill_1 FILLER_24_317 ();
 sg13g2_fill_2 FILLER_24_323 ();
 sg13g2_decap_8 FILLER_24_331 ();
 sg13g2_fill_1 FILLER_24_338 ();
 sg13g2_decap_4 FILLER_24_365 ();
 sg13g2_fill_1 FILLER_24_369 ();
 sg13g2_fill_1 FILLER_24_378 ();
 sg13g2_decap_4 FILLER_25_0 ();
 sg13g2_fill_2 FILLER_25_4 ();
 sg13g2_fill_1 FILLER_25_147 ();
 sg13g2_fill_2 FILLER_25_174 ();
 sg13g2_fill_1 FILLER_25_193 ();
 sg13g2_decap_4 FILLER_25_199 ();
 sg13g2_fill_1 FILLER_25_203 ();
 sg13g2_fill_1 FILLER_25_213 ();
 sg13g2_fill_2 FILLER_25_222 ();
 sg13g2_fill_1 FILLER_25_224 ();
 sg13g2_decap_4 FILLER_25_281 ();
 sg13g2_fill_2 FILLER_25_297 ();
 sg13g2_decap_8 FILLER_25_323 ();
 sg13g2_fill_2 FILLER_25_330 ();
 sg13g2_fill_2 FILLER_25_341 ();
 sg13g2_decap_4 FILLER_25_356 ();
 sg13g2_fill_2 FILLER_25_379 ();
 sg13g2_fill_2 FILLER_25_407 ();
 sg13g2_fill_1 FILLER_26_0 ();
 sg13g2_fill_1 FILLER_26_27 ();
 sg13g2_decap_4 FILLER_26_49 ();
 sg13g2_fill_1 FILLER_26_57 ();
 sg13g2_decap_4 FILLER_26_62 ();
 sg13g2_fill_1 FILLER_26_66 ();
 sg13g2_fill_2 FILLER_26_78 ();
 sg13g2_decap_8 FILLER_26_119 ();
 sg13g2_fill_1 FILLER_26_126 ();
 sg13g2_fill_2 FILLER_26_132 ();
 sg13g2_fill_1 FILLER_26_134 ();
 sg13g2_fill_1 FILLER_26_146 ();
 sg13g2_fill_2 FILLER_26_167 ();
 sg13g2_fill_1 FILLER_26_169 ();
 sg13g2_decap_8 FILLER_26_191 ();
 sg13g2_fill_2 FILLER_26_198 ();
 sg13g2_fill_1 FILLER_26_200 ();
 sg13g2_decap_8 FILLER_26_208 ();
 sg13g2_decap_8 FILLER_26_215 ();
 sg13g2_decap_8 FILLER_26_222 ();
 sg13g2_decap_4 FILLER_26_229 ();
 sg13g2_fill_2 FILLER_26_233 ();
 sg13g2_decap_4 FILLER_26_246 ();
 sg13g2_fill_1 FILLER_26_250 ();
 sg13g2_decap_8 FILLER_26_255 ();
 sg13g2_fill_2 FILLER_26_262 ();
 sg13g2_fill_1 FILLER_26_264 ();
 sg13g2_decap_4 FILLER_26_274 ();
 sg13g2_fill_2 FILLER_26_278 ();
 sg13g2_fill_2 FILLER_26_293 ();
 sg13g2_fill_1 FILLER_26_338 ();
 sg13g2_fill_2 FILLER_26_375 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_fill_2 FILLER_27_7 ();
 sg13g2_fill_2 FILLER_27_73 ();
 sg13g2_fill_1 FILLER_27_121 ();
 sg13g2_fill_2 FILLER_27_148 ();
 sg13g2_fill_1 FILLER_27_150 ();
 sg13g2_decap_8 FILLER_27_169 ();
 sg13g2_fill_2 FILLER_27_211 ();
 sg13g2_fill_2 FILLER_27_234 ();
 sg13g2_fill_1 FILLER_27_266 ();
 sg13g2_fill_2 FILLER_27_271 ();
 sg13g2_fill_1 FILLER_27_273 ();
 sg13g2_fill_1 FILLER_27_306 ();
 sg13g2_fill_1 FILLER_27_311 ();
 sg13g2_decap_8 FILLER_27_317 ();
 sg13g2_fill_2 FILLER_27_324 ();
 sg13g2_decap_4 FILLER_27_354 ();
 sg13g2_fill_2 FILLER_27_407 ();
 sg13g2_decap_4 FILLER_28_0 ();
 sg13g2_fill_2 FILLER_28_30 ();
 sg13g2_fill_1 FILLER_28_65 ();
 sg13g2_fill_2 FILLER_28_75 ();
 sg13g2_fill_1 FILLER_28_77 ();
 sg13g2_fill_2 FILLER_28_100 ();
 sg13g2_fill_2 FILLER_28_139 ();
 sg13g2_fill_1 FILLER_28_141 ();
 sg13g2_fill_2 FILLER_28_146 ();
 sg13g2_fill_1 FILLER_28_148 ();
 sg13g2_decap_8 FILLER_28_190 ();
 sg13g2_decap_8 FILLER_28_214 ();
 sg13g2_decap_4 FILLER_28_221 ();
 sg13g2_fill_2 FILLER_28_258 ();
 sg13g2_fill_1 FILLER_28_299 ();
 sg13g2_fill_1 FILLER_28_326 ();
 sg13g2_fill_2 FILLER_28_351 ();
 sg13g2_fill_2 FILLER_28_359 ();
 sg13g2_fill_2 FILLER_28_375 ();
 sg13g2_fill_1 FILLER_28_377 ();
 sg13g2_fill_2 FILLER_28_390 ();
 sg13g2_fill_1 FILLER_28_392 ();
 sg13g2_fill_2 FILLER_29_0 ();
 sg13g2_fill_1 FILLER_29_2 ();
 sg13g2_fill_2 FILLER_29_29 ();
 sg13g2_fill_1 FILLER_29_36 ();
 sg13g2_fill_1 FILLER_29_89 ();
 sg13g2_fill_1 FILLER_29_102 ();
 sg13g2_fill_1 FILLER_29_112 ();
 sg13g2_fill_2 FILLER_29_157 ();
 sg13g2_fill_2 FILLER_29_185 ();
 sg13g2_fill_1 FILLER_29_200 ();
 sg13g2_fill_1 FILLER_29_236 ();
 sg13g2_fill_1 FILLER_29_260 ();
 sg13g2_fill_1 FILLER_29_274 ();
 sg13g2_fill_1 FILLER_29_296 ();
 sg13g2_fill_2 FILLER_29_320 ();
 sg13g2_fill_2 FILLER_29_332 ();
 sg13g2_fill_2 FILLER_29_343 ();
 sg13g2_fill_1 FILLER_29_345 ();
 sg13g2_fill_2 FILLER_29_384 ();
 sg13g2_fill_1 FILLER_29_386 ();
 sg13g2_decap_4 FILLER_30_0 ();
 sg13g2_fill_2 FILLER_30_68 ();
 sg13g2_fill_2 FILLER_30_82 ();
 sg13g2_fill_1 FILLER_30_97 ();
 sg13g2_fill_2 FILLER_30_133 ();
 sg13g2_fill_2 FILLER_30_246 ();
 sg13g2_fill_1 FILLER_30_248 ();
 sg13g2_fill_1 FILLER_30_254 ();
 sg13g2_fill_2 FILLER_30_264 ();
 sg13g2_fill_1 FILLER_30_271 ();
 sg13g2_fill_2 FILLER_30_298 ();
 sg13g2_fill_1 FILLER_30_300 ();
 sg13g2_fill_2 FILLER_30_357 ();
 sg13g2_fill_1 FILLER_30_372 ();
 sg13g2_fill_2 FILLER_30_391 ();
 sg13g2_fill_2 FILLER_30_406 ();
 sg13g2_fill_1 FILLER_30_408 ();
 sg13g2_fill_1 FILLER_31_0 ();
 sg13g2_fill_2 FILLER_31_36 ();
 sg13g2_fill_1 FILLER_31_47 ();
 sg13g2_fill_1 FILLER_31_62 ();
 sg13g2_fill_1 FILLER_31_74 ();
 sg13g2_fill_1 FILLER_31_101 ();
 sg13g2_fill_1 FILLER_31_107 ();
 sg13g2_fill_1 FILLER_31_127 ();
 sg13g2_fill_1 FILLER_31_186 ();
 sg13g2_fill_1 FILLER_31_191 ();
 sg13g2_fill_1 FILLER_31_228 ();
 sg13g2_fill_1 FILLER_31_238 ();
 sg13g2_fill_2 FILLER_31_296 ();
 sg13g2_fill_2 FILLER_31_347 ();
 sg13g2_fill_1 FILLER_31_349 ();
 sg13g2_fill_2 FILLER_31_358 ();
 sg13g2_fill_1 FILLER_31_360 ();
 sg13g2_fill_2 FILLER_31_377 ();
 sg13g2_fill_2 FILLER_32_0 ();
 sg13g2_fill_1 FILLER_32_28 ();
 sg13g2_fill_1 FILLER_32_34 ();
 sg13g2_fill_1 FILLER_32_83 ();
 sg13g2_fill_1 FILLER_32_110 ();
 sg13g2_fill_1 FILLER_32_131 ();
 sg13g2_fill_1 FILLER_32_201 ();
 sg13g2_fill_2 FILLER_32_220 ();
 sg13g2_fill_1 FILLER_32_222 ();
 sg13g2_fill_1 FILLER_32_323 ();
 sg13g2_fill_1 FILLER_32_340 ();
 sg13g2_fill_2 FILLER_32_360 ();
 sg13g2_fill_1 FILLER_32_408 ();
 sg13g2_fill_2 FILLER_33_0 ();
 sg13g2_fill_1 FILLER_33_103 ();
 sg13g2_fill_2 FILLER_33_187 ();
 sg13g2_fill_2 FILLER_33_226 ();
 sg13g2_fill_2 FILLER_33_249 ();
 sg13g2_fill_1 FILLER_33_251 ();
 sg13g2_fill_2 FILLER_33_264 ();
 sg13g2_decap_4 FILLER_33_301 ();
 sg13g2_fill_2 FILLER_33_326 ();
 sg13g2_fill_2 FILLER_33_380 ();
 sg13g2_fill_1 FILLER_33_382 ();
 sg13g2_fill_1 FILLER_34_0 ();
 sg13g2_fill_2 FILLER_34_125 ();
 sg13g2_fill_1 FILLER_34_141 ();
 sg13g2_fill_2 FILLER_34_147 ();
 sg13g2_fill_1 FILLER_34_163 ();
 sg13g2_fill_2 FILLER_34_169 ();
 sg13g2_decap_4 FILLER_34_250 ();
 sg13g2_fill_2 FILLER_34_263 ();
 sg13g2_fill_1 FILLER_34_265 ();
 sg13g2_fill_1 FILLER_34_276 ();
 sg13g2_fill_1 FILLER_34_333 ();
 sg13g2_fill_1 FILLER_34_354 ();
 sg13g2_fill_1 FILLER_34_364 ();
 sg13g2_fill_1 FILLER_34_408 ();
 sg13g2_decap_4 FILLER_35_0 ();
 sg13g2_fill_2 FILLER_35_105 ();
 sg13g2_fill_1 FILLER_35_133 ();
 sg13g2_fill_2 FILLER_35_173 ();
 sg13g2_fill_2 FILLER_35_200 ();
 sg13g2_decap_4 FILLER_35_211 ();
 sg13g2_fill_1 FILLER_35_256 ();
 sg13g2_fill_2 FILLER_35_269 ();
 sg13g2_decap_4 FILLER_35_281 ();
 sg13g2_fill_1 FILLER_35_295 ();
 sg13g2_fill_1 FILLER_35_339 ();
 sg13g2_fill_2 FILLER_35_353 ();
 sg13g2_fill_1 FILLER_35_408 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_4 FILLER_36_7 ();
 sg13g2_fill_1 FILLER_36_11 ();
 sg13g2_fill_2 FILLER_36_131 ();
 sg13g2_fill_2 FILLER_36_142 ();
 sg13g2_fill_1 FILLER_36_144 ();
 sg13g2_decap_4 FILLER_36_226 ();
 sg13g2_fill_2 FILLER_36_230 ();
 sg13g2_fill_1 FILLER_36_239 ();
 sg13g2_decap_4 FILLER_36_249 ();
 sg13g2_fill_2 FILLER_36_256 ();
 sg13g2_decap_4 FILLER_36_265 ();
 sg13g2_fill_1 FILLER_36_287 ();
 sg13g2_fill_2 FILLER_36_326 ();
 sg13g2_fill_1 FILLER_36_328 ();
 sg13g2_fill_2 FILLER_36_369 ();
 sg13g2_fill_1 FILLER_36_382 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_fill_2 FILLER_37_14 ();
 sg13g2_fill_2 FILLER_37_127 ();
 sg13g2_fill_1 FILLER_37_183 ();
 sg13g2_fill_2 FILLER_37_198 ();
 sg13g2_fill_1 FILLER_37_266 ();
 sg13g2_fill_2 FILLER_37_300 ();
 sg13g2_fill_1 FILLER_37_302 ();
 sg13g2_fill_2 FILLER_37_356 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_fill_1 FILLER_38_21 ();
 sg13g2_fill_1 FILLER_38_68 ();
 sg13g2_decap_8 FILLER_38_217 ();
 sg13g2_fill_1 FILLER_38_224 ();
 sg13g2_decap_8 FILLER_38_229 ();
 sg13g2_decap_8 FILLER_38_236 ();
 sg13g2_fill_2 FILLER_38_243 ();
 sg13g2_decap_4 FILLER_38_249 ();
 sg13g2_fill_1 FILLER_38_273 ();
 sg13g2_fill_1 FILLER_38_292 ();
 sg13g2_fill_1 FILLER_38_408 ();
 assign uio_oe[0] = net13;
 assign uio_oe[1] = net14;
 assign uio_oe[2] = net15;
 assign uio_oe[3] = net16;
 assign uio_oe[4] = net17;
 assign uio_oe[5] = net18;
 assign uio_oe[6] = net137;
 assign uio_oe[7] = net138;
 assign uio_out[0] = net19;
 assign uio_out[1] = net20;
 assign uio_out[2] = net21;
 assign uio_out[3] = net22;
 assign uio_out[4] = net23;
 assign uio_out[5] = net24;
endmodule

module tt_um_whynot (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire \main._w_demo_audio1 ;
 wire \main._w_demo_video_hs ;
 wire \main._w_demo_video_vs ;
 wire \main.demo._d_addr[0] ;
 wire \main.demo._d_addr[1] ;
 wire \main.demo._d_addr[2] ;
 wire \main.demo._d_addr[3] ;
 wire \main.demo._d_addr[4] ;
 wire \main.demo._d_addr[5] ;
 wire \main.demo._d_addr[6] ;
 wire \main.demo._d_addr[7] ;
 wire \main.demo._d_addr[8] ;
 wire \main.demo._d_addr[9] ;
 wire \main.demo._q_addr[0] ;
 wire \main.demo._q_addr[1] ;
 wire \main.demo._q_addr[2] ;
 wire \main.demo._q_addr[3] ;
 wire \main.demo._q_addr[4] ;
 wire \main.demo._q_addr[5] ;
 wire \main.demo._q_addr[6] ;
 wire \main.demo._q_addr[7] ;
 wire \main.demo._q_addr[8] ;
 wire \main.demo._q_addr[9] ;
 wire \main.demo._q_frame[0] ;
 wire \main.demo._q_frame[1] ;
 wire \main.demo._q_frame[2] ;
 wire \main.demo._q_frame[3] ;
 wire \main.demo._q_frame[4] ;
 wire \main.demo._q_frame[5] ;
 wire \main.demo._q_frame[6] ;
 wire \main.demo._q_frame[7] ;
 wire \main.demo._q_frame[8] ;
 wire \main.demo._q_frame[9] ;
 wire \main.demo._q_prev_hs ;
 wire \main.demo._q_prev_vs ;
 wire \main.demo._q_uT[0] ;
 wire \main.demo._q_uT[10] ;
 wire \main.demo._q_uT[11] ;
 wire \main.demo._q_uT[1] ;
 wire \main.demo._q_uT[2] ;
 wire \main.demo._q_uT[3] ;
 wire \main.demo._q_uT[4] ;
 wire \main.demo._q_uT[5] ;
 wire \main.demo._q_uT[6] ;
 wire \main.demo._q_uT[7] ;
 wire \main.demo._q_uT[8] ;
 wire \main.demo._q_uT[9] ;
 wire \main.demo._q_u[0] ;
 wire \main.demo._q_u[1] ;
 wire \main.demo._q_u[2] ;
 wire \main.demo._q_u[3] ;
 wire \main.demo._q_u[4] ;
 wire \main.demo._q_u[5] ;
 wire \main.demo._q_u[6] ;
 wire \main.demo._q_u[7] ;
 wire \main.demo._q_vT[0] ;
 wire \main.demo._q_vT[10] ;
 wire \main.demo._q_vT[11] ;
 wire \main.demo._q_vT[1] ;
 wire \main.demo._q_vT[2] ;
 wire \main.demo._q_vT[3] ;
 wire \main.demo._q_vT[4] ;
 wire \main.demo._q_vT[5] ;
 wire \main.demo._q_vT[6] ;
 wire \main.demo._q_vT[7] ;
 wire \main.demo._q_vT[8] ;
 wire \main.demo._q_vT[9] ;
 wire \main.demo._q_v[0] ;
 wire \main.demo._q_v[1] ;
 wire \main.demo._q_v[2] ;
 wire \main.demo._q_v[3] ;
 wire \main.demo._q_v[4] ;
 wire \main.demo._q_v[5] ;
 wire \main.demo._q_v[6] ;
 wire \main.demo._q_v[7] ;
 wire \main.demo._t___block_1_p4[0] ;
 wire \main.demo._t___block_1_p4[1] ;
 wire \main.demo._t___block_1_p4[2] ;
 wire \main.demo._t___block_1_p4[3] ;
 wire \main.demo._w_vga_active ;
 wire \main.demo.vga._d_active ;
 wire \main.demo.vga._d_vblank ;
 wire \main.demo.vga._q_active_h ;
 wire \main.demo.vga._q_active_v ;
 wire \main.demo.vga._q_xcount[0] ;
 wire \main.demo.vga._q_xcount[10] ;
 wire \main.demo.vga._q_xcount[1] ;
 wire \main.demo.vga._q_xcount[2] ;
 wire \main.demo.vga._q_xcount[3] ;
 wire \main.demo.vga._q_xcount[4] ;
 wire \main.demo.vga._q_xcount[5] ;
 wire \main.demo.vga._q_xcount[6] ;
 wire \main.demo.vga._q_xcount[7] ;
 wire \main.demo.vga._q_xcount[8] ;
 wire \main.demo.vga._q_xcount[9] ;
 wire \main.demo.vga._q_ycount[0] ;
 wire \main.demo.vga._q_ycount[1] ;
 wire \main.demo.vga._q_ycount[2] ;
 wire \main.demo.vga._q_ycount[3] ;
 wire \main.demo.vga._q_ycount[4] ;
 wire \main.demo.vga._q_ycount[5] ;
 wire \main.demo.vga._q_ycount[6] ;
 wire \main.demo.vga._q_ycount[7] ;
 wire \main.demo.vga._q_ycount[8] ;
 wire \main.demo.zic._d_clock_count[0] ;
 wire \main.demo.zic._q_clock_count[0] ;
 wire \main.demo.zic._q_clock_count[1] ;
 wire \main.demo.zic._q_clock_count[2] ;
 wire \main.demo.zic._q_clock_count[3] ;
 wire \main.demo.zic._q_clock_count[4] ;
 wire \main.demo.zic._q_clock_count[5] ;
 wire \main.demo.zic._q_clock_count[6] ;
 wire \main.demo.zic._q_clock_count[7] ;
 wire \main.demo.zic._q_clock_count[8] ;
 wire \main.demo.zic._q_idx[0] ;
 wire \main.demo.zic._q_idx[1] ;
 wire \main.demo.zic._q_idx[2] ;
 wire \main.demo.zic._q_idx[3] ;
 wire \main.demo.zic._q_idx[4] ;
 wire \main.demo.zic._q_qpos[0] ;
 wire \main.demo.zic._q_qpos[10] ;
 wire \main.demo.zic._q_qpos[11] ;
 wire \main.demo.zic._q_qpos[12] ;
 wire \main.demo.zic._q_qpos[1] ;
 wire \main.demo.zic._q_qpos[2] ;
 wire \main.demo.zic._q_qpos[3] ;
 wire \main.demo.zic._q_qpos[4] ;
 wire \main.demo.zic._q_qpos[5] ;
 wire \main.demo.zic._q_qpos[6] ;
 wire \main.demo.zic._q_qpos[7] ;
 wire \main.demo.zic._q_qpos[8] ;
 wire \main.demo.zic._q_qpos[9] ;
 wire \main.demo.zic._q_rythm_count[0] ;
 wire \main.demo.zic._q_rythm_count[10] ;
 wire \main.demo.zic._q_rythm_count[11] ;
 wire \main.demo.zic._q_rythm_count[12] ;
 wire \main.demo.zic._q_rythm_count[1] ;
 wire \main.demo.zic._q_rythm_count[2] ;
 wire \main.demo.zic._q_rythm_count[3] ;
 wire \main.demo.zic._q_rythm_count[4] ;
 wire \main.demo.zic._q_rythm_count[5] ;
 wire \main.demo.zic._q_rythm_count[6] ;
 wire \main.demo.zic._q_rythm_count[7] ;
 wire \main.demo.zic._q_rythm_count[8] ;
 wire \main.demo.zic._q_rythm_count[9] ;
 wire \main.demo.zic._q_squ_env[0] ;
 wire \main.demo.zic._q_squ_env[1] ;
 wire \main.demo.zic._q_squ_env[2] ;
 wire \main.demo.zic._q_squ_env[3] ;
 wire \main.demo.zic._q_squ_env[4] ;
 wire \main.demo.zic._q_squ_env[5] ;
 wire rst_n_q;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire clknet_0_clk;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net1;
 wire net2;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_5_0__leaf_clk;
 wire clknet_5_1__leaf_clk;
 wire clknet_5_2__leaf_clk;
 wire clknet_5_3__leaf_clk;
 wire clknet_5_4__leaf_clk;
 wire clknet_5_5__leaf_clk;
 wire clknet_5_6__leaf_clk;
 wire clknet_5_7__leaf_clk;
 wire clknet_5_8__leaf_clk;
 wire clknet_5_9__leaf_clk;
 wire clknet_5_10__leaf_clk;
 wire clknet_5_11__leaf_clk;
 wire clknet_5_12__leaf_clk;
 wire clknet_5_13__leaf_clk;
 wire clknet_5_14__leaf_clk;
 wire clknet_5_15__leaf_clk;
 wire clknet_5_16__leaf_clk;
 wire clknet_5_17__leaf_clk;
 wire clknet_5_18__leaf_clk;
 wire clknet_5_19__leaf_clk;
 wire clknet_5_20__leaf_clk;
 wire clknet_5_21__leaf_clk;
 wire clknet_5_22__leaf_clk;
 wire clknet_5_23__leaf_clk;
 wire clknet_5_24__leaf_clk;
 wire clknet_5_25__leaf_clk;
 wire clknet_5_26__leaf_clk;
 wire clknet_5_27__leaf_clk;
 wire clknet_5_28__leaf_clk;
 wire clknet_5_29__leaf_clk;
 wire clknet_5_30__leaf_clk;
 wire clknet_5_31__leaf_clk;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;

 sg13g2_inv_1 _1543_ (.Y(_0591_),
    .A(net390));
 sg13g2_inv_1 _1544_ (.Y(_0592_),
    .A(net365));
 sg13g2_inv_1 _1545_ (.Y(_0593_),
    .A(net305));
 sg13g2_inv_1 _1546_ (.Y(_0594_),
    .A(net318));
 sg13g2_inv_1 _1547_ (.Y(_0595_),
    .A(net287));
 sg13g2_inv_1 _1548_ (.Y(_0596_),
    .A(net189));
 sg13g2_inv_1 _1549_ (.Y(_0597_),
    .A(net395));
 sg13g2_inv_1 _1550_ (.Y(_0598_),
    .A(net251));
 sg13g2_inv_1 _1551_ (.Y(_0599_),
    .A(net169));
 sg13g2_inv_1 _1552_ (.Y(_0600_),
    .A(\main.demo.zic._q_idx[3] ));
 sg13g2_inv_1 _1553_ (.Y(_0601_),
    .A(\main.demo.zic._q_idx[2] ));
 sg13g2_inv_1 _1554_ (.Y(_0602_),
    .A(\main.demo.zic._q_idx[4] ));
 sg13g2_inv_1 _1555_ (.Y(_0603_),
    .A(net383));
 sg13g2_inv_1 _1556_ (.Y(_0604_),
    .A(net346));
 sg13g2_inv_1 _1557_ (.Y(_0605_),
    .A(net610));
 sg13g2_inv_1 _1558_ (.Y(_0606_),
    .A(net600));
 sg13g2_inv_2 _1559_ (.Y(_0607_),
    .A(net599));
 sg13g2_inv_1 _1560_ (.Y(_0608_),
    .A(net307));
 sg13g2_inv_1 _1561_ (.Y(_0609_),
    .A(_0002_));
 sg13g2_inv_2 _1562_ (.Y(_0610_),
    .A(\main.demo._q_frame[1] ));
 sg13g2_inv_1 _1563_ (.Y(_0611_),
    .A(\main.demo._q_frame[6] ));
 sg13g2_inv_1 _1564_ (.Y(_0612_),
    .A(_0004_));
 sg13g2_inv_1 _1565_ (.Y(_0613_),
    .A(\main.demo._q_u[6] ));
 sg13g2_inv_1 _1566_ (.Y(_0614_),
    .A(\main.demo._q_uT[2] ));
 sg13g2_or3_2 _1567_ (.A(\main.demo.vga._q_xcount[4] ),
    .B(\main.demo.vga._q_xcount[5] ),
    .C(\main.demo.vga._q_xcount[6] ),
    .X(_0615_));
 sg13g2_nor2_1 _1568_ (.A(\main.demo.vga._q_xcount[8] ),
    .B(\main.demo.vga._q_xcount[10] ),
    .Y(_0616_));
 sg13g2_nand3_1 _1569_ (.B(\main.demo.vga._q_xcount[9] ),
    .C(_0616_),
    .A(net220),
    .Y(_0617_));
 sg13g2_nor2_1 _1570_ (.A(net192),
    .B(net193),
    .Y(_0618_));
 sg13g2_or4_2 _1571_ (.A(\main.demo.vga._q_xcount[0] ),
    .B(\main.demo.vga._q_xcount[1] ),
    .C(\main.demo.vga._q_xcount[2] ),
    .D(\main.demo.vga._q_xcount[3] ),
    .X(_0619_));
 sg13g2_nor3_2 _1572_ (.A(_0615_),
    .B(_0617_),
    .C(_0619_),
    .Y(_0620_));
 sg13g2_or3_2 _1573_ (.A(_0615_),
    .B(_0617_),
    .C(_0619_),
    .X(_0621_));
 sg13g2_nor3_1 _1574_ (.A(_0615_),
    .B(_0617_),
    .C(_0619_),
    .Y(_0622_));
 sg13g2_nor2_1 _1575_ (.A(net220),
    .B(_0619_),
    .Y(_0623_));
 sg13g2_nor4_1 _1576_ (.A(net378),
    .B(net237),
    .C(net353),
    .D(_0615_),
    .Y(_0624_));
 sg13g2_a22oi_1 _1577_ (.Y(_0625_),
    .B1(_0623_),
    .B2(_0624_),
    .A2(_0621_),
    .A1(net223));
 sg13g2_nor4_1 _1578_ (.A(\main.demo.vga._q_ycount[3] ),
    .B(\main.demo.vga._q_ycount[2] ),
    .C(\main.demo.vga._q_ycount[1] ),
    .D(\main.demo.vga._q_ycount[0] ),
    .Y(_0626_));
 sg13g2_nor2_1 _1579_ (.A(\main.demo.vga._q_ycount[4] ),
    .B(net364),
    .Y(_0627_));
 sg13g2_and4_1 _1580_ (.A(\main.demo.vga._q_ycount[8] ),
    .B(\main.demo.vga._q_ycount[7] ),
    .C(\main.demo.vga._q_ycount[6] ),
    .D(\main.demo.vga._q_ycount[5] ),
    .X(_0628_));
 sg13g2_and3_1 _1581_ (.X(_0629_),
    .A(_0626_),
    .B(_0627_),
    .C(_0628_));
 sg13g2_nor4_1 _1582_ (.A(\main.demo.vga._q_ycount[8] ),
    .B(\main.demo.vga._q_ycount[7] ),
    .C(\main.demo.vga._q_ycount[6] ),
    .D(\main.demo.vga._q_ycount[5] ),
    .Y(_0630_));
 sg13g2_nand3_1 _1583_ (.B(_0627_),
    .C(_0630_),
    .A(_0626_),
    .Y(_0631_));
 sg13g2_o21ai_1 _1584_ (.B1(_0631_),
    .Y(_0632_),
    .A1(_0608_),
    .A2(_0629_));
 sg13g2_nor2b_1 _1585_ (.A(net224),
    .B_N(_0632_),
    .Y(\main.demo.vga._d_active ));
 sg13g2_nor3_1 _1586_ (.A(\main.demo.zic._q_squ_env[5] ),
    .B(\main.demo.zic._q_squ_env[4] ),
    .C(\main.demo.zic._q_squ_env[3] ),
    .Y(_0633_));
 sg13g2_nor2_2 _1587_ (.A(\main.demo.zic._q_qpos[12] ),
    .B(_0633_),
    .Y(_0634_));
 sg13g2_nor2_1 _1588_ (.A(_0007_),
    .B(_0008_),
    .Y(_0635_));
 sg13g2_nand4_1 _1589_ (.B(\main.demo.zic._q_clock_count[4] ),
    .C(_0634_),
    .A(\main.demo.zic._q_clock_count[2] ),
    .Y(_0636_),
    .D(_0635_));
 sg13g2_o21ai_1 _1590_ (.B1(\main.demo.zic._q_squ_env[5] ),
    .Y(_0637_),
    .A1(\main.demo.zic._q_squ_env[4] ),
    .A2(\main.demo.zic._q_squ_env[3] ));
 sg13g2_a22oi_1 _1591_ (.Y(_0638_),
    .B1(_0634_),
    .B2(_0637_),
    .A2(_0609_),
    .A1(\main.demo.zic._q_qpos[12] ));
 sg13g2_or2_1 _1592_ (.X(_0639_),
    .B(_0638_),
    .A(\main.demo.zic._q_clock_count[1] ));
 sg13g2_xor2_1 _1593_ (.B(\main.demo.zic._q_squ_env[3] ),
    .A(\main.demo.zic._q_squ_env[4] ),
    .X(_0640_));
 sg13g2_nor2_1 _1594_ (.A(\main.demo.zic._q_qpos[12] ),
    .B(_0640_),
    .Y(_0641_));
 sg13g2_a21oi_1 _1595_ (.A1(\main.demo.zic._q_qpos[12] ),
    .A2(_0001_),
    .Y(_0642_),
    .B1(_0641_));
 sg13g2_nand2_1 _1596_ (.Y(_0643_),
    .A(\main.demo.zic._d_clock_count[0] ),
    .B(_0642_));
 sg13g2_or3_1 _1597_ (.A(\main.demo.zic._q_clock_count[0] ),
    .B(\main.demo.zic._d_clock_count[0] ),
    .C(_0642_),
    .X(_0644_));
 sg13g2_nand3_1 _1598_ (.B(_0643_),
    .C(_0644_),
    .A(_0639_),
    .Y(_0645_));
 sg13g2_nand2_1 _1599_ (.Y(_0646_),
    .A(_0007_),
    .B(_0008_));
 sg13g2_nor4_1 _1600_ (.A(\main.demo.zic._q_clock_count[2] ),
    .B(\main.demo.zic._q_clock_count[4] ),
    .C(_0634_),
    .D(_0646_),
    .Y(_0647_));
 sg13g2_a21oi_1 _1601_ (.A1(_0006_),
    .A2(_0634_),
    .Y(_0648_),
    .B1(_0647_));
 sg13g2_a21oi_1 _1602_ (.A1(\main.demo.zic._q_clock_count[1] ),
    .A2(_0638_),
    .Y(_0649_),
    .B1(_0648_));
 sg13g2_a22oi_1 _1603_ (.Y(_0650_),
    .B1(_0645_),
    .B2(_0649_),
    .A2(_0636_),
    .A1(_0006_));
 sg13g2_inv_1 _1604_ (.Y(\main._w_demo_audio1 ),
    .A(_0650_));
 sg13g2_nand2b_1 _1605_ (.Y(_0651_),
    .B(\main.demo._q_u[4] ),
    .A_N(\main.demo._q_vT[8] ));
 sg13g2_xnor2_1 _1606_ (.Y(_0652_),
    .A(\main.demo._q_vT[8] ),
    .B(\main.demo._q_u[4] ));
 sg13g2_inv_1 _1607_ (.Y(_0653_),
    .A(_0652_));
 sg13g2_nor2b_1 _1608_ (.A(\main.demo._q_vT[7] ),
    .B_N(\main.demo._q_u[3] ),
    .Y(_0654_));
 sg13g2_nand2b_1 _1609_ (.Y(_0655_),
    .B(\main.demo._q_u[3] ),
    .A_N(\main.demo._q_vT[7] ));
 sg13g2_xor2_1 _1610_ (.B(\main.demo._q_u[3] ),
    .A(\main.demo._q_vT[7] ),
    .X(_0656_));
 sg13g2_nor2b_1 _1611_ (.A(\main.demo._q_vT[5] ),
    .B_N(\main.demo._q_u[1] ),
    .Y(_0657_));
 sg13g2_nand2b_1 _1612_ (.Y(_0658_),
    .B(\main.demo._q_vT[4] ),
    .A_N(\main.demo._q_u[0] ));
 sg13g2_nor2_1 _1613_ (.A(_0591_),
    .B(\main.demo._q_u[2] ),
    .Y(_0659_));
 sg13g2_nand2b_1 _1614_ (.Y(_0660_),
    .B(\main.demo._q_vT[5] ),
    .A_N(\main.demo._q_u[1] ));
 sg13g2_a221oi_1 _1615_ (.B2(_0660_),
    .C1(_0657_),
    .B1(_0658_),
    .A1(_0591_),
    .Y(_0661_),
    .A2(\main.demo._q_u[2] ));
 sg13g2_nor3_1 _1616_ (.A(_0656_),
    .B(_0659_),
    .C(_0661_),
    .Y(_0662_));
 sg13g2_or3_1 _1617_ (.A(_0656_),
    .B(_0659_),
    .C(_0661_),
    .X(_0663_));
 sg13g2_a21oi_2 _1618_ (.B1(_0653_),
    .Y(_0664_),
    .A2(_0663_),
    .A1(_0655_));
 sg13g2_o21ai_1 _1619_ (.B1(_0652_),
    .Y(_0665_),
    .A1(_0654_),
    .A2(_0662_));
 sg13g2_nor2b_1 _1620_ (.A(\main.demo._q_vT[9] ),
    .B_N(\main.demo._q_u[5] ),
    .Y(_0666_));
 sg13g2_xor2_1 _1621_ (.B(\main.demo._q_u[5] ),
    .A(\main.demo._q_vT[9] ),
    .X(_0667_));
 sg13g2_a21oi_1 _1622_ (.A1(_0651_),
    .A2(_0665_),
    .Y(_0668_),
    .B1(_0667_));
 sg13g2_a21o_1 _1623_ (.A2(_0665_),
    .A1(_0651_),
    .B1(_0667_),
    .X(_0669_));
 sg13g2_nand3_1 _1624_ (.B(_0665_),
    .C(_0667_),
    .A(_0651_),
    .Y(_0670_));
 sg13g2_nand3_1 _1625_ (.B(_0669_),
    .C(_0670_),
    .A(net400),
    .Y(_0671_));
 sg13g2_nor3_2 _1626_ (.A(_0652_),
    .B(_0654_),
    .C(_0662_),
    .Y(_0672_));
 sg13g2_nor3_1 _1627_ (.A(net344),
    .B(_0664_),
    .C(_0672_),
    .Y(_0673_));
 sg13g2_o21ai_1 _1628_ (.B1(_0656_),
    .Y(_0674_),
    .A1(_0659_),
    .A2(_0661_));
 sg13g2_and2_1 _1629_ (.A(_0663_),
    .B(_0674_),
    .X(_0675_));
 sg13g2_and2_1 _1630_ (.A(net281),
    .B(_0675_),
    .X(_0676_));
 sg13g2_o21ai_1 _1631_ (.B1(net344),
    .Y(_0677_),
    .A1(_0664_),
    .A2(_0672_));
 sg13g2_nor2b_1 _1632_ (.A(_0673_),
    .B_N(_0677_),
    .Y(_0678_));
 sg13g2_a21oi_1 _1633_ (.A1(_0676_),
    .A2(_0677_),
    .Y(_0679_),
    .B1(_0673_));
 sg13g2_a21oi_1 _1634_ (.A1(_0669_),
    .A2(_0670_),
    .Y(_0680_),
    .B1(\main.demo._q_frame[5] ));
 sg13g2_a21o_1 _1635_ (.A2(_0670_),
    .A1(_0669_),
    .B1(\main.demo._q_frame[5] ),
    .X(_0681_));
 sg13g2_nand2_1 _1636_ (.Y(_0682_),
    .A(_0671_),
    .B(_0681_));
 sg13g2_o21ai_1 _1637_ (.B1(_0671_),
    .Y(_0683_),
    .A1(_0679_),
    .A2(_0680_));
 sg13g2_xnor2_1 _1638_ (.Y(_0684_),
    .A(\main.demo._q_vT[10] ),
    .B(\main.demo._q_u[6] ));
 sg13g2_o21ai_1 _1639_ (.B1(_0684_),
    .Y(_0685_),
    .A1(_0666_),
    .A2(_0668_));
 sg13g2_or3_1 _1640_ (.A(_0666_),
    .B(_0668_),
    .C(_0684_),
    .X(_0686_));
 sg13g2_a21oi_1 _1641_ (.A1(_0685_),
    .A2(_0686_),
    .Y(_0687_),
    .B1(_0611_));
 sg13g2_and3_1 _1642_ (.X(_0688_),
    .A(_0611_),
    .B(_0685_),
    .C(_0686_));
 sg13g2_or2_1 _1643_ (.X(_0689_),
    .B(_0688_),
    .A(_0687_));
 sg13g2_o21ai_1 _1644_ (.B1(_0683_),
    .Y(_0690_),
    .A1(_0687_),
    .A2(_0688_));
 sg13g2_xnor2_1 _1645_ (.Y(_0691_),
    .A(_0683_),
    .B(_0689_));
 sg13g2_nand3_1 _1646_ (.B(_0685_),
    .C(_0686_),
    .A(_0612_),
    .Y(_0692_));
 sg13g2_o21ai_1 _1647_ (.B1(_0685_),
    .Y(_0693_),
    .A1(\main.demo._q_vT[10] ),
    .A2(_0613_));
 sg13g2_xnor2_1 _1648_ (.Y(_0694_),
    .A(\main.demo._q_frame[7] ),
    .B(\main.demo._q_u[7] ));
 sg13g2_xnor2_1 _1649_ (.Y(_0695_),
    .A(\main.demo._q_vT[11] ),
    .B(_0694_));
 sg13g2_xnor2_1 _1650_ (.Y(_0696_),
    .A(_0693_),
    .B(_0695_));
 sg13g2_a21oi_1 _1651_ (.A1(_0690_),
    .A2(_0692_),
    .Y(_0697_),
    .B1(_0696_));
 sg13g2_and3_1 _1652_ (.X(_0698_),
    .A(_0690_),
    .B(_0692_),
    .C(_0696_));
 sg13g2_or2_1 _1653_ (.X(_0699_),
    .B(_0698_),
    .A(_0697_));
 sg13g2_nor2b_1 _1654_ (.A(_0691_),
    .B_N(_0699_),
    .Y(_0700_));
 sg13g2_nor2_1 _1655_ (.A(net281),
    .B(_0675_),
    .Y(_0701_));
 sg13g2_nor3_1 _1656_ (.A(_0676_),
    .B(net457),
    .C(_0701_),
    .Y(\main.demo._d_addr[0] ));
 sg13g2_xnor2_1 _1657_ (.Y(_0702_),
    .A(_0676_),
    .B(_0678_));
 sg13g2_nor2_1 _1658_ (.A(net457),
    .B(_0702_),
    .Y(\main.demo._d_addr[1] ));
 sg13g2_xnor2_1 _1659_ (.Y(_0703_),
    .A(_0679_),
    .B(_0682_));
 sg13g2_nor2_1 _1660_ (.A(net457),
    .B(_0703_),
    .Y(\main.demo._d_addr[2] ));
 sg13g2_nand2_1 _1661_ (.Y(_0704_),
    .A(\main.demo._q_v[3] ),
    .B(\main.demo._q_uT[7] ));
 sg13g2_xnor2_1 _1662_ (.Y(_0705_),
    .A(\main.demo._q_v[3] ),
    .B(\main.demo._q_uT[7] ));
 sg13g2_nor2_1 _1663_ (.A(\main.demo._q_v[1] ),
    .B(\main.demo._q_uT[5] ),
    .Y(_0706_));
 sg13g2_nand2_1 _1664_ (.Y(_0707_),
    .A(\main.demo._q_v[0] ),
    .B(\main.demo._q_uT[4] ));
 sg13g2_a22oi_1 _1665_ (.Y(_0708_),
    .B1(\main.demo._q_uT[6] ),
    .B2(\main.demo._q_v[2] ),
    .A2(\main.demo._q_uT[5] ),
    .A1(\main.demo._q_v[1] ));
 sg13g2_o21ai_1 _1666_ (.B1(_0708_),
    .Y(_0709_),
    .A1(_0706_),
    .A2(_0707_));
 sg13g2_o21ai_1 _1667_ (.B1(_0709_),
    .Y(_0710_),
    .A1(\main.demo._q_v[2] ),
    .A2(\main.demo._q_uT[6] ));
 sg13g2_xnor2_1 _1668_ (.Y(_0711_),
    .A(_0705_),
    .B(_0710_));
 sg13g2_or2_1 _1669_ (.X(_0712_),
    .B(_0711_),
    .A(_0691_));
 sg13g2_a21oi_1 _1670_ (.A1(_0691_),
    .A2(_0711_),
    .Y(_0713_),
    .B1(net457));
 sg13g2_and2_1 _1671_ (.A(_0712_),
    .B(_0713_),
    .X(\main.demo._d_addr[3] ));
 sg13g2_and2_1 _1672_ (.A(\main.demo._q_v[4] ),
    .B(\main.demo._q_uT[8] ),
    .X(_0714_));
 sg13g2_or2_1 _1673_ (.X(_0715_),
    .B(\main.demo._q_uT[8] ),
    .A(\main.demo._q_v[4] ));
 sg13g2_nand2b_1 _1674_ (.Y(_0716_),
    .B(_0715_),
    .A_N(_0714_));
 sg13g2_o21ai_1 _1675_ (.B1(_0704_),
    .Y(_0717_),
    .A1(_0705_),
    .A2(_0710_));
 sg13g2_xnor2_1 _1676_ (.Y(_0718_),
    .A(_0716_),
    .B(_0717_));
 sg13g2_nand2b_1 _1677_ (.Y(_0719_),
    .B(_0718_),
    .A_N(_0711_));
 sg13g2_xnor2_1 _1678_ (.Y(_0720_),
    .A(_0711_),
    .B(_0718_));
 sg13g2_o21ai_1 _1679_ (.B1(_0720_),
    .Y(_0721_),
    .A1(_0697_),
    .A2(_0698_));
 sg13g2_xnor2_1 _1680_ (.Y(_0722_),
    .A(_0699_),
    .B(_0720_));
 sg13g2_or2_1 _1681_ (.X(_0723_),
    .B(_0722_),
    .A(_0712_));
 sg13g2_a21oi_1 _1682_ (.A1(_0712_),
    .A2(_0722_),
    .Y(_0724_),
    .B1(net457));
 sg13g2_and2_1 _1683_ (.A(_0723_),
    .B(_0724_),
    .X(\main.demo._d_addr[4] ));
 sg13g2_nand2_1 _1684_ (.Y(_0725_),
    .A(\main.demo._q_v[5] ),
    .B(\main.demo._q_uT[9] ));
 sg13g2_xnor2_1 _1685_ (.Y(_0726_),
    .A(\main.demo._q_v[5] ),
    .B(\main.demo._q_uT[9] ));
 sg13g2_a21oi_2 _1686_ (.B1(_0714_),
    .Y(_0727_),
    .A2(_0717_),
    .A1(_0715_));
 sg13g2_xor2_1 _1687_ (.B(_0727_),
    .A(_0726_),
    .X(_0728_));
 sg13g2_xnor2_1 _1688_ (.Y(_0729_),
    .A(_0726_),
    .B(_0727_));
 sg13g2_nor2_1 _1689_ (.A(_0718_),
    .B(_0729_),
    .Y(_0730_));
 sg13g2_xnor2_1 _1690_ (.Y(_0731_),
    .A(_0718_),
    .B(_0728_));
 sg13g2_a21oi_2 _1691_ (.B1(_0731_),
    .Y(_0732_),
    .A2(_0721_),
    .A1(_0719_));
 sg13g2_and3_1 _1692_ (.X(_0733_),
    .A(_0719_),
    .B(_0721_),
    .C(_0731_));
 sg13g2_nor2_1 _1693_ (.A(_0732_),
    .B(_0733_),
    .Y(_0734_));
 sg13g2_nor4_2 _1694_ (.A(_0712_),
    .B(_0722_),
    .C(_0732_),
    .Y(_0735_),
    .D(_0733_));
 sg13g2_xor2_1 _1695_ (.B(_0734_),
    .A(_0723_),
    .X(_0736_));
 sg13g2_nor2_1 _1696_ (.A(net457),
    .B(_0736_),
    .Y(\main.demo._d_addr[5] ));
 sg13g2_nor2_1 _1697_ (.A(_0732_),
    .B(_0735_),
    .Y(_0737_));
 sg13g2_o21ai_1 _1698_ (.B1(_0725_),
    .Y(_0738_),
    .A1(_0726_),
    .A2(_0727_));
 sg13g2_and2_1 _1699_ (.A(\main.demo._q_v[6] ),
    .B(\main.demo._q_uT[10] ),
    .X(_0739_));
 sg13g2_xor2_1 _1700_ (.B(\main.demo._q_uT[10] ),
    .A(\main.demo._q_v[6] ),
    .X(_0740_));
 sg13g2_xnor2_1 _1701_ (.Y(_0741_),
    .A(_0738_),
    .B(_0740_));
 sg13g2_xnor2_1 _1702_ (.Y(_0742_),
    .A(_0730_),
    .B(_0741_));
 sg13g2_o21ai_1 _1703_ (.B1(_0742_),
    .Y(_0743_),
    .A1(_0732_),
    .A2(_0735_));
 sg13g2_xor2_1 _1704_ (.B(_0742_),
    .A(_0737_),
    .X(_0744_));
 sg13g2_nor2_1 _1705_ (.A(_0700_),
    .B(_0744_),
    .Y(\main.demo._d_addr[6] ));
 sg13g2_nor2_1 _1706_ (.A(_0728_),
    .B(_0741_),
    .Y(_0745_));
 sg13g2_nand3_1 _1707_ (.B(_0728_),
    .C(_0741_),
    .A(_0718_),
    .Y(_0746_));
 sg13g2_and2_1 _1708_ (.A(_0743_),
    .B(_0746_),
    .X(_0747_));
 sg13g2_a21oi_1 _1709_ (.A1(_0738_),
    .A2(_0740_),
    .Y(_0748_),
    .B1(_0739_));
 sg13g2_xor2_1 _1710_ (.B(\main.demo._q_uT[11] ),
    .A(\main.demo._q_v[7] ),
    .X(_0749_));
 sg13g2_xnor2_1 _1711_ (.Y(_0750_),
    .A(_0748_),
    .B(_0749_));
 sg13g2_nand3_1 _1712_ (.B(_0746_),
    .C(_0750_),
    .A(_0743_),
    .Y(_0751_));
 sg13g2_xnor2_1 _1713_ (.Y(_0752_),
    .A(_0745_),
    .B(_0750_));
 sg13g2_xnor2_1 _1714_ (.Y(_0753_),
    .A(_0747_),
    .B(_0752_));
 sg13g2_nor2_1 _1715_ (.A(net457),
    .B(_0753_),
    .Y(\main.demo._d_addr[7] ));
 sg13g2_nand2b_1 _1716_ (.Y(_0754_),
    .B(_0741_),
    .A_N(_0751_));
 sg13g2_o21ai_1 _1717_ (.B1(_0729_),
    .Y(_0755_),
    .A1(_0743_),
    .A2(_0750_));
 sg13g2_nand3b_1 _1718_ (.B(_0751_),
    .C(_0755_),
    .Y(_0756_),
    .A_N(_0741_));
 sg13g2_a21oi_1 _1719_ (.A1(_0754_),
    .A2(_0756_),
    .Y(\main.demo._d_addr[8] ),
    .B1(_0700_));
 sg13g2_nand2b_1 _1720_ (.Y(_0757_),
    .B(_0750_),
    .A_N(net457));
 sg13g2_a21oi_1 _1721_ (.A1(_0741_),
    .A2(_0747_),
    .Y(\main.demo._d_addr[9] ),
    .B1(_0757_));
 sg13g2_nor2b_1 _1722_ (.A(net164),
    .B_N(\main.demo._q_prev_vs ),
    .Y(_0758_));
 sg13g2_o21ai_1 _1723_ (.B1(net613),
    .Y(_0759_),
    .A1(\main.demo._q_frame[0] ),
    .A2(_0758_));
 sg13g2_a21oi_1 _1724_ (.A1(_0599_),
    .A2(_0758_),
    .Y(_0021_),
    .B1(_0759_));
 sg13g2_nor2b_2 _1725_ (.A(\main.demo._q_addr[9] ),
    .B_N(\main.demo._q_addr[8] ),
    .Y(_0760_));
 sg13g2_nand2b_2 _1726_ (.Y(_0761_),
    .B(\main.demo._q_addr[8] ),
    .A_N(\main.demo._q_addr[9] ));
 sg13g2_and2_1 _1727_ (.A(\main.demo._q_addr[5] ),
    .B(\main.demo._q_addr[4] ),
    .X(_0762_));
 sg13g2_nand2_1 _1728_ (.Y(_0763_),
    .A(net601),
    .B(net602));
 sg13g2_nor2b_1 _1729_ (.A(\main.demo._q_addr[6] ),
    .B_N(net599),
    .Y(_0764_));
 sg13g2_nand2b_1 _1730_ (.Y(_0765_),
    .B(net599),
    .A_N(net600));
 sg13g2_nor2_2 _1731_ (.A(net589),
    .B(net586),
    .Y(_0766_));
 sg13g2_nor2_1 _1732_ (.A(net607),
    .B(net608),
    .Y(_0767_));
 sg13g2_or2_1 _1733_ (.X(_0768_),
    .B(net608),
    .A(net606));
 sg13g2_nor2b_1 _1734_ (.A(net605),
    .B_N(\main.demo._q_addr[3] ),
    .Y(_0769_));
 sg13g2_nand2b_2 _1735_ (.Y(_0770_),
    .B(net603),
    .A_N(net604));
 sg13g2_nor2_1 _1736_ (.A(net585),
    .B(_0770_),
    .Y(_0771_));
 sg13g2_nor2b_2 _1737_ (.A(net603),
    .B_N(net605),
    .Y(_0772_));
 sg13g2_nand2b_1 _1738_ (.Y(_0773_),
    .B(net604),
    .A_N(net603));
 sg13g2_nor2b_1 _1739_ (.A(\main.demo._q_addr[0] ),
    .B_N(net607),
    .Y(_0774_));
 sg13g2_nand2b_1 _1740_ (.Y(_0775_),
    .B(net606),
    .A_N(net608));
 sg13g2_nor2_1 _1741_ (.A(net581),
    .B(net578),
    .Y(_0776_));
 sg13g2_nand2b_2 _1742_ (.Y(_0777_),
    .B(net601),
    .A_N(net602));
 sg13g2_nand3b_1 _1743_ (.B(net600),
    .C(\main.demo._q_addr[5] ),
    .Y(_0778_),
    .A_N(\main.demo._q_addr[4] ));
 sg13g2_nor2_1 _1744_ (.A(_0607_),
    .B(_0778_),
    .Y(_0779_));
 sg13g2_a22oi_1 _1745_ (.Y(_0780_),
    .B1(net555),
    .B2(net553),
    .A2(net556),
    .A1(net559));
 sg13g2_nor2_1 _1746_ (.A(net585),
    .B(net583),
    .Y(_0781_));
 sg13g2_nor2_1 _1747_ (.A(net588),
    .B(_0777_),
    .Y(_0782_));
 sg13g2_nor2_1 _1748_ (.A(net604),
    .B(net603),
    .Y(_0783_));
 sg13g2_or2_2 _1749_ (.X(_0784_),
    .B(net603),
    .A(net604));
 sg13g2_nor2b_1 _1750_ (.A(net606),
    .B_N(\main.demo._q_addr[0] ),
    .Y(_0785_));
 sg13g2_nand2b_1 _1751_ (.Y(_0786_),
    .B(net608),
    .A_N(net606));
 sg13g2_nor2_2 _1752_ (.A(net607),
    .B(_0784_),
    .Y(_0787_));
 sg13g2_nor2_1 _1753_ (.A(_0784_),
    .B(net575),
    .Y(_0788_));
 sg13g2_nand3_1 _1754_ (.B(net602),
    .C(net600),
    .A(net601),
    .Y(_0789_));
 sg13g2_nor2_1 _1755_ (.A(_0607_),
    .B(_0789_),
    .Y(_0790_));
 sg13g2_or2_1 _1756_ (.X(_0791_),
    .B(_0789_),
    .A(_0607_));
 sg13g2_a22oi_1 _1757_ (.Y(_0792_),
    .B1(net542),
    .B2(net538),
    .A2(net543),
    .A1(net547));
 sg13g2_or2_2 _1758_ (.X(_0793_),
    .B(net599),
    .A(net600));
 sg13g2_nor2_1 _1759_ (.A(net601),
    .B(net602),
    .Y(_0794_));
 sg13g2_or2_1 _1760_ (.X(_0795_),
    .B(net602),
    .A(net601));
 sg13g2_nor2_2 _1761_ (.A(_0793_),
    .B(net573),
    .Y(_0796_));
 sg13g2_or4_2 _1762_ (.A(net601),
    .B(net602),
    .C(net600),
    .D(net599),
    .X(_0797_));
 sg13g2_and2_1 _1763_ (.A(net606),
    .B(\main.demo._q_addr[0] ),
    .X(_0798_));
 sg13g2_nand2_2 _1764_ (.Y(_0799_),
    .A(net607),
    .B(net608));
 sg13g2_nand2_1 _1765_ (.Y(_0800_),
    .A(net604),
    .B(net603));
 sg13g2_nor2_2 _1766_ (.A(_0799_),
    .B(net571),
    .Y(_0801_));
 sg13g2_nand4_1 _1767_ (.B(net608),
    .C(net604),
    .A(net606),
    .Y(_0802_),
    .D(net603));
 sg13g2_nor2_1 _1768_ (.A(_0797_),
    .B(_0802_),
    .Y(_0803_));
 sg13g2_nand3_1 _1769_ (.B(net608),
    .C(net603),
    .A(net606),
    .Y(_0804_));
 sg13g2_nor2_2 _1770_ (.A(net605),
    .B(_0804_),
    .Y(_0805_));
 sg13g2_nor4_2 _1771_ (.A(net605),
    .B(net590),
    .C(net588),
    .Y(_0806_),
    .D(_0804_));
 sg13g2_nor4_2 _1772_ (.A(net588),
    .B(net583),
    .C(net579),
    .Y(_0807_),
    .D(_0777_));
 sg13g2_nor2_1 _1773_ (.A(net586),
    .B(net573),
    .Y(_0808_));
 sg13g2_nor2_1 _1774_ (.A(net585),
    .B(net571),
    .Y(_0809_));
 sg13g2_nor4_1 _1775_ (.A(net588),
    .B(net585),
    .C(net573),
    .D(net571),
    .Y(_0810_));
 sg13g2_nor2_1 _1776_ (.A(_0807_),
    .B(_0810_),
    .Y(_0811_));
 sg13g2_nand2b_2 _1777_ (.Y(_0812_),
    .B(net602),
    .A_N(net601));
 sg13g2_nor2_2 _1778_ (.A(net574),
    .B(_0812_),
    .Y(_0813_));
 sg13g2_nor3_2 _1779_ (.A(net590),
    .B(net587),
    .C(_0802_),
    .Y(_0814_));
 sg13g2_a221oi_1 _1780_ (.B2(net556),
    .C1(_0814_),
    .B1(net520),
    .A1(net543),
    .Y(_0815_),
    .A2(net542));
 sg13g2_nor4_1 _1781_ (.A(_0803_),
    .B(_0806_),
    .C(_0807_),
    .D(_0810_),
    .Y(_0816_));
 sg13g2_nand4_1 _1782_ (.B(_0792_),
    .C(_0815_),
    .A(_0780_),
    .Y(_0817_),
    .D(_0816_));
 sg13g2_nor3_2 _1783_ (.A(_0606_),
    .B(_0607_),
    .C(net573),
    .Y(_0818_));
 sg13g2_nand3_1 _1784_ (.B(net599),
    .C(_0794_),
    .A(\main.demo._q_addr[6] ),
    .Y(_0819_));
 sg13g2_nor2_1 _1785_ (.A(net576),
    .B(net571),
    .Y(_0820_));
 sg13g2_a22oi_1 _1786_ (.Y(_0821_),
    .B1(net518),
    .B2(net538),
    .A2(net519),
    .A1(net534));
 sg13g2_nor2_1 _1787_ (.A(net581),
    .B(_0799_),
    .Y(_0822_));
 sg13g2_nor2_2 _1788_ (.A(net578),
    .B(net571),
    .Y(_0823_));
 sg13g2_a22oi_1 _1789_ (.Y(_0824_),
    .B1(net513),
    .B2(net519),
    .A2(net515),
    .A1(net553));
 sg13g2_nor2_1 _1790_ (.A(net598),
    .B(_0789_),
    .Y(_0825_));
 sg13g2_a22oi_1 _1791_ (.Y(_0826_),
    .B1(net507),
    .B2(net547),
    .A2(net527),
    .A1(net532));
 sg13g2_nand3b_1 _1792_ (.B(net602),
    .C(net600),
    .Y(_0827_),
    .A_N(net601));
 sg13g2_nor2_2 _1793_ (.A(_0607_),
    .B(_0827_),
    .Y(_0828_));
 sg13g2_nor2_1 _1794_ (.A(_0770_),
    .B(net576),
    .Y(_0829_));
 sg13g2_nand2_1 _1795_ (.Y(_0830_),
    .A(net537),
    .B(net513));
 sg13g2_nor2_1 _1796_ (.A(net579),
    .B(_0784_),
    .Y(_0831_));
 sg13g2_a22oi_1 _1797_ (.Y(_0832_),
    .B1(net500),
    .B2(net545),
    .A2(net521),
    .A1(_0787_));
 sg13g2_nor2_1 _1798_ (.A(_0770_),
    .B(net578),
    .Y(_0833_));
 sg13g2_nor3_2 _1799_ (.A(net577),
    .B(_0797_),
    .C(net572),
    .Y(_0834_));
 sg13g2_nand2_1 _1800_ (.Y(_0835_),
    .A(net539),
    .B(net536));
 sg13g2_nor4_1 _1801_ (.A(net606),
    .B(net608),
    .C(net604),
    .D(\main.demo._q_addr[3] ),
    .Y(_0836_));
 sg13g2_nor4_2 _1802_ (.A(net589),
    .B(net586),
    .C(net581),
    .Y(_0837_),
    .D(_0799_));
 sg13g2_nor2_1 _1803_ (.A(net586),
    .B(_0812_),
    .Y(_0838_));
 sg13g2_nor4_2 _1804_ (.A(net586),
    .B(net575),
    .C(net572),
    .Y(_0839_),
    .D(_0812_));
 sg13g2_nor2_2 _1805_ (.A(_0837_),
    .B(_0839_),
    .Y(_0840_));
 sg13g2_nor2_1 _1806_ (.A(net581),
    .B(net576),
    .Y(_0841_));
 sg13g2_nor2_1 _1807_ (.A(_0784_),
    .B(_0799_),
    .Y(_0842_));
 sg13g2_nand3_1 _1808_ (.B(_0832_),
    .C(_0840_),
    .A(_0826_),
    .Y(_0843_));
 sg13g2_o21ai_1 _1809_ (.B1(net545),
    .Y(_0844_),
    .A1(net497),
    .A2(net489));
 sg13g2_nand3_1 _1810_ (.B(_0830_),
    .C(_0844_),
    .A(_0821_),
    .Y(_0845_));
 sg13g2_a21oi_1 _1811_ (.A1(net505),
    .A2(net503),
    .Y(_0846_),
    .B1(_0834_));
 sg13g2_o21ai_1 _1812_ (.B1(net544),
    .Y(_0847_),
    .A1(net568),
    .A2(net485));
 sg13g2_nand4_1 _1813_ (.B(_0835_),
    .C(_0846_),
    .A(_0824_),
    .Y(_0848_),
    .D(_0847_));
 sg13g2_o21ai_1 _1814_ (.B1(net568),
    .Y(_0849_),
    .A1(net538),
    .A2(net519));
 sg13g2_a22oi_1 _1815_ (.Y(_0850_),
    .B1(net568),
    .B2(net536),
    .A2(net514),
    .A1(net520));
 sg13g2_nand2_1 _1816_ (.Y(_0851_),
    .A(net556),
    .B(net505));
 sg13g2_nor4_1 _1817_ (.A(net581),
    .B(net578),
    .C(net574),
    .D(_0812_),
    .Y(_0852_));
 sg13g2_a221oi_1 _1818_ (.B2(net520),
    .C1(_0852_),
    .B1(net493),
    .A1(net543),
    .Y(_0853_),
    .A2(net514));
 sg13g2_nand4_1 _1819_ (.B(_0850_),
    .C(_0851_),
    .A(_0849_),
    .Y(_0854_),
    .D(_0853_));
 sg13g2_nor4_1 _1820_ (.A(_0843_),
    .B(_0845_),
    .C(_0848_),
    .D(_0854_),
    .Y(_0855_));
 sg13g2_nand2b_1 _1821_ (.Y(_0856_),
    .B(_0855_),
    .A_N(_0817_));
 sg13g2_nor2b_2 _1822_ (.A(\main.demo._q_addr[8] ),
    .B_N(\main.demo._q_addr[9] ),
    .Y(_0857_));
 sg13g2_nand2b_2 _1823_ (.Y(_0858_),
    .B(\main.demo._q_addr[9] ),
    .A_N(\main.demo._q_addr[8] ));
 sg13g2_o21ai_1 _1824_ (.B1(net510),
    .Y(_0859_),
    .A1(net530),
    .A2(net526));
 sg13g2_nor3_1 _1825_ (.A(_0606_),
    .B(net597),
    .C(net573),
    .Y(_0860_));
 sg13g2_nand3_1 _1826_ (.B(_0607_),
    .C(_0794_),
    .A(net600),
    .Y(_0861_));
 sg13g2_o21ai_1 _1827_ (.B1(net490),
    .Y(_0862_),
    .A1(net549),
    .A2(net485));
 sg13g2_o21ai_1 _1828_ (.B1(net522),
    .Y(_0863_),
    .A1(net517),
    .A2(net495));
 sg13g2_nand2_1 _1829_ (.Y(_0864_),
    .A(_0862_),
    .B(_0863_));
 sg13g2_a22oi_1 _1830_ (.Y(_0865_),
    .B1(net479),
    .B2(net516),
    .A2(net495),
    .A1(net535));
 sg13g2_or4_1 _1831_ (.A(net588),
    .B(net584),
    .C(net575),
    .D(_0812_),
    .X(_0866_));
 sg13g2_nor2_1 _1832_ (.A(_0777_),
    .B(net574),
    .Y(_0867_));
 sg13g2_nand2_1 _1833_ (.Y(_0868_),
    .A(net539),
    .B(net475));
 sg13g2_a22oi_1 _1834_ (.Y(_0869_),
    .B1(net502),
    .B2(net535),
    .A2(net513),
    .A1(net523));
 sg13g2_a22oi_1 _1835_ (.Y(_0870_),
    .B1(net479),
    .B2(net530),
    .A2(net487),
    .A1(net490));
 sg13g2_o21ai_1 _1836_ (.B1(net523),
    .Y(_0871_),
    .A1(net554),
    .A2(net502));
 sg13g2_a22oi_1 _1837_ (.Y(_0872_),
    .B1(net477),
    .B2(net540),
    .A2(net479),
    .A1(net525));
 sg13g2_a22oi_1 _1838_ (.Y(_0873_),
    .B1(net479),
    .B2(net496),
    .A2(net490),
    .A1(net499));
 sg13g2_nand4_1 _1839_ (.B(_0870_),
    .C(_0872_),
    .A(_0865_),
    .Y(_0874_),
    .D(_0873_));
 sg13g2_nand3_1 _1840_ (.B(_0869_),
    .C(_0871_),
    .A(_0859_),
    .Y(_0875_));
 sg13g2_or3_1 _1841_ (.A(_0864_),
    .B(_0874_),
    .C(_0875_),
    .X(_0876_));
 sg13g2_nor2_2 _1842_ (.A(\main.demo._q_addr[9] ),
    .B(\main.demo._q_addr[8] ),
    .Y(_0877_));
 sg13g2_or2_2 _1843_ (.X(_0878_),
    .B(\main.demo._q_addr[8] ),
    .A(\main.demo._q_addr[9] ));
 sg13g2_and4_1 _1844_ (.A(\main.demo._q_addr[1] ),
    .B(_0772_),
    .C(net537),
    .D(_0877_),
    .X(_0879_));
 sg13g2_a221oi_1 _1845_ (.B2(_0876_),
    .C1(_0879_),
    .B1(_0857_),
    .A1(_0760_),
    .Y(_0880_),
    .A2(_0856_));
 sg13g2_a22oi_1 _1846_ (.Y(_0881_),
    .B1(net488),
    .B2(net522),
    .A2(net491),
    .A1(net554));
 sg13g2_nand2_1 _1847_ (.Y(_0882_),
    .A(net554),
    .B(net535));
 sg13g2_nand2_1 _1848_ (.Y(_0883_),
    .A(net533),
    .B(net522));
 sg13g2_nand3_1 _1849_ (.B(_0882_),
    .C(_0883_),
    .A(_0881_),
    .Y(_0884_));
 sg13g2_a22oi_1 _1850_ (.Y(_0885_),
    .B1(net475),
    .B2(net513),
    .A2(net491),
    .A1(net540));
 sg13g2_o21ai_1 _1851_ (.B1(net477),
    .Y(_0886_),
    .A1(net554),
    .A2(net498));
 sg13g2_o21ai_1 _1852_ (.B1(_0885_),
    .Y(_0887_),
    .A1(net605),
    .A2(_0886_));
 sg13g2_nand2_1 _1853_ (.Y(_0888_),
    .A(net502),
    .B(net480));
 sg13g2_a22oi_1 _1854_ (.Y(_0889_),
    .B1(net522),
    .B2(net557),
    .A2(_0796_),
    .A1(net540));
 sg13g2_nand2_1 _1855_ (.Y(_0890_),
    .A(_0888_),
    .B(_0889_));
 sg13g2_nor2_1 _1856_ (.A(net589),
    .B(net574),
    .Y(_0891_));
 sg13g2_nor4_2 _1857_ (.A(net590),
    .B(_0770_),
    .C(net577),
    .Y(_0892_),
    .D(_0793_));
 sg13g2_a21o_1 _1858_ (.A2(net481),
    .A1(_0823_),
    .B1(_0892_),
    .X(_0893_));
 sg13g2_or4_1 _1859_ (.A(_0884_),
    .B(_0887_),
    .C(_0890_),
    .D(_0893_),
    .X(_0894_));
 sg13g2_nor2_1 _1860_ (.A(net597),
    .B(_0827_),
    .Y(_0895_));
 sg13g2_a22oi_1 _1861_ (.Y(_0896_),
    .B1(net468),
    .B2(net525),
    .A2(net519),
    .A1(net541));
 sg13g2_a22oi_1 _1862_ (.Y(_0897_),
    .B1(net498),
    .B2(net537),
    .A2(net516),
    .A1(_0766_));
 sg13g2_nand2_1 _1863_ (.Y(_0898_),
    .A(net551),
    .B(net488));
 sg13g2_o21ai_1 _1864_ (.B1(net520),
    .Y(_0899_),
    .A1(net547),
    .A2(net483));
 sg13g2_o21ai_1 _1865_ (.B1(net527),
    .Y(_0900_),
    .A1(net547),
    .A2(net483));
 sg13g2_nand2_1 _1866_ (.Y(_0901_),
    .A(net514),
    .B(net505));
 sg13g2_a22oi_1 _1867_ (.Y(_0902_),
    .B1(net568),
    .B2(net505),
    .A2(net494),
    .A1(net560));
 sg13g2_nor4_2 _1868_ (.A(net589),
    .B(net586),
    .C(net581),
    .Y(_0903_),
    .D(net578));
 sg13g2_a22oi_1 _1869_ (.Y(_0904_),
    .B1(net467),
    .B2(net532),
    .A2(net494),
    .A1(net527));
 sg13g2_and3_1 _1870_ (.X(_0905_),
    .A(_0899_),
    .B(_0900_),
    .C(_0904_));
 sg13g2_a22oi_1 _1871_ (.Y(_0906_),
    .B1(net487),
    .B2(net551),
    .A2(net516),
    .A1(net529));
 sg13g2_and4_2 _1872_ (.A(_0862_),
    .B(_0896_),
    .C(_0897_),
    .D(_0906_),
    .X(_0907_));
 sg13g2_a21oi_1 _1873_ (.A1(net514),
    .A2(net504),
    .Y(_0908_),
    .B1(_0903_));
 sg13g2_nand4_1 _1874_ (.B(_0905_),
    .C(_0907_),
    .A(_0902_),
    .Y(_0909_),
    .D(_0908_));
 sg13g2_a22oi_1 _1875_ (.Y(_0910_),
    .B1(_0909_),
    .B2(_0760_),
    .A2(_0894_),
    .A1(_0857_));
 sg13g2_o21ai_1 _1876_ (.B1(net523),
    .Y(_0911_),
    .A1(net531),
    .A2(net526));
 sg13g2_a22oi_1 _1877_ (.Y(_0912_),
    .B1(net468),
    .B2(net533),
    .A2(net510),
    .A1(net557));
 sg13g2_nor2_1 _1878_ (.A(net598),
    .B(_0778_),
    .Y(_0913_));
 sg13g2_nor3_2 _1879_ (.A(net598),
    .B(_0789_),
    .C(_0802_),
    .Y(_0914_));
 sg13g2_a21oi_1 _1880_ (.A1(net557),
    .A2(net464),
    .Y(_0915_),
    .B1(_0914_));
 sg13g2_and3_1 _1881_ (.X(_0916_),
    .A(_0911_),
    .B(_0912_),
    .C(_0915_));
 sg13g2_a22oi_1 _1882_ (.Y(_0917_),
    .B1(net498),
    .B2(net465),
    .A2(net502),
    .A1(net544));
 sg13g2_nand2_1 _1883_ (.Y(_0918_),
    .A(net514),
    .B(net507));
 sg13g2_o21ai_1 _1884_ (.B1(net508),
    .Y(_0919_),
    .A1(net514),
    .A2(net501));
 sg13g2_nor4_2 _1885_ (.A(net597),
    .B(net580),
    .C(_0778_),
    .Y(_0920_),
    .D(net572));
 sg13g2_nor4_2 _1886_ (.A(net597),
    .B(_0770_),
    .C(net575),
    .Y(_0921_),
    .D(_0827_));
 sg13g2_nor2_2 _1887_ (.A(_0920_),
    .B(_0921_),
    .Y(_0922_));
 sg13g2_a22oi_1 _1888_ (.Y(_0923_),
    .B1(net511),
    .B2(net467),
    .A2(net532),
    .A1(net543));
 sg13g2_a22oi_1 _1889_ (.Y(_0924_),
    .B1(net474),
    .B2(net556),
    .A2(net501),
    .A1(net559));
 sg13g2_nand2_1 _1890_ (.Y(_0925_),
    .A(net487),
    .B(net468));
 sg13g2_a22oi_1 _1891_ (.Y(_0926_),
    .B1(net492),
    .B2(net524),
    .A2(net568),
    .A1(net509));
 sg13g2_nor4_2 _1892_ (.A(net586),
    .B(net578),
    .C(net572),
    .Y(_0927_),
    .D(_0812_));
 sg13g2_a21oi_1 _1893_ (.A1(net534),
    .A2(net474),
    .Y(_0928_),
    .B1(_0927_));
 sg13g2_nand4_1 _1894_ (.B(_0919_),
    .C(_0922_),
    .A(_0917_),
    .Y(_0929_),
    .D(_0926_));
 sg13g2_a22oi_1 _1895_ (.Y(_0930_),
    .B1(net486),
    .B2(net466),
    .A2(net511),
    .A1(net559));
 sg13g2_nand4_1 _1896_ (.B(_0924_),
    .C(_0928_),
    .A(_0923_),
    .Y(_0931_),
    .D(_0930_));
 sg13g2_o21ai_1 _1897_ (.B1(_0760_),
    .Y(_0932_),
    .A1(_0929_),
    .A2(_0931_));
 sg13g2_o21ai_1 _1898_ (.B1(_0932_),
    .Y(_0933_),
    .A1(_0858_),
    .A2(_0916_));
 sg13g2_inv_1 _1899_ (.Y(_0934_),
    .A(_0933_));
 sg13g2_o21ai_1 _1900_ (.B1(net510),
    .Y(_0935_),
    .A1(net555),
    .A2(net540));
 sg13g2_nor2_2 _1901_ (.A(_0761_),
    .B(_0935_),
    .Y(_0936_));
 sg13g2_o21ai_1 _1902_ (.B1(_0802_),
    .Y(_0937_),
    .A1(_0768_),
    .A2(_0770_));
 sg13g2_nor3_1 _1903_ (.A(net598),
    .B(_0778_),
    .C(_0802_),
    .Y(_0938_));
 sg13g2_a221oi_1 _1904_ (.B2(_0937_),
    .C1(_0938_),
    .B1(net466),
    .A1(net556),
    .Y(_0939_),
    .A2(net509));
 sg13g2_a21oi_2 _1905_ (.B1(_0761_),
    .Y(_0940_),
    .A2(_0939_),
    .A1(_0935_));
 sg13g2_nor3_2 _1906_ (.A(net580),
    .B(_0797_),
    .C(net572),
    .Y(_0941_));
 sg13g2_a221oi_1 _1907_ (.B2(net502),
    .C1(_0941_),
    .B1(net522),
    .A1(net560),
    .Y(_0942_),
    .A2(net526));
 sg13g2_nor2_2 _1908_ (.A(net591),
    .B(_0942_),
    .Y(_0943_));
 sg13g2_nor2_1 _1909_ (.A(_0940_),
    .B(_0943_),
    .Y(_0944_));
 sg13g2_nand4_1 _1910_ (.B(_0910_),
    .C(_0934_),
    .A(_0880_),
    .Y(_0945_),
    .D(_0944_));
 sg13g2_inv_1 _1911_ (.Y(_0946_),
    .A(_0945_));
 sg13g2_a22oi_1 _1912_ (.Y(_0947_),
    .B1(net469),
    .B2(net541),
    .A2(net525),
    .A1(net536));
 sg13g2_nor4_1 _1913_ (.A(net585),
    .B(_0777_),
    .C(_0784_),
    .D(net574),
    .Y(_0948_));
 sg13g2_nand2_1 _1914_ (.Y(_0949_),
    .A(net517),
    .B(net476));
 sg13g2_o21ai_1 _1915_ (.B1(net477),
    .Y(_0950_),
    .A1(net518),
    .A2(net568));
 sg13g2_nor4_2 _1916_ (.A(_0606_),
    .B(net597),
    .C(net573),
    .Y(_0951_),
    .D(_0802_));
 sg13g2_nor4_2 _1917_ (.A(net590),
    .B(_0770_),
    .C(net578),
    .Y(_0952_),
    .D(_0793_));
 sg13g2_nor4_2 _1918_ (.A(net588),
    .B(net585),
    .C(_0784_),
    .Y(_0953_),
    .D(_0795_));
 sg13g2_nand3_1 _1919_ (.B(_0794_),
    .C(net569),
    .A(_0764_),
    .Y(_0954_));
 sg13g2_nor4_2 _1920_ (.A(net598),
    .B(net580),
    .C(_0789_),
    .Y(_0955_),
    .D(net572));
 sg13g2_nor4_2 _1921_ (.A(_0951_),
    .B(_0952_),
    .C(_0953_),
    .Y(_0956_),
    .D(_0955_));
 sg13g2_a22oi_1 _1922_ (.Y(_0957_),
    .B1(_0772_),
    .B2(_0798_),
    .A2(_0769_),
    .A1(_0767_));
 sg13g2_nand2b_1 _1923_ (.Y(_0958_),
    .B(net481),
    .A_N(_0957_));
 sg13g2_and2_1 _1924_ (.A(net555),
    .B(net481),
    .X(_0959_));
 sg13g2_a22oi_1 _1925_ (.Y(_0960_),
    .B1(net465),
    .B2(net568),
    .A2(net478),
    .A1(net555));
 sg13g2_nand2_1 _1926_ (.Y(_0961_),
    .A(_0958_),
    .B(_0960_));
 sg13g2_nand3_1 _1927_ (.B(_0958_),
    .C(_0960_),
    .A(_0956_),
    .Y(_0962_));
 sg13g2_nand2b_1 _1928_ (.Y(_0963_),
    .B(net536),
    .A_N(_0957_));
 sg13g2_nor4_2 _1929_ (.A(net597),
    .B(net582),
    .C(_0778_),
    .Y(_0964_),
    .D(_0799_));
 sg13g2_nand4_1 _1930_ (.B(_0919_),
    .C(_0947_),
    .A(_0850_),
    .Y(_0965_),
    .D(_0963_));
 sg13g2_a21oi_1 _1931_ (.A1(net512),
    .A2(net466),
    .Y(_0966_),
    .B1(_0964_));
 sg13g2_a22oi_1 _1932_ (.Y(_0967_),
    .B1(net568),
    .B2(net467),
    .A2(net508),
    .A1(net518));
 sg13g2_a22oi_1 _1933_ (.Y(_0968_),
    .B1(net465),
    .B2(net503),
    .A2(net493),
    .A1(net508));
 sg13g2_nand4_1 _1934_ (.B(_0966_),
    .C(_0967_),
    .A(_0950_),
    .Y(_0969_),
    .D(_0968_));
 sg13g2_or3_1 _1935_ (.A(_0962_),
    .B(_0965_),
    .C(_0969_),
    .X(_0970_));
 sg13g2_nand2_1 _1936_ (.Y(_0971_),
    .A(net556),
    .B(net543));
 sg13g2_o21ai_1 _1937_ (.B1(net545),
    .Y(_0972_),
    .A1(net556),
    .A2(net524));
 sg13g2_a22oi_1 _1938_ (.Y(_0973_),
    .B1(net486),
    .B2(net520),
    .A2(net500),
    .A1(net536));
 sg13g2_a22oi_1 _1939_ (.Y(_0974_),
    .B1(net500),
    .B2(net521),
    .A2(net511),
    .A1(net528));
 sg13g2_a22oi_1 _1940_ (.Y(_0975_),
    .B1(net492),
    .B2(net532),
    .A2(net503),
    .A1(net527));
 sg13g2_a22oi_1 _1941_ (.Y(_0976_),
    .B1(net482),
    .B2(net507),
    .A2(net492),
    .A1(net534));
 sg13g2_o21ai_1 _1942_ (.B1(_0972_),
    .Y(_0977_),
    .A1(_0791_),
    .A2(_0804_));
 sg13g2_nand4_1 _1943_ (.B(_0974_),
    .C(_0975_),
    .A(_0973_),
    .Y(_0978_),
    .D(_0976_));
 sg13g2_or2_1 _1944_ (.X(_0979_),
    .B(_0978_),
    .A(_0977_));
 sg13g2_nand2_1 _1945_ (.Y(_0980_),
    .A(net484),
    .B(net476));
 sg13g2_a22oi_1 _1946_ (.Y(_0981_),
    .B1(net484),
    .B2(net476),
    .A2(net496),
    .A1(net551));
 sg13g2_a22oi_1 _1947_ (.Y(_0982_),
    .B1(net488),
    .B2(net537),
    .A2(net506),
    .A1(net516));
 sg13g2_o21ai_1 _1948_ (.B1(net558),
    .Y(_0983_),
    .A1(net552),
    .A2(net472));
 sg13g2_a22oi_1 _1949_ (.Y(_0984_),
    .B1(net475),
    .B2(net548),
    .A2(net506),
    .A1(net513));
 sg13g2_a22oi_1 _1950_ (.Y(_0985_),
    .B1(net496),
    .B2(net551),
    .A2(net506),
    .A1(net516));
 sg13g2_a22oi_1 _1951_ (.Y(_0986_),
    .B1(net503),
    .B2(net551),
    .A2(net506),
    .A1(net533));
 sg13g2_and3_1 _1952_ (.X(_0987_),
    .A(_0983_),
    .B(_0984_),
    .C(_0985_));
 sg13g2_a21oi_1 _1953_ (.A1(net558),
    .A2(net538),
    .Y(_0988_),
    .B1(_0892_));
 sg13g2_o21ai_1 _1954_ (.B1(net537),
    .Y(_0989_),
    .A1(net533),
    .A2(net488));
 sg13g2_and4_1 _1955_ (.A(_0980_),
    .B(_0986_),
    .C(_0988_),
    .D(_0989_),
    .X(_0990_));
 sg13g2_a21oi_1 _1956_ (.A1(_0987_),
    .A2(_0990_),
    .Y(_0991_),
    .B1(_0878_));
 sg13g2_a221oi_1 _1957_ (.B2(_0760_),
    .C1(_0991_),
    .B1(_0979_),
    .A1(_0857_),
    .Y(_0992_),
    .A2(_0970_));
 sg13g2_nor4_2 _1958_ (.A(net597),
    .B(_0784_),
    .C(_0799_),
    .Y(_0993_),
    .D(_0827_));
 sg13g2_nor4_2 _1959_ (.A(net590),
    .B(net582),
    .C(net575),
    .Y(_0994_),
    .D(net574));
 sg13g2_nor4_2 _1960_ (.A(net589),
    .B(net581),
    .C(net578),
    .Y(_0995_),
    .D(net574));
 sg13g2_nor4_2 _1961_ (.A(net586),
    .B(_0777_),
    .C(net576),
    .Y(_0996_),
    .D(net571));
 sg13g2_nor4_2 _1962_ (.A(_0993_),
    .B(_0994_),
    .C(_0995_),
    .Y(_0997_),
    .D(_0996_));
 sg13g2_nor4_1 _1963_ (.A(net546),
    .B(net532),
    .C(net524),
    .D(net493),
    .Y(_0998_));
 sg13g2_nor2_1 _1964_ (.A(_0791_),
    .B(_0998_),
    .Y(_0999_));
 sg13g2_nor4_2 _1965_ (.A(net604),
    .B(net598),
    .C(_0778_),
    .Y(_1000_),
    .D(_0804_));
 sg13g2_nor4_2 _1966_ (.A(net597),
    .B(_0778_),
    .C(net575),
    .Y(_1001_),
    .D(net571));
 sg13g2_nor4_1 _1967_ (.A(net589),
    .B(net585),
    .C(net574),
    .D(net571),
    .Y(_1002_));
 sg13g2_nor4_2 _1968_ (.A(_0948_),
    .B(_1000_),
    .C(_1001_),
    .Y(_1003_),
    .D(_1002_));
 sg13g2_a22oi_1 _1969_ (.Y(_1004_),
    .B1(net471),
    .B2(net533),
    .A2(net480),
    .A1(net570));
 sg13g2_a22oi_1 _1970_ (.Y(_1005_),
    .B1(net496),
    .B2(net465),
    .A2(_0805_),
    .A1(net553));
 sg13g2_nand2_1 _1971_ (.Y(_1006_),
    .A(_1004_),
    .B(_1005_));
 sg13g2_a22oi_1 _1972_ (.Y(_1007_),
    .B1(net482),
    .B2(net527),
    .A2(net501),
    .A1(net560));
 sg13g2_nor4_1 _1973_ (.A(net589),
    .B(net587),
    .C(net585),
    .D(net581),
    .Y(_1008_));
 sg13g2_a22oi_1 _1974_ (.Y(_1009_),
    .B1(net473),
    .B2(net518),
    .A2(net483),
    .A1(net560));
 sg13g2_nand2b_1 _1975_ (.Y(_1010_),
    .B(net519),
    .A_N(_0957_));
 sg13g2_nor4_2 _1976_ (.A(_0837_),
    .B(_0839_),
    .C(_0903_),
    .Y(_1011_),
    .D(_0927_));
 sg13g2_a22oi_1 _1977_ (.Y(_1012_),
    .B1(net473),
    .B2(net512),
    .A2(net474),
    .A1(net514));
 sg13g2_a221oi_1 _1978_ (.B2(net511),
    .C1(_0964_),
    .B1(net473),
    .A1(net514),
    .Y(_1013_),
    .A2(net474));
 sg13g2_nand2b_1 _1979_ (.Y(_1014_),
    .B(_1012_),
    .A_N(_0964_));
 sg13g2_nor4_2 _1980_ (.A(net588),
    .B(net582),
    .C(_0799_),
    .Y(_1015_),
    .D(_0812_));
 sg13g2_a21o_1 _1981_ (.A2(net466),
    .A1(net546),
    .B1(_1015_),
    .X(_1016_));
 sg13g2_a22oi_1 _1982_ (.Y(_1017_),
    .B1(net506),
    .B2(net525),
    .A2(net519),
    .A1(net547));
 sg13g2_a22oi_1 _1983_ (.Y(_1018_),
    .B1(net569),
    .B2(_0766_),
    .A2(net539),
    .A1(net553));
 sg13g2_o21ai_1 _1984_ (.B1(net465),
    .Y(_1019_),
    .A1(net557),
    .A2(net502));
 sg13g2_nand2_1 _1985_ (.Y(_1020_),
    .A(_1003_),
    .B(_1011_));
 sg13g2_a22oi_1 _1986_ (.Y(_1021_),
    .B1(net478),
    .B2(net511),
    .A2(net492),
    .A1(net534));
 sg13g2_a22oi_1 _1987_ (.Y(_1022_),
    .B1(net466),
    .B2(net546),
    .A2(net482),
    .A1(net504));
 sg13g2_nand4_1 _1988_ (.B(_1007_),
    .C(_1021_),
    .A(_0902_),
    .Y(_1023_),
    .D(_1022_));
 sg13g2_nand4_1 _1989_ (.B(_0821_),
    .C(_1017_),
    .A(_0780_),
    .Y(_1024_),
    .D(_1018_));
 sg13g2_nand3_1 _1990_ (.B(_1010_),
    .C(_1019_),
    .A(_1009_),
    .Y(_1025_));
 sg13g2_nor3_1 _1991_ (.A(_1023_),
    .B(_1024_),
    .C(_1025_),
    .Y(_1026_));
 sg13g2_a221oi_1 _1992_ (.B2(net555),
    .C1(_1015_),
    .B1(net465),
    .A1(net559),
    .Y(_1027_),
    .A2(net546));
 sg13g2_nand4_1 _1993_ (.B(_0997_),
    .C(_1013_),
    .A(_0956_),
    .Y(_1028_),
    .D(_1027_));
 sg13g2_nor4_1 _1994_ (.A(_0999_),
    .B(_1006_),
    .C(_1020_),
    .D(_1028_),
    .Y(_1029_));
 sg13g2_a21o_1 _1995_ (.A2(_1029_),
    .A1(_1026_),
    .B1(_0878_),
    .X(_1030_));
 sg13g2_nand2_2 _1996_ (.Y(_1031_),
    .A(net535),
    .B(net484));
 sg13g2_o21ai_1 _1997_ (.B1(_0858_),
    .Y(_1032_),
    .A1(net591),
    .A2(_1031_));
 sg13g2_nor3_1 _1998_ (.A(_0768_),
    .B(net584),
    .C(_0797_),
    .Y(_1033_));
 sg13g2_nand2_1 _1999_ (.Y(_1034_),
    .A(net549),
    .B(net536));
 sg13g2_and4_1 _2000_ (.A(_0917_),
    .B(_0980_),
    .C(_1031_),
    .D(_1034_),
    .X(_1035_));
 sg13g2_o21ai_1 _2001_ (.B1(net545),
    .Y(_1036_),
    .A1(net530),
    .A2(net495));
 sg13g2_nand2_1 _2002_ (.Y(_1037_),
    .A(net500),
    .B(net473));
 sg13g2_o21ai_1 _2003_ (.B1(net471),
    .Y(_1038_),
    .A1(net499),
    .A2(net484));
 sg13g2_nand2_1 _2004_ (.Y(_1039_),
    .A(net487),
    .B(net464));
 sg13g2_nand4_1 _2005_ (.B(_1036_),
    .C(_1038_),
    .A(_1035_),
    .Y(_1040_),
    .D(_1039_));
 sg13g2_a22oi_1 _2006_ (.Y(_1041_),
    .B1(net471),
    .B2(net548),
    .A2(net530),
    .A1(net535));
 sg13g2_o21ai_1 _2007_ (.B1(net544),
    .Y(_1042_),
    .A1(net525),
    .A2(net513));
 sg13g2_nand2_1 _2008_ (.Y(_1043_),
    .A(_1041_),
    .B(_1042_));
 sg13g2_nand2_1 _2009_ (.Y(_1044_),
    .A(net548),
    .B(net479));
 sg13g2_a22oi_1 _2010_ (.Y(_1045_),
    .B1(net471),
    .B2(net541),
    .A2(net476),
    .A1(net533));
 sg13g2_a22oi_1 _2011_ (.Y(_1046_),
    .B1(net471),
    .B2(net558),
    .A2(net522),
    .A1(net549));
 sg13g2_nand4_1 _2012_ (.B(_1044_),
    .C(_1045_),
    .A(_0997_),
    .Y(_1047_),
    .D(_1046_));
 sg13g2_or2_1 _2013_ (.X(_1048_),
    .B(_1047_),
    .A(_1043_));
 sg13g2_o21ai_1 _2014_ (.B1(_1032_),
    .Y(_1049_),
    .A1(_1040_),
    .A2(_1048_));
 sg13g2_o21ai_1 _2015_ (.B1(_0818_),
    .Y(_1050_),
    .A1(net530),
    .A2(net525));
 sg13g2_a22oi_1 _2016_ (.Y(_1051_),
    .B1(net530),
    .B2(net471),
    .A2(net548),
    .A1(net552));
 sg13g2_nand2_1 _2017_ (.Y(_1052_),
    .A(_1050_),
    .B(_1051_));
 sg13g2_nand2_1 _2018_ (.Y(_1053_),
    .A(net557),
    .B(net490));
 sg13g2_a22oi_1 _2019_ (.Y(_1054_),
    .B1(net484),
    .B2(net480),
    .A2(_0801_),
    .A1(net544));
 sg13g2_nand3_1 _2020_ (.B(_1053_),
    .C(_1054_),
    .A(_1044_),
    .Y(_1055_));
 sg13g2_o21ai_1 _2021_ (.B1(net570),
    .Y(_1056_),
    .A1(net491),
    .A2(net471));
 sg13g2_a22oi_1 _2022_ (.Y(_1057_),
    .B1(net464),
    .B2(net526),
    .A2(net515),
    .A1(net529));
 sg13g2_a22oi_1 _2023_ (.Y(_1058_),
    .B1(net469),
    .B2(net517),
    .A2(net498),
    .A1(net510));
 sg13g2_a22oi_1 _2024_ (.Y(_1059_),
    .B1(net485),
    .B2(net537),
    .A2(net491),
    .A1(net496));
 sg13g2_a22oi_1 _2025_ (.Y(_1060_),
    .B1(net570),
    .B2(net469),
    .A2(net498),
    .A1(net506));
 sg13g2_nand3_1 _2026_ (.B(_1057_),
    .C(_1060_),
    .A(_1017_),
    .Y(_1061_));
 sg13g2_a22oi_1 _2027_ (.Y(_1062_),
    .B1(net493),
    .B2(net466),
    .A2(net504),
    .A1(net532));
 sg13g2_nor3_1 _2028_ (.A(_1014_),
    .B(_1052_),
    .C(_1055_),
    .Y(_1063_));
 sg13g2_a22oi_1 _2029_ (.Y(_1064_),
    .B1(net502),
    .B2(net479),
    .A2(net510),
    .A1(net530));
 sg13g2_nand4_1 _2030_ (.B(_1058_),
    .C(_1059_),
    .A(_1056_),
    .Y(_1065_),
    .D(_1064_));
 sg13g2_a22oi_1 _2031_ (.Y(_1066_),
    .B1(net478),
    .B2(net524),
    .A2(net486),
    .A1(net504));
 sg13g2_a22oi_1 _2032_ (.Y(_1067_),
    .B1(net483),
    .B2(net559),
    .A2(net524),
    .A1(net538));
 sg13g2_a21oi_1 _2033_ (.A1(net507),
    .A2(net486),
    .Y(_1068_),
    .B1(_0996_));
 sg13g2_nand4_1 _2034_ (.B(_1066_),
    .C(_1067_),
    .A(_1062_),
    .Y(_1069_),
    .D(_1068_));
 sg13g2_nor3_1 _2035_ (.A(_1061_),
    .B(_1065_),
    .C(_1069_),
    .Y(_1070_));
 sg13g2_a21o_1 _2036_ (.A2(_1070_),
    .A1(_1063_),
    .B1(net591),
    .X(_1071_));
 sg13g2_nand3_1 _2037_ (.B(_1049_),
    .C(_1071_),
    .A(_1030_),
    .Y(_1072_));
 sg13g2_and4_1 _2038_ (.A(_0992_),
    .B(_1030_),
    .C(_1049_),
    .D(_1071_),
    .X(_1073_));
 sg13g2_o21ai_1 _2039_ (.B1(net527),
    .Y(_1074_),
    .A1(net558),
    .A2(net518));
 sg13g2_nand4_1 _2040_ (.B(_0826_),
    .C(_0904_),
    .A(_0811_),
    .Y(_1075_),
    .D(_1074_));
 sg13g2_a22oi_1 _2041_ (.Y(_1076_),
    .B1(net464),
    .B2(net540),
    .A2(net510),
    .A1(net554));
 sg13g2_nand4_1 _2042_ (.B(_0917_),
    .C(_1058_),
    .A(_0896_),
    .Y(_1077_),
    .D(_1076_));
 sg13g2_nor2_1 _2043_ (.A(_1075_),
    .B(_1077_),
    .Y(_1078_));
 sg13g2_a22oi_1 _2044_ (.Y(_1079_),
    .B1(net494),
    .B2(net478),
    .A2(net501),
    .A1(net504));
 sg13g2_o21ai_1 _2045_ (.B1(net507),
    .Y(_1080_),
    .A1(net501),
    .A2(net494));
 sg13g2_nand2_1 _2046_ (.Y(_1081_),
    .A(_1079_),
    .B(_1080_));
 sg13g2_o21ai_1 _2047_ (.B1(net511),
    .Y(_1082_),
    .A1(net559),
    .A2(net527));
 sg13g2_nand3_1 _2048_ (.B(_1037_),
    .C(_1082_),
    .A(_0792_),
    .Y(_1083_));
 sg13g2_a22oi_1 _2049_ (.Y(_1084_),
    .B1(net477),
    .B2(_0809_),
    .A2(net492),
    .A1(net542));
 sg13g2_a22oi_1 _2050_ (.Y(_1085_),
    .B1(net504),
    .B2(net555),
    .A2(net520),
    .A1(net532));
 sg13g2_nand2_1 _2051_ (.Y(_1086_),
    .A(_1084_),
    .B(_1085_));
 sg13g2_o21ai_1 _2052_ (.B1(net507),
    .Y(_1087_),
    .A1(net486),
    .A2(net482));
 sg13g2_and2_1 _2053_ (.A(net487),
    .B(net479),
    .X(_1088_));
 sg13g2_a22oi_1 _2054_ (.Y(_1089_),
    .B1(net486),
    .B2(net478),
    .A2(net511),
    .A1(net553));
 sg13g2_nand2_1 _2055_ (.Y(_1090_),
    .A(_1087_),
    .B(_1089_));
 sg13g2_nor4_2 _2056_ (.A(_1081_),
    .B(_1083_),
    .C(_1086_),
    .Y(_1091_),
    .D(_1090_));
 sg13g2_a21oi_1 _2057_ (.A1(_1078_),
    .A2(_1091_),
    .Y(_1092_),
    .B1(_0878_));
 sg13g2_a22oi_1 _2058_ (.Y(_1093_),
    .B1(net570),
    .B2(net560),
    .A2(net515),
    .A1(net545));
 sg13g2_nor2_1 _2059_ (.A(_0858_),
    .B(_1093_),
    .Y(_1094_));
 sg13g2_a21oi_1 _2060_ (.A1(_0869_),
    .A2(_0882_),
    .Y(_1095_),
    .B1(net591));
 sg13g2_nor4_1 _2061_ (.A(_0933_),
    .B(_1092_),
    .C(_1094_),
    .D(_1095_),
    .Y(_1096_));
 sg13g2_nand2_1 _2062_ (.Y(_1097_),
    .A(net531),
    .B(net475));
 sg13g2_nand2_1 _2063_ (.Y(_1098_),
    .A(net534),
    .B(net528));
 sg13g2_a22oi_1 _2064_ (.Y(_1099_),
    .B1(net464),
    .B2(net548),
    .A2(net529),
    .A1(net533));
 sg13g2_and2_1 _2065_ (.A(_1097_),
    .B(_1099_),
    .X(_1100_));
 sg13g2_o21ai_1 _2066_ (.B1(_0828_),
    .Y(_1101_),
    .A1(net548),
    .A2(net495));
 sg13g2_o21ai_1 _2067_ (.B1(net499),
    .Y(_1102_),
    .A1(net519),
    .A2(net490));
 sg13g2_nand2_1 _2068_ (.Y(_1103_),
    .A(_1101_),
    .B(_1102_));
 sg13g2_a22oi_1 _2069_ (.Y(_1104_),
    .B1(net472),
    .B2(net515),
    .A2(net485),
    .A1(net551));
 sg13g2_a22oi_1 _2070_ (.Y(_1105_),
    .B1(net506),
    .B2(net541),
    .A2(net517),
    .A1(_0818_));
 sg13g2_nand2_1 _2071_ (.Y(_1106_),
    .A(_1104_),
    .B(_1105_));
 sg13g2_nor4_2 _2072_ (.A(net589),
    .B(net587),
    .C(net582),
    .Y(_1107_),
    .D(net575));
 sg13g2_nor4_2 _2073_ (.A(net587),
    .B(net584),
    .C(net575),
    .Y(_1108_),
    .D(net573));
 sg13g2_nor4_2 _2074_ (.A(net587),
    .B(net582),
    .C(net579),
    .Y(_1109_),
    .D(net573));
 sg13g2_nor4_2 _2075_ (.A(_1008_),
    .B(_1107_),
    .C(_1108_),
    .Y(_1110_),
    .D(_1109_));
 sg13g2_a22oi_1 _2076_ (.Y(_1111_),
    .B1(net513),
    .B2(net475),
    .A2(_0801_),
    .A1(net552));
 sg13g2_a22oi_1 _2077_ (.Y(_1112_),
    .B1(net476),
    .B2(net502),
    .A2(net484),
    .A1(net519));
 sg13g2_and4_1 _2078_ (.A(_1100_),
    .B(_1101_),
    .C(_1102_),
    .D(_1110_),
    .X(_1113_));
 sg13g2_a221oi_1 _2079_ (.B2(net493),
    .C1(_0993_),
    .B1(net509),
    .A1(net536),
    .Y(_1114_),
    .A2(net524));
 sg13g2_nand4_1 _2080_ (.B(_1084_),
    .C(_1085_),
    .A(_1003_),
    .Y(_1115_),
    .D(_1114_));
 sg13g2_a22oi_1 _2081_ (.Y(_1116_),
    .B1(net493),
    .B2(net478),
    .A2(net527),
    .A1(net558));
 sg13g2_a22oi_1 _2082_ (.Y(_1117_),
    .B1(net478),
    .B2(net532),
    .A2(net507),
    .A1(net524));
 sg13g2_a22oi_1 _2083_ (.Y(_1118_),
    .B1(net473),
    .B2(net518),
    .A2(net482),
    .A1(net504));
 sg13g2_a21oi_1 _2084_ (.A1(net546),
    .A2(net538),
    .Y(_1119_),
    .B1(_0951_));
 sg13g2_nand4_1 _2085_ (.B(_1117_),
    .C(_1118_),
    .A(_1116_),
    .Y(_1120_),
    .D(_1119_));
 sg13g2_nand3_1 _2086_ (.B(_1111_),
    .C(_1112_),
    .A(_0983_),
    .Y(_1121_));
 sg13g2_nor4_2 _2087_ (.A(_1106_),
    .B(_1115_),
    .C(_1120_),
    .Y(_1122_),
    .D(_1121_));
 sg13g2_a21oi_1 _2088_ (.A1(_1113_),
    .A2(_1122_),
    .Y(_1123_),
    .B1(net591));
 sg13g2_a21o_1 _2089_ (.A2(_1122_),
    .A1(_1113_),
    .B1(net591),
    .X(_1124_));
 sg13g2_and2_1 _2090_ (.A(net499),
    .B(net468),
    .X(_1125_));
 sg13g2_a221oi_1 _2091_ (.B2(net554),
    .C1(_1125_),
    .B1(net464),
    .A1(net540),
    .Y(_1126_),
    .A2(net529));
 sg13g2_a221oi_1 _2092_ (.B2(net526),
    .C1(_1088_),
    .B1(net475),
    .A1(net535),
    .Y(_1127_),
    .A2(net487));
 sg13g2_a22oi_1 _2093_ (.Y(_1128_),
    .B1(net468),
    .B2(net516),
    .A2(net484),
    .A1(net522));
 sg13g2_a22oi_1 _2094_ (.Y(_1129_),
    .B1(net471),
    .B2(net530),
    .A2(net490),
    .A1(net570));
 sg13g2_and3_1 _2095_ (.X(_1130_),
    .A(_1076_),
    .B(_1128_),
    .C(_1129_));
 sg13g2_a22oi_1 _2096_ (.Y(_1131_),
    .B1(net475),
    .B2(net548),
    .A2(net499),
    .A1(net535));
 sg13g2_a21oi_1 _2097_ (.A1(net495),
    .A2(net464),
    .Y(_1132_),
    .B1(_1015_));
 sg13g2_and4_1 _2098_ (.A(_1126_),
    .B(_1127_),
    .C(_1131_),
    .D(_1132_),
    .X(_1133_));
 sg13g2_a21oi_1 _2099_ (.A1(_1130_),
    .A2(_1133_),
    .Y(_1134_),
    .B1(_0858_));
 sg13g2_a21o_1 _2100_ (.A2(_1133_),
    .A1(_1130_),
    .B1(_0858_),
    .X(_1135_));
 sg13g2_nand2_1 _2101_ (.Y(_1136_),
    .A(net551),
    .B(net498));
 sg13g2_o21ai_1 _2102_ (.B1(_0818_),
    .Y(_1137_),
    .A1(net496),
    .A2(net488));
 sg13g2_a22oi_1 _2103_ (.Y(_1138_),
    .B1(_0785_),
    .B2(_0769_),
    .A2(_0774_),
    .A1(_0772_));
 sg13g2_and2_1 _2104_ (.A(net487),
    .B(net475),
    .X(_1139_));
 sg13g2_nand2_1 _2105_ (.Y(_1140_),
    .A(net486),
    .B(net474));
 sg13g2_o21ai_1 _2106_ (.B1(_0868_),
    .Y(_1141_),
    .A1(_0819_),
    .A2(_1138_));
 sg13g2_a22oi_1 _2107_ (.Y(_1142_),
    .B1(net570),
    .B2(net551),
    .A2(net503),
    .A1(net537));
 sg13g2_nor4_1 _2108_ (.A(_1052_),
    .B(_1106_),
    .C(_1139_),
    .D(_1141_),
    .Y(_1143_));
 sg13g2_nand4_1 _2109_ (.B(_0830_),
    .C(_0898_),
    .A(_0824_),
    .Y(_1144_),
    .D(_1136_));
 sg13g2_nand4_1 _2110_ (.B(_1060_),
    .C(_1137_),
    .A(_0886_),
    .Y(_1145_),
    .D(_1142_));
 sg13g2_nor4_1 _2111_ (.A(_1107_),
    .B(_1125_),
    .C(_1144_),
    .D(_1145_),
    .Y(_1146_));
 sg13g2_a21oi_1 _2112_ (.A1(_1143_),
    .A2(_1146_),
    .Y(_1147_),
    .B1(_0878_));
 sg13g2_a21o_1 _2113_ (.A2(_1146_),
    .A1(_1143_),
    .B1(_0878_),
    .X(_1148_));
 sg13g2_nor4_1 _2114_ (.A(_0940_),
    .B(_1123_),
    .C(_1134_),
    .D(_1147_),
    .Y(_1149_));
 sg13g2_nand3_1 _2115_ (.B(_1096_),
    .C(_1149_),
    .A(_1073_),
    .Y(_1150_));
 sg13g2_nand4_1 _2116_ (.B(_0764_),
    .C(_0774_),
    .A(_0762_),
    .Y(_1151_),
    .D(_0783_));
 sg13g2_a221oi_1 _2117_ (.B2(net560),
    .C1(_0941_),
    .B1(net498),
    .A1(net544),
    .Y(_1152_),
    .A2(_0787_));
 sg13g2_nand2_1 _2118_ (.Y(_1153_),
    .A(net554),
    .B(net468));
 sg13g2_o21ai_1 _2119_ (.B1(net479),
    .Y(_1154_),
    .A1(net540),
    .A2(net499));
 sg13g2_nand4_1 _2120_ (.B(_1152_),
    .C(_1153_),
    .A(_0925_),
    .Y(_1155_),
    .D(_1154_));
 sg13g2_nand3_1 _2121_ (.B(_0926_),
    .C(_0975_),
    .A(_0832_),
    .Y(_1156_));
 sg13g2_nand2_1 _2122_ (.Y(_1157_),
    .A(net559),
    .B(net539));
 sg13g2_a22oi_1 _2123_ (.Y(_1158_),
    .B1(net482),
    .B2(net543),
    .A2(net539),
    .A1(net559));
 sg13g2_a21oi_1 _2124_ (.A1(net539),
    .A2(net509),
    .Y(_1159_),
    .B1(_0938_));
 sg13g2_nand2_2 _2125_ (.Y(_1160_),
    .A(_1158_),
    .B(_1159_));
 sg13g2_a22oi_1 _2126_ (.Y(_1161_),
    .B1(net468),
    .B2(net495),
    .A2(net487),
    .A1(net544));
 sg13g2_nand2b_1 _2127_ (.Y(_1162_),
    .B(net469),
    .A_N(_0957_));
 sg13g2_nand2b_1 _2128_ (.Y(_1163_),
    .B(net474),
    .A_N(_1138_));
 sg13g2_nand2_1 _2129_ (.Y(_1164_),
    .A(net493),
    .B(net477));
 sg13g2_nand4_1 _2130_ (.B(_1057_),
    .C(_1161_),
    .A(_1004_),
    .Y(_1165_),
    .D(_1162_));
 sg13g2_nor4_1 _2131_ (.A(_1075_),
    .B(_1155_),
    .C(_1156_),
    .D(_1165_),
    .Y(_1166_));
 sg13g2_a22oi_1 _2132_ (.Y(_1167_),
    .B1(net493),
    .B2(net492),
    .A2(net500),
    .A1(net507));
 sg13g2_nand2_1 _2133_ (.Y(_1168_),
    .A(_1164_),
    .B(_1167_));
 sg13g2_nand4_1 _2134_ (.B(_1110_),
    .C(_1158_),
    .A(_1011_),
    .Y(_1169_),
    .D(_1159_));
 sg13g2_nand4_1 _2135_ (.B(_0976_),
    .C(_1009_),
    .A(_0900_),
    .Y(_1170_),
    .D(_1012_));
 sg13g2_a21oi_1 _2136_ (.A1(net546),
    .A2(net543),
    .Y(_1171_),
    .B1(_1001_));
 sg13g2_a21oi_1 _2137_ (.A1(net556),
    .A2(net474),
    .Y(_1172_),
    .B1(_0803_));
 sg13g2_nand4_1 _2138_ (.B(_1163_),
    .C(_1171_),
    .A(_0922_),
    .Y(_1173_),
    .D(_1172_));
 sg13g2_nor4_2 _2139_ (.A(_1168_),
    .B(_1169_),
    .C(_1170_),
    .Y(_1174_),
    .D(_1173_));
 sg13g2_a21oi_1 _2140_ (.A1(_1166_),
    .A2(_1174_),
    .Y(_1175_),
    .B1(_0858_));
 sg13g2_nand4_1 _2141_ (.B(_0901_),
    .C(_0918_),
    .A(_0899_),
    .Y(_1176_),
    .D(_0973_));
 sg13g2_a221oi_1 _2142_ (.B2(net512),
    .C1(_0814_),
    .B1(net467),
    .A1(net520),
    .Y(_1177_),
    .A2(net503));
 sg13g2_nand4_1 _2143_ (.B(_1031_),
    .C(_1098_),
    .A(_0971_),
    .Y(_1178_),
    .D(_1177_));
 sg13g2_a21o_1 _2144_ (.A2(net474),
    .A1(net518),
    .B1(_1033_),
    .X(_1179_));
 sg13g2_nand4_1 _2145_ (.B(_1034_),
    .C(_1045_),
    .A(_0949_),
    .Y(_1180_),
    .D(_1056_));
 sg13g2_nor4_1 _2146_ (.A(_0961_),
    .B(_1176_),
    .C(_1178_),
    .D(_1180_),
    .Y(_1181_));
 sg13g2_nand4_1 _2147_ (.B(_0889_),
    .C(_0912_),
    .A(_0888_),
    .Y(_1182_),
    .D(_1111_));
 sg13g2_nor2_1 _2148_ (.A(_0854_),
    .B(_1182_),
    .Y(_1183_));
 sg13g2_a21oi_1 _2149_ (.A1(_1181_),
    .A2(_1183_),
    .Y(_1184_),
    .B1(_0878_));
 sg13g2_a22oi_1 _2150_ (.Y(_1185_),
    .B1(net569),
    .B2(net553),
    .A2(net505),
    .A1(net534));
 sg13g2_o21ai_1 _2151_ (.B1(_1185_),
    .Y(_1186_),
    .A1(_0791_),
    .A2(_1138_));
 sg13g2_a21oi_1 _2152_ (.A1(_0791_),
    .A2(_0819_),
    .Y(_1187_),
    .B1(_0957_));
 sg13g2_nand3_1 _2153_ (.B(_0963_),
    .C(_1018_),
    .A(_0883_),
    .Y(_1188_));
 sg13g2_nor3_1 _2154_ (.A(_1186_),
    .B(_1187_),
    .C(_1188_),
    .Y(_1189_));
 sg13g2_o21ai_1 _2155_ (.B1(_0944_),
    .Y(_1190_),
    .A1(net591),
    .A2(_1189_));
 sg13g2_nor3_1 _2156_ (.A(_1175_),
    .B(_1184_),
    .C(_1190_),
    .Y(_1191_));
 sg13g2_nand3_1 _2157_ (.B(_1038_),
    .C(_1039_),
    .A(_1019_),
    .Y(_1192_));
 sg13g2_a21o_1 _2158_ (.A2(net490),
    .A1(net554),
    .B1(_0914_),
    .X(_1193_));
 sg13g2_nor4_1 _2159_ (.A(_1139_),
    .B(_1141_),
    .C(_1192_),
    .D(_1193_),
    .Y(_1194_));
 sg13g2_a21oi_1 _2160_ (.A1(net543),
    .A2(net511),
    .Y(_1195_),
    .B1(_0995_));
 sg13g2_nand2_1 _2161_ (.Y(_1196_),
    .A(net501),
    .B(net492));
 sg13g2_nand3_1 _2162_ (.B(_1195_),
    .C(_1196_),
    .A(_1157_),
    .Y(_1197_));
 sg13g2_nand2b_1 _2163_ (.Y(_1198_),
    .B(_0984_),
    .A_N(_0893_));
 sg13g2_nor4_2 _2164_ (.A(_0955_),
    .B(_0959_),
    .C(_1197_),
    .Y(_1199_),
    .D(_1198_));
 sg13g2_a21oi_1 _2165_ (.A1(net540),
    .A2(net468),
    .Y(_1200_),
    .B1(_1088_));
 sg13g2_nand2_1 _2166_ (.Y(_1201_),
    .A(net537),
    .B(net495));
 sg13g2_and4_1 _2167_ (.A(_1126_),
    .B(_1154_),
    .C(_1200_),
    .D(_1201_),
    .X(_1202_));
 sg13g2_nand3_1 _2168_ (.B(_1199_),
    .C(_1202_),
    .A(_1194_),
    .Y(_1203_));
 sg13g2_a21oi_1 _2169_ (.A1(net557),
    .A2(net544),
    .Y(_1204_),
    .B1(_0834_));
 sg13g2_a22oi_1 _2170_ (.Y(_1205_),
    .B1(net529),
    .B2(net498),
    .A2(net533),
    .A1(net544));
 sg13g2_a221oi_1 _2171_ (.B2(net524),
    .C1(_1000_),
    .B1(net466),
    .A1(net509),
    .Y(_1206_),
    .A2(net489));
 sg13g2_nand3_1 _2172_ (.B(_1205_),
    .C(_1206_),
    .A(_1204_),
    .Y(_1207_));
 sg13g2_o21ai_1 _2173_ (.B1(net526),
    .Y(_1208_),
    .A1(net552),
    .A2(net523));
 sg13g2_a22oi_1 _2174_ (.Y(_1209_),
    .B1(net499),
    .B2(net529),
    .A2(net510),
    .A1(net517));
 sg13g2_and2_1 _2175_ (.A(_1208_),
    .B(_1209_),
    .X(_1210_));
 sg13g2_nand2_1 _2176_ (.Y(_1211_),
    .A(_1208_),
    .B(_1209_));
 sg13g2_or4_2 _2177_ (.A(net598),
    .B(_0778_),
    .C(_0784_),
    .D(_0799_),
    .X(_1212_));
 sg13g2_nand3_1 _2178_ (.B(_1097_),
    .C(_1212_),
    .A(_1039_),
    .Y(_1213_));
 sg13g2_a21oi_1 _2179_ (.A1(net482),
    .A2(net473),
    .Y(_1214_),
    .B1(_1109_));
 sg13g2_a22oi_1 _2180_ (.Y(_1215_),
    .B1(net501),
    .B2(net492),
    .A2(net528),
    .A1(net539));
 sg13g2_a22oi_1 _2181_ (.Y(_1216_),
    .B1(net521),
    .B2(net534),
    .A2(net528),
    .A1(net546));
 sg13g2_nand4_1 _2182_ (.B(_1214_),
    .C(_1215_),
    .A(_0963_),
    .Y(_1217_),
    .D(_1216_));
 sg13g2_nor3_1 _2183_ (.A(_1211_),
    .B(_1213_),
    .C(_1217_),
    .Y(_1218_));
 sg13g2_nor4_2 _2184_ (.A(_0803_),
    .B(_0806_),
    .C(_0920_),
    .Y(_1219_),
    .D(_0921_));
 sg13g2_nand4_1 _2185_ (.B(_0882_),
    .C(_1112_),
    .A(_0869_),
    .Y(_1220_),
    .D(_1219_));
 sg13g2_nor2_1 _2186_ (.A(_1156_),
    .B(_1220_),
    .Y(_1221_));
 sg13g2_a21oi_1 _2187_ (.A1(_1218_),
    .A2(_1221_),
    .Y(_1222_),
    .B1(_0878_));
 sg13g2_a221oi_1 _2188_ (.B2(_0857_),
    .C1(_1222_),
    .B1(_1207_),
    .A1(_0760_),
    .Y(_1223_),
    .A2(_1203_));
 sg13g2_and4_1 _2189_ (.A(_0910_),
    .B(_1124_),
    .C(_1135_),
    .D(_1148_),
    .X(_1224_));
 sg13g2_and4_1 _2190_ (.A(_0981_),
    .B(_0982_),
    .C(_1004_),
    .D(_1005_),
    .X(_1225_));
 sg13g2_a22oi_1 _2191_ (.Y(_1226_),
    .B1(net495),
    .B2(net476),
    .A2(net516),
    .A1(net552));
 sg13g2_and4_1 _2192_ (.A(_1041_),
    .B(_1136_),
    .C(_1137_),
    .D(_1226_),
    .X(_1227_));
 sg13g2_o21ai_1 _2193_ (.B1(_1212_),
    .Y(_1228_),
    .A1(_0861_),
    .A2(_0957_));
 sg13g2_nand3_1 _2194_ (.B(_0954_),
    .C(_1151_),
    .A(_0866_),
    .Y(_1229_));
 sg13g2_nor4_2 _2195_ (.A(_1016_),
    .B(_1179_),
    .C(_1228_),
    .Y(_1230_),
    .D(_1229_));
 sg13g2_nand4_1 _2196_ (.B(_1225_),
    .C(_1227_),
    .A(_1210_),
    .Y(_1231_),
    .D(_1230_));
 sg13g2_a22oi_1 _2197_ (.Y(_1232_),
    .B1(net464),
    .B2(net548),
    .A2(net506),
    .A1(net531));
 sg13g2_a22oi_1 _2198_ (.Y(_1233_),
    .B1(net476),
    .B2(net557),
    .A2(net491),
    .A1(net549));
 sg13g2_nand4_1 _2199_ (.B(_1059_),
    .C(_1162_),
    .A(_0947_),
    .Y(_1234_),
    .D(_1233_));
 sg13g2_a21oi_1 _2200_ (.A1(net525),
    .A2(net480),
    .Y(_1235_),
    .B1(_0834_));
 sg13g2_nand4_1 _2201_ (.B(_0870_),
    .C(_1232_),
    .A(_0865_),
    .Y(_1236_),
    .D(_1235_));
 sg13g2_or4_1 _2202_ (.A(_1043_),
    .B(_1155_),
    .C(_1234_),
    .D(_1236_),
    .X(_1237_));
 sg13g2_o21ai_1 _2203_ (.B1(net472),
    .Y(_1238_),
    .A1(net526),
    .A2(net570));
 sg13g2_a22oi_1 _2204_ (.Y(_1239_),
    .B1(net472),
    .B2(net515),
    .A2(net490),
    .A1(net557));
 sg13g2_and3_1 _2205_ (.X(_1240_),
    .A(_1212_),
    .B(_1238_),
    .C(_1239_));
 sg13g2_a21oi_1 _2206_ (.A1(_1100_),
    .A2(_1240_),
    .Y(_1241_),
    .B1(_0858_));
 sg13g2_a221oi_1 _2207_ (.B2(_0877_),
    .C1(_1241_),
    .B1(_1237_),
    .A1(_0760_),
    .Y(_1242_),
    .A2(_1231_));
 sg13g2_a22oi_1 _2208_ (.Y(_1243_),
    .B1(net491),
    .B2(net484),
    .A2(net525),
    .A1(net560));
 sg13g2_a22oi_1 _2209_ (.Y(_1244_),
    .B1(net488),
    .B2(net535),
    .A2(net516),
    .A1(net522));
 sg13g2_nor3_1 _2210_ (.A(_1055_),
    .B(_1103_),
    .C(_1160_),
    .Y(_1245_));
 sg13g2_nand4_1 _2211_ (.B(_1036_),
    .C(_1057_),
    .A(_0859_),
    .Y(_1246_),
    .D(_1161_));
 sg13g2_a221oi_1 _2212_ (.B2(net504),
    .C1(_1108_),
    .B1(net486),
    .A1(net520),
    .Y(_1247_),
    .A2(net500));
 sg13g2_nand3_1 _2213_ (.B(_1243_),
    .C(_1247_),
    .A(_0897_),
    .Y(_1248_));
 sg13g2_nand2_1 _2214_ (.Y(_1249_),
    .A(_1226_),
    .B(_1244_));
 sg13g2_nor4_1 _2215_ (.A(_1193_),
    .B(_1246_),
    .C(_1248_),
    .D(_1249_),
    .Y(_1250_));
 sg13g2_a21o_1 _2216_ (.A2(_1250_),
    .A1(_1245_),
    .B1(_0878_),
    .X(_1251_));
 sg13g2_a221oi_1 _2217_ (.B2(net539),
    .C1(_0994_),
    .B1(net473),
    .A1(net553),
    .Y(_1252_),
    .A2(net512));
 sg13g2_a21oi_2 _2218_ (.B1(_0952_),
    .Y(_1253_),
    .A2(net501),
    .A1(net553));
 sg13g2_and4_1 _2219_ (.A(_0865_),
    .B(_0886_),
    .C(_1244_),
    .D(_1253_),
    .X(_1254_));
 sg13g2_a21oi_1 _2220_ (.A1(_1252_),
    .A2(_1254_),
    .Y(_1255_),
    .B1(net591));
 sg13g2_a22oi_1 _2221_ (.Y(_1256_),
    .B1(net466),
    .B2(net546),
    .A2(net478),
    .A1(net482));
 sg13g2_nand4_1 _2222_ (.B(_1140_),
    .C(_1196_),
    .A(_0974_),
    .Y(_1257_),
    .D(_1256_));
 sg13g2_a21oi_1 _2223_ (.A1(_0857_),
    .A2(_1257_),
    .Y(_1258_),
    .B1(_1255_));
 sg13g2_nand2_1 _2224_ (.Y(_1259_),
    .A(_1251_),
    .B(_1258_));
 sg13g2_and3_1 _2225_ (.X(_1260_),
    .A(_1242_),
    .B(_1251_),
    .C(_1258_));
 sg13g2_and3_2 _2226_ (.X(_1261_),
    .A(_0880_),
    .B(_1191_),
    .C(_1224_));
 sg13g2_and4_2 _2227_ (.A(_1073_),
    .B(_1096_),
    .C(_1223_),
    .D(_1260_),
    .X(_1262_));
 sg13g2_and2_1 _2228_ (.A(_1261_),
    .B(_1262_),
    .X(_1263_));
 sg13g2_a21oi_2 _2229_ (.B1(_1150_),
    .Y(_1264_),
    .A2(_1262_),
    .A1(_1261_));
 sg13g2_a21oi_2 _2230_ (.B1(_0945_),
    .Y(_1265_),
    .A2(_1262_),
    .A1(_1261_));
 sg13g2_nand2b_1 _2231_ (.Y(_1266_),
    .B(_0946_),
    .A_N(_1263_));
 sg13g2_and2_1 _2232_ (.A(_0760_),
    .B(_0817_),
    .X(_1267_));
 sg13g2_a21oi_2 _2233_ (.B1(_0858_),
    .Y(_1268_),
    .A2(_0863_),
    .A1(_0862_));
 sg13g2_nor3_1 _2234_ (.A(_0940_),
    .B(_1267_),
    .C(_1268_),
    .Y(_1269_));
 sg13g2_and2_1 _2235_ (.A(_0992_),
    .B(_1269_),
    .X(_1270_));
 sg13g2_and4_1 _2236_ (.A(_1223_),
    .B(_1224_),
    .C(_1242_),
    .D(_1270_),
    .X(_1271_));
 sg13g2_nand4_1 _2237_ (.B(_1224_),
    .C(_1242_),
    .A(_1223_),
    .Y(_1272_),
    .D(_1270_));
 sg13g2_nand2b_1 _2238_ (.Y(_0152_),
    .B(_0910_),
    .A_N(_0936_));
 sg13g2_nor2_1 _2239_ (.A(_0936_),
    .B(_0943_),
    .Y(_0153_));
 sg13g2_nand4_1 _2240_ (.B(_1073_),
    .C(_1260_),
    .A(_0910_),
    .Y(_0154_),
    .D(_0153_));
 sg13g2_a21oi_1 _2241_ (.A1(_1261_),
    .A2(_1262_),
    .Y(_0155_),
    .B1(_0154_));
 sg13g2_and4_2 _2242_ (.A(_0946_),
    .B(_1264_),
    .C(_1271_),
    .D(_0155_),
    .X(_0156_));
 sg13g2_nand4_1 _2243_ (.B(_1264_),
    .C(_1271_),
    .A(_0946_),
    .Y(_0157_),
    .D(_0155_));
 sg13g2_nand2_2 _2244_ (.Y(_0158_),
    .A(net177),
    .B(_0157_));
 sg13g2_and2_1 _2245_ (.A(_1150_),
    .B(_1272_),
    .X(_0159_));
 sg13g2_and2_1 _2246_ (.A(_1265_),
    .B(_0159_),
    .X(_0160_));
 sg13g2_or2_1 _2247_ (.X(_0161_),
    .B(_0160_),
    .A(_1072_));
 sg13g2_or3_1 _2248_ (.A(_1266_),
    .B(_0156_),
    .C(_0161_),
    .X(_0162_));
 sg13g2_xnor2_1 _2249_ (.Y(_0163_),
    .A(\main.demo._t___block_1_p4[2] ),
    .B(\main.demo._t___block_1_p4[0] ));
 sg13g2_xnor2_1 _2250_ (.Y(_0164_),
    .A(net169),
    .B(_0163_));
 sg13g2_inv_2 _2251_ (.Y(_0165_),
    .A(_0164_));
 sg13g2_nand2_1 _2252_ (.Y(_0166_),
    .A(_0162_),
    .B(_0165_));
 sg13g2_xnor2_1 _2253_ (.Y(_0167_),
    .A(_0162_),
    .B(_0164_));
 sg13g2_and2_1 _2254_ (.A(_1272_),
    .B(_0154_),
    .X(_0168_));
 sg13g2_or3_1 _2255_ (.A(_1264_),
    .B(_1265_),
    .C(_0168_),
    .X(_0169_));
 sg13g2_nand2_1 _2256_ (.Y(_0170_),
    .A(_0945_),
    .B(_1264_));
 sg13g2_nand2_2 _2257_ (.Y(_0171_),
    .A(_0169_),
    .B(_0170_));
 sg13g2_nand2_1 _2258_ (.Y(_0172_),
    .A(_1223_),
    .B(_1242_));
 sg13g2_nand3_1 _2259_ (.B(_1223_),
    .C(_1260_),
    .A(_0992_),
    .Y(_0173_));
 sg13g2_or2_1 _2260_ (.X(_0174_),
    .B(_0173_),
    .A(_0171_));
 sg13g2_xor2_1 _2261_ (.B(\main.demo._t___block_1_p4[0] ),
    .A(\main.demo._q_frame[0] ),
    .X(_0175_));
 sg13g2_xnor2_1 _2262_ (.Y(_0176_),
    .A(\main.demo._q_frame[0] ),
    .B(\main.demo._t___block_1_p4[0] ));
 sg13g2_nor2_1 _2263_ (.A(_0174_),
    .B(_0175_),
    .Y(_0177_));
 sg13g2_xnor2_1 _2264_ (.Y(_0178_),
    .A(\main.demo._q_frame[0] ),
    .B(\main.demo._t___block_1_p4[1] ));
 sg13g2_nor2_1 _2265_ (.A(_0156_),
    .B(_0178_),
    .Y(_0179_));
 sg13g2_or2_1 _2266_ (.X(_0180_),
    .B(_0178_),
    .A(_0156_));
 sg13g2_a21oi_1 _2267_ (.A1(_1271_),
    .A2(_0155_),
    .Y(_0181_),
    .B1(_1265_));
 sg13g2_nand2b_1 _2268_ (.Y(_0182_),
    .B(_1264_),
    .A_N(_0168_));
 sg13g2_nand2b_1 _2269_ (.Y(_0183_),
    .B(_0168_),
    .A_N(_1264_));
 sg13g2_o21ai_1 _2270_ (.B1(_0183_),
    .Y(_0184_),
    .A1(_0181_),
    .A2(_0182_));
 sg13g2_xnor2_1 _2271_ (.Y(_0185_),
    .A(\main.demo._t___block_1_p4[3] ),
    .B(_0178_));
 sg13g2_xor2_1 _2272_ (.B(_0178_),
    .A(\main.demo._t___block_1_p4[3] ),
    .X(_0186_));
 sg13g2_o21ai_1 _2273_ (.B1(_0186_),
    .Y(_0187_),
    .A1(_0180_),
    .A2(_0184_));
 sg13g2_nor3_1 _2274_ (.A(\main.demo._t___block_1_p4[3] ),
    .B(_0180_),
    .C(_0184_),
    .Y(_0188_));
 sg13g2_or2_1 _2275_ (.X(_0189_),
    .B(_1263_),
    .A(_0936_));
 sg13g2_nor4_1 _2276_ (.A(_0946_),
    .B(_1150_),
    .C(_1263_),
    .D(_1272_),
    .Y(_0190_));
 sg13g2_nor2_2 _2277_ (.A(_1267_),
    .B(_1268_),
    .Y(_0191_));
 sg13g2_o21ai_1 _2278_ (.B1(_0191_),
    .Y(_0192_),
    .A1(_1266_),
    .A2(_0154_));
 sg13g2_or4_1 _2279_ (.A(_0172_),
    .B(_0189_),
    .C(_0190_),
    .D(_0192_),
    .X(_0193_));
 sg13g2_a221oi_1 _2280_ (.B2(_0193_),
    .C1(_0188_),
    .B1(_0187_),
    .A1(_0174_),
    .Y(_0194_),
    .A2(_0175_));
 sg13g2_nor2_1 _2281_ (.A(_0177_),
    .B(_0194_),
    .Y(_0195_));
 sg13g2_nand2_1 _2282_ (.Y(_0196_),
    .A(_0167_),
    .B(_0195_));
 sg13g2_a21oi_1 _2283_ (.A1(_0166_),
    .A2(_0196_),
    .Y(_0022_),
    .B1(_0158_));
 sg13g2_nand2_1 _2284_ (.Y(_0197_),
    .A(_0165_),
    .B(_0171_));
 sg13g2_or2_1 _2285_ (.X(_0198_),
    .B(_0189_),
    .A(_0943_));
 sg13g2_nor4_2 _2286_ (.A(_0156_),
    .B(_0161_),
    .C(_0172_),
    .Y(_0199_),
    .D(_0198_));
 sg13g2_nor2_1 _2287_ (.A(_0176_),
    .B(_0199_),
    .Y(_0200_));
 sg13g2_or2_1 _2288_ (.X(_0201_),
    .B(_0190_),
    .A(_0160_));
 sg13g2_and2_1 _2289_ (.A(_1260_),
    .B(_0191_),
    .X(_0202_));
 sg13g2_o21ai_1 _2290_ (.B1(_0202_),
    .Y(_0203_),
    .A1(_1264_),
    .A2(_1265_));
 sg13g2_o21ai_1 _2291_ (.B1(_0179_),
    .Y(_0204_),
    .A1(_0201_),
    .A2(_0203_));
 sg13g2_nand2b_1 _2292_ (.Y(_0205_),
    .B(_0191_),
    .A_N(_1263_));
 sg13g2_nor2_1 _2293_ (.A(_1266_),
    .B(_1272_),
    .Y(_0206_));
 sg13g2_nor3_2 _2294_ (.A(_0159_),
    .B(_0205_),
    .C(_0206_),
    .Y(_0207_));
 sg13g2_o21ai_1 _2295_ (.B1(_0204_),
    .Y(_0208_),
    .A1(_0186_),
    .A2(_0207_));
 sg13g2_a22oi_1 _2296_ (.Y(_0209_),
    .B1(_0207_),
    .B2(_0186_),
    .A2(_0199_),
    .A1(_0176_));
 sg13g2_a21oi_2 _2297_ (.B1(_0200_),
    .Y(_0210_),
    .A2(_0209_),
    .A1(_0208_));
 sg13g2_xnor2_1 _2298_ (.Y(_0211_),
    .A(_0165_),
    .B(_0171_));
 sg13g2_or2_1 _2299_ (.X(_0212_),
    .B(_0211_),
    .A(_0210_));
 sg13g2_a21oi_1 _2300_ (.A1(_0197_),
    .A2(_0212_),
    .Y(_0023_),
    .B1(_0158_));
 sg13g2_or2_1 _2301_ (.X(_0213_),
    .B(_0205_),
    .A(_0943_));
 sg13g2_nand2_1 _2302_ (.Y(_0214_),
    .A(_0165_),
    .B(_0213_));
 sg13g2_xnor2_1 _2303_ (.Y(_0215_),
    .A(_0165_),
    .B(_0213_));
 sg13g2_nand3_1 _2304_ (.B(_0157_),
    .C(_0169_),
    .A(_0910_),
    .Y(_0216_));
 sg13g2_nor2_1 _2305_ (.A(_0201_),
    .B(_0216_),
    .Y(_0217_));
 sg13g2_nor2_1 _2306_ (.A(_0176_),
    .B(_0217_),
    .Y(_0218_));
 sg13g2_nor2_1 _2307_ (.A(_0880_),
    .B(_1272_),
    .Y(_0219_));
 sg13g2_nor3_1 _2308_ (.A(_1072_),
    .B(_1263_),
    .C(_0219_),
    .Y(_0220_));
 sg13g2_nand4_1 _2309_ (.B(_1242_),
    .C(_0157_),
    .A(_1223_),
    .Y(_0221_),
    .D(_0220_));
 sg13g2_nor4_1 _2310_ (.A(_0933_),
    .B(_1072_),
    .C(_1259_),
    .D(_0152_),
    .Y(_0222_));
 sg13g2_a21o_1 _2311_ (.A2(_0222_),
    .A1(_0191_),
    .B1(_0180_),
    .X(_0223_));
 sg13g2_nand2_1 _2312_ (.Y(_0224_),
    .A(_0185_),
    .B(_0221_));
 sg13g2_nor2_1 _2313_ (.A(_0185_),
    .B(_0221_),
    .Y(_0225_));
 sg13g2_a221oi_1 _2314_ (.B2(_0224_),
    .C1(_0225_),
    .B1(_0223_),
    .A1(_0176_),
    .Y(_0226_),
    .A2(_0217_));
 sg13g2_nor2_1 _2315_ (.A(_0218_),
    .B(_0226_),
    .Y(_0227_));
 sg13g2_or2_1 _2316_ (.X(_0228_),
    .B(_0227_),
    .A(_0215_));
 sg13g2_a21oi_1 _2317_ (.A1(_0214_),
    .A2(_0228_),
    .Y(_0024_),
    .B1(_0158_));
 sg13g2_or2_1 _2318_ (.X(_0229_),
    .B(_0195_),
    .A(_0167_));
 sg13g2_and4_1 _2319_ (.A(net177),
    .B(_0157_),
    .C(_0196_),
    .D(_0229_),
    .X(_0025_));
 sg13g2_xnor2_1 _2320_ (.Y(_0230_),
    .A(_0210_),
    .B(_0211_));
 sg13g2_nor2_1 _2321_ (.A(_0158_),
    .B(_0230_),
    .Y(_0026_));
 sg13g2_a21oi_1 _2322_ (.A1(_0215_),
    .A2(_0227_),
    .Y(_0231_),
    .B1(_0158_));
 sg13g2_and2_1 _2323_ (.A(_0228_),
    .B(_0231_),
    .X(_0027_));
 sg13g2_nand2_1 _2324_ (.Y(_0232_),
    .A(\main.demo.vga._q_ycount[3] ),
    .B(\main.demo.vga._q_ycount[2] ));
 sg13g2_and2_1 _2325_ (.A(net211),
    .B(_0620_),
    .X(_0233_));
 sg13g2_nand2_2 _2326_ (.Y(_0234_),
    .A(_0620_),
    .B(_0629_));
 sg13g2_nand3_1 _2327_ (.B(net397),
    .C(_0622_),
    .A(\main.demo.vga._q_ycount[1] ),
    .Y(_0235_));
 sg13g2_or2_1 _2328_ (.X(_0236_),
    .B(_0235_),
    .A(_0232_));
 sg13g2_nor2_1 _2329_ (.A(_0597_),
    .B(_0236_),
    .Y(_0237_));
 sg13g2_and4_1 _2330_ (.A(net251),
    .B(\main.demo.vga._q_ycount[2] ),
    .C(\main.demo.vga._q_ycount[1] ),
    .D(\main.demo.vga._q_ycount[0] ),
    .X(_0238_));
 sg13g2_and4_1 _2331_ (.A(\main.demo.vga._q_ycount[5] ),
    .B(\main.demo.vga._q_ycount[4] ),
    .C(_0620_),
    .D(_0238_),
    .X(_0239_));
 sg13g2_and2_1 _2332_ (.A(net279),
    .B(_0239_),
    .X(_0240_));
 sg13g2_nand3_1 _2333_ (.B(net314),
    .C(_0240_),
    .A(net382),
    .Y(_0241_));
 sg13g2_xor2_1 _2334_ (.B(_0241_),
    .A(net349),
    .X(_0242_));
 sg13g2_a21oi_1 _2335_ (.A1(_0234_),
    .A2(net350),
    .Y(_0028_),
    .B1(net595));
 sg13g2_nor2b_1 _2336_ (.A(\main._w_demo_video_hs ),
    .B_N(\main.demo._q_prev_hs ),
    .Y(_0243_));
 sg13g2_nand2b_2 _2337_ (.Y(_0244_),
    .B(\main.demo._q_prev_hs ),
    .A_N(\main._w_demo_video_hs ));
 sg13g2_nor2_1 _2338_ (.A(net166),
    .B(_0244_),
    .Y(_0245_));
 sg13g2_nand2_1 _2339_ (.Y(_0246_),
    .A(net164),
    .B(net612));
 sg13g2_nor2_1 _2340_ (.A(\main.demo._q_v[0] ),
    .B(net566),
    .Y(_0247_));
 sg13g2_nor3_1 _2341_ (.A(_0245_),
    .B(net565),
    .C(_0247_),
    .Y(_0029_));
 sg13g2_and3_1 _2342_ (.X(_0248_),
    .A(net196),
    .B(\main.demo._q_v[0] ),
    .C(net566));
 sg13g2_a21oi_1 _2343_ (.A1(\main.demo._q_v[0] ),
    .A2(net566),
    .Y(_0249_),
    .B1(net196));
 sg13g2_nor3_1 _2344_ (.A(net565),
    .B(_0248_),
    .C(net197),
    .Y(_0030_));
 sg13g2_nor2_1 _2345_ (.A(net255),
    .B(_0248_),
    .Y(_0250_));
 sg13g2_and2_1 _2346_ (.A(net255),
    .B(_0248_),
    .X(_0251_));
 sg13g2_nor3_1 _2347_ (.A(net564),
    .B(net256),
    .C(_0251_),
    .Y(_0031_));
 sg13g2_nor2_1 _2348_ (.A(net286),
    .B(_0251_),
    .Y(_0252_));
 sg13g2_and2_1 _2349_ (.A(net286),
    .B(_0251_),
    .X(_0253_));
 sg13g2_nor3_1 _2350_ (.A(net564),
    .B(_0252_),
    .C(_0253_),
    .Y(_0032_));
 sg13g2_nor2_1 _2351_ (.A(net244),
    .B(_0253_),
    .Y(_0254_));
 sg13g2_and2_1 _2352_ (.A(net244),
    .B(_0253_),
    .X(_0255_));
 sg13g2_nor3_1 _2353_ (.A(net564),
    .B(net245),
    .C(_0255_),
    .Y(_0033_));
 sg13g2_xnor2_1 _2354_ (.Y(_0256_),
    .A(net317),
    .B(_0255_));
 sg13g2_nor2_1 _2355_ (.A(net564),
    .B(_0256_),
    .Y(_0034_));
 sg13g2_a21oi_1 _2356_ (.A1(\main.demo._q_v[5] ),
    .A2(_0255_),
    .Y(_0257_),
    .B1(net234));
 sg13g2_and3_1 _2357_ (.X(_0258_),
    .A(net234),
    .B(net402),
    .C(_0255_));
 sg13g2_nor3_1 _2358_ (.A(net565),
    .B(net235),
    .C(_0258_),
    .Y(_0035_));
 sg13g2_nor2b_1 _2359_ (.A(net224),
    .B_N(net192),
    .Y(_0036_));
 sg13g2_nor2b_1 _2360_ (.A(_0625_),
    .B_N(net193),
    .Y(_0037_));
 sg13g2_and2_1 _2361_ (.A(net612),
    .B(_0632_),
    .X(_0038_));
 sg13g2_nand4_1 _2362_ (.B(\main.demo.vga._q_ycount[7] ),
    .C(\main.demo.vga._q_ycount[6] ),
    .A(\main.demo.vga._q_ycount[8] ),
    .Y(_0259_),
    .D(\main.demo.vga._d_vblank ));
 sg13g2_or3_1 _2363_ (.A(\main.demo.vga._q_ycount[5] ),
    .B(_0597_),
    .C(_0259_),
    .X(_0260_));
 sg13g2_nor3_1 _2364_ (.A(net211),
    .B(_0232_),
    .C(_0260_),
    .Y(_0261_));
 sg13g2_a21oi_1 _2365_ (.A1(\main.demo.vga._q_ycount[1] ),
    .A2(_0261_),
    .Y(_0262_),
    .B1(net164));
 sg13g2_nor3_1 _2366_ (.A(\main.demo.vga._q_ycount[1] ),
    .B(_0232_),
    .C(_0260_),
    .Y(_0263_));
 sg13g2_a21oi_1 _2367_ (.A1(net211),
    .A2(_0263_),
    .Y(_0039_),
    .B1(_0262_));
 sg13g2_and2_1 _2368_ (.A(net192),
    .B(net193),
    .X(_0264_));
 sg13g2_and3_2 _2369_ (.X(_0265_),
    .A(net282),
    .B(net183),
    .C(_0264_));
 sg13g2_nand3_1 _2370_ (.B(net237),
    .C(\main.demo.vga._q_xcount[10] ),
    .A(\main.demo.vga._q_xcount[8] ),
    .Y(_0266_));
 sg13g2_nand2_1 _2371_ (.Y(_0267_),
    .A(\main.demo.vga._q_xcount[6] ),
    .B(net220));
 sg13g2_nor4_1 _2372_ (.A(\main.demo.vga._q_xcount[4] ),
    .B(net336),
    .C(_0266_),
    .D(_0267_),
    .Y(_0268_));
 sg13g2_a21oi_1 _2373_ (.A1(_0265_),
    .A2(net337),
    .Y(_0269_),
    .B1(net173));
 sg13g2_nand3_1 _2374_ (.B(net336),
    .C(\main.demo.vga._q_xcount[6] ),
    .A(\main.demo.vga._q_xcount[4] ),
    .Y(_0270_));
 sg13g2_nor2_1 _2375_ (.A(_0266_),
    .B(_0270_),
    .Y(_0271_));
 sg13g2_a21oi_1 _2376_ (.A1(_0623_),
    .A2(_0271_),
    .Y(_0040_),
    .B1(_0269_));
 sg13g2_nor2_1 _2377_ (.A(net595),
    .B(_0625_),
    .Y(_0041_));
 sg13g2_nor2_1 _2378_ (.A(net192),
    .B(net595),
    .Y(_0042_));
 sg13g2_and3_1 _2379_ (.X(_0272_),
    .A(\main.demo.vga._q_xcount[4] ),
    .B(\main.demo.vga._q_xcount[5] ),
    .C(_0265_));
 sg13g2_a21oi_1 _2380_ (.A1(net339),
    .A2(_0265_),
    .Y(_0273_),
    .B1(net336));
 sg13g2_o21ai_1 _2381_ (.B1(_0621_),
    .Y(_0274_),
    .A1(_0272_),
    .A2(_0273_));
 sg13g2_and2_1 _2382_ (.A(net613),
    .B(_0274_),
    .X(_0043_));
 sg13g2_xnor2_1 _2383_ (.Y(_0275_),
    .A(net362),
    .B(_0272_));
 sg13g2_a21oi_1 _2384_ (.A1(_0621_),
    .A2(net363),
    .Y(_0044_),
    .B1(net596));
 sg13g2_nor2b_2 _2385_ (.A(_0267_),
    .B_N(_0272_),
    .Y(_0276_));
 sg13g2_xnor2_1 _2386_ (.Y(_0277_),
    .A(net378),
    .B(_0276_));
 sg13g2_a21oi_1 _2387_ (.A1(_0621_),
    .A2(_0277_),
    .Y(_0045_),
    .B1(net596));
 sg13g2_a21oi_1 _2388_ (.A1(\main.demo.vga._q_xcount[8] ),
    .A2(_0276_),
    .Y(_0278_),
    .B1(net237));
 sg13g2_nand3_1 _2389_ (.B(net237),
    .C(_0276_),
    .A(net401),
    .Y(_0279_));
 sg13g2_nand2_1 _2390_ (.Y(_0280_),
    .A(net612),
    .B(_0279_));
 sg13g2_nor2_1 _2391_ (.A(net238),
    .B(_0280_),
    .Y(_0046_));
 sg13g2_xor2_1 _2392_ (.B(_0279_),
    .A(net353),
    .X(_0281_));
 sg13g2_a21oi_1 _2393_ (.A1(_0621_),
    .A2(_0281_),
    .Y(_0047_),
    .B1(net596));
 sg13g2_nand2_1 _2394_ (.Y(_0282_),
    .A(net613),
    .B(_0234_));
 sg13g2_nor2_1 _2395_ (.A(net211),
    .B(_0620_),
    .Y(_0283_));
 sg13g2_nor3_1 _2396_ (.A(_0233_),
    .B(_0282_),
    .C(_0283_),
    .Y(_0048_));
 sg13g2_or2_1 _2397_ (.X(_0284_),
    .B(_0233_),
    .A(net308));
 sg13g2_and3_1 _2398_ (.X(_0049_),
    .A(net612),
    .B(_0235_),
    .C(_0284_));
 sg13g2_nand3_1 _2399_ (.B(\main.demo.vga._q_ycount[1] ),
    .C(_0233_),
    .A(\main.demo.vga._q_ycount[2] ),
    .Y(_0285_));
 sg13g2_xor2_1 _2400_ (.B(_0235_),
    .A(net373),
    .X(_0286_));
 sg13g2_a21oi_1 _2401_ (.A1(_0234_),
    .A2(net374),
    .Y(_0050_),
    .B1(net595));
 sg13g2_a221oi_1 _2402_ (.B2(_0598_),
    .C1(net595),
    .B1(_0285_),
    .A1(_0620_),
    .Y(_0051_),
    .A2(_0238_));
 sg13g2_xnor2_1 _2403_ (.Y(_0287_),
    .A(_0597_),
    .B(_0236_));
 sg13g2_a21oi_1 _2404_ (.A1(_0234_),
    .A2(_0287_),
    .Y(_0052_),
    .B1(net595));
 sg13g2_xnor2_1 _2405_ (.Y(_0288_),
    .A(net329),
    .B(_0237_));
 sg13g2_nor2_1 _2406_ (.A(_0282_),
    .B(net330),
    .Y(_0053_));
 sg13g2_nor2_1 _2407_ (.A(net279),
    .B(_0239_),
    .Y(_0289_));
 sg13g2_nor3_1 _2408_ (.A(net595),
    .B(_0240_),
    .C(net280),
    .Y(_0054_));
 sg13g2_xnor2_1 _2409_ (.Y(_0290_),
    .A(net314),
    .B(_0240_));
 sg13g2_nor2_1 _2410_ (.A(net595),
    .B(_0290_),
    .Y(_0055_));
 sg13g2_a21o_1 _2411_ (.A2(_0240_),
    .A1(net314),
    .B1(net382),
    .X(_0291_));
 sg13g2_and3_1 _2412_ (.X(_0056_),
    .A(net612),
    .B(_0241_),
    .C(_0291_));
 sg13g2_a21oi_1 _2413_ (.A1(net303),
    .A2(_0258_),
    .Y(_0292_),
    .B1(net565));
 sg13g2_o21ai_1 _2414_ (.B1(_0292_),
    .Y(_0293_),
    .A1(net303),
    .A2(_0258_));
 sg13g2_inv_1 _2415_ (.Y(_0057_),
    .A(_0293_));
 sg13g2_nor3_1 _2416_ (.A(\main.demo.zic._q_clock_count[7] ),
    .B(\main.demo.zic._q_clock_count[6] ),
    .C(\main.demo.zic._q_clock_count[8] ),
    .Y(_0294_));
 sg13g2_nor2_1 _2417_ (.A(\main.demo.zic._q_clock_count[1] ),
    .B(net357),
    .Y(_0295_));
 sg13g2_nor4_1 _2418_ (.A(\main.demo.zic._q_clock_count[3] ),
    .B(\main.demo.zic._q_clock_count[2] ),
    .C(\main.demo.zic._q_clock_count[5] ),
    .D(\main.demo.zic._q_clock_count[4] ),
    .Y(_0296_));
 sg13g2_and3_1 _2419_ (.X(_0297_),
    .A(_0294_),
    .B(_0295_),
    .C(_0296_));
 sg13g2_nand3_1 _2420_ (.B(_0295_),
    .C(_0296_),
    .A(_0294_),
    .Y(_0298_));
 sg13g2_nor2_1 _2421_ (.A(\main.demo.zic._q_idx[4] ),
    .B(_0015_),
    .Y(_0299_));
 sg13g2_nand2b_1 _2422_ (.Y(_0300_),
    .B(\main.demo.zic._q_idx[0] ),
    .A_N(\main.demo.zic._q_idx[1] ));
 sg13g2_xnor2_1 _2423_ (.Y(_0301_),
    .A(\main.demo.zic._q_idx[0] ),
    .B(\main.demo.zic._q_idx[1] ));
 sg13g2_xor2_1 _2424_ (.B(\main.demo.zic._q_idx[1] ),
    .A(\main.demo.zic._q_idx[0] ),
    .X(_0302_));
 sg13g2_nand2_1 _2425_ (.Y(_0303_),
    .A(\main.demo.zic._q_idx[0] ),
    .B(\main.demo.zic._q_idx[1] ));
 sg13g2_nand3b_1 _2426_ (.B(\main.demo.zic._q_idx[1] ),
    .C(_0015_),
    .Y(_0304_),
    .A_N(\main.demo.zic._q_idx[0] ));
 sg13g2_o21ai_1 _2427_ (.B1(_0304_),
    .Y(_0305_),
    .A1(\main.demo.zic._q_idx[4] ),
    .A2(_0303_));
 sg13g2_nand2b_1 _2428_ (.Y(_0306_),
    .B(\main.demo.zic._q_idx[3] ),
    .A_N(\main.demo.zic._q_idx[2] ));
 sg13g2_a21oi_1 _2429_ (.A1(\main.demo.zic._q_idx[0] ),
    .A2(_0299_),
    .Y(_0307_),
    .B1(_0306_));
 sg13g2_and2_1 _2430_ (.A(_0301_),
    .B(_0307_),
    .X(_0308_));
 sg13g2_nor2_1 _2431_ (.A(_0600_),
    .B(_0601_),
    .Y(_0309_));
 sg13g2_nand2_1 _2432_ (.Y(_0310_),
    .A(\main.demo.zic._q_idx[3] ),
    .B(\main.demo.zic._q_idx[2] ));
 sg13g2_a21o_1 _2433_ (.A2(_0309_),
    .A1(_0305_),
    .B1(_0308_),
    .X(_0311_));
 sg13g2_or4_1 _2434_ (.A(\main.demo.zic._q_idx[3] ),
    .B(_0601_),
    .C(_0299_),
    .D(_0300_),
    .X(_0312_));
 sg13g2_inv_1 _2435_ (.Y(_0313_),
    .A(_0312_));
 sg13g2_and4_1 _2436_ (.A(_0600_),
    .B(_0601_),
    .C(_0300_),
    .D(_0302_),
    .X(_0314_));
 sg13g2_a22oi_1 _2437_ (.Y(_0315_),
    .B1(_0302_),
    .B2(_0601_),
    .A2(_0300_),
    .A1(_0600_));
 sg13g2_or3_1 _2438_ (.A(_0299_),
    .B(_0314_),
    .C(_0315_),
    .X(_0316_));
 sg13g2_nor3_1 _2439_ (.A(\main.demo.zic._q_idx[1] ),
    .B(_0603_),
    .C(_0310_),
    .Y(_0317_));
 sg13g2_a221oi_1 _2440_ (.B2(_0305_),
    .C1(_0317_),
    .B1(_0309_),
    .A1(_0301_),
    .Y(_0318_),
    .A2(_0307_));
 sg13g2_and2_1 _2441_ (.A(_0316_),
    .B(_0318_),
    .X(_0319_));
 sg13g2_nand3_1 _2442_ (.B(_0316_),
    .C(_0318_),
    .A(_0312_),
    .Y(_0320_));
 sg13g2_a21oi_1 _2443_ (.A1(_0602_),
    .A2(_0303_),
    .Y(_0321_),
    .B1(_0310_));
 sg13g2_o21ai_1 _2444_ (.B1(_0321_),
    .Y(_0322_),
    .A1(_0603_),
    .A2(_0303_));
 sg13g2_and4_1 _2445_ (.A(_0312_),
    .B(_0316_),
    .C(_0318_),
    .D(_0322_),
    .X(_0323_));
 sg13g2_or2_1 _2446_ (.X(_0324_),
    .B(_0323_),
    .A(_0311_));
 sg13g2_a21oi_1 _2447_ (.A1(net463),
    .A2(_0324_),
    .Y(_0325_),
    .B1(net174));
 sg13g2_o21ai_1 _2448_ (.B1(net174),
    .Y(_0326_),
    .A1(_0311_),
    .A2(_0323_));
 sg13g2_o21ai_1 _2449_ (.B1(net610),
    .Y(_0327_),
    .A1(_0298_),
    .A2(_0326_));
 sg13g2_nor2_1 _2450_ (.A(_0325_),
    .B(_0327_),
    .Y(_0058_));
 sg13g2_nor2b_1 _2451_ (.A(_0009_),
    .B_N(_0320_),
    .Y(_0328_));
 sg13g2_xor2_1 _2452_ (.B(_0320_),
    .A(_0009_),
    .X(_0329_));
 sg13g2_nor2_1 _2453_ (.A(_0326_),
    .B(_0329_),
    .Y(_0330_));
 sg13g2_xnor2_1 _2454_ (.Y(_0331_),
    .A(_0326_),
    .B(_0329_));
 sg13g2_o21ai_1 _2455_ (.B1(net609),
    .Y(_0332_),
    .A1(net216),
    .A2(net463));
 sg13g2_a21oi_1 _2456_ (.A1(net462),
    .A2(_0331_),
    .Y(_0059_),
    .B1(_0332_));
 sg13g2_nand2_1 _2457_ (.Y(_0333_),
    .A(\main.demo.zic._q_qpos[2] ),
    .B(_0324_));
 sg13g2_xor2_1 _2458_ (.B(_0324_),
    .A(\main.demo.zic._q_qpos[2] ),
    .X(_0334_));
 sg13g2_o21ai_1 _2459_ (.B1(_0334_),
    .Y(_0335_),
    .A1(_0328_),
    .A2(_0330_));
 sg13g2_or3_1 _2460_ (.A(_0328_),
    .B(_0330_),
    .C(_0334_),
    .X(_0336_));
 sg13g2_nand2_1 _2461_ (.Y(_0337_),
    .A(_0335_),
    .B(_0336_));
 sg13g2_o21ai_1 _2462_ (.B1(net609),
    .Y(_0338_),
    .A1(net313),
    .A2(net463));
 sg13g2_a21oi_1 _2463_ (.A1(net462),
    .A2(_0337_),
    .Y(_0060_),
    .B1(_0338_));
 sg13g2_xnor2_1 _2464_ (.Y(_0339_),
    .A(_0010_),
    .B(_0319_));
 sg13g2_a21o_1 _2465_ (.A2(_0335_),
    .A1(_0333_),
    .B1(_0339_),
    .X(_0340_));
 sg13g2_nand3_1 _2466_ (.B(_0335_),
    .C(_0339_),
    .A(_0333_),
    .Y(_0341_));
 sg13g2_nand2_1 _2467_ (.Y(_0342_),
    .A(_0340_),
    .B(_0341_));
 sg13g2_o21ai_1 _2468_ (.B1(net609),
    .Y(_0343_),
    .A1(net218),
    .A2(net462));
 sg13g2_a21oi_1 _2469_ (.A1(net462),
    .A2(_0342_),
    .Y(_0061_),
    .B1(_0343_));
 sg13g2_nor2_1 _2470_ (.A(_0313_),
    .B(_0323_),
    .Y(_0344_));
 sg13g2_nor2b_1 _2471_ (.A(_0344_),
    .B_N(\main.demo.zic._q_qpos[4] ),
    .Y(_0345_));
 sg13g2_xnor2_1 _2472_ (.Y(_0346_),
    .A(\main.demo.zic._q_qpos[4] ),
    .B(_0344_));
 sg13g2_o21ai_1 _2473_ (.B1(_0340_),
    .Y(_0347_),
    .A1(_0010_),
    .A2(_0319_));
 sg13g2_xnor2_1 _2474_ (.Y(_0348_),
    .A(_0346_),
    .B(_0347_));
 sg13g2_o21ai_1 _2475_ (.B1(net609),
    .Y(_0349_),
    .A1(net309),
    .A2(net462));
 sg13g2_a21oi_1 _2476_ (.A1(net462),
    .A2(_0348_),
    .Y(_0062_),
    .B1(_0349_));
 sg13g2_a21oi_2 _2477_ (.B1(_0345_),
    .Y(_0350_),
    .A2(_0347_),
    .A1(_0346_));
 sg13g2_nor3_2 _2478_ (.A(_0011_),
    .B(_0298_),
    .C(_0350_),
    .Y(_0351_));
 sg13g2_and3_1 _2479_ (.X(_0352_),
    .A(_0011_),
    .B(net462),
    .C(_0350_));
 sg13g2_o21ai_1 _2480_ (.B1(net611),
    .Y(_0353_),
    .A1(net228),
    .A2(net462));
 sg13g2_nor3_1 _2481_ (.A(_0011_),
    .B(_0298_),
    .C(_0350_),
    .Y(_0354_));
 sg13g2_nor3_1 _2482_ (.A(_0351_),
    .B(_0352_),
    .C(net229),
    .Y(_0063_));
 sg13g2_nand2_1 _2483_ (.Y(_0355_),
    .A(net319),
    .B(_0351_));
 sg13g2_o21ai_1 _2484_ (.B1(net609),
    .Y(_0356_),
    .A1(net319),
    .A2(_0351_));
 sg13g2_nor2b_1 _2485_ (.A(net320),
    .B_N(_0355_),
    .Y(_0064_));
 sg13g2_a21oi_1 _2486_ (.A1(\main.demo.zic._q_qpos[6] ),
    .A2(_0351_),
    .Y(_0357_),
    .B1(net189));
 sg13g2_and3_1 _2487_ (.X(_0358_),
    .A(net189),
    .B(\main.demo.zic._q_qpos[6] ),
    .C(_0354_));
 sg13g2_nor3_1 _2488_ (.A(net592),
    .B(net190),
    .C(_0358_),
    .Y(_0065_));
 sg13g2_nor2_1 _2489_ (.A(net287),
    .B(_0358_),
    .Y(_0359_));
 sg13g2_nor3_1 _2490_ (.A(_0595_),
    .B(_0596_),
    .C(_0355_),
    .Y(_0360_));
 sg13g2_nor3_1 _2491_ (.A(net592),
    .B(net288),
    .C(_0360_),
    .Y(_0066_));
 sg13g2_or2_1 _2492_ (.X(_0361_),
    .B(_0360_),
    .A(net381));
 sg13g2_nand3_1 _2493_ (.B(net287),
    .C(_0358_),
    .A(net381),
    .Y(_0362_));
 sg13g2_and3_1 _2494_ (.X(_0067_),
    .A(net609),
    .B(_0361_),
    .C(_0362_));
 sg13g2_nand2b_1 _2495_ (.Y(_0363_),
    .B(_0362_),
    .A_N(net341));
 sg13g2_nand4_1 _2496_ (.B(\main.demo.zic._q_qpos[9] ),
    .C(net287),
    .A(net341),
    .Y(_0364_),
    .D(_0358_));
 sg13g2_and3_1 _2497_ (.X(_0068_),
    .A(net609),
    .B(net342),
    .C(_0364_));
 sg13g2_nor2b_1 _2498_ (.A(net178),
    .B_N(_0364_),
    .Y(_0365_));
 sg13g2_and4_1 _2499_ (.A(net178),
    .B(\main.demo.zic._q_qpos[10] ),
    .C(\main.demo.zic._q_qpos[9] ),
    .D(_0360_),
    .X(_0366_));
 sg13g2_nor3_1 _2500_ (.A(net592),
    .B(net179),
    .C(_0366_),
    .Y(_0069_));
 sg13g2_o21ai_1 _2501_ (.B1(net609),
    .Y(_0367_),
    .A1(net327),
    .A2(_0366_));
 sg13g2_a21oi_1 _2502_ (.A1(net327),
    .A2(_0366_),
    .Y(_0070_),
    .B1(_0367_));
 sg13g2_nor2_1 _2503_ (.A(net171),
    .B(_0298_),
    .Y(_0368_));
 sg13g2_nor2_1 _2504_ (.A(\main.demo.zic._q_rythm_count[10] ),
    .B(\main.demo.zic._q_rythm_count[9] ),
    .Y(_0369_));
 sg13g2_and4_1 _2505_ (.A(net186),
    .B(net253),
    .C(net273),
    .D(_0369_),
    .X(_0370_));
 sg13g2_or2_1 _2506_ (.X(_0371_),
    .B(net461),
    .A(_0016_));
 sg13g2_nor2_1 _2507_ (.A(\main.demo.zic._q_rythm_count[0] ),
    .B(_0297_),
    .Y(_0372_));
 sg13g2_nor3_1 _2508_ (.A(_0368_),
    .B(net459),
    .C(_0372_),
    .Y(_0071_));
 sg13g2_a21oi_1 _2509_ (.A1(\main.demo.zic._q_rythm_count[0] ),
    .A2(net463),
    .Y(_0373_),
    .B1(net213));
 sg13g2_and3_1 _2510_ (.X(_0374_),
    .A(net213),
    .B(\main.demo.zic._q_rythm_count[0] ),
    .C(net463));
 sg13g2_nor3_1 _2511_ (.A(net459),
    .B(net214),
    .C(_0374_),
    .Y(_0072_));
 sg13g2_nor2_1 _2512_ (.A(net266),
    .B(_0374_),
    .Y(_0375_));
 sg13g2_and4_1 _2513_ (.A(net266),
    .B(net213),
    .C(\main.demo.zic._q_rythm_count[0] ),
    .D(net463),
    .X(_0376_));
 sg13g2_nor3_1 _2514_ (.A(net459),
    .B(net267),
    .C(_0376_),
    .Y(_0073_));
 sg13g2_nor2_1 _2515_ (.A(net260),
    .B(_0376_),
    .Y(_0377_));
 sg13g2_and3_1 _2516_ (.X(_0378_),
    .A(net260),
    .B(net266),
    .C(_0374_));
 sg13g2_nor3_1 _2517_ (.A(net459),
    .B(net261),
    .C(_0378_),
    .Y(_0074_));
 sg13g2_nor2_1 _2518_ (.A(net304),
    .B(_0378_),
    .Y(_0379_));
 sg13g2_and2_1 _2519_ (.A(net304),
    .B(_0378_),
    .X(_0380_));
 sg13g2_nor3_1 _2520_ (.A(net459),
    .B(_0379_),
    .C(_0380_),
    .Y(_0075_));
 sg13g2_nor2_1 _2521_ (.A(net269),
    .B(_0380_),
    .Y(_0381_));
 sg13g2_and4_1 _2522_ (.A(net269),
    .B(\main.demo.zic._q_rythm_count[4] ),
    .C(net260),
    .D(_0376_),
    .X(_0382_));
 sg13g2_nor3_1 _2523_ (.A(net459),
    .B(net270),
    .C(_0382_),
    .Y(_0076_));
 sg13g2_xnor2_1 _2524_ (.Y(_0383_),
    .A(net295),
    .B(_0382_));
 sg13g2_nor2_1 _2525_ (.A(net460),
    .B(net296),
    .Y(_0077_));
 sg13g2_a21oi_1 _2526_ (.A1(\main.demo.zic._q_rythm_count[6] ),
    .A2(_0382_),
    .Y(_0384_),
    .B1(net204));
 sg13g2_and4_1 _2527_ (.A(net204),
    .B(\main.demo.zic._q_rythm_count[6] ),
    .C(net269),
    .D(_0380_),
    .X(_0385_));
 sg13g2_nor3_1 _2528_ (.A(net459),
    .B(net205),
    .C(_0385_),
    .Y(_0078_));
 sg13g2_nor2_1 _2529_ (.A(net273),
    .B(_0385_),
    .Y(_0386_));
 sg13g2_and4_1 _2530_ (.A(net273),
    .B(net204),
    .C(\main.demo.zic._q_rythm_count[6] ),
    .D(_0382_),
    .X(_0387_));
 sg13g2_nor3_1 _2531_ (.A(net460),
    .B(net274),
    .C(_0387_),
    .Y(_0079_));
 sg13g2_nor2_1 _2532_ (.A(net276),
    .B(_0387_),
    .Y(_0388_));
 sg13g2_and2_1 _2533_ (.A(net276),
    .B(_0387_),
    .X(_0389_));
 sg13g2_nor3_1 _2534_ (.A(net460),
    .B(net277),
    .C(_0389_),
    .Y(_0080_));
 sg13g2_nor2_1 _2535_ (.A(net263),
    .B(_0389_),
    .Y(_0390_));
 sg13g2_and4_2 _2536_ (.A(net263),
    .B(\main.demo.zic._q_rythm_count[9] ),
    .C(\main.demo.zic._q_rythm_count[8] ),
    .D(_0385_),
    .X(_0391_));
 sg13g2_nor3_1 _2537_ (.A(net460),
    .B(net264),
    .C(_0391_),
    .Y(_0081_));
 sg13g2_nor2_1 _2538_ (.A(net253),
    .B(_0391_),
    .Y(_0392_));
 sg13g2_a21oi_1 _2539_ (.A1(net253),
    .A2(_0391_),
    .Y(_0393_),
    .B1(net460));
 sg13g2_nor2b_1 _2540_ (.A(net254),
    .B_N(_0393_),
    .Y(_0082_));
 sg13g2_a21oi_1 _2541_ (.A1(\main.demo.zic._q_rythm_count[11] ),
    .A2(_0391_),
    .Y(_0394_),
    .B1(net186));
 sg13g2_and3_1 _2542_ (.X(_0395_),
    .A(net186),
    .B(\main.demo.zic._q_rythm_count[11] ),
    .C(_0391_));
 sg13g2_nor3_1 _2543_ (.A(net459),
    .B(net187),
    .C(_0395_),
    .Y(_0083_));
 sg13g2_xnor2_1 _2544_ (.Y(_0396_),
    .A(net379),
    .B(_0370_));
 sg13g2_nor2_1 _2545_ (.A(net593),
    .B(net380),
    .Y(_0084_));
 sg13g2_nor2_1 _2546_ (.A(net168),
    .B(net461),
    .Y(_0397_));
 sg13g2_a21oi_1 _2547_ (.A1(_0302_),
    .A2(net461),
    .Y(_0398_),
    .B1(_0397_));
 sg13g2_nor2_1 _2548_ (.A(net593),
    .B(_0398_),
    .Y(_0085_));
 sg13g2_nand2b_1 _2549_ (.Y(_0399_),
    .B(net461),
    .A_N(_0303_));
 sg13g2_nor2_1 _2550_ (.A(net195),
    .B(_0399_),
    .Y(_0400_));
 sg13g2_and2_1 _2551_ (.A(net195),
    .B(_0399_),
    .X(_0401_));
 sg13g2_nor3_1 _2552_ (.A(net594),
    .B(_0400_),
    .C(_0401_),
    .Y(_0086_));
 sg13g2_xor2_1 _2553_ (.B(_0400_),
    .A(net210),
    .X(_0402_));
 sg13g2_nor2_1 _2554_ (.A(net592),
    .B(_0402_),
    .Y(_0087_));
 sg13g2_nor2_1 _2555_ (.A(_0310_),
    .B(_0399_),
    .Y(_0403_));
 sg13g2_xnor2_1 _2556_ (.Y(_0404_),
    .A(_0603_),
    .B(_0403_));
 sg13g2_nor2_1 _2557_ (.A(net592),
    .B(net384),
    .Y(_0088_));
 sg13g2_and2_1 _2558_ (.A(net211),
    .B(_0632_),
    .X(_0089_));
 sg13g2_and2_1 _2559_ (.A(net308),
    .B(_0632_),
    .X(_0090_));
 sg13g2_nor4_1 _2560_ (.A(_0012_),
    .B(_0400_),
    .C(_0401_),
    .D(_0404_),
    .Y(_0405_));
 sg13g2_nand2b_2 _2561_ (.Y(_0406_),
    .B(net461),
    .A_N(_0405_));
 sg13g2_nor4_1 _2562_ (.A(\main.demo.zic._q_rythm_count[7] ),
    .B(\main.demo.zic._q_rythm_count[6] ),
    .C(\main.demo.zic._q_rythm_count[5] ),
    .D(\main.demo.zic._q_rythm_count[4] ),
    .Y(_0407_));
 sg13g2_nor4_1 _2563_ (.A(\main.demo.zic._q_rythm_count[3] ),
    .B(\main.demo.zic._q_rythm_count[2] ),
    .C(\main.demo.zic._q_rythm_count[1] ),
    .D(\main.demo.zic._q_rythm_count[0] ),
    .Y(_0408_));
 sg13g2_and3_1 _2564_ (.X(_0409_),
    .A(net463),
    .B(_0407_),
    .C(_0408_));
 sg13g2_nor2_2 _2565_ (.A(net461),
    .B(_0409_),
    .Y(_0410_));
 sg13g2_or2_1 _2566_ (.X(_0411_),
    .B(_0409_),
    .A(net461));
 sg13g2_nor2_1 _2567_ (.A(\main.demo.zic._q_squ_env[1] ),
    .B(\main.demo.zic._q_squ_env[0] ),
    .Y(_0412_));
 sg13g2_nor4_2 _2568_ (.A(\main.demo.zic._q_squ_env[3] ),
    .B(net283),
    .C(\main.demo.zic._q_squ_env[1] ),
    .Y(_0413_),
    .D(\main.demo.zic._q_squ_env[0] ));
 sg13g2_nor2b_1 _2569_ (.A(\main.demo.zic._q_squ_env[4] ),
    .B_N(_0413_),
    .Y(_0414_));
 sg13g2_a21oi_2 _2570_ (.B1(net461),
    .Y(_0415_),
    .A2(_0414_),
    .A1(_0593_));
 sg13g2_a21oi_1 _2571_ (.A1(_0594_),
    .A2(_0415_),
    .Y(_0416_),
    .B1(_0410_));
 sg13g2_a221oi_1 _2572_ (.B2(_0406_),
    .C1(net594),
    .B1(_0416_),
    .A1(_0594_),
    .Y(_0091_),
    .A2(_0410_));
 sg13g2_xnor2_1 _2573_ (.Y(_0417_),
    .A(\main.demo.zic._q_squ_env[1] ),
    .B(net318));
 sg13g2_a21oi_1 _2574_ (.A1(_0415_),
    .A2(_0417_),
    .Y(_0418_),
    .B1(_0410_));
 sg13g2_o21ai_1 _2575_ (.B1(net611),
    .Y(_0419_),
    .A1(net347),
    .A2(_0411_));
 sg13g2_a21oi_1 _2576_ (.A1(_0406_),
    .A2(_0418_),
    .Y(_0092_),
    .B1(_0419_));
 sg13g2_xnor2_1 _2577_ (.Y(_0420_),
    .A(_0000_),
    .B(_0412_));
 sg13g2_and2_1 _2578_ (.A(_0409_),
    .B(_0415_),
    .X(_0421_));
 sg13g2_a22oi_1 _2579_ (.Y(_0422_),
    .B1(_0420_),
    .B2(_0421_),
    .A2(_0410_),
    .A1(net283));
 sg13g2_a21oi_1 _2580_ (.A1(_0406_),
    .A2(net284),
    .Y(_0093_),
    .B1(net594));
 sg13g2_nand3_1 _2581_ (.B(_0411_),
    .C(_0412_),
    .A(net385),
    .Y(_0423_));
 sg13g2_xnor2_1 _2582_ (.Y(_0424_),
    .A(\main.demo.zic._q_squ_env[3] ),
    .B(_0423_));
 sg13g2_o21ai_1 _2583_ (.B1(net386),
    .Y(_0425_),
    .A1(_0410_),
    .A2(_0415_));
 sg13g2_a21oi_1 _2584_ (.A1(_0406_),
    .A2(_0425_),
    .Y(_0094_),
    .B1(net593));
 sg13g2_xnor2_1 _2585_ (.Y(_0426_),
    .A(_0001_),
    .B(_0413_));
 sg13g2_a22oi_1 _2586_ (.Y(_0427_),
    .B1(_0421_),
    .B2(_0426_),
    .A2(_0410_),
    .A1(net354));
 sg13g2_a21oi_1 _2587_ (.A1(_0406_),
    .A2(net355),
    .Y(_0095_),
    .B1(net593));
 sg13g2_xnor2_1 _2588_ (.Y(_0428_),
    .A(_0002_),
    .B(_0414_));
 sg13g2_a21oi_1 _2589_ (.A1(_0415_),
    .A2(_0428_),
    .Y(_0429_),
    .B1(_0410_));
 sg13g2_a221oi_1 _2590_ (.B2(_0406_),
    .C1(net593),
    .B1(_0429_),
    .A1(_0593_),
    .Y(_0096_),
    .A2(_0410_));
 sg13g2_and2_1 _2591_ (.A(net610),
    .B(net165),
    .X(_0097_));
 sg13g2_and2_1 _2592_ (.A(\main.demo.zic._q_clock_count[1] ),
    .B(net357),
    .X(_0430_));
 sg13g2_nor3_1 _2593_ (.A(net592),
    .B(_0295_),
    .C(net358),
    .Y(_0098_));
 sg13g2_nor2_1 _2594_ (.A(net301),
    .B(_0430_),
    .Y(_0431_));
 sg13g2_nand2_1 _2595_ (.Y(_0432_),
    .A(net301),
    .B(_0430_));
 sg13g2_nand2_1 _2596_ (.Y(_0433_),
    .A(net610),
    .B(_0432_));
 sg13g2_nor2_1 _2597_ (.A(net302),
    .B(_0433_),
    .Y(_0099_));
 sg13g2_and2_1 _2598_ (.A(_0604_),
    .B(_0432_),
    .X(_0434_));
 sg13g2_nor2_1 _2599_ (.A(_0604_),
    .B(_0432_),
    .Y(_0435_));
 sg13g2_nor3_1 _2600_ (.A(net592),
    .B(_0434_),
    .C(_0435_),
    .Y(_0100_));
 sg13g2_and2_1 _2601_ (.A(net322),
    .B(_0435_),
    .X(_0436_));
 sg13g2_o21ai_1 _2602_ (.B1(net610),
    .Y(_0437_),
    .A1(net322),
    .A2(_0435_));
 sg13g2_nor2_1 _2603_ (.A(_0436_),
    .B(net323),
    .Y(_0101_));
 sg13g2_nor2_1 _2604_ (.A(net242),
    .B(_0436_),
    .Y(_0438_));
 sg13g2_and2_1 _2605_ (.A(net242),
    .B(_0436_),
    .X(_0439_));
 sg13g2_nor3_1 _2606_ (.A(net592),
    .B(net243),
    .C(_0439_),
    .Y(_0102_));
 sg13g2_o21ai_1 _2607_ (.B1(net610),
    .Y(_0440_),
    .A1(net181),
    .A2(_0439_));
 sg13g2_a21oi_1 _2608_ (.A1(net181),
    .A2(_0439_),
    .Y(_0103_),
    .B1(_0440_));
 sg13g2_nor2b_1 _2609_ (.A(_0006_),
    .B_N(_0439_),
    .Y(_0441_));
 sg13g2_o21ai_1 _2610_ (.B1(net610),
    .Y(_0442_),
    .A1(net199),
    .A2(_0441_));
 sg13g2_a21oi_1 _2611_ (.A1(net199),
    .A2(_0441_),
    .Y(_0104_),
    .B1(_0442_));
 sg13g2_and3_1 _2612_ (.X(_0443_),
    .A(\main.demo.zic._q_clock_count[7] ),
    .B(\main.demo.zic._q_clock_count[6] ),
    .C(_0439_));
 sg13g2_o21ai_1 _2613_ (.B1(net610),
    .Y(_0444_),
    .A1(net175),
    .A2(_0443_));
 sg13g2_a21oi_1 _2614_ (.A1(net175),
    .A2(_0443_),
    .Y(_0105_),
    .B1(_0444_));
 sg13g2_nand3b_1 _2615_ (.B(\main.demo._q_frame[0] ),
    .C(\main.demo._q_prev_vs ),
    .Y(_0445_),
    .A_N(\main._w_demo_video_vs ));
 sg13g2_nor2_1 _2616_ (.A(_0610_),
    .B(_0445_),
    .Y(_0446_));
 sg13g2_xnor2_1 _2617_ (.Y(_0447_),
    .A(net360),
    .B(_0445_));
 sg13g2_nand2_1 _2618_ (.Y(_0448_),
    .A(\main.demo._q_frame[2] ),
    .B(\main.demo._q_frame[3] ));
 sg13g2_nor3_2 _2619_ (.A(_0610_),
    .B(_0445_),
    .C(_0448_),
    .Y(_0449_));
 sg13g2_nand2_1 _2620_ (.Y(_0450_),
    .A(net315),
    .B(\main.demo._q_frame[5] ));
 sg13g2_nor4_2 _2621_ (.A(_0610_),
    .B(_0445_),
    .C(_0448_),
    .Y(_0451_),
    .D(_0450_));
 sg13g2_and2_1 _2622_ (.A(\main.demo._q_frame[6] ),
    .B(\main.demo._q_frame[7] ),
    .X(_0452_));
 sg13g2_nand3_1 _2623_ (.B(_0451_),
    .C(_0452_),
    .A(net361),
    .Y(_0453_));
 sg13g2_xor2_1 _2624_ (.B(_0453_),
    .A(_0005_),
    .X(_0454_));
 sg13g2_xor2_1 _2625_ (.B(net458),
    .A(_0447_),
    .X(_0455_));
 sg13g2_nand2_1 _2626_ (.Y(_0456_),
    .A(net567),
    .B(_0455_));
 sg13g2_xor2_1 _2627_ (.B(_0456_),
    .A(net272),
    .X(_0457_));
 sg13g2_nor2_1 _2628_ (.A(net564),
    .B(_0457_),
    .Y(_0106_));
 sg13g2_nand2_1 _2629_ (.Y(_0458_),
    .A(\main.demo._q_vT[0] ),
    .B(_0455_));
 sg13g2_xnor2_1 _2630_ (.Y(_0459_),
    .A(net369),
    .B(_0446_));
 sg13g2_xnor2_1 _2631_ (.Y(_0460_),
    .A(net458),
    .B(_0459_));
 sg13g2_nand2_1 _2632_ (.Y(_0461_),
    .A(\main.demo._q_vT[1] ),
    .B(_0460_));
 sg13g2_xnor2_1 _2633_ (.Y(_0462_),
    .A(\main.demo._q_vT[1] ),
    .B(_0460_));
 sg13g2_xor2_1 _2634_ (.B(_0462_),
    .A(_0458_),
    .X(_0463_));
 sg13g2_nor2_1 _2635_ (.A(_0244_),
    .B(_0463_),
    .Y(_0464_));
 sg13g2_nor2_1 _2636_ (.A(net249),
    .B(net567),
    .Y(_0465_));
 sg13g2_nor3_1 _2637_ (.A(net564),
    .B(_0464_),
    .C(_0465_),
    .Y(_0107_));
 sg13g2_a21o_1 _2638_ (.A2(_0446_),
    .A1(net369),
    .B1(net281),
    .X(_0466_));
 sg13g2_nand2b_1 _2639_ (.Y(_0467_),
    .B(_0466_),
    .A_N(_0449_));
 sg13g2_xor2_1 _2640_ (.B(_0467_),
    .A(net458),
    .X(_0468_));
 sg13g2_nor2_1 _2641_ (.A(_0592_),
    .B(_0468_),
    .Y(_0469_));
 sg13g2_xnor2_1 _2642_ (.Y(_0470_),
    .A(net365),
    .B(_0468_));
 sg13g2_o21ai_1 _2643_ (.B1(_0461_),
    .Y(_0471_),
    .A1(_0458_),
    .A2(_0462_));
 sg13g2_xnor2_1 _2644_ (.Y(_0472_),
    .A(_0470_),
    .B(_0471_));
 sg13g2_a21o_1 _2645_ (.A2(_0244_),
    .A1(_0592_),
    .B1(net564),
    .X(_0473_));
 sg13g2_a21oi_1 _2646_ (.A1(net567),
    .A2(_0472_),
    .Y(_0108_),
    .B1(net366));
 sg13g2_xnor2_1 _2647_ (.Y(_0474_),
    .A(net315),
    .B(_0449_));
 sg13g2_xnor2_1 _2648_ (.Y(_0475_),
    .A(_0454_),
    .B(_0474_));
 sg13g2_nand2_1 _2649_ (.Y(_0476_),
    .A(\main.demo._q_vT[3] ),
    .B(_0475_));
 sg13g2_nor2_1 _2650_ (.A(\main.demo._q_vT[3] ),
    .B(_0475_),
    .Y(_0477_));
 sg13g2_xor2_1 _2651_ (.B(_0475_),
    .A(\main.demo._q_vT[3] ),
    .X(_0478_));
 sg13g2_a21oi_1 _2652_ (.A1(_0470_),
    .A2(_0471_),
    .Y(_0479_),
    .B1(_0469_));
 sg13g2_xnor2_1 _2653_ (.Y(_0480_),
    .A(_0478_),
    .B(_0479_));
 sg13g2_nor2_1 _2654_ (.A(_0244_),
    .B(_0480_),
    .Y(_0481_));
 sg13g2_nor2_1 _2655_ (.A(net293),
    .B(net567),
    .Y(_0482_));
 sg13g2_nor3_1 _2656_ (.A(net564),
    .B(_0481_),
    .C(_0482_),
    .Y(_0109_));
 sg13g2_nor2b_1 _2657_ (.A(net344),
    .B_N(_0449_),
    .Y(_0483_));
 sg13g2_xnor2_1 _2658_ (.Y(_0484_),
    .A(\main.demo._q_frame[5] ),
    .B(_0483_));
 sg13g2_xnor2_1 _2659_ (.Y(_0485_),
    .A(net458),
    .B(_0484_));
 sg13g2_and2_1 _2660_ (.A(\main.demo._q_vT[4] ),
    .B(_0485_),
    .X(_0486_));
 sg13g2_xor2_1 _2661_ (.B(_0485_),
    .A(\main.demo._q_vT[4] ),
    .X(_0487_));
 sg13g2_o21ai_1 _2662_ (.B1(_0476_),
    .Y(_0488_),
    .A1(_0477_),
    .A2(_0479_));
 sg13g2_xor2_1 _2663_ (.B(_0488_),
    .A(_0487_),
    .X(_0489_));
 sg13g2_nor2_1 _2664_ (.A(_0244_),
    .B(_0489_),
    .Y(_0490_));
 sg13g2_nor2_1 _2665_ (.A(net294),
    .B(net566),
    .Y(_0491_));
 sg13g2_nor3_1 _2666_ (.A(net563),
    .B(_0490_),
    .C(_0491_),
    .Y(_0110_));
 sg13g2_a21oi_1 _2667_ (.A1(_0487_),
    .A2(_0488_),
    .Y(_0492_),
    .B1(_0486_));
 sg13g2_xnor2_1 _2668_ (.Y(_0493_),
    .A(net325),
    .B(_0451_));
 sg13g2_xnor2_1 _2669_ (.Y(_0494_),
    .A(net458),
    .B(_0493_));
 sg13g2_nor2_1 _2670_ (.A(\main.demo._q_vT[5] ),
    .B(_0494_),
    .Y(_0495_));
 sg13g2_xor2_1 _2671_ (.B(_0494_),
    .A(\main.demo._q_vT[5] ),
    .X(_0496_));
 sg13g2_o21ai_1 _2672_ (.B1(net566),
    .Y(_0497_),
    .A1(_0492_),
    .A2(_0496_));
 sg13g2_a21oi_1 _2673_ (.A1(_0492_),
    .A2(_0496_),
    .Y(_0498_),
    .B1(_0497_));
 sg13g2_nor2_1 _2674_ (.A(net324),
    .B(net566),
    .Y(_0499_));
 sg13g2_nor3_1 _2675_ (.A(net563),
    .B(_0498_),
    .C(_0499_),
    .Y(_0111_));
 sg13g2_nand2_1 _2676_ (.Y(_0500_),
    .A(_0612_),
    .B(_0451_));
 sg13g2_xor2_1 _2677_ (.B(_0500_),
    .A(net388),
    .X(_0501_));
 sg13g2_xnor2_1 _2678_ (.Y(_0502_),
    .A(net458),
    .B(_0501_));
 sg13g2_and2_1 _2679_ (.A(\main.demo._q_vT[6] ),
    .B(_0502_),
    .X(_0503_));
 sg13g2_xnor2_1 _2680_ (.Y(_0504_),
    .A(_0591_),
    .B(_0502_));
 sg13g2_inv_1 _2681_ (.Y(_0505_),
    .A(_0504_));
 sg13g2_a221oi_1 _2682_ (.B2(\main.demo._q_vT[5] ),
    .C1(_0486_),
    .B1(_0494_),
    .A1(_0487_),
    .Y(_0506_),
    .A2(_0488_));
 sg13g2_nor3_1 _2683_ (.A(_0495_),
    .B(_0505_),
    .C(_0506_),
    .Y(_0507_));
 sg13g2_o21ai_1 _2684_ (.B1(_0505_),
    .Y(_0508_),
    .A1(_0495_),
    .A2(_0506_));
 sg13g2_nand2b_1 _2685_ (.Y(_0509_),
    .B(_0508_),
    .A_N(_0507_));
 sg13g2_a21o_1 _2686_ (.A2(_0244_),
    .A1(_0591_),
    .B1(net563),
    .X(_0510_));
 sg13g2_a21oi_1 _2687_ (.A1(net566),
    .A2(_0509_),
    .Y(_0112_),
    .B1(net391));
 sg13g2_a21o_1 _2688_ (.A2(_0452_),
    .A1(_0451_),
    .B1(net361),
    .X(_0511_));
 sg13g2_nand2_1 _2689_ (.Y(_0512_),
    .A(_0453_),
    .B(_0511_));
 sg13g2_mux2_2 _2690_ (.A0(_0005_),
    .A1(net458),
    .S(_0512_),
    .X(_0513_));
 sg13g2_nand2_1 _2691_ (.Y(_0514_),
    .A(\main.demo._q_vT[7] ),
    .B(_0513_));
 sg13g2_xor2_1 _2692_ (.B(_0513_),
    .A(\main.demo._q_vT[7] ),
    .X(_0515_));
 sg13g2_o21ai_1 _2693_ (.B1(_0515_),
    .Y(_0516_),
    .A1(_0503_),
    .A2(_0507_));
 sg13g2_or3_1 _2694_ (.A(_0503_),
    .B(_0507_),
    .C(_0515_),
    .X(_0517_));
 sg13g2_a21o_1 _2695_ (.A2(_0517_),
    .A1(_0516_),
    .B1(_0244_),
    .X(_0518_));
 sg13g2_o21ai_1 _2696_ (.B1(_0518_),
    .Y(_0519_),
    .A1(net372),
    .A2(net566));
 sg13g2_nor2_1 _2697_ (.A(net563),
    .B(_0519_),
    .Y(_0113_));
 sg13g2_a21oi_2 _2698_ (.B1(_0244_),
    .Y(_0520_),
    .A2(_0516_),
    .A1(_0514_));
 sg13g2_xnor2_1 _2699_ (.Y(_0521_),
    .A(net352),
    .B(_0520_));
 sg13g2_nor2_1 _2700_ (.A(net563),
    .B(_0521_),
    .Y(_0114_));
 sg13g2_a21oi_1 _2701_ (.A1(net352),
    .A2(_0520_),
    .Y(_0522_),
    .B1(net371));
 sg13g2_nand3_1 _2702_ (.B(net352),
    .C(_0520_),
    .A(net371),
    .Y(_0523_));
 sg13g2_nor2_1 _2703_ (.A(net563),
    .B(_0522_),
    .Y(_0524_));
 sg13g2_and2_1 _2704_ (.A(_0523_),
    .B(_0524_),
    .X(_0115_));
 sg13g2_nor2b_1 _2705_ (.A(net257),
    .B_N(_0523_),
    .Y(_0525_));
 sg13g2_and4_1 _2706_ (.A(net257),
    .B(\main.demo._q_vT[9] ),
    .C(\main.demo._q_vT[8] ),
    .D(_0520_),
    .X(_0526_));
 sg13g2_nor3_1 _2707_ (.A(net563),
    .B(net258),
    .C(_0526_),
    .Y(_0116_));
 sg13g2_xnor2_1 _2708_ (.Y(_0527_),
    .A(net240),
    .B(_0526_));
 sg13g2_nor2_1 _2709_ (.A(net563),
    .B(net241),
    .Y(_0117_));
 sg13g2_nor3_1 _2710_ (.A(net233),
    .B(_0618_),
    .C(_0264_),
    .Y(_0118_));
 sg13g2_nand2b_2 _2711_ (.Y(_0528_),
    .B(_0621_),
    .A_N(net233));
 sg13g2_xnor2_1 _2712_ (.Y(_0529_),
    .A(net282),
    .B(_0264_));
 sg13g2_nor2_1 _2713_ (.A(_0528_),
    .B(_0529_),
    .Y(_0119_));
 sg13g2_a21oi_1 _2714_ (.A1(\main.demo.vga._q_xcount[2] ),
    .A2(_0264_),
    .Y(_0530_),
    .B1(net183));
 sg13g2_nor3_1 _2715_ (.A(_0265_),
    .B(_0528_),
    .C(net184),
    .Y(_0120_));
 sg13g2_xnor2_1 _2716_ (.Y(_0531_),
    .A(net339),
    .B(_0265_));
 sg13g2_nor2_1 _2717_ (.A(_0528_),
    .B(_0531_),
    .Y(_0121_));
 sg13g2_a21oi_1 _2718_ (.A1(\main.demo.vga._q_xcount[6] ),
    .A2(_0272_),
    .Y(_0532_),
    .B1(net220));
 sg13g2_nor3_1 _2719_ (.A(_0276_),
    .B(_0528_),
    .C(net221),
    .Y(_0122_));
 sg13g2_or2_1 _2720_ (.X(_0533_),
    .B(_0455_),
    .A(net290));
 sg13g2_and2_1 _2721_ (.A(net173),
    .B(net612),
    .X(_0534_));
 sg13g2_nand2_2 _2722_ (.Y(_0535_),
    .A(net173),
    .B(net612));
 sg13g2_nand2_1 _2723_ (.Y(_0536_),
    .A(net290),
    .B(_0455_));
 sg13g2_and3_1 _2724_ (.X(_0123_),
    .A(_0533_),
    .B(_0534_),
    .C(_0536_));
 sg13g2_nand2_1 _2725_ (.Y(_0537_),
    .A(net392),
    .B(_0460_));
 sg13g2_xnor2_1 _2726_ (.Y(_0538_),
    .A(\main.demo._q_uT[1] ),
    .B(_0460_));
 sg13g2_o21ai_1 _2727_ (.B1(_0534_),
    .Y(_0539_),
    .A1(_0536_),
    .A2(_0538_));
 sg13g2_a21oi_1 _2728_ (.A1(_0536_),
    .A2(_0538_),
    .Y(_0124_),
    .B1(_0539_));
 sg13g2_nor2_1 _2729_ (.A(_0614_),
    .B(_0468_),
    .Y(_0540_));
 sg13g2_xnor2_1 _2730_ (.Y(_0541_),
    .A(_0614_),
    .B(_0468_));
 sg13g2_inv_1 _2731_ (.Y(_0542_),
    .A(_0541_));
 sg13g2_o21ai_1 _2732_ (.B1(_0537_),
    .Y(_0543_),
    .A1(_0536_),
    .A2(_0538_));
 sg13g2_nor2_1 _2733_ (.A(_0542_),
    .B(_0543_),
    .Y(_0544_));
 sg13g2_a21oi_1 _2734_ (.A1(_0542_),
    .A2(_0543_),
    .Y(_0545_),
    .B1(_0535_));
 sg13g2_nor2b_1 _2735_ (.A(net393),
    .B_N(_0545_),
    .Y(_0125_));
 sg13g2_nand2_1 _2736_ (.Y(_0546_),
    .A(\main.demo._q_uT[3] ),
    .B(_0475_));
 sg13g2_xnor2_1 _2737_ (.Y(_0547_),
    .A(net376),
    .B(_0475_));
 sg13g2_a21oi_2 _2738_ (.B1(_0540_),
    .Y(_0548_),
    .A2(_0543_),
    .A1(_0542_));
 sg13g2_o21ai_1 _2739_ (.B1(net562),
    .Y(_0549_),
    .A1(_0547_),
    .A2(_0548_));
 sg13g2_a21oi_1 _2740_ (.A1(_0547_),
    .A2(_0548_),
    .Y(_0126_),
    .B1(_0549_));
 sg13g2_nand2_1 _2741_ (.Y(_0550_),
    .A(\main.demo._q_uT[4] ),
    .B(_0485_));
 sg13g2_inv_1 _2742_ (.Y(_0551_),
    .A(_0550_));
 sg13g2_xor2_1 _2743_ (.B(_0485_),
    .A(\main.demo._q_uT[4] ),
    .X(_0552_));
 sg13g2_o21ai_1 _2744_ (.B1(_0546_),
    .Y(_0553_),
    .A1(_0547_),
    .A2(_0548_));
 sg13g2_or2_1 _2745_ (.X(_0554_),
    .B(_0553_),
    .A(_0552_));
 sg13g2_nand2_1 _2746_ (.Y(_0555_),
    .A(_0552_),
    .B(_0553_));
 sg13g2_and3_1 _2747_ (.X(_0127_),
    .A(net562),
    .B(_0554_),
    .C(_0555_));
 sg13g2_nand2_1 _2748_ (.Y(_0556_),
    .A(_0550_),
    .B(_0555_));
 sg13g2_nor2_1 _2749_ (.A(net403),
    .B(_0494_),
    .Y(_0557_));
 sg13g2_xnor2_1 _2750_ (.Y(_0558_),
    .A(net398),
    .B(_0494_));
 sg13g2_xor2_1 _2751_ (.B(_0558_),
    .A(_0556_),
    .X(_0559_));
 sg13g2_nor2_1 _2752_ (.A(net561),
    .B(net399),
    .Y(_0128_));
 sg13g2_nand2_1 _2753_ (.Y(_0560_),
    .A(net394),
    .B(_0502_));
 sg13g2_xor2_1 _2754_ (.B(_0502_),
    .A(\main.demo._q_uT[6] ),
    .X(_0561_));
 sg13g2_inv_1 _2755_ (.Y(_0562_),
    .A(_0561_));
 sg13g2_a221oi_1 _2756_ (.B2(_0553_),
    .C1(_0551_),
    .B1(_0552_),
    .A1(\main.demo._q_uT[5] ),
    .Y(_0563_),
    .A2(_0494_));
 sg13g2_o21ai_1 _2757_ (.B1(_0562_),
    .Y(_0564_),
    .A1(_0557_),
    .A2(_0563_));
 sg13g2_or3_1 _2758_ (.A(_0557_),
    .B(_0562_),
    .C(_0563_),
    .X(_0565_));
 sg13g2_and3_1 _2759_ (.X(_0129_),
    .A(net562),
    .B(_0564_),
    .C(_0565_));
 sg13g2_nand2_1 _2760_ (.Y(_0566_),
    .A(\main.demo._q_uT[7] ),
    .B(_0513_));
 sg13g2_xor2_1 _2761_ (.B(_0513_),
    .A(\main.demo._q_uT[7] ),
    .X(_0567_));
 sg13g2_inv_1 _2762_ (.Y(_0568_),
    .A(_0567_));
 sg13g2_nand3_1 _2763_ (.B(_0565_),
    .C(_0568_),
    .A(_0560_),
    .Y(_0569_));
 sg13g2_a21o_1 _2764_ (.A2(_0565_),
    .A1(_0560_),
    .B1(_0568_),
    .X(_0570_));
 sg13g2_and3_1 _2765_ (.X(_0130_),
    .A(net562),
    .B(_0569_),
    .C(_0570_));
 sg13g2_nand2_2 _2766_ (.Y(_0571_),
    .A(_0566_),
    .B(_0570_));
 sg13g2_o21ai_1 _2767_ (.B1(net562),
    .Y(_0572_),
    .A1(net231),
    .A2(_0571_));
 sg13g2_a21oi_1 _2768_ (.A1(net231),
    .A2(_0571_),
    .Y(_0131_),
    .B1(_0572_));
 sg13g2_a21oi_1 _2769_ (.A1(\main.demo._q_uT[8] ),
    .A2(_0571_),
    .Y(_0573_),
    .B1(net207));
 sg13g2_and3_2 _2770_ (.X(_0574_),
    .A(net231),
    .B(net207),
    .C(_0571_));
 sg13g2_nor3_1 _2771_ (.A(net561),
    .B(net208),
    .C(_0574_),
    .Y(_0132_));
 sg13g2_o21ai_1 _2772_ (.B1(net562),
    .Y(_0575_),
    .A1(net292),
    .A2(_0574_));
 sg13g2_a21oi_1 _2773_ (.A1(net292),
    .A2(_0574_),
    .Y(_0133_),
    .B1(_0575_));
 sg13g2_a21oi_1 _2774_ (.A1(\main.demo._q_uT[10] ),
    .A2(_0574_),
    .Y(_0576_),
    .B1(net201));
 sg13g2_and3_1 _2775_ (.X(_0577_),
    .A(\main.demo._q_uT[10] ),
    .B(net201),
    .C(_0574_));
 sg13g2_nor3_1 _2776_ (.A(_0535_),
    .B(net202),
    .C(_0577_),
    .Y(_0134_));
 sg13g2_and2_1 _2777_ (.A(net163),
    .B(net562),
    .X(_0135_));
 sg13g2_nor2_1 _2778_ (.A(net225),
    .B(\main.demo._q_u[1] ),
    .Y(_0578_));
 sg13g2_and2_1 _2779_ (.A(net225),
    .B(\main.demo._q_u[1] ),
    .X(_0579_));
 sg13g2_nor3_1 _2780_ (.A(net561),
    .B(net226),
    .C(_0579_),
    .Y(_0136_));
 sg13g2_a21oi_1 _2781_ (.A1(net367),
    .A2(_0579_),
    .Y(_0580_),
    .B1(net561));
 sg13g2_o21ai_1 _2782_ (.B1(_0580_),
    .Y(_0581_),
    .A1(net367),
    .A2(_0579_));
 sg13g2_inv_1 _2783_ (.Y(_0137_),
    .A(net368));
 sg13g2_a21oi_1 _2784_ (.A1(\main.demo._q_u[2] ),
    .A2(_0579_),
    .Y(_0582_),
    .B1(net298));
 sg13g2_and3_1 _2785_ (.X(_0583_),
    .A(\main.demo._q_u[2] ),
    .B(net298),
    .C(_0579_));
 sg13g2_nor3_1 _2786_ (.A(net561),
    .B(net299),
    .C(_0583_),
    .Y(_0138_));
 sg13g2_and2_1 _2787_ (.A(net332),
    .B(_0583_),
    .X(_0584_));
 sg13g2_o21ai_1 _2788_ (.B1(net562),
    .Y(_0585_),
    .A1(net332),
    .A2(_0583_));
 sg13g2_nor2_1 _2789_ (.A(_0584_),
    .B(net333),
    .Y(_0139_));
 sg13g2_xnor2_1 _2790_ (.Y(_0586_),
    .A(net340),
    .B(_0584_));
 sg13g2_nor2_1 _2791_ (.A(net561),
    .B(_0586_),
    .Y(_0140_));
 sg13g2_a21oi_1 _2792_ (.A1(\main.demo._q_u[5] ),
    .A2(_0584_),
    .Y(_0587_),
    .B1(net246));
 sg13g2_and3_1 _2793_ (.X(_0588_),
    .A(\main.demo._q_u[5] ),
    .B(net246),
    .C(_0584_));
 sg13g2_nor3_1 _2794_ (.A(net561),
    .B(net247),
    .C(_0588_),
    .Y(_0141_));
 sg13g2_a21oi_1 _2795_ (.A1(net311),
    .A2(_0588_),
    .Y(_0589_),
    .B1(net561));
 sg13g2_o21ai_1 _2796_ (.B1(_0589_),
    .Y(_0590_),
    .A1(net311),
    .A2(_0588_));
 sg13g2_inv_1 _2797_ (.Y(_0142_),
    .A(net312));
 sg13g2_and2_1 _2798_ (.A(net612),
    .B(_0447_),
    .X(_0143_));
 sg13g2_nor2_1 _2799_ (.A(net596),
    .B(net370),
    .Y(_0144_));
 sg13g2_nor2_1 _2800_ (.A(net596),
    .B(_0467_),
    .Y(_0145_));
 sg13g2_nor2_1 _2801_ (.A(net596),
    .B(net316),
    .Y(_0146_));
 sg13g2_nor2_1 _2802_ (.A(net596),
    .B(net345),
    .Y(_0147_));
 sg13g2_nor2_1 _2803_ (.A(net593),
    .B(net326),
    .Y(_0148_));
 sg13g2_nor2_1 _2804_ (.A(net593),
    .B(net389),
    .Y(_0149_));
 sg13g2_nor2_1 _2805_ (.A(net593),
    .B(_0512_),
    .Y(_0150_));
 sg13g2_and2_1 _2806_ (.A(net611),
    .B(net458),
    .X(_0151_));
 sg13g2_dfrbp_1 _2807_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net34),
    .D(net170),
    .Q_N(_0020_),
    .Q(\main.demo._q_frame[0] ));
 sg13g2_dfrbp_1 _2808_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net46),
    .D(_0022_),
    .Q_N(_1383_),
    .Q(uo_out[0]));
 sg13g2_dfrbp_1 _2809_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net45),
    .D(_0023_),
    .Q_N(_1382_),
    .Q(uo_out[1]));
 sg13g2_dfrbp_1 _2810_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net44),
    .D(_0024_),
    .Q_N(_1381_),
    .Q(uo_out[2]));
 sg13g2_dfrbp_1 _2811_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net43),
    .D(_0025_),
    .Q_N(_1380_),
    .Q(uo_out[4]));
 sg13g2_dfrbp_1 _2812_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net42),
    .D(_0026_),
    .Q_N(_1379_),
    .Q(uo_out[5]));
 sg13g2_dfrbp_1 _2813_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net41),
    .D(_0027_),
    .Q_N(_1378_),
    .Q(uo_out[6]));
 sg13g2_dfrbp_1 _2814_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net40),
    .D(net351),
    .Q_N(_1377_),
    .Q(\main.demo.vga._d_vblank ));
 sg13g2_dfrbp_1 _2815_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net38),
    .D(net167),
    .Q_N(_0019_),
    .Q(\main.demo._q_v[0] ));
 sg13g2_dfrbp_1 _2816_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net36),
    .D(net198),
    .Q_N(_1376_),
    .Q(\main.demo._q_v[1] ));
 sg13g2_dfrbp_1 _2817_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net33),
    .D(_0031_),
    .Q_N(_1375_),
    .Q(\main.demo._q_v[2] ));
 sg13g2_dfrbp_1 _2818_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net31),
    .D(_0032_),
    .Q_N(_1374_),
    .Q(\main.demo._q_v[3] ));
 sg13g2_dfrbp_1 _2819_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net29),
    .D(_0033_),
    .Q_N(_1373_),
    .Q(\main.demo._q_v[4] ));
 sg13g2_dfrbp_1 _2820_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net27),
    .D(_0034_),
    .Q_N(_1372_),
    .Q(\main.demo._q_v[5] ));
 sg13g2_dfrbp_1 _2821_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net25),
    .D(net236),
    .Q_N(_1371_),
    .Q(\main.demo._q_v[6] ));
 sg13g2_dfrbp_1 _2822_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net23),
    .D(_0036_),
    .Q_N(_1370_),
    .Q(\main.demo._t___block_1_p4[0] ));
 sg13g2_dfrbp_1 _2823_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net22),
    .D(net194),
    .Q_N(_1369_),
    .Q(\main.demo._t___block_1_p4[1] ));
 sg13g2_dfrbp_1 _2824_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net93),
    .D(_0038_),
    .Q_N(_1384_),
    .Q(\main.demo.vga._q_active_v ));
 sg13g2_dfrbp_1 _2825_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net21),
    .D(\main.demo.vga._d_active ),
    .Q_N(_1368_),
    .Q(\main.demo._w_vga_active ));
 sg13g2_dfrbp_1 _2826_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net20),
    .D(net212),
    .Q_N(_1367_),
    .Q(\main._w_demo_video_vs ));
 sg13g2_dfrbp_1 _2827_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net18),
    .D(net338),
    .Q_N(_1366_),
    .Q(\main._w_demo_video_hs ));
 sg13g2_dfrbp_1 _2828_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net16),
    .D(_0041_),
    .Q_N(_1365_),
    .Q(\main.demo.vga._q_active_h ));
 sg13g2_dfrbp_1 _2829_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net158),
    .D(_0042_),
    .Q_N(_1364_),
    .Q(\main.demo.vga._q_xcount[0] ));
 sg13g2_dfrbp_1 _2830_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net157),
    .D(_0043_),
    .Q_N(_1363_),
    .Q(\main.demo.vga._q_xcount[5] ));
 sg13g2_dfrbp_1 _2831_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net156),
    .D(_0044_),
    .Q_N(_1362_),
    .Q(\main.demo.vga._q_xcount[6] ));
 sg13g2_dfrbp_1 _2832_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net155),
    .D(_0045_),
    .Q_N(_1361_),
    .Q(\main.demo.vga._q_xcount[8] ));
 sg13g2_dfrbp_1 _2833_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net154),
    .D(net239),
    .Q_N(_1360_),
    .Q(\main.demo.vga._q_xcount[9] ));
 sg13g2_dfrbp_1 _2834_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net153),
    .D(_0047_),
    .Q_N(_1359_),
    .Q(\main.demo.vga._q_xcount[10] ));
 sg13g2_dfrbp_1 _2835_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net152),
    .D(net335),
    .Q_N(_1358_),
    .Q(\main.demo.vga._q_ycount[0] ));
 sg13g2_dfrbp_1 _2836_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net150),
    .D(_0049_),
    .Q_N(_1357_),
    .Q(\main.demo.vga._q_ycount[1] ));
 sg13g2_dfrbp_1 _2837_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net148),
    .D(net375),
    .Q_N(_1356_),
    .Q(\main.demo.vga._q_ycount[2] ));
 sg13g2_dfrbp_1 _2838_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net146),
    .D(net252),
    .Q_N(_1355_),
    .Q(\main.demo.vga._q_ycount[3] ));
 sg13g2_dfrbp_1 _2839_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net144),
    .D(net396),
    .Q_N(_1354_),
    .Q(\main.demo.vga._q_ycount[4] ));
 sg13g2_dfrbp_1 _2840_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net142),
    .D(net331),
    .Q_N(_1353_),
    .Q(\main.demo.vga._q_ycount[5] ));
 sg13g2_dfrbp_1 _2841_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net140),
    .D(_0054_),
    .Q_N(_1352_),
    .Q(\main.demo.vga._q_ycount[6] ));
 sg13g2_dfrbp_1 _2842_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net138),
    .D(_0055_),
    .Q_N(_1351_),
    .Q(\main.demo.vga._q_ycount[7] ));
 sg13g2_dfrbp_1 _2843_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net136),
    .D(_0056_),
    .Q_N(_1350_),
    .Q(\main.demo.vga._q_ycount[8] ));
 sg13g2_dfrbp_1 _2844_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net134),
    .D(_0057_),
    .Q_N(_1349_),
    .Q(\main.demo._q_v[7] ));
 sg13g2_dfrbp_1 _2845_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net132),
    .D(_0058_),
    .Q_N(_1348_),
    .Q(\main.demo.zic._q_qpos[0] ));
 sg13g2_dfrbp_1 _2846_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net130),
    .D(net217),
    .Q_N(_0009_),
    .Q(\main.demo.zic._q_qpos[1] ));
 sg13g2_dfrbp_1 _2847_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net128),
    .D(_0060_),
    .Q_N(_1347_),
    .Q(\main.demo.zic._q_qpos[2] ));
 sg13g2_dfrbp_1 _2848_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net126),
    .D(net219),
    .Q_N(_0010_),
    .Q(\main.demo.zic._q_qpos[3] ));
 sg13g2_dfrbp_1 _2849_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net124),
    .D(net310),
    .Q_N(_1346_),
    .Q(\main.demo.zic._q_qpos[4] ));
 sg13g2_dfrbp_1 _2850_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net122),
    .D(net230),
    .Q_N(_0011_),
    .Q(\main.demo.zic._q_qpos[5] ));
 sg13g2_dfrbp_1 _2851_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net120),
    .D(net321),
    .Q_N(_1345_),
    .Q(\main.demo.zic._q_qpos[6] ));
 sg13g2_dfrbp_1 _2852_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net118),
    .D(net191),
    .Q_N(_1344_),
    .Q(\main.demo.zic._q_qpos[7] ));
 sg13g2_dfrbp_1 _2853_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net116),
    .D(net289),
    .Q_N(_1343_),
    .Q(\main.demo.zic._q_qpos[8] ));
 sg13g2_dfrbp_1 _2854_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net114),
    .D(_0067_),
    .Q_N(_1342_),
    .Q(\main.demo.zic._q_qpos[9] ));
 sg13g2_dfrbp_1 _2855_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net102),
    .D(net343),
    .Q_N(_1341_),
    .Q(\main.demo.zic._q_qpos[10] ));
 sg13g2_dfrbp_1 _2856_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net100),
    .D(net180),
    .Q_N(_1340_),
    .Q(\main.demo.zic._q_qpos[11] ));
 sg13g2_dfrbp_1 _2857_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net98),
    .D(net328),
    .Q_N(_1339_),
    .Q(\main.demo.zic._q_qpos[12] ));
 sg13g2_dfrbp_1 _2858_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net96),
    .D(net172),
    .Q_N(_0018_),
    .Q(\main.demo.zic._q_rythm_count[0] ));
 sg13g2_dfrbp_1 _2859_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net94),
    .D(net215),
    .Q_N(_1338_),
    .Q(\main.demo.zic._q_rythm_count[1] ));
 sg13g2_dfrbp_1 _2860_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net91),
    .D(net268),
    .Q_N(_1337_),
    .Q(\main.demo.zic._q_rythm_count[2] ));
 sg13g2_dfrbp_1 _2861_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net89),
    .D(net262),
    .Q_N(_1336_),
    .Q(\main.demo.zic._q_rythm_count[3] ));
 sg13g2_dfrbp_1 _2862_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net87),
    .D(_0075_),
    .Q_N(_1335_),
    .Q(\main.demo.zic._q_rythm_count[4] ));
 sg13g2_dfrbp_1 _2863_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net85),
    .D(net271),
    .Q_N(_1334_),
    .Q(\main.demo.zic._q_rythm_count[5] ));
 sg13g2_dfrbp_1 _2864_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net83),
    .D(net297),
    .Q_N(_1333_),
    .Q(\main.demo.zic._q_rythm_count[6] ));
 sg13g2_dfrbp_1 _2865_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net81),
    .D(net206),
    .Q_N(_1332_),
    .Q(\main.demo.zic._q_rythm_count[7] ));
 sg13g2_dfrbp_1 _2866_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net79),
    .D(net275),
    .Q_N(_1331_),
    .Q(\main.demo.zic._q_rythm_count[8] ));
 sg13g2_dfrbp_1 _2867_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net77),
    .D(net278),
    .Q_N(_1330_),
    .Q(\main.demo.zic._q_rythm_count[9] ));
 sg13g2_dfrbp_1 _2868_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net75),
    .D(net265),
    .Q_N(_1329_),
    .Q(\main.demo.zic._q_rythm_count[10] ));
 sg13g2_dfrbp_1 _2869_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net73),
    .D(_0082_),
    .Q_N(_1328_),
    .Q(\main.demo.zic._q_rythm_count[11] ));
 sg13g2_dfrbp_1 _2870_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net71),
    .D(net188),
    .Q_N(_1327_),
    .Q(\main.demo.zic._q_rythm_count[12] ));
 sg13g2_dfrbp_1 _2871_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net69),
    .D(_0084_),
    .Q_N(_1326_),
    .Q(\main.demo.zic._q_idx[0] ));
 sg13g2_dfrbp_1 _2872_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net68),
    .D(_0085_),
    .Q_N(_0014_),
    .Q(\main.demo.zic._q_idx[1] ));
 sg13g2_dfrbp_1 _2873_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net67),
    .D(_0086_),
    .Q_N(_0013_),
    .Q(\main.demo.zic._q_idx[2] ));
 sg13g2_dfrbp_1 _2874_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net66),
    .D(_0087_),
    .Q_N(_0012_),
    .Q(\main.demo.zic._q_idx[3] ));
 sg13g2_dfrbp_1 _2875_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net65),
    .D(_0088_),
    .Q_N(_0015_),
    .Q(\main.demo.zic._q_idx[4] ));
 sg13g2_dfrbp_1 _2876_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net64),
    .D(_0089_),
    .Q_N(_1325_),
    .Q(\main.demo._t___block_1_p4[2] ));
 sg13g2_dfrbp_1 _2877_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net63),
    .D(_0090_),
    .Q_N(_1324_),
    .Q(\main.demo._t___block_1_p4[3] ));
 sg13g2_dfrbp_1 _2878_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net62),
    .D(_0091_),
    .Q_N(_1323_),
    .Q(\main.demo.zic._q_squ_env[0] ));
 sg13g2_dfrbp_1 _2879_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net60),
    .D(net348),
    .Q_N(_1322_),
    .Q(\main.demo.zic._q_squ_env[1] ));
 sg13g2_dfrbp_1 _2880_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net58),
    .D(net285),
    .Q_N(_0000_),
    .Q(\main.demo.zic._q_squ_env[2] ));
 sg13g2_dfrbp_1 _2881_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net56),
    .D(net387),
    .Q_N(_1321_),
    .Q(\main.demo.zic._q_squ_env[3] ));
 sg13g2_dfrbp_1 _2882_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net54),
    .D(net356),
    .Q_N(_0001_),
    .Q(\main.demo.zic._q_squ_env[4] ));
 sg13g2_dfrbp_1 _2883_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net103),
    .D(net306),
    .Q_N(_0002_),
    .Q(\main.demo.zic._q_squ_env[5] ));
 sg13g2_dfrbp_1 _2884_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net52),
    .D(net1),
    .Q_N(_0016_),
    .Q(rst_n_q));
 sg13g2_dfrbp_1 _2885_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net50),
    .D(_0097_),
    .Q_N(\main.demo.zic._d_clock_count[0] ),
    .Q(\main.demo.zic._q_clock_count[0] ));
 sg13g2_dfrbp_1 _2886_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net49),
    .D(net359),
    .Q_N(_1320_),
    .Q(\main.demo.zic._q_clock_count[1] ));
 sg13g2_dfrbp_1 _2887_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net48),
    .D(_0099_),
    .Q_N(_1319_),
    .Q(\main.demo.zic._q_clock_count[2] ));
 sg13g2_dfrbp_1 _2888_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net47),
    .D(_0100_),
    .Q_N(_0008_),
    .Q(\main.demo.zic._q_clock_count[3] ));
 sg13g2_dfrbp_1 _2889_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net39),
    .D(_0101_),
    .Q_N(_1318_),
    .Q(\main.demo.zic._q_clock_count[4] ));
 sg13g2_dfrbp_1 _2890_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net37),
    .D(_0102_),
    .Q_N(_0007_),
    .Q(\main.demo.zic._q_clock_count[5] ));
 sg13g2_dfrbp_1 _2891_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net35),
    .D(net182),
    .Q_N(_0006_),
    .Q(\main.demo.zic._q_clock_count[6] ));
 sg13g2_dfrbp_1 _2892_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net32),
    .D(net200),
    .Q_N(_1317_),
    .Q(\main.demo.zic._q_clock_count[7] ));
 sg13g2_dfrbp_1 _2893_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net104),
    .D(net176),
    .Q_N(_1385_),
    .Q(\main.demo.zic._q_clock_count[8] ));
 sg13g2_dfrbp_1 _2894_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net105),
    .D(\main.demo._d_addr[0] ),
    .Q_N(_1386_),
    .Q(\main.demo._q_addr[0] ));
 sg13g2_dfrbp_1 _2895_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net106),
    .D(\main.demo._d_addr[1] ),
    .Q_N(_1387_),
    .Q(\main.demo._q_addr[1] ));
 sg13g2_dfrbp_1 _2896_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net107),
    .D(\main.demo._d_addr[2] ),
    .Q_N(_1388_),
    .Q(\main.demo._q_addr[2] ));
 sg13g2_dfrbp_1 _2897_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net108),
    .D(\main.demo._d_addr[3] ),
    .Q_N(_1389_),
    .Q(\main.demo._q_addr[3] ));
 sg13g2_dfrbp_1 _2898_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net109),
    .D(\main.demo._d_addr[4] ),
    .Q_N(_1390_),
    .Q(\main.demo._q_addr[4] ));
 sg13g2_dfrbp_1 _2899_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net110),
    .D(\main.demo._d_addr[5] ),
    .Q_N(_1391_),
    .Q(\main.demo._q_addr[5] ));
 sg13g2_dfrbp_1 _2900_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net111),
    .D(\main.demo._d_addr[6] ),
    .Q_N(_1392_),
    .Q(\main.demo._q_addr[6] ));
 sg13g2_dfrbp_1 _2901_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net112),
    .D(\main.demo._d_addr[7] ),
    .Q_N(_1393_),
    .Q(\main.demo._q_addr[7] ));
 sg13g2_dfrbp_1 _2902_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net159),
    .D(\main.demo._d_addr[8] ),
    .Q_N(_1394_),
    .Q(\main.demo._q_addr[8] ));
 sg13g2_dfrbp_1 _2903_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net30),
    .D(\main.demo._d_addr[9] ),
    .Q_N(_1316_),
    .Q(\main.demo._q_addr[9] ));
 sg13g2_dfrbp_1 _2904_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net28),
    .D(_0106_),
    .Q_N(_1315_),
    .Q(\main.demo._q_vT[0] ));
 sg13g2_dfrbp_1 _2905_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net24),
    .D(net250),
    .Q_N(_1314_),
    .Q(\main.demo._q_vT[1] ));
 sg13g2_dfrbp_1 _2906_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net17),
    .D(_0108_),
    .Q_N(_1313_),
    .Q(\main.demo._q_vT[2] ));
 sg13g2_dfrbp_1 _2907_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net149),
    .D(_0109_),
    .Q_N(_1312_),
    .Q(\main.demo._q_vT[3] ));
 sg13g2_dfrbp_1 _2908_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net145),
    .D(_0110_),
    .Q_N(_1311_),
    .Q(\main.demo._q_vT[4] ));
 sg13g2_dfrbp_1 _2909_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net141),
    .D(_0111_),
    .Q_N(_1310_),
    .Q(\main.demo._q_vT[5] ));
 sg13g2_dfrbp_1 _2910_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net137),
    .D(_0112_),
    .Q_N(_1309_),
    .Q(\main.demo._q_vT[6] ));
 sg13g2_dfrbp_1 _2911_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net133),
    .D(_0113_),
    .Q_N(_1308_),
    .Q(\main.demo._q_vT[7] ));
 sg13g2_dfrbp_1 _2912_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net129),
    .D(_0114_),
    .Q_N(_1307_),
    .Q(\main.demo._q_vT[8] ));
 sg13g2_dfrbp_1 _2913_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net125),
    .D(_0115_),
    .Q_N(_1306_),
    .Q(\main.demo._q_vT[9] ));
 sg13g2_dfrbp_1 _2914_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net121),
    .D(net259),
    .Q_N(_1305_),
    .Q(\main.demo._q_vT[10] ));
 sg13g2_dfrbp_1 _2915_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net117),
    .D(_0117_),
    .Q_N(_1304_),
    .Q(\main.demo._q_vT[11] ));
 sg13g2_dfrbp_1 _2916_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net113),
    .D(_0118_),
    .Q_N(_1303_),
    .Q(\main.demo.vga._q_xcount[1] ));
 sg13g2_dfrbp_1 _2917_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net101),
    .D(_0119_),
    .Q_N(_1302_),
    .Q(\main.demo.vga._q_xcount[2] ));
 sg13g2_dfrbp_1 _2918_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net99),
    .D(net185),
    .Q_N(_1301_),
    .Q(\main.demo.vga._q_xcount[3] ));
 sg13g2_dfrbp_1 _2919_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net97),
    .D(_0121_),
    .Q_N(_1300_),
    .Q(\main.demo.vga._q_xcount[4] ));
 sg13g2_dfrbp_1 _2920_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net95),
    .D(net222),
    .Q_N(_1299_),
    .Q(\main.demo.vga._q_xcount[7] ));
 sg13g2_dfrbp_1 _2921_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net92),
    .D(_0123_),
    .Q_N(_1298_),
    .Q(\main.demo._q_uT[0] ));
 sg13g2_dfrbp_1 _2922_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net90),
    .D(net291),
    .Q_N(_1297_),
    .Q(\main.demo._q_uT[1] ));
 sg13g2_dfrbp_1 _2923_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net88),
    .D(_0125_),
    .Q_N(_1296_),
    .Q(\main.demo._q_uT[2] ));
 sg13g2_dfrbp_1 _2924_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net86),
    .D(net377),
    .Q_N(_1295_),
    .Q(\main.demo._q_uT[3] ));
 sg13g2_dfrbp_1 _2925_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net84),
    .D(_0127_),
    .Q_N(_1294_),
    .Q(\main.demo._q_uT[4] ));
 sg13g2_dfrbp_1 _2926_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net82),
    .D(_0128_),
    .Q_N(_1293_),
    .Q(\main.demo._q_uT[5] ));
 sg13g2_dfrbp_1 _2927_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net80),
    .D(_0129_),
    .Q_N(_1292_),
    .Q(\main.demo._q_uT[6] ));
 sg13g2_dfrbp_1 _2928_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net78),
    .D(_0130_),
    .Q_N(_1291_),
    .Q(\main.demo._q_uT[7] ));
 sg13g2_dfrbp_1 _2929_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net76),
    .D(net232),
    .Q_N(_1290_),
    .Q(\main.demo._q_uT[8] ));
 sg13g2_dfrbp_1 _2930_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net74),
    .D(net209),
    .Q_N(_1289_),
    .Q(\main.demo._q_uT[9] ));
 sg13g2_dfrbp_1 _2931_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net72),
    .D(_0133_),
    .Q_N(_1288_),
    .Q(\main.demo._q_uT[10] ));
 sg13g2_dfrbp_1 _2932_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net70),
    .D(net203),
    .Q_N(_1287_),
    .Q(\main.demo._q_uT[11] ));
 sg13g2_dfrbp_1 _2933_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net61),
    .D(_0135_),
    .Q_N(_0017_),
    .Q(\main.demo._q_u[0] ));
 sg13g2_dfrbp_1 _2934_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net59),
    .D(net227),
    .Q_N(_1286_),
    .Q(\main.demo._q_u[1] ));
 sg13g2_dfrbp_1 _2935_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net57),
    .D(_0137_),
    .Q_N(_1285_),
    .Q(\main.demo._q_u[2] ));
 sg13g2_dfrbp_1 _2936_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net55),
    .D(net300),
    .Q_N(_1284_),
    .Q(\main.demo._q_u[3] ));
 sg13g2_dfrbp_1 _2937_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net53),
    .D(_0139_),
    .Q_N(_1283_),
    .Q(\main.demo._q_u[4] ));
 sg13g2_dfrbp_1 _2938_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net51),
    .D(_0140_),
    .Q_N(_1282_),
    .Q(\main.demo._q_u[5] ));
 sg13g2_dfrbp_1 _2939_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net26),
    .D(net248),
    .Q_N(_1281_),
    .Q(\main.demo._q_u[6] ));
 sg13g2_dfrbp_1 _2940_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net19),
    .D(_0142_),
    .Q_N(_1280_),
    .Q(\main.demo._q_u[7] ));
 sg13g2_dfrbp_1 _2941_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net151),
    .D(_0143_),
    .Q_N(_1279_),
    .Q(\main.demo._q_frame[1] ));
 sg13g2_dfrbp_1 _2942_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net147),
    .D(_0144_),
    .Q_N(_1278_),
    .Q(\main.demo._q_frame[2] ));
 sg13g2_dfrbp_1 _2943_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net143),
    .D(_0145_),
    .Q_N(_1277_),
    .Q(\main.demo._q_frame[3] ));
 sg13g2_dfrbp_1 _2944_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net139),
    .D(_0146_),
    .Q_N(_0003_),
    .Q(\main.demo._q_frame[4] ));
 sg13g2_dfrbp_1 _2945_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net135),
    .D(_0147_),
    .Q_N(_1276_),
    .Q(\main.demo._q_frame[5] ));
 sg13g2_dfrbp_1 _2946_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net131),
    .D(_0148_),
    .Q_N(_0004_),
    .Q(\main.demo._q_frame[6] ));
 sg13g2_dfrbp_1 _2947_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net127),
    .D(_0149_),
    .Q_N(_1275_),
    .Q(\main.demo._q_frame[7] ));
 sg13g2_dfrbp_1 _2948_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net123),
    .D(_0150_),
    .Q_N(_1274_),
    .Q(\main.demo._q_frame[8] ));
 sg13g2_dfrbp_1 _2949_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net160),
    .D(_0151_),
    .Q_N(_0005_),
    .Q(\main.demo._q_frame[9] ));
 sg13g2_dfrbp_1 _2950_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net161),
    .D(net164),
    .Q_N(_1395_),
    .Q(\main.demo._q_prev_vs ));
 sg13g2_dfrbp_1 _2951_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net115),
    .D(net173),
    .Q_N(_1396_),
    .Q(\main.demo._q_prev_hs ));
 sg13g2_dfrbp_1 _2952_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net119),
    .D(\main._w_demo_audio1 ),
    .Q_N(_1273_),
    .Q(uio_out[7]));
 sg13g2_tiehi _2906__17 (.L_HI(net17));
 sg13g2_tiehi _2827__18 (.L_HI(net18));
 sg13g2_tiehi _2940__19 (.L_HI(net19));
 sg13g2_tiehi _2826__20 (.L_HI(net20));
 sg13g2_tiehi _2825__21 (.L_HI(net21));
 sg13g2_tiehi _2823__22 (.L_HI(net22));
 sg13g2_tiehi _2822__23 (.L_HI(net23));
 sg13g2_tiehi _2905__24 (.L_HI(net24));
 sg13g2_tiehi _2821__25 (.L_HI(net25));
 sg13g2_tiehi _2939__26 (.L_HI(net26));
 sg13g2_tiehi _2820__27 (.L_HI(net27));
 sg13g2_tiehi _2904__28 (.L_HI(net28));
 sg13g2_tiehi _2819__29 (.L_HI(net29));
 sg13g2_tiehi _2903__30 (.L_HI(net30));
 sg13g2_tiehi _2818__31 (.L_HI(net31));
 sg13g2_tiehi _2892__32 (.L_HI(net32));
 sg13g2_tiehi _2817__33 (.L_HI(net33));
 sg13g2_tiehi _2807__34 (.L_HI(net34));
 sg13g2_tiehi _2891__35 (.L_HI(net35));
 sg13g2_tiehi _2816__36 (.L_HI(net36));
 sg13g2_tiehi _2890__37 (.L_HI(net37));
 sg13g2_tiehi _2815__38 (.L_HI(net38));
 sg13g2_tiehi _2889__39 (.L_HI(net39));
 sg13g2_tiehi _2814__40 (.L_HI(net40));
 sg13g2_tiehi _2813__41 (.L_HI(net41));
 sg13g2_tiehi _2812__42 (.L_HI(net42));
 sg13g2_tiehi _2811__43 (.L_HI(net43));
 sg13g2_tiehi _2810__44 (.L_HI(net44));
 sg13g2_tiehi _2809__45 (.L_HI(net45));
 sg13g2_tiehi _2808__46 (.L_HI(net46));
 sg13g2_tiehi _2888__47 (.L_HI(net47));
 sg13g2_tiehi _2887__48 (.L_HI(net48));
 sg13g2_tiehi _2886__49 (.L_HI(net49));
 sg13g2_tiehi _2885__50 (.L_HI(net50));
 sg13g2_tiehi _2938__51 (.L_HI(net51));
 sg13g2_tiehi _2884__52 (.L_HI(net52));
 sg13g2_tiehi _2937__53 (.L_HI(net53));
 sg13g2_tiehi _2882__54 (.L_HI(net54));
 sg13g2_tiehi _2936__55 (.L_HI(net55));
 sg13g2_tiehi _2881__56 (.L_HI(net56));
 sg13g2_tiehi _2935__57 (.L_HI(net57));
 sg13g2_tiehi _2880__58 (.L_HI(net58));
 sg13g2_tiehi _2934__59 (.L_HI(net59));
 sg13g2_tiehi _2879__60 (.L_HI(net60));
 sg13g2_tiehi _2933__61 (.L_HI(net61));
 sg13g2_tiehi _2878__62 (.L_HI(net62));
 sg13g2_tiehi _2877__63 (.L_HI(net63));
 sg13g2_tiehi _2876__64 (.L_HI(net64));
 sg13g2_tiehi _2875__65 (.L_HI(net65));
 sg13g2_tiehi _2874__66 (.L_HI(net66));
 sg13g2_tiehi _2873__67 (.L_HI(net67));
 sg13g2_tiehi _2872__68 (.L_HI(net68));
 sg13g2_tiehi _2871__69 (.L_HI(net69));
 sg13g2_tiehi _2932__70 (.L_HI(net70));
 sg13g2_tiehi _2870__71 (.L_HI(net71));
 sg13g2_tiehi _2931__72 (.L_HI(net72));
 sg13g2_tiehi _2869__73 (.L_HI(net73));
 sg13g2_tiehi _2930__74 (.L_HI(net74));
 sg13g2_tiehi _2868__75 (.L_HI(net75));
 sg13g2_tiehi _2929__76 (.L_HI(net76));
 sg13g2_tiehi _2867__77 (.L_HI(net77));
 sg13g2_tiehi _2928__78 (.L_HI(net78));
 sg13g2_tiehi _2866__79 (.L_HI(net79));
 sg13g2_tiehi _2927__80 (.L_HI(net80));
 sg13g2_tiehi _2865__81 (.L_HI(net81));
 sg13g2_tiehi _2926__82 (.L_HI(net82));
 sg13g2_tiehi _2864__83 (.L_HI(net83));
 sg13g2_tiehi _2925__84 (.L_HI(net84));
 sg13g2_tiehi _2863__85 (.L_HI(net85));
 sg13g2_tiehi _2924__86 (.L_HI(net86));
 sg13g2_tiehi _2862__87 (.L_HI(net87));
 sg13g2_tiehi _2923__88 (.L_HI(net88));
 sg13g2_tiehi _2861__89 (.L_HI(net89));
 sg13g2_tiehi _2922__90 (.L_HI(net90));
 sg13g2_tiehi _2860__91 (.L_HI(net91));
 sg13g2_tiehi _2921__92 (.L_HI(net92));
 sg13g2_tiehi _2824__93 (.L_HI(net93));
 sg13g2_tiehi _2859__94 (.L_HI(net94));
 sg13g2_tiehi _2920__95 (.L_HI(net95));
 sg13g2_tiehi _2858__96 (.L_HI(net96));
 sg13g2_tiehi _2919__97 (.L_HI(net97));
 sg13g2_tiehi _2857__98 (.L_HI(net98));
 sg13g2_tiehi _2918__99 (.L_HI(net99));
 sg13g2_tiehi _2856__100 (.L_HI(net100));
 sg13g2_tiehi _2917__101 (.L_HI(net101));
 sg13g2_tiehi _2855__102 (.L_HI(net102));
 sg13g2_tiehi _2883__103 (.L_HI(net103));
 sg13g2_tiehi _2893__104 (.L_HI(net104));
 sg13g2_tiehi _2894__105 (.L_HI(net105));
 sg13g2_tiehi _2895__106 (.L_HI(net106));
 sg13g2_tiehi _2896__107 (.L_HI(net107));
 sg13g2_tiehi _2897__108 (.L_HI(net108));
 sg13g2_tiehi _2898__109 (.L_HI(net109));
 sg13g2_tiehi _2899__110 (.L_HI(net110));
 sg13g2_tiehi _2900__111 (.L_HI(net111));
 sg13g2_tiehi _2901__112 (.L_HI(net112));
 sg13g2_tiehi _2916__113 (.L_HI(net113));
 sg13g2_tiehi _2854__114 (.L_HI(net114));
 sg13g2_tiehi _2951__115 (.L_HI(net115));
 sg13g2_tiehi _2853__116 (.L_HI(net116));
 sg13g2_tiehi _2915__117 (.L_HI(net117));
 sg13g2_tiehi _2852__118 (.L_HI(net118));
 sg13g2_tiehi _2952__119 (.L_HI(net119));
 sg13g2_tiehi _2851__120 (.L_HI(net120));
 sg13g2_tiehi _2914__121 (.L_HI(net121));
 sg13g2_tiehi _2850__122 (.L_HI(net122));
 sg13g2_tiehi _2948__123 (.L_HI(net123));
 sg13g2_tiehi _2849__124 (.L_HI(net124));
 sg13g2_tiehi _2913__125 (.L_HI(net125));
 sg13g2_tiehi _2848__126 (.L_HI(net126));
 sg13g2_tiehi _2947__127 (.L_HI(net127));
 sg13g2_tiehi _2847__128 (.L_HI(net128));
 sg13g2_tiehi _2912__129 (.L_HI(net129));
 sg13g2_tiehi _2846__130 (.L_HI(net130));
 sg13g2_tiehi _2946__131 (.L_HI(net131));
 sg13g2_tiehi _2845__132 (.L_HI(net132));
 sg13g2_tiehi _2911__133 (.L_HI(net133));
 sg13g2_tiehi _2844__134 (.L_HI(net134));
 sg13g2_tiehi _2945__135 (.L_HI(net135));
 sg13g2_tiehi _2843__136 (.L_HI(net136));
 sg13g2_tiehi _2910__137 (.L_HI(net137));
 sg13g2_tiehi _2842__138 (.L_HI(net138));
 sg13g2_tiehi _2944__139 (.L_HI(net139));
 sg13g2_tiehi _2841__140 (.L_HI(net140));
 sg13g2_tiehi _2909__141 (.L_HI(net141));
 sg13g2_tiehi _2840__142 (.L_HI(net142));
 sg13g2_tiehi _2943__143 (.L_HI(net143));
 sg13g2_tiehi _2839__144 (.L_HI(net144));
 sg13g2_tiehi _2908__145 (.L_HI(net145));
 sg13g2_tiehi _2838__146 (.L_HI(net146));
 sg13g2_tiehi _2942__147 (.L_HI(net147));
 sg13g2_tiehi _2837__148 (.L_HI(net148));
 sg13g2_tiehi _2907__149 (.L_HI(net149));
 sg13g2_tiehi _2836__150 (.L_HI(net150));
 sg13g2_tiehi _2941__151 (.L_HI(net151));
 sg13g2_tiehi _2835__152 (.L_HI(net152));
 sg13g2_tiehi _2834__153 (.L_HI(net153));
 sg13g2_tiehi _2833__154 (.L_HI(net154));
 sg13g2_tiehi _2832__155 (.L_HI(net155));
 sg13g2_tiehi _2831__156 (.L_HI(net156));
 sg13g2_tiehi _2830__157 (.L_HI(net157));
 sg13g2_tiehi _2829__158 (.L_HI(net158));
 sg13g2_tiehi _2902__159 (.L_HI(net159));
 sg13g2_tiehi _2949__160 (.L_HI(net160));
 sg13g2_tiehi _2950__161 (.L_HI(net161));
 sg13g2_tiehi tt_um_whynot_162 (.L_HI(net162));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_whynot_3 (.L_LO(net3));
 sg13g2_tielo tt_um_whynot_4 (.L_LO(net4));
 sg13g2_tielo tt_um_whynot_5 (.L_LO(net5));
 sg13g2_tielo tt_um_whynot_6 (.L_LO(net6));
 sg13g2_tielo tt_um_whynot_7 (.L_LO(net7));
 sg13g2_tielo tt_um_whynot_8 (.L_LO(net8));
 sg13g2_tielo tt_um_whynot_9 (.L_LO(net9));
 sg13g2_tielo tt_um_whynot_10 (.L_LO(net10));
 sg13g2_tielo tt_um_whynot_11 (.L_LO(net11));
 sg13g2_tielo tt_um_whynot_12 (.L_LO(net12));
 sg13g2_tielo tt_um_whynot_13 (.L_LO(net13));
 sg13g2_tielo tt_um_whynot_14 (.L_LO(net14));
 sg13g2_tielo tt_um_whynot_15 (.L_LO(net15));
 sg13g2_tiehi _2828__16 (.L_HI(net16));
 sg13g2_buf_1 _3114_ (.A(\main.demo._q_prev_vs ),
    .X(uo_out[3]));
 sg13g2_buf_2 _3115_ (.A(\main.demo._q_prev_hs ),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout457 (.A(_0700_),
    .X(net457));
 sg13g2_buf_4 fanout458 (.X(net458),
    .A(_0454_));
 sg13g2_buf_2 fanout459 (.A(_0371_),
    .X(net459));
 sg13g2_buf_1 fanout460 (.A(_0371_),
    .X(net460));
 sg13g2_buf_4 fanout461 (.X(net461),
    .A(_0370_));
 sg13g2_buf_2 fanout462 (.A(net463),
    .X(net462));
 sg13g2_buf_2 fanout463 (.A(_0297_),
    .X(net463));
 sg13g2_buf_4 fanout464 (.X(net464),
    .A(net465));
 sg13g2_buf_4 fanout465 (.X(net465),
    .A(_0913_));
 sg13g2_buf_2 fanout466 (.A(net470),
    .X(net466));
 sg13g2_buf_2 fanout467 (.A(net470),
    .X(net467));
 sg13g2_buf_4 fanout468 (.X(net468),
    .A(net470));
 sg13g2_buf_1 fanout469 (.A(net470),
    .X(net469));
 sg13g2_buf_2 fanout470 (.A(_0895_),
    .X(net470));
 sg13g2_buf_2 fanout471 (.A(net472),
    .X(net471));
 sg13g2_buf_2 fanout472 (.A(net473),
    .X(net472));
 sg13g2_buf_4 fanout473 (.X(net473),
    .A(_0891_));
 sg13g2_buf_2 fanout474 (.A(net477),
    .X(net474));
 sg13g2_buf_4 fanout475 (.X(net475),
    .A(net476));
 sg13g2_buf_2 fanout476 (.A(net477),
    .X(net476));
 sg13g2_buf_4 fanout477 (.X(net477),
    .A(_0867_));
 sg13g2_buf_4 fanout478 (.X(net478),
    .A(net481));
 sg13g2_buf_2 fanout479 (.A(net480),
    .X(net479));
 sg13g2_buf_2 fanout480 (.A(net481),
    .X(net480));
 sg13g2_buf_2 fanout481 (.A(_0860_),
    .X(net481));
 sg13g2_buf_2 fanout482 (.A(net485),
    .X(net482));
 sg13g2_buf_1 fanout483 (.A(net485),
    .X(net483));
 sg13g2_buf_4 fanout484 (.X(net484),
    .A(net485));
 sg13g2_buf_4 fanout485 (.X(net485),
    .A(_0842_));
 sg13g2_buf_2 fanout486 (.A(net489),
    .X(net486));
 sg13g2_buf_2 fanout487 (.A(net488),
    .X(net487));
 sg13g2_buf_2 fanout488 (.A(net489),
    .X(net488));
 sg13g2_buf_2 fanout489 (.A(_0841_),
    .X(net489));
 sg13g2_buf_2 fanout490 (.A(net491),
    .X(net490));
 sg13g2_buf_4 fanout491 (.X(net491),
    .A(_0838_));
 sg13g2_buf_4 fanout492 (.X(net492),
    .A(_0838_));
 sg13g2_buf_4 fanout493 (.X(net493),
    .A(net497));
 sg13g2_buf_1 fanout494 (.A(net497),
    .X(net494));
 sg13g2_buf_2 fanout495 (.A(net496),
    .X(net495));
 sg13g2_buf_2 fanout496 (.A(net497),
    .X(net496));
 sg13g2_buf_2 fanout497 (.A(_0833_),
    .X(net497));
 sg13g2_buf_2 fanout498 (.A(net500),
    .X(net498));
 sg13g2_buf_2 fanout499 (.A(net500),
    .X(net499));
 sg13g2_buf_4 fanout500 (.X(net500),
    .A(_0831_));
 sg13g2_buf_4 fanout501 (.X(net501),
    .A(net503));
 sg13g2_buf_4 fanout502 (.X(net502),
    .A(net503));
 sg13g2_buf_4 fanout503 (.X(net503),
    .A(_0829_));
 sg13g2_buf_2 fanout504 (.A(net505),
    .X(net504));
 sg13g2_buf_2 fanout505 (.A(_0828_),
    .X(net505));
 sg13g2_buf_2 fanout506 (.A(_0828_),
    .X(net506));
 sg13g2_buf_2 fanout507 (.A(net508),
    .X(net507));
 sg13g2_buf_1 fanout508 (.A(net509),
    .X(net508));
 sg13g2_buf_2 fanout509 (.A(net510),
    .X(net509));
 sg13g2_buf_4 fanout510 (.X(net510),
    .A(_0825_));
 sg13g2_buf_2 fanout511 (.A(net512),
    .X(net511));
 sg13g2_buf_1 fanout512 (.A(net513),
    .X(net512));
 sg13g2_buf_4 fanout513 (.X(net513),
    .A(_0823_));
 sg13g2_buf_2 fanout514 (.A(_0822_),
    .X(net514));
 sg13g2_buf_4 fanout515 (.X(net515),
    .A(_0822_));
 sg13g2_buf_2 fanout516 (.A(net517),
    .X(net516));
 sg13g2_buf_2 fanout517 (.A(net518),
    .X(net517));
 sg13g2_buf_4 fanout518 (.X(net518),
    .A(_0820_));
 sg13g2_buf_4 fanout519 (.X(net519),
    .A(_0818_));
 sg13g2_buf_2 fanout520 (.A(net521),
    .X(net520));
 sg13g2_buf_1 fanout521 (.A(_0813_),
    .X(net521));
 sg13g2_buf_4 fanout522 (.X(net522),
    .A(_0813_));
 sg13g2_buf_2 fanout523 (.A(_0813_),
    .X(net523));
 sg13g2_buf_2 fanout524 (.A(_0809_),
    .X(net524));
 sg13g2_buf_2 fanout525 (.A(net526),
    .X(net525));
 sg13g2_buf_4 fanout526 (.X(net526),
    .A(_0809_));
 sg13g2_buf_2 fanout527 (.A(net528),
    .X(net527));
 sg13g2_buf_2 fanout528 (.A(net529),
    .X(net528));
 sg13g2_buf_4 fanout529 (.X(net529),
    .A(_0808_));
 sg13g2_buf_2 fanout530 (.A(net531),
    .X(net530));
 sg13g2_buf_2 fanout531 (.A(_0805_),
    .X(net531));
 sg13g2_buf_2 fanout532 (.A(_0805_),
    .X(net532));
 sg13g2_buf_4 fanout533 (.X(net533),
    .A(net534));
 sg13g2_buf_4 fanout534 (.X(net534),
    .A(_0801_));
 sg13g2_buf_4 fanout535 (.X(net535),
    .A(net536));
 sg13g2_buf_4 fanout536 (.X(net536),
    .A(_0796_));
 sg13g2_buf_4 fanout537 (.X(net537),
    .A(net538));
 sg13g2_buf_4 fanout538 (.X(net538),
    .A(_0790_));
 sg13g2_buf_2 fanout539 (.A(net542),
    .X(net539));
 sg13g2_buf_4 fanout540 (.X(net540),
    .A(net542));
 sg13g2_buf_2 fanout541 (.A(net542),
    .X(net541));
 sg13g2_buf_4 fanout542 (.X(net542),
    .A(_0788_));
 sg13g2_buf_4 fanout543 (.X(net543),
    .A(net545));
 sg13g2_buf_2 fanout544 (.A(net545),
    .X(net544));
 sg13g2_buf_4 fanout545 (.X(net545),
    .A(_0782_));
 sg13g2_buf_4 fanout546 (.X(net546),
    .A(net550));
 sg13g2_buf_2 fanout547 (.A(net550),
    .X(net547));
 sg13g2_buf_4 fanout548 (.X(net548),
    .A(net550));
 sg13g2_buf_1 fanout549 (.A(net550),
    .X(net549));
 sg13g2_buf_4 fanout550 (.X(net550),
    .A(_0781_));
 sg13g2_buf_2 fanout551 (.A(net552),
    .X(net551));
 sg13g2_buf_2 fanout552 (.A(_0779_),
    .X(net552));
 sg13g2_buf_4 fanout553 (.X(net553),
    .A(_0779_));
 sg13g2_buf_4 fanout554 (.X(net554),
    .A(net555));
 sg13g2_buf_4 fanout555 (.X(net555),
    .A(_0776_));
 sg13g2_buf_4 fanout556 (.X(net556),
    .A(net558));
 sg13g2_buf_4 fanout557 (.X(net557),
    .A(net558));
 sg13g2_buf_4 fanout558 (.X(net558),
    .A(_0771_));
 sg13g2_buf_2 fanout559 (.A(net560),
    .X(net559));
 sg13g2_buf_4 fanout560 (.X(net560),
    .A(_0766_));
 sg13g2_buf_4 fanout561 (.X(net561),
    .A(_0535_));
 sg13g2_buf_4 fanout562 (.X(net562),
    .A(_0534_));
 sg13g2_buf_2 fanout563 (.A(net565),
    .X(net563));
 sg13g2_buf_2 fanout564 (.A(net565),
    .X(net564));
 sg13g2_buf_2 fanout565 (.A(_0246_),
    .X(net565));
 sg13g2_buf_2 fanout566 (.A(_0243_),
    .X(net566));
 sg13g2_buf_1 fanout567 (.A(_0243_),
    .X(net567));
 sg13g2_buf_2 fanout568 (.A(net569),
    .X(net568));
 sg13g2_buf_2 fanout569 (.A(net570),
    .X(net569));
 sg13g2_buf_4 fanout570 (.X(net570),
    .A(_0836_));
 sg13g2_buf_2 fanout571 (.A(net572),
    .X(net571));
 sg13g2_buf_4 fanout572 (.X(net572),
    .A(_0800_));
 sg13g2_buf_4 fanout573 (.X(net573),
    .A(_0795_));
 sg13g2_buf_2 fanout574 (.A(_0793_),
    .X(net574));
 sg13g2_buf_4 fanout575 (.X(net575),
    .A(net577));
 sg13g2_buf_1 fanout576 (.A(net577),
    .X(net576));
 sg13g2_buf_2 fanout577 (.A(_0786_),
    .X(net577));
 sg13g2_buf_4 fanout578 (.X(net578),
    .A(net579));
 sg13g2_buf_2 fanout579 (.A(net580),
    .X(net579));
 sg13g2_buf_2 fanout580 (.A(_0775_),
    .X(net580));
 sg13g2_buf_2 fanout581 (.A(net583),
    .X(net581));
 sg13g2_buf_2 fanout582 (.A(net583),
    .X(net582));
 sg13g2_buf_1 fanout583 (.A(net584),
    .X(net583));
 sg13g2_buf_2 fanout584 (.A(_0773_),
    .X(net584));
 sg13g2_buf_2 fanout585 (.A(_0768_),
    .X(net585));
 sg13g2_buf_4 fanout586 (.X(net586),
    .A(_0765_));
 sg13g2_buf_2 fanout587 (.A(net588),
    .X(net587));
 sg13g2_buf_4 fanout588 (.X(net588),
    .A(_0765_));
 sg13g2_buf_4 fanout589 (.X(net589),
    .A(_0763_));
 sg13g2_buf_2 fanout590 (.A(_0763_),
    .X(net590));
 sg13g2_buf_2 fanout591 (.A(_0761_),
    .X(net591));
 sg13g2_buf_2 fanout592 (.A(net594),
    .X(net592));
 sg13g2_buf_2 fanout593 (.A(net594),
    .X(net593));
 sg13g2_buf_2 fanout594 (.A(_0605_),
    .X(net594));
 sg13g2_buf_2 fanout595 (.A(net596),
    .X(net595));
 sg13g2_buf_4 fanout596 (.X(net596),
    .A(_0605_));
 sg13g2_buf_4 fanout597 (.X(net597),
    .A(net599));
 sg13g2_buf_2 fanout598 (.A(net599),
    .X(net598));
 sg13g2_buf_2 fanout599 (.A(\main.demo._q_addr[7] ),
    .X(net599));
 sg13g2_buf_2 fanout600 (.A(\main.demo._q_addr[6] ),
    .X(net600));
 sg13g2_buf_2 fanout601 (.A(\main.demo._q_addr[5] ),
    .X(net601));
 sg13g2_buf_2 fanout602 (.A(\main.demo._q_addr[4] ),
    .X(net602));
 sg13g2_buf_2 fanout603 (.A(\main.demo._q_addr[3] ),
    .X(net603));
 sg13g2_buf_2 fanout604 (.A(net605),
    .X(net604));
 sg13g2_buf_2 fanout605 (.A(\main.demo._q_addr[2] ),
    .X(net605));
 sg13g2_buf_2 fanout606 (.A(net607),
    .X(net606));
 sg13g2_buf_2 fanout607 (.A(\main.demo._q_addr[1] ),
    .X(net607));
 sg13g2_buf_2 fanout608 (.A(\main.demo._q_addr[0] ),
    .X(net608));
 sg13g2_buf_2 fanout609 (.A(net611),
    .X(net609));
 sg13g2_buf_2 fanout610 (.A(net611),
    .X(net610));
 sg13g2_buf_2 fanout611 (.A(net334),
    .X(net611));
 sg13g2_buf_4 fanout612 (.X(net612),
    .A(net613));
 sg13g2_buf_2 fanout613 (.A(net334),
    .X(net613));
 sg13g2_buf_2 input1 (.A(rst_n),
    .X(net1));
 sg13g2_tielo tt_um_whynot_2 (.L_LO(net2));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_buf_2 clkbuf_5_0__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_0__leaf_clk));
 sg13g2_buf_2 clkbuf_5_1__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_1__leaf_clk));
 sg13g2_buf_2 clkbuf_5_2__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_2__leaf_clk));
 sg13g2_buf_2 clkbuf_5_3__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_3__leaf_clk));
 sg13g2_buf_2 clkbuf_5_4__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_4__leaf_clk));
 sg13g2_buf_2 clkbuf_5_5__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_5__leaf_clk));
 sg13g2_buf_2 clkbuf_5_6__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_6__leaf_clk));
 sg13g2_buf_2 clkbuf_5_7__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_7__leaf_clk));
 sg13g2_buf_2 clkbuf_5_8__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_8__leaf_clk));
 sg13g2_buf_2 clkbuf_5_9__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_9__leaf_clk));
 sg13g2_buf_2 clkbuf_5_10__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_10__leaf_clk));
 sg13g2_buf_2 clkbuf_5_11__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_11__leaf_clk));
 sg13g2_buf_2 clkbuf_5_12__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_12__leaf_clk));
 sg13g2_buf_2 clkbuf_5_13__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_13__leaf_clk));
 sg13g2_buf_2 clkbuf_5_14__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_14__leaf_clk));
 sg13g2_buf_2 clkbuf_5_15__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_15__leaf_clk));
 sg13g2_buf_2 clkbuf_5_16__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_16__leaf_clk));
 sg13g2_buf_2 clkbuf_5_17__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_17__leaf_clk));
 sg13g2_buf_2 clkbuf_5_18__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_18__leaf_clk));
 sg13g2_buf_2 clkbuf_5_19__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_19__leaf_clk));
 sg13g2_buf_2 clkbuf_5_20__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_20__leaf_clk));
 sg13g2_buf_2 clkbuf_5_21__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_21__leaf_clk));
 sg13g2_buf_2 clkbuf_5_22__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_22__leaf_clk));
 sg13g2_buf_2 clkbuf_5_23__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_23__leaf_clk));
 sg13g2_buf_2 clkbuf_5_24__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_24__leaf_clk));
 sg13g2_buf_2 clkbuf_5_25__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_25__leaf_clk));
 sg13g2_buf_2 clkbuf_5_26__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_26__leaf_clk));
 sg13g2_buf_2 clkbuf_5_27__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_27__leaf_clk));
 sg13g2_buf_2 clkbuf_5_28__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_28__leaf_clk));
 sg13g2_buf_2 clkbuf_5_29__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_29__leaf_clk));
 sg13g2_buf_2 clkbuf_5_30__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_30__leaf_clk));
 sg13g2_buf_2 clkbuf_5_31__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_31__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_5_3__leaf_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_5_5__leaf_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_5_7__leaf_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_5_9__leaf_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_5_11__leaf_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_5_13__leaf_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_5_15__leaf_clk));
 sg13g2_inv_1 clkload7 (.A(clknet_5_19__leaf_clk));
 sg13g2_inv_1 clkload8 (.A(clknet_5_21__leaf_clk));
 sg13g2_inv_1 clkload9 (.A(clknet_5_23__leaf_clk));
 sg13g2_inv_1 clkload10 (.A(clknet_5_25__leaf_clk));
 sg13g2_inv_1 clkload11 (.A(clknet_5_27__leaf_clk));
 sg13g2_inv_1 clkload12 (.A(clknet_5_29__leaf_clk));
 sg13g2_inv_1 clkload13 (.A(clknet_5_31__leaf_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(_0017_),
    .X(net163));
 sg13g2_dlygate4sd3_1 hold2 (.A(\main._w_demo_video_vs ),
    .X(net164));
 sg13g2_dlygate4sd3_1 hold3 (.A(\main.demo.zic._d_clock_count[0] ),
    .X(net165));
 sg13g2_dlygate4sd3_1 hold4 (.A(_0019_),
    .X(net166));
 sg13g2_dlygate4sd3_1 hold5 (.A(_0029_),
    .X(net167));
 sg13g2_dlygate4sd3_1 hold6 (.A(_0014_),
    .X(net168));
 sg13g2_dlygate4sd3_1 hold7 (.A(_0020_),
    .X(net169));
 sg13g2_dlygate4sd3_1 hold8 (.A(_0021_),
    .X(net170));
 sg13g2_dlygate4sd3_1 hold9 (.A(_0018_),
    .X(net171));
 sg13g2_dlygate4sd3_1 hold10 (.A(_0071_),
    .X(net172));
 sg13g2_dlygate4sd3_1 hold11 (.A(\main._w_demo_video_hs ),
    .X(net173));
 sg13g2_dlygate4sd3_1 hold12 (.A(\main.demo.zic._q_qpos[0] ),
    .X(net174));
 sg13g2_dlygate4sd3_1 hold13 (.A(\main.demo.zic._q_clock_count[8] ),
    .X(net175));
 sg13g2_dlygate4sd3_1 hold14 (.A(_0105_),
    .X(net176));
 sg13g2_dlygate4sd3_1 hold15 (.A(\main.demo._w_vga_active ),
    .X(net177));
 sg13g2_dlygate4sd3_1 hold16 (.A(\main.demo.zic._q_qpos[11] ),
    .X(net178));
 sg13g2_dlygate4sd3_1 hold17 (.A(_0365_),
    .X(net179));
 sg13g2_dlygate4sd3_1 hold18 (.A(_0069_),
    .X(net180));
 sg13g2_dlygate4sd3_1 hold19 (.A(\main.demo.zic._q_clock_count[6] ),
    .X(net181));
 sg13g2_dlygate4sd3_1 hold20 (.A(_0103_),
    .X(net182));
 sg13g2_dlygate4sd3_1 hold21 (.A(\main.demo.vga._q_xcount[3] ),
    .X(net183));
 sg13g2_dlygate4sd3_1 hold22 (.A(_0530_),
    .X(net184));
 sg13g2_dlygate4sd3_1 hold23 (.A(_0120_),
    .X(net185));
 sg13g2_dlygate4sd3_1 hold24 (.A(\main.demo.zic._q_rythm_count[12] ),
    .X(net186));
 sg13g2_dlygate4sd3_1 hold25 (.A(_0394_),
    .X(net187));
 sg13g2_dlygate4sd3_1 hold26 (.A(_0083_),
    .X(net188));
 sg13g2_dlygate4sd3_1 hold27 (.A(\main.demo.zic._q_qpos[7] ),
    .X(net189));
 sg13g2_dlygate4sd3_1 hold28 (.A(_0357_),
    .X(net190));
 sg13g2_dlygate4sd3_1 hold29 (.A(_0065_),
    .X(net191));
 sg13g2_dlygate4sd3_1 hold30 (.A(\main.demo.vga._q_xcount[0] ),
    .X(net192));
 sg13g2_dlygate4sd3_1 hold31 (.A(\main.demo.vga._q_xcount[1] ),
    .X(net193));
 sg13g2_dlygate4sd3_1 hold32 (.A(_0037_),
    .X(net194));
 sg13g2_dlygate4sd3_1 hold33 (.A(_0013_),
    .X(net195));
 sg13g2_dlygate4sd3_1 hold34 (.A(\main.demo._q_v[1] ),
    .X(net196));
 sg13g2_dlygate4sd3_1 hold35 (.A(_0249_),
    .X(net197));
 sg13g2_dlygate4sd3_1 hold36 (.A(_0030_),
    .X(net198));
 sg13g2_dlygate4sd3_1 hold37 (.A(\main.demo.zic._q_clock_count[7] ),
    .X(net199));
 sg13g2_dlygate4sd3_1 hold38 (.A(_0104_),
    .X(net200));
 sg13g2_dlygate4sd3_1 hold39 (.A(\main.demo._q_uT[11] ),
    .X(net201));
 sg13g2_dlygate4sd3_1 hold40 (.A(_0576_),
    .X(net202));
 sg13g2_dlygate4sd3_1 hold41 (.A(_0134_),
    .X(net203));
 sg13g2_dlygate4sd3_1 hold42 (.A(\main.demo.zic._q_rythm_count[7] ),
    .X(net204));
 sg13g2_dlygate4sd3_1 hold43 (.A(_0384_),
    .X(net205));
 sg13g2_dlygate4sd3_1 hold44 (.A(_0078_),
    .X(net206));
 sg13g2_dlygate4sd3_1 hold45 (.A(\main.demo._q_uT[9] ),
    .X(net207));
 sg13g2_dlygate4sd3_1 hold46 (.A(_0573_),
    .X(net208));
 sg13g2_dlygate4sd3_1 hold47 (.A(_0132_),
    .X(net209));
 sg13g2_dlygate4sd3_1 hold48 (.A(_0012_),
    .X(net210));
 sg13g2_dlygate4sd3_1 hold49 (.A(\main.demo.vga._q_ycount[0] ),
    .X(net211));
 sg13g2_dlygate4sd3_1 hold50 (.A(_0039_),
    .X(net212));
 sg13g2_dlygate4sd3_1 hold51 (.A(\main.demo.zic._q_rythm_count[1] ),
    .X(net213));
 sg13g2_dlygate4sd3_1 hold52 (.A(_0373_),
    .X(net214));
 sg13g2_dlygate4sd3_1 hold53 (.A(_0072_),
    .X(net215));
 sg13g2_dlygate4sd3_1 hold54 (.A(\main.demo.zic._q_qpos[1] ),
    .X(net216));
 sg13g2_dlygate4sd3_1 hold55 (.A(_0059_),
    .X(net217));
 sg13g2_dlygate4sd3_1 hold56 (.A(\main.demo.zic._q_qpos[3] ),
    .X(net218));
 sg13g2_dlygate4sd3_1 hold57 (.A(_0061_),
    .X(net219));
 sg13g2_dlygate4sd3_1 hold58 (.A(\main.demo.vga._q_xcount[7] ),
    .X(net220));
 sg13g2_dlygate4sd3_1 hold59 (.A(_0532_),
    .X(net221));
 sg13g2_dlygate4sd3_1 hold60 (.A(_0122_),
    .X(net222));
 sg13g2_dlygate4sd3_1 hold61 (.A(\main.demo.vga._q_active_h ),
    .X(net223));
 sg13g2_dlygate4sd3_1 hold62 (.A(_0625_),
    .X(net224));
 sg13g2_dlygate4sd3_1 hold63 (.A(\main.demo._q_u[0] ),
    .X(net225));
 sg13g2_dlygate4sd3_1 hold64 (.A(_0578_),
    .X(net226));
 sg13g2_dlygate4sd3_1 hold65 (.A(_0136_),
    .X(net227));
 sg13g2_dlygate4sd3_1 hold66 (.A(\main.demo.zic._q_qpos[5] ),
    .X(net228));
 sg13g2_dlygate4sd3_1 hold67 (.A(_0353_),
    .X(net229));
 sg13g2_dlygate4sd3_1 hold68 (.A(_0063_),
    .X(net230));
 sg13g2_dlygate4sd3_1 hold69 (.A(\main.demo._q_uT[8] ),
    .X(net231));
 sg13g2_dlygate4sd3_1 hold70 (.A(_0131_),
    .X(net232));
 sg13g2_dlygate4sd3_1 hold71 (.A(_0016_),
    .X(net233));
 sg13g2_dlygate4sd3_1 hold72 (.A(\main.demo._q_v[6] ),
    .X(net234));
 sg13g2_dlygate4sd3_1 hold73 (.A(_0257_),
    .X(net235));
 sg13g2_dlygate4sd3_1 hold74 (.A(_0035_),
    .X(net236));
 sg13g2_dlygate4sd3_1 hold75 (.A(\main.demo.vga._q_xcount[9] ),
    .X(net237));
 sg13g2_dlygate4sd3_1 hold76 (.A(_0278_),
    .X(net238));
 sg13g2_dlygate4sd3_1 hold77 (.A(_0046_),
    .X(net239));
 sg13g2_dlygate4sd3_1 hold78 (.A(\main.demo._q_vT[11] ),
    .X(net240));
 sg13g2_dlygate4sd3_1 hold79 (.A(_0527_),
    .X(net241));
 sg13g2_dlygate4sd3_1 hold80 (.A(\main.demo.zic._q_clock_count[5] ),
    .X(net242));
 sg13g2_dlygate4sd3_1 hold81 (.A(_0438_),
    .X(net243));
 sg13g2_dlygate4sd3_1 hold82 (.A(\main.demo._q_v[4] ),
    .X(net244));
 sg13g2_dlygate4sd3_1 hold83 (.A(_0254_),
    .X(net245));
 sg13g2_dlygate4sd3_1 hold84 (.A(\main.demo._q_u[6] ),
    .X(net246));
 sg13g2_dlygate4sd3_1 hold85 (.A(_0587_),
    .X(net247));
 sg13g2_dlygate4sd3_1 hold86 (.A(_0141_),
    .X(net248));
 sg13g2_dlygate4sd3_1 hold87 (.A(\main.demo._q_vT[1] ),
    .X(net249));
 sg13g2_dlygate4sd3_1 hold88 (.A(_0107_),
    .X(net250));
 sg13g2_dlygate4sd3_1 hold89 (.A(\main.demo.vga._q_ycount[3] ),
    .X(net251));
 sg13g2_dlygate4sd3_1 hold90 (.A(_0051_),
    .X(net252));
 sg13g2_dlygate4sd3_1 hold91 (.A(\main.demo.zic._q_rythm_count[11] ),
    .X(net253));
 sg13g2_dlygate4sd3_1 hold92 (.A(_0392_),
    .X(net254));
 sg13g2_dlygate4sd3_1 hold93 (.A(\main.demo._q_v[2] ),
    .X(net255));
 sg13g2_dlygate4sd3_1 hold94 (.A(_0250_),
    .X(net256));
 sg13g2_dlygate4sd3_1 hold95 (.A(\main.demo._q_vT[10] ),
    .X(net257));
 sg13g2_dlygate4sd3_1 hold96 (.A(_0525_),
    .X(net258));
 sg13g2_dlygate4sd3_1 hold97 (.A(_0116_),
    .X(net259));
 sg13g2_dlygate4sd3_1 hold98 (.A(\main.demo.zic._q_rythm_count[3] ),
    .X(net260));
 sg13g2_dlygate4sd3_1 hold99 (.A(_0377_),
    .X(net261));
 sg13g2_dlygate4sd3_1 hold100 (.A(_0074_),
    .X(net262));
 sg13g2_dlygate4sd3_1 hold101 (.A(\main.demo.zic._q_rythm_count[10] ),
    .X(net263));
 sg13g2_dlygate4sd3_1 hold102 (.A(_0390_),
    .X(net264));
 sg13g2_dlygate4sd3_1 hold103 (.A(_0081_),
    .X(net265));
 sg13g2_dlygate4sd3_1 hold104 (.A(\main.demo.zic._q_rythm_count[2] ),
    .X(net266));
 sg13g2_dlygate4sd3_1 hold105 (.A(_0375_),
    .X(net267));
 sg13g2_dlygate4sd3_1 hold106 (.A(_0073_),
    .X(net268));
 sg13g2_dlygate4sd3_1 hold107 (.A(\main.demo.zic._q_rythm_count[5] ),
    .X(net269));
 sg13g2_dlygate4sd3_1 hold108 (.A(_0381_),
    .X(net270));
 sg13g2_dlygate4sd3_1 hold109 (.A(_0076_),
    .X(net271));
 sg13g2_dlygate4sd3_1 hold110 (.A(\main.demo._q_vT[0] ),
    .X(net272));
 sg13g2_dlygate4sd3_1 hold111 (.A(\main.demo.zic._q_rythm_count[8] ),
    .X(net273));
 sg13g2_dlygate4sd3_1 hold112 (.A(_0386_),
    .X(net274));
 sg13g2_dlygate4sd3_1 hold113 (.A(_0079_),
    .X(net275));
 sg13g2_dlygate4sd3_1 hold114 (.A(\main.demo.zic._q_rythm_count[9] ),
    .X(net276));
 sg13g2_dlygate4sd3_1 hold115 (.A(_0388_),
    .X(net277));
 sg13g2_dlygate4sd3_1 hold116 (.A(_0080_),
    .X(net278));
 sg13g2_dlygate4sd3_1 hold117 (.A(\main.demo.vga._q_ycount[6] ),
    .X(net279));
 sg13g2_dlygate4sd3_1 hold118 (.A(_0289_),
    .X(net280));
 sg13g2_dlygate4sd3_1 hold119 (.A(\main.demo._q_frame[3] ),
    .X(net281));
 sg13g2_dlygate4sd3_1 hold120 (.A(\main.demo.vga._q_xcount[2] ),
    .X(net282));
 sg13g2_dlygate4sd3_1 hold121 (.A(\main.demo.zic._q_squ_env[2] ),
    .X(net283));
 sg13g2_dlygate4sd3_1 hold122 (.A(_0422_),
    .X(net284));
 sg13g2_dlygate4sd3_1 hold123 (.A(_0093_),
    .X(net285));
 sg13g2_dlygate4sd3_1 hold124 (.A(\main.demo._q_v[3] ),
    .X(net286));
 sg13g2_dlygate4sd3_1 hold125 (.A(\main.demo.zic._q_qpos[8] ),
    .X(net287));
 sg13g2_dlygate4sd3_1 hold126 (.A(_0359_),
    .X(net288));
 sg13g2_dlygate4sd3_1 hold127 (.A(_0066_),
    .X(net289));
 sg13g2_dlygate4sd3_1 hold128 (.A(\main.demo._q_uT[0] ),
    .X(net290));
 sg13g2_dlygate4sd3_1 hold129 (.A(_0124_),
    .X(net291));
 sg13g2_dlygate4sd3_1 hold130 (.A(\main.demo._q_uT[10] ),
    .X(net292));
 sg13g2_dlygate4sd3_1 hold131 (.A(\main.demo._q_vT[3] ),
    .X(net293));
 sg13g2_dlygate4sd3_1 hold132 (.A(\main.demo._q_vT[4] ),
    .X(net294));
 sg13g2_dlygate4sd3_1 hold133 (.A(\main.demo.zic._q_rythm_count[6] ),
    .X(net295));
 sg13g2_dlygate4sd3_1 hold134 (.A(_0383_),
    .X(net296));
 sg13g2_dlygate4sd3_1 hold135 (.A(_0077_),
    .X(net297));
 sg13g2_dlygate4sd3_1 hold136 (.A(\main.demo._q_u[3] ),
    .X(net298));
 sg13g2_dlygate4sd3_1 hold137 (.A(_0582_),
    .X(net299));
 sg13g2_dlygate4sd3_1 hold138 (.A(_0138_),
    .X(net300));
 sg13g2_dlygate4sd3_1 hold139 (.A(\main.demo.zic._q_clock_count[2] ),
    .X(net301));
 sg13g2_dlygate4sd3_1 hold140 (.A(_0431_),
    .X(net302));
 sg13g2_dlygate4sd3_1 hold141 (.A(\main.demo._q_v[7] ),
    .X(net303));
 sg13g2_dlygate4sd3_1 hold142 (.A(\main.demo.zic._q_rythm_count[4] ),
    .X(net304));
 sg13g2_dlygate4sd3_1 hold143 (.A(\main.demo.zic._q_squ_env[5] ),
    .X(net305));
 sg13g2_dlygate4sd3_1 hold144 (.A(_0096_),
    .X(net306));
 sg13g2_dlygate4sd3_1 hold145 (.A(\main.demo.vga._q_active_v ),
    .X(net307));
 sg13g2_dlygate4sd3_1 hold146 (.A(\main.demo.vga._q_ycount[1] ),
    .X(net308));
 sg13g2_dlygate4sd3_1 hold147 (.A(\main.demo.zic._q_qpos[4] ),
    .X(net309));
 sg13g2_dlygate4sd3_1 hold148 (.A(_0062_),
    .X(net310));
 sg13g2_dlygate4sd3_1 hold149 (.A(\main.demo._q_u[7] ),
    .X(net311));
 sg13g2_dlygate4sd3_1 hold150 (.A(_0590_),
    .X(net312));
 sg13g2_dlygate4sd3_1 hold151 (.A(\main.demo.zic._q_qpos[2] ),
    .X(net313));
 sg13g2_dlygate4sd3_1 hold152 (.A(\main.demo.vga._q_ycount[7] ),
    .X(net314));
 sg13g2_dlygate4sd3_1 hold153 (.A(\main.demo._q_frame[4] ),
    .X(net315));
 sg13g2_dlygate4sd3_1 hold154 (.A(_0474_),
    .X(net316));
 sg13g2_dlygate4sd3_1 hold155 (.A(\main.demo._q_v[5] ),
    .X(net317));
 sg13g2_dlygate4sd3_1 hold156 (.A(\main.demo.zic._q_squ_env[0] ),
    .X(net318));
 sg13g2_dlygate4sd3_1 hold157 (.A(\main.demo.zic._q_qpos[6] ),
    .X(net319));
 sg13g2_dlygate4sd3_1 hold158 (.A(_0356_),
    .X(net320));
 sg13g2_dlygate4sd3_1 hold159 (.A(_0064_),
    .X(net321));
 sg13g2_dlygate4sd3_1 hold160 (.A(\main.demo.zic._q_clock_count[4] ),
    .X(net322));
 sg13g2_dlygate4sd3_1 hold161 (.A(_0437_),
    .X(net323));
 sg13g2_dlygate4sd3_1 hold162 (.A(\main.demo._q_vT[5] ),
    .X(net324));
 sg13g2_dlygate4sd3_1 hold163 (.A(\main.demo._q_frame[6] ),
    .X(net325));
 sg13g2_dlygate4sd3_1 hold164 (.A(_0493_),
    .X(net326));
 sg13g2_dlygate4sd3_1 hold165 (.A(\main.demo.zic._q_qpos[12] ),
    .X(net327));
 sg13g2_dlygate4sd3_1 hold166 (.A(_0070_),
    .X(net328));
 sg13g2_dlygate4sd3_1 hold167 (.A(\main.demo.vga._q_ycount[5] ),
    .X(net329));
 sg13g2_dlygate4sd3_1 hold168 (.A(_0288_),
    .X(net330));
 sg13g2_dlygate4sd3_1 hold169 (.A(_0053_),
    .X(net331));
 sg13g2_dlygate4sd3_1 hold170 (.A(\main.demo._q_u[4] ),
    .X(net332));
 sg13g2_dlygate4sd3_1 hold171 (.A(_0585_),
    .X(net333));
 sg13g2_dlygate4sd3_1 hold172 (.A(rst_n_q),
    .X(net334));
 sg13g2_dlygate4sd3_1 hold173 (.A(_0048_),
    .X(net335));
 sg13g2_dlygate4sd3_1 hold174 (.A(\main.demo.vga._q_xcount[5] ),
    .X(net336));
 sg13g2_dlygate4sd3_1 hold175 (.A(_0268_),
    .X(net337));
 sg13g2_dlygate4sd3_1 hold176 (.A(_0040_),
    .X(net338));
 sg13g2_dlygate4sd3_1 hold177 (.A(\main.demo.vga._q_xcount[4] ),
    .X(net339));
 sg13g2_dlygate4sd3_1 hold178 (.A(\main.demo._q_u[5] ),
    .X(net340));
 sg13g2_dlygate4sd3_1 hold179 (.A(\main.demo.zic._q_qpos[10] ),
    .X(net341));
 sg13g2_dlygate4sd3_1 hold180 (.A(_0363_),
    .X(net342));
 sg13g2_dlygate4sd3_1 hold181 (.A(_0068_),
    .X(net343));
 sg13g2_dlygate4sd3_1 hold182 (.A(_0003_),
    .X(net344));
 sg13g2_dlygate4sd3_1 hold183 (.A(_0484_),
    .X(net345));
 sg13g2_dlygate4sd3_1 hold184 (.A(\main.demo.zic._q_clock_count[3] ),
    .X(net346));
 sg13g2_dlygate4sd3_1 hold185 (.A(\main.demo.zic._q_squ_env[1] ),
    .X(net347));
 sg13g2_dlygate4sd3_1 hold186 (.A(_0092_),
    .X(net348));
 sg13g2_dlygate4sd3_1 hold187 (.A(\main.demo.vga._d_vblank ),
    .X(net349));
 sg13g2_dlygate4sd3_1 hold188 (.A(_0242_),
    .X(net350));
 sg13g2_dlygate4sd3_1 hold189 (.A(_0028_),
    .X(net351));
 sg13g2_dlygate4sd3_1 hold190 (.A(\main.demo._q_vT[8] ),
    .X(net352));
 sg13g2_dlygate4sd3_1 hold191 (.A(\main.demo.vga._q_xcount[10] ),
    .X(net353));
 sg13g2_dlygate4sd3_1 hold192 (.A(\main.demo.zic._q_squ_env[4] ),
    .X(net354));
 sg13g2_dlygate4sd3_1 hold193 (.A(_0427_),
    .X(net355));
 sg13g2_dlygate4sd3_1 hold194 (.A(_0095_),
    .X(net356));
 sg13g2_dlygate4sd3_1 hold195 (.A(\main.demo.zic._q_clock_count[0] ),
    .X(net357));
 sg13g2_dlygate4sd3_1 hold196 (.A(_0430_),
    .X(net358));
 sg13g2_dlygate4sd3_1 hold197 (.A(_0098_),
    .X(net359));
 sg13g2_dlygate4sd3_1 hold198 (.A(\main.demo._q_frame[1] ),
    .X(net360));
 sg13g2_dlygate4sd3_1 hold199 (.A(\main.demo._q_frame[8] ),
    .X(net361));
 sg13g2_dlygate4sd3_1 hold200 (.A(\main.demo.vga._q_xcount[6] ),
    .X(net362));
 sg13g2_dlygate4sd3_1 hold201 (.A(_0275_),
    .X(net363));
 sg13g2_dlygate4sd3_1 hold202 (.A(\main.demo.vga._d_vblank ),
    .X(net364));
 sg13g2_dlygate4sd3_1 hold203 (.A(\main.demo._q_vT[2] ),
    .X(net365));
 sg13g2_dlygate4sd3_1 hold204 (.A(_0473_),
    .X(net366));
 sg13g2_dlygate4sd3_1 hold205 (.A(\main.demo._q_u[2] ),
    .X(net367));
 sg13g2_dlygate4sd3_1 hold206 (.A(_0581_),
    .X(net368));
 sg13g2_dlygate4sd3_1 hold207 (.A(\main.demo._q_frame[2] ),
    .X(net369));
 sg13g2_dlygate4sd3_1 hold208 (.A(_0459_),
    .X(net370));
 sg13g2_dlygate4sd3_1 hold209 (.A(\main.demo._q_vT[9] ),
    .X(net371));
 sg13g2_dlygate4sd3_1 hold210 (.A(\main.demo._q_vT[7] ),
    .X(net372));
 sg13g2_dlygate4sd3_1 hold211 (.A(\main.demo.vga._q_ycount[2] ),
    .X(net373));
 sg13g2_dlygate4sd3_1 hold212 (.A(_0286_),
    .X(net374));
 sg13g2_dlygate4sd3_1 hold213 (.A(_0050_),
    .X(net375));
 sg13g2_dlygate4sd3_1 hold214 (.A(\main.demo._q_uT[3] ),
    .X(net376));
 sg13g2_dlygate4sd3_1 hold215 (.A(_0126_),
    .X(net377));
 sg13g2_dlygate4sd3_1 hold216 (.A(\main.demo.vga._q_xcount[8] ),
    .X(net378));
 sg13g2_dlygate4sd3_1 hold217 (.A(\main.demo.zic._q_idx[0] ),
    .X(net379));
 sg13g2_dlygate4sd3_1 hold218 (.A(_0396_),
    .X(net380));
 sg13g2_dlygate4sd3_1 hold219 (.A(\main.demo.zic._q_qpos[9] ),
    .X(net381));
 sg13g2_dlygate4sd3_1 hold220 (.A(\main.demo.vga._q_ycount[8] ),
    .X(net382));
 sg13g2_dlygate4sd3_1 hold221 (.A(_0015_),
    .X(net383));
 sg13g2_dlygate4sd3_1 hold222 (.A(_0404_),
    .X(net384));
 sg13g2_dlygate4sd3_1 hold223 (.A(_0000_),
    .X(net385));
 sg13g2_dlygate4sd3_1 hold224 (.A(_0424_),
    .X(net386));
 sg13g2_dlygate4sd3_1 hold225 (.A(_0094_),
    .X(net387));
 sg13g2_dlygate4sd3_1 hold226 (.A(\main.demo._q_frame[7] ),
    .X(net388));
 sg13g2_dlygate4sd3_1 hold227 (.A(_0501_),
    .X(net389));
 sg13g2_dlygate4sd3_1 hold228 (.A(\main.demo._q_vT[6] ),
    .X(net390));
 sg13g2_dlygate4sd3_1 hold229 (.A(_0510_),
    .X(net391));
 sg13g2_dlygate4sd3_1 hold230 (.A(\main.demo._q_uT[1] ),
    .X(net392));
 sg13g2_dlygate4sd3_1 hold231 (.A(_0544_),
    .X(net393));
 sg13g2_dlygate4sd3_1 hold232 (.A(\main.demo._q_uT[6] ),
    .X(net394));
 sg13g2_dlygate4sd3_1 hold233 (.A(\main.demo.vga._q_ycount[4] ),
    .X(net395));
 sg13g2_dlygate4sd3_1 hold234 (.A(_0052_),
    .X(net396));
 sg13g2_dlygate4sd3_1 hold235 (.A(\main.demo.vga._q_ycount[0] ),
    .X(net397));
 sg13g2_dlygate4sd3_1 hold236 (.A(\main.demo._q_uT[5] ),
    .X(net398));
 sg13g2_dlygate4sd3_1 hold237 (.A(_0559_),
    .X(net399));
 sg13g2_dlygate4sd3_1 hold238 (.A(\main.demo._q_frame[5] ),
    .X(net400));
 sg13g2_dlygate4sd3_1 hold239 (.A(\main.demo.vga._q_xcount[8] ),
    .X(net401));
 sg13g2_dlygate4sd3_1 hold240 (.A(\main.demo._q_v[5] ),
    .X(net402));
 sg13g2_dlygate4sd3_1 hold241 (.A(\main.demo._q_uT[5] ),
    .X(net403));
 sg13g2_antennanp ANTENNA_1 (.A(clk));
 sg13g2_antennanp ANTENNA_2 (.A(clk));
 sg13g2_antennanp ANTENNA_3 (.A(net1));
 sg13g2_antennanp ANTENNA_4 (.A(clk));
 sg13g2_antennanp ANTENNA_5 (.A(net1));
 sg13g2_antennanp ANTENNA_6 (.A(net1));
 sg13g2_antennanp ANTENNA_7 (.A(net1));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_fill_1 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_166 ();
 sg13g2_decap_8 FILLER_2_173 ();
 sg13g2_decap_8 FILLER_2_180 ();
 sg13g2_decap_8 FILLER_2_187 ();
 sg13g2_decap_8 FILLER_2_194 ();
 sg13g2_decap_8 FILLER_2_201 ();
 sg13g2_decap_8 FILLER_2_208 ();
 sg13g2_decap_8 FILLER_2_215 ();
 sg13g2_decap_8 FILLER_2_222 ();
 sg13g2_decap_8 FILLER_2_229 ();
 sg13g2_decap_8 FILLER_2_236 ();
 sg13g2_decap_8 FILLER_2_243 ();
 sg13g2_decap_8 FILLER_2_250 ();
 sg13g2_decap_8 FILLER_2_257 ();
 sg13g2_decap_8 FILLER_2_264 ();
 sg13g2_decap_8 FILLER_2_271 ();
 sg13g2_decap_8 FILLER_2_278 ();
 sg13g2_decap_8 FILLER_2_285 ();
 sg13g2_decap_8 FILLER_2_292 ();
 sg13g2_decap_8 FILLER_2_299 ();
 sg13g2_decap_8 FILLER_2_306 ();
 sg13g2_decap_8 FILLER_2_313 ();
 sg13g2_decap_8 FILLER_2_320 ();
 sg13g2_decap_8 FILLER_2_327 ();
 sg13g2_decap_8 FILLER_2_334 ();
 sg13g2_decap_8 FILLER_2_341 ();
 sg13g2_decap_8 FILLER_2_348 ();
 sg13g2_decap_8 FILLER_2_355 ();
 sg13g2_decap_8 FILLER_2_362 ();
 sg13g2_decap_8 FILLER_2_369 ();
 sg13g2_decap_8 FILLER_2_376 ();
 sg13g2_decap_8 FILLER_2_383 ();
 sg13g2_decap_8 FILLER_2_390 ();
 sg13g2_decap_8 FILLER_2_397 ();
 sg13g2_decap_4 FILLER_2_404 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_181 ();
 sg13g2_decap_8 FILLER_3_188 ();
 sg13g2_decap_8 FILLER_3_195 ();
 sg13g2_decap_8 FILLER_3_202 ();
 sg13g2_fill_2 FILLER_3_209 ();
 sg13g2_fill_1 FILLER_3_211 ();
 sg13g2_decap_8 FILLER_3_221 ();
 sg13g2_decap_8 FILLER_3_228 ();
 sg13g2_decap_8 FILLER_3_235 ();
 sg13g2_decap_8 FILLER_3_242 ();
 sg13g2_decap_8 FILLER_3_249 ();
 sg13g2_decap_8 FILLER_3_256 ();
 sg13g2_decap_8 FILLER_3_263 ();
 sg13g2_decap_8 FILLER_3_270 ();
 sg13g2_decap_8 FILLER_3_277 ();
 sg13g2_decap_8 FILLER_3_284 ();
 sg13g2_decap_8 FILLER_3_291 ();
 sg13g2_decap_8 FILLER_3_298 ();
 sg13g2_decap_8 FILLER_3_305 ();
 sg13g2_decap_8 FILLER_3_312 ();
 sg13g2_decap_8 FILLER_3_319 ();
 sg13g2_decap_8 FILLER_3_326 ();
 sg13g2_decap_8 FILLER_3_333 ();
 sg13g2_decap_8 FILLER_3_340 ();
 sg13g2_decap_8 FILLER_3_347 ();
 sg13g2_decap_8 FILLER_3_354 ();
 sg13g2_decap_8 FILLER_3_361 ();
 sg13g2_decap_8 FILLER_3_368 ();
 sg13g2_decap_8 FILLER_3_375 ();
 sg13g2_decap_8 FILLER_3_382 ();
 sg13g2_decap_8 FILLER_3_389 ();
 sg13g2_decap_8 FILLER_3_396 ();
 sg13g2_decap_4 FILLER_3_403 ();
 sg13g2_fill_2 FILLER_3_407 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_4 FILLER_4_133 ();
 sg13g2_fill_1 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_188 ();
 sg13g2_fill_2 FILLER_4_195 ();
 sg13g2_fill_2 FILLER_4_207 ();
 sg13g2_fill_1 FILLER_4_209 ();
 sg13g2_decap_8 FILLER_4_229 ();
 sg13g2_decap_8 FILLER_4_236 ();
 sg13g2_decap_8 FILLER_4_243 ();
 sg13g2_decap_8 FILLER_4_250 ();
 sg13g2_decap_8 FILLER_4_257 ();
 sg13g2_decap_8 FILLER_4_264 ();
 sg13g2_decap_8 FILLER_4_271 ();
 sg13g2_decap_8 FILLER_4_278 ();
 sg13g2_decap_8 FILLER_4_285 ();
 sg13g2_decap_8 FILLER_4_292 ();
 sg13g2_decap_8 FILLER_4_299 ();
 sg13g2_decap_8 FILLER_4_306 ();
 sg13g2_decap_8 FILLER_4_313 ();
 sg13g2_decap_8 FILLER_4_320 ();
 sg13g2_decap_8 FILLER_4_327 ();
 sg13g2_decap_8 FILLER_4_334 ();
 sg13g2_decap_8 FILLER_4_341 ();
 sg13g2_decap_8 FILLER_4_348 ();
 sg13g2_decap_8 FILLER_4_355 ();
 sg13g2_decap_8 FILLER_4_362 ();
 sg13g2_decap_8 FILLER_4_369 ();
 sg13g2_decap_8 FILLER_4_376 ();
 sg13g2_decap_8 FILLER_4_383 ();
 sg13g2_decap_8 FILLER_4_390 ();
 sg13g2_decap_8 FILLER_4_397 ();
 sg13g2_decap_4 FILLER_4_404 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_4 FILLER_5_126 ();
 sg13g2_fill_1 FILLER_5_130 ();
 sg13g2_fill_1 FILLER_5_157 ();
 sg13g2_decap_8 FILLER_5_251 ();
 sg13g2_decap_8 FILLER_5_258 ();
 sg13g2_decap_8 FILLER_5_265 ();
 sg13g2_decap_8 FILLER_5_272 ();
 sg13g2_decap_8 FILLER_5_279 ();
 sg13g2_decap_8 FILLER_5_286 ();
 sg13g2_decap_8 FILLER_5_293 ();
 sg13g2_decap_8 FILLER_5_300 ();
 sg13g2_decap_8 FILLER_5_307 ();
 sg13g2_decap_8 FILLER_5_314 ();
 sg13g2_decap_8 FILLER_5_321 ();
 sg13g2_decap_8 FILLER_5_328 ();
 sg13g2_decap_8 FILLER_5_335 ();
 sg13g2_decap_8 FILLER_5_342 ();
 sg13g2_decap_8 FILLER_5_349 ();
 sg13g2_decap_8 FILLER_5_356 ();
 sg13g2_decap_8 FILLER_5_363 ();
 sg13g2_decap_8 FILLER_5_370 ();
 sg13g2_decap_8 FILLER_5_377 ();
 sg13g2_decap_8 FILLER_5_384 ();
 sg13g2_decap_8 FILLER_5_391 ();
 sg13g2_decap_8 FILLER_5_398 ();
 sg13g2_decap_4 FILLER_5_405 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_fill_2 FILLER_6_223 ();
 sg13g2_decap_8 FILLER_6_251 ();
 sg13g2_decap_8 FILLER_6_258 ();
 sg13g2_decap_8 FILLER_6_265 ();
 sg13g2_decap_8 FILLER_6_272 ();
 sg13g2_decap_8 FILLER_6_279 ();
 sg13g2_decap_8 FILLER_6_286 ();
 sg13g2_decap_8 FILLER_6_293 ();
 sg13g2_decap_8 FILLER_6_300 ();
 sg13g2_decap_8 FILLER_6_307 ();
 sg13g2_decap_8 FILLER_6_314 ();
 sg13g2_decap_8 FILLER_6_321 ();
 sg13g2_decap_8 FILLER_6_328 ();
 sg13g2_decap_8 FILLER_6_335 ();
 sg13g2_decap_8 FILLER_6_342 ();
 sg13g2_decap_8 FILLER_6_349 ();
 sg13g2_decap_8 FILLER_6_356 ();
 sg13g2_decap_8 FILLER_6_363 ();
 sg13g2_decap_8 FILLER_6_370 ();
 sg13g2_decap_8 FILLER_6_377 ();
 sg13g2_decap_8 FILLER_6_384 ();
 sg13g2_decap_8 FILLER_6_391 ();
 sg13g2_decap_8 FILLER_6_398 ();
 sg13g2_decap_4 FILLER_6_405 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_fill_2 FILLER_7_119 ();
 sg13g2_fill_1 FILLER_7_121 ();
 sg13g2_fill_1 FILLER_7_161 ();
 sg13g2_fill_2 FILLER_7_189 ();
 sg13g2_fill_2 FILLER_7_209 ();
 sg13g2_fill_1 FILLER_7_219 ();
 sg13g2_fill_2 FILLER_7_243 ();
 sg13g2_decap_8 FILLER_7_262 ();
 sg13g2_decap_8 FILLER_7_269 ();
 sg13g2_decap_8 FILLER_7_276 ();
 sg13g2_decap_8 FILLER_7_283 ();
 sg13g2_decap_8 FILLER_7_290 ();
 sg13g2_decap_8 FILLER_7_297 ();
 sg13g2_decap_8 FILLER_7_304 ();
 sg13g2_decap_8 FILLER_7_311 ();
 sg13g2_decap_8 FILLER_7_318 ();
 sg13g2_decap_8 FILLER_7_325 ();
 sg13g2_decap_8 FILLER_7_332 ();
 sg13g2_decap_8 FILLER_7_339 ();
 sg13g2_decap_8 FILLER_7_346 ();
 sg13g2_decap_8 FILLER_7_353 ();
 sg13g2_decap_8 FILLER_7_360 ();
 sg13g2_decap_8 FILLER_7_367 ();
 sg13g2_decap_8 FILLER_7_374 ();
 sg13g2_decap_8 FILLER_7_381 ();
 sg13g2_decap_8 FILLER_7_388 ();
 sg13g2_decap_8 FILLER_7_395 ();
 sg13g2_decap_8 FILLER_7_402 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_4 FILLER_8_119 ();
 sg13g2_fill_2 FILLER_8_170 ();
 sg13g2_fill_1 FILLER_8_197 ();
 sg13g2_fill_2 FILLER_8_216 ();
 sg13g2_decap_8 FILLER_8_249 ();
 sg13g2_decap_8 FILLER_8_256 ();
 sg13g2_decap_8 FILLER_8_263 ();
 sg13g2_decap_8 FILLER_8_270 ();
 sg13g2_decap_8 FILLER_8_277 ();
 sg13g2_decap_8 FILLER_8_284 ();
 sg13g2_decap_8 FILLER_8_291 ();
 sg13g2_decap_8 FILLER_8_298 ();
 sg13g2_decap_8 FILLER_8_305 ();
 sg13g2_decap_8 FILLER_8_312 ();
 sg13g2_decap_8 FILLER_8_319 ();
 sg13g2_decap_8 FILLER_8_326 ();
 sg13g2_decap_8 FILLER_8_333 ();
 sg13g2_decap_8 FILLER_8_340 ();
 sg13g2_decap_8 FILLER_8_347 ();
 sg13g2_decap_8 FILLER_8_354 ();
 sg13g2_decap_8 FILLER_8_361 ();
 sg13g2_decap_8 FILLER_8_368 ();
 sg13g2_decap_8 FILLER_8_375 ();
 sg13g2_decap_8 FILLER_8_382 ();
 sg13g2_decap_8 FILLER_8_389 ();
 sg13g2_decap_8 FILLER_8_396 ();
 sg13g2_decap_4 FILLER_8_403 ();
 sg13g2_fill_2 FILLER_8_407 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_4 FILLER_9_126 ();
 sg13g2_fill_1 FILLER_9_156 ();
 sg13g2_fill_1 FILLER_9_174 ();
 sg13g2_fill_2 FILLER_9_214 ();
 sg13g2_decap_8 FILLER_9_233 ();
 sg13g2_decap_8 FILLER_9_240 ();
 sg13g2_decap_8 FILLER_9_247 ();
 sg13g2_decap_8 FILLER_9_254 ();
 sg13g2_decap_8 FILLER_9_261 ();
 sg13g2_decap_8 FILLER_9_268 ();
 sg13g2_decap_8 FILLER_9_275 ();
 sg13g2_decap_8 FILLER_9_282 ();
 sg13g2_decap_8 FILLER_9_289 ();
 sg13g2_decap_8 FILLER_9_296 ();
 sg13g2_decap_8 FILLER_9_303 ();
 sg13g2_decap_8 FILLER_9_310 ();
 sg13g2_decap_8 FILLER_9_317 ();
 sg13g2_decap_8 FILLER_9_324 ();
 sg13g2_decap_8 FILLER_9_331 ();
 sg13g2_decap_8 FILLER_9_338 ();
 sg13g2_decap_8 FILLER_9_345 ();
 sg13g2_decap_8 FILLER_9_352 ();
 sg13g2_decap_8 FILLER_9_359 ();
 sg13g2_decap_8 FILLER_9_366 ();
 sg13g2_decap_8 FILLER_9_373 ();
 sg13g2_decap_8 FILLER_9_380 ();
 sg13g2_decap_8 FILLER_9_387 ();
 sg13g2_decap_8 FILLER_9_394 ();
 sg13g2_decap_8 FILLER_9_401 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_fill_1 FILLER_10_183 ();
 sg13g2_fill_1 FILLER_10_216 ();
 sg13g2_fill_2 FILLER_10_226 ();
 sg13g2_decap_8 FILLER_10_246 ();
 sg13g2_decap_8 FILLER_10_253 ();
 sg13g2_decap_8 FILLER_10_260 ();
 sg13g2_decap_8 FILLER_10_267 ();
 sg13g2_decap_8 FILLER_10_274 ();
 sg13g2_decap_8 FILLER_10_281 ();
 sg13g2_decap_8 FILLER_10_288 ();
 sg13g2_decap_8 FILLER_10_295 ();
 sg13g2_decap_8 FILLER_10_302 ();
 sg13g2_decap_8 FILLER_10_309 ();
 sg13g2_decap_8 FILLER_10_316 ();
 sg13g2_decap_8 FILLER_10_323 ();
 sg13g2_decap_8 FILLER_10_330 ();
 sg13g2_decap_8 FILLER_10_337 ();
 sg13g2_decap_8 FILLER_10_344 ();
 sg13g2_decap_8 FILLER_10_351 ();
 sg13g2_decap_8 FILLER_10_358 ();
 sg13g2_decap_8 FILLER_10_365 ();
 sg13g2_decap_8 FILLER_10_372 ();
 sg13g2_decap_8 FILLER_10_379 ();
 sg13g2_decap_8 FILLER_10_386 ();
 sg13g2_decap_8 FILLER_10_393 ();
 sg13g2_decap_8 FILLER_10_400 ();
 sg13g2_fill_2 FILLER_10_407 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_fill_1 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_250 ();
 sg13g2_decap_8 FILLER_11_257 ();
 sg13g2_decap_8 FILLER_11_264 ();
 sg13g2_decap_8 FILLER_11_271 ();
 sg13g2_decap_8 FILLER_11_278 ();
 sg13g2_decap_8 FILLER_11_285 ();
 sg13g2_decap_8 FILLER_11_292 ();
 sg13g2_decap_8 FILLER_11_299 ();
 sg13g2_decap_8 FILLER_11_306 ();
 sg13g2_decap_8 FILLER_11_313 ();
 sg13g2_decap_8 FILLER_11_320 ();
 sg13g2_decap_8 FILLER_11_327 ();
 sg13g2_decap_8 FILLER_11_334 ();
 sg13g2_decap_8 FILLER_11_341 ();
 sg13g2_decap_8 FILLER_11_348 ();
 sg13g2_decap_8 FILLER_11_355 ();
 sg13g2_decap_8 FILLER_11_362 ();
 sg13g2_decap_8 FILLER_11_369 ();
 sg13g2_decap_8 FILLER_11_376 ();
 sg13g2_decap_8 FILLER_11_383 ();
 sg13g2_decap_8 FILLER_11_390 ();
 sg13g2_decap_8 FILLER_11_397 ();
 sg13g2_decap_4 FILLER_11_404 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_4 FILLER_12_140 ();
 sg13g2_fill_1 FILLER_12_144 ();
 sg13g2_fill_2 FILLER_12_159 ();
 sg13g2_fill_1 FILLER_12_161 ();
 sg13g2_fill_2 FILLER_12_197 ();
 sg13g2_fill_2 FILLER_12_208 ();
 sg13g2_fill_2 FILLER_12_242 ();
 sg13g2_fill_1 FILLER_12_244 ();
 sg13g2_decap_8 FILLER_12_254 ();
 sg13g2_decap_8 FILLER_12_261 ();
 sg13g2_decap_8 FILLER_12_268 ();
 sg13g2_decap_8 FILLER_12_275 ();
 sg13g2_decap_8 FILLER_12_282 ();
 sg13g2_decap_8 FILLER_12_289 ();
 sg13g2_decap_8 FILLER_12_296 ();
 sg13g2_decap_8 FILLER_12_303 ();
 sg13g2_decap_8 FILLER_12_310 ();
 sg13g2_decap_8 FILLER_12_317 ();
 sg13g2_decap_8 FILLER_12_324 ();
 sg13g2_decap_8 FILLER_12_331 ();
 sg13g2_decap_8 FILLER_12_338 ();
 sg13g2_decap_8 FILLER_12_345 ();
 sg13g2_decap_8 FILLER_12_352 ();
 sg13g2_decap_8 FILLER_12_359 ();
 sg13g2_decap_8 FILLER_12_366 ();
 sg13g2_decap_8 FILLER_12_373 ();
 sg13g2_decap_8 FILLER_12_380 ();
 sg13g2_decap_8 FILLER_12_387 ();
 sg13g2_decap_8 FILLER_12_394 ();
 sg13g2_decap_8 FILLER_12_401 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_fill_2 FILLER_13_126 ();
 sg13g2_fill_1 FILLER_13_154 ();
 sg13g2_decap_4 FILLER_13_225 ();
 sg13g2_fill_1 FILLER_13_229 ();
 sg13g2_decap_8 FILLER_13_234 ();
 sg13g2_decap_8 FILLER_13_241 ();
 sg13g2_decap_8 FILLER_13_248 ();
 sg13g2_decap_8 FILLER_13_255 ();
 sg13g2_decap_8 FILLER_13_262 ();
 sg13g2_decap_8 FILLER_13_269 ();
 sg13g2_decap_8 FILLER_13_276 ();
 sg13g2_decap_8 FILLER_13_283 ();
 sg13g2_decap_8 FILLER_13_290 ();
 sg13g2_decap_8 FILLER_13_297 ();
 sg13g2_decap_8 FILLER_13_304 ();
 sg13g2_decap_8 FILLER_13_311 ();
 sg13g2_decap_8 FILLER_13_318 ();
 sg13g2_decap_8 FILLER_13_325 ();
 sg13g2_decap_8 FILLER_13_332 ();
 sg13g2_decap_8 FILLER_13_339 ();
 sg13g2_decap_8 FILLER_13_346 ();
 sg13g2_decap_8 FILLER_13_353 ();
 sg13g2_decap_8 FILLER_13_360 ();
 sg13g2_decap_8 FILLER_13_367 ();
 sg13g2_decap_8 FILLER_13_374 ();
 sg13g2_decap_8 FILLER_13_381 ();
 sg13g2_decap_8 FILLER_13_388 ();
 sg13g2_decap_8 FILLER_13_395 ();
 sg13g2_decap_8 FILLER_13_402 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_4 FILLER_14_119 ();
 sg13g2_fill_1 FILLER_14_123 ();
 sg13g2_fill_2 FILLER_14_162 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_fill_2 FILLER_14_406 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_4 FILLER_15_119 ();
 sg13g2_fill_1 FILLER_15_123 ();
 sg13g2_fill_2 FILLER_15_152 ();
 sg13g2_fill_1 FILLER_15_154 ();
 sg13g2_fill_2 FILLER_15_197 ();
 sg13g2_decap_8 FILLER_15_234 ();
 sg13g2_decap_8 FILLER_15_241 ();
 sg13g2_decap_8 FILLER_15_248 ();
 sg13g2_decap_8 FILLER_15_255 ();
 sg13g2_decap_8 FILLER_15_262 ();
 sg13g2_decap_8 FILLER_15_269 ();
 sg13g2_decap_8 FILLER_15_276 ();
 sg13g2_decap_8 FILLER_15_283 ();
 sg13g2_decap_8 FILLER_15_290 ();
 sg13g2_decap_8 FILLER_15_297 ();
 sg13g2_decap_8 FILLER_15_304 ();
 sg13g2_decap_8 FILLER_15_311 ();
 sg13g2_decap_8 FILLER_15_318 ();
 sg13g2_decap_8 FILLER_15_325 ();
 sg13g2_decap_8 FILLER_15_332 ();
 sg13g2_decap_8 FILLER_15_339 ();
 sg13g2_decap_8 FILLER_15_346 ();
 sg13g2_decap_8 FILLER_15_353 ();
 sg13g2_decap_8 FILLER_15_360 ();
 sg13g2_decap_8 FILLER_15_367 ();
 sg13g2_decap_8 FILLER_15_374 ();
 sg13g2_decap_8 FILLER_15_381 ();
 sg13g2_decap_8 FILLER_15_388 ();
 sg13g2_decap_8 FILLER_15_395 ();
 sg13g2_decap_8 FILLER_15_402 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_4 FILLER_16_112 ();
 sg13g2_fill_1 FILLER_16_142 ();
 sg13g2_fill_1 FILLER_16_206 ();
 sg13g2_decap_8 FILLER_16_241 ();
 sg13g2_decap_8 FILLER_16_248 ();
 sg13g2_decap_8 FILLER_16_255 ();
 sg13g2_decap_8 FILLER_16_262 ();
 sg13g2_decap_8 FILLER_16_269 ();
 sg13g2_decap_8 FILLER_16_276 ();
 sg13g2_decap_8 FILLER_16_283 ();
 sg13g2_decap_8 FILLER_16_290 ();
 sg13g2_decap_8 FILLER_16_297 ();
 sg13g2_decap_8 FILLER_16_304 ();
 sg13g2_decap_8 FILLER_16_311 ();
 sg13g2_decap_8 FILLER_16_318 ();
 sg13g2_decap_8 FILLER_16_325 ();
 sg13g2_decap_8 FILLER_16_332 ();
 sg13g2_decap_8 FILLER_16_339 ();
 sg13g2_decap_8 FILLER_16_346 ();
 sg13g2_decap_8 FILLER_16_353 ();
 sg13g2_decap_8 FILLER_16_360 ();
 sg13g2_decap_8 FILLER_16_367 ();
 sg13g2_decap_8 FILLER_16_374 ();
 sg13g2_decap_8 FILLER_16_381 ();
 sg13g2_decap_8 FILLER_16_388 ();
 sg13g2_decap_8 FILLER_16_395 ();
 sg13g2_decap_8 FILLER_16_402 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_fill_1 FILLER_17_119 ();
 sg13g2_fill_2 FILLER_17_173 ();
 sg13g2_fill_1 FILLER_17_175 ();
 sg13g2_fill_1 FILLER_17_202 ();
 sg13g2_decap_8 FILLER_17_233 ();
 sg13g2_decap_8 FILLER_17_240 ();
 sg13g2_decap_8 FILLER_17_247 ();
 sg13g2_decap_8 FILLER_17_254 ();
 sg13g2_decap_8 FILLER_17_261 ();
 sg13g2_decap_8 FILLER_17_268 ();
 sg13g2_decap_8 FILLER_17_275 ();
 sg13g2_decap_8 FILLER_17_282 ();
 sg13g2_decap_8 FILLER_17_289 ();
 sg13g2_decap_8 FILLER_17_296 ();
 sg13g2_decap_8 FILLER_17_303 ();
 sg13g2_decap_8 FILLER_17_310 ();
 sg13g2_decap_8 FILLER_17_317 ();
 sg13g2_decap_8 FILLER_17_324 ();
 sg13g2_decap_8 FILLER_17_331 ();
 sg13g2_decap_8 FILLER_17_338 ();
 sg13g2_decap_8 FILLER_17_345 ();
 sg13g2_decap_8 FILLER_17_352 ();
 sg13g2_decap_8 FILLER_17_359 ();
 sg13g2_decap_8 FILLER_17_366 ();
 sg13g2_decap_8 FILLER_17_373 ();
 sg13g2_decap_8 FILLER_17_380 ();
 sg13g2_decap_8 FILLER_17_387 ();
 sg13g2_decap_8 FILLER_17_394 ();
 sg13g2_decap_8 FILLER_17_401 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_4 FILLER_18_119 ();
 sg13g2_fill_1 FILLER_18_158 ();
 sg13g2_fill_1 FILLER_18_173 ();
 sg13g2_fill_1 FILLER_18_187 ();
 sg13g2_fill_1 FILLER_18_206 ();
 sg13g2_decap_8 FILLER_18_224 ();
 sg13g2_decap_8 FILLER_18_231 ();
 sg13g2_decap_8 FILLER_18_238 ();
 sg13g2_decap_8 FILLER_18_245 ();
 sg13g2_decap_8 FILLER_18_252 ();
 sg13g2_decap_8 FILLER_18_259 ();
 sg13g2_decap_8 FILLER_18_266 ();
 sg13g2_decap_8 FILLER_18_273 ();
 sg13g2_decap_8 FILLER_18_280 ();
 sg13g2_decap_8 FILLER_18_287 ();
 sg13g2_decap_8 FILLER_18_294 ();
 sg13g2_decap_8 FILLER_18_301 ();
 sg13g2_decap_8 FILLER_18_308 ();
 sg13g2_decap_8 FILLER_18_315 ();
 sg13g2_decap_8 FILLER_18_322 ();
 sg13g2_decap_8 FILLER_18_329 ();
 sg13g2_decap_8 FILLER_18_336 ();
 sg13g2_decap_8 FILLER_18_343 ();
 sg13g2_decap_8 FILLER_18_350 ();
 sg13g2_decap_8 FILLER_18_357 ();
 sg13g2_decap_8 FILLER_18_364 ();
 sg13g2_decap_8 FILLER_18_371 ();
 sg13g2_decap_8 FILLER_18_378 ();
 sg13g2_decap_8 FILLER_18_385 ();
 sg13g2_decap_8 FILLER_18_392 ();
 sg13g2_decap_8 FILLER_18_399 ();
 sg13g2_fill_2 FILLER_18_406 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_4 FILLER_19_112 ();
 sg13g2_fill_2 FILLER_19_116 ();
 sg13g2_fill_2 FILLER_19_148 ();
 sg13g2_fill_2 FILLER_19_165 ();
 sg13g2_fill_2 FILLER_19_174 ();
 sg13g2_fill_2 FILLER_19_198 ();
 sg13g2_decap_4 FILLER_19_209 ();
 sg13g2_decap_4 FILLER_19_216 ();
 sg13g2_fill_1 FILLER_19_220 ();
 sg13g2_decap_8 FILLER_19_231 ();
 sg13g2_decap_8 FILLER_19_238 ();
 sg13g2_decap_8 FILLER_19_245 ();
 sg13g2_decap_8 FILLER_19_252 ();
 sg13g2_decap_8 FILLER_19_259 ();
 sg13g2_decap_8 FILLER_19_266 ();
 sg13g2_decap_8 FILLER_19_273 ();
 sg13g2_decap_8 FILLER_19_280 ();
 sg13g2_decap_8 FILLER_19_287 ();
 sg13g2_decap_8 FILLER_19_294 ();
 sg13g2_decap_8 FILLER_19_301 ();
 sg13g2_decap_8 FILLER_19_308 ();
 sg13g2_decap_8 FILLER_19_315 ();
 sg13g2_decap_8 FILLER_19_322 ();
 sg13g2_decap_8 FILLER_19_329 ();
 sg13g2_decap_8 FILLER_19_336 ();
 sg13g2_decap_8 FILLER_19_343 ();
 sg13g2_decap_8 FILLER_19_350 ();
 sg13g2_decap_8 FILLER_19_357 ();
 sg13g2_decap_8 FILLER_19_364 ();
 sg13g2_decap_8 FILLER_19_371 ();
 sg13g2_decap_8 FILLER_19_378 ();
 sg13g2_decap_8 FILLER_19_385 ();
 sg13g2_decap_8 FILLER_19_392 ();
 sg13g2_decap_8 FILLER_19_399 ();
 sg13g2_fill_2 FILLER_19_406 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_4 FILLER_20_119 ();
 sg13g2_fill_1 FILLER_20_123 ();
 sg13g2_decap_8 FILLER_20_194 ();
 sg13g2_fill_2 FILLER_20_201 ();
 sg13g2_fill_1 FILLER_20_203 ();
 sg13g2_decap_8 FILLER_20_247 ();
 sg13g2_decap_8 FILLER_20_254 ();
 sg13g2_decap_8 FILLER_20_261 ();
 sg13g2_decap_8 FILLER_20_268 ();
 sg13g2_decap_8 FILLER_20_275 ();
 sg13g2_decap_8 FILLER_20_282 ();
 sg13g2_decap_8 FILLER_20_289 ();
 sg13g2_decap_8 FILLER_20_296 ();
 sg13g2_decap_8 FILLER_20_303 ();
 sg13g2_decap_8 FILLER_20_310 ();
 sg13g2_decap_8 FILLER_20_317 ();
 sg13g2_decap_8 FILLER_20_324 ();
 sg13g2_decap_8 FILLER_20_331 ();
 sg13g2_decap_8 FILLER_20_338 ();
 sg13g2_decap_8 FILLER_20_345 ();
 sg13g2_decap_8 FILLER_20_352 ();
 sg13g2_decap_8 FILLER_20_359 ();
 sg13g2_decap_8 FILLER_20_366 ();
 sg13g2_decap_8 FILLER_20_373 ();
 sg13g2_decap_8 FILLER_20_380 ();
 sg13g2_decap_8 FILLER_20_387 ();
 sg13g2_decap_8 FILLER_20_394 ();
 sg13g2_decap_8 FILLER_20_401 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_decap_8 FILLER_21_119 ();
 sg13g2_fill_1 FILLER_21_126 ();
 sg13g2_fill_2 FILLER_21_178 ();
 sg13g2_fill_2 FILLER_21_222 ();
 sg13g2_decap_8 FILLER_21_250 ();
 sg13g2_decap_8 FILLER_21_257 ();
 sg13g2_decap_8 FILLER_21_264 ();
 sg13g2_decap_8 FILLER_21_271 ();
 sg13g2_decap_8 FILLER_21_278 ();
 sg13g2_decap_8 FILLER_21_285 ();
 sg13g2_decap_8 FILLER_21_292 ();
 sg13g2_decap_8 FILLER_21_299 ();
 sg13g2_decap_8 FILLER_21_306 ();
 sg13g2_decap_8 FILLER_21_313 ();
 sg13g2_decap_8 FILLER_21_320 ();
 sg13g2_decap_8 FILLER_21_327 ();
 sg13g2_decap_8 FILLER_21_334 ();
 sg13g2_decap_8 FILLER_21_341 ();
 sg13g2_decap_8 FILLER_21_348 ();
 sg13g2_decap_8 FILLER_21_355 ();
 sg13g2_decap_8 FILLER_21_362 ();
 sg13g2_decap_8 FILLER_21_369 ();
 sg13g2_decap_8 FILLER_21_376 ();
 sg13g2_decap_8 FILLER_21_383 ();
 sg13g2_decap_8 FILLER_21_390 ();
 sg13g2_decap_8 FILLER_21_397 ();
 sg13g2_decap_4 FILLER_21_404 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_8 FILLER_22_105 ();
 sg13g2_decap_8 FILLER_22_112 ();
 sg13g2_fill_1 FILLER_22_159 ();
 sg13g2_fill_2 FILLER_22_223 ();
 sg13g2_decap_8 FILLER_22_260 ();
 sg13g2_decap_8 FILLER_22_267 ();
 sg13g2_decap_8 FILLER_22_274 ();
 sg13g2_decap_8 FILLER_22_281 ();
 sg13g2_decap_8 FILLER_22_288 ();
 sg13g2_decap_8 FILLER_22_295 ();
 sg13g2_decap_8 FILLER_22_302 ();
 sg13g2_decap_8 FILLER_22_309 ();
 sg13g2_decap_8 FILLER_22_316 ();
 sg13g2_decap_8 FILLER_22_323 ();
 sg13g2_decap_8 FILLER_22_330 ();
 sg13g2_decap_8 FILLER_22_337 ();
 sg13g2_decap_8 FILLER_22_344 ();
 sg13g2_decap_8 FILLER_22_351 ();
 sg13g2_decap_8 FILLER_22_358 ();
 sg13g2_decap_8 FILLER_22_365 ();
 sg13g2_decap_8 FILLER_22_372 ();
 sg13g2_decap_8 FILLER_22_379 ();
 sg13g2_decap_8 FILLER_22_386 ();
 sg13g2_decap_8 FILLER_22_393 ();
 sg13g2_decap_8 FILLER_22_400 ();
 sg13g2_fill_2 FILLER_22_407 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_98 ();
 sg13g2_fill_2 FILLER_23_105 ();
 sg13g2_fill_1 FILLER_23_107 ();
 sg13g2_fill_1 FILLER_23_138 ();
 sg13g2_decap_4 FILLER_23_151 ();
 sg13g2_fill_2 FILLER_23_187 ();
 sg13g2_fill_1 FILLER_23_189 ();
 sg13g2_fill_1 FILLER_23_226 ();
 sg13g2_decap_8 FILLER_23_270 ();
 sg13g2_decap_8 FILLER_23_277 ();
 sg13g2_decap_8 FILLER_23_284 ();
 sg13g2_decap_8 FILLER_23_291 ();
 sg13g2_decap_8 FILLER_23_298 ();
 sg13g2_decap_8 FILLER_23_305 ();
 sg13g2_decap_8 FILLER_23_312 ();
 sg13g2_decap_8 FILLER_23_319 ();
 sg13g2_decap_8 FILLER_23_326 ();
 sg13g2_decap_8 FILLER_23_333 ();
 sg13g2_decap_8 FILLER_23_340 ();
 sg13g2_decap_8 FILLER_23_347 ();
 sg13g2_decap_8 FILLER_23_354 ();
 sg13g2_decap_8 FILLER_23_361 ();
 sg13g2_decap_8 FILLER_23_368 ();
 sg13g2_decap_8 FILLER_23_375 ();
 sg13g2_decap_8 FILLER_23_382 ();
 sg13g2_decap_8 FILLER_23_389 ();
 sg13g2_decap_8 FILLER_23_396 ();
 sg13g2_decap_4 FILLER_23_403 ();
 sg13g2_fill_2 FILLER_23_407 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_fill_2 FILLER_24_107 ();
 sg13g2_fill_1 FILLER_24_109 ();
 sg13g2_fill_1 FILLER_24_118 ();
 sg13g2_fill_1 FILLER_24_138 ();
 sg13g2_fill_1 FILLER_24_169 ();
 sg13g2_fill_2 FILLER_24_193 ();
 sg13g2_fill_2 FILLER_24_215 ();
 sg13g2_fill_1 FILLER_24_217 ();
 sg13g2_fill_1 FILLER_24_231 ();
 sg13g2_decap_8 FILLER_24_265 ();
 sg13g2_decap_8 FILLER_24_272 ();
 sg13g2_decap_8 FILLER_24_279 ();
 sg13g2_decap_8 FILLER_24_286 ();
 sg13g2_decap_8 FILLER_24_293 ();
 sg13g2_decap_8 FILLER_24_300 ();
 sg13g2_decap_8 FILLER_24_307 ();
 sg13g2_decap_8 FILLER_24_314 ();
 sg13g2_decap_8 FILLER_24_321 ();
 sg13g2_decap_8 FILLER_24_328 ();
 sg13g2_decap_8 FILLER_24_335 ();
 sg13g2_decap_8 FILLER_24_342 ();
 sg13g2_decap_8 FILLER_24_349 ();
 sg13g2_decap_8 FILLER_24_356 ();
 sg13g2_decap_8 FILLER_24_363 ();
 sg13g2_decap_8 FILLER_24_370 ();
 sg13g2_decap_8 FILLER_24_377 ();
 sg13g2_decap_8 FILLER_24_384 ();
 sg13g2_decap_8 FILLER_24_391 ();
 sg13g2_decap_8 FILLER_24_398 ();
 sg13g2_decap_4 FILLER_24_405 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_fill_1 FILLER_25_170 ();
 sg13g2_fill_2 FILLER_25_197 ();
 sg13g2_fill_1 FILLER_25_225 ();
 sg13g2_fill_1 FILLER_25_234 ();
 sg13g2_decap_8 FILLER_25_266 ();
 sg13g2_decap_8 FILLER_25_273 ();
 sg13g2_decap_8 FILLER_25_280 ();
 sg13g2_decap_8 FILLER_25_287 ();
 sg13g2_decap_8 FILLER_25_294 ();
 sg13g2_decap_8 FILLER_25_301 ();
 sg13g2_decap_8 FILLER_25_308 ();
 sg13g2_decap_8 FILLER_25_315 ();
 sg13g2_decap_8 FILLER_25_322 ();
 sg13g2_decap_8 FILLER_25_329 ();
 sg13g2_decap_8 FILLER_25_336 ();
 sg13g2_decap_8 FILLER_25_343 ();
 sg13g2_decap_8 FILLER_25_350 ();
 sg13g2_decap_8 FILLER_25_357 ();
 sg13g2_decap_8 FILLER_25_364 ();
 sg13g2_decap_8 FILLER_25_371 ();
 sg13g2_decap_8 FILLER_25_378 ();
 sg13g2_decap_8 FILLER_25_385 ();
 sg13g2_decap_8 FILLER_25_392 ();
 sg13g2_decap_8 FILLER_25_399 ();
 sg13g2_fill_2 FILLER_25_406 ();
 sg13g2_fill_1 FILLER_25_408 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_4 FILLER_26_70 ();
 sg13g2_fill_1 FILLER_26_126 ();
 sg13g2_fill_2 FILLER_26_153 ();
 sg13g2_fill_2 FILLER_26_159 ();
 sg13g2_fill_2 FILLER_26_166 ();
 sg13g2_fill_1 FILLER_26_172 ();
 sg13g2_fill_1 FILLER_26_202 ();
 sg13g2_fill_2 FILLER_26_226 ();
 sg13g2_decap_8 FILLER_26_269 ();
 sg13g2_decap_8 FILLER_26_276 ();
 sg13g2_decap_8 FILLER_26_283 ();
 sg13g2_decap_8 FILLER_26_290 ();
 sg13g2_decap_8 FILLER_26_297 ();
 sg13g2_decap_8 FILLER_26_304 ();
 sg13g2_decap_8 FILLER_26_311 ();
 sg13g2_decap_8 FILLER_26_318 ();
 sg13g2_decap_8 FILLER_26_325 ();
 sg13g2_decap_8 FILLER_26_332 ();
 sg13g2_decap_8 FILLER_26_339 ();
 sg13g2_decap_8 FILLER_26_346 ();
 sg13g2_decap_8 FILLER_26_353 ();
 sg13g2_decap_8 FILLER_26_360 ();
 sg13g2_decap_8 FILLER_26_367 ();
 sg13g2_decap_8 FILLER_26_374 ();
 sg13g2_decap_8 FILLER_26_381 ();
 sg13g2_decap_8 FILLER_26_388 ();
 sg13g2_decap_8 FILLER_26_395 ();
 sg13g2_decap_8 FILLER_26_402 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_fill_1 FILLER_27_63 ();
 sg13g2_fill_2 FILLER_27_72 ();
 sg13g2_fill_1 FILLER_27_74 ();
 sg13g2_fill_2 FILLER_27_140 ();
 sg13g2_fill_1 FILLER_27_164 ();
 sg13g2_fill_1 FILLER_27_203 ();
 sg13g2_fill_1 FILLER_27_234 ();
 sg13g2_decap_8 FILLER_27_265 ();
 sg13g2_decap_8 FILLER_27_272 ();
 sg13g2_decap_8 FILLER_27_279 ();
 sg13g2_decap_8 FILLER_27_286 ();
 sg13g2_decap_8 FILLER_27_293 ();
 sg13g2_decap_8 FILLER_27_300 ();
 sg13g2_decap_8 FILLER_27_307 ();
 sg13g2_decap_8 FILLER_27_314 ();
 sg13g2_decap_8 FILLER_27_321 ();
 sg13g2_decap_8 FILLER_27_328 ();
 sg13g2_decap_8 FILLER_27_335 ();
 sg13g2_decap_8 FILLER_27_342 ();
 sg13g2_decap_8 FILLER_27_349 ();
 sg13g2_decap_8 FILLER_27_356 ();
 sg13g2_decap_8 FILLER_27_363 ();
 sg13g2_decap_8 FILLER_27_370 ();
 sg13g2_decap_8 FILLER_27_377 ();
 sg13g2_decap_8 FILLER_27_384 ();
 sg13g2_decap_8 FILLER_27_391 ();
 sg13g2_decap_8 FILLER_27_398 ();
 sg13g2_decap_4 FILLER_27_405 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_fill_2 FILLER_28_56 ();
 sg13g2_fill_1 FILLER_28_58 ();
 sg13g2_fill_2 FILLER_28_196 ();
 sg13g2_fill_1 FILLER_28_198 ();
 sg13g2_decap_8 FILLER_28_269 ();
 sg13g2_decap_8 FILLER_28_276 ();
 sg13g2_decap_8 FILLER_28_283 ();
 sg13g2_decap_8 FILLER_28_290 ();
 sg13g2_decap_8 FILLER_28_297 ();
 sg13g2_decap_8 FILLER_28_304 ();
 sg13g2_decap_8 FILLER_28_311 ();
 sg13g2_decap_8 FILLER_28_318 ();
 sg13g2_decap_8 FILLER_28_325 ();
 sg13g2_decap_8 FILLER_28_332 ();
 sg13g2_decap_8 FILLER_28_339 ();
 sg13g2_decap_8 FILLER_28_346 ();
 sg13g2_decap_8 FILLER_28_353 ();
 sg13g2_decap_8 FILLER_28_360 ();
 sg13g2_decap_8 FILLER_28_367 ();
 sg13g2_decap_8 FILLER_28_374 ();
 sg13g2_decap_8 FILLER_28_381 ();
 sg13g2_decap_8 FILLER_28_388 ();
 sg13g2_decap_8 FILLER_28_395 ();
 sg13g2_decap_8 FILLER_28_402 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_fill_2 FILLER_29_93 ();
 sg13g2_fill_1 FILLER_29_95 ();
 sg13g2_fill_2 FILLER_29_105 ();
 sg13g2_fill_1 FILLER_29_107 ();
 sg13g2_fill_1 FILLER_29_117 ();
 sg13g2_fill_2 FILLER_29_174 ();
 sg13g2_fill_2 FILLER_29_214 ();
 sg13g2_fill_1 FILLER_29_247 ();
 sg13g2_decap_8 FILLER_29_278 ();
 sg13g2_decap_8 FILLER_29_285 ();
 sg13g2_decap_8 FILLER_29_292 ();
 sg13g2_decap_8 FILLER_29_299 ();
 sg13g2_decap_8 FILLER_29_306 ();
 sg13g2_decap_8 FILLER_29_313 ();
 sg13g2_decap_8 FILLER_29_320 ();
 sg13g2_decap_8 FILLER_29_327 ();
 sg13g2_decap_8 FILLER_29_334 ();
 sg13g2_decap_8 FILLER_29_341 ();
 sg13g2_decap_8 FILLER_29_348 ();
 sg13g2_decap_8 FILLER_29_355 ();
 sg13g2_decap_8 FILLER_29_362 ();
 sg13g2_decap_8 FILLER_29_369 ();
 sg13g2_decap_8 FILLER_29_376 ();
 sg13g2_decap_8 FILLER_29_383 ();
 sg13g2_decap_8 FILLER_29_390 ();
 sg13g2_decap_8 FILLER_29_397 ();
 sg13g2_decap_4 FILLER_29_404 ();
 sg13g2_fill_1 FILLER_29_408 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_4 FILLER_30_49 ();
 sg13g2_fill_1 FILLER_30_187 ();
 sg13g2_fill_1 FILLER_30_199 ();
 sg13g2_fill_2 FILLER_30_269 ();
 sg13g2_fill_1 FILLER_30_271 ();
 sg13g2_fill_1 FILLER_30_281 ();
 sg13g2_decap_4 FILLER_30_288 ();
 sg13g2_fill_1 FILLER_30_292 ();
 sg13g2_decap_8 FILLER_30_297 ();
 sg13g2_decap_8 FILLER_30_304 ();
 sg13g2_decap_8 FILLER_30_311 ();
 sg13g2_decap_8 FILLER_30_318 ();
 sg13g2_decap_8 FILLER_30_325 ();
 sg13g2_decap_8 FILLER_30_332 ();
 sg13g2_decap_8 FILLER_30_339 ();
 sg13g2_decap_8 FILLER_30_346 ();
 sg13g2_decap_8 FILLER_30_353 ();
 sg13g2_decap_8 FILLER_30_360 ();
 sg13g2_decap_8 FILLER_30_367 ();
 sg13g2_decap_8 FILLER_30_374 ();
 sg13g2_decap_8 FILLER_30_381 ();
 sg13g2_decap_8 FILLER_30_388 ();
 sg13g2_decap_8 FILLER_30_395 ();
 sg13g2_decap_8 FILLER_30_402 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_fill_2 FILLER_31_56 ();
 sg13g2_fill_1 FILLER_31_71 ();
 sg13g2_fill_1 FILLER_31_202 ();
 sg13g2_fill_1 FILLER_31_237 ();
 sg13g2_fill_1 FILLER_31_252 ();
 sg13g2_fill_2 FILLER_31_297 ();
 sg13g2_decap_8 FILLER_31_319 ();
 sg13g2_decap_8 FILLER_31_326 ();
 sg13g2_decap_8 FILLER_31_333 ();
 sg13g2_decap_8 FILLER_31_340 ();
 sg13g2_decap_8 FILLER_31_347 ();
 sg13g2_decap_8 FILLER_31_354 ();
 sg13g2_decap_8 FILLER_31_361 ();
 sg13g2_decap_8 FILLER_31_368 ();
 sg13g2_decap_8 FILLER_31_375 ();
 sg13g2_decap_8 FILLER_31_382 ();
 sg13g2_decap_8 FILLER_31_389 ();
 sg13g2_decap_8 FILLER_31_396 ();
 sg13g2_decap_4 FILLER_31_403 ();
 sg13g2_fill_2 FILLER_31_407 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_4 FILLER_32_49 ();
 sg13g2_fill_1 FILLER_32_53 ();
 sg13g2_fill_1 FILLER_32_106 ();
 sg13g2_fill_1 FILLER_32_115 ();
 sg13g2_fill_2 FILLER_32_220 ();
 sg13g2_fill_2 FILLER_32_248 ();
 sg13g2_fill_1 FILLER_32_250 ();
 sg13g2_fill_2 FILLER_32_263 ();
 sg13g2_fill_1 FILLER_32_265 ();
 sg13g2_decap_8 FILLER_32_332 ();
 sg13g2_decap_8 FILLER_32_339 ();
 sg13g2_decap_8 FILLER_32_346 ();
 sg13g2_decap_8 FILLER_32_353 ();
 sg13g2_decap_8 FILLER_32_360 ();
 sg13g2_decap_8 FILLER_32_367 ();
 sg13g2_decap_8 FILLER_32_374 ();
 sg13g2_decap_8 FILLER_32_381 ();
 sg13g2_decap_8 FILLER_32_388 ();
 sg13g2_decap_8 FILLER_32_395 ();
 sg13g2_decap_8 FILLER_32_402 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_fill_1 FILLER_33_70 ();
 sg13g2_fill_1 FILLER_33_75 ();
 sg13g2_fill_2 FILLER_33_98 ();
 sg13g2_fill_2 FILLER_33_142 ();
 sg13g2_fill_2 FILLER_33_303 ();
 sg13g2_fill_1 FILLER_33_305 ();
 sg13g2_decap_8 FILLER_33_330 ();
 sg13g2_decap_8 FILLER_33_337 ();
 sg13g2_decap_8 FILLER_33_344 ();
 sg13g2_decap_8 FILLER_33_351 ();
 sg13g2_decap_8 FILLER_33_358 ();
 sg13g2_decap_8 FILLER_33_365 ();
 sg13g2_decap_8 FILLER_33_372 ();
 sg13g2_decap_8 FILLER_33_379 ();
 sg13g2_decap_8 FILLER_33_386 ();
 sg13g2_decap_8 FILLER_33_393 ();
 sg13g2_decap_8 FILLER_33_400 ();
 sg13g2_fill_2 FILLER_33_407 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_fill_1 FILLER_34_87 ();
 sg13g2_fill_1 FILLER_34_109 ();
 sg13g2_fill_2 FILLER_34_136 ();
 sg13g2_fill_2 FILLER_34_146 ();
 sg13g2_fill_1 FILLER_34_177 ();
 sg13g2_decap_8 FILLER_34_284 ();
 sg13g2_decap_4 FILLER_34_291 ();
 sg13g2_fill_1 FILLER_34_295 ();
 sg13g2_decap_4 FILLER_34_313 ();
 sg13g2_fill_1 FILLER_34_317 ();
 sg13g2_decap_8 FILLER_34_322 ();
 sg13g2_decap_8 FILLER_34_329 ();
 sg13g2_decap_8 FILLER_34_336 ();
 sg13g2_decap_8 FILLER_34_343 ();
 sg13g2_decap_8 FILLER_34_350 ();
 sg13g2_decap_8 FILLER_34_357 ();
 sg13g2_decap_8 FILLER_34_364 ();
 sg13g2_decap_8 FILLER_34_371 ();
 sg13g2_decap_8 FILLER_34_378 ();
 sg13g2_decap_8 FILLER_34_385 ();
 sg13g2_decap_8 FILLER_34_392 ();
 sg13g2_decap_8 FILLER_34_399 ();
 sg13g2_fill_2 FILLER_34_406 ();
 sg13g2_fill_1 FILLER_34_408 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_fill_1 FILLER_35_132 ();
 sg13g2_fill_1 FILLER_35_147 ();
 sg13g2_fill_2 FILLER_35_165 ();
 sg13g2_decap_4 FILLER_35_275 ();
 sg13g2_fill_2 FILLER_35_311 ();
 sg13g2_fill_1 FILLER_35_313 ();
 sg13g2_decap_8 FILLER_35_332 ();
 sg13g2_decap_8 FILLER_35_339 ();
 sg13g2_decap_8 FILLER_35_346 ();
 sg13g2_decap_8 FILLER_35_353 ();
 sg13g2_decap_8 FILLER_35_360 ();
 sg13g2_decap_8 FILLER_35_367 ();
 sg13g2_decap_8 FILLER_35_374 ();
 sg13g2_decap_8 FILLER_35_381 ();
 sg13g2_decap_8 FILLER_35_388 ();
 sg13g2_decap_8 FILLER_35_395 ();
 sg13g2_decap_8 FILLER_35_402 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_fill_2 FILLER_36_49 ();
 sg13g2_fill_1 FILLER_36_85 ();
 sg13g2_fill_2 FILLER_36_121 ();
 sg13g2_fill_1 FILLER_36_123 ();
 sg13g2_fill_1 FILLER_36_131 ();
 sg13g2_fill_1 FILLER_36_214 ();
 sg13g2_decap_4 FILLER_36_270 ();
 sg13g2_fill_1 FILLER_36_280 ();
 sg13g2_fill_2 FILLER_36_293 ();
 sg13g2_fill_1 FILLER_36_295 ();
 sg13g2_decap_8 FILLER_36_338 ();
 sg13g2_decap_8 FILLER_36_345 ();
 sg13g2_decap_8 FILLER_36_352 ();
 sg13g2_decap_8 FILLER_36_359 ();
 sg13g2_decap_8 FILLER_36_366 ();
 sg13g2_decap_8 FILLER_36_373 ();
 sg13g2_decap_8 FILLER_36_380 ();
 sg13g2_decap_8 FILLER_36_387 ();
 sg13g2_decap_8 FILLER_36_394 ();
 sg13g2_decap_8 FILLER_36_401 ();
 sg13g2_fill_1 FILLER_36_408 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_4 FILLER_37_56 ();
 sg13g2_fill_1 FILLER_37_94 ();
 sg13g2_fill_2 FILLER_37_131 ();
 sg13g2_fill_1 FILLER_37_133 ();
 sg13g2_fill_2 FILLER_37_139 ();
 sg13g2_fill_1 FILLER_37_163 ();
 sg13g2_fill_1 FILLER_37_173 ();
 sg13g2_fill_1 FILLER_37_244 ();
 sg13g2_decap_8 FILLER_37_337 ();
 sg13g2_decap_8 FILLER_37_344 ();
 sg13g2_decap_8 FILLER_37_351 ();
 sg13g2_decap_8 FILLER_37_358 ();
 sg13g2_decap_8 FILLER_37_365 ();
 sg13g2_decap_8 FILLER_37_372 ();
 sg13g2_decap_8 FILLER_37_379 ();
 sg13g2_decap_8 FILLER_37_386 ();
 sg13g2_decap_8 FILLER_37_393 ();
 sg13g2_decap_8 FILLER_37_400 ();
 sg13g2_fill_2 FILLER_37_407 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_8 FILLER_38_56 ();
 sg13g2_decap_8 FILLER_38_63 ();
 sg13g2_decap_4 FILLER_38_70 ();
 sg13g2_fill_1 FILLER_38_74 ();
 sg13g2_decap_4 FILLER_38_93 ();
 sg13g2_fill_1 FILLER_38_97 ();
 sg13g2_decap_4 FILLER_38_102 ();
 sg13g2_fill_2 FILLER_38_106 ();
 sg13g2_decap_8 FILLER_38_126 ();
 sg13g2_fill_2 FILLER_38_133 ();
 sg13g2_fill_1 FILLER_38_135 ();
 sg13g2_fill_2 FILLER_38_179 ();
 sg13g2_fill_2 FILLER_38_197 ();
 sg13g2_fill_1 FILLER_38_270 ();
 sg13g2_fill_2 FILLER_38_288 ();
 sg13g2_fill_1 FILLER_38_290 ();
 sg13g2_fill_2 FILLER_38_295 ();
 sg13g2_fill_1 FILLER_38_297 ();
 sg13g2_fill_2 FILLER_38_321 ();
 sg13g2_decap_8 FILLER_38_344 ();
 sg13g2_decap_8 FILLER_38_351 ();
 sg13g2_decap_8 FILLER_38_358 ();
 sg13g2_decap_8 FILLER_38_365 ();
 sg13g2_decap_8 FILLER_38_372 ();
 sg13g2_decap_8 FILLER_38_379 ();
 sg13g2_decap_8 FILLER_38_386 ();
 sg13g2_decap_8 FILLER_38_393 ();
 sg13g2_decap_8 FILLER_38_400 ();
 sg13g2_fill_2 FILLER_38_407 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_14 ();
 sg13g2_decap_8 FILLER_39_21 ();
 sg13g2_decap_8 FILLER_39_28 ();
 sg13g2_decap_8 FILLER_39_35 ();
 sg13g2_decap_8 FILLER_39_42 ();
 sg13g2_decap_8 FILLER_39_49 ();
 sg13g2_decap_8 FILLER_39_56 ();
 sg13g2_decap_8 FILLER_39_63 ();
 sg13g2_decap_4 FILLER_39_70 ();
 sg13g2_fill_1 FILLER_39_74 ();
 sg13g2_decap_8 FILLER_39_79 ();
 sg13g2_decap_8 FILLER_39_90 ();
 sg13g2_decap_8 FILLER_39_97 ();
 sg13g2_decap_8 FILLER_39_104 ();
 sg13g2_fill_2 FILLER_39_111 ();
 sg13g2_fill_1 FILLER_39_173 ();
 sg13g2_fill_1 FILLER_39_184 ();
 sg13g2_decap_8 FILLER_39_190 ();
 sg13g2_decap_8 FILLER_39_197 ();
 sg13g2_decap_4 FILLER_39_204 ();
 sg13g2_fill_2 FILLER_39_208 ();
 sg13g2_fill_1 FILLER_39_214 ();
 sg13g2_fill_1 FILLER_39_219 ();
 sg13g2_decap_8 FILLER_39_262 ();
 sg13g2_fill_2 FILLER_39_269 ();
 sg13g2_fill_1 FILLER_39_271 ();
 sg13g2_fill_2 FILLER_39_295 ();
 sg13g2_fill_2 FILLER_39_305 ();
 sg13g2_decap_8 FILLER_39_351 ();
 sg13g2_decap_8 FILLER_39_358 ();
 sg13g2_decap_8 FILLER_39_365 ();
 sg13g2_decap_8 FILLER_39_372 ();
 sg13g2_decap_8 FILLER_39_379 ();
 sg13g2_decap_8 FILLER_39_386 ();
 sg13g2_decap_8 FILLER_39_393 ();
 sg13g2_decap_8 FILLER_39_400 ();
 sg13g2_fill_2 FILLER_39_407 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_14 ();
 sg13g2_decap_8 FILLER_40_21 ();
 sg13g2_decap_8 FILLER_40_28 ();
 sg13g2_decap_8 FILLER_40_35 ();
 sg13g2_decap_8 FILLER_40_42 ();
 sg13g2_decap_8 FILLER_40_49 ();
 sg13g2_decap_4 FILLER_40_56 ();
 sg13g2_fill_2 FILLER_40_94 ();
 sg13g2_decap_8 FILLER_40_107 ();
 sg13g2_fill_2 FILLER_40_152 ();
 sg13g2_fill_1 FILLER_40_175 ();
 sg13g2_fill_1 FILLER_40_190 ();
 sg13g2_decap_8 FILLER_40_201 ();
 sg13g2_decap_4 FILLER_40_208 ();
 sg13g2_fill_2 FILLER_40_212 ();
 sg13g2_decap_8 FILLER_40_222 ();
 sg13g2_decap_8 FILLER_40_229 ();
 sg13g2_decap_8 FILLER_40_236 ();
 sg13g2_decap_8 FILLER_40_243 ();
 sg13g2_fill_1 FILLER_40_250 ();
 sg13g2_decap_8 FILLER_40_261 ();
 sg13g2_fill_2 FILLER_40_268 ();
 sg13g2_fill_1 FILLER_40_270 ();
 sg13g2_fill_1 FILLER_40_280 ();
 sg13g2_decap_4 FILLER_40_287 ();
 sg13g2_fill_2 FILLER_40_295 ();
 sg13g2_decap_4 FILLER_40_309 ();
 sg13g2_decap_8 FILLER_40_318 ();
 sg13g2_decap_4 FILLER_40_325 ();
 sg13g2_decap_8 FILLER_40_340 ();
 sg13g2_decap_8 FILLER_40_347 ();
 sg13g2_decap_8 FILLER_40_354 ();
 sg13g2_decap_8 FILLER_40_361 ();
 sg13g2_decap_8 FILLER_40_368 ();
 sg13g2_decap_8 FILLER_40_375 ();
 sg13g2_decap_8 FILLER_40_382 ();
 sg13g2_decap_8 FILLER_40_389 ();
 sg13g2_decap_8 FILLER_40_396 ();
 sg13g2_decap_4 FILLER_40_403 ();
 sg13g2_fill_2 FILLER_40_407 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_8 FILLER_41_14 ();
 sg13g2_decap_8 FILLER_41_21 ();
 sg13g2_decap_8 FILLER_41_28 ();
 sg13g2_decap_8 FILLER_41_35 ();
 sg13g2_decap_8 FILLER_41_42 ();
 sg13g2_decap_4 FILLER_41_49 ();
 sg13g2_fill_2 FILLER_41_116 ();
 sg13g2_decap_4 FILLER_41_198 ();
 sg13g2_fill_1 FILLER_41_202 ();
 sg13g2_decap_8 FILLER_41_207 ();
 sg13g2_decap_8 FILLER_41_214 ();
 sg13g2_decap_8 FILLER_41_221 ();
 sg13g2_fill_2 FILLER_41_228 ();
 sg13g2_fill_1 FILLER_41_230 ();
 sg13g2_fill_2 FILLER_41_295 ();
 sg13g2_fill_2 FILLER_41_309 ();
 sg13g2_fill_2 FILLER_41_323 ();
 sg13g2_decap_8 FILLER_41_337 ();
 sg13g2_decap_8 FILLER_41_344 ();
 sg13g2_decap_8 FILLER_41_351 ();
 sg13g2_decap_8 FILLER_41_358 ();
 sg13g2_decap_8 FILLER_41_365 ();
 sg13g2_decap_8 FILLER_41_372 ();
 sg13g2_decap_8 FILLER_41_379 ();
 sg13g2_decap_8 FILLER_41_386 ();
 sg13g2_decap_8 FILLER_41_393 ();
 sg13g2_decap_8 FILLER_41_400 ();
 sg13g2_fill_2 FILLER_41_407 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_decap_8 FILLER_42_14 ();
 sg13g2_decap_8 FILLER_42_21 ();
 sg13g2_decap_8 FILLER_42_28 ();
 sg13g2_decap_8 FILLER_42_35 ();
 sg13g2_decap_4 FILLER_42_42 ();
 sg13g2_fill_2 FILLER_42_46 ();
 sg13g2_fill_1 FILLER_42_74 ();
 sg13g2_fill_2 FILLER_42_92 ();
 sg13g2_fill_1 FILLER_42_94 ();
 sg13g2_fill_2 FILLER_42_120 ();
 sg13g2_fill_2 FILLER_42_145 ();
 sg13g2_fill_1 FILLER_42_147 ();
 sg13g2_fill_1 FILLER_42_163 ();
 sg13g2_decap_4 FILLER_42_179 ();
 sg13g2_decap_4 FILLER_42_187 ();
 sg13g2_fill_1 FILLER_42_191 ();
 sg13g2_fill_2 FILLER_42_223 ();
 sg13g2_fill_2 FILLER_42_230 ();
 sg13g2_fill_1 FILLER_42_252 ();
 sg13g2_fill_2 FILLER_42_270 ();
 sg13g2_fill_1 FILLER_42_272 ();
 sg13g2_fill_2 FILLER_42_313 ();
 sg13g2_fill_1 FILLER_42_315 ();
 sg13g2_fill_2 FILLER_42_327 ();
 sg13g2_fill_1 FILLER_42_329 ();
 sg13g2_decap_8 FILLER_42_355 ();
 sg13g2_decap_8 FILLER_42_362 ();
 sg13g2_decap_8 FILLER_42_369 ();
 sg13g2_decap_8 FILLER_42_376 ();
 sg13g2_decap_8 FILLER_42_383 ();
 sg13g2_decap_8 FILLER_42_390 ();
 sg13g2_decap_8 FILLER_42_397 ();
 sg13g2_decap_4 FILLER_42_404 ();
 sg13g2_fill_1 FILLER_42_408 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_decap_8 FILLER_43_14 ();
 sg13g2_decap_8 FILLER_43_21 ();
 sg13g2_decap_8 FILLER_43_28 ();
 sg13g2_decap_8 FILLER_43_35 ();
 sg13g2_decap_8 FILLER_43_42 ();
 sg13g2_decap_8 FILLER_43_49 ();
 sg13g2_fill_2 FILLER_43_56 ();
 sg13g2_fill_1 FILLER_43_58 ();
 sg13g2_fill_2 FILLER_43_85 ();
 sg13g2_fill_1 FILLER_43_103 ();
 sg13g2_fill_2 FILLER_43_111 ();
 sg13g2_decap_4 FILLER_43_128 ();
 sg13g2_fill_1 FILLER_43_132 ();
 sg13g2_fill_1 FILLER_43_160 ();
 sg13g2_decap_4 FILLER_43_173 ();
 sg13g2_decap_4 FILLER_43_186 ();
 sg13g2_fill_1 FILLER_43_224 ();
 sg13g2_fill_2 FILLER_43_242 ();
 sg13g2_fill_1 FILLER_43_244 ();
 sg13g2_decap_4 FILLER_43_270 ();
 sg13g2_fill_2 FILLER_43_274 ();
 sg13g2_decap_4 FILLER_43_282 ();
 sg13g2_fill_2 FILLER_43_294 ();
 sg13g2_fill_1 FILLER_43_296 ();
 sg13g2_decap_4 FILLER_43_333 ();
 sg13g2_decap_8 FILLER_43_358 ();
 sg13g2_decap_8 FILLER_43_365 ();
 sg13g2_decap_8 FILLER_43_372 ();
 sg13g2_decap_8 FILLER_43_379 ();
 sg13g2_decap_8 FILLER_43_386 ();
 sg13g2_decap_8 FILLER_43_393 ();
 sg13g2_decap_8 FILLER_43_400 ();
 sg13g2_fill_2 FILLER_43_407 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_decap_8 FILLER_44_14 ();
 sg13g2_decap_8 FILLER_44_21 ();
 sg13g2_decap_8 FILLER_44_28 ();
 sg13g2_decap_8 FILLER_44_35 ();
 sg13g2_decap_8 FILLER_44_42 ();
 sg13g2_decap_8 FILLER_44_49 ();
 sg13g2_decap_4 FILLER_44_56 ();
 sg13g2_fill_1 FILLER_44_60 ();
 sg13g2_fill_1 FILLER_44_88 ();
 sg13g2_fill_2 FILLER_44_94 ();
 sg13g2_fill_1 FILLER_44_96 ();
 sg13g2_fill_1 FILLER_44_104 ();
 sg13g2_fill_1 FILLER_44_161 ();
 sg13g2_fill_1 FILLER_44_172 ();
 sg13g2_fill_2 FILLER_44_196 ();
 sg13g2_fill_2 FILLER_44_224 ();
 sg13g2_fill_2 FILLER_44_240 ();
 sg13g2_fill_2 FILLER_44_247 ();
 sg13g2_decap_4 FILLER_44_261 ();
 sg13g2_fill_2 FILLER_44_265 ();
 sg13g2_fill_1 FILLER_44_277 ();
 sg13g2_decap_4 FILLER_44_306 ();
 sg13g2_fill_1 FILLER_44_310 ();
 sg13g2_fill_1 FILLER_44_316 ();
 sg13g2_fill_1 FILLER_44_341 ();
 sg13g2_decap_8 FILLER_44_364 ();
 sg13g2_decap_8 FILLER_44_371 ();
 sg13g2_decap_8 FILLER_44_378 ();
 sg13g2_decap_8 FILLER_44_385 ();
 sg13g2_decap_8 FILLER_44_392 ();
 sg13g2_decap_8 FILLER_44_399 ();
 sg13g2_fill_2 FILLER_44_406 ();
 sg13g2_fill_1 FILLER_44_408 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_7 ();
 sg13g2_decap_8 FILLER_45_14 ();
 sg13g2_decap_8 FILLER_45_21 ();
 sg13g2_decap_8 FILLER_45_28 ();
 sg13g2_decap_8 FILLER_45_35 ();
 sg13g2_decap_8 FILLER_45_42 ();
 sg13g2_fill_2 FILLER_45_49 ();
 sg13g2_fill_1 FILLER_45_97 ();
 sg13g2_fill_2 FILLER_45_108 ();
 sg13g2_fill_1 FILLER_45_110 ();
 sg13g2_fill_2 FILLER_45_134 ();
 sg13g2_fill_1 FILLER_45_136 ();
 sg13g2_fill_2 FILLER_45_184 ();
 sg13g2_decap_8 FILLER_45_201 ();
 sg13g2_fill_1 FILLER_45_208 ();
 sg13g2_decap_8 FILLER_45_213 ();
 sg13g2_decap_8 FILLER_45_220 ();
 sg13g2_decap_4 FILLER_45_231 ();
 sg13g2_fill_2 FILLER_45_252 ();
 sg13g2_fill_1 FILLER_45_254 ();
 sg13g2_fill_1 FILLER_45_288 ();
 sg13g2_fill_2 FILLER_45_295 ();
 sg13g2_fill_2 FILLER_45_301 ();
 sg13g2_fill_1 FILLER_45_303 ();
 sg13g2_fill_2 FILLER_45_316 ();
 sg13g2_fill_1 FILLER_45_318 ();
 sg13g2_decap_4 FILLER_45_325 ();
 sg13g2_fill_1 FILLER_45_329 ();
 sg13g2_decap_8 FILLER_45_353 ();
 sg13g2_decap_8 FILLER_45_360 ();
 sg13g2_decap_8 FILLER_45_367 ();
 sg13g2_decap_8 FILLER_45_374 ();
 sg13g2_decap_8 FILLER_45_381 ();
 sg13g2_decap_8 FILLER_45_388 ();
 sg13g2_decap_8 FILLER_45_395 ();
 sg13g2_decap_8 FILLER_45_402 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_7 ();
 sg13g2_decap_8 FILLER_46_14 ();
 sg13g2_decap_8 FILLER_46_21 ();
 sg13g2_decap_8 FILLER_46_28 ();
 sg13g2_decap_8 FILLER_46_35 ();
 sg13g2_decap_8 FILLER_46_42 ();
 sg13g2_decap_4 FILLER_46_49 ();
 sg13g2_fill_1 FILLER_46_53 ();
 sg13g2_fill_2 FILLER_46_89 ();
 sg13g2_fill_1 FILLER_46_91 ();
 sg13g2_fill_2 FILLER_46_101 ();
 sg13g2_fill_2 FILLER_46_112 ();
 sg13g2_fill_1 FILLER_46_114 ();
 sg13g2_fill_1 FILLER_46_162 ();
 sg13g2_fill_1 FILLER_46_195 ();
 sg13g2_decap_8 FILLER_46_237 ();
 sg13g2_decap_8 FILLER_46_244 ();
 sg13g2_decap_8 FILLER_46_251 ();
 sg13g2_fill_2 FILLER_46_258 ();
 sg13g2_fill_2 FILLER_46_283 ();
 sg13g2_fill_1 FILLER_46_285 ();
 sg13g2_fill_1 FILLER_46_311 ();
 sg13g2_decap_8 FILLER_46_324 ();
 sg13g2_decap_8 FILLER_46_331 ();
 sg13g2_decap_8 FILLER_46_338 ();
 sg13g2_decap_8 FILLER_46_345 ();
 sg13g2_decap_8 FILLER_46_352 ();
 sg13g2_decap_8 FILLER_46_359 ();
 sg13g2_decap_8 FILLER_46_366 ();
 sg13g2_decap_8 FILLER_46_373 ();
 sg13g2_decap_8 FILLER_46_380 ();
 sg13g2_decap_8 FILLER_46_387 ();
 sg13g2_decap_8 FILLER_46_394 ();
 sg13g2_decap_8 FILLER_46_401 ();
 sg13g2_fill_1 FILLER_46_408 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_7 ();
 sg13g2_decap_8 FILLER_47_14 ();
 sg13g2_decap_8 FILLER_47_21 ();
 sg13g2_decap_8 FILLER_47_28 ();
 sg13g2_decap_8 FILLER_47_35 ();
 sg13g2_decap_4 FILLER_47_42 ();
 sg13g2_fill_2 FILLER_47_46 ();
 sg13g2_decap_4 FILLER_47_126 ();
 sg13g2_fill_1 FILLER_47_260 ();
 sg13g2_decap_4 FILLER_47_270 ();
 sg13g2_decap_8 FILLER_47_286 ();
 sg13g2_fill_1 FILLER_47_293 ();
 sg13g2_fill_2 FILLER_47_302 ();
 sg13g2_fill_1 FILLER_47_304 ();
 sg13g2_fill_2 FILLER_47_311 ();
 sg13g2_decap_4 FILLER_47_323 ();
 sg13g2_fill_2 FILLER_47_327 ();
 sg13g2_fill_1 FILLER_47_340 ();
 sg13g2_decap_8 FILLER_47_351 ();
 sg13g2_decap_8 FILLER_47_358 ();
 sg13g2_decap_8 FILLER_47_365 ();
 sg13g2_decap_8 FILLER_47_372 ();
 sg13g2_decap_8 FILLER_47_379 ();
 sg13g2_decap_8 FILLER_47_386 ();
 sg13g2_decap_8 FILLER_47_393 ();
 sg13g2_decap_8 FILLER_47_400 ();
 sg13g2_fill_2 FILLER_47_407 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_decap_8 FILLER_48_14 ();
 sg13g2_decap_8 FILLER_48_21 ();
 sg13g2_decap_8 FILLER_48_28 ();
 sg13g2_decap_8 FILLER_48_35 ();
 sg13g2_decap_8 FILLER_48_42 ();
 sg13g2_decap_8 FILLER_48_49 ();
 sg13g2_decap_4 FILLER_48_56 ();
 sg13g2_decap_4 FILLER_48_74 ();
 sg13g2_decap_4 FILLER_48_82 ();
 sg13g2_fill_1 FILLER_48_110 ();
 sg13g2_fill_1 FILLER_48_124 ();
 sg13g2_fill_2 FILLER_48_151 ();
 sg13g2_fill_1 FILLER_48_153 ();
 sg13g2_decap_4 FILLER_48_158 ();
 sg13g2_decap_8 FILLER_48_167 ();
 sg13g2_decap_8 FILLER_48_174 ();
 sg13g2_decap_8 FILLER_48_186 ();
 sg13g2_decap_8 FILLER_48_193 ();
 sg13g2_fill_2 FILLER_48_200 ();
 sg13g2_fill_1 FILLER_48_202 ();
 sg13g2_fill_2 FILLER_48_208 ();
 sg13g2_fill_2 FILLER_48_218 ();
 sg13g2_fill_2 FILLER_48_248 ();
 sg13g2_fill_1 FILLER_48_250 ();
 sg13g2_decap_8 FILLER_48_255 ();
 sg13g2_fill_2 FILLER_48_262 ();
 sg13g2_fill_1 FILLER_48_264 ();
 sg13g2_decap_8 FILLER_48_275 ();
 sg13g2_decap_8 FILLER_48_282 ();
 sg13g2_decap_8 FILLER_48_289 ();
 sg13g2_decap_4 FILLER_48_296 ();
 sg13g2_fill_2 FILLER_48_300 ();
 sg13g2_fill_2 FILLER_48_316 ();
 sg13g2_fill_1 FILLER_48_318 ();
 sg13g2_decap_8 FILLER_48_359 ();
 sg13g2_decap_8 FILLER_48_366 ();
 sg13g2_decap_8 FILLER_48_373 ();
 sg13g2_decap_8 FILLER_48_380 ();
 sg13g2_decap_8 FILLER_48_387 ();
 sg13g2_decap_8 FILLER_48_394 ();
 sg13g2_decap_8 FILLER_48_401 ();
 sg13g2_fill_1 FILLER_48_408 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_7 ();
 sg13g2_decap_8 FILLER_49_14 ();
 sg13g2_decap_8 FILLER_49_21 ();
 sg13g2_decap_8 FILLER_49_28 ();
 sg13g2_decap_8 FILLER_49_35 ();
 sg13g2_decap_4 FILLER_49_42 ();
 sg13g2_fill_1 FILLER_49_46 ();
 sg13g2_fill_2 FILLER_49_81 ();
 sg13g2_fill_2 FILLER_49_87 ();
 sg13g2_fill_1 FILLER_49_89 ();
 sg13g2_fill_1 FILLER_49_102 ();
 sg13g2_fill_2 FILLER_49_120 ();
 sg13g2_fill_1 FILLER_49_122 ();
 sg13g2_fill_1 FILLER_49_128 ();
 sg13g2_decap_4 FILLER_49_150 ();
 sg13g2_fill_1 FILLER_49_183 ();
 sg13g2_decap_8 FILLER_49_196 ();
 sg13g2_decap_4 FILLER_49_203 ();
 sg13g2_fill_1 FILLER_49_207 ();
 sg13g2_decap_4 FILLER_49_212 ();
 sg13g2_decap_4 FILLER_49_220 ();
 sg13g2_decap_4 FILLER_49_229 ();
 sg13g2_fill_2 FILLER_49_233 ();
 sg13g2_fill_2 FILLER_49_282 ();
 sg13g2_fill_2 FILLER_49_296 ();
 sg13g2_fill_2 FILLER_49_325 ();
 sg13g2_fill_1 FILLER_49_327 ();
 sg13g2_decap_8 FILLER_49_352 ();
 sg13g2_decap_8 FILLER_49_359 ();
 sg13g2_decap_8 FILLER_49_366 ();
 sg13g2_decap_8 FILLER_49_373 ();
 sg13g2_decap_8 FILLER_49_380 ();
 sg13g2_decap_8 FILLER_49_387 ();
 sg13g2_decap_8 FILLER_49_394 ();
 sg13g2_decap_8 FILLER_49_401 ();
 sg13g2_fill_1 FILLER_49_408 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_8 FILLER_50_7 ();
 sg13g2_decap_8 FILLER_50_14 ();
 sg13g2_decap_8 FILLER_50_21 ();
 sg13g2_decap_8 FILLER_50_28 ();
 sg13g2_decap_8 FILLER_50_35 ();
 sg13g2_decap_8 FILLER_50_42 ();
 sg13g2_fill_2 FILLER_50_49 ();
 sg13g2_fill_1 FILLER_50_92 ();
 sg13g2_fill_1 FILLER_50_141 ();
 sg13g2_decap_4 FILLER_50_168 ();
 sg13g2_fill_2 FILLER_50_172 ();
 sg13g2_fill_1 FILLER_50_178 ();
 sg13g2_fill_2 FILLER_50_188 ();
 sg13g2_fill_2 FILLER_50_194 ();
 sg13g2_fill_1 FILLER_50_196 ();
 sg13g2_decap_8 FILLER_50_223 ();
 sg13g2_fill_1 FILLER_50_240 ();
 sg13g2_fill_1 FILLER_50_256 ();
 sg13g2_fill_2 FILLER_50_269 ();
 sg13g2_fill_1 FILLER_50_271 ();
 sg13g2_fill_2 FILLER_50_278 ();
 sg13g2_fill_2 FILLER_50_285 ();
 sg13g2_fill_2 FILLER_50_314 ();
 sg13g2_fill_1 FILLER_50_334 ();
 sg13g2_decap_8 FILLER_50_361 ();
 sg13g2_decap_8 FILLER_50_368 ();
 sg13g2_decap_8 FILLER_50_375 ();
 sg13g2_decap_8 FILLER_50_382 ();
 sg13g2_decap_8 FILLER_50_389 ();
 sg13g2_decap_8 FILLER_50_396 ();
 sg13g2_decap_4 FILLER_50_403 ();
 sg13g2_fill_2 FILLER_50_407 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_decap_8 FILLER_51_7 ();
 sg13g2_decap_8 FILLER_51_14 ();
 sg13g2_decap_8 FILLER_51_21 ();
 sg13g2_decap_8 FILLER_51_28 ();
 sg13g2_decap_8 FILLER_51_35 ();
 sg13g2_decap_8 FILLER_51_42 ();
 sg13g2_fill_2 FILLER_51_67 ();
 sg13g2_fill_2 FILLER_51_120 ();
 sg13g2_fill_1 FILLER_51_122 ();
 sg13g2_fill_1 FILLER_51_140 ();
 sg13g2_fill_1 FILLER_51_162 ();
 sg13g2_fill_1 FILLER_51_184 ();
 sg13g2_fill_2 FILLER_51_190 ();
 sg13g2_fill_1 FILLER_51_197 ();
 sg13g2_decap_8 FILLER_51_229 ();
 sg13g2_fill_1 FILLER_51_236 ();
 sg13g2_fill_2 FILLER_51_275 ();
 sg13g2_fill_1 FILLER_51_277 ();
 sg13g2_fill_2 FILLER_51_286 ();
 sg13g2_fill_2 FILLER_51_306 ();
 sg13g2_fill_1 FILLER_51_308 ();
 sg13g2_fill_2 FILLER_51_315 ();
 sg13g2_fill_1 FILLER_51_317 ();
 sg13g2_decap_4 FILLER_51_337 ();
 sg13g2_decap_8 FILLER_51_351 ();
 sg13g2_decap_8 FILLER_51_358 ();
 sg13g2_decap_8 FILLER_51_365 ();
 sg13g2_decap_8 FILLER_51_372 ();
 sg13g2_decap_8 FILLER_51_379 ();
 sg13g2_decap_8 FILLER_51_386 ();
 sg13g2_decap_8 FILLER_51_393 ();
 sg13g2_decap_8 FILLER_51_400 ();
 sg13g2_fill_2 FILLER_51_407 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_decap_8 FILLER_52_7 ();
 sg13g2_decap_8 FILLER_52_14 ();
 sg13g2_decap_8 FILLER_52_21 ();
 sg13g2_decap_8 FILLER_52_28 ();
 sg13g2_decap_8 FILLER_52_35 ();
 sg13g2_decap_8 FILLER_52_42 ();
 sg13g2_decap_4 FILLER_52_49 ();
 sg13g2_fill_2 FILLER_52_53 ();
 sg13g2_fill_1 FILLER_52_71 ();
 sg13g2_fill_2 FILLER_52_128 ();
 sg13g2_fill_1 FILLER_52_130 ();
 sg13g2_fill_2 FILLER_52_144 ();
 sg13g2_fill_2 FILLER_52_159 ();
 sg13g2_decap_4 FILLER_52_237 ();
 sg13g2_fill_1 FILLER_52_241 ();
 sg13g2_fill_2 FILLER_52_246 ();
 sg13g2_fill_1 FILLER_52_252 ();
 sg13g2_fill_2 FILLER_52_262 ();
 sg13g2_fill_1 FILLER_52_264 ();
 sg13g2_fill_2 FILLER_52_289 ();
 sg13g2_fill_2 FILLER_52_307 ();
 sg13g2_fill_2 FILLER_52_333 ();
 sg13g2_decap_8 FILLER_52_356 ();
 sg13g2_decap_8 FILLER_52_363 ();
 sg13g2_decap_8 FILLER_52_370 ();
 sg13g2_decap_8 FILLER_52_377 ();
 sg13g2_decap_8 FILLER_52_384 ();
 sg13g2_decap_8 FILLER_52_391 ();
 sg13g2_decap_8 FILLER_52_398 ();
 sg13g2_decap_4 FILLER_52_405 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_decap_8 FILLER_53_7 ();
 sg13g2_decap_8 FILLER_53_14 ();
 sg13g2_decap_8 FILLER_53_21 ();
 sg13g2_decap_8 FILLER_53_28 ();
 sg13g2_decap_8 FILLER_53_35 ();
 sg13g2_decap_8 FILLER_53_42 ();
 sg13g2_fill_2 FILLER_53_68 ();
 sg13g2_fill_2 FILLER_53_79 ();
 sg13g2_fill_1 FILLER_53_86 ();
 sg13g2_fill_1 FILLER_53_116 ();
 sg13g2_fill_2 FILLER_53_139 ();
 sg13g2_fill_1 FILLER_53_141 ();
 sg13g2_fill_2 FILLER_53_168 ();
 sg13g2_fill_1 FILLER_53_170 ();
 sg13g2_decap_8 FILLER_53_198 ();
 sg13g2_decap_4 FILLER_53_205 ();
 sg13g2_decap_8 FILLER_53_217 ();
 sg13g2_decap_8 FILLER_53_224 ();
 sg13g2_decap_4 FILLER_53_231 ();
 sg13g2_fill_1 FILLER_53_235 ();
 sg13g2_decap_8 FILLER_53_241 ();
 sg13g2_decap_4 FILLER_53_248 ();
 sg13g2_decap_4 FILLER_53_257 ();
 sg13g2_fill_2 FILLER_53_276 ();
 sg13g2_decap_8 FILLER_53_283 ();
 sg13g2_fill_1 FILLER_53_290 ();
 sg13g2_decap_4 FILLER_53_299 ();
 sg13g2_fill_1 FILLER_53_303 ();
 sg13g2_decap_8 FILLER_53_314 ();
 sg13g2_fill_2 FILLER_53_321 ();
 sg13g2_decap_8 FILLER_53_345 ();
 sg13g2_decap_8 FILLER_53_352 ();
 sg13g2_decap_8 FILLER_53_359 ();
 sg13g2_decap_8 FILLER_53_366 ();
 sg13g2_decap_8 FILLER_53_373 ();
 sg13g2_decap_8 FILLER_53_380 ();
 sg13g2_decap_8 FILLER_53_387 ();
 sg13g2_decap_8 FILLER_53_394 ();
 sg13g2_decap_8 FILLER_53_401 ();
 sg13g2_fill_1 FILLER_53_408 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_decap_8 FILLER_54_7 ();
 sg13g2_decap_8 FILLER_54_14 ();
 sg13g2_decap_8 FILLER_54_21 ();
 sg13g2_decap_8 FILLER_54_28 ();
 sg13g2_decap_8 FILLER_54_35 ();
 sg13g2_decap_4 FILLER_54_42 ();
 sg13g2_fill_2 FILLER_54_80 ();
 sg13g2_fill_2 FILLER_54_169 ();
 sg13g2_fill_1 FILLER_54_180 ();
 sg13g2_fill_2 FILLER_54_186 ();
 sg13g2_decap_4 FILLER_54_193 ();
 sg13g2_fill_1 FILLER_54_197 ();
 sg13g2_decap_8 FILLER_54_224 ();
 sg13g2_decap_4 FILLER_54_231 ();
 sg13g2_decap_8 FILLER_54_241 ();
 sg13g2_decap_4 FILLER_54_248 ();
 sg13g2_fill_2 FILLER_54_252 ();
 sg13g2_fill_1 FILLER_54_259 ();
 sg13g2_fill_2 FILLER_54_270 ();
 sg13g2_fill_1 FILLER_54_272 ();
 sg13g2_decap_4 FILLER_54_283 ();
 sg13g2_decap_8 FILLER_54_292 ();
 sg13g2_decap_4 FILLER_54_304 ();
 sg13g2_decap_8 FILLER_54_320 ();
 sg13g2_decap_8 FILLER_54_327 ();
 sg13g2_decap_8 FILLER_54_343 ();
 sg13g2_decap_8 FILLER_54_350 ();
 sg13g2_decap_8 FILLER_54_357 ();
 sg13g2_decap_8 FILLER_54_364 ();
 sg13g2_decap_8 FILLER_54_371 ();
 sg13g2_decap_8 FILLER_54_378 ();
 sg13g2_decap_8 FILLER_54_385 ();
 sg13g2_decap_8 FILLER_54_392 ();
 sg13g2_decap_8 FILLER_54_399 ();
 sg13g2_fill_2 FILLER_54_406 ();
 sg13g2_fill_1 FILLER_54_408 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_decap_8 FILLER_55_7 ();
 sg13g2_decap_8 FILLER_55_14 ();
 sg13g2_decap_8 FILLER_55_21 ();
 sg13g2_decap_8 FILLER_55_28 ();
 sg13g2_decap_8 FILLER_55_35 ();
 sg13g2_decap_8 FILLER_55_42 ();
 sg13g2_fill_2 FILLER_55_49 ();
 sg13g2_fill_1 FILLER_55_51 ();
 sg13g2_fill_2 FILLER_55_61 ();
 sg13g2_fill_1 FILLER_55_98 ();
 sg13g2_fill_2 FILLER_55_129 ();
 sg13g2_fill_2 FILLER_55_139 ();
 sg13g2_fill_1 FILLER_55_155 ();
 sg13g2_decap_8 FILLER_55_182 ();
 sg13g2_decap_8 FILLER_55_189 ();
 sg13g2_fill_2 FILLER_55_196 ();
 sg13g2_decap_4 FILLER_55_224 ();
 sg13g2_fill_2 FILLER_55_228 ();
 sg13g2_fill_2 FILLER_55_244 ();
 sg13g2_fill_1 FILLER_55_246 ();
 sg13g2_decap_4 FILLER_55_260 ();
 sg13g2_fill_1 FILLER_55_277 ();
 sg13g2_decap_4 FILLER_55_297 ();
 sg13g2_decap_8 FILLER_55_345 ();
 sg13g2_decap_8 FILLER_55_352 ();
 sg13g2_decap_8 FILLER_55_359 ();
 sg13g2_decap_8 FILLER_55_366 ();
 sg13g2_decap_8 FILLER_55_373 ();
 sg13g2_decap_8 FILLER_55_380 ();
 sg13g2_decap_8 FILLER_55_387 ();
 sg13g2_decap_8 FILLER_55_394 ();
 sg13g2_decap_8 FILLER_55_401 ();
 sg13g2_fill_1 FILLER_55_408 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_decap_8 FILLER_56_7 ();
 sg13g2_decap_8 FILLER_56_14 ();
 sg13g2_decap_8 FILLER_56_21 ();
 sg13g2_decap_8 FILLER_56_28 ();
 sg13g2_decap_8 FILLER_56_35 ();
 sg13g2_decap_8 FILLER_56_42 ();
 sg13g2_fill_2 FILLER_56_49 ();
 sg13g2_fill_1 FILLER_56_51 ();
 sg13g2_fill_2 FILLER_56_98 ();
 sg13g2_fill_2 FILLER_56_126 ();
 sg13g2_fill_2 FILLER_56_155 ();
 sg13g2_fill_2 FILLER_56_191 ();
 sg13g2_fill_1 FILLER_56_193 ();
 sg13g2_decap_4 FILLER_56_203 ();
 sg13g2_fill_2 FILLER_56_207 ();
 sg13g2_decap_8 FILLER_56_217 ();
 sg13g2_fill_2 FILLER_56_261 ();
 sg13g2_fill_1 FILLER_56_291 ();
 sg13g2_fill_2 FILLER_56_300 ();
 sg13g2_fill_1 FILLER_56_302 ();
 sg13g2_fill_2 FILLER_56_327 ();
 sg13g2_fill_1 FILLER_56_329 ();
 sg13g2_decap_8 FILLER_56_354 ();
 sg13g2_decap_8 FILLER_56_361 ();
 sg13g2_decap_8 FILLER_56_368 ();
 sg13g2_decap_8 FILLER_56_375 ();
 sg13g2_decap_8 FILLER_56_382 ();
 sg13g2_decap_8 FILLER_56_389 ();
 sg13g2_decap_8 FILLER_56_396 ();
 sg13g2_decap_4 FILLER_56_403 ();
 sg13g2_fill_2 FILLER_56_407 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_decap_8 FILLER_57_7 ();
 sg13g2_decap_8 FILLER_57_14 ();
 sg13g2_decap_8 FILLER_57_21 ();
 sg13g2_decap_8 FILLER_57_28 ();
 sg13g2_decap_8 FILLER_57_35 ();
 sg13g2_decap_8 FILLER_57_42 ();
 sg13g2_decap_8 FILLER_57_49 ();
 sg13g2_fill_1 FILLER_57_60 ();
 sg13g2_fill_2 FILLER_57_66 ();
 sg13g2_fill_2 FILLER_57_99 ();
 sg13g2_fill_2 FILLER_57_161 ();
 sg13g2_fill_2 FILLER_57_171 ();
 sg13g2_fill_1 FILLER_57_173 ();
 sg13g2_decap_8 FILLER_57_212 ();
 sg13g2_decap_8 FILLER_57_219 ();
 sg13g2_decap_4 FILLER_57_226 ();
 sg13g2_fill_2 FILLER_57_230 ();
 sg13g2_fill_2 FILLER_57_257 ();
 sg13g2_decap_4 FILLER_57_266 ();
 sg13g2_fill_2 FILLER_57_292 ();
 sg13g2_fill_1 FILLER_57_322 ();
 sg13g2_fill_2 FILLER_57_329 ();
 sg13g2_decap_8 FILLER_57_353 ();
 sg13g2_decap_8 FILLER_57_360 ();
 sg13g2_decap_8 FILLER_57_367 ();
 sg13g2_decap_8 FILLER_57_374 ();
 sg13g2_decap_8 FILLER_57_381 ();
 sg13g2_decap_8 FILLER_57_388 ();
 sg13g2_decap_8 FILLER_57_395 ();
 sg13g2_decap_8 FILLER_57_402 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_decap_8 FILLER_58_7 ();
 sg13g2_decap_8 FILLER_58_14 ();
 sg13g2_decap_8 FILLER_58_21 ();
 sg13g2_decap_8 FILLER_58_28 ();
 sg13g2_decap_8 FILLER_58_35 ();
 sg13g2_decap_8 FILLER_58_42 ();
 sg13g2_decap_4 FILLER_58_49 ();
 sg13g2_fill_1 FILLER_58_53 ();
 sg13g2_fill_2 FILLER_58_90 ();
 sg13g2_fill_1 FILLER_58_92 ();
 sg13g2_fill_1 FILLER_58_124 ();
 sg13g2_fill_2 FILLER_58_142 ();
 sg13g2_fill_1 FILLER_58_144 ();
 sg13g2_decap_8 FILLER_58_221 ();
 sg13g2_fill_2 FILLER_58_228 ();
 sg13g2_fill_1 FILLER_58_236 ();
 sg13g2_fill_2 FILLER_58_255 ();
 sg13g2_fill_1 FILLER_58_257 ();
 sg13g2_fill_2 FILLER_58_295 ();
 sg13g2_fill_1 FILLER_58_297 ();
 sg13g2_decap_8 FILLER_58_306 ();
 sg13g2_decap_8 FILLER_58_342 ();
 sg13g2_decap_8 FILLER_58_349 ();
 sg13g2_decap_8 FILLER_58_356 ();
 sg13g2_decap_8 FILLER_58_363 ();
 sg13g2_decap_8 FILLER_58_370 ();
 sg13g2_decap_8 FILLER_58_377 ();
 sg13g2_decap_8 FILLER_58_384 ();
 sg13g2_decap_8 FILLER_58_391 ();
 sg13g2_decap_8 FILLER_58_398 ();
 sg13g2_decap_4 FILLER_58_405 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_decap_8 FILLER_59_7 ();
 sg13g2_decap_8 FILLER_59_14 ();
 sg13g2_decap_8 FILLER_59_21 ();
 sg13g2_decap_8 FILLER_59_28 ();
 sg13g2_decap_8 FILLER_59_35 ();
 sg13g2_decap_4 FILLER_59_42 ();
 sg13g2_fill_2 FILLER_59_46 ();
 sg13g2_fill_1 FILLER_59_98 ();
 sg13g2_fill_2 FILLER_59_121 ();
 sg13g2_decap_8 FILLER_59_211 ();
 sg13g2_decap_8 FILLER_59_218 ();
 sg13g2_fill_2 FILLER_59_225 ();
 sg13g2_fill_2 FILLER_59_231 ();
 sg13g2_decap_8 FILLER_59_240 ();
 sg13g2_fill_2 FILLER_59_247 ();
 sg13g2_decap_4 FILLER_59_254 ();
 sg13g2_fill_1 FILLER_59_273 ();
 sg13g2_fill_1 FILLER_59_285 ();
 sg13g2_decap_4 FILLER_59_292 ();
 sg13g2_fill_1 FILLER_59_296 ();
 sg13g2_decap_8 FILLER_59_302 ();
 sg13g2_decap_8 FILLER_59_309 ();
 sg13g2_decap_4 FILLER_59_316 ();
 sg13g2_fill_1 FILLER_59_320 ();
 sg13g2_decap_8 FILLER_59_337 ();
 sg13g2_decap_8 FILLER_59_344 ();
 sg13g2_decap_8 FILLER_59_351 ();
 sg13g2_decap_8 FILLER_59_358 ();
 sg13g2_decap_8 FILLER_59_365 ();
 sg13g2_decap_8 FILLER_59_372 ();
 sg13g2_decap_8 FILLER_59_379 ();
 sg13g2_decap_8 FILLER_59_386 ();
 sg13g2_decap_8 FILLER_59_393 ();
 sg13g2_decap_8 FILLER_59_400 ();
 sg13g2_fill_2 FILLER_59_407 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_decap_8 FILLER_60_7 ();
 sg13g2_decap_8 FILLER_60_14 ();
 sg13g2_decap_8 FILLER_60_21 ();
 sg13g2_decap_8 FILLER_60_28 ();
 sg13g2_decap_8 FILLER_60_35 ();
 sg13g2_decap_8 FILLER_60_42 ();
 sg13g2_fill_2 FILLER_60_107 ();
 sg13g2_fill_2 FILLER_60_121 ();
 sg13g2_fill_1 FILLER_60_123 ();
 sg13g2_fill_1 FILLER_60_177 ();
 sg13g2_decap_4 FILLER_60_242 ();
 sg13g2_fill_2 FILLER_60_246 ();
 sg13g2_decap_4 FILLER_60_283 ();
 sg13g2_fill_2 FILLER_60_298 ();
 sg13g2_fill_1 FILLER_60_300 ();
 sg13g2_fill_2 FILLER_60_317 ();
 sg13g2_fill_1 FILLER_60_319 ();
 sg13g2_decap_8 FILLER_60_339 ();
 sg13g2_decap_8 FILLER_60_346 ();
 sg13g2_decap_8 FILLER_60_353 ();
 sg13g2_decap_8 FILLER_60_360 ();
 sg13g2_decap_8 FILLER_60_367 ();
 sg13g2_decap_8 FILLER_60_374 ();
 sg13g2_decap_8 FILLER_60_381 ();
 sg13g2_decap_8 FILLER_60_388 ();
 sg13g2_decap_8 FILLER_60_395 ();
 sg13g2_decap_8 FILLER_60_402 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_decap_8 FILLER_61_7 ();
 sg13g2_decap_8 FILLER_61_14 ();
 sg13g2_decap_8 FILLER_61_21 ();
 sg13g2_decap_8 FILLER_61_28 ();
 sg13g2_decap_8 FILLER_61_35 ();
 sg13g2_fill_1 FILLER_61_42 ();
 sg13g2_fill_2 FILLER_61_61 ();
 sg13g2_fill_1 FILLER_61_63 ();
 sg13g2_fill_1 FILLER_61_86 ();
 sg13g2_fill_2 FILLER_61_165 ();
 sg13g2_fill_1 FILLER_61_167 ();
 sg13g2_fill_2 FILLER_61_207 ();
 sg13g2_fill_1 FILLER_61_222 ();
 sg13g2_fill_2 FILLER_61_253 ();
 sg13g2_fill_1 FILLER_61_255 ();
 sg13g2_decap_8 FILLER_61_279 ();
 sg13g2_decap_4 FILLER_61_286 ();
 sg13g2_fill_1 FILLER_61_290 ();
 sg13g2_fill_2 FILLER_61_329 ();
 sg13g2_fill_1 FILLER_61_331 ();
 sg13g2_decap_8 FILLER_61_345 ();
 sg13g2_decap_8 FILLER_61_352 ();
 sg13g2_decap_8 FILLER_61_359 ();
 sg13g2_decap_8 FILLER_61_366 ();
 sg13g2_decap_8 FILLER_61_373 ();
 sg13g2_decap_8 FILLER_61_380 ();
 sg13g2_decap_8 FILLER_61_387 ();
 sg13g2_decap_8 FILLER_61_394 ();
 sg13g2_decap_8 FILLER_61_401 ();
 sg13g2_fill_1 FILLER_61_408 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_decap_8 FILLER_62_7 ();
 sg13g2_decap_8 FILLER_62_14 ();
 sg13g2_decap_8 FILLER_62_21 ();
 sg13g2_decap_8 FILLER_62_28 ();
 sg13g2_decap_8 FILLER_62_35 ();
 sg13g2_decap_8 FILLER_62_42 ();
 sg13g2_fill_1 FILLER_62_49 ();
 sg13g2_fill_2 FILLER_62_65 ();
 sg13g2_fill_2 FILLER_62_84 ();
 sg13g2_fill_2 FILLER_62_108 ();
 sg13g2_fill_1 FILLER_62_110 ();
 sg13g2_fill_1 FILLER_62_120 ();
 sg13g2_fill_1 FILLER_62_204 ();
 sg13g2_fill_2 FILLER_62_244 ();
 sg13g2_decap_4 FILLER_62_265 ();
 sg13g2_fill_1 FILLER_62_269 ();
 sg13g2_fill_2 FILLER_62_285 ();
 sg13g2_fill_1 FILLER_62_287 ();
 sg13g2_fill_1 FILLER_62_334 ();
 sg13g2_decap_8 FILLER_62_343 ();
 sg13g2_decap_8 FILLER_62_350 ();
 sg13g2_decap_8 FILLER_62_357 ();
 sg13g2_decap_8 FILLER_62_364 ();
 sg13g2_decap_8 FILLER_62_371 ();
 sg13g2_decap_8 FILLER_62_378 ();
 sg13g2_decap_8 FILLER_62_385 ();
 sg13g2_decap_8 FILLER_62_392 ();
 sg13g2_decap_8 FILLER_62_399 ();
 sg13g2_fill_2 FILLER_62_406 ();
 sg13g2_fill_1 FILLER_62_408 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_decap_8 FILLER_63_7 ();
 sg13g2_decap_8 FILLER_63_14 ();
 sg13g2_decap_8 FILLER_63_21 ();
 sg13g2_decap_8 FILLER_63_28 ();
 sg13g2_decap_8 FILLER_63_35 ();
 sg13g2_decap_8 FILLER_63_42 ();
 sg13g2_decap_8 FILLER_63_49 ();
 sg13g2_fill_2 FILLER_63_56 ();
 sg13g2_fill_1 FILLER_63_58 ();
 sg13g2_fill_2 FILLER_63_133 ();
 sg13g2_fill_1 FILLER_63_156 ();
 sg13g2_fill_2 FILLER_63_181 ();
 sg13g2_fill_1 FILLER_63_183 ();
 sg13g2_fill_1 FILLER_63_211 ();
 sg13g2_fill_2 FILLER_63_256 ();
 sg13g2_fill_2 FILLER_63_279 ();
 sg13g2_fill_1 FILLER_63_281 ();
 sg13g2_fill_1 FILLER_63_318 ();
 sg13g2_decap_8 FILLER_63_341 ();
 sg13g2_decap_8 FILLER_63_348 ();
 sg13g2_decap_8 FILLER_63_355 ();
 sg13g2_decap_8 FILLER_63_362 ();
 sg13g2_decap_8 FILLER_63_369 ();
 sg13g2_decap_8 FILLER_63_376 ();
 sg13g2_decap_8 FILLER_63_383 ();
 sg13g2_decap_8 FILLER_63_390 ();
 sg13g2_decap_8 FILLER_63_397 ();
 sg13g2_decap_4 FILLER_63_404 ();
 sg13g2_fill_1 FILLER_63_408 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_8 FILLER_64_7 ();
 sg13g2_decap_8 FILLER_64_14 ();
 sg13g2_decap_8 FILLER_64_21 ();
 sg13g2_decap_8 FILLER_64_28 ();
 sg13g2_decap_8 FILLER_64_35 ();
 sg13g2_decap_8 FILLER_64_42 ();
 sg13g2_decap_8 FILLER_64_49 ();
 sg13g2_decap_8 FILLER_64_56 ();
 sg13g2_decap_4 FILLER_64_63 ();
 sg13g2_fill_1 FILLER_64_67 ();
 sg13g2_fill_2 FILLER_64_94 ();
 sg13g2_fill_1 FILLER_64_96 ();
 sg13g2_fill_1 FILLER_64_155 ();
 sg13g2_fill_2 FILLER_64_198 ();
 sg13g2_fill_1 FILLER_64_200 ();
 sg13g2_decap_8 FILLER_64_210 ();
 sg13g2_fill_2 FILLER_64_227 ();
 sg13g2_fill_1 FILLER_64_229 ();
 sg13g2_decap_4 FILLER_64_283 ();
 sg13g2_decap_8 FILLER_64_300 ();
 sg13g2_decap_8 FILLER_64_307 ();
 sg13g2_decap_4 FILLER_64_314 ();
 sg13g2_fill_1 FILLER_64_318 ();
 sg13g2_decap_8 FILLER_64_334 ();
 sg13g2_decap_8 FILLER_64_341 ();
 sg13g2_decap_8 FILLER_64_348 ();
 sg13g2_decap_8 FILLER_64_355 ();
 sg13g2_decap_8 FILLER_64_362 ();
 sg13g2_decap_8 FILLER_64_369 ();
 sg13g2_decap_8 FILLER_64_376 ();
 sg13g2_decap_8 FILLER_64_383 ();
 sg13g2_decap_8 FILLER_64_390 ();
 sg13g2_decap_8 FILLER_64_397 ();
 sg13g2_decap_4 FILLER_64_404 ();
 sg13g2_fill_1 FILLER_64_408 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_8 FILLER_65_7 ();
 sg13g2_decap_8 FILLER_65_14 ();
 sg13g2_decap_8 FILLER_65_21 ();
 sg13g2_decap_8 FILLER_65_28 ();
 sg13g2_decap_8 FILLER_65_35 ();
 sg13g2_decap_8 FILLER_65_42 ();
 sg13g2_decap_8 FILLER_65_49 ();
 sg13g2_decap_8 FILLER_65_56 ();
 sg13g2_decap_8 FILLER_65_63 ();
 sg13g2_decap_8 FILLER_65_70 ();
 sg13g2_fill_2 FILLER_65_77 ();
 sg13g2_decap_4 FILLER_65_83 ();
 sg13g2_fill_1 FILLER_65_103 ();
 sg13g2_fill_2 FILLER_65_122 ();
 sg13g2_fill_1 FILLER_65_150 ();
 sg13g2_decap_8 FILLER_65_196 ();
 sg13g2_fill_2 FILLER_65_203 ();
 sg13g2_fill_2 FILLER_65_247 ();
 sg13g2_fill_1 FILLER_65_249 ();
 sg13g2_decap_4 FILLER_65_255 ();
 sg13g2_decap_4 FILLER_65_276 ();
 sg13g2_decap_8 FILLER_65_285 ();
 sg13g2_decap_8 FILLER_65_292 ();
 sg13g2_decap_4 FILLER_65_316 ();
 sg13g2_fill_1 FILLER_65_320 ();
 sg13g2_decap_8 FILLER_65_342 ();
 sg13g2_decap_8 FILLER_65_349 ();
 sg13g2_decap_8 FILLER_65_356 ();
 sg13g2_decap_8 FILLER_65_363 ();
 sg13g2_decap_8 FILLER_65_370 ();
 sg13g2_decap_8 FILLER_65_377 ();
 sg13g2_decap_8 FILLER_65_384 ();
 sg13g2_decap_8 FILLER_65_391 ();
 sg13g2_decap_8 FILLER_65_398 ();
 sg13g2_decap_4 FILLER_65_405 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_8 FILLER_66_7 ();
 sg13g2_decap_8 FILLER_66_14 ();
 sg13g2_decap_8 FILLER_66_21 ();
 sg13g2_decap_8 FILLER_66_28 ();
 sg13g2_decap_8 FILLER_66_35 ();
 sg13g2_decap_8 FILLER_66_42 ();
 sg13g2_decap_8 FILLER_66_49 ();
 sg13g2_decap_8 FILLER_66_56 ();
 sg13g2_decap_8 FILLER_66_63 ();
 sg13g2_decap_8 FILLER_66_70 ();
 sg13g2_decap_8 FILLER_66_77 ();
 sg13g2_decap_8 FILLER_66_84 ();
 sg13g2_decap_8 FILLER_66_91 ();
 sg13g2_fill_2 FILLER_66_172 ();
 sg13g2_decap_8 FILLER_66_200 ();
 sg13g2_fill_1 FILLER_66_207 ();
 sg13g2_decap_8 FILLER_66_249 ();
 sg13g2_decap_4 FILLER_66_256 ();
 sg13g2_fill_1 FILLER_66_264 ();
 sg13g2_fill_1 FILLER_66_270 ();
 sg13g2_decap_4 FILLER_66_287 ();
 sg13g2_fill_2 FILLER_66_303 ();
 sg13g2_fill_1 FILLER_66_305 ();
 sg13g2_fill_1 FILLER_66_318 ();
 sg13g2_decap_8 FILLER_66_341 ();
 sg13g2_decap_8 FILLER_66_348 ();
 sg13g2_decap_8 FILLER_66_355 ();
 sg13g2_decap_8 FILLER_66_362 ();
 sg13g2_decap_8 FILLER_66_369 ();
 sg13g2_decap_8 FILLER_66_376 ();
 sg13g2_decap_8 FILLER_66_383 ();
 sg13g2_decap_8 FILLER_66_390 ();
 sg13g2_decap_8 FILLER_66_397 ();
 sg13g2_decap_4 FILLER_66_404 ();
 sg13g2_fill_1 FILLER_66_408 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_8 FILLER_67_7 ();
 sg13g2_decap_8 FILLER_67_14 ();
 sg13g2_decap_8 FILLER_67_21 ();
 sg13g2_decap_8 FILLER_67_28 ();
 sg13g2_decap_8 FILLER_67_35 ();
 sg13g2_decap_8 FILLER_67_42 ();
 sg13g2_decap_8 FILLER_67_49 ();
 sg13g2_decap_8 FILLER_67_56 ();
 sg13g2_decap_8 FILLER_67_63 ();
 sg13g2_decap_8 FILLER_67_70 ();
 sg13g2_decap_8 FILLER_67_77 ();
 sg13g2_decap_8 FILLER_67_84 ();
 sg13g2_decap_8 FILLER_67_91 ();
 sg13g2_decap_8 FILLER_67_98 ();
 sg13g2_fill_1 FILLER_67_108 ();
 sg13g2_decap_8 FILLER_67_113 ();
 sg13g2_fill_1 FILLER_67_120 ();
 sg13g2_fill_2 FILLER_67_171 ();
 sg13g2_decap_4 FILLER_67_208 ();
 sg13g2_fill_2 FILLER_67_212 ();
 sg13g2_decap_8 FILLER_67_241 ();
 sg13g2_fill_1 FILLER_67_253 ();
 sg13g2_fill_1 FILLER_67_259 ();
 sg13g2_fill_1 FILLER_67_271 ();
 sg13g2_fill_1 FILLER_67_294 ();
 sg13g2_decap_8 FILLER_67_341 ();
 sg13g2_decap_8 FILLER_67_348 ();
 sg13g2_decap_8 FILLER_67_355 ();
 sg13g2_decap_8 FILLER_67_362 ();
 sg13g2_decap_8 FILLER_67_369 ();
 sg13g2_decap_8 FILLER_67_376 ();
 sg13g2_decap_8 FILLER_67_383 ();
 sg13g2_decap_8 FILLER_67_390 ();
 sg13g2_decap_8 FILLER_67_397 ();
 sg13g2_decap_4 FILLER_67_404 ();
 sg13g2_fill_1 FILLER_67_408 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_8 FILLER_68_7 ();
 sg13g2_decap_8 FILLER_68_14 ();
 sg13g2_decap_8 FILLER_68_21 ();
 sg13g2_decap_8 FILLER_68_28 ();
 sg13g2_decap_8 FILLER_68_35 ();
 sg13g2_decap_8 FILLER_68_42 ();
 sg13g2_decap_8 FILLER_68_49 ();
 sg13g2_decap_8 FILLER_68_56 ();
 sg13g2_decap_8 FILLER_68_63 ();
 sg13g2_decap_8 FILLER_68_70 ();
 sg13g2_decap_8 FILLER_68_77 ();
 sg13g2_decap_8 FILLER_68_84 ();
 sg13g2_decap_8 FILLER_68_91 ();
 sg13g2_decap_8 FILLER_68_98 ();
 sg13g2_decap_8 FILLER_68_105 ();
 sg13g2_decap_4 FILLER_68_112 ();
 sg13g2_fill_1 FILLER_68_116 ();
 sg13g2_fill_1 FILLER_68_122 ();
 sg13g2_fill_2 FILLER_68_127 ();
 sg13g2_fill_1 FILLER_68_151 ();
 sg13g2_fill_2 FILLER_68_169 ();
 sg13g2_decap_8 FILLER_68_206 ();
 sg13g2_fill_2 FILLER_68_213 ();
 sg13g2_fill_1 FILLER_68_215 ();
 sg13g2_decap_4 FILLER_68_220 ();
 sg13g2_fill_1 FILLER_68_224 ();
 sg13g2_decap_8 FILLER_68_230 ();
 sg13g2_decap_4 FILLER_68_237 ();
 sg13g2_fill_2 FILLER_68_241 ();
 sg13g2_fill_1 FILLER_68_264 ();
 sg13g2_fill_2 FILLER_68_276 ();
 sg13g2_fill_1 FILLER_68_278 ();
 sg13g2_fill_1 FILLER_68_285 ();
 sg13g2_fill_2 FILLER_68_318 ();
 sg13g2_decap_8 FILLER_68_342 ();
 sg13g2_decap_8 FILLER_68_349 ();
 sg13g2_decap_8 FILLER_68_356 ();
 sg13g2_decap_8 FILLER_68_363 ();
 sg13g2_decap_8 FILLER_68_370 ();
 sg13g2_decap_8 FILLER_68_377 ();
 sg13g2_decap_8 FILLER_68_384 ();
 sg13g2_decap_8 FILLER_68_391 ();
 sg13g2_decap_8 FILLER_68_398 ();
 sg13g2_decap_4 FILLER_68_405 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_8 FILLER_69_7 ();
 sg13g2_decap_8 FILLER_69_14 ();
 sg13g2_decap_8 FILLER_69_21 ();
 sg13g2_decap_8 FILLER_69_28 ();
 sg13g2_decap_8 FILLER_69_35 ();
 sg13g2_decap_8 FILLER_69_42 ();
 sg13g2_decap_8 FILLER_69_49 ();
 sg13g2_decap_8 FILLER_69_56 ();
 sg13g2_decap_8 FILLER_69_63 ();
 sg13g2_decap_8 FILLER_69_70 ();
 sg13g2_decap_8 FILLER_69_77 ();
 sg13g2_decap_8 FILLER_69_84 ();
 sg13g2_decap_8 FILLER_69_91 ();
 sg13g2_decap_8 FILLER_69_98 ();
 sg13g2_decap_4 FILLER_69_105 ();
 sg13g2_fill_1 FILLER_69_109 ();
 sg13g2_fill_1 FILLER_69_140 ();
 sg13g2_decap_8 FILLER_69_157 ();
 sg13g2_fill_2 FILLER_69_164 ();
 sg13g2_fill_1 FILLER_69_166 ();
 sg13g2_decap_4 FILLER_69_197 ();
 sg13g2_fill_1 FILLER_69_209 ();
 sg13g2_decap_8 FILLER_69_237 ();
 sg13g2_fill_2 FILLER_69_244 ();
 sg13g2_fill_2 FILLER_69_265 ();
 sg13g2_fill_2 FILLER_69_278 ();
 sg13g2_decap_4 FILLER_69_306 ();
 sg13g2_fill_1 FILLER_69_310 ();
 sg13g2_decap_8 FILLER_69_334 ();
 sg13g2_decap_8 FILLER_69_341 ();
 sg13g2_decap_8 FILLER_69_348 ();
 sg13g2_decap_8 FILLER_69_355 ();
 sg13g2_decap_8 FILLER_69_362 ();
 sg13g2_decap_8 FILLER_69_369 ();
 sg13g2_decap_8 FILLER_69_376 ();
 sg13g2_decap_8 FILLER_69_383 ();
 sg13g2_decap_8 FILLER_69_390 ();
 sg13g2_decap_8 FILLER_69_397 ();
 sg13g2_decap_4 FILLER_69_404 ();
 sg13g2_fill_1 FILLER_69_408 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_decap_8 FILLER_70_14 ();
 sg13g2_decap_8 FILLER_70_21 ();
 sg13g2_decap_8 FILLER_70_28 ();
 sg13g2_decap_8 FILLER_70_35 ();
 sg13g2_decap_8 FILLER_70_42 ();
 sg13g2_decap_8 FILLER_70_49 ();
 sg13g2_decap_8 FILLER_70_56 ();
 sg13g2_decap_8 FILLER_70_63 ();
 sg13g2_decap_8 FILLER_70_70 ();
 sg13g2_decap_8 FILLER_70_77 ();
 sg13g2_decap_8 FILLER_70_84 ();
 sg13g2_decap_8 FILLER_70_91 ();
 sg13g2_fill_2 FILLER_70_98 ();
 sg13g2_fill_1 FILLER_70_100 ();
 sg13g2_fill_2 FILLER_70_124 ();
 sg13g2_fill_1 FILLER_70_178 ();
 sg13g2_fill_2 FILLER_70_205 ();
 sg13g2_fill_2 FILLER_70_246 ();
 sg13g2_fill_2 FILLER_70_255 ();
 sg13g2_decap_8 FILLER_70_282 ();
 sg13g2_fill_2 FILLER_70_289 ();
 sg13g2_fill_2 FILLER_70_296 ();
 sg13g2_fill_1 FILLER_70_298 ();
 sg13g2_fill_2 FILLER_70_305 ();
 sg13g2_fill_2 FILLER_70_313 ();
 sg13g2_fill_1 FILLER_70_315 ();
 sg13g2_decap_8 FILLER_70_330 ();
 sg13g2_decap_8 FILLER_70_337 ();
 sg13g2_decap_8 FILLER_70_344 ();
 sg13g2_decap_8 FILLER_70_351 ();
 sg13g2_decap_8 FILLER_70_358 ();
 sg13g2_decap_8 FILLER_70_365 ();
 sg13g2_decap_8 FILLER_70_372 ();
 sg13g2_decap_8 FILLER_70_379 ();
 sg13g2_decap_8 FILLER_70_386 ();
 sg13g2_decap_8 FILLER_70_393 ();
 sg13g2_decap_8 FILLER_70_400 ();
 sg13g2_fill_2 FILLER_70_407 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_decap_8 FILLER_71_7 ();
 sg13g2_decap_8 FILLER_71_14 ();
 sg13g2_decap_8 FILLER_71_21 ();
 sg13g2_decap_8 FILLER_71_28 ();
 sg13g2_decap_8 FILLER_71_35 ();
 sg13g2_decap_8 FILLER_71_42 ();
 sg13g2_decap_8 FILLER_71_49 ();
 sg13g2_decap_8 FILLER_71_56 ();
 sg13g2_decap_8 FILLER_71_63 ();
 sg13g2_decap_8 FILLER_71_70 ();
 sg13g2_decap_8 FILLER_71_77 ();
 sg13g2_decap_8 FILLER_71_84 ();
 sg13g2_decap_8 FILLER_71_91 ();
 sg13g2_fill_2 FILLER_71_98 ();
 sg13g2_fill_1 FILLER_71_126 ();
 sg13g2_fill_1 FILLER_71_141 ();
 sg13g2_fill_1 FILLER_71_203 ();
 sg13g2_fill_2 FILLER_71_238 ();
 sg13g2_fill_1 FILLER_71_240 ();
 sg13g2_decap_4 FILLER_71_266 ();
 sg13g2_fill_1 FILLER_71_270 ();
 sg13g2_fill_1 FILLER_71_276 ();
 sg13g2_fill_1 FILLER_71_291 ();
 sg13g2_fill_2 FILLER_71_304 ();
 sg13g2_fill_2 FILLER_71_325 ();
 sg13g2_decap_8 FILLER_71_335 ();
 sg13g2_decap_8 FILLER_71_342 ();
 sg13g2_decap_8 FILLER_71_349 ();
 sg13g2_decap_8 FILLER_71_356 ();
 sg13g2_decap_8 FILLER_71_363 ();
 sg13g2_decap_8 FILLER_71_370 ();
 sg13g2_decap_8 FILLER_71_377 ();
 sg13g2_decap_8 FILLER_71_384 ();
 sg13g2_decap_8 FILLER_71_391 ();
 sg13g2_decap_8 FILLER_71_398 ();
 sg13g2_decap_4 FILLER_71_405 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_decap_8 FILLER_72_14 ();
 sg13g2_decap_8 FILLER_72_21 ();
 sg13g2_decap_8 FILLER_72_28 ();
 sg13g2_decap_8 FILLER_72_35 ();
 sg13g2_decap_8 FILLER_72_42 ();
 sg13g2_decap_8 FILLER_72_49 ();
 sg13g2_decap_8 FILLER_72_56 ();
 sg13g2_decap_8 FILLER_72_63 ();
 sg13g2_decap_8 FILLER_72_70 ();
 sg13g2_decap_8 FILLER_72_77 ();
 sg13g2_decap_8 FILLER_72_84 ();
 sg13g2_fill_1 FILLER_72_117 ();
 sg13g2_fill_1 FILLER_72_140 ();
 sg13g2_fill_2 FILLER_72_150 ();
 sg13g2_fill_1 FILLER_72_170 ();
 sg13g2_fill_1 FILLER_72_198 ();
 sg13g2_fill_1 FILLER_72_208 ();
 sg13g2_fill_1 FILLER_72_221 ();
 sg13g2_fill_1 FILLER_72_226 ();
 sg13g2_fill_2 FILLER_72_235 ();
 sg13g2_decap_8 FILLER_72_241 ();
 sg13g2_fill_1 FILLER_72_248 ();
 sg13g2_decap_8 FILLER_72_253 ();
 sg13g2_decap_4 FILLER_72_260 ();
 sg13g2_fill_1 FILLER_72_300 ();
 sg13g2_decap_8 FILLER_72_333 ();
 sg13g2_decap_8 FILLER_72_340 ();
 sg13g2_decap_8 FILLER_72_347 ();
 sg13g2_decap_8 FILLER_72_354 ();
 sg13g2_decap_8 FILLER_72_361 ();
 sg13g2_decap_8 FILLER_72_368 ();
 sg13g2_decap_8 FILLER_72_375 ();
 sg13g2_decap_8 FILLER_72_382 ();
 sg13g2_decap_8 FILLER_72_389 ();
 sg13g2_decap_8 FILLER_72_396 ();
 sg13g2_decap_4 FILLER_72_403 ();
 sg13g2_fill_2 FILLER_72_407 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_decap_8 FILLER_73_14 ();
 sg13g2_decap_8 FILLER_73_21 ();
 sg13g2_decap_8 FILLER_73_28 ();
 sg13g2_decap_8 FILLER_73_35 ();
 sg13g2_decap_8 FILLER_73_42 ();
 sg13g2_decap_8 FILLER_73_49 ();
 sg13g2_decap_8 FILLER_73_56 ();
 sg13g2_decap_8 FILLER_73_63 ();
 sg13g2_decap_8 FILLER_73_70 ();
 sg13g2_decap_8 FILLER_73_77 ();
 sg13g2_decap_4 FILLER_73_84 ();
 sg13g2_fill_2 FILLER_73_188 ();
 sg13g2_decap_4 FILLER_73_194 ();
 sg13g2_decap_8 FILLER_73_209 ();
 sg13g2_decap_8 FILLER_73_216 ();
 sg13g2_decap_8 FILLER_73_223 ();
 sg13g2_fill_2 FILLER_73_230 ();
 sg13g2_fill_1 FILLER_73_232 ();
 sg13g2_decap_8 FILLER_73_236 ();
 sg13g2_decap_8 FILLER_73_243 ();
 sg13g2_decap_4 FILLER_73_250 ();
 sg13g2_fill_2 FILLER_73_254 ();
 sg13g2_decap_4 FILLER_73_310 ();
 sg13g2_fill_2 FILLER_73_314 ();
 sg13g2_decap_8 FILLER_73_326 ();
 sg13g2_decap_8 FILLER_73_333 ();
 sg13g2_decap_8 FILLER_73_340 ();
 sg13g2_decap_8 FILLER_73_347 ();
 sg13g2_decap_8 FILLER_73_354 ();
 sg13g2_decap_8 FILLER_73_361 ();
 sg13g2_decap_8 FILLER_73_368 ();
 sg13g2_decap_8 FILLER_73_375 ();
 sg13g2_decap_8 FILLER_73_382 ();
 sg13g2_decap_8 FILLER_73_389 ();
 sg13g2_decap_8 FILLER_73_396 ();
 sg13g2_decap_4 FILLER_73_403 ();
 sg13g2_fill_2 FILLER_73_407 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_decap_8 FILLER_74_14 ();
 sg13g2_decap_8 FILLER_74_21 ();
 sg13g2_decap_8 FILLER_74_28 ();
 sg13g2_decap_8 FILLER_74_35 ();
 sg13g2_decap_8 FILLER_74_42 ();
 sg13g2_decap_8 FILLER_74_49 ();
 sg13g2_decap_8 FILLER_74_56 ();
 sg13g2_decap_8 FILLER_74_63 ();
 sg13g2_decap_8 FILLER_74_70 ();
 sg13g2_decap_8 FILLER_74_77 ();
 sg13g2_decap_4 FILLER_74_84 ();
 sg13g2_fill_2 FILLER_74_88 ();
 sg13g2_fill_1 FILLER_74_120 ();
 sg13g2_decap_8 FILLER_74_208 ();
 sg13g2_fill_2 FILLER_74_258 ();
 sg13g2_decap_8 FILLER_74_311 ();
 sg13g2_decap_8 FILLER_74_318 ();
 sg13g2_decap_8 FILLER_74_325 ();
 sg13g2_decap_8 FILLER_74_332 ();
 sg13g2_decap_8 FILLER_74_339 ();
 sg13g2_decap_8 FILLER_74_346 ();
 sg13g2_decap_8 FILLER_74_353 ();
 sg13g2_decap_8 FILLER_74_360 ();
 sg13g2_decap_8 FILLER_74_367 ();
 sg13g2_decap_8 FILLER_74_374 ();
 sg13g2_decap_8 FILLER_74_381 ();
 sg13g2_decap_8 FILLER_74_388 ();
 sg13g2_decap_8 FILLER_74_395 ();
 sg13g2_decap_8 FILLER_74_402 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_14 ();
 sg13g2_decap_8 FILLER_75_21 ();
 sg13g2_decap_8 FILLER_75_28 ();
 sg13g2_decap_8 FILLER_75_35 ();
 sg13g2_decap_8 FILLER_75_42 ();
 sg13g2_decap_8 FILLER_75_49 ();
 sg13g2_decap_8 FILLER_75_56 ();
 sg13g2_decap_8 FILLER_75_63 ();
 sg13g2_decap_8 FILLER_75_70 ();
 sg13g2_decap_8 FILLER_75_77 ();
 sg13g2_decap_8 FILLER_75_84 ();
 sg13g2_fill_2 FILLER_75_114 ();
 sg13g2_fill_1 FILLER_75_116 ();
 sg13g2_fill_2 FILLER_75_132 ();
 sg13g2_fill_1 FILLER_75_134 ();
 sg13g2_fill_2 FILLER_75_181 ();
 sg13g2_fill_2 FILLER_75_231 ();
 sg13g2_decap_8 FILLER_75_259 ();
 sg13g2_decap_4 FILLER_75_266 ();
 sg13g2_fill_2 FILLER_75_270 ();
 sg13g2_decap_4 FILLER_75_277 ();
 sg13g2_fill_1 FILLER_75_281 ();
 sg13g2_decap_4 FILLER_75_287 ();
 sg13g2_decap_8 FILLER_75_301 ();
 sg13g2_decap_8 FILLER_75_308 ();
 sg13g2_decap_8 FILLER_75_315 ();
 sg13g2_decap_8 FILLER_75_322 ();
 sg13g2_decap_8 FILLER_75_329 ();
 sg13g2_decap_8 FILLER_75_336 ();
 sg13g2_decap_8 FILLER_75_343 ();
 sg13g2_decap_8 FILLER_75_350 ();
 sg13g2_decap_8 FILLER_75_357 ();
 sg13g2_decap_8 FILLER_75_364 ();
 sg13g2_decap_8 FILLER_75_371 ();
 sg13g2_decap_8 FILLER_75_378 ();
 sg13g2_decap_8 FILLER_75_385 ();
 sg13g2_decap_8 FILLER_75_392 ();
 sg13g2_decap_8 FILLER_75_399 ();
 sg13g2_fill_2 FILLER_75_406 ();
 sg13g2_fill_1 FILLER_75_408 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_8 FILLER_76_21 ();
 sg13g2_decap_8 FILLER_76_28 ();
 sg13g2_decap_8 FILLER_76_35 ();
 sg13g2_decap_8 FILLER_76_42 ();
 sg13g2_decap_8 FILLER_76_49 ();
 sg13g2_decap_8 FILLER_76_56 ();
 sg13g2_decap_8 FILLER_76_63 ();
 sg13g2_decap_8 FILLER_76_70 ();
 sg13g2_decap_8 FILLER_76_77 ();
 sg13g2_decap_4 FILLER_76_84 ();
 sg13g2_fill_2 FILLER_76_88 ();
 sg13g2_fill_2 FILLER_76_141 ();
 sg13g2_fill_1 FILLER_76_211 ();
 sg13g2_fill_1 FILLER_76_220 ();
 sg13g2_decap_8 FILLER_76_260 ();
 sg13g2_decap_8 FILLER_76_267 ();
 sg13g2_decap_8 FILLER_76_274 ();
 sg13g2_decap_8 FILLER_76_281 ();
 sg13g2_decap_8 FILLER_76_288 ();
 sg13g2_decap_8 FILLER_76_295 ();
 sg13g2_decap_8 FILLER_76_302 ();
 sg13g2_decap_8 FILLER_76_309 ();
 sg13g2_decap_8 FILLER_76_316 ();
 sg13g2_decap_8 FILLER_76_323 ();
 sg13g2_decap_8 FILLER_76_330 ();
 sg13g2_decap_8 FILLER_76_337 ();
 sg13g2_decap_8 FILLER_76_344 ();
 sg13g2_decap_8 FILLER_76_351 ();
 sg13g2_decap_8 FILLER_76_358 ();
 sg13g2_decap_8 FILLER_76_365 ();
 sg13g2_decap_8 FILLER_76_372 ();
 sg13g2_decap_8 FILLER_76_379 ();
 sg13g2_decap_8 FILLER_76_386 ();
 sg13g2_decap_8 FILLER_76_393 ();
 sg13g2_decap_8 FILLER_76_400 ();
 sg13g2_fill_2 FILLER_76_407 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_decap_8 FILLER_77_28 ();
 sg13g2_decap_8 FILLER_77_35 ();
 sg13g2_decap_8 FILLER_77_42 ();
 sg13g2_decap_8 FILLER_77_49 ();
 sg13g2_decap_8 FILLER_77_56 ();
 sg13g2_decap_8 FILLER_77_63 ();
 sg13g2_decap_8 FILLER_77_70 ();
 sg13g2_decap_8 FILLER_77_77 ();
 sg13g2_decap_8 FILLER_77_84 ();
 sg13g2_decap_8 FILLER_77_91 ();
 sg13g2_fill_1 FILLER_77_98 ();
 sg13g2_fill_2 FILLER_77_185 ();
 sg13g2_decap_4 FILLER_77_213 ();
 sg13g2_fill_1 FILLER_77_217 ();
 sg13g2_fill_2 FILLER_77_237 ();
 sg13g2_fill_1 FILLER_77_239 ();
 sg13g2_decap_8 FILLER_77_266 ();
 sg13g2_decap_8 FILLER_77_273 ();
 sg13g2_decap_8 FILLER_77_280 ();
 sg13g2_decap_8 FILLER_77_287 ();
 sg13g2_decap_8 FILLER_77_294 ();
 sg13g2_decap_8 FILLER_77_301 ();
 sg13g2_decap_8 FILLER_77_308 ();
 sg13g2_decap_8 FILLER_77_315 ();
 sg13g2_decap_8 FILLER_77_322 ();
 sg13g2_decap_8 FILLER_77_329 ();
 sg13g2_decap_8 FILLER_77_336 ();
 sg13g2_decap_8 FILLER_77_343 ();
 sg13g2_decap_8 FILLER_77_350 ();
 sg13g2_decap_8 FILLER_77_357 ();
 sg13g2_decap_8 FILLER_77_364 ();
 sg13g2_decap_8 FILLER_77_371 ();
 sg13g2_decap_8 FILLER_77_378 ();
 sg13g2_decap_8 FILLER_77_385 ();
 sg13g2_decap_8 FILLER_77_392 ();
 sg13g2_decap_8 FILLER_77_399 ();
 sg13g2_fill_2 FILLER_77_406 ();
 sg13g2_fill_1 FILLER_77_408 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_decap_8 FILLER_78_28 ();
 sg13g2_decap_8 FILLER_78_35 ();
 sg13g2_decap_8 FILLER_78_42 ();
 sg13g2_decap_8 FILLER_78_49 ();
 sg13g2_decap_8 FILLER_78_56 ();
 sg13g2_decap_8 FILLER_78_63 ();
 sg13g2_decap_8 FILLER_78_70 ();
 sg13g2_decap_8 FILLER_78_77 ();
 sg13g2_decap_8 FILLER_78_84 ();
 sg13g2_decap_8 FILLER_78_91 ();
 sg13g2_decap_8 FILLER_78_98 ();
 sg13g2_fill_2 FILLER_78_131 ();
 sg13g2_decap_8 FILLER_78_190 ();
 sg13g2_fill_2 FILLER_78_201 ();
 sg13g2_fill_1 FILLER_78_203 ();
 sg13g2_fill_2 FILLER_78_221 ();
 sg13g2_fill_1 FILLER_78_223 ();
 sg13g2_fill_2 FILLER_78_229 ();
 sg13g2_decap_8 FILLER_78_262 ();
 sg13g2_decap_8 FILLER_78_269 ();
 sg13g2_decap_8 FILLER_78_276 ();
 sg13g2_decap_8 FILLER_78_283 ();
 sg13g2_decap_8 FILLER_78_290 ();
 sg13g2_decap_8 FILLER_78_297 ();
 sg13g2_decap_8 FILLER_78_304 ();
 sg13g2_decap_8 FILLER_78_311 ();
 sg13g2_decap_8 FILLER_78_318 ();
 sg13g2_decap_8 FILLER_78_325 ();
 sg13g2_decap_8 FILLER_78_332 ();
 sg13g2_decap_8 FILLER_78_339 ();
 sg13g2_decap_8 FILLER_78_346 ();
 sg13g2_decap_8 FILLER_78_353 ();
 sg13g2_decap_8 FILLER_78_360 ();
 sg13g2_decap_8 FILLER_78_367 ();
 sg13g2_decap_8 FILLER_78_374 ();
 sg13g2_decap_8 FILLER_78_381 ();
 sg13g2_decap_8 FILLER_78_388 ();
 sg13g2_decap_8 FILLER_78_395 ();
 sg13g2_decap_8 FILLER_78_402 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_decap_8 FILLER_79_35 ();
 sg13g2_decap_8 FILLER_79_42 ();
 sg13g2_decap_8 FILLER_79_49 ();
 sg13g2_decap_8 FILLER_79_56 ();
 sg13g2_decap_8 FILLER_79_63 ();
 sg13g2_decap_8 FILLER_79_70 ();
 sg13g2_decap_8 FILLER_79_77 ();
 sg13g2_decap_8 FILLER_79_84 ();
 sg13g2_decap_8 FILLER_79_91 ();
 sg13g2_decap_4 FILLER_79_98 ();
 sg13g2_fill_1 FILLER_79_102 ();
 sg13g2_fill_1 FILLER_79_145 ();
 sg13g2_fill_2 FILLER_79_198 ();
 sg13g2_fill_1 FILLER_79_200 ();
 sg13g2_decap_8 FILLER_79_261 ();
 sg13g2_decap_8 FILLER_79_268 ();
 sg13g2_decap_8 FILLER_79_275 ();
 sg13g2_decap_8 FILLER_79_282 ();
 sg13g2_decap_8 FILLER_79_289 ();
 sg13g2_decap_8 FILLER_79_296 ();
 sg13g2_decap_8 FILLER_79_303 ();
 sg13g2_decap_8 FILLER_79_310 ();
 sg13g2_decap_8 FILLER_79_317 ();
 sg13g2_decap_8 FILLER_79_324 ();
 sg13g2_decap_8 FILLER_79_331 ();
 sg13g2_decap_8 FILLER_79_338 ();
 sg13g2_decap_8 FILLER_79_345 ();
 sg13g2_decap_8 FILLER_79_352 ();
 sg13g2_decap_8 FILLER_79_359 ();
 sg13g2_decap_8 FILLER_79_366 ();
 sg13g2_decap_8 FILLER_79_373 ();
 sg13g2_decap_8 FILLER_79_380 ();
 sg13g2_decap_8 FILLER_79_387 ();
 sg13g2_decap_8 FILLER_79_394 ();
 sg13g2_decap_8 FILLER_79_401 ();
 sg13g2_fill_1 FILLER_79_408 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_42 ();
 sg13g2_decap_8 FILLER_80_49 ();
 sg13g2_decap_4 FILLER_80_60 ();
 sg13g2_decap_4 FILLER_80_68 ();
 sg13g2_decap_4 FILLER_80_76 ();
 sg13g2_decap_4 FILLER_80_84 ();
 sg13g2_fill_2 FILLER_80_156 ();
 sg13g2_fill_2 FILLER_80_174 ();
 sg13g2_decap_8 FILLER_80_192 ();
 sg13g2_decap_8 FILLER_80_199 ();
 sg13g2_decap_4 FILLER_80_206 ();
 sg13g2_fill_1 FILLER_80_210 ();
 sg13g2_decap_8 FILLER_80_215 ();
 sg13g2_decap_8 FILLER_80_222 ();
 sg13g2_decap_8 FILLER_80_238 ();
 sg13g2_decap_8 FILLER_80_245 ();
 sg13g2_decap_8 FILLER_80_252 ();
 sg13g2_decap_8 FILLER_80_259 ();
 sg13g2_decap_8 FILLER_80_266 ();
 sg13g2_decap_8 FILLER_80_273 ();
 sg13g2_decap_8 FILLER_80_280 ();
 sg13g2_decap_8 FILLER_80_287 ();
 sg13g2_decap_8 FILLER_80_294 ();
 sg13g2_decap_8 FILLER_80_301 ();
 sg13g2_decap_8 FILLER_80_308 ();
 sg13g2_decap_8 FILLER_80_315 ();
 sg13g2_decap_8 FILLER_80_322 ();
 sg13g2_decap_8 FILLER_80_329 ();
 sg13g2_decap_8 FILLER_80_336 ();
 sg13g2_decap_8 FILLER_80_343 ();
 sg13g2_decap_8 FILLER_80_350 ();
 sg13g2_decap_8 FILLER_80_357 ();
 sg13g2_decap_8 FILLER_80_364 ();
 sg13g2_decap_4 FILLER_80_371 ();
 sg13g2_fill_1 FILLER_80_375 ();
 sg13g2_decap_8 FILLER_80_381 ();
 sg13g2_decap_8 FILLER_80_388 ();
 sg13g2_decap_8 FILLER_80_395 ();
 sg13g2_decap_8 FILLER_80_402 ();
 assign uio_oe[0] = net2;
 assign uio_oe[1] = net3;
 assign uio_oe[2] = net4;
 assign uio_oe[3] = net5;
 assign uio_oe[4] = net6;
 assign uio_oe[5] = net7;
 assign uio_oe[6] = net8;
 assign uio_oe[7] = net162;
 assign uio_out[0] = net9;
 assign uio_out[1] = net10;
 assign uio_out[2] = net11;
 assign uio_out[3] = net12;
 assign uio_out[4] = net13;
 assign uio_out[5] = net14;
 assign uio_out[6] = net15;
endmodule

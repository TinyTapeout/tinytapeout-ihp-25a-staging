module tt_um_project_tt09 (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire clknet_0_clk;
 wire \div[0] ;
 wire \div[10] ;
 wire \div[11] ;
 wire \div[12] ;
 wire \div[13] ;
 wire \div[14] ;
 wire \div[15] ;
 wire \div[16] ;
 wire \div[17] ;
 wire \div[18] ;
 wire \div[19] ;
 wire \div[1] ;
 wire \div[20] ;
 wire \div[21] ;
 wire \div[22] ;
 wire \div[23] ;
 wire \div[24] ;
 wire \div[25] ;
 wire \div[2] ;
 wire \div[3] ;
 wire \div[4] ;
 wire \div[5] ;
 wire \div[6] ;
 wire \div[7] ;
 wire \div[8] ;
 wire \div[9] ;
 wire indicator;
 wire \lif1.U[0] ;
 wire \lif1.U[1] ;
 wire \lif1.U[2] ;
 wire \lif1.U[3] ;
 wire \lif1.U[4] ;
 wire \lif1.U[5] ;
 wire \lif1.U[6] ;
 wire \lif1.U[7] ;
 wire \lif1.spike ;
 wire \lif1.timer[0] ;
 wire \lif1.timer[1] ;
 wire \lif1.timer[2] ;
 wire \lif1.timer[3] ;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net33;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;

 sg13g2_inv_1 _282_ (.Y(_198_),
    .A(net112));
 sg13g2_inv_1 _283_ (.Y(_199_),
    .A(\lif1.U[4] ));
 sg13g2_inv_1 _284_ (.Y(_200_),
    .A(net32));
 sg13g2_nand4_1 _285_ (.B(\lif1.U[2] ),
    .C(\lif1.U[1] ),
    .A(\lif1.U[3] ),
    .Y(_201_),
    .D(\lif1.U[0] ));
 sg13g2_nand3_1 _286_ (.B(\lif1.U[6] ),
    .C(\lif1.U[5] ),
    .A(\lif1.U[7] ),
    .Y(_202_));
 sg13g2_a21oi_2 _287_ (.B1(_202_),
    .Y(\lif1.spike ),
    .A2(_201_),
    .A1(_199_));
 sg13g2_nand3_1 _288_ (.B(net85),
    .C(net133),
    .A(\div[0] ),
    .Y(_203_));
 sg13g2_and4_2 _289_ (.A(\div[0] ),
    .B(net85),
    .C(net80),
    .D(\div[2] ),
    .X(_204_));
 sg13g2_nand3_1 _290_ (.B(net97),
    .C(_204_),
    .A(net132),
    .Y(_205_));
 sg13g2_and4_1 _291_ (.A(\div[5] ),
    .B(net97),
    .C(net78),
    .D(_204_),
    .X(_041_));
 sg13g2_nor4_1 _292_ (.A(\div[7] ),
    .B(\div[9] ),
    .C(\div[8] ),
    .D(\div[11] ),
    .Y(_042_));
 sg13g2_nor2b_1 _293_ (.A(\div[10] ),
    .B_N(\div[12] ),
    .Y(_043_));
 sg13g2_nand4_1 _294_ (.B(\div[15] ),
    .C(_042_),
    .A(\div[13] ),
    .Y(_044_),
    .D(_043_));
 sg13g2_and4_1 _295_ (.A(\div[21] ),
    .B(\div[20] ),
    .C(\div[22] ),
    .D(\div[23] ),
    .X(_045_));
 sg13g2_nand4_1 _296_ (.B(\div[17] ),
    .C(\div[19] ),
    .A(\div[14] ),
    .Y(_046_),
    .D(\div[25] ));
 sg13g2_nor4_1 _297_ (.A(\div[16] ),
    .B(\div[18] ),
    .C(\div[24] ),
    .D(_046_),
    .Y(_047_));
 sg13g2_nor2b_1 _298_ (.A(_044_),
    .B_N(_047_),
    .Y(_048_));
 sg13g2_and3_1 _299_ (.X(_049_),
    .A(_041_),
    .B(_045_),
    .C(_048_));
 sg13g2_mux2_1 _300_ (.A0(indicator),
    .A1(net73),
    .S(net29),
    .X(_002_));
 sg13g2_nor2b_1 _301_ (.A(net28),
    .B_N(net72),
    .Y(_003_));
 sg13g2_xor2_1 _302_ (.B(net85),
    .A(\div[0] ),
    .X(_004_));
 sg13g2_a21o_1 _303_ (.A2(net85),
    .A1(\div[0] ),
    .B1(net133),
    .X(_050_));
 sg13g2_and2_1 _304_ (.A(_203_),
    .B(net134),
    .X(_005_));
 sg13g2_xnor2_1 _305_ (.Y(_006_),
    .A(net80),
    .B(_203_));
 sg13g2_xor2_1 _306_ (.B(_204_),
    .A(net97),
    .X(_007_));
 sg13g2_a21o_1 _307_ (.A2(_204_),
    .A1(net97),
    .B1(net132),
    .X(_051_));
 sg13g2_and2_1 _308_ (.A(_205_),
    .B(_051_),
    .X(_008_));
 sg13g2_xnor2_1 _309_ (.Y(_009_),
    .A(net78),
    .B(_205_));
 sg13g2_nor2_1 _310_ (.A(net124),
    .B(_041_),
    .Y(_052_));
 sg13g2_and2_1 _311_ (.A(net124),
    .B(_041_),
    .X(_053_));
 sg13g2_nor3_1 _312_ (.A(net28),
    .B(net125),
    .C(_053_),
    .Y(_010_));
 sg13g2_and2_1 _313_ (.A(net95),
    .B(_053_),
    .X(_054_));
 sg13g2_xor2_1 _314_ (.B(_053_),
    .A(net95),
    .X(_011_));
 sg13g2_xor2_1 _315_ (.B(_054_),
    .A(net123),
    .X(_012_));
 sg13g2_a21oi_1 _316_ (.A1(\div[9] ),
    .A2(_054_),
    .Y(_055_),
    .B1(net87));
 sg13g2_nand3_1 _317_ (.B(net87),
    .C(_054_),
    .A(\div[9] ),
    .Y(_056_));
 sg13g2_nor2b_1 _318_ (.A(net88),
    .B_N(_056_),
    .Y(_013_));
 sg13g2_and3_1 _319_ (.X(_057_),
    .A(\div[9] ),
    .B(\div[11] ),
    .C(\div[10] ));
 sg13g2_and4_1 _320_ (.A(net124),
    .B(net95),
    .C(_041_),
    .D(_057_),
    .X(_058_));
 sg13g2_xnor2_1 _321_ (.Y(_014_),
    .A(net93),
    .B(_056_));
 sg13g2_nor2_1 _322_ (.A(net126),
    .B(_058_),
    .Y(_059_));
 sg13g2_and2_1 _323_ (.A(net126),
    .B(_058_),
    .X(_060_));
 sg13g2_nor3_1 _324_ (.A(net28),
    .B(_059_),
    .C(_060_),
    .Y(_015_));
 sg13g2_nor2_1 _325_ (.A(net127),
    .B(_060_),
    .Y(_061_));
 sg13g2_and2_1 _326_ (.A(net127),
    .B(_060_),
    .X(_062_));
 sg13g2_nor3_1 _327_ (.A(net28),
    .B(_061_),
    .C(_062_),
    .Y(_016_));
 sg13g2_nor2_1 _328_ (.A(net118),
    .B(_062_),
    .Y(_063_));
 sg13g2_and4_1 _329_ (.A(\div[13] ),
    .B(\div[12] ),
    .C(net118),
    .D(_058_),
    .X(_064_));
 sg13g2_nor3_1 _330_ (.A(net28),
    .B(net119),
    .C(_064_),
    .Y(_017_));
 sg13g2_nor2_1 _331_ (.A(net121),
    .B(_064_),
    .Y(_065_));
 sg13g2_and2_1 _332_ (.A(net121),
    .B(_064_),
    .X(_066_));
 sg13g2_nor3_1 _333_ (.A(net28),
    .B(net122),
    .C(_066_),
    .Y(_018_));
 sg13g2_xor2_1 _334_ (.B(_066_),
    .A(net99),
    .X(_019_));
 sg13g2_a21oi_1 _335_ (.A1(\div[16] ),
    .A2(_066_),
    .Y(_067_),
    .B1(net82));
 sg13g2_and4_2 _336_ (.A(\div[15] ),
    .B(net99),
    .C(net82),
    .D(_064_),
    .X(_068_));
 sg13g2_nor3_1 _337_ (.A(net28),
    .B(net83),
    .C(_068_),
    .Y(_020_));
 sg13g2_xor2_1 _338_ (.B(_068_),
    .A(net110),
    .X(_021_));
 sg13g2_a21oi_1 _339_ (.A1(\div[18] ),
    .A2(_068_),
    .Y(_069_),
    .B1(net105));
 sg13g2_and3_2 _340_ (.X(_070_),
    .A(net110),
    .B(net105),
    .C(_068_));
 sg13g2_nor3_1 _341_ (.A(net29),
    .B(net106),
    .C(_070_),
    .Y(_022_));
 sg13g2_nor2_1 _342_ (.A(net128),
    .B(_070_),
    .Y(_071_));
 sg13g2_and2_1 _343_ (.A(net128),
    .B(_070_),
    .X(_072_));
 sg13g2_nor3_1 _344_ (.A(net29),
    .B(_071_),
    .C(_072_),
    .Y(_023_));
 sg13g2_nor2_1 _345_ (.A(net115),
    .B(_072_),
    .Y(_073_));
 sg13g2_and3_1 _346_ (.X(_074_),
    .A(net115),
    .B(\div[20] ),
    .C(_070_));
 sg13g2_nor3_1 _347_ (.A(net29),
    .B(net116),
    .C(_074_),
    .Y(_024_));
 sg13g2_nor2_1 _348_ (.A(net102),
    .B(_074_),
    .Y(_075_));
 sg13g2_and4_1 _349_ (.A(net143),
    .B(\div[20] ),
    .C(net102),
    .D(_070_),
    .X(_076_));
 sg13g2_nor3_1 _350_ (.A(net29),
    .B(net103),
    .C(_076_),
    .Y(_025_));
 sg13g2_nor2_1 _351_ (.A(net108),
    .B(_076_),
    .Y(_077_));
 sg13g2_and2_1 _352_ (.A(net108),
    .B(_076_),
    .X(_078_));
 sg13g2_nor3_1 _353_ (.A(net28),
    .B(net109),
    .C(_078_),
    .Y(_026_));
 sg13g2_and2_1 _354_ (.A(\div[24] ),
    .B(_045_),
    .X(_079_));
 sg13g2_and4_2 _355_ (.A(net110),
    .B(net105),
    .C(_068_),
    .D(_079_),
    .X(_080_));
 sg13g2_a21oi_1 _356_ (.A1(_045_),
    .A2(_070_),
    .Y(_081_),
    .B1(net75));
 sg13g2_nor2_1 _357_ (.A(_080_),
    .B(net76),
    .Y(_027_));
 sg13g2_nor2_1 _358_ (.A(net130),
    .B(_080_),
    .Y(_082_));
 sg13g2_and2_1 _359_ (.A(\div[25] ),
    .B(_080_),
    .X(_083_));
 sg13g2_nand2_2 _360_ (.Y(_084_),
    .A(net130),
    .B(_080_));
 sg13g2_nor3_1 _361_ (.A(net29),
    .B(_082_),
    .C(net27),
    .Y(_028_));
 sg13g2_or2_1 _362_ (.X(_085_),
    .B(\lif1.timer[1] ),
    .A(net90));
 sg13g2_nor3_2 _363_ (.A(\lif1.timer[3] ),
    .B(\lif1.timer[0] ),
    .C(_085_),
    .Y(_086_));
 sg13g2_and2_2 _364_ (.A(\lif1.spike ),
    .B(_086_),
    .X(_087_));
 sg13g2_nand2_1 _365_ (.Y(_088_),
    .A(\lif1.spike ),
    .B(_086_));
 sg13g2_nor2_1 _366_ (.A(\lif1.U[1] ),
    .B(_087_),
    .Y(_089_));
 sg13g2_a21oi_1 _367_ (.A1(net131),
    .A2(_087_),
    .Y(_090_),
    .B1(_089_));
 sg13g2_xnor2_1 _368_ (.Y(_091_),
    .A(net2),
    .B(_090_));
 sg13g2_o21ai_1 _369_ (.B1(net1),
    .Y(_092_),
    .A1(net131),
    .A2(net27));
 sg13g2_a21oi_1 _370_ (.A1(net27),
    .A2(_091_),
    .Y(_029_),
    .B1(_092_));
 sg13g2_nor2_2 _371_ (.A(\lif1.U[0] ),
    .B(net2),
    .Y(_093_));
 sg13g2_and2_1 _372_ (.A(\lif1.U[1] ),
    .B(net3),
    .X(_094_));
 sg13g2_nand2_1 _373_ (.Y(_095_),
    .A(\lif1.U[1] ),
    .B(net3));
 sg13g2_nor2_1 _374_ (.A(\lif1.U[1] ),
    .B(net3),
    .Y(_096_));
 sg13g2_nor2_1 _375_ (.A(_094_),
    .B(_096_),
    .Y(_097_));
 sg13g2_nand2b_1 _376_ (.Y(_098_),
    .B(_097_),
    .A_N(_093_));
 sg13g2_xnor2_1 _377_ (.Y(_099_),
    .A(_093_),
    .B(_097_));
 sg13g2_nand2_1 _378_ (.Y(_100_),
    .A(\lif1.U[1] ),
    .B(net2));
 sg13g2_nand2_1 _379_ (.Y(_101_),
    .A(\lif1.U[2] ),
    .B(net3));
 sg13g2_xnor2_1 _380_ (.Y(_102_),
    .A(\lif1.U[2] ),
    .B(net3));
 sg13g2_or2_1 _381_ (.X(_103_),
    .B(_102_),
    .A(_100_));
 sg13g2_a21oi_1 _382_ (.A1(_100_),
    .A2(_102_),
    .Y(_104_),
    .B1(_087_));
 sg13g2_a22oi_1 _383_ (.Y(_105_),
    .B1(_103_),
    .B2(_104_),
    .A2(_099_),
    .A1(_087_));
 sg13g2_o21ai_1 _384_ (.B1(net32),
    .Y(_106_),
    .A1(net138),
    .A2(net26));
 sg13g2_a21oi_1 _385_ (.A1(net26),
    .A2(_105_),
    .Y(_030_),
    .B1(_106_));
 sg13g2_and2_1 _386_ (.A(\lif1.U[3] ),
    .B(net4),
    .X(_107_));
 sg13g2_or2_1 _387_ (.X(_108_),
    .B(net4),
    .A(\lif1.U[3] ));
 sg13g2_nor2b_1 _388_ (.A(_107_),
    .B_N(_108_),
    .Y(_109_));
 sg13g2_o21ai_1 _389_ (.B1(_101_),
    .Y(_110_),
    .A1(_100_),
    .A2(_102_));
 sg13g2_nand2_1 _390_ (.Y(_111_),
    .A(\lif1.U[2] ),
    .B(net4));
 sg13g2_xnor2_1 _391_ (.Y(_112_),
    .A(\lif1.U[2] ),
    .B(net4));
 sg13g2_nor2_1 _392_ (.A(_095_),
    .B(_112_),
    .Y(_113_));
 sg13g2_xnor2_1 _393_ (.Y(_114_),
    .A(_094_),
    .B(_112_));
 sg13g2_nor4_2 _394_ (.A(_093_),
    .B(_094_),
    .C(_096_),
    .Y(_115_),
    .D(_112_));
 sg13g2_xnor2_1 _395_ (.Y(_116_),
    .A(_098_),
    .B(_114_));
 sg13g2_xnor2_1 _396_ (.Y(_117_),
    .A(_109_),
    .B(_110_));
 sg13g2_nand2_1 _397_ (.Y(_118_),
    .A(_088_),
    .B(_117_));
 sg13g2_o21ai_1 _398_ (.B1(_118_),
    .Y(_119_),
    .A1(_088_),
    .A2(_116_));
 sg13g2_o21ai_1 _399_ (.B1(net32),
    .Y(_120_),
    .A1(net139),
    .A2(net26));
 sg13g2_a21oi_1 _400_ (.A1(net26),
    .A2(_119_),
    .Y(_031_),
    .B1(_120_));
 sg13g2_nand2_1 _401_ (.Y(_121_),
    .A(\lif1.U[4] ),
    .B(net5));
 sg13g2_nor2_1 _402_ (.A(\lif1.U[4] ),
    .B(net5),
    .Y(_122_));
 sg13g2_xor2_1 _403_ (.B(net5),
    .A(\lif1.U[4] ),
    .X(_123_));
 sg13g2_a21oi_1 _404_ (.A1(_108_),
    .A2(_110_),
    .Y(_124_),
    .B1(_107_));
 sg13g2_xnor2_1 _405_ (.Y(_125_),
    .A(_123_),
    .B(_124_));
 sg13g2_nand2_1 _406_ (.Y(_126_),
    .A(\lif1.U[3] ),
    .B(net5));
 sg13g2_xor2_1 _407_ (.B(net5),
    .A(\lif1.U[3] ),
    .X(_127_));
 sg13g2_xnor2_1 _408_ (.Y(_128_),
    .A(_111_),
    .B(_127_));
 sg13g2_o21ai_1 _409_ (.B1(_128_),
    .Y(_129_),
    .A1(_113_),
    .A2(_115_));
 sg13g2_nor3_1 _410_ (.A(_113_),
    .B(_115_),
    .C(_128_),
    .Y(_130_));
 sg13g2_nor2_1 _411_ (.A(net30),
    .B(_130_),
    .Y(_131_));
 sg13g2_a22oi_1 _412_ (.Y(_132_),
    .B1(_129_),
    .B2(_131_),
    .A2(_125_),
    .A1(net30));
 sg13g2_o21ai_1 _413_ (.B1(net32),
    .Y(_133_),
    .A1(net137),
    .A2(net26));
 sg13g2_a21oi_1 _414_ (.A1(net26),
    .A2(_132_),
    .Y(_032_),
    .B1(_133_));
 sg13g2_and2_1 _415_ (.A(\lif1.U[5] ),
    .B(net6),
    .X(_134_));
 sg13g2_xor2_1 _416_ (.B(net6),
    .A(\lif1.U[5] ),
    .X(_135_));
 sg13g2_o21ai_1 _417_ (.B1(_121_),
    .Y(_136_),
    .A1(_122_),
    .A2(_124_));
 sg13g2_xor2_1 _418_ (.B(_136_),
    .A(_135_),
    .X(_137_));
 sg13g2_o21ai_1 _419_ (.B1(_111_),
    .Y(_138_),
    .A1(_095_),
    .A2(_112_));
 sg13g2_a22oi_1 _420_ (.Y(_139_),
    .B1(_138_),
    .B2(_127_),
    .A2(_128_),
    .A1(_115_));
 sg13g2_nor2_1 _421_ (.A(\lif1.U[4] ),
    .B(net6),
    .Y(_140_));
 sg13g2_xor2_1 _422_ (.B(net6),
    .A(\lif1.U[4] ),
    .X(_141_));
 sg13g2_or2_1 _423_ (.X(_142_),
    .B(_141_),
    .A(_126_));
 sg13g2_xnor2_1 _424_ (.Y(_143_),
    .A(_126_),
    .B(_141_));
 sg13g2_nor2_1 _425_ (.A(_139_),
    .B(_143_),
    .Y(_144_));
 sg13g2_inv_1 _426_ (.Y(_145_),
    .A(_144_));
 sg13g2_a21oi_1 _427_ (.A1(_139_),
    .A2(_143_),
    .Y(_146_),
    .B1(net30));
 sg13g2_a22oi_1 _428_ (.Y(_147_),
    .B1(_145_),
    .B2(_146_),
    .A2(_137_),
    .A1(net30));
 sg13g2_o21ai_1 _429_ (.B1(net32),
    .Y(_148_),
    .A1(net142),
    .A2(net26));
 sg13g2_a21oi_1 _430_ (.A1(net26),
    .A2(_147_),
    .Y(_033_),
    .B1(_148_));
 sg13g2_nand2_1 _431_ (.Y(_149_),
    .A(\lif1.U[5] ),
    .B(net7));
 sg13g2_xor2_1 _432_ (.B(net7),
    .A(\lif1.U[5] ),
    .X(_150_));
 sg13g2_nor2b_1 _433_ (.A(_150_),
    .B_N(_140_),
    .Y(_151_));
 sg13g2_nor2b_1 _434_ (.A(_140_),
    .B_N(_150_),
    .Y(_152_));
 sg13g2_or2_1 _435_ (.X(_153_),
    .B(_152_),
    .A(_151_));
 sg13g2_a21oi_1 _436_ (.A1(_135_),
    .A2(_136_),
    .Y(_154_),
    .B1(_134_));
 sg13g2_nor2_1 _437_ (.A(\lif1.U[6] ),
    .B(net7),
    .Y(_155_));
 sg13g2_xor2_1 _438_ (.B(net7),
    .A(\lif1.U[6] ),
    .X(_156_));
 sg13g2_xnor2_1 _439_ (.Y(_157_),
    .A(_154_),
    .B(_156_));
 sg13g2_nand3_1 _440_ (.B(_145_),
    .C(_153_),
    .A(_142_),
    .Y(_158_));
 sg13g2_a21oi_1 _441_ (.A1(_142_),
    .A2(_145_),
    .Y(_159_),
    .B1(_153_));
 sg13g2_nor2_1 _442_ (.A(net30),
    .B(_159_),
    .Y(_160_));
 sg13g2_a221oi_1 _443_ (.B2(_160_),
    .C1(_084_),
    .B1(_158_),
    .A1(net30),
    .Y(_161_),
    .A2(_157_));
 sg13g2_o21ai_1 _444_ (.B1(net32),
    .Y(_162_),
    .A1(net140),
    .A2(net27));
 sg13g2_nor2_1 _445_ (.A(_161_),
    .B(_162_),
    .Y(_034_));
 sg13g2_and2_1 _446_ (.A(\lif1.U[7] ),
    .B(net8),
    .X(_163_));
 sg13g2_xnor2_1 _447_ (.Y(_164_),
    .A(\lif1.U[7] ),
    .B(net8));
 sg13g2_a221oi_1 _448_ (.B2(_136_),
    .C1(_134_),
    .B1(_135_),
    .A1(\lif1.U[6] ),
    .Y(_165_),
    .A2(net7));
 sg13g2_or2_1 _449_ (.X(_166_),
    .B(_165_),
    .A(_155_));
 sg13g2_nor3_1 _450_ (.A(_155_),
    .B(_164_),
    .C(_165_),
    .Y(_167_));
 sg13g2_a221oi_1 _451_ (.B2(_166_),
    .C1(_167_),
    .B1(_164_),
    .A1(\lif1.spike ),
    .Y(_168_),
    .A2(_086_));
 sg13g2_nor3_1 _452_ (.A(_139_),
    .B(_143_),
    .C(_153_),
    .Y(_169_));
 sg13g2_nor2_1 _453_ (.A(_142_),
    .B(_151_),
    .Y(_170_));
 sg13g2_or2_1 _454_ (.X(_171_),
    .B(_170_),
    .A(_152_));
 sg13g2_nand2_1 _455_ (.Y(_172_),
    .A(\lif1.U[6] ),
    .B(net8));
 sg13g2_xor2_1 _456_ (.B(net8),
    .A(\lif1.U[6] ),
    .X(_173_));
 sg13g2_xnor2_1 _457_ (.Y(_174_),
    .A(_149_),
    .B(_173_));
 sg13g2_or3_1 _458_ (.A(_169_),
    .B(_171_),
    .C(_174_),
    .X(_175_));
 sg13g2_o21ai_1 _459_ (.B1(_174_),
    .Y(_176_),
    .A1(_169_),
    .A2(_171_));
 sg13g2_and3_1 _460_ (.X(_177_),
    .A(_087_),
    .B(_175_),
    .C(_176_));
 sg13g2_nor3_1 _461_ (.A(_084_),
    .B(_168_),
    .C(_177_),
    .Y(_178_));
 sg13g2_o21ai_1 _462_ (.B1(net32),
    .Y(_179_),
    .A1(net141),
    .A2(net27));
 sg13g2_nor2_1 _463_ (.A(_178_),
    .B(_179_),
    .Y(_035_));
 sg13g2_o21ai_1 _464_ (.B1(net9),
    .Y(_180_),
    .A1(_163_),
    .A2(_167_));
 sg13g2_or3_1 _465_ (.A(net9),
    .B(_163_),
    .C(_167_),
    .X(_181_));
 sg13g2_nand3_1 _466_ (.B(_180_),
    .C(_181_),
    .A(net30),
    .Y(_182_));
 sg13g2_nand3_1 _467_ (.B(_175_),
    .C(_176_),
    .A(net8),
    .Y(_183_));
 sg13g2_xor2_1 _468_ (.B(net9),
    .A(\lif1.U[7] ),
    .X(_184_));
 sg13g2_xnor2_1 _469_ (.Y(_185_),
    .A(_172_),
    .B(_184_));
 sg13g2_or2_1 _470_ (.X(_186_),
    .B(_185_),
    .A(_183_));
 sg13g2_a21oi_1 _471_ (.A1(_183_),
    .A2(_185_),
    .Y(_187_),
    .B1(net30));
 sg13g2_o21ai_1 _472_ (.B1(net32),
    .Y(_188_),
    .A1(net136),
    .A2(net27));
 sg13g2_a21oi_1 _473_ (.A1(_186_),
    .A2(_187_),
    .Y(_189_),
    .B1(_084_));
 sg13g2_a21oi_1 _474_ (.A1(_182_),
    .A2(_189_),
    .Y(_036_),
    .B1(_188_));
 sg13g2_nand2b_1 _475_ (.Y(_190_),
    .B(_086_),
    .A_N(net31));
 sg13g2_nand4_1 _476_ (.B(\div[25] ),
    .C(_080_),
    .A(_198_),
    .Y(_191_),
    .D(_190_));
 sg13g2_nand2_1 _477_ (.Y(_192_),
    .A(net112),
    .B(_084_));
 sg13g2_a21oi_1 _478_ (.A1(_191_),
    .A2(net113),
    .Y(_037_),
    .B1(_200_));
 sg13g2_xor2_1 _479_ (.B(_191_),
    .A(net129),
    .X(_193_));
 sg13g2_nor2_1 _480_ (.A(_200_),
    .B(_193_),
    .Y(_038_));
 sg13g2_o21ai_1 _481_ (.B1(net90),
    .Y(_194_),
    .A1(\lif1.timer[1] ),
    .A2(_191_));
 sg13g2_or2_1 _482_ (.X(_195_),
    .B(_191_),
    .A(_085_));
 sg13g2_a21oi_1 _483_ (.A1(net91),
    .A2(_195_),
    .Y(_039_),
    .B1(_200_));
 sg13g2_o21ai_1 _484_ (.B1(net101),
    .Y(_196_),
    .A1(_085_),
    .A2(_191_));
 sg13g2_nand2_1 _485_ (.Y(_197_),
    .A(net27),
    .B(_087_));
 sg13g2_a21oi_1 _486_ (.A1(_196_),
    .A2(_197_),
    .Y(_040_),
    .B1(_200_));
 sg13g2_dfrbp_1 _487_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net59),
    .D(net74),
    .Q_N(_000_),
    .Q(indicator));
 sg13g2_dfrbp_1 _488_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net55),
    .D(_003_),
    .Q_N(_001_),
    .Q(\div[0] ));
 sg13g2_dfrbp_1 _489_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net54),
    .D(net86),
    .Q_N(_242_),
    .Q(\div[1] ));
 sg13g2_dfrbp_1 _490_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net53),
    .D(net135),
    .Q_N(_241_),
    .Q(\div[2] ));
 sg13g2_dfrbp_1 _491_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net52),
    .D(net81),
    .Q_N(_240_),
    .Q(\div[3] ));
 sg13g2_dfrbp_1 _492_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net51),
    .D(net98),
    .Q_N(_239_),
    .Q(\div[4] ));
 sg13g2_dfrbp_1 _493_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net50),
    .D(_008_),
    .Q_N(_238_),
    .Q(\div[5] ));
 sg13g2_dfrbp_1 _494_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net49),
    .D(net79),
    .Q_N(_237_),
    .Q(\div[6] ));
 sg13g2_dfrbp_1 _495_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net48),
    .D(_010_),
    .Q_N(_236_),
    .Q(\div[7] ));
 sg13g2_dfrbp_1 _496_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net47),
    .D(net96),
    .Q_N(_235_),
    .Q(\div[8] ));
 sg13g2_dfrbp_1 _497_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net46),
    .D(_012_),
    .Q_N(_234_),
    .Q(\div[9] ));
 sg13g2_dfrbp_1 _498_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net45),
    .D(net89),
    .Q_N(_233_),
    .Q(\div[10] ));
 sg13g2_dfrbp_1 _499_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net44),
    .D(net94),
    .Q_N(_232_),
    .Q(\div[11] ));
 sg13g2_dfrbp_1 _500_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net43),
    .D(_015_),
    .Q_N(_231_),
    .Q(\div[12] ));
 sg13g2_dfrbp_1 _501_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net42),
    .D(_016_),
    .Q_N(_230_),
    .Q(\div[13] ));
 sg13g2_dfrbp_1 _502_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net41),
    .D(net120),
    .Q_N(_229_),
    .Q(\div[14] ));
 sg13g2_dfrbp_1 _503_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net40),
    .D(_018_),
    .Q_N(_228_),
    .Q(\div[15] ));
 sg13g2_dfrbp_1 _504_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net39),
    .D(net100),
    .Q_N(_227_),
    .Q(\div[16] ));
 sg13g2_dfrbp_1 _505_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net38),
    .D(net84),
    .Q_N(_226_),
    .Q(\div[17] ));
 sg13g2_dfrbp_1 _506_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net37),
    .D(net111),
    .Q_N(_225_),
    .Q(\div[18] ));
 sg13g2_dfrbp_1 _507_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net36),
    .D(net107),
    .Q_N(_224_),
    .Q(\div[19] ));
 sg13g2_dfrbp_1 _508_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net35),
    .D(_023_),
    .Q_N(_223_),
    .Q(\div[20] ));
 sg13g2_dfrbp_1 _509_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net34),
    .D(net117),
    .Q_N(_222_),
    .Q(\div[21] ));
 sg13g2_dfrbp_1 _510_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net33),
    .D(net104),
    .Q_N(_221_),
    .Q(\div[22] ));
 sg13g2_dfrbp_1 _511_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net71),
    .D(_026_),
    .Q_N(_220_),
    .Q(\div[23] ));
 sg13g2_dfrbp_1 _512_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net70),
    .D(net77),
    .Q_N(_219_),
    .Q(\div[24] ));
 sg13g2_dfrbp_1 _513_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net69),
    .D(_028_),
    .Q_N(_218_),
    .Q(\div[25] ));
 sg13g2_dfrbp_1 _514_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net68),
    .D(_029_),
    .Q_N(_217_),
    .Q(\lif1.U[0] ));
 sg13g2_dfrbp_1 _515_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net66),
    .D(_030_),
    .Q_N(_216_),
    .Q(\lif1.U[1] ));
 sg13g2_dfrbp_1 _516_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net64),
    .D(_031_),
    .Q_N(_215_),
    .Q(\lif1.U[2] ));
 sg13g2_dfrbp_1 _517_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net62),
    .D(_032_),
    .Q_N(_214_),
    .Q(\lif1.U[3] ));
 sg13g2_dfrbp_1 _518_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net60),
    .D(_033_),
    .Q_N(_213_),
    .Q(\lif1.U[4] ));
 sg13g2_dfrbp_1 _519_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net58),
    .D(_034_),
    .Q_N(_212_),
    .Q(\lif1.U[5] ));
 sg13g2_dfrbp_1 _520_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net56),
    .D(_035_),
    .Q_N(_211_),
    .Q(\lif1.U[6] ));
 sg13g2_dfrbp_1 _521_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net65),
    .D(_036_),
    .Q_N(_210_),
    .Q(\lif1.U[7] ));
 sg13g2_dfrbp_1 _522_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net61),
    .D(net114),
    .Q_N(_209_),
    .Q(\lif1.timer[0] ));
 sg13g2_dfrbp_1 _523_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net57),
    .D(_038_),
    .Q_N(_208_),
    .Q(\lif1.timer[1] ));
 sg13g2_dfrbp_1 _524_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net63),
    .D(net92),
    .Q_N(_207_),
    .Q(\lif1.timer[2] ));
 sg13g2_dfrbp_1 _525_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net67),
    .D(_040_),
    .Q_N(_206_),
    .Q(\lif1.timer[3] ));
 sg13g2_tiehi _509__27 (.L_HI(net34));
 sg13g2_tiehi _508__28 (.L_HI(net35));
 sg13g2_tiehi _507__29 (.L_HI(net36));
 sg13g2_tiehi _506__30 (.L_HI(net37));
 sg13g2_tiehi _505__31 (.L_HI(net38));
 sg13g2_tiehi _504__32 (.L_HI(net39));
 sg13g2_tiehi _503__33 (.L_HI(net40));
 sg13g2_tiehi _502__34 (.L_HI(net41));
 sg13g2_tiehi _501__35 (.L_HI(net42));
 sg13g2_tiehi _500__36 (.L_HI(net43));
 sg13g2_tiehi _499__37 (.L_HI(net44));
 sg13g2_tiehi _498__38 (.L_HI(net45));
 sg13g2_tiehi _497__39 (.L_HI(net46));
 sg13g2_tiehi _496__40 (.L_HI(net47));
 sg13g2_tiehi _495__41 (.L_HI(net48));
 sg13g2_tiehi _494__42 (.L_HI(net49));
 sg13g2_tiehi _493__43 (.L_HI(net50));
 sg13g2_tiehi _492__44 (.L_HI(net51));
 sg13g2_tiehi _491__45 (.L_HI(net52));
 sg13g2_tiehi _490__46 (.L_HI(net53));
 sg13g2_tiehi _489__47 (.L_HI(net54));
 sg13g2_tiehi _488__48 (.L_HI(net55));
 sg13g2_tiehi _520__49 (.L_HI(net56));
 sg13g2_tiehi _523__50 (.L_HI(net57));
 sg13g2_tiehi _519__51 (.L_HI(net58));
 sg13g2_tiehi _487__52 (.L_HI(net59));
 sg13g2_tiehi _518__53 (.L_HI(net60));
 sg13g2_tiehi _522__54 (.L_HI(net61));
 sg13g2_tiehi _517__55 (.L_HI(net62));
 sg13g2_tiehi _524__56 (.L_HI(net63));
 sg13g2_tiehi _516__57 (.L_HI(net64));
 sg13g2_tiehi _521__58 (.L_HI(net65));
 sg13g2_tiehi _515__59 (.L_HI(net66));
 sg13g2_tiehi _525__60 (.L_HI(net67));
 sg13g2_tiehi _514__61 (.L_HI(net68));
 sg13g2_tiehi _513__62 (.L_HI(net69));
 sg13g2_tiehi _512__63 (.L_HI(net70));
 sg13g2_tiehi _511__64 (.L_HI(net71));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_project_tt09_11 (.L_LO(net11));
 sg13g2_tielo tt_um_project_tt09_12 (.L_LO(net12));
 sg13g2_tielo tt_um_project_tt09_13 (.L_LO(net13));
 sg13g2_tielo tt_um_project_tt09_14 (.L_LO(net14));
 sg13g2_tielo tt_um_project_tt09_15 (.L_LO(net15));
 sg13g2_tielo tt_um_project_tt09_16 (.L_LO(net16));
 sg13g2_tielo tt_um_project_tt09_17 (.L_LO(net17));
 sg13g2_tielo tt_um_project_tt09_18 (.L_LO(net18));
 sg13g2_tielo tt_um_project_tt09_19 (.L_LO(net19));
 sg13g2_tielo tt_um_project_tt09_20 (.L_LO(net20));
 sg13g2_tielo tt_um_project_tt09_21 (.L_LO(net21));
 sg13g2_tielo tt_um_project_tt09_22 (.L_LO(net22));
 sg13g2_tielo tt_um_project_tt09_23 (.L_LO(net23));
 sg13g2_tielo tt_um_project_tt09_24 (.L_LO(net24));
 sg13g2_tielo tt_um_project_tt09_25 (.L_LO(net25));
 sg13g2_tiehi _510__26 (.L_HI(net33));
 sg13g2_buf_1 _581_ (.A(net31),
    .X(uo_out[0]));
 sg13g2_buf_1 _582_ (.A(net31),
    .X(uo_out[1]));
 sg13g2_buf_1 _583_ (.A(net31),
    .X(uo_out[2]));
 sg13g2_buf_1 _584_ (.A(net31),
    .X(uo_out[3]));
 sg13g2_buf_1 _585_ (.A(net31),
    .X(uo_out[4]));
 sg13g2_buf_1 _586_ (.A(net31),
    .X(uo_out[5]));
 sg13g2_buf_1 _587_ (.A(net31),
    .X(uo_out[6]));
 sg13g2_buf_1 _588_ (.A(indicator),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout26 (.A(net27),
    .X(net26));
 sg13g2_buf_2 fanout27 (.A(_083_),
    .X(net27));
 sg13g2_buf_2 fanout28 (.A(_049_),
    .X(net28));
 sg13g2_buf_2 fanout29 (.A(_049_),
    .X(net29));
 sg13g2_buf_2 fanout30 (.A(_088_),
    .X(net30));
 sg13g2_buf_2 fanout31 (.A(\lif1.spike ),
    .X(net31));
 sg13g2_buf_2 fanout32 (.A(net1),
    .X(net32));
 sg13g2_buf_1 input1 (.A(rst_n),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[0]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[1]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[2]),
    .X(net4));
 sg13g2_buf_2 input5 (.A(ui_in[3]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[4]),
    .X(net6));
 sg13g2_buf_2 input7 (.A(ui_in[5]),
    .X(net7));
 sg13g2_buf_2 input8 (.A(ui_in[6]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(ui_in[7]),
    .X(net9));
 sg13g2_tielo tt_um_project_tt09_10 (.L_LO(net10));
 sg13g2_buf_2 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sg13g2_buf_2 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sg13g2_buf_2 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sg13g2_buf_2 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sg13g2_buf_2 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sg13g2_buf_2 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sg13g2_buf_2 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sg13g2_buf_2 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_3_7__leaf_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(_001_),
    .X(net72));
 sg13g2_dlygate4sd3_1 hold2 (.A(_000_),
    .X(net73));
 sg13g2_dlygate4sd3_1 hold3 (.A(_002_),
    .X(net74));
 sg13g2_dlygate4sd3_1 hold4 (.A(\div[24] ),
    .X(net75));
 sg13g2_dlygate4sd3_1 hold5 (.A(_081_),
    .X(net76));
 sg13g2_dlygate4sd3_1 hold6 (.A(_027_),
    .X(net77));
 sg13g2_dlygate4sd3_1 hold7 (.A(\div[6] ),
    .X(net78));
 sg13g2_dlygate4sd3_1 hold8 (.A(_009_),
    .X(net79));
 sg13g2_dlygate4sd3_1 hold9 (.A(\div[3] ),
    .X(net80));
 sg13g2_dlygate4sd3_1 hold10 (.A(_006_),
    .X(net81));
 sg13g2_dlygate4sd3_1 hold11 (.A(\div[17] ),
    .X(net82));
 sg13g2_dlygate4sd3_1 hold12 (.A(_067_),
    .X(net83));
 sg13g2_dlygate4sd3_1 hold13 (.A(_020_),
    .X(net84));
 sg13g2_dlygate4sd3_1 hold14 (.A(\div[1] ),
    .X(net85));
 sg13g2_dlygate4sd3_1 hold15 (.A(_004_),
    .X(net86));
 sg13g2_dlygate4sd3_1 hold16 (.A(\div[10] ),
    .X(net87));
 sg13g2_dlygate4sd3_1 hold17 (.A(_055_),
    .X(net88));
 sg13g2_dlygate4sd3_1 hold18 (.A(_013_),
    .X(net89));
 sg13g2_dlygate4sd3_1 hold19 (.A(\lif1.timer[2] ),
    .X(net90));
 sg13g2_dlygate4sd3_1 hold20 (.A(_194_),
    .X(net91));
 sg13g2_dlygate4sd3_1 hold21 (.A(_039_),
    .X(net92));
 sg13g2_dlygate4sd3_1 hold22 (.A(\div[11] ),
    .X(net93));
 sg13g2_dlygate4sd3_1 hold23 (.A(_014_),
    .X(net94));
 sg13g2_dlygate4sd3_1 hold24 (.A(\div[8] ),
    .X(net95));
 sg13g2_dlygate4sd3_1 hold25 (.A(_011_),
    .X(net96));
 sg13g2_dlygate4sd3_1 hold26 (.A(\div[4] ),
    .X(net97));
 sg13g2_dlygate4sd3_1 hold27 (.A(_007_),
    .X(net98));
 sg13g2_dlygate4sd3_1 hold28 (.A(\div[16] ),
    .X(net99));
 sg13g2_dlygate4sd3_1 hold29 (.A(_019_),
    .X(net100));
 sg13g2_dlygate4sd3_1 hold30 (.A(\lif1.timer[3] ),
    .X(net101));
 sg13g2_dlygate4sd3_1 hold31 (.A(\div[22] ),
    .X(net102));
 sg13g2_dlygate4sd3_1 hold32 (.A(_075_),
    .X(net103));
 sg13g2_dlygate4sd3_1 hold33 (.A(_025_),
    .X(net104));
 sg13g2_dlygate4sd3_1 hold34 (.A(\div[19] ),
    .X(net105));
 sg13g2_dlygate4sd3_1 hold35 (.A(_069_),
    .X(net106));
 sg13g2_dlygate4sd3_1 hold36 (.A(_022_),
    .X(net107));
 sg13g2_dlygate4sd3_1 hold37 (.A(\div[23] ),
    .X(net108));
 sg13g2_dlygate4sd3_1 hold38 (.A(_077_),
    .X(net109));
 sg13g2_dlygate4sd3_1 hold39 (.A(\div[18] ),
    .X(net110));
 sg13g2_dlygate4sd3_1 hold40 (.A(_021_),
    .X(net111));
 sg13g2_dlygate4sd3_1 hold41 (.A(\lif1.timer[0] ),
    .X(net112));
 sg13g2_dlygate4sd3_1 hold42 (.A(_192_),
    .X(net113));
 sg13g2_dlygate4sd3_1 hold43 (.A(_037_),
    .X(net114));
 sg13g2_dlygate4sd3_1 hold44 (.A(\div[21] ),
    .X(net115));
 sg13g2_dlygate4sd3_1 hold45 (.A(_073_),
    .X(net116));
 sg13g2_dlygate4sd3_1 hold46 (.A(_024_),
    .X(net117));
 sg13g2_dlygate4sd3_1 hold47 (.A(\div[14] ),
    .X(net118));
 sg13g2_dlygate4sd3_1 hold48 (.A(_063_),
    .X(net119));
 sg13g2_dlygate4sd3_1 hold49 (.A(_017_),
    .X(net120));
 sg13g2_dlygate4sd3_1 hold50 (.A(\div[15] ),
    .X(net121));
 sg13g2_dlygate4sd3_1 hold51 (.A(_065_),
    .X(net122));
 sg13g2_dlygate4sd3_1 hold52 (.A(\div[9] ),
    .X(net123));
 sg13g2_dlygate4sd3_1 hold53 (.A(\div[7] ),
    .X(net124));
 sg13g2_dlygate4sd3_1 hold54 (.A(_052_),
    .X(net125));
 sg13g2_dlygate4sd3_1 hold55 (.A(\div[12] ),
    .X(net126));
 sg13g2_dlygate4sd3_1 hold56 (.A(\div[13] ),
    .X(net127));
 sg13g2_dlygate4sd3_1 hold57 (.A(\div[20] ),
    .X(net128));
 sg13g2_dlygate4sd3_1 hold58 (.A(\lif1.timer[1] ),
    .X(net129));
 sg13g2_dlygate4sd3_1 hold59 (.A(\div[25] ),
    .X(net130));
 sg13g2_dlygate4sd3_1 hold60 (.A(\lif1.U[0] ),
    .X(net131));
 sg13g2_dlygate4sd3_1 hold61 (.A(\div[5] ),
    .X(net132));
 sg13g2_dlygate4sd3_1 hold62 (.A(\div[2] ),
    .X(net133));
 sg13g2_dlygate4sd3_1 hold63 (.A(_050_),
    .X(net134));
 sg13g2_dlygate4sd3_1 hold64 (.A(_005_),
    .X(net135));
 sg13g2_dlygate4sd3_1 hold65 (.A(\lif1.U[7] ),
    .X(net136));
 sg13g2_dlygate4sd3_1 hold66 (.A(\lif1.U[3] ),
    .X(net137));
 sg13g2_dlygate4sd3_1 hold67 (.A(\lif1.U[1] ),
    .X(net138));
 sg13g2_dlygate4sd3_1 hold68 (.A(\lif1.U[2] ),
    .X(net139));
 sg13g2_dlygate4sd3_1 hold69 (.A(\lif1.U[5] ),
    .X(net140));
 sg13g2_dlygate4sd3_1 hold70 (.A(\lif1.U[6] ),
    .X(net141));
 sg13g2_dlygate4sd3_1 hold71 (.A(\lif1.U[4] ),
    .X(net142));
 sg13g2_dlygate4sd3_1 hold72 (.A(\div[21] ),
    .X(net143));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_fill_2 FILLER_14_406 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_252 ();
 sg13g2_decap_8 FILLER_15_259 ();
 sg13g2_decap_8 FILLER_15_266 ();
 sg13g2_decap_8 FILLER_15_273 ();
 sg13g2_decap_8 FILLER_15_280 ();
 sg13g2_decap_8 FILLER_15_287 ();
 sg13g2_decap_8 FILLER_15_294 ();
 sg13g2_decap_8 FILLER_15_301 ();
 sg13g2_decap_8 FILLER_15_308 ();
 sg13g2_decap_8 FILLER_15_315 ();
 sg13g2_decap_8 FILLER_15_322 ();
 sg13g2_decap_8 FILLER_15_329 ();
 sg13g2_decap_8 FILLER_15_336 ();
 sg13g2_decap_8 FILLER_15_343 ();
 sg13g2_decap_8 FILLER_15_350 ();
 sg13g2_decap_8 FILLER_15_357 ();
 sg13g2_decap_8 FILLER_15_364 ();
 sg13g2_decap_8 FILLER_15_371 ();
 sg13g2_decap_8 FILLER_15_378 ();
 sg13g2_decap_8 FILLER_15_385 ();
 sg13g2_decap_8 FILLER_15_392 ();
 sg13g2_decap_8 FILLER_15_399 ();
 sg13g2_fill_2 FILLER_15_406 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_decap_8 FILLER_16_217 ();
 sg13g2_decap_8 FILLER_16_224 ();
 sg13g2_decap_8 FILLER_16_231 ();
 sg13g2_decap_8 FILLER_16_238 ();
 sg13g2_decap_8 FILLER_16_245 ();
 sg13g2_decap_8 FILLER_16_252 ();
 sg13g2_decap_8 FILLER_16_259 ();
 sg13g2_decap_8 FILLER_16_266 ();
 sg13g2_decap_8 FILLER_16_273 ();
 sg13g2_decap_8 FILLER_16_280 ();
 sg13g2_decap_8 FILLER_16_287 ();
 sg13g2_decap_8 FILLER_16_294 ();
 sg13g2_decap_8 FILLER_16_301 ();
 sg13g2_decap_8 FILLER_16_308 ();
 sg13g2_decap_8 FILLER_16_315 ();
 sg13g2_decap_8 FILLER_16_322 ();
 sg13g2_decap_8 FILLER_16_329 ();
 sg13g2_decap_8 FILLER_16_336 ();
 sg13g2_decap_8 FILLER_16_343 ();
 sg13g2_decap_8 FILLER_16_350 ();
 sg13g2_decap_8 FILLER_16_357 ();
 sg13g2_decap_8 FILLER_16_364 ();
 sg13g2_decap_8 FILLER_16_371 ();
 sg13g2_decap_8 FILLER_16_378 ();
 sg13g2_decap_8 FILLER_16_385 ();
 sg13g2_decap_8 FILLER_16_392 ();
 sg13g2_decap_8 FILLER_16_399 ();
 sg13g2_fill_2 FILLER_16_406 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_fill_1 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_163 ();
 sg13g2_decap_8 FILLER_17_170 ();
 sg13g2_decap_8 FILLER_17_177 ();
 sg13g2_decap_8 FILLER_17_184 ();
 sg13g2_decap_8 FILLER_17_191 ();
 sg13g2_decap_8 FILLER_17_198 ();
 sg13g2_decap_8 FILLER_17_205 ();
 sg13g2_decap_8 FILLER_17_212 ();
 sg13g2_decap_8 FILLER_17_219 ();
 sg13g2_fill_1 FILLER_17_226 ();
 sg13g2_decap_8 FILLER_17_231 ();
 sg13g2_decap_8 FILLER_17_238 ();
 sg13g2_decap_8 FILLER_17_245 ();
 sg13g2_decap_8 FILLER_17_252 ();
 sg13g2_decap_8 FILLER_17_259 ();
 sg13g2_decap_8 FILLER_17_266 ();
 sg13g2_decap_8 FILLER_17_273 ();
 sg13g2_decap_8 FILLER_17_280 ();
 sg13g2_decap_8 FILLER_17_287 ();
 sg13g2_decap_8 FILLER_17_294 ();
 sg13g2_decap_8 FILLER_17_301 ();
 sg13g2_decap_8 FILLER_17_308 ();
 sg13g2_decap_8 FILLER_17_315 ();
 sg13g2_decap_8 FILLER_17_322 ();
 sg13g2_decap_8 FILLER_17_329 ();
 sg13g2_decap_8 FILLER_17_336 ();
 sg13g2_decap_8 FILLER_17_343 ();
 sg13g2_decap_8 FILLER_17_350 ();
 sg13g2_decap_8 FILLER_17_357 ();
 sg13g2_decap_8 FILLER_17_364 ();
 sg13g2_decap_8 FILLER_17_371 ();
 sg13g2_decap_8 FILLER_17_378 ();
 sg13g2_decap_8 FILLER_17_385 ();
 sg13g2_decap_8 FILLER_17_392 ();
 sg13g2_decap_8 FILLER_17_399 ();
 sg13g2_fill_2 FILLER_17_406 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_fill_2 FILLER_18_147 ();
 sg13g2_fill_1 FILLER_18_149 ();
 sg13g2_decap_4 FILLER_18_159 ();
 sg13g2_fill_1 FILLER_18_172 ();
 sg13g2_decap_8 FILLER_18_199 ();
 sg13g2_fill_2 FILLER_18_206 ();
 sg13g2_fill_1 FILLER_18_208 ();
 sg13g2_fill_2 FILLER_18_226 ();
 sg13g2_decap_8 FILLER_18_237 ();
 sg13g2_decap_8 FILLER_18_244 ();
 sg13g2_decap_8 FILLER_18_251 ();
 sg13g2_decap_8 FILLER_18_258 ();
 sg13g2_decap_8 FILLER_18_265 ();
 sg13g2_decap_8 FILLER_18_272 ();
 sg13g2_decap_8 FILLER_18_279 ();
 sg13g2_decap_8 FILLER_18_286 ();
 sg13g2_decap_8 FILLER_18_293 ();
 sg13g2_decap_8 FILLER_18_300 ();
 sg13g2_decap_8 FILLER_18_307 ();
 sg13g2_decap_8 FILLER_18_314 ();
 sg13g2_decap_8 FILLER_18_321 ();
 sg13g2_decap_8 FILLER_18_328 ();
 sg13g2_decap_8 FILLER_18_335 ();
 sg13g2_decap_8 FILLER_18_342 ();
 sg13g2_decap_8 FILLER_18_349 ();
 sg13g2_decap_8 FILLER_18_356 ();
 sg13g2_decap_8 FILLER_18_363 ();
 sg13g2_decap_8 FILLER_18_370 ();
 sg13g2_decap_8 FILLER_18_377 ();
 sg13g2_decap_8 FILLER_18_384 ();
 sg13g2_decap_8 FILLER_18_391 ();
 sg13g2_decap_8 FILLER_18_398 ();
 sg13g2_decap_4 FILLER_18_405 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_decap_8 FILLER_19_166 ();
 sg13g2_fill_1 FILLER_19_182 ();
 sg13g2_fill_1 FILLER_19_187 ();
 sg13g2_decap_8 FILLER_19_247 ();
 sg13g2_decap_8 FILLER_19_254 ();
 sg13g2_decap_8 FILLER_19_261 ();
 sg13g2_decap_8 FILLER_19_268 ();
 sg13g2_decap_8 FILLER_19_275 ();
 sg13g2_decap_8 FILLER_19_282 ();
 sg13g2_decap_8 FILLER_19_289 ();
 sg13g2_decap_8 FILLER_19_296 ();
 sg13g2_decap_8 FILLER_19_303 ();
 sg13g2_decap_8 FILLER_19_310 ();
 sg13g2_decap_8 FILLER_19_317 ();
 sg13g2_decap_8 FILLER_19_324 ();
 sg13g2_decap_8 FILLER_19_331 ();
 sg13g2_decap_8 FILLER_19_338 ();
 sg13g2_decap_8 FILLER_19_345 ();
 sg13g2_decap_8 FILLER_19_352 ();
 sg13g2_decap_8 FILLER_19_359 ();
 sg13g2_decap_8 FILLER_19_366 ();
 sg13g2_decap_8 FILLER_19_373 ();
 sg13g2_decap_8 FILLER_19_380 ();
 sg13g2_decap_8 FILLER_19_387 ();
 sg13g2_decap_8 FILLER_19_394 ();
 sg13g2_decap_8 FILLER_19_401 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_decap_8 FILLER_20_126 ();
 sg13g2_decap_8 FILLER_20_133 ();
 sg13g2_decap_8 FILLER_20_140 ();
 sg13g2_decap_4 FILLER_20_147 ();
 sg13g2_fill_2 FILLER_20_155 ();
 sg13g2_fill_1 FILLER_20_157 ();
 sg13g2_fill_2 FILLER_20_180 ();
 sg13g2_fill_1 FILLER_20_182 ();
 sg13g2_fill_2 FILLER_20_223 ();
 sg13g2_fill_1 FILLER_20_225 ();
 sg13g2_decap_4 FILLER_20_252 ();
 sg13g2_decap_8 FILLER_20_264 ();
 sg13g2_decap_8 FILLER_20_271 ();
 sg13g2_decap_8 FILLER_20_278 ();
 sg13g2_decap_8 FILLER_20_285 ();
 sg13g2_decap_8 FILLER_20_292 ();
 sg13g2_decap_8 FILLER_20_299 ();
 sg13g2_decap_8 FILLER_20_306 ();
 sg13g2_decap_8 FILLER_20_313 ();
 sg13g2_decap_8 FILLER_20_320 ();
 sg13g2_decap_8 FILLER_20_327 ();
 sg13g2_decap_8 FILLER_20_334 ();
 sg13g2_decap_8 FILLER_20_341 ();
 sg13g2_decap_8 FILLER_20_348 ();
 sg13g2_decap_8 FILLER_20_355 ();
 sg13g2_decap_8 FILLER_20_362 ();
 sg13g2_decap_8 FILLER_20_369 ();
 sg13g2_decap_8 FILLER_20_376 ();
 sg13g2_decap_8 FILLER_20_383 ();
 sg13g2_decap_8 FILLER_20_390 ();
 sg13g2_decap_8 FILLER_20_397 ();
 sg13g2_decap_4 FILLER_20_404 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_decap_8 FILLER_21_119 ();
 sg13g2_decap_8 FILLER_21_126 ();
 sg13g2_fill_2 FILLER_21_133 ();
 sg13g2_fill_1 FILLER_21_135 ();
 sg13g2_fill_1 FILLER_21_162 ();
 sg13g2_fill_2 FILLER_21_197 ();
 sg13g2_fill_1 FILLER_21_217 ();
 sg13g2_fill_1 FILLER_21_240 ();
 sg13g2_fill_1 FILLER_21_250 ();
 sg13g2_decap_8 FILLER_21_277 ();
 sg13g2_decap_8 FILLER_21_284 ();
 sg13g2_decap_8 FILLER_21_291 ();
 sg13g2_decap_8 FILLER_21_298 ();
 sg13g2_decap_8 FILLER_21_305 ();
 sg13g2_decap_8 FILLER_21_312 ();
 sg13g2_decap_8 FILLER_21_319 ();
 sg13g2_decap_8 FILLER_21_326 ();
 sg13g2_decap_8 FILLER_21_333 ();
 sg13g2_decap_8 FILLER_21_340 ();
 sg13g2_decap_8 FILLER_21_347 ();
 sg13g2_decap_8 FILLER_21_354 ();
 sg13g2_decap_8 FILLER_21_361 ();
 sg13g2_decap_8 FILLER_21_368 ();
 sg13g2_decap_8 FILLER_21_375 ();
 sg13g2_decap_8 FILLER_21_382 ();
 sg13g2_decap_8 FILLER_21_389 ();
 sg13g2_decap_8 FILLER_21_396 ();
 sg13g2_decap_4 FILLER_21_403 ();
 sg13g2_fill_2 FILLER_21_407 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_8 FILLER_22_105 ();
 sg13g2_decap_8 FILLER_22_112 ();
 sg13g2_decap_8 FILLER_22_119 ();
 sg13g2_decap_8 FILLER_22_126 ();
 sg13g2_decap_8 FILLER_22_133 ();
 sg13g2_fill_2 FILLER_22_180 ();
 sg13g2_fill_2 FILLER_22_221 ();
 sg13g2_decap_8 FILLER_22_297 ();
 sg13g2_decap_8 FILLER_22_304 ();
 sg13g2_decap_8 FILLER_22_311 ();
 sg13g2_decap_8 FILLER_22_318 ();
 sg13g2_decap_8 FILLER_22_325 ();
 sg13g2_decap_8 FILLER_22_332 ();
 sg13g2_decap_8 FILLER_22_339 ();
 sg13g2_decap_8 FILLER_22_346 ();
 sg13g2_decap_8 FILLER_22_353 ();
 sg13g2_decap_8 FILLER_22_360 ();
 sg13g2_decap_8 FILLER_22_367 ();
 sg13g2_decap_8 FILLER_22_374 ();
 sg13g2_decap_8 FILLER_22_381 ();
 sg13g2_decap_8 FILLER_22_388 ();
 sg13g2_decap_8 FILLER_22_395 ();
 sg13g2_decap_8 FILLER_22_402 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_98 ();
 sg13g2_decap_8 FILLER_23_105 ();
 sg13g2_decap_8 FILLER_23_112 ();
 sg13g2_decap_8 FILLER_23_119 ();
 sg13g2_decap_8 FILLER_23_126 ();
 sg13g2_decap_8 FILLER_23_133 ();
 sg13g2_decap_4 FILLER_23_140 ();
 sg13g2_fill_1 FILLER_23_144 ();
 sg13g2_fill_2 FILLER_23_182 ();
 sg13g2_fill_1 FILLER_23_184 ();
 sg13g2_fill_2 FILLER_23_211 ();
 sg13g2_fill_1 FILLER_23_223 ();
 sg13g2_fill_1 FILLER_23_232 ();
 sg13g2_decap_4 FILLER_23_251 ();
 sg13g2_decap_8 FILLER_23_294 ();
 sg13g2_decap_8 FILLER_23_301 ();
 sg13g2_decap_8 FILLER_23_308 ();
 sg13g2_decap_8 FILLER_23_315 ();
 sg13g2_decap_8 FILLER_23_322 ();
 sg13g2_decap_8 FILLER_23_329 ();
 sg13g2_decap_8 FILLER_23_336 ();
 sg13g2_decap_8 FILLER_23_343 ();
 sg13g2_decap_8 FILLER_23_350 ();
 sg13g2_decap_8 FILLER_23_357 ();
 sg13g2_decap_8 FILLER_23_364 ();
 sg13g2_decap_8 FILLER_23_371 ();
 sg13g2_decap_8 FILLER_23_378 ();
 sg13g2_decap_8 FILLER_23_385 ();
 sg13g2_decap_8 FILLER_23_392 ();
 sg13g2_decap_8 FILLER_23_399 ();
 sg13g2_fill_2 FILLER_23_406 ();
 sg13g2_fill_1 FILLER_23_408 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_decap_8 FILLER_24_98 ();
 sg13g2_decap_8 FILLER_24_105 ();
 sg13g2_decap_8 FILLER_24_112 ();
 sg13g2_decap_8 FILLER_24_119 ();
 sg13g2_decap_8 FILLER_24_126 ();
 sg13g2_decap_8 FILLER_24_133 ();
 sg13g2_decap_8 FILLER_24_140 ();
 sg13g2_decap_4 FILLER_24_147 ();
 sg13g2_fill_1 FILLER_24_160 ();
 sg13g2_fill_2 FILLER_24_174 ();
 sg13g2_fill_2 FILLER_24_220 ();
 sg13g2_fill_1 FILLER_24_222 ();
 sg13g2_fill_2 FILLER_24_242 ();
 sg13g2_fill_1 FILLER_24_244 ();
 sg13g2_decap_8 FILLER_24_282 ();
 sg13g2_decap_8 FILLER_24_289 ();
 sg13g2_decap_8 FILLER_24_296 ();
 sg13g2_decap_8 FILLER_24_303 ();
 sg13g2_decap_8 FILLER_24_310 ();
 sg13g2_decap_8 FILLER_24_317 ();
 sg13g2_decap_8 FILLER_24_324 ();
 sg13g2_decap_8 FILLER_24_331 ();
 sg13g2_decap_8 FILLER_24_338 ();
 sg13g2_decap_8 FILLER_24_345 ();
 sg13g2_decap_8 FILLER_24_352 ();
 sg13g2_decap_8 FILLER_24_359 ();
 sg13g2_decap_8 FILLER_24_366 ();
 sg13g2_decap_8 FILLER_24_373 ();
 sg13g2_decap_8 FILLER_24_380 ();
 sg13g2_decap_8 FILLER_24_387 ();
 sg13g2_decap_8 FILLER_24_394 ();
 sg13g2_decap_8 FILLER_24_401 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_8 FILLER_25_91 ();
 sg13g2_decap_8 FILLER_25_98 ();
 sg13g2_decap_8 FILLER_25_105 ();
 sg13g2_decap_8 FILLER_25_112 ();
 sg13g2_decap_8 FILLER_25_119 ();
 sg13g2_decap_8 FILLER_25_126 ();
 sg13g2_decap_8 FILLER_25_133 ();
 sg13g2_fill_2 FILLER_25_140 ();
 sg13g2_fill_1 FILLER_25_142 ();
 sg13g2_fill_2 FILLER_25_192 ();
 sg13g2_fill_1 FILLER_25_194 ();
 sg13g2_fill_2 FILLER_25_199 ();
 sg13g2_fill_2 FILLER_25_210 ();
 sg13g2_fill_1 FILLER_25_212 ();
 sg13g2_fill_1 FILLER_25_227 ();
 sg13g2_decap_4 FILLER_25_278 ();
 sg13g2_decap_8 FILLER_25_287 ();
 sg13g2_decap_8 FILLER_25_294 ();
 sg13g2_decap_8 FILLER_25_305 ();
 sg13g2_decap_8 FILLER_25_312 ();
 sg13g2_decap_8 FILLER_25_319 ();
 sg13g2_decap_8 FILLER_25_326 ();
 sg13g2_decap_8 FILLER_25_333 ();
 sg13g2_decap_8 FILLER_25_340 ();
 sg13g2_decap_8 FILLER_25_347 ();
 sg13g2_decap_8 FILLER_25_354 ();
 sg13g2_decap_8 FILLER_25_361 ();
 sg13g2_decap_8 FILLER_25_368 ();
 sg13g2_decap_8 FILLER_25_375 ();
 sg13g2_decap_8 FILLER_25_382 ();
 sg13g2_decap_8 FILLER_25_389 ();
 sg13g2_decap_8 FILLER_25_396 ();
 sg13g2_decap_4 FILLER_25_403 ();
 sg13g2_fill_2 FILLER_25_407 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_decap_8 FILLER_26_91 ();
 sg13g2_decap_8 FILLER_26_98 ();
 sg13g2_decap_8 FILLER_26_105 ();
 sg13g2_decap_8 FILLER_26_112 ();
 sg13g2_decap_8 FILLER_26_119 ();
 sg13g2_decap_8 FILLER_26_126 ();
 sg13g2_decap_4 FILLER_26_133 ();
 sg13g2_fill_2 FILLER_26_137 ();
 sg13g2_fill_2 FILLER_26_165 ();
 sg13g2_fill_1 FILLER_26_167 ();
 sg13g2_fill_2 FILLER_26_177 ();
 sg13g2_fill_1 FILLER_26_188 ();
 sg13g2_decap_4 FILLER_26_284 ();
 sg13g2_fill_2 FILLER_26_288 ();
 sg13g2_fill_2 FILLER_26_301 ();
 sg13g2_fill_1 FILLER_26_303 ();
 sg13g2_decap_4 FILLER_26_313 ();
 sg13g2_fill_1 FILLER_26_317 ();
 sg13g2_decap_8 FILLER_26_323 ();
 sg13g2_decap_8 FILLER_26_330 ();
 sg13g2_decap_8 FILLER_26_337 ();
 sg13g2_decap_8 FILLER_26_344 ();
 sg13g2_decap_8 FILLER_26_351 ();
 sg13g2_decap_8 FILLER_26_358 ();
 sg13g2_decap_8 FILLER_26_365 ();
 sg13g2_decap_8 FILLER_26_372 ();
 sg13g2_decap_8 FILLER_26_379 ();
 sg13g2_decap_8 FILLER_26_386 ();
 sg13g2_decap_8 FILLER_26_393 ();
 sg13g2_decap_8 FILLER_26_400 ();
 sg13g2_fill_2 FILLER_26_407 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_decap_8 FILLER_27_84 ();
 sg13g2_decap_8 FILLER_27_91 ();
 sg13g2_decap_8 FILLER_27_98 ();
 sg13g2_decap_8 FILLER_27_105 ();
 sg13g2_decap_8 FILLER_27_112 ();
 sg13g2_decap_8 FILLER_27_119 ();
 sg13g2_decap_8 FILLER_27_126 ();
 sg13g2_fill_2 FILLER_27_133 ();
 sg13g2_fill_2 FILLER_27_170 ();
 sg13g2_fill_2 FILLER_27_194 ();
 sg13g2_fill_2 FILLER_27_214 ();
 sg13g2_fill_2 FILLER_27_230 ();
 sg13g2_fill_1 FILLER_27_232 ();
 sg13g2_fill_1 FILLER_27_261 ();
 sg13g2_fill_2 FILLER_27_288 ();
 sg13g2_fill_2 FILLER_27_316 ();
 sg13g2_decap_8 FILLER_27_349 ();
 sg13g2_decap_8 FILLER_27_356 ();
 sg13g2_decap_8 FILLER_27_363 ();
 sg13g2_decap_8 FILLER_27_370 ();
 sg13g2_decap_8 FILLER_27_377 ();
 sg13g2_decap_8 FILLER_27_384 ();
 sg13g2_decap_8 FILLER_27_391 ();
 sg13g2_decap_8 FILLER_27_398 ();
 sg13g2_decap_4 FILLER_27_405 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_decap_8 FILLER_28_84 ();
 sg13g2_decap_8 FILLER_28_91 ();
 sg13g2_decap_8 FILLER_28_98 ();
 sg13g2_decap_8 FILLER_28_105 ();
 sg13g2_decap_8 FILLER_28_112 ();
 sg13g2_decap_8 FILLER_28_119 ();
 sg13g2_decap_8 FILLER_28_126 ();
 sg13g2_fill_1 FILLER_28_133 ();
 sg13g2_fill_1 FILLER_28_243 ();
 sg13g2_fill_1 FILLER_28_293 ();
 sg13g2_decap_8 FILLER_28_353 ();
 sg13g2_decap_8 FILLER_28_360 ();
 sg13g2_decap_8 FILLER_28_367 ();
 sg13g2_decap_8 FILLER_28_374 ();
 sg13g2_decap_8 FILLER_28_381 ();
 sg13g2_decap_8 FILLER_28_388 ();
 sg13g2_decap_8 FILLER_28_395 ();
 sg13g2_decap_8 FILLER_28_402 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_decap_8 FILLER_29_84 ();
 sg13g2_decap_8 FILLER_29_91 ();
 sg13g2_decap_8 FILLER_29_98 ();
 sg13g2_decap_8 FILLER_29_105 ();
 sg13g2_decap_8 FILLER_29_112 ();
 sg13g2_decap_8 FILLER_29_119 ();
 sg13g2_decap_8 FILLER_29_126 ();
 sg13g2_decap_4 FILLER_29_133 ();
 sg13g2_fill_2 FILLER_29_137 ();
 sg13g2_fill_2 FILLER_29_183 ();
 sg13g2_fill_1 FILLER_29_185 ();
 sg13g2_fill_1 FILLER_29_212 ();
 sg13g2_fill_2 FILLER_29_242 ();
 sg13g2_fill_1 FILLER_29_244 ();
 sg13g2_fill_2 FILLER_29_275 ();
 sg13g2_fill_1 FILLER_29_283 ();
 sg13g2_fill_1 FILLER_29_329 ();
 sg13g2_decap_4 FILLER_29_356 ();
 sg13g2_decap_8 FILLER_29_386 ();
 sg13g2_decap_8 FILLER_29_393 ();
 sg13g2_decap_8 FILLER_29_400 ();
 sg13g2_fill_2 FILLER_29_407 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_77 ();
 sg13g2_decap_8 FILLER_30_84 ();
 sg13g2_decap_8 FILLER_30_91 ();
 sg13g2_decap_8 FILLER_30_98 ();
 sg13g2_decap_8 FILLER_30_105 ();
 sg13g2_decap_8 FILLER_30_112 ();
 sg13g2_decap_8 FILLER_30_119 ();
 sg13g2_decap_8 FILLER_30_126 ();
 sg13g2_decap_8 FILLER_30_133 ();
 sg13g2_decap_4 FILLER_30_140 ();
 sg13g2_fill_1 FILLER_30_144 ();
 sg13g2_fill_1 FILLER_30_167 ();
 sg13g2_fill_1 FILLER_30_180 ();
 sg13g2_decap_4 FILLER_30_225 ();
 sg13g2_fill_2 FILLER_30_264 ();
 sg13g2_fill_2 FILLER_30_281 ();
 sg13g2_fill_1 FILLER_30_305 ();
 sg13g2_fill_2 FILLER_30_315 ();
 sg13g2_fill_1 FILLER_30_327 ();
 sg13g2_decap_4 FILLER_30_350 ();
 sg13g2_fill_2 FILLER_30_354 ();
 sg13g2_fill_2 FILLER_30_359 ();
 sg13g2_fill_1 FILLER_30_361 ();
 sg13g2_decap_4 FILLER_30_390 ();
 sg13g2_decap_8 FILLER_30_398 ();
 sg13g2_decap_4 FILLER_30_405 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_decap_8 FILLER_31_84 ();
 sg13g2_decap_8 FILLER_31_91 ();
 sg13g2_decap_8 FILLER_31_98 ();
 sg13g2_decap_8 FILLER_31_105 ();
 sg13g2_decap_8 FILLER_31_112 ();
 sg13g2_decap_8 FILLER_31_119 ();
 sg13g2_decap_8 FILLER_31_126 ();
 sg13g2_decap_8 FILLER_31_133 ();
 sg13g2_decap_8 FILLER_31_140 ();
 sg13g2_fill_2 FILLER_31_147 ();
 sg13g2_fill_1 FILLER_31_149 ();
 sg13g2_fill_2 FILLER_31_191 ();
 sg13g2_fill_1 FILLER_31_193 ();
 sg13g2_decap_8 FILLER_31_203 ();
 sg13g2_decap_4 FILLER_31_210 ();
 sg13g2_fill_1 FILLER_31_269 ();
 sg13g2_fill_2 FILLER_31_274 ();
 sg13g2_fill_2 FILLER_31_318 ();
 sg13g2_fill_1 FILLER_31_320 ();
 sg13g2_fill_2 FILLER_31_327 ();
 sg13g2_fill_1 FILLER_31_329 ();
 sg13g2_fill_1 FILLER_31_370 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_8 FILLER_32_84 ();
 sg13g2_decap_8 FILLER_32_91 ();
 sg13g2_decap_8 FILLER_32_98 ();
 sg13g2_decap_8 FILLER_32_105 ();
 sg13g2_decap_8 FILLER_32_112 ();
 sg13g2_decap_8 FILLER_32_119 ();
 sg13g2_decap_8 FILLER_32_126 ();
 sg13g2_decap_8 FILLER_32_133 ();
 sg13g2_decap_8 FILLER_32_140 ();
 sg13g2_decap_8 FILLER_32_147 ();
 sg13g2_decap_4 FILLER_32_154 ();
 sg13g2_fill_1 FILLER_32_158 ();
 sg13g2_decap_8 FILLER_32_189 ();
 sg13g2_decap_8 FILLER_32_196 ();
 sg13g2_decap_8 FILLER_32_203 ();
 sg13g2_decap_4 FILLER_32_210 ();
 sg13g2_fill_1 FILLER_32_214 ();
 sg13g2_decap_4 FILLER_32_233 ();
 sg13g2_fill_2 FILLER_32_237 ();
 sg13g2_fill_1 FILLER_32_274 ();
 sg13g2_decap_4 FILLER_32_328 ();
 sg13g2_fill_1 FILLER_32_347 ();
 sg13g2_decap_4 FILLER_32_366 ();
 sg13g2_fill_2 FILLER_32_370 ();
 sg13g2_fill_2 FILLER_32_377 ();
 sg13g2_decap_4 FILLER_32_384 ();
 sg13g2_fill_2 FILLER_32_388 ();
 sg13g2_decap_4 FILLER_32_403 ();
 sg13g2_fill_2 FILLER_32_407 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_decap_8 FILLER_33_91 ();
 sg13g2_decap_8 FILLER_33_98 ();
 sg13g2_decap_8 FILLER_33_105 ();
 sg13g2_decap_8 FILLER_33_112 ();
 sg13g2_decap_8 FILLER_33_119 ();
 sg13g2_decap_8 FILLER_33_126 ();
 sg13g2_decap_8 FILLER_33_133 ();
 sg13g2_decap_8 FILLER_33_140 ();
 sg13g2_decap_8 FILLER_33_147 ();
 sg13g2_decap_8 FILLER_33_154 ();
 sg13g2_decap_8 FILLER_33_161 ();
 sg13g2_decap_4 FILLER_33_168 ();
 sg13g2_fill_2 FILLER_33_172 ();
 sg13g2_decap_8 FILLER_33_178 ();
 sg13g2_decap_8 FILLER_33_185 ();
 sg13g2_decap_8 FILLER_33_192 ();
 sg13g2_decap_8 FILLER_33_199 ();
 sg13g2_decap_8 FILLER_33_206 ();
 sg13g2_decap_8 FILLER_33_213 ();
 sg13g2_decap_8 FILLER_33_220 ();
 sg13g2_decap_8 FILLER_33_227 ();
 sg13g2_decap_8 FILLER_33_234 ();
 sg13g2_decap_8 FILLER_33_241 ();
 sg13g2_fill_2 FILLER_33_248 ();
 sg13g2_fill_1 FILLER_33_254 ();
 sg13g2_fill_1 FILLER_33_279 ();
 sg13g2_fill_2 FILLER_33_298 ();
 sg13g2_fill_1 FILLER_33_322 ();
 sg13g2_fill_1 FILLER_33_338 ();
 sg13g2_fill_1 FILLER_33_376 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_decap_8 FILLER_34_91 ();
 sg13g2_decap_8 FILLER_34_98 ();
 sg13g2_decap_8 FILLER_34_105 ();
 sg13g2_decap_8 FILLER_34_112 ();
 sg13g2_decap_8 FILLER_34_119 ();
 sg13g2_decap_8 FILLER_34_126 ();
 sg13g2_decap_8 FILLER_34_133 ();
 sg13g2_decap_8 FILLER_34_140 ();
 sg13g2_decap_8 FILLER_34_147 ();
 sg13g2_decap_8 FILLER_34_154 ();
 sg13g2_decap_8 FILLER_34_161 ();
 sg13g2_decap_8 FILLER_34_168 ();
 sg13g2_decap_8 FILLER_34_175 ();
 sg13g2_decap_8 FILLER_34_182 ();
 sg13g2_decap_8 FILLER_34_189 ();
 sg13g2_decap_8 FILLER_34_196 ();
 sg13g2_decap_8 FILLER_34_203 ();
 sg13g2_decap_8 FILLER_34_210 ();
 sg13g2_decap_8 FILLER_34_217 ();
 sg13g2_decap_8 FILLER_34_224 ();
 sg13g2_decap_8 FILLER_34_231 ();
 sg13g2_decap_8 FILLER_34_238 ();
 sg13g2_decap_8 FILLER_34_245 ();
 sg13g2_fill_2 FILLER_34_277 ();
 sg13g2_fill_1 FILLER_34_279 ();
 sg13g2_decap_4 FILLER_34_297 ();
 sg13g2_fill_2 FILLER_34_301 ();
 sg13g2_decap_8 FILLER_34_319 ();
 sg13g2_decap_8 FILLER_34_326 ();
 sg13g2_decap_8 FILLER_34_333 ();
 sg13g2_decap_4 FILLER_34_350 ();
 sg13g2_fill_2 FILLER_34_354 ();
 sg13g2_fill_2 FILLER_34_365 ();
 sg13g2_fill_1 FILLER_34_376 ();
 sg13g2_fill_2 FILLER_34_382 ();
 sg13g2_fill_1 FILLER_34_408 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_decap_8 FILLER_35_98 ();
 sg13g2_decap_8 FILLER_35_105 ();
 sg13g2_decap_8 FILLER_35_112 ();
 sg13g2_decap_8 FILLER_35_119 ();
 sg13g2_decap_8 FILLER_35_126 ();
 sg13g2_decap_8 FILLER_35_133 ();
 sg13g2_decap_8 FILLER_35_140 ();
 sg13g2_decap_8 FILLER_35_147 ();
 sg13g2_decap_8 FILLER_35_154 ();
 sg13g2_decap_8 FILLER_35_161 ();
 sg13g2_decap_8 FILLER_35_168 ();
 sg13g2_decap_8 FILLER_35_175 ();
 sg13g2_decap_8 FILLER_35_182 ();
 sg13g2_decap_8 FILLER_35_189 ();
 sg13g2_decap_8 FILLER_35_196 ();
 sg13g2_decap_8 FILLER_35_203 ();
 sg13g2_decap_8 FILLER_35_210 ();
 sg13g2_decap_8 FILLER_35_217 ();
 sg13g2_decap_8 FILLER_35_224 ();
 sg13g2_decap_8 FILLER_35_231 ();
 sg13g2_decap_8 FILLER_35_238 ();
 sg13g2_decap_8 FILLER_35_245 ();
 sg13g2_decap_8 FILLER_35_252 ();
 sg13g2_fill_2 FILLER_35_259 ();
 sg13g2_decap_4 FILLER_35_279 ();
 sg13g2_decap_8 FILLER_35_295 ();
 sg13g2_decap_4 FILLER_35_302 ();
 sg13g2_fill_2 FILLER_35_306 ();
 sg13g2_decap_4 FILLER_35_316 ();
 sg13g2_fill_2 FILLER_35_336 ();
 sg13g2_fill_1 FILLER_35_338 ();
 sg13g2_decap_8 FILLER_35_359 ();
 sg13g2_fill_2 FILLER_35_366 ();
 sg13g2_fill_1 FILLER_35_381 ();
 sg13g2_fill_2 FILLER_35_387 ();
 sg13g2_decap_4 FILLER_35_405 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_decap_8 FILLER_36_112 ();
 sg13g2_decap_8 FILLER_36_119 ();
 sg13g2_decap_8 FILLER_36_126 ();
 sg13g2_decap_8 FILLER_36_133 ();
 sg13g2_decap_8 FILLER_36_140 ();
 sg13g2_decap_8 FILLER_36_147 ();
 sg13g2_decap_8 FILLER_36_154 ();
 sg13g2_decap_8 FILLER_36_161 ();
 sg13g2_decap_8 FILLER_36_168 ();
 sg13g2_decap_8 FILLER_36_175 ();
 sg13g2_decap_8 FILLER_36_182 ();
 sg13g2_decap_8 FILLER_36_189 ();
 sg13g2_decap_8 FILLER_36_196 ();
 sg13g2_decap_8 FILLER_36_203 ();
 sg13g2_decap_8 FILLER_36_210 ();
 sg13g2_decap_8 FILLER_36_217 ();
 sg13g2_decap_8 FILLER_36_224 ();
 sg13g2_decap_8 FILLER_36_231 ();
 sg13g2_decap_8 FILLER_36_238 ();
 sg13g2_decap_8 FILLER_36_245 ();
 sg13g2_decap_8 FILLER_36_252 ();
 sg13g2_decap_4 FILLER_36_259 ();
 sg13g2_fill_2 FILLER_36_263 ();
 sg13g2_fill_2 FILLER_36_269 ();
 sg13g2_fill_2 FILLER_36_326 ();
 sg13g2_decap_4 FILLER_36_334 ();
 sg13g2_fill_2 FILLER_36_338 ();
 sg13g2_fill_2 FILLER_36_358 ();
 sg13g2_fill_1 FILLER_36_360 ();
 sg13g2_fill_2 FILLER_36_380 ();
 sg13g2_fill_1 FILLER_36_408 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_8 FILLER_37_112 ();
 sg13g2_decap_8 FILLER_37_119 ();
 sg13g2_decap_8 FILLER_37_126 ();
 sg13g2_decap_8 FILLER_37_133 ();
 sg13g2_decap_8 FILLER_37_140 ();
 sg13g2_decap_8 FILLER_37_147 ();
 sg13g2_decap_8 FILLER_37_154 ();
 sg13g2_decap_8 FILLER_37_161 ();
 sg13g2_decap_8 FILLER_37_168 ();
 sg13g2_decap_8 FILLER_37_175 ();
 sg13g2_decap_8 FILLER_37_182 ();
 sg13g2_decap_8 FILLER_37_189 ();
 sg13g2_decap_8 FILLER_37_196 ();
 sg13g2_decap_8 FILLER_37_203 ();
 sg13g2_decap_8 FILLER_37_210 ();
 sg13g2_decap_8 FILLER_37_217 ();
 sg13g2_decap_8 FILLER_37_224 ();
 sg13g2_decap_8 FILLER_37_231 ();
 sg13g2_decap_8 FILLER_37_238 ();
 sg13g2_decap_8 FILLER_37_245 ();
 sg13g2_decap_8 FILLER_37_252 ();
 sg13g2_decap_8 FILLER_37_259 ();
 sg13g2_decap_8 FILLER_37_266 ();
 sg13g2_decap_8 FILLER_37_273 ();
 sg13g2_decap_8 FILLER_37_280 ();
 sg13g2_decap_8 FILLER_37_287 ();
 sg13g2_fill_2 FILLER_37_307 ();
 sg13g2_fill_1 FILLER_37_309 ();
 sg13g2_fill_1 FILLER_37_366 ();
 sg13g2_fill_2 FILLER_37_380 ();
 sg13g2_fill_1 FILLER_37_408 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_4 FILLER_38_60 ();
 sg13g2_decap_4 FILLER_38_68 ();
 sg13g2_decap_4 FILLER_38_76 ();
 sg13g2_decap_4 FILLER_38_84 ();
 sg13g2_decap_4 FILLER_38_92 ();
 sg13g2_decap_4 FILLER_38_100 ();
 sg13g2_decap_4 FILLER_38_108 ();
 sg13g2_decap_4 FILLER_38_116 ();
 sg13g2_decap_4 FILLER_38_124 ();
 sg13g2_decap_4 FILLER_38_132 ();
 sg13g2_decap_4 FILLER_38_140 ();
 sg13g2_decap_4 FILLER_38_148 ();
 sg13g2_decap_4 FILLER_38_156 ();
 sg13g2_decap_4 FILLER_38_164 ();
 sg13g2_decap_4 FILLER_38_172 ();
 sg13g2_decap_8 FILLER_38_180 ();
 sg13g2_decap_8 FILLER_38_187 ();
 sg13g2_decap_8 FILLER_38_194 ();
 sg13g2_decap_8 FILLER_38_201 ();
 sg13g2_decap_8 FILLER_38_208 ();
 sg13g2_decap_8 FILLER_38_215 ();
 sg13g2_decap_8 FILLER_38_222 ();
 sg13g2_decap_8 FILLER_38_229 ();
 sg13g2_decap_8 FILLER_38_236 ();
 sg13g2_decap_8 FILLER_38_243 ();
 sg13g2_decap_8 FILLER_38_250 ();
 sg13g2_decap_8 FILLER_38_257 ();
 sg13g2_decap_8 FILLER_38_264 ();
 sg13g2_decap_8 FILLER_38_271 ();
 sg13g2_decap_8 FILLER_38_278 ();
 sg13g2_decap_8 FILLER_38_285 ();
 sg13g2_decap_8 FILLER_38_292 ();
 sg13g2_fill_1 FILLER_38_299 ();
 sg13g2_fill_2 FILLER_38_341 ();
 sg13g2_fill_1 FILLER_38_343 ();
 sg13g2_fill_2 FILLER_38_353 ();
 sg13g2_fill_1 FILLER_38_355 ();
 sg13g2_fill_2 FILLER_38_387 ();
 sg13g2_decap_8 FILLER_38_401 ();
 sg13g2_fill_1 FILLER_38_408 ();
 assign uio_oe[0] = net10;
 assign uio_oe[1] = net11;
 assign uio_oe[2] = net12;
 assign uio_oe[3] = net13;
 assign uio_oe[4] = net14;
 assign uio_oe[5] = net15;
 assign uio_oe[6] = net16;
 assign uio_oe[7] = net17;
 assign uio_out[0] = net18;
 assign uio_out[1] = net19;
 assign uio_out[2] = net20;
 assign uio_out[3] = net21;
 assign uio_out[4] = net22;
 assign uio_out[5] = net23;
 assign uio_out[6] = net24;
 assign uio_out[7] = net25;
endmodule

module tt_um_ran_DanielZhu (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire inverterringout;
 wire ran16out;
 wire ranbitstring;
 wire \tt_16bitran.connection[10] ;
 wire \tt_16bitran.connection[11] ;
 wire \tt_16bitran.connection[12] ;
 wire \tt_16bitran.connection[13] ;
 wire \tt_16bitran.connection[14] ;
 wire \tt_16bitran.connection[15] ;
 wire \tt_16bitran.connection[1] ;
 wire \tt_16bitran.connection[2] ;
 wire \tt_16bitran.connection[3] ;
 wire \tt_16bitran.connection[4] ;
 wire \tt_16bitran.connection[5] ;
 wire \tt_16bitran.connection[6] ;
 wire \tt_16bitran.connection[7] ;
 wire \tt_16bitran.connection[8] ;
 wire \tt_16bitran.connection[9] ;
 wire \tt_finalprocess.genblk1[0].multblock.multblockout ;
 wire \tt_finalprocess.genblk1[1].multblock.multblockout ;
 wire \tt_finalprocess.genblk1[2].multblock.multblockout ;
 wire \tt_finalprocess.genblk1[3].multblock.multblockout ;
 wire \tt_finalprocess.genblk1[4].multblock.multblockout ;
 wire \tt_finalprocess.genblk1[5].multblock.multblockout ;
 wire \tt_finalprocess.genblk1[6].multblock.multblockout ;
 wire \tt_finalprocess.genblk1[7].multblock.multblockout ;
 wire \tt_finalprocess.num2[0] ;
 wire \tt_finalprocess.num2[1] ;
 wire \tt_finalprocess.num2[2] ;
 wire \tt_finalprocess.num2[3] ;
 wire \tt_invring1.ringosc1[10].inv.cnt_bit_I.Y ;
 wire \tt_invring1.ringosc2[18].inv.cnt_bit_I.Y ;
 wire \tt_invring1.ringosc3[22].inv.cnt_bit_I.Y ;
 wire \tt_invring1.ringosc4[28].inv.cnt_bit_I.Y ;
 wire \tt_invring1.ringosc5[36].inv.cnt_bit_I.Y ;
 wire \tt_invring1.ringosc6[40].inv.cnt_bit_I.Y ;
 wire \tt_invring1.ringosc7[46].inv.cnt_bit_I.Y ;
 wire \tt_invring1.ringosc8[38].inv.cnt_bit_I.Y ;
 wire \tt_invring1.ringoutsam[0] ;
 wire \tt_invring1.ringoutsam[1] ;
 wire \tt_invring1.ringoutsam[2] ;
 wire \tt_invring1.ringoutsam[3] ;
 wire \tt_invring1.ringoutsam[4] ;
 wire \tt_invring1.ringoutsam[5] ;
 wire \tt_invring1.ringoutsam[6] ;
 wire \tt_invring1.ringoutsam[7] ;
 wire \tt_invring2.ringosc1[10].inv.cnt_bit_I.Y ;
 wire \tt_invring2.ringosc2[18].inv.cnt_bit_I.Y ;
 wire \tt_invring2.ringosc3[22].inv.cnt_bit_I.Y ;
 wire \tt_invring2.ringosc4[28].inv.cnt_bit_I.Y ;
 wire \tt_invring2.ringosc5[36].inv.cnt_bit_I.Y ;
 wire \tt_invring2.ringosc6[40].inv.cnt_bit_I.Y ;
 wire \tt_invring2.ringosc7[46].inv.cnt_bit_I.Y ;
 wire \tt_invring2.ringosc8[38].inv.cnt_bit_I.Y ;
 wire \tt_invring2.ringoutsam[0] ;
 wire \tt_invring2.ringoutsam[1] ;
 wire \tt_invring2.ringoutsam[2] ;
 wire \tt_invring2.ringoutsam[3] ;
 wire \tt_invring2.ringoutsam[4] ;
 wire \tt_invring2.ringoutsam[5] ;
 wire \tt_invring2.ringoutsam[6] ;
 wire \tt_invring2.ringoutsam[7] ;
 wire \tt_process.bitsadjacent[0] ;
 wire \tt_process.bitsadjacent[1] ;
 wire \tt_process.bitsadjacent[2] ;
 wire \tt_process.bitsgroup[0] ;
 wire \tt_process.bitsgroup[1] ;
 wire \tt_process.clk_half ;
 wire \tt_process.tt_13n.connection[0] ;
 wire \tt_process.tt_13n.connection[10] ;
 wire \tt_process.tt_13n.connection[11] ;
 wire \tt_process.tt_13n.connection[12] ;
 wire \tt_process.tt_13n.connection[13] ;
 wire \tt_process.tt_13n.connection[1] ;
 wire \tt_process.tt_13n.connection[2] ;
 wire \tt_process.tt_13n.connection[3] ;
 wire \tt_process.tt_13n.connection[4] ;
 wire \tt_process.tt_13n.connection[5] ;
 wire \tt_process.tt_13n.connection[6] ;
 wire \tt_process.tt_13n.connection[7] ;
 wire \tt_process.tt_13n.connection[8] ;
 wire \tt_process.tt_13n.connection[9] ;
 wire \tt_samplekey.bitsadjacent[0] ;
 wire \tt_samplekey.bitsadjacent[1] ;
 wire \tt_samplekey.bitsadjacent[2] ;
 wire \tt_samplekey.bitsadjacent[3] ;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire clknet_0_clk;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;

 sg13g2_inv_1 _165_ (.Y(_012_),
    .A(\tt_samplekey.bitsadjacent[3] ));
 sg13g2_inv_1 _166_ (.Y(_013_),
    .A(\tt_samplekey.bitsadjacent[0] ));
 sg13g2_inv_1 _167_ (.Y(_014_),
    .A(\tt_finalprocess.num2[3] ));
 sg13g2_inv_1 _168_ (.Y(_015_),
    .A(\tt_finalprocess.genblk1[0].multblock.multblockout ));
 sg13g2_inv_1 _169_ (.Y(_016_),
    .A(\tt_finalprocess.genblk1[1].multblock.multblockout ));
 sg13g2_inv_1 _170_ (.Y(_017_),
    .A(\tt_finalprocess.genblk1[2].multblock.multblockout ));
 sg13g2_inv_1 _171_ (.Y(_018_),
    .A(\tt_finalprocess.genblk1[3].multblock.multblockout ));
 sg13g2_xor2_1 _172_ (.B(net64),
    .A(net56),
    .X(_019_));
 sg13g2_xor2_1 _173_ (.B(net65),
    .A(net71),
    .X(_020_));
 sg13g2_xnor2_1 _174_ (.Y(_011_),
    .A(_019_),
    .B(_020_));
 sg13g2_nor2_1 _175_ (.A(_009_),
    .B(_012_),
    .Y(_021_));
 sg13g2_or2_1 _176_ (.X(_022_),
    .B(_021_),
    .A(net31));
 sg13g2_nand2_1 _177_ (.Y(_023_),
    .A(\tt_samplekey.bitsadjacent[3] ),
    .B(net31));
 sg13g2_and2_1 _178_ (.A(\tt_samplekey.bitsadjacent[0] ),
    .B(_023_),
    .X(_024_));
 sg13g2_nand2b_1 _179_ (.Y(_025_),
    .B(\tt_samplekey.bitsadjacent[0] ),
    .A_N(net31));
 sg13g2_nor2_1 _180_ (.A(\tt_samplekey.bitsadjacent[3] ),
    .B(_013_),
    .Y(_026_));
 sg13g2_a22oi_1 _181_ (.Y(_001_),
    .B1(_022_),
    .B2(_024_),
    .A2(_012_),
    .A1(_009_));
 sg13g2_nor3_1 _182_ (.A(\tt_samplekey.bitsadjacent[1] ),
    .B(_013_),
    .C(\tt_samplekey.bitsadjacent[2] ),
    .Y(_027_));
 sg13g2_nor2_2 _183_ (.A(\tt_samplekey.bitsadjacent[3] ),
    .B(net31),
    .Y(_028_));
 sg13g2_inv_1 _184_ (.Y(_029_),
    .A(_028_));
 sg13g2_nor3_1 _185_ (.A(_026_),
    .B(_027_),
    .C(_028_),
    .Y(_002_));
 sg13g2_a21oi_1 _186_ (.A1(\tt_samplekey.bitsadjacent[0] ),
    .A2(\tt_samplekey.bitsadjacent[2] ),
    .Y(_030_),
    .B1(_029_));
 sg13g2_nor2_1 _187_ (.A(\tt_samplekey.bitsadjacent[0] ),
    .B(\tt_samplekey.bitsadjacent[2] ),
    .Y(_031_));
 sg13g2_nor2b_1 _188_ (.A(_023_),
    .B_N(_031_),
    .Y(_032_));
 sg13g2_and3_1 _189_ (.X(_033_),
    .A(net31),
    .B(\tt_samplekey.bitsadjacent[0] ),
    .C(\tt_samplekey.bitsadjacent[2] ));
 sg13g2_nor3_1 _190_ (.A(_030_),
    .B(_032_),
    .C(_033_),
    .Y(_003_));
 sg13g2_a22oi_1 _191_ (.Y(_004_),
    .B1(_031_),
    .B2(_012_),
    .A2(_025_),
    .A1(_021_));
 sg13g2_nand2_1 _192_ (.Y(_034_),
    .A(\tt_samplekey.bitsadjacent[2] ),
    .B(_028_));
 sg13g2_a21oi_1 _193_ (.A1(_023_),
    .A2(_034_),
    .Y(_035_),
    .B1(_013_));
 sg13g2_xor2_1 _194_ (.B(_028_),
    .A(\tt_samplekey.bitsadjacent[2] ),
    .X(_036_));
 sg13g2_a21oi_1 _195_ (.A1(_013_),
    .A2(_036_),
    .Y(_005_),
    .B1(_035_));
 sg13g2_xnor2_1 _196_ (.Y(_037_),
    .A(net31),
    .B(\tt_samplekey.bitsadjacent[2] ));
 sg13g2_nor3_1 _197_ (.A(_012_),
    .B(_013_),
    .C(_037_),
    .Y(_038_));
 sg13g2_nor2_1 _198_ (.A(_030_),
    .B(_038_),
    .Y(_006_));
 sg13g2_nand2b_1 _199_ (.Y(\tt_finalprocess.genblk1[4].multblock.multblockout ),
    .B(net4),
    .A_N(\tt_finalprocess.genblk1[4].multblock.multblockout ));
 sg13g2_nand2_1 _200_ (.Y(\tt_finalprocess.genblk1[0].multblock.multblockout ),
    .A(net4),
    .B(_015_));
 sg13g2_nand2b_1 _201_ (.Y(\tt_finalprocess.genblk1[5].multblock.multblockout ),
    .B(net4),
    .A_N(\tt_finalprocess.genblk1[5].multblock.multblockout ));
 sg13g2_nand2_1 _202_ (.Y(\tt_finalprocess.genblk1[1].multblock.multblockout ),
    .A(net4),
    .B(_016_));
 sg13g2_nand2b_1 _203_ (.Y(\tt_finalprocess.genblk1[6].multblock.multblockout ),
    .B(net4),
    .A_N(\tt_finalprocess.genblk1[6].multblock.multblockout ));
 sg13g2_nand2_1 _204_ (.Y(\tt_finalprocess.genblk1[2].multblock.multblockout ),
    .A(net4),
    .B(_017_));
 sg13g2_nand2b_1 _205_ (.Y(\tt_finalprocess.genblk1[7].multblock.multblockout ),
    .B(net4),
    .A_N(\tt_finalprocess.genblk1[7].multblock.multblockout ));
 sg13g2_nand2_1 _206_ (.Y(\tt_finalprocess.genblk1[3].multblock.multblockout ),
    .A(net4),
    .B(_018_));
 sg13g2_nand2_1 _207_ (.Y(\tt_invring1.ringosc8[38].inv.cnt_bit_I.Y ),
    .A(net33),
    .B(\tt_invring1.ringosc8[38].inv.cnt_bit_I.Y ));
 sg13g2_nand2_1 _208_ (.Y(\tt_invring1.ringosc7[46].inv.cnt_bit_I.Y ),
    .A(net33),
    .B(\tt_invring1.ringosc7[46].inv.cnt_bit_I.Y ));
 sg13g2_nand2_1 _209_ (.Y(\tt_invring1.ringosc6[40].inv.cnt_bit_I.Y ),
    .A(net33),
    .B(\tt_invring1.ringosc6[40].inv.cnt_bit_I.Y ));
 sg13g2_nand2_1 _210_ (.Y(\tt_invring1.ringosc5[36].inv.cnt_bit_I.Y ),
    .A(net32),
    .B(\tt_invring1.ringosc5[36].inv.cnt_bit_I.Y ));
 sg13g2_nand2_1 _211_ (.Y(\tt_invring1.ringosc4[28].inv.cnt_bit_I.Y ),
    .A(net32),
    .B(\tt_invring1.ringosc4[28].inv.cnt_bit_I.Y ));
 sg13g2_nand2_1 _212_ (.Y(\tt_invring1.ringosc3[22].inv.cnt_bit_I.Y ),
    .A(net32),
    .B(\tt_invring1.ringosc3[22].inv.cnt_bit_I.Y ));
 sg13g2_nand2_1 _213_ (.Y(\tt_invring1.ringosc2[18].inv.cnt_bit_I.Y ),
    .A(net32),
    .B(\tt_invring1.ringosc2[18].inv.cnt_bit_I.Y ));
 sg13g2_nand2_1 _214_ (.Y(\tt_invring1.ringosc1[10].inv.cnt_bit_I.Y ),
    .A(net32),
    .B(\tt_invring1.ringosc1[10].inv.cnt_bit_I.Y ));
 sg13g2_nand2_1 _215_ (.Y(\tt_invring2.ringosc8[38].inv.cnt_bit_I.Y ),
    .A(net33),
    .B(\tt_invring2.ringosc8[38].inv.cnt_bit_I.Y ));
 sg13g2_nand2_1 _216_ (.Y(\tt_invring2.ringosc7[46].inv.cnt_bit_I.Y ),
    .A(net33),
    .B(\tt_invring2.ringosc7[46].inv.cnt_bit_I.Y ));
 sg13g2_nand2_1 _217_ (.Y(\tt_invring2.ringosc6[40].inv.cnt_bit_I.Y ),
    .A(net33),
    .B(\tt_invring2.ringosc6[40].inv.cnt_bit_I.Y ));
 sg13g2_nand2_1 _218_ (.Y(\tt_invring2.ringosc5[36].inv.cnt_bit_I.Y ),
    .A(net33),
    .B(\tt_invring2.ringosc5[36].inv.cnt_bit_I.Y ));
 sg13g2_nand2_1 _219_ (.Y(\tt_invring2.ringosc4[28].inv.cnt_bit_I.Y ),
    .A(net32),
    .B(\tt_invring2.ringosc4[28].inv.cnt_bit_I.Y ));
 sg13g2_nand2_1 _220_ (.Y(\tt_invring2.ringosc3[22].inv.cnt_bit_I.Y ),
    .A(net33),
    .B(\tt_invring2.ringosc3[22].inv.cnt_bit_I.Y ));
 sg13g2_nand2_1 _221_ (.Y(\tt_invring2.ringosc2[18].inv.cnt_bit_I.Y ),
    .A(net32),
    .B(\tt_invring2.ringosc2[18].inv.cnt_bit_I.Y ));
 sg13g2_nand2_1 _222_ (.Y(\tt_invring2.ringosc1[10].inv.cnt_bit_I.Y ),
    .A(net32),
    .B(\tt_invring2.ringosc1[10].inv.cnt_bit_I.Y ));
 sg13g2_nand2b_1 _223_ (.Y(_039_),
    .B(\tt_process.bitsgroup[0] ),
    .A_N(\tt_process.bitsgroup[1] ));
 sg13g2_xor2_1 _224_ (.B(\tt_process.tt_13n.connection[11] ),
    .A(\tt_process.tt_13n.connection[4] ),
    .X(_040_));
 sg13g2_xnor2_1 _225_ (.Y(_041_),
    .A(\tt_process.tt_13n.connection[3] ),
    .B(_040_));
 sg13g2_xor2_1 _226_ (.B(\tt_process.tt_13n.connection[9] ),
    .A(\tt_process.tt_13n.connection[7] ),
    .X(_042_));
 sg13g2_xnor2_1 _227_ (.Y(_043_),
    .A(\tt_process.tt_13n.connection[13] ),
    .B(_042_));
 sg13g2_xnor2_1 _228_ (.Y(_044_),
    .A(_041_),
    .B(_043_));
 sg13g2_xor2_1 _229_ (.B(\tt_process.tt_13n.connection[10] ),
    .A(\tt_process.tt_13n.connection[6] ),
    .X(_045_));
 sg13g2_xnor2_1 _230_ (.Y(_046_),
    .A(\tt_process.tt_13n.connection[8] ),
    .B(\tt_process.tt_13n.connection[12] ));
 sg13g2_xor2_1 _231_ (.B(\tt_process.tt_13n.connection[1] ),
    .A(\tt_process.tt_13n.connection[2] ),
    .X(_047_));
 sg13g2_xnor2_1 _232_ (.Y(_048_),
    .A(_045_),
    .B(_047_));
 sg13g2_xnor2_1 _233_ (.Y(_049_),
    .A(\tt_process.tt_13n.connection[5] ),
    .B(_046_));
 sg13g2_xnor2_1 _234_ (.Y(_050_),
    .A(_048_),
    .B(_049_));
 sg13g2_nor2b_1 _235_ (.A(\tt_process.bitsgroup[0] ),
    .B_N(\tt_process.bitsgroup[1] ),
    .Y(_051_));
 sg13g2_xnor2_1 _236_ (.Y(_052_),
    .A(_044_),
    .B(_050_));
 sg13g2_o21ai_1 _237_ (.B1(_039_),
    .Y(_053_),
    .A1(_051_),
    .A2(_052_));
 sg13g2_xnor2_1 _238_ (.Y(ranbitstring),
    .A(net71),
    .B(_053_));
 sg13g2_xnor2_1 _239_ (.Y(_054_),
    .A(\tt_invring2.ringoutsam[6] ),
    .B(\tt_invring2.ringoutsam[7] ));
 sg13g2_xnor2_1 _240_ (.Y(_055_),
    .A(\tt_invring2.ringoutsam[5] ),
    .B(_054_));
 sg13g2_xor2_1 _241_ (.B(\tt_invring2.ringoutsam[0] ),
    .A(\tt_invring2.ringoutsam[1] ),
    .X(_056_));
 sg13g2_xor2_1 _242_ (.B(\tt_invring2.ringoutsam[2] ),
    .A(\tt_invring2.ringoutsam[4] ),
    .X(_057_));
 sg13g2_xnor2_1 _243_ (.Y(_058_),
    .A(\tt_invring2.ringoutsam[3] ),
    .B(_057_));
 sg13g2_xnor2_1 _244_ (.Y(_059_),
    .A(_056_),
    .B(_058_));
 sg13g2_nor2_1 _245_ (.A(net1),
    .B(_008_),
    .Y(_060_));
 sg13g2_a21oi_1 _246_ (.A1(net1),
    .A2(_059_),
    .Y(_061_),
    .B1(_060_));
 sg13g2_xnor2_1 _247_ (.Y(_062_),
    .A(_055_),
    .B(_061_));
 sg13g2_xnor2_1 _248_ (.Y(_063_),
    .A(\tt_invring1.ringoutsam[6] ),
    .B(\tt_invring1.ringoutsam[7] ));
 sg13g2_xnor2_1 _249_ (.Y(_064_),
    .A(\tt_invring1.ringoutsam[5] ),
    .B(_063_));
 sg13g2_xor2_1 _250_ (.B(\tt_invring1.ringoutsam[0] ),
    .A(\tt_invring1.ringoutsam[1] ),
    .X(_065_));
 sg13g2_xor2_1 _251_ (.B(\tt_invring1.ringoutsam[2] ),
    .A(\tt_invring1.ringoutsam[4] ),
    .X(_066_));
 sg13g2_xnor2_1 _252_ (.Y(_067_),
    .A(\tt_invring1.ringoutsam[3] ),
    .B(_066_));
 sg13g2_xnor2_1 _253_ (.Y(_068_),
    .A(_065_),
    .B(_067_));
 sg13g2_nor2_1 _254_ (.A(net73),
    .B(net1),
    .Y(_069_));
 sg13g2_a21oi_1 _255_ (.A1(net1),
    .A2(_068_),
    .Y(_070_),
    .B1(_069_));
 sg13g2_xnor2_1 _256_ (.Y(_071_),
    .A(_064_),
    .B(_070_));
 sg13g2_mux2_1 _257_ (.A0(_071_),
    .A1(_062_),
    .S(net2),
    .X(inverterringout));
 sg13g2_o21ai_1 _258_ (.B1(net34),
    .Y(_072_),
    .A1(net5),
    .A2(\tt_finalprocess.genblk1[6].multblock.multblockout ));
 sg13g2_a21oi_2 _259_ (.B1(_072_),
    .Y(\tt_finalprocess.num2[2] ),
    .A2(_017_),
    .A1(net5));
 sg13g2_o21ai_1 _260_ (.B1(net34),
    .Y(_073_),
    .A1(net5),
    .A2(\tt_finalprocess.genblk1[5].multblock.multblockout ));
 sg13g2_a21oi_2 _261_ (.B1(_073_),
    .Y(\tt_finalprocess.num2[1] ),
    .A2(_016_),
    .A1(net5));
 sg13g2_o21ai_1 _262_ (.B1(net35),
    .Y(_074_),
    .A1(net5),
    .A2(\tt_finalprocess.genblk1[4].multblock.multblockout ));
 sg13g2_a21oi_2 _263_ (.B1(_074_),
    .Y(\tt_finalprocess.num2[0] ),
    .A2(_015_),
    .A1(net5));
 sg13g2_o21ai_1 _264_ (.B1(net35),
    .Y(_075_),
    .A1(net5),
    .A2(\tt_finalprocess.genblk1[7].multblock.multblockout ));
 sg13g2_a21oi_2 _265_ (.B1(_075_),
    .Y(\tt_finalprocess.num2[3] ),
    .A2(_018_),
    .A1(net5));
 sg13g2_nand2b_2 _266_ (.Y(_076_),
    .B(\tt_finalprocess.num2[0] ),
    .A_N(\tt_finalprocess.num2[1] ));
 sg13g2_inv_1 _267_ (.Y(_077_),
    .A(_076_));
 sg13g2_nand2b_1 _268_ (.Y(_078_),
    .B(_076_),
    .A_N(net44));
 sg13g2_nand2_1 _269_ (.Y(_079_),
    .A(\tt_finalprocess.num2[1] ),
    .B(\tt_finalprocess.num2[0] ));
 sg13g2_a21oi_1 _270_ (.A1(net44),
    .A2(_079_),
    .Y(_080_),
    .B1(\tt_finalprocess.num2[3] ));
 sg13g2_nor2_1 _271_ (.A(\tt_finalprocess.num2[1] ),
    .B(\tt_finalprocess.num2[0] ),
    .Y(_081_));
 sg13g2_and2_1 _272_ (.A(net44),
    .B(\tt_finalprocess.num2[3] ),
    .X(_082_));
 sg13g2_a22oi_1 _273_ (.Y(uio_out[0]),
    .B1(_081_),
    .B2(_082_),
    .A2(_080_),
    .A1(_078_));
 sg13g2_a21oi_1 _274_ (.A1(_077_),
    .A2(_082_),
    .Y(uio_out[1]),
    .B1(_080_));
 sg13g2_nand2b_1 _275_ (.Y(_083_),
    .B(\tt_finalprocess.num2[1] ),
    .A_N(\tt_finalprocess.num2[0] ));
 sg13g2_nor2_1 _276_ (.A(\tt_finalprocess.num2[2] ),
    .B(\tt_finalprocess.num2[1] ),
    .Y(_084_));
 sg13g2_a22oi_1 _277_ (.Y(uio_out[2]),
    .B1(_084_),
    .B2(\tt_finalprocess.num2[0] ),
    .A2(_083_),
    .A1(_014_));
 sg13g2_nand3_1 _278_ (.B(_076_),
    .C(_083_),
    .A(net44),
    .Y(_085_));
 sg13g2_nor2_1 _279_ (.A(\tt_finalprocess.num2[3] ),
    .B(_084_),
    .Y(_086_));
 sg13g2_mux2_1 _280_ (.A0(_083_),
    .A1(_079_),
    .S(\tt_finalprocess.num2[2] ),
    .X(_087_));
 sg13g2_a22oi_1 _281_ (.Y(_088_),
    .B1(_087_),
    .B2(\tt_finalprocess.num2[3] ),
    .A2(_086_),
    .A1(_085_));
 sg13g2_inv_1 _282_ (.Y(uio_out[3]),
    .A(_088_));
 sg13g2_nor2_1 _283_ (.A(net44),
    .B(\tt_finalprocess.num2[0] ),
    .Y(_089_));
 sg13g2_a22oi_1 _284_ (.Y(uio_out[4]),
    .B1(_089_),
    .B2(_014_),
    .A2(_082_),
    .A1(_076_));
 sg13g2_nor2_1 _285_ (.A(net44),
    .B(_081_),
    .Y(_090_));
 sg13g2_nor2_1 _286_ (.A(\tt_finalprocess.num2[3] ),
    .B(_090_),
    .Y(_091_));
 sg13g2_a21oi_1 _287_ (.A1(\tt_finalprocess.num2[1] ),
    .A2(\tt_finalprocess.num2[0] ),
    .Y(_092_),
    .B1(net44));
 sg13g2_nor2_1 _288_ (.A(_014_),
    .B(_092_),
    .Y(_093_));
 sg13g2_a22oi_1 _289_ (.Y(uio_out[5]),
    .B1(_093_),
    .B2(_076_),
    .A2(_091_),
    .A1(_085_));
 sg13g2_nand2b_1 _290_ (.Y(_094_),
    .B(_086_),
    .A_N(_081_));
 sg13g2_a21oi_1 _291_ (.A1(net44),
    .A2(_076_),
    .Y(_095_),
    .B1(_092_));
 sg13g2_o21ai_1 _292_ (.B1(_094_),
    .Y(uio_out[6]),
    .A1(_014_),
    .A2(_095_));
 sg13g2_nor2_1 _293_ (.A(net31),
    .B(\tt_samplekey.bitsadjacent[0] ),
    .Y(_096_));
 sg13g2_a22oi_1 _294_ (.Y(_000_),
    .B1(_096_),
    .B2(_021_),
    .A2(_037_),
    .A1(_026_));
 sg13g2_dfrbp_1 _295_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net40),
    .D(\tt_invring1.ringosc1[10].inv.cnt_bit_I.Y ),
    .Q_N(_100_),
    .Q(\tt_invring1.ringoutsam[0] ));
 sg13g2_dfrbp_1 _296_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net40),
    .D(\tt_invring1.ringosc2[18].inv.cnt_bit_I.Y ),
    .Q_N(_101_),
    .Q(\tt_invring1.ringoutsam[1] ));
 sg13g2_dfrbp_1 _297_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net40),
    .D(\tt_invring1.ringosc3[22].inv.cnt_bit_I.Y ),
    .Q_N(_102_),
    .Q(\tt_invring1.ringoutsam[2] ));
 sg13g2_dfrbp_1 _298_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net40),
    .D(\tt_invring1.ringosc4[28].inv.cnt_bit_I.Y ),
    .Q_N(_103_),
    .Q(\tt_invring1.ringoutsam[3] ));
 sg13g2_dfrbp_1 _299_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net40),
    .D(\tt_invring1.ringosc5[36].inv.cnt_bit_I.Y ),
    .Q_N(_007_),
    .Q(\tt_invring1.ringoutsam[4] ));
 sg13g2_dfrbp_1 _300_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net38),
    .D(\tt_invring1.ringosc6[40].inv.cnt_bit_I.Y ),
    .Q_N(_104_),
    .Q(\tt_invring1.ringoutsam[5] ));
 sg13g2_dfrbp_1 _301_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net38),
    .D(\tt_invring1.ringosc7[46].inv.cnt_bit_I.Y ),
    .Q_N(_105_),
    .Q(\tt_invring1.ringoutsam[6] ));
 sg13g2_dfrbp_1 _302_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net38),
    .D(\tt_invring1.ringosc8[38].inv.cnt_bit_I.Y ),
    .Q_N(_106_),
    .Q(\tt_invring1.ringoutsam[7] ));
 sg13g2_dfrbp_1 _303_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net40),
    .D(\tt_invring2.ringosc1[10].inv.cnt_bit_I.Y ),
    .Q_N(_107_),
    .Q(\tt_invring2.ringoutsam[0] ));
 sg13g2_dfrbp_1 _304_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net40),
    .D(\tt_invring2.ringosc2[18].inv.cnt_bit_I.Y ),
    .Q_N(_108_),
    .Q(\tt_invring2.ringoutsam[1] ));
 sg13g2_dfrbp_1 _305_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net41),
    .D(\tt_invring2.ringosc3[22].inv.cnt_bit_I.Y ),
    .Q_N(_109_),
    .Q(\tt_invring2.ringoutsam[2] ));
 sg13g2_dfrbp_1 _306_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net41),
    .D(\tt_invring2.ringosc4[28].inv.cnt_bit_I.Y ),
    .Q_N(_110_),
    .Q(\tt_invring2.ringoutsam[3] ));
 sg13g2_dfrbp_1 _307_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net40),
    .D(\tt_invring2.ringosc5[36].inv.cnt_bit_I.Y ),
    .Q_N(_008_),
    .Q(\tt_invring2.ringoutsam[4] ));
 sg13g2_dfrbp_1 _308_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net38),
    .D(\tt_invring2.ringosc6[40].inv.cnt_bit_I.Y ),
    .Q_N(_111_),
    .Q(\tt_invring2.ringoutsam[5] ));
 sg13g2_dfrbp_1 _309_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net42),
    .D(\tt_invring2.ringosc7[46].inv.cnt_bit_I.Y ),
    .Q_N(_112_),
    .Q(\tt_invring2.ringoutsam[6] ));
 sg13g2_dfrbp_1 _310_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net42),
    .D(\tt_invring2.ringosc8[38].inv.cnt_bit_I.Y ),
    .Q_N(_113_),
    .Q(\tt_invring2.ringoutsam[7] ));
 sg13g2_dfrbp_1 _311_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net38),
    .D(net27),
    .Q_N(_114_),
    .Q(\tt_process.tt_13n.connection[0] ));
 sg13g2_dfrbp_1 _312_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net38),
    .D(net51),
    .Q_N(_115_),
    .Q(\tt_process.tt_13n.connection[1] ));
 sg13g2_dfrbp_1 _313_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net38),
    .D(net54),
    .Q_N(_116_),
    .Q(\tt_process.tt_13n.connection[2] ));
 sg13g2_dfrbp_1 _314_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net38),
    .D(net67),
    .Q_N(_117_),
    .Q(\tt_process.tt_13n.connection[3] ));
 sg13g2_dfrbp_1 _315_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net39),
    .D(net68),
    .Q_N(_118_),
    .Q(\tt_process.tt_13n.connection[4] ));
 sg13g2_dfrbp_1 _316_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net39),
    .D(net61),
    .Q_N(_119_),
    .Q(\tt_process.tt_13n.connection[5] ));
 sg13g2_dfrbp_1 _317_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net39),
    .D(net62),
    .Q_N(_120_),
    .Q(\tt_process.tt_13n.connection[6] ));
 sg13g2_dfrbp_1 _318_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net41),
    .D(net58),
    .Q_N(_121_),
    .Q(\tt_process.tt_13n.connection[7] ));
 sg13g2_dfrbp_1 _319_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net41),
    .D(net60),
    .Q_N(_122_),
    .Q(\tt_process.tt_13n.connection[8] ));
 sg13g2_dfrbp_1 _320_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net39),
    .D(net63),
    .Q_N(_123_),
    .Q(\tt_process.tt_13n.connection[9] ));
 sg13g2_dfrbp_1 _321_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net39),
    .D(net66),
    .Q_N(_124_),
    .Q(\tt_process.tt_13n.connection[10] ));
 sg13g2_dfrbp_1 _322_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net39),
    .D(net59),
    .Q_N(_125_),
    .Q(\tt_process.tt_13n.connection[11] ));
 sg13g2_dfrbp_1 _323_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net39),
    .D(net55),
    .Q_N(_126_),
    .Q(\tt_process.tt_13n.connection[12] ));
 sg13g2_dfrbp_1 _324_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net39),
    .D(net57),
    .Q_N(_127_),
    .Q(\tt_process.tt_13n.connection[13] ));
 sg13g2_dfrbp_1 _325_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net37),
    .D(net24),
    .Q_N(_097_),
    .Q(\tt_process.clk_half ));
 sg13g2_dfrbp_1 _326_ (.CLK(\tt_process.clk_half ),
    .RESET_B(net7),
    .D(\tt_process.bitsadjacent[0] ),
    .Q_N(_128_),
    .Q(\tt_process.bitsgroup[0] ));
 sg13g2_dfrbp_1 _327_ (.CLK(\tt_process.clk_half ),
    .RESET_B(net8),
    .D(\tt_process.bitsadjacent[1] ),
    .Q_N(_129_),
    .Q(\tt_process.bitsgroup[1] ));
 sg13g2_dfrbp_1 _328_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net37),
    .D(net74),
    .Q_N(_130_),
    .Q(\tt_process.bitsadjacent[0] ));
 sg13g2_dfrbp_1 _329_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net37),
    .D(net53),
    .Q_N(_131_),
    .Q(\tt_process.bitsadjacent[1] ));
 sg13g2_dfrbp_1 _330_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net37),
    .D(net50),
    .Q_N(_099_),
    .Q(\tt_process.bitsadjacent[2] ));
 sg13g2_dfrbp_1 _331_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net34),
    .D(_011_),
    .Q_N(\tt_16bitran.connection[1] ),
    .Q(_010_));
 sg13g2_dfrbp_1 _332_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net34),
    .D(net23),
    .Q_N(_132_),
    .Q(\tt_16bitran.connection[2] ));
 sg13g2_dfrbp_1 _333_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net34),
    .D(net28),
    .Q_N(_133_),
    .Q(\tt_16bitran.connection[3] ));
 sg13g2_dfrbp_1 _334_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net34),
    .D(net45),
    .Q_N(_134_),
    .Q(\tt_16bitran.connection[4] ));
 sg13g2_dfrbp_1 _335_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net34),
    .D(net56),
    .Q_N(_135_),
    .Q(\tt_16bitran.connection[5] ));
 sg13g2_dfrbp_1 _336_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net34),
    .D(net49),
    .Q_N(_136_),
    .Q(\tt_16bitran.connection[6] ));
 sg13g2_dfrbp_1 _337_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net36),
    .D(net25),
    .Q_N(_137_),
    .Q(\tt_16bitran.connection[7] ));
 sg13g2_dfrbp_1 _338_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net36),
    .D(net26),
    .Q_N(_138_),
    .Q(\tt_16bitran.connection[8] ));
 sg13g2_dfrbp_1 _339_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net36),
    .D(net47),
    .Q_N(_139_),
    .Q(\tt_16bitran.connection[9] ));
 sg13g2_dfrbp_1 _340_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net36),
    .D(net46),
    .Q_N(_140_),
    .Q(\tt_16bitran.connection[10] ));
 sg13g2_dfrbp_1 _341_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net37),
    .D(net29),
    .Q_N(_141_),
    .Q(\tt_16bitran.connection[11] ));
 sg13g2_dfrbp_1 _342_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net37),
    .D(net30),
    .Q_N(_142_),
    .Q(\tt_16bitran.connection[12] ));
 sg13g2_dfrbp_1 _343_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net36),
    .D(net52),
    .Q_N(_143_),
    .Q(\tt_16bitran.connection[13] ));
 sg13g2_dfrbp_1 _344_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net36),
    .D(net65),
    .Q_N(_144_),
    .Q(\tt_16bitran.connection[14] ));
 sg13g2_dfrbp_1 _345_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net36),
    .D(net48),
    .Q_N(_145_),
    .Q(\tt_16bitran.connection[15] ));
 sg13g2_dfrbp_1 _346_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net36),
    .D(net64),
    .Q_N(_146_),
    .Q(ran16out));
 sg13g2_dfrbp_1 _347_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net35),
    .D(ranbitstring),
    .Q_N(_147_),
    .Q(\tt_samplekey.bitsadjacent[0] ));
 sg13g2_dfrbp_1 _348_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net35),
    .D(net69),
    .Q_N(_148_),
    .Q(\tt_samplekey.bitsadjacent[1] ));
 sg13g2_dfrbp_1 _349_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net35),
    .D(net31),
    .Q_N(_009_),
    .Q(\tt_samplekey.bitsadjacent[2] ));
 sg13g2_dfrbp_1 _350_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net35),
    .D(net70),
    .Q_N(_149_),
    .Q(\tt_samplekey.bitsadjacent[3] ));
 sg13g2_dfrbp_1 _351_ (.CLK(net3),
    .RESET_B(net10),
    .D(_000_),
    .Q_N(_150_),
    .Q(uo_out[0]));
 sg13g2_dfrbp_1 _352_ (.CLK(net3),
    .RESET_B(net11),
    .D(_001_),
    .Q_N(_151_),
    .Q(uo_out[1]));
 sg13g2_dfrbp_1 _353_ (.CLK(net3),
    .RESET_B(net12),
    .D(_002_),
    .Q_N(_152_),
    .Q(uo_out[2]));
 sg13g2_dfrbp_1 _354_ (.CLK(net3),
    .RESET_B(net13),
    .D(_003_),
    .Q_N(_153_),
    .Q(uo_out[3]));
 sg13g2_dfrbp_1 _355_ (.CLK(net3),
    .RESET_B(net14),
    .D(_004_),
    .Q_N(_154_),
    .Q(uo_out[4]));
 sg13g2_dfrbp_1 _356_ (.CLK(net3),
    .RESET_B(net6),
    .D(_005_),
    .Q_N(_155_),
    .Q(uo_out[5]));
 sg13g2_dfrbp_1 _357_ (.CLK(net3),
    .RESET_B(net9),
    .D(_006_),
    .Q_N(_098_),
    .Q(uo_out[6]));
 sg13g2_tiehi _326__7 (.L_HI(net7));
 sg13g2_tiehi _327__8 (.L_HI(net8));
 sg13g2_tiehi _357__9 (.L_HI(net9));
 sg13g2_tiehi _351__10 (.L_HI(net10));
 sg13g2_tiehi _352__11 (.L_HI(net11));
 sg13g2_tiehi _353__12 (.L_HI(net12));
 sg13g2_tiehi _354__13 (.L_HI(net13));
 sg13g2_tiehi _355__14 (.L_HI(net14));
 sg13g2_tiehi tt_um_ran_DanielZhu_15 (.L_HI(net15));
 sg13g2_tiehi tt_um_ran_DanielZhu_16 (.L_HI(net16));
 sg13g2_tiehi tt_um_ran_DanielZhu_17 (.L_HI(net17));
 sg13g2_tiehi tt_um_ran_DanielZhu_18 (.L_HI(net18));
 sg13g2_tiehi tt_um_ran_DanielZhu_19 (.L_HI(net19));
 sg13g2_tiehi tt_um_ran_DanielZhu_20 (.L_HI(net20));
 sg13g2_tiehi tt_um_ran_DanielZhu_21 (.L_HI(net21));
 sg13g2_tiehi tt_um_ran_DanielZhu_22 (.L_HI(net22));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_1 _375_ (.A(ranbitstring),
    .X(uio_out[7]));
 sg13g2_buf_1 _376_ (.A(inverterringout),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout31 (.A(net72),
    .X(net31));
 sg13g2_buf_2 fanout32 (.A(ui_in[0]),
    .X(net32));
 sg13g2_buf_2 fanout33 (.A(ui_in[0]),
    .X(net33));
 sg13g2_buf_4 fanout34 (.X(net34),
    .A(net43));
 sg13g2_buf_2 fanout35 (.A(net43),
    .X(net35));
 sg13g2_buf_4 fanout36 (.X(net36),
    .A(net37));
 sg13g2_buf_4 fanout37 (.X(net37),
    .A(net43));
 sg13g2_buf_4 fanout38 (.X(net38),
    .A(net42));
 sg13g2_buf_4 fanout39 (.X(net39),
    .A(net41));
 sg13g2_buf_4 fanout40 (.X(net40),
    .A(net41));
 sg13g2_buf_4 fanout41 (.X(net41),
    .A(net42));
 sg13g2_buf_2 fanout42 (.A(net43),
    .X(net42));
 sg13g2_buf_2 fanout43 (.A(rst_n),
    .X(net43));
 sg13g2_buf_2 fanout44 (.A(\tt_finalprocess.num2[2] ),
    .X(net44));
 sg13g2_buf_1 input1 (.A(ui_in[1]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[2]),
    .X(net2));
 sg13g2_buf_2 input3 (.A(ui_in[3]),
    .X(net3));
 sg13g2_buf_2 input4 (.A(ui_in[4]),
    .X(net4));
 sg13g2_buf_4 input5 (.X(net5),
    .A(ui_in[5]));
 sg13g2_tiehi _356__6 (.L_HI(net6));
 sg13g2_buf_2 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sg13g2_buf_2 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sg13g2_buf_2 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sg13g2_buf_2 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sg13g2_buf_2 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sg13g2_buf_2 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sg13g2_buf_2 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sg13g2_buf_2 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_3_3__leaf_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_3_7__leaf_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\tt_16bitran.connection[1] ),
    .X(net23));
 sg13g2_dlygate4sd3_1 hold2 (.A(_097_),
    .X(net24));
 sg13g2_dlygate4sd3_1 hold3 (.A(\tt_16bitran.connection[6] ),
    .X(net25));
 sg13g2_dlygate4sd3_1 hold4 (.A(\tt_16bitran.connection[7] ),
    .X(net26));
 sg13g2_dlygate4sd3_1 hold5 (.A(\tt_process.bitsadjacent[2] ),
    .X(net27));
 sg13g2_dlygate4sd3_1 hold6 (.A(\tt_16bitran.connection[2] ),
    .X(net28));
 sg13g2_dlygate4sd3_1 hold7 (.A(\tt_16bitran.connection[10] ),
    .X(net29));
 sg13g2_dlygate4sd3_1 hold8 (.A(\tt_16bitran.connection[11] ),
    .X(net30));
 sg13g2_dlygate4sd3_1 hold9 (.A(\tt_16bitran.connection[3] ),
    .X(net45));
 sg13g2_dlygate4sd3_1 hold10 (.A(\tt_16bitran.connection[9] ),
    .X(net46));
 sg13g2_dlygate4sd3_1 hold11 (.A(\tt_16bitran.connection[8] ),
    .X(net47));
 sg13g2_dlygate4sd3_1 hold12 (.A(\tt_16bitran.connection[14] ),
    .X(net48));
 sg13g2_dlygate4sd3_1 hold13 (.A(\tt_16bitran.connection[5] ),
    .X(net49));
 sg13g2_dlygate4sd3_1 hold14 (.A(\tt_process.bitsadjacent[1] ),
    .X(net50));
 sg13g2_dlygate4sd3_1 hold15 (.A(\tt_process.tt_13n.connection[0] ),
    .X(net51));
 sg13g2_dlygate4sd3_1 hold16 (.A(\tt_16bitran.connection[12] ),
    .X(net52));
 sg13g2_dlygate4sd3_1 hold17 (.A(\tt_process.bitsadjacent[0] ),
    .X(net53));
 sg13g2_dlygate4sd3_1 hold18 (.A(\tt_process.tt_13n.connection[1] ),
    .X(net54));
 sg13g2_dlygate4sd3_1 hold19 (.A(\tt_process.tt_13n.connection[11] ),
    .X(net55));
 sg13g2_dlygate4sd3_1 hold20 (.A(\tt_16bitran.connection[4] ),
    .X(net56));
 sg13g2_dlygate4sd3_1 hold21 (.A(\tt_process.tt_13n.connection[12] ),
    .X(net57));
 sg13g2_dlygate4sd3_1 hold22 (.A(\tt_process.tt_13n.connection[6] ),
    .X(net58));
 sg13g2_dlygate4sd3_1 hold23 (.A(\tt_process.tt_13n.connection[10] ),
    .X(net59));
 sg13g2_dlygate4sd3_1 hold24 (.A(\tt_process.tt_13n.connection[7] ),
    .X(net60));
 sg13g2_dlygate4sd3_1 hold25 (.A(\tt_process.tt_13n.connection[4] ),
    .X(net61));
 sg13g2_dlygate4sd3_1 hold26 (.A(\tt_process.tt_13n.connection[5] ),
    .X(net62));
 sg13g2_dlygate4sd3_1 hold27 (.A(\tt_process.tt_13n.connection[8] ),
    .X(net63));
 sg13g2_dlygate4sd3_1 hold28 (.A(\tt_16bitran.connection[15] ),
    .X(net64));
 sg13g2_dlygate4sd3_1 hold29 (.A(\tt_16bitran.connection[13] ),
    .X(net65));
 sg13g2_dlygate4sd3_1 hold30 (.A(\tt_process.tt_13n.connection[9] ),
    .X(net66));
 sg13g2_dlygate4sd3_1 hold31 (.A(\tt_process.tt_13n.connection[2] ),
    .X(net67));
 sg13g2_dlygate4sd3_1 hold32 (.A(\tt_process.tt_13n.connection[3] ),
    .X(net68));
 sg13g2_dlygate4sd3_1 hold33 (.A(\tt_samplekey.bitsadjacent[0] ),
    .X(net69));
 sg13g2_dlygate4sd3_1 hold34 (.A(\tt_samplekey.bitsadjacent[2] ),
    .X(net70));
 sg13g2_dlygate4sd3_1 hold35 (.A(ran16out),
    .X(net71));
 sg13g2_dlygate4sd3_1 hold36 (.A(\tt_samplekey.bitsadjacent[1] ),
    .X(net72));
 sg13g2_dlygate4sd3_1 hold37 (.A(_007_),
    .X(net73));
 sg13g2_dlygate4sd3_1 hold38 (.A(inverterringout),
    .X(net74));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_fill_2 FILLER_14_406 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_252 ();
 sg13g2_decap_8 FILLER_15_259 ();
 sg13g2_decap_8 FILLER_15_266 ();
 sg13g2_decap_8 FILLER_15_273 ();
 sg13g2_decap_8 FILLER_15_280 ();
 sg13g2_decap_8 FILLER_15_287 ();
 sg13g2_decap_8 FILLER_15_294 ();
 sg13g2_decap_8 FILLER_15_301 ();
 sg13g2_decap_8 FILLER_15_308 ();
 sg13g2_decap_8 FILLER_15_315 ();
 sg13g2_decap_8 FILLER_15_322 ();
 sg13g2_decap_8 FILLER_15_329 ();
 sg13g2_decap_8 FILLER_15_336 ();
 sg13g2_decap_8 FILLER_15_343 ();
 sg13g2_decap_8 FILLER_15_350 ();
 sg13g2_decap_8 FILLER_15_357 ();
 sg13g2_decap_8 FILLER_15_364 ();
 sg13g2_decap_8 FILLER_15_371 ();
 sg13g2_decap_8 FILLER_15_378 ();
 sg13g2_decap_8 FILLER_15_385 ();
 sg13g2_decap_8 FILLER_15_392 ();
 sg13g2_decap_8 FILLER_15_399 ();
 sg13g2_fill_2 FILLER_15_406 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_decap_8 FILLER_16_217 ();
 sg13g2_decap_8 FILLER_16_224 ();
 sg13g2_decap_8 FILLER_16_231 ();
 sg13g2_decap_8 FILLER_16_238 ();
 sg13g2_decap_8 FILLER_16_245 ();
 sg13g2_decap_8 FILLER_16_252 ();
 sg13g2_decap_8 FILLER_16_259 ();
 sg13g2_decap_8 FILLER_16_266 ();
 sg13g2_decap_8 FILLER_16_273 ();
 sg13g2_decap_8 FILLER_16_280 ();
 sg13g2_decap_8 FILLER_16_287 ();
 sg13g2_decap_8 FILLER_16_294 ();
 sg13g2_decap_8 FILLER_16_301 ();
 sg13g2_decap_8 FILLER_16_308 ();
 sg13g2_decap_8 FILLER_16_315 ();
 sg13g2_decap_8 FILLER_16_322 ();
 sg13g2_decap_8 FILLER_16_329 ();
 sg13g2_decap_8 FILLER_16_336 ();
 sg13g2_decap_8 FILLER_16_343 ();
 sg13g2_decap_8 FILLER_16_350 ();
 sg13g2_decap_8 FILLER_16_357 ();
 sg13g2_decap_8 FILLER_16_364 ();
 sg13g2_decap_8 FILLER_16_371 ();
 sg13g2_decap_8 FILLER_16_378 ();
 sg13g2_decap_8 FILLER_16_385 ();
 sg13g2_decap_8 FILLER_16_392 ();
 sg13g2_decap_8 FILLER_16_399 ();
 sg13g2_fill_2 FILLER_16_406 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_decap_8 FILLER_17_168 ();
 sg13g2_decap_8 FILLER_17_175 ();
 sg13g2_decap_8 FILLER_17_182 ();
 sg13g2_decap_8 FILLER_17_189 ();
 sg13g2_decap_8 FILLER_17_196 ();
 sg13g2_decap_8 FILLER_17_203 ();
 sg13g2_decap_8 FILLER_17_210 ();
 sg13g2_decap_8 FILLER_17_217 ();
 sg13g2_decap_8 FILLER_17_224 ();
 sg13g2_decap_8 FILLER_17_231 ();
 sg13g2_decap_8 FILLER_17_238 ();
 sg13g2_decap_8 FILLER_17_245 ();
 sg13g2_decap_8 FILLER_17_252 ();
 sg13g2_decap_8 FILLER_17_259 ();
 sg13g2_decap_8 FILLER_17_266 ();
 sg13g2_decap_8 FILLER_17_273 ();
 sg13g2_decap_8 FILLER_17_280 ();
 sg13g2_decap_8 FILLER_17_287 ();
 sg13g2_decap_8 FILLER_17_294 ();
 sg13g2_decap_8 FILLER_17_301 ();
 sg13g2_decap_8 FILLER_17_308 ();
 sg13g2_decap_8 FILLER_17_315 ();
 sg13g2_decap_8 FILLER_17_322 ();
 sg13g2_decap_8 FILLER_17_329 ();
 sg13g2_decap_8 FILLER_17_336 ();
 sg13g2_decap_8 FILLER_17_343 ();
 sg13g2_decap_8 FILLER_17_350 ();
 sg13g2_decap_8 FILLER_17_357 ();
 sg13g2_decap_8 FILLER_17_364 ();
 sg13g2_decap_8 FILLER_17_371 ();
 sg13g2_decap_8 FILLER_17_378 ();
 sg13g2_decap_8 FILLER_17_385 ();
 sg13g2_decap_8 FILLER_17_392 ();
 sg13g2_decap_8 FILLER_17_399 ();
 sg13g2_fill_2 FILLER_17_406 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_decap_8 FILLER_18_147 ();
 sg13g2_decap_8 FILLER_18_154 ();
 sg13g2_decap_8 FILLER_18_161 ();
 sg13g2_decap_8 FILLER_18_168 ();
 sg13g2_decap_8 FILLER_18_175 ();
 sg13g2_decap_8 FILLER_18_182 ();
 sg13g2_decap_8 FILLER_18_189 ();
 sg13g2_decap_8 FILLER_18_196 ();
 sg13g2_decap_8 FILLER_18_203 ();
 sg13g2_decap_8 FILLER_18_210 ();
 sg13g2_decap_8 FILLER_18_217 ();
 sg13g2_decap_8 FILLER_18_224 ();
 sg13g2_decap_8 FILLER_18_231 ();
 sg13g2_decap_8 FILLER_18_238 ();
 sg13g2_decap_8 FILLER_18_245 ();
 sg13g2_decap_8 FILLER_18_252 ();
 sg13g2_decap_8 FILLER_18_259 ();
 sg13g2_decap_8 FILLER_18_266 ();
 sg13g2_decap_8 FILLER_18_273 ();
 sg13g2_decap_8 FILLER_18_280 ();
 sg13g2_decap_8 FILLER_18_287 ();
 sg13g2_decap_8 FILLER_18_294 ();
 sg13g2_decap_8 FILLER_18_301 ();
 sg13g2_decap_8 FILLER_18_308 ();
 sg13g2_decap_8 FILLER_18_315 ();
 sg13g2_decap_8 FILLER_18_322 ();
 sg13g2_decap_8 FILLER_18_329 ();
 sg13g2_decap_8 FILLER_18_336 ();
 sg13g2_decap_8 FILLER_18_343 ();
 sg13g2_decap_8 FILLER_18_350 ();
 sg13g2_decap_8 FILLER_18_357 ();
 sg13g2_decap_8 FILLER_18_364 ();
 sg13g2_decap_8 FILLER_18_371 ();
 sg13g2_decap_8 FILLER_18_378 ();
 sg13g2_decap_8 FILLER_18_385 ();
 sg13g2_decap_8 FILLER_18_392 ();
 sg13g2_decap_8 FILLER_18_399 ();
 sg13g2_fill_2 FILLER_18_406 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_decap_8 FILLER_19_140 ();
 sg13g2_decap_8 FILLER_19_147 ();
 sg13g2_decap_8 FILLER_19_154 ();
 sg13g2_decap_8 FILLER_19_161 ();
 sg13g2_decap_8 FILLER_19_168 ();
 sg13g2_decap_8 FILLER_19_175 ();
 sg13g2_decap_8 FILLER_19_182 ();
 sg13g2_decap_8 FILLER_19_189 ();
 sg13g2_decap_8 FILLER_19_196 ();
 sg13g2_decap_8 FILLER_19_203 ();
 sg13g2_decap_8 FILLER_19_210 ();
 sg13g2_decap_8 FILLER_19_217 ();
 sg13g2_decap_8 FILLER_19_224 ();
 sg13g2_decap_8 FILLER_19_231 ();
 sg13g2_decap_8 FILLER_19_238 ();
 sg13g2_decap_8 FILLER_19_245 ();
 sg13g2_decap_8 FILLER_19_252 ();
 sg13g2_decap_8 FILLER_19_259 ();
 sg13g2_decap_8 FILLER_19_266 ();
 sg13g2_decap_8 FILLER_19_273 ();
 sg13g2_decap_8 FILLER_19_280 ();
 sg13g2_decap_8 FILLER_19_287 ();
 sg13g2_decap_8 FILLER_19_294 ();
 sg13g2_decap_8 FILLER_19_301 ();
 sg13g2_decap_8 FILLER_19_308 ();
 sg13g2_decap_8 FILLER_19_315 ();
 sg13g2_decap_8 FILLER_19_322 ();
 sg13g2_decap_8 FILLER_19_329 ();
 sg13g2_decap_8 FILLER_19_336 ();
 sg13g2_decap_8 FILLER_19_343 ();
 sg13g2_decap_8 FILLER_19_350 ();
 sg13g2_decap_8 FILLER_19_357 ();
 sg13g2_decap_8 FILLER_19_364 ();
 sg13g2_decap_8 FILLER_19_371 ();
 sg13g2_decap_8 FILLER_19_378 ();
 sg13g2_decap_8 FILLER_19_385 ();
 sg13g2_decap_8 FILLER_19_392 ();
 sg13g2_decap_8 FILLER_19_399 ();
 sg13g2_fill_2 FILLER_19_406 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_decap_8 FILLER_20_126 ();
 sg13g2_decap_8 FILLER_20_133 ();
 sg13g2_decap_8 FILLER_20_140 ();
 sg13g2_decap_8 FILLER_20_147 ();
 sg13g2_decap_8 FILLER_20_154 ();
 sg13g2_decap_8 FILLER_20_161 ();
 sg13g2_decap_8 FILLER_20_168 ();
 sg13g2_decap_8 FILLER_20_175 ();
 sg13g2_decap_8 FILLER_20_182 ();
 sg13g2_decap_8 FILLER_20_189 ();
 sg13g2_decap_8 FILLER_20_196 ();
 sg13g2_decap_8 FILLER_20_203 ();
 sg13g2_decap_8 FILLER_20_210 ();
 sg13g2_decap_8 FILLER_20_217 ();
 sg13g2_decap_8 FILLER_20_224 ();
 sg13g2_decap_8 FILLER_20_231 ();
 sg13g2_decap_8 FILLER_20_238 ();
 sg13g2_decap_8 FILLER_20_245 ();
 sg13g2_decap_8 FILLER_20_252 ();
 sg13g2_decap_8 FILLER_20_259 ();
 sg13g2_decap_8 FILLER_20_266 ();
 sg13g2_decap_8 FILLER_20_273 ();
 sg13g2_decap_8 FILLER_20_280 ();
 sg13g2_decap_8 FILLER_20_287 ();
 sg13g2_decap_8 FILLER_20_294 ();
 sg13g2_decap_8 FILLER_20_301 ();
 sg13g2_decap_8 FILLER_20_308 ();
 sg13g2_decap_8 FILLER_20_315 ();
 sg13g2_decap_8 FILLER_20_322 ();
 sg13g2_decap_8 FILLER_20_329 ();
 sg13g2_decap_8 FILLER_20_336 ();
 sg13g2_decap_8 FILLER_20_343 ();
 sg13g2_decap_8 FILLER_20_350 ();
 sg13g2_decap_8 FILLER_20_357 ();
 sg13g2_decap_8 FILLER_20_364 ();
 sg13g2_decap_8 FILLER_20_371 ();
 sg13g2_decap_8 FILLER_20_378 ();
 sg13g2_decap_8 FILLER_20_385 ();
 sg13g2_decap_8 FILLER_20_392 ();
 sg13g2_decap_8 FILLER_20_399 ();
 sg13g2_fill_2 FILLER_20_406 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_decap_8 FILLER_21_119 ();
 sg13g2_decap_8 FILLER_21_126 ();
 sg13g2_decap_8 FILLER_21_133 ();
 sg13g2_decap_8 FILLER_21_140 ();
 sg13g2_decap_8 FILLER_21_147 ();
 sg13g2_decap_8 FILLER_21_154 ();
 sg13g2_decap_8 FILLER_21_161 ();
 sg13g2_decap_8 FILLER_21_168 ();
 sg13g2_decap_8 FILLER_21_175 ();
 sg13g2_decap_8 FILLER_21_182 ();
 sg13g2_decap_8 FILLER_21_189 ();
 sg13g2_decap_8 FILLER_21_196 ();
 sg13g2_decap_8 FILLER_21_203 ();
 sg13g2_decap_8 FILLER_21_210 ();
 sg13g2_decap_8 FILLER_21_217 ();
 sg13g2_decap_8 FILLER_21_224 ();
 sg13g2_decap_8 FILLER_21_231 ();
 sg13g2_decap_8 FILLER_21_238 ();
 sg13g2_decap_8 FILLER_21_245 ();
 sg13g2_decap_8 FILLER_21_252 ();
 sg13g2_decap_8 FILLER_21_259 ();
 sg13g2_decap_8 FILLER_21_266 ();
 sg13g2_decap_8 FILLER_21_273 ();
 sg13g2_decap_8 FILLER_21_280 ();
 sg13g2_decap_8 FILLER_21_287 ();
 sg13g2_decap_8 FILLER_21_294 ();
 sg13g2_decap_8 FILLER_21_301 ();
 sg13g2_decap_8 FILLER_21_308 ();
 sg13g2_decap_8 FILLER_21_315 ();
 sg13g2_decap_8 FILLER_21_322 ();
 sg13g2_decap_8 FILLER_21_329 ();
 sg13g2_decap_8 FILLER_21_336 ();
 sg13g2_decap_8 FILLER_21_343 ();
 sg13g2_decap_8 FILLER_21_350 ();
 sg13g2_decap_8 FILLER_21_357 ();
 sg13g2_decap_8 FILLER_21_364 ();
 sg13g2_decap_8 FILLER_21_371 ();
 sg13g2_decap_8 FILLER_21_378 ();
 sg13g2_decap_8 FILLER_21_385 ();
 sg13g2_decap_8 FILLER_21_392 ();
 sg13g2_decap_8 FILLER_21_399 ();
 sg13g2_fill_2 FILLER_21_406 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_8 FILLER_22_105 ();
 sg13g2_decap_8 FILLER_22_112 ();
 sg13g2_decap_8 FILLER_22_119 ();
 sg13g2_decap_8 FILLER_22_126 ();
 sg13g2_decap_8 FILLER_22_133 ();
 sg13g2_decap_8 FILLER_22_140 ();
 sg13g2_decap_8 FILLER_22_147 ();
 sg13g2_decap_8 FILLER_22_154 ();
 sg13g2_decap_8 FILLER_22_161 ();
 sg13g2_decap_8 FILLER_22_168 ();
 sg13g2_decap_8 FILLER_22_175 ();
 sg13g2_decap_8 FILLER_22_182 ();
 sg13g2_decap_8 FILLER_22_189 ();
 sg13g2_decap_8 FILLER_22_196 ();
 sg13g2_decap_8 FILLER_22_203 ();
 sg13g2_decap_8 FILLER_22_210 ();
 sg13g2_decap_8 FILLER_22_217 ();
 sg13g2_decap_8 FILLER_22_224 ();
 sg13g2_decap_8 FILLER_22_231 ();
 sg13g2_decap_8 FILLER_22_238 ();
 sg13g2_decap_8 FILLER_22_245 ();
 sg13g2_decap_8 FILLER_22_252 ();
 sg13g2_decap_8 FILLER_22_259 ();
 sg13g2_decap_8 FILLER_22_266 ();
 sg13g2_decap_8 FILLER_22_273 ();
 sg13g2_decap_8 FILLER_22_280 ();
 sg13g2_decap_8 FILLER_22_287 ();
 sg13g2_decap_8 FILLER_22_294 ();
 sg13g2_decap_8 FILLER_22_301 ();
 sg13g2_decap_8 FILLER_22_308 ();
 sg13g2_decap_8 FILLER_22_315 ();
 sg13g2_decap_8 FILLER_22_322 ();
 sg13g2_decap_8 FILLER_22_329 ();
 sg13g2_decap_8 FILLER_22_336 ();
 sg13g2_decap_8 FILLER_22_343 ();
 sg13g2_decap_8 FILLER_22_350 ();
 sg13g2_decap_8 FILLER_22_357 ();
 sg13g2_decap_8 FILLER_22_364 ();
 sg13g2_decap_8 FILLER_22_371 ();
 sg13g2_decap_8 FILLER_22_378 ();
 sg13g2_decap_8 FILLER_22_385 ();
 sg13g2_decap_8 FILLER_22_392 ();
 sg13g2_decap_8 FILLER_22_399 ();
 sg13g2_fill_2 FILLER_22_406 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_98 ();
 sg13g2_decap_8 FILLER_23_105 ();
 sg13g2_decap_8 FILLER_23_112 ();
 sg13g2_decap_8 FILLER_23_119 ();
 sg13g2_decap_8 FILLER_23_126 ();
 sg13g2_decap_8 FILLER_23_133 ();
 sg13g2_decap_8 FILLER_23_140 ();
 sg13g2_decap_8 FILLER_23_147 ();
 sg13g2_decap_8 FILLER_23_154 ();
 sg13g2_decap_8 FILLER_23_161 ();
 sg13g2_decap_8 FILLER_23_168 ();
 sg13g2_decap_8 FILLER_23_175 ();
 sg13g2_decap_8 FILLER_23_182 ();
 sg13g2_decap_8 FILLER_23_189 ();
 sg13g2_decap_8 FILLER_23_196 ();
 sg13g2_decap_8 FILLER_23_203 ();
 sg13g2_decap_8 FILLER_23_210 ();
 sg13g2_decap_8 FILLER_23_217 ();
 sg13g2_decap_8 FILLER_23_224 ();
 sg13g2_decap_8 FILLER_23_231 ();
 sg13g2_decap_8 FILLER_23_238 ();
 sg13g2_decap_8 FILLER_23_245 ();
 sg13g2_fill_2 FILLER_23_252 ();
 sg13g2_fill_1 FILLER_23_254 ();
 sg13g2_decap_8 FILLER_23_264 ();
 sg13g2_decap_8 FILLER_23_271 ();
 sg13g2_decap_8 FILLER_23_278 ();
 sg13g2_decap_8 FILLER_23_285 ();
 sg13g2_decap_8 FILLER_23_292 ();
 sg13g2_decap_8 FILLER_23_299 ();
 sg13g2_decap_8 FILLER_23_306 ();
 sg13g2_decap_8 FILLER_23_313 ();
 sg13g2_decap_8 FILLER_23_320 ();
 sg13g2_decap_8 FILLER_23_327 ();
 sg13g2_decap_8 FILLER_23_334 ();
 sg13g2_decap_8 FILLER_23_341 ();
 sg13g2_decap_8 FILLER_23_348 ();
 sg13g2_decap_8 FILLER_23_355 ();
 sg13g2_decap_8 FILLER_23_362 ();
 sg13g2_decap_8 FILLER_23_369 ();
 sg13g2_decap_8 FILLER_23_376 ();
 sg13g2_decap_8 FILLER_23_383 ();
 sg13g2_decap_8 FILLER_23_390 ();
 sg13g2_decap_8 FILLER_23_397 ();
 sg13g2_decap_4 FILLER_23_404 ();
 sg13g2_fill_1 FILLER_23_408 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_decap_8 FILLER_24_98 ();
 sg13g2_decap_8 FILLER_24_105 ();
 sg13g2_decap_8 FILLER_24_112 ();
 sg13g2_decap_8 FILLER_24_119 ();
 sg13g2_decap_8 FILLER_24_126 ();
 sg13g2_decap_8 FILLER_24_133 ();
 sg13g2_decap_8 FILLER_24_140 ();
 sg13g2_decap_8 FILLER_24_147 ();
 sg13g2_decap_8 FILLER_24_154 ();
 sg13g2_fill_2 FILLER_24_161 ();
 sg13g2_decap_8 FILLER_24_189 ();
 sg13g2_decap_8 FILLER_24_196 ();
 sg13g2_decap_8 FILLER_24_203 ();
 sg13g2_decap_8 FILLER_24_210 ();
 sg13g2_decap_4 FILLER_24_217 ();
 sg13g2_decap_8 FILLER_24_282 ();
 sg13g2_decap_8 FILLER_24_289 ();
 sg13g2_decap_8 FILLER_24_296 ();
 sg13g2_decap_8 FILLER_24_303 ();
 sg13g2_decap_8 FILLER_24_310 ();
 sg13g2_decap_8 FILLER_24_331 ();
 sg13g2_decap_8 FILLER_24_338 ();
 sg13g2_decap_8 FILLER_24_345 ();
 sg13g2_decap_8 FILLER_24_352 ();
 sg13g2_decap_8 FILLER_24_359 ();
 sg13g2_decap_8 FILLER_24_366 ();
 sg13g2_decap_8 FILLER_24_373 ();
 sg13g2_decap_8 FILLER_24_380 ();
 sg13g2_decap_8 FILLER_24_387 ();
 sg13g2_decap_8 FILLER_24_394 ();
 sg13g2_decap_8 FILLER_24_401 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_8 FILLER_25_91 ();
 sg13g2_decap_8 FILLER_25_98 ();
 sg13g2_decap_8 FILLER_25_105 ();
 sg13g2_decap_8 FILLER_25_112 ();
 sg13g2_decap_8 FILLER_25_119 ();
 sg13g2_decap_8 FILLER_25_126 ();
 sg13g2_decap_8 FILLER_25_133 ();
 sg13g2_decap_8 FILLER_25_140 ();
 sg13g2_fill_2 FILLER_25_147 ();
 sg13g2_fill_1 FILLER_25_149 ();
 sg13g2_fill_1 FILLER_25_289 ();
 sg13g2_decap_4 FILLER_25_298 ();
 sg13g2_fill_2 FILLER_25_302 ();
 sg13g2_decap_8 FILLER_25_338 ();
 sg13g2_fill_2 FILLER_25_345 ();
 sg13g2_decap_4 FILLER_25_373 ();
 sg13g2_fill_1 FILLER_25_377 ();
 sg13g2_decap_4 FILLER_25_404 ();
 sg13g2_fill_1 FILLER_25_408 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_decap_8 FILLER_26_91 ();
 sg13g2_decap_8 FILLER_26_98 ();
 sg13g2_decap_8 FILLER_26_105 ();
 sg13g2_decap_8 FILLER_26_112 ();
 sg13g2_decap_8 FILLER_26_119 ();
 sg13g2_decap_8 FILLER_26_126 ();
 sg13g2_decap_8 FILLER_26_133 ();
 sg13g2_decap_8 FILLER_26_140 ();
 sg13g2_decap_8 FILLER_26_147 ();
 sg13g2_fill_2 FILLER_26_154 ();
 sg13g2_fill_1 FILLER_26_156 ();
 sg13g2_decap_4 FILLER_26_209 ();
 sg13g2_fill_2 FILLER_26_213 ();
 sg13g2_fill_2 FILLER_26_290 ();
 sg13g2_decap_4 FILLER_26_301 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_decap_8 FILLER_27_84 ();
 sg13g2_decap_8 FILLER_27_91 ();
 sg13g2_decap_8 FILLER_27_98 ();
 sg13g2_decap_8 FILLER_27_105 ();
 sg13g2_decap_8 FILLER_27_112 ();
 sg13g2_decap_8 FILLER_27_119 ();
 sg13g2_decap_8 FILLER_27_126 ();
 sg13g2_decap_8 FILLER_27_133 ();
 sg13g2_decap_8 FILLER_27_140 ();
 sg13g2_decap_8 FILLER_27_147 ();
 sg13g2_decap_8 FILLER_27_154 ();
 sg13g2_fill_1 FILLER_27_240 ();
 sg13g2_decap_8 FILLER_27_250 ();
 sg13g2_decap_8 FILLER_27_257 ();
 sg13g2_decap_4 FILLER_27_264 ();
 sg13g2_fill_2 FILLER_27_268 ();
 sg13g2_decap_8 FILLER_27_305 ();
 sg13g2_fill_1 FILLER_27_312 ();
 sg13g2_fill_1 FILLER_27_339 ();
 sg13g2_decap_4 FILLER_27_357 ();
 sg13g2_fill_1 FILLER_27_361 ();
 sg13g2_fill_2 FILLER_27_406 ();
 sg13g2_fill_1 FILLER_27_408 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_decap_8 FILLER_28_84 ();
 sg13g2_decap_8 FILLER_28_91 ();
 sg13g2_decap_8 FILLER_28_98 ();
 sg13g2_decap_8 FILLER_28_105 ();
 sg13g2_decap_8 FILLER_28_112 ();
 sg13g2_decap_8 FILLER_28_119 ();
 sg13g2_decap_8 FILLER_28_126 ();
 sg13g2_decap_8 FILLER_28_133 ();
 sg13g2_decap_8 FILLER_28_140 ();
 sg13g2_decap_8 FILLER_28_147 ();
 sg13g2_decap_8 FILLER_28_154 ();
 sg13g2_decap_8 FILLER_28_161 ();
 sg13g2_fill_2 FILLER_28_168 ();
 sg13g2_decap_4 FILLER_28_195 ();
 sg13g2_fill_2 FILLER_28_204 ();
 sg13g2_decap_4 FILLER_28_214 ();
 sg13g2_fill_1 FILLER_28_218 ();
 sg13g2_decap_4 FILLER_28_228 ();
 sg13g2_decap_8 FILLER_28_249 ();
 sg13g2_decap_4 FILLER_28_256 ();
 sg13g2_fill_1 FILLER_28_260 ();
 sg13g2_decap_4 FILLER_28_296 ();
 sg13g2_fill_2 FILLER_28_300 ();
 sg13g2_decap_4 FILLER_28_335 ();
 sg13g2_fill_2 FILLER_28_339 ();
 sg13g2_decap_4 FILLER_28_393 ();
 sg13g2_decap_4 FILLER_28_405 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_decap_8 FILLER_29_84 ();
 sg13g2_decap_8 FILLER_29_91 ();
 sg13g2_decap_8 FILLER_29_98 ();
 sg13g2_decap_8 FILLER_29_105 ();
 sg13g2_decap_8 FILLER_29_112 ();
 sg13g2_decap_8 FILLER_29_119 ();
 sg13g2_decap_8 FILLER_29_126 ();
 sg13g2_decap_8 FILLER_29_133 ();
 sg13g2_decap_8 FILLER_29_140 ();
 sg13g2_decap_8 FILLER_29_147 ();
 sg13g2_decap_8 FILLER_29_154 ();
 sg13g2_fill_2 FILLER_29_165 ();
 sg13g2_fill_1 FILLER_29_167 ();
 sg13g2_decap_8 FILLER_29_191 ();
 sg13g2_decap_8 FILLER_29_198 ();
 sg13g2_fill_2 FILLER_29_205 ();
 sg13g2_fill_1 FILLER_29_228 ();
 sg13g2_fill_1 FILLER_29_255 ();
 sg13g2_decap_8 FILLER_29_297 ();
 sg13g2_decap_8 FILLER_29_304 ();
 sg13g2_fill_2 FILLER_29_320 ();
 sg13g2_fill_1 FILLER_29_330 ();
 sg13g2_fill_2 FILLER_29_357 ();
 sg13g2_decap_8 FILLER_29_397 ();
 sg13g2_decap_4 FILLER_29_404 ();
 sg13g2_fill_1 FILLER_29_408 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_77 ();
 sg13g2_decap_8 FILLER_30_84 ();
 sg13g2_decap_8 FILLER_30_91 ();
 sg13g2_decap_8 FILLER_30_98 ();
 sg13g2_decap_8 FILLER_30_105 ();
 sg13g2_decap_8 FILLER_30_112 ();
 sg13g2_decap_8 FILLER_30_119 ();
 sg13g2_decap_8 FILLER_30_126 ();
 sg13g2_decap_8 FILLER_30_133 ();
 sg13g2_decap_8 FILLER_30_140 ();
 sg13g2_decap_4 FILLER_30_147 ();
 sg13g2_fill_1 FILLER_30_151 ();
 sg13g2_fill_2 FILLER_30_258 ();
 sg13g2_fill_1 FILLER_30_260 ();
 sg13g2_fill_2 FILLER_30_299 ();
 sg13g2_fill_1 FILLER_30_327 ();
 sg13g2_fill_2 FILLER_30_349 ();
 sg13g2_fill_1 FILLER_30_351 ();
 sg13g2_decap_8 FILLER_30_378 ();
 sg13g2_decap_8 FILLER_30_385 ();
 sg13g2_decap_8 FILLER_30_392 ();
 sg13g2_decap_8 FILLER_30_399 ();
 sg13g2_fill_2 FILLER_30_406 ();
 sg13g2_fill_1 FILLER_30_408 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_decap_8 FILLER_31_84 ();
 sg13g2_decap_8 FILLER_31_91 ();
 sg13g2_decap_8 FILLER_31_98 ();
 sg13g2_decap_8 FILLER_31_105 ();
 sg13g2_decap_8 FILLER_31_112 ();
 sg13g2_decap_8 FILLER_31_119 ();
 sg13g2_decap_8 FILLER_31_126 ();
 sg13g2_decap_8 FILLER_31_133 ();
 sg13g2_decap_4 FILLER_31_140 ();
 sg13g2_decap_8 FILLER_31_198 ();
 sg13g2_fill_2 FILLER_31_205 ();
 sg13g2_decap_8 FILLER_31_225 ();
 sg13g2_fill_2 FILLER_31_232 ();
 sg13g2_fill_1 FILLER_31_373 ();
 sg13g2_decap_4 FILLER_31_404 ();
 sg13g2_fill_1 FILLER_31_408 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_8 FILLER_32_84 ();
 sg13g2_decap_8 FILLER_32_91 ();
 sg13g2_decap_8 FILLER_32_98 ();
 sg13g2_decap_8 FILLER_32_105 ();
 sg13g2_decap_8 FILLER_32_112 ();
 sg13g2_decap_8 FILLER_32_119 ();
 sg13g2_decap_8 FILLER_32_126 ();
 sg13g2_fill_2 FILLER_32_133 ();
 sg13g2_fill_2 FILLER_32_177 ();
 sg13g2_decap_8 FILLER_32_188 ();
 sg13g2_decap_8 FILLER_32_195 ();
 sg13g2_decap_4 FILLER_32_202 ();
 sg13g2_fill_2 FILLER_32_232 ();
 sg13g2_fill_1 FILLER_32_234 ();
 sg13g2_fill_2 FILLER_32_256 ();
 sg13g2_fill_1 FILLER_32_258 ();
 sg13g2_fill_2 FILLER_32_267 ();
 sg13g2_fill_2 FILLER_32_278 ();
 sg13g2_fill_1 FILLER_32_280 ();
 sg13g2_decap_4 FILLER_32_291 ();
 sg13g2_fill_1 FILLER_32_304 ();
 sg13g2_fill_2 FILLER_32_339 ();
 sg13g2_fill_1 FILLER_32_341 ();
 sg13g2_fill_2 FILLER_32_372 ();
 sg13g2_decap_4 FILLER_32_404 ();
 sg13g2_fill_1 FILLER_32_408 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_decap_8 FILLER_33_91 ();
 sg13g2_decap_8 FILLER_33_98 ();
 sg13g2_decap_8 FILLER_33_105 ();
 sg13g2_decap_8 FILLER_33_112 ();
 sg13g2_decap_8 FILLER_33_119 ();
 sg13g2_decap_8 FILLER_33_126 ();
 sg13g2_decap_8 FILLER_33_133 ();
 sg13g2_fill_2 FILLER_33_140 ();
 sg13g2_fill_1 FILLER_33_142 ();
 sg13g2_decap_4 FILLER_33_181 ();
 sg13g2_fill_2 FILLER_33_185 ();
 sg13g2_fill_1 FILLER_33_213 ();
 sg13g2_fill_2 FILLER_33_227 ();
 sg13g2_fill_2 FILLER_33_248 ();
 sg13g2_fill_1 FILLER_33_250 ();
 sg13g2_decap_8 FILLER_33_277 ();
 sg13g2_fill_1 FILLER_33_284 ();
 sg13g2_decap_4 FILLER_33_349 ();
 sg13g2_fill_1 FILLER_33_353 ();
 sg13g2_decap_4 FILLER_33_358 ();
 sg13g2_fill_1 FILLER_33_362 ();
 sg13g2_decap_8 FILLER_33_402 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_decap_8 FILLER_34_91 ();
 sg13g2_decap_8 FILLER_34_98 ();
 sg13g2_decap_8 FILLER_34_105 ();
 sg13g2_decap_8 FILLER_34_112 ();
 sg13g2_decap_8 FILLER_34_119 ();
 sg13g2_decap_8 FILLER_34_126 ();
 sg13g2_decap_8 FILLER_34_133 ();
 sg13g2_decap_8 FILLER_34_140 ();
 sg13g2_fill_2 FILLER_34_147 ();
 sg13g2_fill_1 FILLER_34_149 ();
 sg13g2_decap_8 FILLER_34_171 ();
 sg13g2_decap_8 FILLER_34_178 ();
 sg13g2_decap_8 FILLER_34_185 ();
 sg13g2_decap_8 FILLER_34_192 ();
 sg13g2_fill_2 FILLER_34_199 ();
 sg13g2_fill_1 FILLER_34_201 ();
 sg13g2_decap_8 FILLER_34_283 ();
 sg13g2_decap_8 FILLER_34_328 ();
 sg13g2_decap_8 FILLER_34_335 ();
 sg13g2_fill_1 FILLER_34_342 ();
 sg13g2_decap_8 FILLER_34_351 ();
 sg13g2_fill_1 FILLER_34_358 ();
 sg13g2_fill_1 FILLER_34_363 ();
 sg13g2_fill_1 FILLER_34_369 ();
 sg13g2_fill_2 FILLER_34_375 ();
 sg13g2_decap_4 FILLER_34_403 ();
 sg13g2_fill_2 FILLER_34_407 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_decap_8 FILLER_35_98 ();
 sg13g2_decap_8 FILLER_35_105 ();
 sg13g2_decap_8 FILLER_35_112 ();
 sg13g2_decap_8 FILLER_35_119 ();
 sg13g2_decap_8 FILLER_35_126 ();
 sg13g2_decap_8 FILLER_35_133 ();
 sg13g2_decap_8 FILLER_35_140 ();
 sg13g2_decap_8 FILLER_35_147 ();
 sg13g2_decap_8 FILLER_35_154 ();
 sg13g2_decap_8 FILLER_35_161 ();
 sg13g2_decap_8 FILLER_35_168 ();
 sg13g2_decap_8 FILLER_35_175 ();
 sg13g2_decap_8 FILLER_35_182 ();
 sg13g2_decap_8 FILLER_35_189 ();
 sg13g2_decap_8 FILLER_35_196 ();
 sg13g2_decap_8 FILLER_35_279 ();
 sg13g2_decap_8 FILLER_35_286 ();
 sg13g2_fill_2 FILLER_35_293 ();
 sg13g2_fill_1 FILLER_35_295 ();
 sg13g2_fill_2 FILLER_35_300 ();
 sg13g2_fill_2 FILLER_35_340 ();
 sg13g2_fill_2 FILLER_35_357 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_decap_8 FILLER_36_112 ();
 sg13g2_decap_8 FILLER_36_119 ();
 sg13g2_decap_8 FILLER_36_126 ();
 sg13g2_decap_8 FILLER_36_133 ();
 sg13g2_decap_8 FILLER_36_140 ();
 sg13g2_decap_8 FILLER_36_147 ();
 sg13g2_decap_8 FILLER_36_154 ();
 sg13g2_decap_8 FILLER_36_161 ();
 sg13g2_decap_8 FILLER_36_168 ();
 sg13g2_decap_8 FILLER_36_175 ();
 sg13g2_decap_8 FILLER_36_182 ();
 sg13g2_decap_8 FILLER_36_189 ();
 sg13g2_decap_8 FILLER_36_196 ();
 sg13g2_decap_8 FILLER_36_203 ();
 sg13g2_fill_1 FILLER_36_210 ();
 sg13g2_decap_4 FILLER_36_265 ();
 sg13g2_fill_1 FILLER_36_269 ();
 sg13g2_decap_8 FILLER_36_278 ();
 sg13g2_decap_8 FILLER_36_285 ();
 sg13g2_decap_4 FILLER_36_404 ();
 sg13g2_fill_1 FILLER_36_408 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_8 FILLER_37_112 ();
 sg13g2_decap_8 FILLER_37_119 ();
 sg13g2_decap_8 FILLER_37_126 ();
 sg13g2_decap_8 FILLER_37_133 ();
 sg13g2_decap_8 FILLER_37_140 ();
 sg13g2_decap_8 FILLER_37_147 ();
 sg13g2_decap_8 FILLER_37_154 ();
 sg13g2_decap_8 FILLER_37_161 ();
 sg13g2_decap_8 FILLER_37_168 ();
 sg13g2_decap_8 FILLER_37_175 ();
 sg13g2_decap_8 FILLER_37_182 ();
 sg13g2_decap_8 FILLER_37_189 ();
 sg13g2_decap_8 FILLER_37_196 ();
 sg13g2_decap_8 FILLER_37_203 ();
 sg13g2_decap_8 FILLER_37_210 ();
 sg13g2_fill_1 FILLER_37_217 ();
 sg13g2_fill_1 FILLER_37_237 ();
 sg13g2_decap_8 FILLER_37_290 ();
 sg13g2_fill_2 FILLER_37_297 ();
 sg13g2_fill_1 FILLER_37_299 ();
 sg13g2_fill_2 FILLER_37_342 ();
 sg13g2_fill_2 FILLER_37_361 ();
 sg13g2_decap_4 FILLER_37_403 ();
 sg13g2_fill_2 FILLER_37_407 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_4 FILLER_38_60 ();
 sg13g2_decap_4 FILLER_38_68 ();
 sg13g2_decap_4 FILLER_38_76 ();
 sg13g2_decap_4 FILLER_38_84 ();
 sg13g2_decap_4 FILLER_38_92 ();
 sg13g2_decap_4 FILLER_38_100 ();
 sg13g2_decap_4 FILLER_38_108 ();
 sg13g2_decap_8 FILLER_38_116 ();
 sg13g2_decap_8 FILLER_38_123 ();
 sg13g2_decap_8 FILLER_38_130 ();
 sg13g2_decap_8 FILLER_38_137 ();
 sg13g2_decap_8 FILLER_38_144 ();
 sg13g2_decap_8 FILLER_38_151 ();
 sg13g2_decap_8 FILLER_38_158 ();
 sg13g2_decap_8 FILLER_38_165 ();
 sg13g2_decap_8 FILLER_38_172 ();
 sg13g2_decap_8 FILLER_38_179 ();
 sg13g2_decap_8 FILLER_38_186 ();
 sg13g2_decap_8 FILLER_38_193 ();
 sg13g2_decap_8 FILLER_38_200 ();
 sg13g2_decap_8 FILLER_38_207 ();
 sg13g2_decap_8 FILLER_38_214 ();
 sg13g2_decap_4 FILLER_38_221 ();
 sg13g2_fill_2 FILLER_38_225 ();
 sg13g2_decap_8 FILLER_38_236 ();
 sg13g2_fill_2 FILLER_38_243 ();
 sg13g2_fill_2 FILLER_38_257 ();
 sg13g2_fill_1 FILLER_38_259 ();
 sg13g2_decap_8 FILLER_38_286 ();
 sg13g2_decap_8 FILLER_38_293 ();
 sg13g2_decap_8 FILLER_38_300 ();
 sg13g2_decap_4 FILLER_38_307 ();
 sg13g2_fill_1 FILLER_38_311 ();
 sg13g2_decap_8 FILLER_38_321 ();
 sg13g2_fill_2 FILLER_38_341 ();
 sg13g2_fill_1 FILLER_38_343 ();
 sg13g2_fill_2 FILLER_38_349 ();
 sg13g2_fill_1 FILLER_38_351 ();
 sg13g2_decap_4 FILLER_38_356 ();
 sg13g2_decap_4 FILLER_38_364 ();
 sg13g2_fill_1 FILLER_38_368 ();
 sg13g2_fill_2 FILLER_38_385 ();
 sg13g2_decap_8 FILLER_38_395 ();
 sg13g2_decap_8 FILLER_38_402 ();
 assign uio_oe[0] = net15;
 assign uio_oe[1] = net16;
 assign uio_oe[2] = net17;
 assign uio_oe[3] = net18;
 assign uio_oe[4] = net19;
 assign uio_oe[5] = net20;
 assign uio_oe[6] = net21;
 assign uio_oe[7] = net22;
endmodule

module tt_um_jun1okamura_test0 (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire net4;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire clk2;
 wire clk2d;
 wire \counter[0] ;
 wire \counter[10] ;
 wire \counter[11] ;
 wire \counter[12] ;
 wire \counter[13] ;
 wire \counter[14] ;
 wire \counter[15] ;
 wire \counter[1] ;
 wire \counter[2] ;
 wire \counter[3] ;
 wire \counter[4] ;
 wire \counter[5] ;
 wire \counter[6] ;
 wire \counter[7] ;
 wire \counter[8] ;
 wire \counter[9] ;
 wire \data[0] ;
 wire \data[1] ;
 wire \data[2] ;
 wire \data[3] ;
 wire \lfsr_mod.data.lfsr_out[0] ;
 wire \lfsr_mod.data.lfsr_out[10] ;
 wire \lfsr_mod.data.lfsr_out[11] ;
 wire \lfsr_mod.data.lfsr_out[12] ;
 wire \lfsr_mod.data.lfsr_out[13] ;
 wire \lfsr_mod.data.lfsr_out[14] ;
 wire \lfsr_mod.data.lfsr_out[15] ;
 wire \lfsr_mod.data.lfsr_out[1] ;
 wire \lfsr_mod.data.lfsr_out[2] ;
 wire \lfsr_mod.data.lfsr_out[3] ;
 wire \lfsr_mod.data.lfsr_out[4] ;
 wire \lfsr_mod.data.lfsr_out[5] ;
 wire \lfsr_mod.data.lfsr_out[6] ;
 wire \lfsr_mod.data.lfsr_out[7] ;
 wire \lfsr_mod.data.lfsr_out[8] ;
 wire \lfsr_mod.data.lfsr_out[9] ;
 wire \lfsr_mod.mux1.sel8[0] ;
 wire \lfsr_mod.mux1.sel8[1] ;
 wire \lfsr_mod.mux1.sel8[2] ;
 wire \lfsr_mod.mux1.sel8[3] ;
 wire \lfsr_mod.mux1.sel8[4] ;
 wire \lfsr_mod.mux1.sel8[5] ;
 wire \lfsr_mod.mux1.sel8[6] ;
 wire \lfsr_mod.mux1.sel8[7] ;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire clknet_0_clk;
 wire net3;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net1;
 wire net2;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net104;
 wire net105;

 sg13g2_inv_1 _235_ (.Y(_057_),
    .A(\counter[8] ));
 sg13g2_inv_1 _236_ (.Y(_058_),
    .A(\counter[9] ));
 sg13g2_inv_1 _237_ (.Y(_059_),
    .A(net14));
 sg13g2_inv_2 _238_ (.Y(_060_),
    .A(net92));
 sg13g2_inv_1 _239_ (.Y(_061_),
    .A(net91));
 sg13g2_inv_2 _240_ (.Y(_062_),
    .A(net89));
 sg13g2_inv_1 _241_ (.Y(_063_),
    .A(net95));
 sg13g2_mux2_2 _242_ (.A0(\lfsr_mod.data.lfsr_out[8] ),
    .A1(\lfsr_mod.data.lfsr_out[9] ),
    .S(\lfsr_mod.mux1.sel8[4] ),
    .X(uio_out[4]));
 sg13g2_o21ai_1 _243_ (.B1(_058_),
    .Y(_064_),
    .A1(_063_),
    .A2(uio_out[4]));
 sg13g2_mux2_2 _244_ (.A0(\lfsr_mod.data.lfsr_out[6] ),
    .A1(\lfsr_mod.data.lfsr_out[7] ),
    .S(\lfsr_mod.mux1.sel8[3] ),
    .X(uio_out[3]));
 sg13g2_o21ai_1 _245_ (.B1(_057_),
    .Y(_065_),
    .A1(_063_),
    .A2(uio_out[3]));
 sg13g2_nand2_1 _246_ (.Y(_066_),
    .A(_064_),
    .B(_065_));
 sg13g2_nand3b_1 _247_ (.B(net95),
    .C(\counter[9] ),
    .Y(_067_),
    .A_N(uio_out[4]));
 sg13g2_nand3b_1 _248_ (.B(net95),
    .C(\counter[8] ),
    .Y(_068_),
    .A_N(uio_out[3]));
 sg13g2_and4_1 _249_ (.A(_064_),
    .B(_065_),
    .C(_067_),
    .D(_068_),
    .X(_069_));
 sg13g2_mux2_2 _250_ (.A0(\lfsr_mod.data.lfsr_out[14] ),
    .A1(\lfsr_mod.data.lfsr_out[15] ),
    .S(\lfsr_mod.mux1.sel8[7] ),
    .X(uio_out[7]));
 sg13g2_and3_1 _251_ (.X(_070_),
    .A(net95),
    .B(_025_),
    .C(uio_out[7]));
 sg13g2_a21oi_1 _252_ (.A1(net95),
    .A2(uio_out[7]),
    .Y(_071_),
    .B1(_025_));
 sg13g2_nor2_1 _253_ (.A(\counter[14] ),
    .B(\counter[15] ),
    .Y(_072_));
 sg13g2_or2_1 _254_ (.X(_073_),
    .B(\counter[15] ),
    .A(\counter[14] ));
 sg13g2_nor4_2 _255_ (.A(_026_),
    .B(_070_),
    .C(_071_),
    .Y(_074_),
    .D(_073_));
 sg13g2_mux2_2 _256_ (.A0(\lfsr_mod.data.lfsr_out[12] ),
    .A1(\lfsr_mod.data.lfsr_out[13] ),
    .S(\lfsr_mod.mux1.sel8[6] ),
    .X(uio_out[6]));
 sg13g2_a21o_1 _257_ (.A2(uio_out[6]),
    .A1(net95),
    .B1(_024_),
    .X(_075_));
 sg13g2_nand3_1 _258_ (.B(net95),
    .C(uio_out[6]),
    .A(_024_),
    .Y(_076_));
 sg13g2_mux2_2 _259_ (.A0(\lfsr_mod.data.lfsr_out[10] ),
    .A1(\lfsr_mod.data.lfsr_out[11] ),
    .S(\lfsr_mod.mux1.sel8[5] ),
    .X(uio_out[5]));
 sg13g2_nor2_1 _260_ (.A(_063_),
    .B(uio_out[5]),
    .Y(_077_));
 sg13g2_or3_1 _261_ (.A(_023_),
    .B(_063_),
    .C(uio_out[5]),
    .X(_078_));
 sg13g2_o21ai_1 _262_ (.B1(_023_),
    .Y(_079_),
    .A1(_063_),
    .A2(uio_out[5]));
 sg13g2_and4_1 _263_ (.A(_075_),
    .B(_076_),
    .C(_078_),
    .D(_079_),
    .X(_080_));
 sg13g2_nand3_1 _264_ (.B(_074_),
    .C(_080_),
    .A(_069_),
    .Y(_081_));
 sg13g2_mux2_2 _265_ (.A0(\lfsr_mod.data.lfsr_out[4] ),
    .A1(\lfsr_mod.data.lfsr_out[5] ),
    .S(\lfsr_mod.mux1.sel8[2] ),
    .X(uio_out[2]));
 sg13g2_nand2_2 _266_ (.Y(_082_),
    .A(net96),
    .B(uio_out[2]));
 sg13g2_xor2_1 _267_ (.B(_082_),
    .A(_022_),
    .X(_083_));
 sg13g2_xnor2_1 _268_ (.Y(_084_),
    .A(_022_),
    .B(_082_));
 sg13g2_mux2_1 _269_ (.A0(\lfsr_mod.data.lfsr_out[2] ),
    .A1(\lfsr_mod.data.lfsr_out[3] ),
    .S(\lfsr_mod.mux1.sel8[1] ),
    .X(uio_out[1]));
 sg13g2_nand2_1 _270_ (.Y(_085_),
    .A(net95),
    .B(uio_out[1]));
 sg13g2_xor2_1 _271_ (.B(_085_),
    .A(_021_),
    .X(_086_));
 sg13g2_mux2_2 _272_ (.A0(\lfsr_mod.data.lfsr_out[0] ),
    .A1(\lfsr_mod.data.lfsr_out[1] ),
    .S(\lfsr_mod.mux1.sel8[0] ),
    .X(uio_out[0]));
 sg13g2_and2_1 _273_ (.A(net96),
    .B(uio_out[0]),
    .X(_087_));
 sg13g2_nor2_1 _274_ (.A(\counter[4] ),
    .B(net96),
    .Y(_088_));
 sg13g2_o21ai_1 _275_ (.B1(_020_),
    .Y(_089_),
    .A1(_087_),
    .A2(_088_));
 sg13g2_or3_1 _276_ (.A(_083_),
    .B(_086_),
    .C(_089_),
    .X(_090_));
 sg13g2_nor2_1 _277_ (.A(\counter[7] ),
    .B(_082_),
    .Y(_091_));
 sg13g2_nor2_1 _278_ (.A(\counter[6] ),
    .B(_085_),
    .Y(_092_));
 sg13g2_a21oi_1 _279_ (.A1(_084_),
    .A2(_092_),
    .Y(_093_),
    .B1(_091_));
 sg13g2_a21oi_1 _280_ (.A1(_090_),
    .A2(_093_),
    .Y(_094_),
    .B1(_081_));
 sg13g2_nand4_1 _281_ (.B(_067_),
    .C(_074_),
    .A(_066_),
    .Y(_095_),
    .D(_080_));
 sg13g2_o21ai_1 _282_ (.B1(_072_),
    .Y(_096_),
    .A1(_059_),
    .A2(_070_));
 sg13g2_o21ai_1 _283_ (.B1(_076_),
    .Y(_097_),
    .A1(\counter[10] ),
    .A2(_077_));
 sg13g2_nand3_1 _284_ (.B(_075_),
    .C(_097_),
    .A(_074_),
    .Y(_098_));
 sg13g2_nand3_1 _285_ (.B(_096_),
    .C(_098_),
    .A(_095_),
    .Y(_099_));
 sg13g2_or2_1 _286_ (.X(_100_),
    .B(\counter[1] ),
    .A(\counter[0] ));
 sg13g2_nor3_1 _287_ (.A(\counter[2] ),
    .B(\counter[3] ),
    .C(_088_),
    .Y(_101_));
 sg13g2_a221oi_1 _288_ (.B2(_020_),
    .C1(_100_),
    .B1(_087_),
    .A1(\counter[4] ),
    .Y(_102_),
    .A2(net96));
 sg13g2_o21ai_1 _289_ (.B1(_101_),
    .Y(_103_),
    .A1(_020_),
    .A2(_087_));
 sg13g2_nor3_1 _290_ (.A(_083_),
    .B(_086_),
    .C(_103_),
    .Y(_104_));
 sg13g2_nand3b_1 _291_ (.B(_102_),
    .C(_104_),
    .Y(_105_),
    .A_N(_081_));
 sg13g2_o21ai_1 _292_ (.B1(_105_),
    .Y(_106_),
    .A1(_094_),
    .A2(_099_));
 sg13g2_nor2_1 _293_ (.A(net32),
    .B(net80),
    .Y(_000_));
 sg13g2_xnor2_1 _294_ (.Y(_107_),
    .A(net32),
    .B(net66));
 sg13g2_nor2_1 _295_ (.A(net80),
    .B(_107_),
    .Y(_007_));
 sg13g2_and3_1 _296_ (.X(_108_),
    .A(net32),
    .B(net66),
    .C(net25));
 sg13g2_a21oi_1 _297_ (.A1(\counter[0] ),
    .A2(\counter[1] ),
    .Y(_109_),
    .B1(net25));
 sg13g2_nor3_1 _298_ (.A(net80),
    .B(_108_),
    .C(net26),
    .Y(_008_));
 sg13g2_nor2_1 _299_ (.A(net71),
    .B(_108_),
    .Y(_110_));
 sg13g2_and4_1 _300_ (.A(net32),
    .B(net66),
    .C(net25),
    .D(net71),
    .X(_111_));
 sg13g2_nor3_1 _301_ (.A(net80),
    .B(_110_),
    .C(_111_),
    .Y(_009_));
 sg13g2_nor2_1 _302_ (.A(net72),
    .B(_111_),
    .Y(_112_));
 sg13g2_and2_1 _303_ (.A(net72),
    .B(_111_),
    .X(_113_));
 sg13g2_nor3_1 _304_ (.A(net80),
    .B(_112_),
    .C(_113_),
    .Y(_010_));
 sg13g2_xor2_1 _305_ (.B(_113_),
    .A(net69),
    .X(_114_));
 sg13g2_nor2_1 _306_ (.A(net80),
    .B(net70),
    .Y(_011_));
 sg13g2_and3_1 _307_ (.X(_115_),
    .A(\counter[4] ),
    .B(\counter[5] ),
    .C(_111_));
 sg13g2_nand2b_1 _308_ (.Y(_116_),
    .B(_115_),
    .A_N(net58));
 sg13g2_xor2_1 _309_ (.B(_115_),
    .A(net58),
    .X(_117_));
 sg13g2_nor2_1 _310_ (.A(net79),
    .B(net59),
    .Y(_012_));
 sg13g2_xnor2_1 _311_ (.Y(_118_),
    .A(net74),
    .B(_116_));
 sg13g2_nor2_1 _312_ (.A(net80),
    .B(net75),
    .Y(_013_));
 sg13g2_and2_1 _313_ (.A(\counter[7] ),
    .B(\counter[6] ),
    .X(_119_));
 sg13g2_a21oi_1 _314_ (.A1(_115_),
    .A2(_119_),
    .Y(_120_),
    .B1(net33));
 sg13g2_and4_1 _315_ (.A(\counter[7] ),
    .B(\counter[6] ),
    .C(net33),
    .D(_115_),
    .X(_121_));
 sg13g2_nor3_1 _316_ (.A(net79),
    .B(net34),
    .C(_121_),
    .Y(_014_));
 sg13g2_nor2_1 _317_ (.A(net67),
    .B(_121_),
    .Y(_122_));
 sg13g2_and2_1 _318_ (.A(net67),
    .B(_121_),
    .X(_123_));
 sg13g2_nor3_1 _319_ (.A(net79),
    .B(net68),
    .C(_123_),
    .Y(_015_));
 sg13g2_nor2b_1 _320_ (.A(net61),
    .B_N(_123_),
    .Y(_124_));
 sg13g2_nor2b_1 _321_ (.A(_123_),
    .B_N(net61),
    .Y(_125_));
 sg13g2_nor3_1 _322_ (.A(net79),
    .B(_124_),
    .C(net62),
    .Y(_001_));
 sg13g2_xor2_1 _323_ (.B(_124_),
    .A(net47),
    .X(_126_));
 sg13g2_nor2_1 _324_ (.A(net79),
    .B(net48),
    .Y(_002_));
 sg13g2_nand3_1 _325_ (.B(\counter[10] ),
    .C(_123_),
    .A(\counter[11] ),
    .Y(_127_));
 sg13g2_nand4_1 _326_ (.B(\counter[10] ),
    .C(\counter[12] ),
    .A(\counter[11] ),
    .Y(_128_),
    .D(_123_));
 sg13g2_xor2_1 _327_ (.B(_127_),
    .A(net56),
    .X(_129_));
 sg13g2_nor2_1 _328_ (.A(net81),
    .B(net57),
    .Y(_003_));
 sg13g2_xnor2_1 _329_ (.Y(_130_),
    .A(net39),
    .B(_128_));
 sg13g2_nor2_1 _330_ (.A(net79),
    .B(net40),
    .Y(_004_));
 sg13g2_nor3_1 _331_ (.A(_059_),
    .B(net79),
    .C(_128_),
    .Y(_005_));
 sg13g2_nand2_1 _332_ (.Y(_131_),
    .A(\data[0] ),
    .B(\data[1] ));
 sg13g2_a21oi_1 _333_ (.A1(\data[0] ),
    .A2(net91),
    .Y(_132_),
    .B1(net89));
 sg13g2_o21ai_1 _334_ (.B1(net87),
    .Y(_133_),
    .A1(_062_),
    .A2(_018_));
 sg13g2_nor2_2 _335_ (.A(net91),
    .B(_062_),
    .Y(_134_));
 sg13g2_nor2_1 _336_ (.A(net92),
    .B(net86),
    .Y(_135_));
 sg13g2_a21oi_1 _337_ (.A1(_134_),
    .A2(_135_),
    .Y(_136_),
    .B1(net93));
 sg13g2_nor2_2 _338_ (.A(_060_),
    .B(net91),
    .Y(_137_));
 sg13g2_nand2_2 _339_ (.Y(_138_),
    .A(net92),
    .B(_061_));
 sg13g2_nand2_1 _340_ (.Y(_139_),
    .A(net92),
    .B(_062_));
 sg13g2_nor3_1 _341_ (.A(net89),
    .B(net87),
    .C(_138_),
    .Y(_140_));
 sg13g2_o21ai_1 _342_ (.B1(_136_),
    .Y(_141_),
    .A1(_132_),
    .A2(_133_));
 sg13g2_nor2_1 _343_ (.A(_140_),
    .B(_141_),
    .Y(_142_));
 sg13g2_nand2_2 _344_ (.Y(_143_),
    .A(_060_),
    .B(net91));
 sg13g2_o21ai_1 _345_ (.B1(net86),
    .Y(_144_),
    .A1(net89),
    .A2(_143_));
 sg13g2_a21oi_1 _346_ (.A1(_060_),
    .A2(_134_),
    .Y(_145_),
    .B1(_144_));
 sg13g2_nand2_1 _347_ (.Y(_146_),
    .A(net91),
    .B(_135_));
 sg13g2_o21ai_1 _348_ (.B1(net94),
    .Y(_147_),
    .A1(_017_),
    .A2(_146_));
 sg13g2_nor2_1 _349_ (.A(_145_),
    .B(_147_),
    .Y(_148_));
 sg13g2_nor2_1 _350_ (.A(_142_),
    .B(_148_),
    .Y(uo_out[0]));
 sg13g2_nor2_2 _351_ (.A(net90),
    .B(_137_),
    .Y(_149_));
 sg13g2_inv_1 _352_ (.Y(_150_),
    .A(_149_));
 sg13g2_nand2_1 _353_ (.Y(_151_),
    .A(_138_),
    .B(_143_));
 sg13g2_nand2_1 _354_ (.Y(_152_),
    .A(_143_),
    .B(_149_));
 sg13g2_a21oi_1 _355_ (.A1(net92),
    .A2(net89),
    .Y(_153_),
    .B1(net86));
 sg13g2_inv_1 _356_ (.Y(_154_),
    .A(_153_));
 sg13g2_nand2_1 _357_ (.Y(_155_),
    .A(_152_),
    .B(_153_));
 sg13g2_nand2_1 _358_ (.Y(_156_),
    .A(net86),
    .B(_149_));
 sg13g2_nand3_1 _359_ (.B(_155_),
    .C(_156_),
    .A(net94),
    .Y(_157_));
 sg13g2_a21oi_1 _360_ (.A1(net90),
    .A2(_151_),
    .Y(_158_),
    .B1(net88));
 sg13g2_a21oi_1 _361_ (.A1(net86),
    .A2(_137_),
    .Y(_159_),
    .B1(_132_));
 sg13g2_nand2b_1 _362_ (.Y(_160_),
    .B(_159_),
    .A_N(net94));
 sg13g2_o21ai_1 _363_ (.B1(_157_),
    .Y(uo_out[1]),
    .A1(_158_),
    .A2(_160_));
 sg13g2_a21oi_1 _364_ (.A1(_017_),
    .A2(_138_),
    .Y(_161_),
    .B1(net86));
 sg13g2_o21ai_1 _365_ (.B1(net86),
    .Y(_162_),
    .A1(_134_),
    .A2(_149_));
 sg13g2_nand2b_1 _366_ (.Y(_163_),
    .B(_162_),
    .A_N(_161_));
 sg13g2_a21oi_1 _367_ (.A1(_062_),
    .A2(_146_),
    .Y(_164_),
    .B1(_137_));
 sg13g2_nor2_1 _368_ (.A(net94),
    .B(_164_),
    .Y(_165_));
 sg13g2_nor2_1 _369_ (.A(net87),
    .B(net93),
    .Y(_166_));
 sg13g2_a221oi_1 _370_ (.B2(net89),
    .C1(_165_),
    .B1(_166_),
    .A1(net94),
    .Y(uo_out[2]),
    .A2(_163_));
 sg13g2_nand2_1 _371_ (.Y(_167_),
    .A(net90),
    .B(_131_));
 sg13g2_nand3_1 _372_ (.B(_152_),
    .C(_167_),
    .A(_146_),
    .Y(_168_));
 sg13g2_a221oi_1 _373_ (.B2(_060_),
    .C1(net88),
    .B1(_134_),
    .A1(_062_),
    .Y(_169_),
    .A2(_019_));
 sg13g2_a21o_1 _374_ (.A2(_134_),
    .A1(net87),
    .B1(_169_),
    .X(_170_));
 sg13g2_a22oi_1 _375_ (.Y(uo_out[3]),
    .B1(_170_),
    .B2(net93),
    .A2(_168_),
    .A1(_136_));
 sg13g2_nor2_1 _376_ (.A(net92),
    .B(_134_),
    .Y(_171_));
 sg13g2_nor2_1 _377_ (.A(net87),
    .B(_171_),
    .Y(_172_));
 sg13g2_and3_1 _378_ (.X(_173_),
    .A(_062_),
    .B(net88),
    .C(_137_));
 sg13g2_nand3_1 _379_ (.B(_139_),
    .C(_151_),
    .A(net86),
    .Y(_174_));
 sg13g2_nor3_1 _380_ (.A(net92),
    .B(net91),
    .C(net89),
    .Y(_175_));
 sg13g2_o21ai_1 _381_ (.B1(_174_),
    .Y(_176_),
    .A1(_154_),
    .A2(_175_));
 sg13g2_nor3_1 _382_ (.A(net93),
    .B(_172_),
    .C(_173_),
    .Y(_177_));
 sg13g2_a21oi_1 _383_ (.A1(net93),
    .A2(_176_),
    .Y(uo_out[4]),
    .B1(_177_));
 sg13g2_a21oi_1 _384_ (.A1(_060_),
    .A2(_061_),
    .Y(_178_),
    .B1(net87));
 sg13g2_a221oi_1 _385_ (.B2(_178_),
    .C1(net93),
    .B1(_167_),
    .A1(net87),
    .Y(_179_),
    .A2(_134_));
 sg13g2_a21oi_1 _386_ (.A1(net92),
    .A2(net87),
    .Y(_180_),
    .B1(_175_));
 sg13g2_a21oi_1 _387_ (.A1(net93),
    .A2(_180_),
    .Y(uo_out[5]),
    .B1(_179_));
 sg13g2_a21oi_1 _388_ (.A1(_143_),
    .A2(_150_),
    .Y(_181_),
    .B1(_144_));
 sg13g2_o21ai_1 _389_ (.B1(_166_),
    .Y(_182_),
    .A1(net89),
    .A2(_018_));
 sg13g2_nand2b_1 _390_ (.Y(_183_),
    .B(_167_),
    .A_N(_182_));
 sg13g2_o21ai_1 _391_ (.B1(net93),
    .Y(_184_),
    .A1(_140_),
    .A2(_181_));
 sg13g2_nand2_1 _392_ (.Y(uo_out[6]),
    .A(_183_),
    .B(_184_));
 sg13g2_xor2_1 _393_ (.B(clk2d),
    .A(clk2),
    .X(_185_));
 sg13g2_xnor2_1 _394_ (.Y(_186_),
    .A(clk2),
    .B(clk2d));
 sg13g2_nand2_1 _395_ (.Y(_187_),
    .A(net30),
    .B(net83));
 sg13g2_xnor2_1 _396_ (.Y(_188_),
    .A(\lfsr_mod.mux1.sel8[7] ),
    .B(\lfsr_mod.mux1.sel8[5] ));
 sg13g2_xor2_1 _397_ (.B(\lfsr_mod.mux1.sel8[3] ),
    .A(\lfsr_mod.mux1.sel8[4] ),
    .X(_189_));
 sg13g2_xnor2_1 _398_ (.Y(_190_),
    .A(_188_),
    .B(_189_));
 sg13g2_o21ai_1 _399_ (.B1(_187_),
    .Y(_028_),
    .A1(net82),
    .A2(_190_));
 sg13g2_mux2_1 _400_ (.A0(net60),
    .A1(net30),
    .S(net85),
    .X(_029_));
 sg13g2_mux2_1 _401_ (.A0(net45),
    .A1(\lfsr_mod.mux1.sel8[1] ),
    .S(net85),
    .X(_030_));
 sg13g2_mux2_1 _402_ (.A0(net53),
    .A1(net45),
    .S(net84),
    .X(_031_));
 sg13g2_mux2_1 _403_ (.A0(net73),
    .A1(net53),
    .S(net84),
    .X(_032_));
 sg13g2_mux2_1 _404_ (.A0(net63),
    .A1(\lfsr_mod.mux1.sel8[4] ),
    .S(net84),
    .X(_033_));
 sg13g2_mux2_1 _405_ (.A0(net63),
    .A1(net65),
    .S(net82),
    .X(_034_));
 sg13g2_mux2_1 _406_ (.A0(net51),
    .A1(\lfsr_mod.mux1.sel8[6] ),
    .S(net84),
    .X(_035_));
 sg13g2_xnor2_1 _407_ (.Y(_036_),
    .A(_060_),
    .B(net81));
 sg13g2_a21oi_1 _408_ (.A1(_138_),
    .A2(_143_),
    .Y(_191_),
    .B1(_173_));
 sg13g2_mux2_1 _409_ (.A0(net91),
    .A1(_191_),
    .S(net81),
    .X(_037_));
 sg13g2_nor2_1 _410_ (.A(_017_),
    .B(_131_),
    .Y(_192_));
 sg13g2_and2_1 _411_ (.A(_017_),
    .B(_131_),
    .X(_193_));
 sg13g2_nor3_1 _412_ (.A(_173_),
    .B(_192_),
    .C(_193_),
    .Y(_194_));
 sg13g2_mux2_1 _413_ (.A0(net90),
    .A1(_194_),
    .S(net80),
    .X(_038_));
 sg13g2_xor2_1 _414_ (.B(_192_),
    .A(_027_),
    .X(_195_));
 sg13g2_nor2_1 _415_ (.A(_173_),
    .B(_195_),
    .Y(_196_));
 sg13g2_mux2_1 _416_ (.A0(net88),
    .A1(_196_),
    .S(net81),
    .X(_039_));
 sg13g2_mux2_1 _417_ (.A0(net12),
    .A1(net13),
    .S(net79),
    .X(_040_));
 sg13g2_nand2_1 _418_ (.Y(_197_),
    .A(net16),
    .B(net83));
 sg13g2_xnor2_1 _419_ (.Y(_198_),
    .A(\lfsr_mod.data.lfsr_out[15] ),
    .B(\lfsr_mod.data.lfsr_out[14] ));
 sg13g2_xor2_1 _420_ (.B(\lfsr_mod.data.lfsr_out[10] ),
    .A(\lfsr_mod.data.lfsr_out[12] ),
    .X(_199_));
 sg13g2_xnor2_1 _421_ (.Y(_200_),
    .A(_198_),
    .B(_199_));
 sg13g2_o21ai_1 _422_ (.B1(_197_),
    .Y(_041_),
    .A1(net83),
    .A2(_200_));
 sg13g2_mux2_1 _423_ (.A0(net16),
    .A1(net20),
    .S(net83),
    .X(_042_));
 sg13g2_mux2_1 _424_ (.A0(net18),
    .A1(net20),
    .S(net85),
    .X(_043_));
 sg13g2_mux2_1 _425_ (.A0(net18),
    .A1(\lfsr_mod.data.lfsr_out[3] ),
    .S(net83),
    .X(_044_));
 sg13g2_mux2_1 _426_ (.A0(net21),
    .A1(net29),
    .S(net84),
    .X(_045_));
 sg13g2_mux2_1 _427_ (.A0(net21),
    .A1(\lfsr_mod.data.lfsr_out[5] ),
    .S(net82),
    .X(_046_));
 sg13g2_mux2_1 _428_ (.A0(net38),
    .A1(net36),
    .S(net82),
    .X(_047_));
 sg13g2_mux2_1 _429_ (.A0(net36),
    .A1(\lfsr_mod.data.lfsr_out[7] ),
    .S(net82),
    .X(_048_));
 sg13g2_mux2_1 _430_ (.A0(net23),
    .A1(\lfsr_mod.data.lfsr_out[7] ),
    .S(net84),
    .X(_049_));
 sg13g2_mux2_1 _431_ (.A0(net23),
    .A1(net28),
    .S(net82),
    .X(_050_));
 sg13g2_mux2_1 _432_ (.A0(net41),
    .A1(net28),
    .S(net84),
    .X(_051_));
 sg13g2_mux2_1 _433_ (.A0(net41),
    .A1(net42),
    .S(net82),
    .X(_052_));
 sg13g2_mux2_1 _434_ (.A0(net43),
    .A1(net42),
    .S(net84),
    .X(_053_));
 sg13g2_mux2_1 _435_ (.A0(net43),
    .A1(\lfsr_mod.data.lfsr_out[13] ),
    .S(net82),
    .X(_054_));
 sg13g2_mux2_1 _436_ (.A0(\lfsr_mod.data.lfsr_out[14] ),
    .A1(net49),
    .S(net85),
    .X(_055_));
 sg13g2_mux2_1 _437_ (.A0(net54),
    .A1(\lfsr_mod.data.lfsr_out[14] ),
    .S(net85),
    .X(_056_));
 sg13g2_dfrbp_1 _438_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net102),
    .D(_000_),
    .Q_N(_227_),
    .Q(\counter[0] ));
 sg13g2_dfrbp_1 _439_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net102),
    .D(_007_),
    .Q_N(_228_),
    .Q(\counter[1] ));
 sg13g2_dfrbp_1 _440_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net102),
    .D(net27),
    .Q_N(_229_),
    .Q(\counter[2] ));
 sg13g2_dfrbp_1 _441_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net102),
    .D(_009_),
    .Q_N(_230_),
    .Q(\counter[3] ));
 sg13g2_dfrbp_1 _442_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net102),
    .D(_010_),
    .Q_N(_231_),
    .Q(\counter[4] ));
 sg13g2_dfrbp_1 _443_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net102),
    .D(_011_),
    .Q_N(_020_),
    .Q(\counter[5] ));
 sg13g2_dfrbp_1 _444_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net103),
    .D(_012_),
    .Q_N(_021_),
    .Q(\counter[6] ));
 sg13g2_dfrbp_1 _445_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net103),
    .D(_013_),
    .Q_N(_022_),
    .Q(\counter[7] ));
 sg13g2_dfrbp_1 _446_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net103),
    .D(net35),
    .Q_N(_232_),
    .Q(\counter[8] ));
 sg13g2_dfrbp_1 _447_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net103),
    .D(_015_),
    .Q_N(_233_),
    .Q(\counter[9] ));
 sg13g2_dfrbp_1 _448_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net99),
    .D(_001_),
    .Q_N(_023_),
    .Q(\counter[10] ));
 sg13g2_dfrbp_1 _449_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net99),
    .D(_002_),
    .Q_N(_024_),
    .Q(\counter[11] ));
 sg13g2_dfrbp_1 _450_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net99),
    .D(_003_),
    .Q_N(_025_),
    .Q(\counter[12] ));
 sg13g2_dfrbp_1 _451_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net99),
    .D(_004_),
    .Q_N(_026_),
    .Q(\counter[13] ));
 sg13g2_dfrbp_1 _452_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net103),
    .D(net15),
    .Q_N(_234_),
    .Q(\counter[14] ));
 sg13g2_dfrbp_1 _453_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net103),
    .D(net3),
    .Q_N(_226_),
    .Q(\counter[15] ));
 sg13g2_dfrbp_1 _454_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net101),
    .D(net31),
    .Q_N(_225_),
    .Q(\lfsr_mod.mux1.sel8[0] ));
 sg13g2_dfrbp_1 _455_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net100),
    .D(_029_),
    .Q_N(_224_),
    .Q(\lfsr_mod.mux1.sel8[1] ));
 sg13g2_dfrbp_1 _456_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net97),
    .D(net46),
    .Q_N(_223_),
    .Q(\lfsr_mod.mux1.sel8[2] ));
 sg13g2_dfrbp_1 _457_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net97),
    .D(_031_),
    .Q_N(_222_),
    .Q(\lfsr_mod.mux1.sel8[3] ));
 sg13g2_dfrbp_1 _458_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net97),
    .D(_032_),
    .Q_N(_221_),
    .Q(\lfsr_mod.mux1.sel8[4] ));
 sg13g2_dfrbp_1 _459_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net98),
    .D(net64),
    .Q_N(_220_),
    .Q(\lfsr_mod.mux1.sel8[5] ));
 sg13g2_dfrbp_1 _460_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net98),
    .D(_034_),
    .Q_N(_219_),
    .Q(\lfsr_mod.mux1.sel8[6] ));
 sg13g2_dfrbp_1 _461_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net98),
    .D(net52),
    .Q_N(_218_),
    .Q(\lfsr_mod.mux1.sel8[7] ));
 sg13g2_dfrbp_1 _462_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net1),
    .D(_036_),
    .Q_N(_019_),
    .Q(\data[0] ));
 sg13g2_dfrbp_1 _463_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net103),
    .D(_037_),
    .Q_N(_018_),
    .Q(\data[1] ));
 sg13g2_dfrbp_1 _464_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net102),
    .D(net104),
    .Q_N(_017_),
    .Q(\data[2] ));
 sg13g2_dfrbp_1 _465_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net102),
    .D(net77),
    .Q_N(_027_),
    .Q(\data[3] ));
 sg13g2_dfrbp_1 _466_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net99),
    .D(net12),
    .Q_N(_217_),
    .Q(clk2d));
 sg13g2_dfrbp_1 _467_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net99),
    .D(_040_),
    .Q_N(_016_),
    .Q(clk2));
 sg13g2_dfrbp_1 _468_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net100),
    .D(net17),
    .Q_N(_216_),
    .Q(\lfsr_mod.data.lfsr_out[0] ));
 sg13g2_dfrbp_1 _469_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net100),
    .D(_042_),
    .Q_N(_215_),
    .Q(\lfsr_mod.data.lfsr_out[1] ));
 sg13g2_dfrbp_1 _470_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net100),
    .D(_043_),
    .Q_N(_214_),
    .Q(\lfsr_mod.data.lfsr_out[2] ));
 sg13g2_dfrbp_1 _471_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net99),
    .D(net19),
    .Q_N(_213_),
    .Q(\lfsr_mod.data.lfsr_out[3] ));
 sg13g2_dfrbp_1 _472_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net100),
    .D(_045_),
    .Q_N(_212_),
    .Q(\lfsr_mod.data.lfsr_out[4] ));
 sg13g2_dfrbp_1 _473_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net97),
    .D(net22),
    .Q_N(_211_),
    .Q(\lfsr_mod.data.lfsr_out[5] ));
 sg13g2_dfrbp_1 _474_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net97),
    .D(_047_),
    .Q_N(_210_),
    .Q(\lfsr_mod.data.lfsr_out[6] ));
 sg13g2_dfrbp_1 _475_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net97),
    .D(net37),
    .Q_N(_209_),
    .Q(\lfsr_mod.data.lfsr_out[7] ));
 sg13g2_dfrbp_1 _476_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net97),
    .D(net24),
    .Q_N(_208_),
    .Q(\lfsr_mod.data.lfsr_out[8] ));
 sg13g2_dfrbp_1 _477_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net97),
    .D(_050_),
    .Q_N(_207_),
    .Q(\lfsr_mod.data.lfsr_out[9] ));
 sg13g2_dfrbp_1 _478_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net98),
    .D(_051_),
    .Q_N(_206_),
    .Q(\lfsr_mod.data.lfsr_out[10] ));
 sg13g2_dfrbp_1 _479_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net98),
    .D(_052_),
    .Q_N(_205_),
    .Q(\lfsr_mod.data.lfsr_out[11] ));
 sg13g2_dfrbp_1 _480_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net98),
    .D(_053_),
    .Q_N(_204_),
    .Q(\lfsr_mod.data.lfsr_out[12] ));
 sg13g2_dfrbp_1 _481_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net98),
    .D(net44),
    .Q_N(_203_),
    .Q(\lfsr_mod.data.lfsr_out[13] ));
 sg13g2_dfrbp_1 _482_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net98),
    .D(net50),
    .Q_N(_202_),
    .Q(\lfsr_mod.data.lfsr_out[14] ));
 sg13g2_dfrbp_1 _483_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net99),
    .D(net55),
    .Q_N(_201_),
    .Q(\lfsr_mod.data.lfsr_out[15] ));
 sg13g2_tiehi tt_um_jun1okamura_test0_5 (.L_HI(net5));
 sg13g2_tiehi tt_um_jun1okamura_test0_6 (.L_HI(net6));
 sg13g2_tiehi tt_um_jun1okamura_test0_7 (.L_HI(net7));
 sg13g2_tiehi tt_um_jun1okamura_test0_8 (.L_HI(net8));
 sg13g2_tiehi tt_um_jun1okamura_test0_9 (.L_HI(net9));
 sg13g2_tiehi tt_um_jun1okamura_test0_10 (.L_HI(net10));
 sg13g2_tiehi tt_um_jun1okamura_test0_11 (.L_HI(net11));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo _453__3 (.L_LO(net3));
 sg13g2_tiehi tt_um_jun1okamura_test0_4 (.L_HI(net4));
 sg13g2_buf_2 fanout79 (.A(net81),
    .X(net79));
 sg13g2_buf_2 fanout80 (.A(net81),
    .X(net80));
 sg13g2_buf_2 fanout81 (.A(_106_),
    .X(net81));
 sg13g2_buf_4 fanout82 (.X(net82),
    .A(_186_));
 sg13g2_buf_2 fanout83 (.A(_186_),
    .X(net83));
 sg13g2_buf_4 fanout84 (.X(net84),
    .A(_185_));
 sg13g2_buf_2 fanout85 (.A(_185_),
    .X(net85));
 sg13g2_buf_2 fanout86 (.A(net88),
    .X(net86));
 sg13g2_buf_2 fanout87 (.A(net88),
    .X(net87));
 sg13g2_buf_2 fanout88 (.A(net76),
    .X(net88));
 sg13g2_buf_2 fanout89 (.A(\data[2] ),
    .X(net89));
 sg13g2_buf_1 fanout90 (.A(net78),
    .X(net90));
 sg13g2_buf_2 fanout91 (.A(net105),
    .X(net91));
 sg13g2_buf_2 fanout92 (.A(\data[0] ),
    .X(net92));
 sg13g2_buf_2 fanout93 (.A(net94),
    .X(net93));
 sg13g2_buf_2 fanout94 (.A(ui_in[1]),
    .X(net94));
 sg13g2_buf_2 fanout95 (.A(net96),
    .X(net95));
 sg13g2_buf_2 fanout96 (.A(ui_in[0]),
    .X(net96));
 sg13g2_buf_4 fanout97 (.X(net97),
    .A(net101));
 sg13g2_buf_4 fanout98 (.X(net98),
    .A(net101));
 sg13g2_buf_4 fanout99 (.X(net99),
    .A(net101));
 sg13g2_buf_2 fanout100 (.A(net101),
    .X(net100));
 sg13g2_buf_2 fanout101 (.A(net1),
    .X(net101));
 sg13g2_buf_4 fanout102 (.X(net102),
    .A(net103));
 sg13g2_buf_4 fanout103 (.X(net103),
    .A(net1));
 sg13g2_buf_2 input1 (.A(rst_n),
    .X(net1));
 sg13g2_tielo tt_um_jun1okamura_test0_2 (.L_LO(net2));
 sg13g2_buf_2 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sg13g2_buf_2 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sg13g2_buf_2 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sg13g2_buf_2 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sg13g2_buf_2 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sg13g2_buf_2 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sg13g2_buf_2 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sg13g2_buf_2 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_3_3__leaf_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_3_7__leaf_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(clk2),
    .X(net12));
 sg13g2_dlygate4sd3_1 hold2 (.A(_016_),
    .X(net13));
 sg13g2_dlygate4sd3_1 hold3 (.A(\counter[13] ),
    .X(net14));
 sg13g2_dlygate4sd3_1 hold4 (.A(_005_),
    .X(net15));
 sg13g2_dlygate4sd3_1 hold5 (.A(\lfsr_mod.data.lfsr_out[0] ),
    .X(net16));
 sg13g2_dlygate4sd3_1 hold6 (.A(_041_),
    .X(net17));
 sg13g2_dlygate4sd3_1 hold7 (.A(\lfsr_mod.data.lfsr_out[2] ),
    .X(net18));
 sg13g2_dlygate4sd3_1 hold8 (.A(_044_),
    .X(net19));
 sg13g2_dlygate4sd3_1 hold9 (.A(\lfsr_mod.data.lfsr_out[1] ),
    .X(net20));
 sg13g2_dlygate4sd3_1 hold10 (.A(\lfsr_mod.data.lfsr_out[4] ),
    .X(net21));
 sg13g2_dlygate4sd3_1 hold11 (.A(_046_),
    .X(net22));
 sg13g2_dlygate4sd3_1 hold12 (.A(\lfsr_mod.data.lfsr_out[8] ),
    .X(net23));
 sg13g2_dlygate4sd3_1 hold13 (.A(_049_),
    .X(net24));
 sg13g2_dlygate4sd3_1 hold14 (.A(\counter[2] ),
    .X(net25));
 sg13g2_dlygate4sd3_1 hold15 (.A(_109_),
    .X(net26));
 sg13g2_dlygate4sd3_1 hold16 (.A(_008_),
    .X(net27));
 sg13g2_dlygate4sd3_1 hold17 (.A(\lfsr_mod.data.lfsr_out[9] ),
    .X(net28));
 sg13g2_dlygate4sd3_1 hold18 (.A(\lfsr_mod.data.lfsr_out[3] ),
    .X(net29));
 sg13g2_dlygate4sd3_1 hold19 (.A(\lfsr_mod.mux1.sel8[0] ),
    .X(net30));
 sg13g2_dlygate4sd3_1 hold20 (.A(_028_),
    .X(net31));
 sg13g2_dlygate4sd3_1 hold21 (.A(\counter[0] ),
    .X(net32));
 sg13g2_dlygate4sd3_1 hold22 (.A(\counter[8] ),
    .X(net33));
 sg13g2_dlygate4sd3_1 hold23 (.A(_120_),
    .X(net34));
 sg13g2_dlygate4sd3_1 hold24 (.A(_014_),
    .X(net35));
 sg13g2_dlygate4sd3_1 hold25 (.A(\lfsr_mod.data.lfsr_out[6] ),
    .X(net36));
 sg13g2_dlygate4sd3_1 hold26 (.A(_048_),
    .X(net37));
 sg13g2_dlygate4sd3_1 hold27 (.A(\lfsr_mod.data.lfsr_out[5] ),
    .X(net38));
 sg13g2_dlygate4sd3_1 hold28 (.A(_026_),
    .X(net39));
 sg13g2_dlygate4sd3_1 hold29 (.A(_130_),
    .X(net40));
 sg13g2_dlygate4sd3_1 hold30 (.A(\lfsr_mod.data.lfsr_out[10] ),
    .X(net41));
 sg13g2_dlygate4sd3_1 hold31 (.A(\lfsr_mod.data.lfsr_out[11] ),
    .X(net42));
 sg13g2_dlygate4sd3_1 hold32 (.A(\lfsr_mod.data.lfsr_out[12] ),
    .X(net43));
 sg13g2_dlygate4sd3_1 hold33 (.A(_054_),
    .X(net44));
 sg13g2_dlygate4sd3_1 hold34 (.A(\lfsr_mod.mux1.sel8[2] ),
    .X(net45));
 sg13g2_dlygate4sd3_1 hold35 (.A(_030_),
    .X(net46));
 sg13g2_dlygate4sd3_1 hold36 (.A(_024_),
    .X(net47));
 sg13g2_dlygate4sd3_1 hold37 (.A(_126_),
    .X(net48));
 sg13g2_dlygate4sd3_1 hold38 (.A(\lfsr_mod.data.lfsr_out[13] ),
    .X(net49));
 sg13g2_dlygate4sd3_1 hold39 (.A(_055_),
    .X(net50));
 sg13g2_dlygate4sd3_1 hold40 (.A(\lfsr_mod.mux1.sel8[7] ),
    .X(net51));
 sg13g2_dlygate4sd3_1 hold41 (.A(_035_),
    .X(net52));
 sg13g2_dlygate4sd3_1 hold42 (.A(\lfsr_mod.mux1.sel8[3] ),
    .X(net53));
 sg13g2_dlygate4sd3_1 hold43 (.A(\lfsr_mod.data.lfsr_out[15] ),
    .X(net54));
 sg13g2_dlygate4sd3_1 hold44 (.A(_056_),
    .X(net55));
 sg13g2_dlygate4sd3_1 hold45 (.A(\counter[12] ),
    .X(net56));
 sg13g2_dlygate4sd3_1 hold46 (.A(_129_),
    .X(net57));
 sg13g2_dlygate4sd3_1 hold47 (.A(_021_),
    .X(net58));
 sg13g2_dlygate4sd3_1 hold48 (.A(_117_),
    .X(net59));
 sg13g2_dlygate4sd3_1 hold49 (.A(\lfsr_mod.mux1.sel8[1] ),
    .X(net60));
 sg13g2_dlygate4sd3_1 hold50 (.A(_023_),
    .X(net61));
 sg13g2_dlygate4sd3_1 hold51 (.A(_125_),
    .X(net62));
 sg13g2_dlygate4sd3_1 hold52 (.A(\lfsr_mod.mux1.sel8[5] ),
    .X(net63));
 sg13g2_dlygate4sd3_1 hold53 (.A(_033_),
    .X(net64));
 sg13g2_dlygate4sd3_1 hold54 (.A(\lfsr_mod.mux1.sel8[6] ),
    .X(net65));
 sg13g2_dlygate4sd3_1 hold55 (.A(\counter[1] ),
    .X(net66));
 sg13g2_dlygate4sd3_1 hold56 (.A(\counter[9] ),
    .X(net67));
 sg13g2_dlygate4sd3_1 hold57 (.A(_122_),
    .X(net68));
 sg13g2_dlygate4sd3_1 hold58 (.A(_020_),
    .X(net69));
 sg13g2_dlygate4sd3_1 hold59 (.A(_114_),
    .X(net70));
 sg13g2_dlygate4sd3_1 hold60 (.A(\counter[3] ),
    .X(net71));
 sg13g2_dlygate4sd3_1 hold61 (.A(\counter[4] ),
    .X(net72));
 sg13g2_dlygate4sd3_1 hold62 (.A(\lfsr_mod.mux1.sel8[4] ),
    .X(net73));
 sg13g2_dlygate4sd3_1 hold63 (.A(_022_),
    .X(net74));
 sg13g2_dlygate4sd3_1 hold64 (.A(_118_),
    .X(net75));
 sg13g2_dlygate4sd3_1 hold65 (.A(\data[3] ),
    .X(net76));
 sg13g2_dlygate4sd3_1 hold66 (.A(_039_),
    .X(net77));
 sg13g2_dlygate4sd3_1 hold67 (.A(\data[2] ),
    .X(net78));
 sg13g2_dlygate4sd3_1 hold68 (.A(_038_),
    .X(net104));
 sg13g2_dlygate4sd3_1 hold69 (.A(\data[1] ),
    .X(net105));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_fill_2 FILLER_14_406 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_252 ();
 sg13g2_decap_8 FILLER_15_259 ();
 sg13g2_decap_8 FILLER_15_266 ();
 sg13g2_decap_8 FILLER_15_273 ();
 sg13g2_decap_8 FILLER_15_280 ();
 sg13g2_decap_8 FILLER_15_287 ();
 sg13g2_decap_8 FILLER_15_294 ();
 sg13g2_decap_8 FILLER_15_301 ();
 sg13g2_decap_8 FILLER_15_308 ();
 sg13g2_decap_8 FILLER_15_315 ();
 sg13g2_decap_8 FILLER_15_322 ();
 sg13g2_decap_8 FILLER_15_329 ();
 sg13g2_decap_8 FILLER_15_336 ();
 sg13g2_decap_8 FILLER_15_343 ();
 sg13g2_decap_8 FILLER_15_350 ();
 sg13g2_decap_8 FILLER_15_357 ();
 sg13g2_decap_8 FILLER_15_364 ();
 sg13g2_decap_8 FILLER_15_371 ();
 sg13g2_decap_8 FILLER_15_378 ();
 sg13g2_decap_8 FILLER_15_385 ();
 sg13g2_decap_8 FILLER_15_392 ();
 sg13g2_decap_8 FILLER_15_399 ();
 sg13g2_fill_2 FILLER_15_406 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_decap_8 FILLER_16_217 ();
 sg13g2_decap_8 FILLER_16_224 ();
 sg13g2_decap_8 FILLER_16_231 ();
 sg13g2_decap_8 FILLER_16_238 ();
 sg13g2_decap_8 FILLER_16_245 ();
 sg13g2_decap_8 FILLER_16_252 ();
 sg13g2_decap_8 FILLER_16_259 ();
 sg13g2_decap_8 FILLER_16_266 ();
 sg13g2_decap_8 FILLER_16_273 ();
 sg13g2_decap_8 FILLER_16_280 ();
 sg13g2_decap_8 FILLER_16_287 ();
 sg13g2_decap_8 FILLER_16_294 ();
 sg13g2_decap_8 FILLER_16_301 ();
 sg13g2_decap_8 FILLER_16_308 ();
 sg13g2_decap_8 FILLER_16_315 ();
 sg13g2_decap_8 FILLER_16_322 ();
 sg13g2_decap_8 FILLER_16_329 ();
 sg13g2_decap_8 FILLER_16_336 ();
 sg13g2_decap_8 FILLER_16_343 ();
 sg13g2_decap_8 FILLER_16_350 ();
 sg13g2_decap_8 FILLER_16_357 ();
 sg13g2_decap_8 FILLER_16_364 ();
 sg13g2_decap_8 FILLER_16_371 ();
 sg13g2_decap_8 FILLER_16_378 ();
 sg13g2_decap_8 FILLER_16_385 ();
 sg13g2_decap_8 FILLER_16_392 ();
 sg13g2_decap_8 FILLER_16_399 ();
 sg13g2_fill_2 FILLER_16_406 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_decap_8 FILLER_17_168 ();
 sg13g2_decap_8 FILLER_17_175 ();
 sg13g2_decap_8 FILLER_17_182 ();
 sg13g2_decap_8 FILLER_17_189 ();
 sg13g2_decap_8 FILLER_17_196 ();
 sg13g2_decap_8 FILLER_17_203 ();
 sg13g2_decap_8 FILLER_17_210 ();
 sg13g2_decap_8 FILLER_17_217 ();
 sg13g2_decap_8 FILLER_17_224 ();
 sg13g2_decap_8 FILLER_17_231 ();
 sg13g2_decap_8 FILLER_17_238 ();
 sg13g2_decap_8 FILLER_17_245 ();
 sg13g2_decap_8 FILLER_17_252 ();
 sg13g2_decap_8 FILLER_17_259 ();
 sg13g2_decap_8 FILLER_17_266 ();
 sg13g2_decap_8 FILLER_17_273 ();
 sg13g2_decap_8 FILLER_17_280 ();
 sg13g2_decap_8 FILLER_17_287 ();
 sg13g2_decap_8 FILLER_17_294 ();
 sg13g2_decap_8 FILLER_17_301 ();
 sg13g2_decap_8 FILLER_17_308 ();
 sg13g2_decap_8 FILLER_17_315 ();
 sg13g2_decap_8 FILLER_17_322 ();
 sg13g2_decap_8 FILLER_17_329 ();
 sg13g2_decap_8 FILLER_17_336 ();
 sg13g2_decap_8 FILLER_17_343 ();
 sg13g2_decap_8 FILLER_17_350 ();
 sg13g2_decap_8 FILLER_17_357 ();
 sg13g2_decap_8 FILLER_17_364 ();
 sg13g2_decap_8 FILLER_17_371 ();
 sg13g2_decap_8 FILLER_17_378 ();
 sg13g2_decap_8 FILLER_17_385 ();
 sg13g2_decap_8 FILLER_17_392 ();
 sg13g2_decap_8 FILLER_17_399 ();
 sg13g2_fill_2 FILLER_17_406 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_decap_8 FILLER_18_147 ();
 sg13g2_decap_8 FILLER_18_154 ();
 sg13g2_decap_8 FILLER_18_161 ();
 sg13g2_decap_8 FILLER_18_168 ();
 sg13g2_decap_8 FILLER_18_175 ();
 sg13g2_decap_8 FILLER_18_182 ();
 sg13g2_decap_8 FILLER_18_189 ();
 sg13g2_decap_8 FILLER_18_196 ();
 sg13g2_decap_8 FILLER_18_203 ();
 sg13g2_decap_8 FILLER_18_210 ();
 sg13g2_decap_8 FILLER_18_217 ();
 sg13g2_decap_8 FILLER_18_224 ();
 sg13g2_decap_8 FILLER_18_231 ();
 sg13g2_decap_8 FILLER_18_238 ();
 sg13g2_decap_8 FILLER_18_245 ();
 sg13g2_decap_8 FILLER_18_252 ();
 sg13g2_decap_8 FILLER_18_259 ();
 sg13g2_decap_8 FILLER_18_266 ();
 sg13g2_decap_8 FILLER_18_273 ();
 sg13g2_decap_8 FILLER_18_280 ();
 sg13g2_decap_8 FILLER_18_287 ();
 sg13g2_decap_8 FILLER_18_294 ();
 sg13g2_decap_8 FILLER_18_301 ();
 sg13g2_decap_8 FILLER_18_308 ();
 sg13g2_decap_8 FILLER_18_315 ();
 sg13g2_decap_8 FILLER_18_322 ();
 sg13g2_decap_8 FILLER_18_329 ();
 sg13g2_decap_8 FILLER_18_336 ();
 sg13g2_decap_8 FILLER_18_343 ();
 sg13g2_decap_8 FILLER_18_350 ();
 sg13g2_decap_8 FILLER_18_357 ();
 sg13g2_decap_8 FILLER_18_364 ();
 sg13g2_decap_8 FILLER_18_371 ();
 sg13g2_decap_8 FILLER_18_378 ();
 sg13g2_decap_8 FILLER_18_385 ();
 sg13g2_decap_8 FILLER_18_392 ();
 sg13g2_decap_8 FILLER_18_399 ();
 sg13g2_fill_2 FILLER_18_406 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_decap_8 FILLER_19_140 ();
 sg13g2_decap_8 FILLER_19_147 ();
 sg13g2_decap_8 FILLER_19_154 ();
 sg13g2_decap_8 FILLER_19_161 ();
 sg13g2_decap_8 FILLER_19_168 ();
 sg13g2_decap_8 FILLER_19_175 ();
 sg13g2_decap_8 FILLER_19_182 ();
 sg13g2_decap_8 FILLER_19_189 ();
 sg13g2_decap_8 FILLER_19_196 ();
 sg13g2_decap_8 FILLER_19_203 ();
 sg13g2_decap_8 FILLER_19_210 ();
 sg13g2_decap_8 FILLER_19_217 ();
 sg13g2_decap_8 FILLER_19_224 ();
 sg13g2_decap_8 FILLER_19_231 ();
 sg13g2_decap_8 FILLER_19_238 ();
 sg13g2_decap_8 FILLER_19_245 ();
 sg13g2_decap_8 FILLER_19_252 ();
 sg13g2_decap_8 FILLER_19_259 ();
 sg13g2_decap_8 FILLER_19_266 ();
 sg13g2_decap_8 FILLER_19_273 ();
 sg13g2_decap_8 FILLER_19_280 ();
 sg13g2_decap_8 FILLER_19_287 ();
 sg13g2_decap_8 FILLER_19_294 ();
 sg13g2_decap_8 FILLER_19_301 ();
 sg13g2_decap_8 FILLER_19_308 ();
 sg13g2_decap_8 FILLER_19_315 ();
 sg13g2_decap_8 FILLER_19_322 ();
 sg13g2_decap_8 FILLER_19_329 ();
 sg13g2_decap_8 FILLER_19_336 ();
 sg13g2_decap_8 FILLER_19_343 ();
 sg13g2_decap_8 FILLER_19_350 ();
 sg13g2_decap_8 FILLER_19_357 ();
 sg13g2_decap_8 FILLER_19_364 ();
 sg13g2_decap_8 FILLER_19_371 ();
 sg13g2_decap_8 FILLER_19_378 ();
 sg13g2_decap_8 FILLER_19_385 ();
 sg13g2_decap_8 FILLER_19_392 ();
 sg13g2_decap_8 FILLER_19_399 ();
 sg13g2_fill_2 FILLER_19_406 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_decap_8 FILLER_20_126 ();
 sg13g2_decap_8 FILLER_20_133 ();
 sg13g2_decap_8 FILLER_20_140 ();
 sg13g2_decap_8 FILLER_20_147 ();
 sg13g2_decap_8 FILLER_20_154 ();
 sg13g2_decap_8 FILLER_20_161 ();
 sg13g2_decap_8 FILLER_20_168 ();
 sg13g2_decap_8 FILLER_20_175 ();
 sg13g2_decap_8 FILLER_20_182 ();
 sg13g2_decap_8 FILLER_20_189 ();
 sg13g2_decap_8 FILLER_20_196 ();
 sg13g2_decap_8 FILLER_20_203 ();
 sg13g2_decap_8 FILLER_20_210 ();
 sg13g2_decap_8 FILLER_20_217 ();
 sg13g2_decap_8 FILLER_20_224 ();
 sg13g2_decap_8 FILLER_20_231 ();
 sg13g2_decap_8 FILLER_20_238 ();
 sg13g2_decap_8 FILLER_20_245 ();
 sg13g2_decap_8 FILLER_20_252 ();
 sg13g2_decap_8 FILLER_20_259 ();
 sg13g2_decap_8 FILLER_20_266 ();
 sg13g2_decap_8 FILLER_20_273 ();
 sg13g2_decap_8 FILLER_20_280 ();
 sg13g2_decap_8 FILLER_20_287 ();
 sg13g2_decap_8 FILLER_20_294 ();
 sg13g2_decap_8 FILLER_20_301 ();
 sg13g2_decap_8 FILLER_20_308 ();
 sg13g2_decap_8 FILLER_20_315 ();
 sg13g2_decap_8 FILLER_20_322 ();
 sg13g2_decap_8 FILLER_20_329 ();
 sg13g2_decap_8 FILLER_20_336 ();
 sg13g2_decap_8 FILLER_20_343 ();
 sg13g2_decap_8 FILLER_20_350 ();
 sg13g2_decap_8 FILLER_20_357 ();
 sg13g2_decap_8 FILLER_20_364 ();
 sg13g2_decap_8 FILLER_20_371 ();
 sg13g2_decap_8 FILLER_20_378 ();
 sg13g2_decap_8 FILLER_20_385 ();
 sg13g2_decap_8 FILLER_20_392 ();
 sg13g2_decap_8 FILLER_20_399 ();
 sg13g2_fill_2 FILLER_20_406 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_decap_8 FILLER_21_119 ();
 sg13g2_decap_8 FILLER_21_126 ();
 sg13g2_decap_8 FILLER_21_133 ();
 sg13g2_decap_8 FILLER_21_140 ();
 sg13g2_decap_8 FILLER_21_147 ();
 sg13g2_decap_8 FILLER_21_154 ();
 sg13g2_decap_8 FILLER_21_161 ();
 sg13g2_decap_8 FILLER_21_168 ();
 sg13g2_decap_8 FILLER_21_175 ();
 sg13g2_decap_8 FILLER_21_182 ();
 sg13g2_decap_8 FILLER_21_189 ();
 sg13g2_decap_8 FILLER_21_196 ();
 sg13g2_decap_8 FILLER_21_203 ();
 sg13g2_decap_8 FILLER_21_210 ();
 sg13g2_decap_8 FILLER_21_217 ();
 sg13g2_decap_8 FILLER_21_224 ();
 sg13g2_decap_8 FILLER_21_231 ();
 sg13g2_decap_8 FILLER_21_238 ();
 sg13g2_decap_8 FILLER_21_245 ();
 sg13g2_decap_8 FILLER_21_252 ();
 sg13g2_decap_8 FILLER_21_259 ();
 sg13g2_decap_8 FILLER_21_266 ();
 sg13g2_decap_8 FILLER_21_273 ();
 sg13g2_decap_8 FILLER_21_280 ();
 sg13g2_decap_8 FILLER_21_287 ();
 sg13g2_decap_8 FILLER_21_294 ();
 sg13g2_decap_8 FILLER_21_301 ();
 sg13g2_decap_8 FILLER_21_308 ();
 sg13g2_decap_8 FILLER_21_315 ();
 sg13g2_decap_8 FILLER_21_322 ();
 sg13g2_decap_8 FILLER_21_329 ();
 sg13g2_decap_8 FILLER_21_336 ();
 sg13g2_decap_8 FILLER_21_343 ();
 sg13g2_decap_8 FILLER_21_350 ();
 sg13g2_decap_8 FILLER_21_357 ();
 sg13g2_decap_8 FILLER_21_364 ();
 sg13g2_decap_8 FILLER_21_371 ();
 sg13g2_decap_8 FILLER_21_378 ();
 sg13g2_decap_8 FILLER_21_385 ();
 sg13g2_decap_8 FILLER_21_392 ();
 sg13g2_decap_8 FILLER_21_399 ();
 sg13g2_fill_2 FILLER_21_406 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_8 FILLER_22_105 ();
 sg13g2_decap_8 FILLER_22_112 ();
 sg13g2_decap_8 FILLER_22_119 ();
 sg13g2_decap_8 FILLER_22_126 ();
 sg13g2_decap_8 FILLER_22_133 ();
 sg13g2_decap_8 FILLER_22_140 ();
 sg13g2_decap_8 FILLER_22_147 ();
 sg13g2_decap_8 FILLER_22_154 ();
 sg13g2_decap_8 FILLER_22_161 ();
 sg13g2_decap_8 FILLER_22_168 ();
 sg13g2_decap_8 FILLER_22_175 ();
 sg13g2_decap_8 FILLER_22_182 ();
 sg13g2_decap_8 FILLER_22_189 ();
 sg13g2_decap_8 FILLER_22_196 ();
 sg13g2_decap_8 FILLER_22_203 ();
 sg13g2_decap_8 FILLER_22_210 ();
 sg13g2_decap_8 FILLER_22_217 ();
 sg13g2_decap_8 FILLER_22_224 ();
 sg13g2_decap_8 FILLER_22_231 ();
 sg13g2_decap_8 FILLER_22_238 ();
 sg13g2_decap_8 FILLER_22_245 ();
 sg13g2_decap_8 FILLER_22_252 ();
 sg13g2_decap_8 FILLER_22_259 ();
 sg13g2_decap_8 FILLER_22_266 ();
 sg13g2_decap_8 FILLER_22_273 ();
 sg13g2_decap_8 FILLER_22_280 ();
 sg13g2_decap_8 FILLER_22_287 ();
 sg13g2_decap_8 FILLER_22_294 ();
 sg13g2_decap_8 FILLER_22_301 ();
 sg13g2_decap_8 FILLER_22_308 ();
 sg13g2_decap_8 FILLER_22_315 ();
 sg13g2_decap_8 FILLER_22_322 ();
 sg13g2_decap_8 FILLER_22_329 ();
 sg13g2_decap_8 FILLER_22_336 ();
 sg13g2_decap_8 FILLER_22_343 ();
 sg13g2_decap_8 FILLER_22_350 ();
 sg13g2_decap_8 FILLER_22_357 ();
 sg13g2_decap_8 FILLER_22_364 ();
 sg13g2_decap_8 FILLER_22_371 ();
 sg13g2_decap_8 FILLER_22_378 ();
 sg13g2_decap_8 FILLER_22_385 ();
 sg13g2_decap_8 FILLER_22_392 ();
 sg13g2_decap_8 FILLER_22_399 ();
 sg13g2_fill_2 FILLER_22_406 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_fill_2 FILLER_23_84 ();
 sg13g2_fill_1 FILLER_23_86 ();
 sg13g2_decap_4 FILLER_23_96 ();
 sg13g2_fill_1 FILLER_23_100 ();
 sg13g2_decap_8 FILLER_23_111 ();
 sg13g2_fill_2 FILLER_23_118 ();
 sg13g2_fill_1 FILLER_23_120 ();
 sg13g2_fill_1 FILLER_23_147 ();
 sg13g2_decap_8 FILLER_23_153 ();
 sg13g2_decap_8 FILLER_23_160 ();
 sg13g2_decap_8 FILLER_23_167 ();
 sg13g2_decap_8 FILLER_23_174 ();
 sg13g2_decap_8 FILLER_23_181 ();
 sg13g2_decap_8 FILLER_23_188 ();
 sg13g2_decap_8 FILLER_23_195 ();
 sg13g2_decap_8 FILLER_23_202 ();
 sg13g2_decap_8 FILLER_23_209 ();
 sg13g2_decap_8 FILLER_23_216 ();
 sg13g2_decap_8 FILLER_23_223 ();
 sg13g2_decap_8 FILLER_23_230 ();
 sg13g2_decap_8 FILLER_23_237 ();
 sg13g2_decap_8 FILLER_23_244 ();
 sg13g2_decap_8 FILLER_23_251 ();
 sg13g2_decap_8 FILLER_23_258 ();
 sg13g2_decap_8 FILLER_23_265 ();
 sg13g2_decap_8 FILLER_23_272 ();
 sg13g2_decap_8 FILLER_23_279 ();
 sg13g2_decap_8 FILLER_23_286 ();
 sg13g2_decap_8 FILLER_23_293 ();
 sg13g2_decap_8 FILLER_23_300 ();
 sg13g2_decap_8 FILLER_23_307 ();
 sg13g2_decap_8 FILLER_23_314 ();
 sg13g2_decap_8 FILLER_23_321 ();
 sg13g2_decap_8 FILLER_23_328 ();
 sg13g2_decap_8 FILLER_23_335 ();
 sg13g2_decap_8 FILLER_23_342 ();
 sg13g2_decap_8 FILLER_23_349 ();
 sg13g2_decap_8 FILLER_23_356 ();
 sg13g2_decap_8 FILLER_23_363 ();
 sg13g2_decap_8 FILLER_23_370 ();
 sg13g2_decap_8 FILLER_23_377 ();
 sg13g2_decap_8 FILLER_23_384 ();
 sg13g2_decap_8 FILLER_23_391 ();
 sg13g2_decap_8 FILLER_23_398 ();
 sg13g2_decap_4 FILLER_23_405 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_4 FILLER_24_56 ();
 sg13g2_fill_1 FILLER_24_60 ();
 sg13g2_decap_8 FILLER_24_113 ();
 sg13g2_decap_4 FILLER_24_120 ();
 sg13g2_fill_1 FILLER_24_124 ();
 sg13g2_decap_4 FILLER_24_135 ();
 sg13g2_decap_8 FILLER_24_165 ();
 sg13g2_fill_2 FILLER_24_172 ();
 sg13g2_fill_1 FILLER_24_174 ();
 sg13g2_fill_2 FILLER_24_183 ();
 sg13g2_decap_8 FILLER_24_194 ();
 sg13g2_decap_8 FILLER_24_201 ();
 sg13g2_fill_1 FILLER_24_208 ();
 sg13g2_decap_8 FILLER_24_213 ();
 sg13g2_fill_2 FILLER_24_220 ();
 sg13g2_decap_8 FILLER_24_231 ();
 sg13g2_decap_8 FILLER_24_238 ();
 sg13g2_decap_8 FILLER_24_245 ();
 sg13g2_decap_8 FILLER_24_252 ();
 sg13g2_decap_8 FILLER_24_259 ();
 sg13g2_decap_8 FILLER_24_266 ();
 sg13g2_decap_8 FILLER_24_273 ();
 sg13g2_decap_8 FILLER_24_280 ();
 sg13g2_decap_8 FILLER_24_287 ();
 sg13g2_decap_8 FILLER_24_294 ();
 sg13g2_decap_8 FILLER_24_301 ();
 sg13g2_decap_8 FILLER_24_308 ();
 sg13g2_decap_8 FILLER_24_315 ();
 sg13g2_decap_8 FILLER_24_322 ();
 sg13g2_decap_8 FILLER_24_329 ();
 sg13g2_decap_8 FILLER_24_336 ();
 sg13g2_decap_8 FILLER_24_343 ();
 sg13g2_decap_8 FILLER_24_350 ();
 sg13g2_decap_8 FILLER_24_357 ();
 sg13g2_decap_8 FILLER_24_364 ();
 sg13g2_decap_8 FILLER_24_371 ();
 sg13g2_decap_8 FILLER_24_378 ();
 sg13g2_decap_8 FILLER_24_385 ();
 sg13g2_decap_8 FILLER_24_392 ();
 sg13g2_decap_8 FILLER_24_399 ();
 sg13g2_fill_2 FILLER_24_406 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_fill_1 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_27 ();
 sg13g2_decap_8 FILLER_25_34 ();
 sg13g2_fill_2 FILLER_25_41 ();
 sg13g2_fill_1 FILLER_25_43 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_4 FILLER_25_77 ();
 sg13g2_fill_2 FILLER_25_81 ();
 sg13g2_decap_8 FILLER_25_108 ();
 sg13g2_fill_2 FILLER_25_115 ();
 sg13g2_fill_1 FILLER_25_117 ();
 sg13g2_fill_1 FILLER_25_131 ();
 sg13g2_fill_1 FILLER_25_155 ();
 sg13g2_decap_4 FILLER_25_235 ();
 sg13g2_decap_8 FILLER_25_248 ();
 sg13g2_decap_8 FILLER_25_255 ();
 sg13g2_decap_8 FILLER_25_262 ();
 sg13g2_decap_8 FILLER_25_269 ();
 sg13g2_decap_8 FILLER_25_276 ();
 sg13g2_decap_8 FILLER_25_283 ();
 sg13g2_decap_8 FILLER_25_290 ();
 sg13g2_decap_8 FILLER_25_297 ();
 sg13g2_decap_8 FILLER_25_304 ();
 sg13g2_decap_8 FILLER_25_311 ();
 sg13g2_decap_8 FILLER_25_318 ();
 sg13g2_decap_8 FILLER_25_325 ();
 sg13g2_decap_8 FILLER_25_332 ();
 sg13g2_decap_8 FILLER_25_339 ();
 sg13g2_decap_8 FILLER_25_346 ();
 sg13g2_decap_8 FILLER_25_353 ();
 sg13g2_decap_8 FILLER_25_360 ();
 sg13g2_decap_8 FILLER_25_367 ();
 sg13g2_decap_8 FILLER_25_374 ();
 sg13g2_decap_8 FILLER_25_381 ();
 sg13g2_decap_8 FILLER_25_388 ();
 sg13g2_decap_8 FILLER_25_395 ();
 sg13g2_decap_8 FILLER_25_402 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_4 FILLER_26_7 ();
 sg13g2_fill_2 FILLER_26_11 ();
 sg13g2_fill_2 FILLER_26_75 ();
 sg13g2_fill_1 FILLER_26_85 ();
 sg13g2_fill_1 FILLER_26_99 ();
 sg13g2_decap_8 FILLER_26_254 ();
 sg13g2_decap_8 FILLER_26_261 ();
 sg13g2_decap_8 FILLER_26_268 ();
 sg13g2_decap_8 FILLER_26_275 ();
 sg13g2_decap_8 FILLER_26_282 ();
 sg13g2_decap_8 FILLER_26_289 ();
 sg13g2_decap_8 FILLER_26_296 ();
 sg13g2_decap_8 FILLER_26_303 ();
 sg13g2_decap_8 FILLER_26_310 ();
 sg13g2_decap_8 FILLER_26_317 ();
 sg13g2_decap_8 FILLER_26_324 ();
 sg13g2_decap_8 FILLER_26_331 ();
 sg13g2_decap_8 FILLER_26_338 ();
 sg13g2_decap_8 FILLER_26_345 ();
 sg13g2_decap_8 FILLER_26_352 ();
 sg13g2_decap_8 FILLER_26_359 ();
 sg13g2_decap_8 FILLER_26_366 ();
 sg13g2_decap_8 FILLER_26_373 ();
 sg13g2_decap_8 FILLER_26_380 ();
 sg13g2_decap_8 FILLER_26_387 ();
 sg13g2_decap_8 FILLER_26_394 ();
 sg13g2_decap_8 FILLER_26_401 ();
 sg13g2_fill_1 FILLER_26_408 ();
 sg13g2_decap_4 FILLER_27_0 ();
 sg13g2_fill_1 FILLER_27_4 ();
 sg13g2_fill_2 FILLER_27_15 ();
 sg13g2_fill_1 FILLER_27_17 ();
 sg13g2_fill_2 FILLER_27_32 ();
 sg13g2_fill_1 FILLER_27_34 ();
 sg13g2_decap_8 FILLER_27_44 ();
 sg13g2_fill_1 FILLER_27_51 ();
 sg13g2_decap_8 FILLER_27_61 ();
 sg13g2_fill_2 FILLER_27_68 ();
 sg13g2_fill_2 FILLER_27_89 ();
 sg13g2_fill_1 FILLER_27_91 ();
 sg13g2_decap_4 FILLER_27_97 ();
 sg13g2_decap_4 FILLER_27_140 ();
 sg13g2_fill_1 FILLER_27_147 ();
 sg13g2_fill_1 FILLER_27_175 ();
 sg13g2_fill_2 FILLER_27_189 ();
 sg13g2_fill_1 FILLER_27_191 ();
 sg13g2_decap_8 FILLER_27_249 ();
 sg13g2_decap_8 FILLER_27_256 ();
 sg13g2_decap_8 FILLER_27_263 ();
 sg13g2_decap_8 FILLER_27_270 ();
 sg13g2_decap_8 FILLER_27_277 ();
 sg13g2_decap_8 FILLER_27_284 ();
 sg13g2_decap_8 FILLER_27_291 ();
 sg13g2_decap_8 FILLER_27_298 ();
 sg13g2_decap_8 FILLER_27_305 ();
 sg13g2_decap_8 FILLER_27_312 ();
 sg13g2_decap_8 FILLER_27_319 ();
 sg13g2_decap_8 FILLER_27_326 ();
 sg13g2_decap_8 FILLER_27_333 ();
 sg13g2_decap_8 FILLER_27_340 ();
 sg13g2_decap_8 FILLER_27_347 ();
 sg13g2_decap_8 FILLER_27_354 ();
 sg13g2_decap_8 FILLER_27_361 ();
 sg13g2_decap_8 FILLER_27_368 ();
 sg13g2_decap_8 FILLER_27_375 ();
 sg13g2_decap_8 FILLER_27_382 ();
 sg13g2_decap_8 FILLER_27_389 ();
 sg13g2_decap_8 FILLER_27_396 ();
 sg13g2_decap_4 FILLER_27_403 ();
 sg13g2_fill_2 FILLER_27_407 ();
 sg13g2_decap_4 FILLER_28_0 ();
 sg13g2_fill_1 FILLER_28_14 ();
 sg13g2_fill_2 FILLER_28_115 ();
 sg13g2_fill_1 FILLER_28_137 ();
 sg13g2_fill_2 FILLER_28_150 ();
 sg13g2_decap_4 FILLER_28_162 ();
 sg13g2_fill_2 FILLER_28_166 ();
 sg13g2_fill_2 FILLER_28_176 ();
 sg13g2_fill_1 FILLER_28_186 ();
 sg13g2_fill_2 FILLER_28_195 ();
 sg13g2_fill_2 FILLER_28_202 ();
 sg13g2_fill_1 FILLER_28_213 ();
 sg13g2_fill_2 FILLER_28_219 ();
 sg13g2_decap_8 FILLER_28_255 ();
 sg13g2_decap_8 FILLER_28_262 ();
 sg13g2_decap_8 FILLER_28_269 ();
 sg13g2_decap_8 FILLER_28_276 ();
 sg13g2_decap_8 FILLER_28_283 ();
 sg13g2_decap_8 FILLER_28_290 ();
 sg13g2_decap_8 FILLER_28_297 ();
 sg13g2_decap_8 FILLER_28_304 ();
 sg13g2_decap_8 FILLER_28_311 ();
 sg13g2_decap_8 FILLER_28_318 ();
 sg13g2_decap_8 FILLER_28_325 ();
 sg13g2_decap_8 FILLER_28_332 ();
 sg13g2_decap_8 FILLER_28_339 ();
 sg13g2_decap_8 FILLER_28_346 ();
 sg13g2_decap_8 FILLER_28_353 ();
 sg13g2_decap_8 FILLER_28_360 ();
 sg13g2_decap_8 FILLER_28_367 ();
 sg13g2_decap_8 FILLER_28_374 ();
 sg13g2_decap_8 FILLER_28_381 ();
 sg13g2_decap_8 FILLER_28_388 ();
 sg13g2_decap_8 FILLER_28_395 ();
 sg13g2_decap_8 FILLER_28_402 ();
 sg13g2_decap_4 FILLER_29_52 ();
 sg13g2_fill_2 FILLER_29_56 ();
 sg13g2_decap_4 FILLER_29_67 ();
 sg13g2_fill_2 FILLER_29_71 ();
 sg13g2_fill_1 FILLER_29_88 ();
 sg13g2_fill_1 FILLER_29_145 ();
 sg13g2_fill_2 FILLER_29_168 ();
 sg13g2_fill_2 FILLER_29_194 ();
 sg13g2_fill_2 FILLER_29_204 ();
 sg13g2_fill_1 FILLER_29_235 ();
 sg13g2_decap_8 FILLER_29_255 ();
 sg13g2_decap_8 FILLER_29_262 ();
 sg13g2_decap_8 FILLER_29_269 ();
 sg13g2_decap_8 FILLER_29_276 ();
 sg13g2_decap_8 FILLER_29_283 ();
 sg13g2_decap_8 FILLER_29_290 ();
 sg13g2_decap_8 FILLER_29_297 ();
 sg13g2_decap_8 FILLER_29_304 ();
 sg13g2_decap_8 FILLER_29_311 ();
 sg13g2_decap_8 FILLER_29_318 ();
 sg13g2_decap_8 FILLER_29_325 ();
 sg13g2_decap_8 FILLER_29_332 ();
 sg13g2_decap_8 FILLER_29_339 ();
 sg13g2_decap_8 FILLER_29_346 ();
 sg13g2_decap_8 FILLER_29_353 ();
 sg13g2_decap_8 FILLER_29_360 ();
 sg13g2_decap_8 FILLER_29_367 ();
 sg13g2_decap_8 FILLER_29_374 ();
 sg13g2_decap_8 FILLER_29_381 ();
 sg13g2_decap_8 FILLER_29_388 ();
 sg13g2_decap_8 FILLER_29_395 ();
 sg13g2_decap_8 FILLER_29_402 ();
 sg13g2_decap_4 FILLER_30_0 ();
 sg13g2_decap_4 FILLER_30_34 ();
 sg13g2_fill_1 FILLER_30_74 ();
 sg13g2_decap_8 FILLER_30_86 ();
 sg13g2_fill_2 FILLER_30_93 ();
 sg13g2_fill_1 FILLER_30_108 ();
 sg13g2_fill_2 FILLER_30_180 ();
 sg13g2_fill_1 FILLER_30_182 ();
 sg13g2_decap_4 FILLER_30_188 ();
 sg13g2_fill_1 FILLER_30_197 ();
 sg13g2_fill_2 FILLER_30_203 ();
 sg13g2_fill_1 FILLER_30_205 ();
 sg13g2_decap_8 FILLER_30_267 ();
 sg13g2_decap_8 FILLER_30_274 ();
 sg13g2_decap_8 FILLER_30_281 ();
 sg13g2_decap_8 FILLER_30_288 ();
 sg13g2_decap_8 FILLER_30_295 ();
 sg13g2_decap_8 FILLER_30_302 ();
 sg13g2_decap_8 FILLER_30_309 ();
 sg13g2_decap_8 FILLER_30_316 ();
 sg13g2_decap_8 FILLER_30_323 ();
 sg13g2_decap_8 FILLER_30_330 ();
 sg13g2_decap_8 FILLER_30_337 ();
 sg13g2_decap_8 FILLER_30_344 ();
 sg13g2_decap_8 FILLER_30_351 ();
 sg13g2_decap_8 FILLER_30_358 ();
 sg13g2_decap_8 FILLER_30_365 ();
 sg13g2_decap_8 FILLER_30_372 ();
 sg13g2_decap_8 FILLER_30_379 ();
 sg13g2_decap_8 FILLER_30_386 ();
 sg13g2_decap_8 FILLER_30_393 ();
 sg13g2_decap_8 FILLER_30_400 ();
 sg13g2_fill_2 FILLER_30_407 ();
 sg13g2_fill_1 FILLER_31_0 ();
 sg13g2_fill_2 FILLER_31_27 ();
 sg13g2_fill_1 FILLER_31_29 ();
 sg13g2_fill_1 FILLER_31_73 ();
 sg13g2_fill_2 FILLER_31_135 ();
 sg13g2_fill_1 FILLER_31_137 ();
 sg13g2_fill_2 FILLER_31_147 ();
 sg13g2_decap_4 FILLER_31_169 ();
 sg13g2_decap_8 FILLER_31_193 ();
 sg13g2_fill_1 FILLER_31_205 ();
 sg13g2_fill_2 FILLER_31_224 ();
 sg13g2_fill_1 FILLER_31_226 ();
 sg13g2_decap_4 FILLER_31_236 ();
 sg13g2_decap_8 FILLER_31_253 ();
 sg13g2_decap_8 FILLER_31_260 ();
 sg13g2_decap_8 FILLER_31_267 ();
 sg13g2_decap_8 FILLER_31_274 ();
 sg13g2_decap_8 FILLER_31_281 ();
 sg13g2_decap_8 FILLER_31_288 ();
 sg13g2_decap_8 FILLER_31_295 ();
 sg13g2_decap_8 FILLER_31_302 ();
 sg13g2_decap_8 FILLER_31_309 ();
 sg13g2_decap_8 FILLER_31_316 ();
 sg13g2_decap_8 FILLER_31_323 ();
 sg13g2_decap_8 FILLER_31_330 ();
 sg13g2_decap_8 FILLER_31_337 ();
 sg13g2_decap_8 FILLER_31_344 ();
 sg13g2_decap_8 FILLER_31_351 ();
 sg13g2_decap_8 FILLER_31_358 ();
 sg13g2_decap_8 FILLER_31_365 ();
 sg13g2_decap_8 FILLER_31_372 ();
 sg13g2_decap_8 FILLER_31_379 ();
 sg13g2_decap_8 FILLER_31_386 ();
 sg13g2_decap_8 FILLER_31_393 ();
 sg13g2_decap_8 FILLER_31_400 ();
 sg13g2_fill_2 FILLER_31_407 ();
 sg13g2_decap_4 FILLER_32_0 ();
 sg13g2_fill_1 FILLER_32_13 ();
 sg13g2_decap_8 FILLER_32_33 ();
 sg13g2_fill_1 FILLER_32_40 ();
 sg13g2_fill_1 FILLER_32_67 ();
 sg13g2_fill_1 FILLER_32_85 ();
 sg13g2_fill_2 FILLER_32_104 ();
 sg13g2_fill_1 FILLER_32_106 ();
 sg13g2_fill_2 FILLER_32_121 ();
 sg13g2_fill_1 FILLER_32_123 ();
 sg13g2_fill_2 FILLER_32_150 ();
 sg13g2_decap_4 FILLER_32_175 ();
 sg13g2_fill_1 FILLER_32_179 ();
 sg13g2_fill_2 FILLER_32_215 ();
 sg13g2_decap_8 FILLER_32_267 ();
 sg13g2_decap_8 FILLER_32_274 ();
 sg13g2_decap_8 FILLER_32_281 ();
 sg13g2_decap_8 FILLER_32_288 ();
 sg13g2_decap_8 FILLER_32_295 ();
 sg13g2_decap_8 FILLER_32_302 ();
 sg13g2_decap_8 FILLER_32_309 ();
 sg13g2_decap_8 FILLER_32_316 ();
 sg13g2_decap_8 FILLER_32_323 ();
 sg13g2_decap_8 FILLER_32_330 ();
 sg13g2_decap_8 FILLER_32_337 ();
 sg13g2_decap_8 FILLER_32_344 ();
 sg13g2_decap_8 FILLER_32_351 ();
 sg13g2_decap_8 FILLER_32_358 ();
 sg13g2_decap_8 FILLER_32_365 ();
 sg13g2_decap_8 FILLER_32_372 ();
 sg13g2_decap_8 FILLER_32_379 ();
 sg13g2_decap_8 FILLER_32_386 ();
 sg13g2_decap_8 FILLER_32_393 ();
 sg13g2_decap_8 FILLER_32_400 ();
 sg13g2_fill_2 FILLER_32_407 ();
 sg13g2_decap_4 FILLER_33_0 ();
 sg13g2_fill_2 FILLER_33_59 ();
 sg13g2_fill_1 FILLER_33_61 ();
 sg13g2_fill_2 FILLER_33_131 ();
 sg13g2_fill_1 FILLER_33_133 ();
 sg13g2_fill_1 FILLER_33_148 ();
 sg13g2_decap_8 FILLER_33_175 ();
 sg13g2_fill_2 FILLER_33_182 ();
 sg13g2_decap_8 FILLER_33_193 ();
 sg13g2_fill_2 FILLER_33_200 ();
 sg13g2_decap_4 FILLER_33_206 ();
 sg13g2_fill_2 FILLER_33_210 ();
 sg13g2_decap_8 FILLER_33_231 ();
 sg13g2_decap_4 FILLER_33_238 ();
 sg13g2_fill_2 FILLER_33_242 ();
 sg13g2_fill_2 FILLER_33_255 ();
 sg13g2_fill_1 FILLER_33_257 ();
 sg13g2_decap_8 FILLER_33_263 ();
 sg13g2_decap_8 FILLER_33_270 ();
 sg13g2_decap_8 FILLER_33_277 ();
 sg13g2_decap_8 FILLER_33_284 ();
 sg13g2_decap_8 FILLER_33_291 ();
 sg13g2_decap_8 FILLER_33_298 ();
 sg13g2_decap_8 FILLER_33_305 ();
 sg13g2_decap_8 FILLER_33_312 ();
 sg13g2_decap_8 FILLER_33_319 ();
 sg13g2_decap_8 FILLER_33_326 ();
 sg13g2_decap_8 FILLER_33_333 ();
 sg13g2_decap_8 FILLER_33_340 ();
 sg13g2_decap_8 FILLER_33_347 ();
 sg13g2_decap_8 FILLER_33_354 ();
 sg13g2_decap_8 FILLER_33_361 ();
 sg13g2_decap_8 FILLER_33_368 ();
 sg13g2_decap_8 FILLER_33_375 ();
 sg13g2_decap_8 FILLER_33_382 ();
 sg13g2_decap_8 FILLER_33_389 ();
 sg13g2_decap_8 FILLER_33_396 ();
 sg13g2_decap_4 FILLER_33_403 ();
 sg13g2_fill_2 FILLER_33_407 ();
 sg13g2_fill_2 FILLER_34_0 ();
 sg13g2_fill_1 FILLER_34_2 ();
 sg13g2_decap_4 FILLER_34_29 ();
 sg13g2_fill_1 FILLER_34_53 ();
 sg13g2_fill_2 FILLER_34_67 ();
 sg13g2_fill_2 FILLER_34_104 ();
 sg13g2_fill_1 FILLER_34_106 ();
 sg13g2_fill_2 FILLER_34_144 ();
 sg13g2_fill_2 FILLER_34_190 ();
 sg13g2_fill_1 FILLER_34_192 ();
 sg13g2_decap_8 FILLER_34_209 ();
 sg13g2_fill_1 FILLER_34_216 ();
 sg13g2_fill_2 FILLER_34_234 ();
 sg13g2_fill_2 FILLER_34_255 ();
 sg13g2_fill_1 FILLER_34_257 ();
 sg13g2_decap_8 FILLER_34_272 ();
 sg13g2_decap_8 FILLER_34_279 ();
 sg13g2_decap_8 FILLER_34_286 ();
 sg13g2_decap_8 FILLER_34_293 ();
 sg13g2_decap_8 FILLER_34_300 ();
 sg13g2_decap_8 FILLER_34_307 ();
 sg13g2_decap_8 FILLER_34_314 ();
 sg13g2_decap_8 FILLER_34_321 ();
 sg13g2_decap_8 FILLER_34_328 ();
 sg13g2_decap_8 FILLER_34_335 ();
 sg13g2_decap_8 FILLER_34_342 ();
 sg13g2_decap_8 FILLER_34_349 ();
 sg13g2_decap_8 FILLER_34_356 ();
 sg13g2_decap_8 FILLER_34_363 ();
 sg13g2_decap_8 FILLER_34_370 ();
 sg13g2_decap_8 FILLER_34_377 ();
 sg13g2_decap_8 FILLER_34_384 ();
 sg13g2_decap_8 FILLER_34_391 ();
 sg13g2_decap_8 FILLER_34_398 ();
 sg13g2_decap_4 FILLER_34_405 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_fill_1 FILLER_35_7 ();
 sg13g2_fill_1 FILLER_35_39 ();
 sg13g2_fill_2 FILLER_35_66 ();
 sg13g2_fill_1 FILLER_35_87 ();
 sg13g2_fill_2 FILLER_35_98 ();
 sg13g2_fill_1 FILLER_35_100 ();
 sg13g2_decap_4 FILLER_35_152 ();
 sg13g2_decap_8 FILLER_35_172 ();
 sg13g2_decap_4 FILLER_35_179 ();
 sg13g2_fill_2 FILLER_35_191 ();
 sg13g2_fill_1 FILLER_35_193 ();
 sg13g2_fill_2 FILLER_35_204 ();
 sg13g2_fill_2 FILLER_35_217 ();
 sg13g2_fill_1 FILLER_35_219 ();
 sg13g2_fill_1 FILLER_35_237 ();
 sg13g2_fill_2 FILLER_35_243 ();
 sg13g2_fill_1 FILLER_35_245 ();
 sg13g2_decap_4 FILLER_35_250 ();
 sg13g2_decap_8 FILLER_35_277 ();
 sg13g2_decap_8 FILLER_35_284 ();
 sg13g2_decap_8 FILLER_35_291 ();
 sg13g2_decap_8 FILLER_35_298 ();
 sg13g2_decap_8 FILLER_35_305 ();
 sg13g2_decap_8 FILLER_35_312 ();
 sg13g2_decap_8 FILLER_35_319 ();
 sg13g2_decap_8 FILLER_35_326 ();
 sg13g2_decap_8 FILLER_35_333 ();
 sg13g2_decap_8 FILLER_35_340 ();
 sg13g2_decap_8 FILLER_35_347 ();
 sg13g2_decap_8 FILLER_35_354 ();
 sg13g2_decap_8 FILLER_35_361 ();
 sg13g2_decap_8 FILLER_35_368 ();
 sg13g2_decap_8 FILLER_35_375 ();
 sg13g2_decap_8 FILLER_35_382 ();
 sg13g2_decap_8 FILLER_35_389 ();
 sg13g2_decap_8 FILLER_35_396 ();
 sg13g2_decap_4 FILLER_35_403 ();
 sg13g2_fill_2 FILLER_35_407 ();
 sg13g2_decap_4 FILLER_36_0 ();
 sg13g2_fill_1 FILLER_36_4 ();
 sg13g2_fill_1 FILLER_36_24 ();
 sg13g2_fill_2 FILLER_36_34 ();
 sg13g2_fill_2 FILLER_36_46 ();
 sg13g2_fill_2 FILLER_36_83 ();
 sg13g2_fill_1 FILLER_36_119 ();
 sg13g2_decap_4 FILLER_36_165 ();
 sg13g2_decap_4 FILLER_36_179 ();
 sg13g2_fill_2 FILLER_36_183 ();
 sg13g2_decap_4 FILLER_36_197 ();
 sg13g2_fill_2 FILLER_36_201 ();
 sg13g2_decap_4 FILLER_36_207 ();
 sg13g2_fill_2 FILLER_36_226 ();
 sg13g2_fill_2 FILLER_36_232 ();
 sg13g2_fill_1 FILLER_36_254 ();
 sg13g2_fill_2 FILLER_36_260 ();
 sg13g2_decap_8 FILLER_36_275 ();
 sg13g2_decap_8 FILLER_36_282 ();
 sg13g2_decap_8 FILLER_36_289 ();
 sg13g2_decap_8 FILLER_36_296 ();
 sg13g2_decap_8 FILLER_36_303 ();
 sg13g2_decap_8 FILLER_36_310 ();
 sg13g2_decap_8 FILLER_36_317 ();
 sg13g2_decap_8 FILLER_36_324 ();
 sg13g2_decap_8 FILLER_36_331 ();
 sg13g2_decap_8 FILLER_36_338 ();
 sg13g2_decap_8 FILLER_36_345 ();
 sg13g2_decap_8 FILLER_36_352 ();
 sg13g2_decap_8 FILLER_36_359 ();
 sg13g2_decap_8 FILLER_36_366 ();
 sg13g2_decap_8 FILLER_36_373 ();
 sg13g2_decap_8 FILLER_36_380 ();
 sg13g2_decap_8 FILLER_36_387 ();
 sg13g2_decap_8 FILLER_36_394 ();
 sg13g2_decap_8 FILLER_36_401 ();
 sg13g2_fill_1 FILLER_36_408 ();
 sg13g2_decap_4 FILLER_37_0 ();
 sg13g2_fill_2 FILLER_37_40 ();
 sg13g2_fill_1 FILLER_37_42 ();
 sg13g2_fill_2 FILLER_37_117 ();
 sg13g2_decap_8 FILLER_37_171 ();
 sg13g2_decap_8 FILLER_37_178 ();
 sg13g2_fill_1 FILLER_37_185 ();
 sg13g2_fill_1 FILLER_37_196 ();
 sg13g2_fill_2 FILLER_37_206 ();
 sg13g2_fill_2 FILLER_37_232 ();
 sg13g2_fill_1 FILLER_37_234 ();
 sg13g2_fill_2 FILLER_37_245 ();
 sg13g2_fill_1 FILLER_37_247 ();
 sg13g2_decap_8 FILLER_37_274 ();
 sg13g2_decap_8 FILLER_37_281 ();
 sg13g2_decap_8 FILLER_37_288 ();
 sg13g2_decap_8 FILLER_37_295 ();
 sg13g2_decap_8 FILLER_37_302 ();
 sg13g2_decap_8 FILLER_37_309 ();
 sg13g2_decap_8 FILLER_37_316 ();
 sg13g2_decap_8 FILLER_37_323 ();
 sg13g2_decap_8 FILLER_37_330 ();
 sg13g2_decap_8 FILLER_37_337 ();
 sg13g2_decap_8 FILLER_37_344 ();
 sg13g2_decap_8 FILLER_37_351 ();
 sg13g2_decap_8 FILLER_37_358 ();
 sg13g2_decap_8 FILLER_37_365 ();
 sg13g2_decap_8 FILLER_37_372 ();
 sg13g2_decap_8 FILLER_37_379 ();
 sg13g2_decap_8 FILLER_37_386 ();
 sg13g2_decap_8 FILLER_37_393 ();
 sg13g2_decap_8 FILLER_37_400 ();
 sg13g2_fill_2 FILLER_37_407 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_4 FILLER_38_28 ();
 sg13g2_fill_1 FILLER_38_32 ();
 sg13g2_fill_2 FILLER_38_58 ();
 sg13g2_fill_1 FILLER_38_60 ();
 sg13g2_fill_1 FILLER_38_79 ();
 sg13g2_decap_8 FILLER_38_150 ();
 sg13g2_fill_2 FILLER_38_157 ();
 sg13g2_decap_8 FILLER_38_167 ();
 sg13g2_fill_1 FILLER_38_174 ();
 sg13g2_fill_2 FILLER_38_210 ();
 sg13g2_fill_1 FILLER_38_217 ();
 sg13g2_decap_8 FILLER_38_226 ();
 sg13g2_decap_8 FILLER_38_233 ();
 sg13g2_decap_4 FILLER_38_240 ();
 sg13g2_fill_1 FILLER_38_244 ();
 sg13g2_fill_2 FILLER_38_249 ();
 sg13g2_fill_1 FILLER_38_251 ();
 sg13g2_fill_2 FILLER_38_262 ();
 sg13g2_decap_8 FILLER_38_268 ();
 sg13g2_decap_8 FILLER_38_275 ();
 sg13g2_decap_8 FILLER_38_282 ();
 sg13g2_decap_8 FILLER_38_289 ();
 sg13g2_decap_8 FILLER_38_296 ();
 sg13g2_decap_8 FILLER_38_303 ();
 sg13g2_decap_8 FILLER_38_310 ();
 sg13g2_decap_8 FILLER_38_317 ();
 sg13g2_decap_8 FILLER_38_324 ();
 sg13g2_decap_8 FILLER_38_331 ();
 sg13g2_decap_8 FILLER_38_338 ();
 sg13g2_decap_8 FILLER_38_345 ();
 sg13g2_decap_8 FILLER_38_352 ();
 sg13g2_decap_8 FILLER_38_359 ();
 sg13g2_decap_8 FILLER_38_366 ();
 sg13g2_fill_2 FILLER_38_373 ();
 sg13g2_fill_1 FILLER_38_375 ();
 sg13g2_decap_8 FILLER_38_381 ();
 sg13g2_decap_8 FILLER_38_388 ();
 sg13g2_decap_8 FILLER_38_395 ();
 sg13g2_decap_8 FILLER_38_402 ();
 assign uio_oe[0] = net4;
 assign uio_oe[1] = net5;
 assign uio_oe[2] = net6;
 assign uio_oe[3] = net7;
 assign uio_oe[4] = net8;
 assign uio_oe[5] = net9;
 assign uio_oe[6] = net10;
 assign uio_oe[7] = net11;
 assign uo_out[7] = net2;
endmodule

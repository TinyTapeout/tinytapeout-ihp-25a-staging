module tt_um_lif_tk (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire _297_;
 wire _298_;
 wire _299_;
 wire _300_;
 wire _301_;
 wire _302_;
 wire _303_;
 wire _304_;
 wire _305_;
 wire _306_;
 wire _307_;
 wire _308_;
 wire _309_;
 wire _310_;
 wire _311_;
 wire _312_;
 wire _313_;
 wire _314_;
 wire _315_;
 wire _316_;
 wire _317_;
 wire _318_;
 wire _319_;
 wire _320_;
 wire _321_;
 wire _322_;
 wire _323_;
 wire _324_;
 wire _325_;
 wire _326_;
 wire _327_;
 wire _328_;
 wire _329_;
 wire _330_;
 wire _331_;
 wire _332_;
 wire _333_;
 wire _334_;
 wire _335_;
 wire _336_;
 wire _337_;
 wire _338_;
 wire _339_;
 wire _340_;
 wire _341_;
 wire _342_;
 wire _343_;
 wire _344_;
 wire _345_;
 wire _346_;
 wire _347_;
 wire _348_;
 wire _349_;
 wire _350_;
 wire _351_;
 wire _352_;
 wire _353_;
 wire _354_;
 wire _355_;
 wire _356_;
 wire _357_;
 wire _358_;
 wire _359_;
 wire _360_;
 wire _361_;
 wire _362_;
 wire _363_;
 wire _364_;
 wire _365_;
 wire _366_;
 wire _367_;
 wire _368_;
 wire _369_;
 wire _370_;
 wire _371_;
 wire _372_;
 wire _373_;
 wire _374_;
 wire _375_;
 wire _376_;
 wire _377_;
 wire _378_;
 wire _379_;
 wire _380_;
 wire _381_;
 wire _382_;
 wire _383_;
 wire _384_;
 wire _385_;
 wire _386_;
 wire _387_;
 wire _388_;
 wire _389_;
 wire _390_;
 wire _391_;
 wire _392_;
 wire _393_;
 wire _394_;
 wire _395_;
 wire _396_;
 wire _397_;
 wire _398_;
 wire _399_;
 wire _400_;
 wire _401_;
 wire _402_;
 wire _403_;
 wire _404_;
 wire _405_;
 wire _406_;
 wire _407_;
 wire _408_;
 wire _409_;
 wire _410_;
 wire _411_;
 wire _412_;
 wire _413_;
 wire _414_;
 wire _415_;
 wire _416_;
 wire _417_;
 wire _418_;
 wire _419_;
 wire _420_;
 wire _421_;
 wire _422_;
 wire _423_;
 wire _424_;
 wire _425_;
 wire _426_;
 wire _427_;
 wire _428_;
 wire _429_;
 wire _430_;
 wire _431_;
 wire _432_;
 wire _433_;
 wire _434_;
 wire _435_;
 wire _436_;
 wire _437_;
 wire _438_;
 wire _439_;
 wire _440_;
 wire _441_;
 wire _442_;
 wire _443_;
 wire _444_;
 wire _445_;
 wire _446_;
 wire _447_;
 wire _448_;
 wire _449_;
 wire _450_;
 wire _451_;
 wire _452_;
 wire _453_;
 wire _454_;
 wire _455_;
 wire _456_;
 wire _457_;
 wire _458_;
 wire _459_;
 wire \neuron1.refractory_counter[0] ;
 wire \neuron1.refractory_counter[1] ;
 wire \neuron1.refractory_counter[2] ;
 wire \neuron1.refractory_counter[3] ;
 wire \neuron1.spike ;
 wire \neuron2.membrane_potential[0] ;
 wire \neuron2.membrane_potential[1] ;
 wire \neuron2.membrane_potential[2] ;
 wire \neuron2.membrane_potential[3] ;
 wire \neuron2.membrane_potential[4] ;
 wire \neuron2.membrane_potential[5] ;
 wire \neuron2.membrane_potential[6] ;
 wire \neuron2.membrane_potential[7] ;
 wire \neuron2.phase_counter[0] ;
 wire \neuron2.phase_counter[1] ;
 wire \neuron2.phase_counter[2] ;
 wire \neuron2.phase_counter[3] ;
 wire \neuron2.phase_counter[4] ;
 wire \neuron2.phase_counter[5] ;
 wire \neuron2.phase_counter[6] ;
 wire \neuron2.phase_counter[7] ;
 wire \neuron2.refractory_counter[0] ;
 wire \neuron2.refractory_counter[1] ;
 wire \neuron2.refractory_counter[2] ;
 wire \neuron2.refractory_counter[3] ;
 wire \neuron2.spike ;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire clknet_0_clk;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;

 sg13g2_inv_1 _460_ (.Y(_436_),
    .A(net35));
 sg13g2_inv_1 _461_ (.Y(_437_),
    .A(net50));
 sg13g2_inv_1 _462_ (.Y(_046_),
    .A(\neuron2.membrane_potential[1] ));
 sg13g2_inv_1 _463_ (.Y(_047_),
    .A(net72));
 sg13g2_inv_1 _464_ (.Y(_048_),
    .A(net60));
 sg13g2_inv_1 _465_ (.Y(_049_),
    .A(uio_out[5]));
 sg13g2_inv_1 _466_ (.Y(_050_),
    .A(net82));
 sg13g2_inv_1 _467_ (.Y(_051_),
    .A(net1));
 sg13g2_inv_1 _468_ (.Y(_052_),
    .A(net46));
 sg13g2_inv_1 _469_ (.Y(_053_),
    .A(net118));
 sg13g2_inv_1 _470_ (.Y(_054_),
    .A(net38));
 sg13g2_inv_1 _471_ (.Y(_055_),
    .A(net40));
 sg13g2_mux2_1 _472_ (.A0(\neuron2.phase_counter[0] ),
    .A1(net28),
    .S(net130),
    .X(_012_));
 sg13g2_nand3_1 _473_ (.B(net75),
    .C(net131),
    .A(\neuron2.phase_counter[0] ),
    .Y(_056_));
 sg13g2_a21o_1 _474_ (.A2(net131),
    .A1(\neuron2.phase_counter[0] ),
    .B1(net75),
    .X(_057_));
 sg13g2_and2_1 _475_ (.A(_056_),
    .B(net76),
    .X(_013_));
 sg13g2_nand4_1 _476_ (.B(net44),
    .C(\neuron2.phase_counter[1] ),
    .A(\neuron2.phase_counter[0] ),
    .Y(_058_),
    .D(net130));
 sg13g2_xnor2_1 _477_ (.Y(_014_),
    .A(net44),
    .B(_056_));
 sg13g2_nor2_2 _478_ (.A(_054_),
    .B(_058_),
    .Y(_059_));
 sg13g2_xnor2_1 _479_ (.Y(_015_),
    .A(net38),
    .B(_058_));
 sg13g2_xor2_1 _480_ (.B(_059_),
    .A(net54),
    .X(_016_));
 sg13g2_nand3_1 _481_ (.B(net74),
    .C(_059_),
    .A(net54),
    .Y(_060_));
 sg13g2_a21o_1 _482_ (.A2(_059_),
    .A1(net54),
    .B1(net74),
    .X(_061_));
 sg13g2_and2_1 _483_ (.A(_060_),
    .B(_061_),
    .X(_017_));
 sg13g2_and2_1 _484_ (.A(net36),
    .B(\neuron2.phase_counter[5] ),
    .X(_062_));
 sg13g2_nand3_1 _485_ (.B(_059_),
    .C(_062_),
    .A(\neuron2.phase_counter[4] ),
    .Y(_063_));
 sg13g2_xnor2_1 _486_ (.Y(_018_),
    .A(net36),
    .B(_060_));
 sg13g2_xnor2_1 _487_ (.Y(_019_),
    .A(net42),
    .B(_063_));
 sg13g2_nor2_1 _488_ (.A(\neuron1.refractory_counter[1] ),
    .B(\neuron1.refractory_counter[0] ),
    .Y(_064_));
 sg13g2_nor4_2 _489_ (.A(\neuron1.refractory_counter[1] ),
    .B(net62),
    .C(net46),
    .Y(_065_),
    .D(\neuron1.refractory_counter[2] ));
 sg13g2_or3_1 _490_ (.A(uio_out[3]),
    .B(uio_out[5]),
    .C(uio_out[4]),
    .X(_066_));
 sg13g2_nand3_1 _491_ (.B(uio_out[6]),
    .C(_066_),
    .A(uio_out[7]),
    .Y(_067_));
 sg13g2_and2_1 _492_ (.A(net126),
    .B(_067_),
    .X(_068_));
 sg13g2_nand2_1 _493_ (.Y(_069_),
    .A(net127),
    .B(_067_));
 sg13g2_and2_2 _494_ (.A(_065_),
    .B(_068_),
    .X(_070_));
 sg13g2_nand2_1 _495_ (.Y(_071_),
    .A(_065_),
    .B(_068_));
 sg13g2_nand2b_2 _496_ (.Y(_072_),
    .B(net2),
    .A_N(net3));
 sg13g2_nand2b_1 _497_ (.Y(_073_),
    .B(net1),
    .A_N(net3));
 sg13g2_nor2_2 _498_ (.A(_051_),
    .B(_072_),
    .Y(_074_));
 sg13g2_nand3b_1 _499_ (.B(net1),
    .C(net2),
    .Y(_075_),
    .A_N(net3));
 sg13g2_nand2_2 _500_ (.Y(_076_),
    .A(net7),
    .B(net104));
 sg13g2_nor2_1 _501_ (.A(net111),
    .B(_076_),
    .Y(_077_));
 sg13g2_nand3_1 _502_ (.B(net113),
    .C(net103),
    .A(net4),
    .Y(_078_));
 sg13g2_xnor2_1 _503_ (.Y(_079_),
    .A(net4),
    .B(_077_));
 sg13g2_or2_1 _504_ (.X(_080_),
    .B(_079_),
    .A(_047_));
 sg13g2_xnor2_1 _505_ (.Y(_081_),
    .A(_047_),
    .B(_079_));
 sg13g2_a21oi_1 _506_ (.A1(uio_out[1]),
    .A2(uio_out[2]),
    .Y(_082_),
    .B1(uio_out[7]));
 sg13g2_nor4_1 _507_ (.A(uio_out[3]),
    .B(uio_out[5]),
    .C(uio_out[4]),
    .D(uio_out[6]),
    .Y(_083_));
 sg13g2_and2_1 _508_ (.A(_082_),
    .B(_083_),
    .X(_084_));
 sg13g2_inv_1 _509_ (.Y(_085_),
    .A(_084_));
 sg13g2_xnor2_1 _510_ (.Y(_086_),
    .A(_081_),
    .B(_085_));
 sg13g2_nand2_1 _511_ (.Y(_087_),
    .A(_070_),
    .B(_086_));
 sg13g2_o21ai_1 _512_ (.B1(_087_),
    .Y(_020_),
    .A1(_047_),
    .A2(net127));
 sg13g2_nand2b_1 _513_ (.Y(_088_),
    .B(net31),
    .A_N(net129));
 sg13g2_and2_1 _514_ (.A(net103),
    .B(net112),
    .X(_089_));
 sg13g2_nand2_1 _515_ (.Y(_090_),
    .A(net103),
    .B(net112));
 sg13g2_a21oi_1 _516_ (.A1(net103),
    .A2(net8),
    .Y(_091_),
    .B1(net5));
 sg13g2_nand3_1 _517_ (.B(net120),
    .C(net112),
    .A(net103),
    .Y(_092_));
 sg13g2_nand2b_1 _518_ (.Y(_093_),
    .B(_092_),
    .A_N(_091_));
 sg13g2_xnor2_1 _519_ (.Y(_094_),
    .A(_078_),
    .B(_093_));
 sg13g2_nor2b_1 _520_ (.A(net120),
    .B_N(net111),
    .Y(_095_));
 sg13g2_nor2_1 _521_ (.A(net2),
    .B(_073_),
    .Y(_096_));
 sg13g2_or2_2 _522_ (.X(_097_),
    .B(_073_),
    .A(net2));
 sg13g2_and2_1 _523_ (.A(net103),
    .B(net6),
    .X(_098_));
 sg13g2_nand2_2 _524_ (.Y(_099_),
    .A(net103),
    .B(net6));
 sg13g2_a221oi_1 _525_ (.B2(_098_),
    .C1(_095_),
    .B1(net101),
    .A1(_074_),
    .Y(_100_),
    .A2(_094_));
 sg13g2_nor4_2 _526_ (.A(net2),
    .B(net120),
    .C(_073_),
    .Y(_101_),
    .D(_099_));
 sg13g2_o21ai_1 _527_ (.B1(uio_out[1]),
    .Y(_102_),
    .A1(_100_),
    .A2(_101_));
 sg13g2_nor3_1 _528_ (.A(uio_out[1]),
    .B(_100_),
    .C(_101_),
    .Y(_103_));
 sg13g2_or3_1 _529_ (.A(uio_out[1]),
    .B(_100_),
    .C(_101_),
    .X(_104_));
 sg13g2_nand2_1 _530_ (.Y(_105_),
    .A(_102_),
    .B(_104_));
 sg13g2_xnor2_1 _531_ (.Y(_106_),
    .A(_080_),
    .B(_105_));
 sg13g2_nand2_1 _532_ (.Y(_107_),
    .A(_081_),
    .B(_106_));
 sg13g2_a21oi_1 _533_ (.A1(_081_),
    .A2(_085_),
    .Y(_108_),
    .B1(_106_));
 sg13g2_o21ai_1 _534_ (.B1(_070_),
    .Y(_109_),
    .A1(_084_),
    .A2(_107_));
 sg13g2_o21ai_1 _535_ (.B1(_088_),
    .Y(_021_),
    .A1(_108_),
    .A2(_109_));
 sg13g2_o21ai_1 _536_ (.B1(_102_),
    .Y(_110_),
    .A1(_080_),
    .A2(_103_));
 sg13g2_a21o_1 _537_ (.A2(net104),
    .A1(net113),
    .B1(net119),
    .X(_111_));
 sg13g2_nand3_1 _538_ (.B(net104),
    .C(net119),
    .A(net113),
    .Y(_112_));
 sg13g2_and2_1 _539_ (.A(_111_),
    .B(_112_),
    .X(_113_));
 sg13g2_nand4_1 _540_ (.B(_098_),
    .C(_111_),
    .A(net5),
    .Y(_114_),
    .D(_112_));
 sg13g2_a21o_1 _541_ (.A2(_098_),
    .A1(net120),
    .B1(_113_),
    .X(_115_));
 sg13g2_a21oi_2 _542_ (.B1(_097_),
    .Y(_116_),
    .A2(_115_),
    .A1(_114_));
 sg13g2_o21ai_1 _543_ (.B1(_092_),
    .Y(_117_),
    .A1(_078_),
    .A2(_091_));
 sg13g2_nand2_2 _544_ (.Y(_118_),
    .A(net103),
    .B(net9));
 sg13g2_nor2_1 _545_ (.A(_053_),
    .B(_118_),
    .Y(_119_));
 sg13g2_xnor2_1 _546_ (.Y(_120_),
    .A(net119),
    .B(_118_));
 sg13g2_xnor2_1 _547_ (.Y(_121_),
    .A(_117_),
    .B(_120_));
 sg13g2_and2_1 _548_ (.A(_053_),
    .B(net111),
    .X(_122_));
 sg13g2_nor2_2 _549_ (.A(net1),
    .B(_072_),
    .Y(_123_));
 sg13g2_nand2b_2 _550_ (.Y(_124_),
    .B(_051_),
    .A_N(_072_));
 sg13g2_a221oi_1 _551_ (.B2(_098_),
    .C1(_122_),
    .B1(_123_),
    .A1(_074_),
    .Y(_125_),
    .A2(_121_));
 sg13g2_nor4_1 _552_ (.A(net1),
    .B(net118),
    .C(_072_),
    .D(_099_),
    .Y(_126_));
 sg13g2_nor3_2 _553_ (.A(net101),
    .B(_125_),
    .C(_126_),
    .Y(_127_));
 sg13g2_nor3_1 _554_ (.A(_000_),
    .B(_116_),
    .C(_127_),
    .Y(_128_));
 sg13g2_o21ai_1 _555_ (.B1(_000_),
    .Y(_129_),
    .A1(_116_),
    .A2(_127_));
 sg13g2_nor2b_1 _556_ (.A(_128_),
    .B_N(_129_),
    .Y(_130_));
 sg13g2_xor2_1 _557_ (.B(_130_),
    .A(_110_),
    .X(_131_));
 sg13g2_a21oi_1 _558_ (.A1(_081_),
    .A2(_106_),
    .Y(_132_),
    .B1(_084_));
 sg13g2_a21oi_1 _559_ (.A1(_131_),
    .A2(_132_),
    .Y(_133_),
    .B1(_071_));
 sg13g2_o21ai_1 _560_ (.B1(_133_),
    .Y(_134_),
    .A1(_131_),
    .A2(_132_));
 sg13g2_o21ai_1 _561_ (.B1(_134_),
    .Y(_022_),
    .A1(_048_),
    .A2(net127));
 sg13g2_a21oi_1 _562_ (.A1(_110_),
    .A2(_129_),
    .Y(_135_),
    .B1(_128_));
 sg13g2_a21oi_2 _563_ (.B1(_119_),
    .Y(_136_),
    .A2(_120_),
    .A1(_117_));
 sg13g2_nand2_2 _564_ (.Y(_137_),
    .A(net102),
    .B(net10));
 sg13g2_nand3_1 _565_ (.B(net116),
    .C(net10),
    .A(net102),
    .Y(_138_));
 sg13g2_xor2_1 _566_ (.B(_137_),
    .A(net116),
    .X(_139_));
 sg13g2_xor2_1 _567_ (.B(_139_),
    .A(_136_),
    .X(_140_));
 sg13g2_a21o_1 _568_ (.A2(_072_),
    .A1(net116),
    .B1(_074_),
    .X(_141_));
 sg13g2_o21ai_1 _569_ (.B1(_141_),
    .Y(_142_),
    .A1(net110),
    .A2(_140_));
 sg13g2_nand2_1 _570_ (.Y(_143_),
    .A(net117),
    .B(_076_));
 sg13g2_xor2_1 _571_ (.B(_076_),
    .A(net116),
    .X(_144_));
 sg13g2_o21ai_1 _572_ (.B1(_144_),
    .Y(_145_),
    .A1(net119),
    .A2(_099_));
 sg13g2_nor3_1 _573_ (.A(net118),
    .B(_099_),
    .C(_144_),
    .Y(_146_));
 sg13g2_nor2_1 _574_ (.A(_124_),
    .B(_146_),
    .Y(_147_));
 sg13g2_a21oi_1 _575_ (.A1(_145_),
    .A2(_147_),
    .Y(_148_),
    .B1(net101));
 sg13g2_xnor2_1 _576_ (.Y(_149_),
    .A(net117),
    .B(_089_));
 sg13g2_a21oi_1 _577_ (.A1(_112_),
    .A2(_114_),
    .Y(_150_),
    .B1(_149_));
 sg13g2_nand3_1 _578_ (.B(_114_),
    .C(_149_),
    .A(_112_),
    .Y(_151_));
 sg13g2_nand2b_1 _579_ (.Y(_152_),
    .B(_151_),
    .A_N(_150_));
 sg13g2_a22oi_1 _580_ (.Y(_153_),
    .B1(_152_),
    .B2(net101),
    .A2(_148_),
    .A1(_142_));
 sg13g2_nand2_1 _581_ (.Y(_154_),
    .A(uio_out[3]),
    .B(_153_));
 sg13g2_xnor2_1 _582_ (.Y(_155_),
    .A(uio_out[3]),
    .B(_153_));
 sg13g2_xor2_1 _583_ (.B(_155_),
    .A(_135_),
    .X(_156_));
 sg13g2_a21oi_1 _584_ (.A1(_107_),
    .A2(_131_),
    .Y(_157_),
    .B1(_084_));
 sg13g2_a221oi_1 _585_ (.B2(_131_),
    .C1(_156_),
    .B1(_107_),
    .A1(_082_),
    .Y(_158_),
    .A2(_083_));
 sg13g2_xnor2_1 _586_ (.Y(_159_),
    .A(_156_),
    .B(_157_));
 sg13g2_nand2b_1 _587_ (.Y(_160_),
    .B(net68),
    .A_N(net126));
 sg13g2_o21ai_1 _588_ (.B1(_160_),
    .Y(_023_),
    .A1(_071_),
    .A2(_159_));
 sg13g2_nand2b_1 _589_ (.Y(_161_),
    .B(net30),
    .A_N(net126));
 sg13g2_o21ai_1 _590_ (.B1(_154_),
    .Y(_162_),
    .A1(_135_),
    .A2(_155_));
 sg13g2_nand3_1 _591_ (.B(net9),
    .C(net114),
    .A(net105),
    .Y(_163_));
 sg13g2_xor2_1 _592_ (.B(_118_),
    .A(net114),
    .X(_164_));
 sg13g2_a21oi_1 _593_ (.A1(net116),
    .A2(_089_),
    .Y(_165_),
    .B1(_150_));
 sg13g2_xnor2_1 _594_ (.Y(_166_),
    .A(_164_),
    .B(_165_));
 sg13g2_nand2_2 _595_ (.Y(_167_),
    .A(net102),
    .B(net11));
 sg13g2_nand3_1 _596_ (.B(net114),
    .C(net11),
    .A(net102),
    .Y(_168_));
 sg13g2_xor2_1 _597_ (.B(_167_),
    .A(net114),
    .X(_169_));
 sg13g2_o21ai_1 _598_ (.B1(_138_),
    .Y(_170_),
    .A1(_136_),
    .A2(_139_));
 sg13g2_nand2b_1 _599_ (.Y(_171_),
    .B(_170_),
    .A_N(_169_));
 sg13g2_xnor2_1 _600_ (.Y(_172_),
    .A(_169_),
    .B(_170_));
 sg13g2_a21o_1 _601_ (.A2(_072_),
    .A1(net114),
    .B1(_074_),
    .X(_173_));
 sg13g2_o21ai_1 _602_ (.B1(_173_),
    .Y(_174_),
    .A1(net110),
    .A2(_172_));
 sg13g2_nand2_1 _603_ (.Y(_175_),
    .A(net115),
    .B(_090_));
 sg13g2_xnor2_1 _604_ (.Y(_176_),
    .A(net115),
    .B(_090_));
 sg13g2_a21o_1 _605_ (.A2(_145_),
    .A1(_143_),
    .B1(_176_),
    .X(_177_));
 sg13g2_nand3_1 _606_ (.B(_145_),
    .C(_176_),
    .A(_143_),
    .Y(_178_));
 sg13g2_nand3_1 _607_ (.B(_177_),
    .C(_178_),
    .A(net99),
    .Y(_179_));
 sg13g2_and2_1 _608_ (.A(_097_),
    .B(_179_),
    .X(_180_));
 sg13g2_a22oi_1 _609_ (.Y(_181_),
    .B1(_174_),
    .B2(_180_),
    .A2(_166_),
    .A1(net100));
 sg13g2_and2_1 _610_ (.A(uio_out[4]),
    .B(_181_),
    .X(_182_));
 sg13g2_xor2_1 _611_ (.B(_181_),
    .A(uio_out[4]),
    .X(_183_));
 sg13g2_xnor2_1 _612_ (.Y(_184_),
    .A(_162_),
    .B(_183_));
 sg13g2_and2_1 _613_ (.A(_158_),
    .B(_184_),
    .X(_185_));
 sg13g2_o21ai_1 _614_ (.B1(_070_),
    .Y(_186_),
    .A1(_158_),
    .A2(_184_));
 sg13g2_o21ai_1 _615_ (.B1(_161_),
    .Y(_024_),
    .A1(_185_),
    .A2(_186_));
 sg13g2_nand2b_1 _616_ (.Y(_187_),
    .B(net34),
    .A_N(net126));
 sg13g2_a21oi_1 _617_ (.A1(_162_),
    .A2(_183_),
    .Y(_188_),
    .B1(_182_));
 sg13g2_nand2_1 _618_ (.Y(_189_),
    .A(net102),
    .B(net12));
 sg13g2_nand3_1 _619_ (.B(_171_),
    .C(_189_),
    .A(_168_),
    .Y(_190_));
 sg13g2_a21oi_1 _620_ (.A1(_168_),
    .A2(_171_),
    .Y(_191_),
    .B1(_189_));
 sg13g2_nor2_1 _621_ (.A(net110),
    .B(_191_),
    .Y(_192_));
 sg13g2_nand2_1 _622_ (.Y(_193_),
    .A(_175_),
    .B(_177_));
 sg13g2_and2_1 _623_ (.A(_118_),
    .B(_193_),
    .X(_194_));
 sg13g2_o21ai_1 _624_ (.B1(net99),
    .Y(_195_),
    .A1(_118_),
    .A2(_193_));
 sg13g2_nor2_1 _625_ (.A(_194_),
    .B(_195_),
    .Y(_196_));
 sg13g2_o21ai_1 _626_ (.B1(_163_),
    .Y(_197_),
    .A1(_164_),
    .A2(_165_));
 sg13g2_nand2b_1 _627_ (.Y(_198_),
    .B(_197_),
    .A_N(_137_));
 sg13g2_xnor2_1 _628_ (.Y(_199_),
    .A(_137_),
    .B(_197_));
 sg13g2_a221oi_1 _629_ (.B2(net100),
    .C1(_196_),
    .B1(_199_),
    .A1(_190_),
    .Y(_200_),
    .A2(_192_));
 sg13g2_or2_1 _630_ (.X(_201_),
    .B(_200_),
    .A(_049_));
 sg13g2_and2_1 _631_ (.A(_049_),
    .B(_200_),
    .X(_202_));
 sg13g2_xnor2_1 _632_ (.Y(_203_),
    .A(uio_out[5]),
    .B(_200_));
 sg13g2_xnor2_1 _633_ (.Y(_204_),
    .A(_188_),
    .B(_203_));
 sg13g2_nor2b_1 _634_ (.A(_204_),
    .B_N(_185_),
    .Y(_205_));
 sg13g2_nand2b_1 _635_ (.Y(_206_),
    .B(_204_),
    .A_N(_185_));
 sg13g2_nand2_1 _636_ (.Y(_207_),
    .A(_070_),
    .B(_206_));
 sg13g2_o21ai_1 _637_ (.B1(_187_),
    .Y(_025_),
    .A1(_205_),
    .A2(_207_));
 sg13g2_o21ai_1 _638_ (.B1(_201_),
    .Y(_208_),
    .A1(_188_),
    .A2(_202_));
 sg13g2_nand2_1 _639_ (.Y(_209_),
    .A(_167_),
    .B(_198_));
 sg13g2_nand4_1 _640_ (.B(net10),
    .C(net11),
    .A(net102),
    .Y(_210_),
    .D(_197_));
 sg13g2_nand2_1 _641_ (.Y(_211_),
    .A(net13),
    .B(_191_));
 sg13g2_a21oi_1 _642_ (.A1(net102),
    .A2(net13),
    .Y(_212_),
    .B1(_191_));
 sg13g2_nor2_1 _643_ (.A(net110),
    .B(_212_),
    .Y(_213_));
 sg13g2_nand2_1 _644_ (.Y(_214_),
    .A(_137_),
    .B(_194_));
 sg13g2_nor2_1 _645_ (.A(_137_),
    .B(_194_),
    .Y(_215_));
 sg13g2_nor2_1 _646_ (.A(_124_),
    .B(_215_),
    .Y(_216_));
 sg13g2_and3_1 _647_ (.X(_217_),
    .A(net100),
    .B(_209_),
    .C(_210_));
 sg13g2_a221oi_1 _648_ (.B2(_216_),
    .C1(_217_),
    .B1(_214_),
    .A1(_211_),
    .Y(_218_),
    .A2(_213_));
 sg13g2_nor2_1 _649_ (.A(_050_),
    .B(_218_),
    .Y(_219_));
 sg13g2_nand2_1 _650_ (.Y(_220_),
    .A(_050_),
    .B(_218_));
 sg13g2_xnor2_1 _651_ (.Y(_221_),
    .A(uio_out[6]),
    .B(_218_));
 sg13g2_xnor2_1 _652_ (.Y(_222_),
    .A(_208_),
    .B(_221_));
 sg13g2_and2_1 _653_ (.A(_205_),
    .B(_222_),
    .X(_223_));
 sg13g2_nor2_1 _654_ (.A(_205_),
    .B(_222_),
    .Y(_224_));
 sg13g2_o21ai_1 _655_ (.B1(_070_),
    .Y(_225_),
    .A1(_223_),
    .A2(_224_));
 sg13g2_o21ai_1 _656_ (.B1(_225_),
    .Y(_026_),
    .A1(_050_),
    .A2(net126));
 sg13g2_nand2b_1 _657_ (.Y(_226_),
    .B(net65),
    .A_N(net126));
 sg13g2_a21oi_1 _658_ (.A1(_208_),
    .A2(_220_),
    .Y(_227_),
    .B1(_219_));
 sg13g2_xnor2_1 _659_ (.Y(_228_),
    .A(_167_),
    .B(_214_));
 sg13g2_a21oi_1 _660_ (.A1(net1),
    .A2(_211_),
    .Y(_229_),
    .B1(_072_));
 sg13g2_o21ai_1 _661_ (.B1(_229_),
    .Y(_230_),
    .A1(_124_),
    .A2(_228_));
 sg13g2_a21oi_1 _662_ (.A1(_189_),
    .A2(_210_),
    .Y(_231_),
    .B1(_097_));
 sg13g2_o21ai_1 _663_ (.B1(_231_),
    .Y(_232_),
    .A1(_189_),
    .A2(_210_));
 sg13g2_nand2_1 _664_ (.Y(_233_),
    .A(_230_),
    .B(_232_));
 sg13g2_xor2_1 _665_ (.B(_233_),
    .A(uio_out[7]),
    .X(_234_));
 sg13g2_xnor2_1 _666_ (.Y(_235_),
    .A(_227_),
    .B(_234_));
 sg13g2_and2_1 _667_ (.A(_223_),
    .B(_235_),
    .X(_236_));
 sg13g2_o21ai_1 _668_ (.B1(_070_),
    .Y(_237_),
    .A1(_223_),
    .A2(_235_));
 sg13g2_o21ai_1 _669_ (.B1(_226_),
    .Y(_027_),
    .A1(_236_),
    .A2(_237_));
 sg13g2_o21ai_1 _670_ (.B1(_069_),
    .Y(_238_),
    .A1(net109),
    .A2(net126));
 sg13g2_inv_1 _671_ (.Y(_028_),
    .A(_238_));
 sg13g2_nor2_1 _672_ (.A(_065_),
    .B(_069_),
    .Y(_239_));
 sg13g2_nor2_1 _673_ (.A(net62),
    .B(_239_),
    .Y(_240_));
 sg13g2_a21oi_1 _674_ (.A1(net62),
    .A2(net127),
    .Y(_029_),
    .B1(_240_));
 sg13g2_xor2_1 _675_ (.B(net62),
    .A(net70),
    .X(_241_));
 sg13g2_o21ai_1 _676_ (.B1(_071_),
    .Y(_242_),
    .A1(net70),
    .A2(net126));
 sg13g2_a21oi_1 _677_ (.A1(_068_),
    .A2(_241_),
    .Y(_030_),
    .B1(net71));
 sg13g2_xnor2_1 _678_ (.Y(_243_),
    .A(_001_),
    .B(_064_));
 sg13g2_nor2b_1 _679_ (.A(net127),
    .B_N(net78),
    .Y(_244_));
 sg13g2_a21o_1 _680_ (.A2(_243_),
    .A1(_239_),
    .B1(_244_),
    .X(_031_));
 sg13g2_nand4_1 _681_ (.B(\neuron1.refractory_counter[2] ),
    .C(_001_),
    .A(_052_),
    .Y(_245_),
    .D(_064_));
 sg13g2_nand2_1 _682_ (.Y(_246_),
    .A(_067_),
    .B(_245_));
 sg13g2_nand3_1 _683_ (.B(net127),
    .C(_064_),
    .A(_001_),
    .Y(_247_));
 sg13g2_a22oi_1 _684_ (.Y(_248_),
    .B1(_247_),
    .B2(net46),
    .A2(_246_),
    .A1(net127));
 sg13g2_inv_1 _685_ (.Y(_032_),
    .A(net47));
 sg13g2_nor2_1 _686_ (.A(\neuron2.refractory_counter[0] ),
    .B(\neuron2.refractory_counter[1] ),
    .Y(_249_));
 sg13g2_nor4_2 _687_ (.A(\neuron2.refractory_counter[0] ),
    .B(\neuron2.refractory_counter[1] ),
    .C(net40),
    .Y(_250_),
    .D(net86));
 sg13g2_or3_1 _688_ (.A(\neuron2.membrane_potential[3] ),
    .B(\neuron2.membrane_potential[4] ),
    .C(\neuron2.membrane_potential[5] ),
    .X(_251_));
 sg13g2_nand3_1 _689_ (.B(net56),
    .C(_251_),
    .A(net52),
    .Y(_252_));
 sg13g2_and2_1 _690_ (.A(net129),
    .B(_252_),
    .X(_253_));
 sg13g2_nand2_1 _691_ (.Y(_254_),
    .A(net128),
    .B(_252_));
 sg13g2_and2_1 _692_ (.A(_250_),
    .B(_253_),
    .X(_255_));
 sg13g2_nand2_2 _693_ (.Y(_256_),
    .A(_250_),
    .B(_253_));
 sg13g2_or3_1 _694_ (.A(\neuron2.phase_counter[3] ),
    .B(\neuron2.phase_counter[2] ),
    .C(\neuron2.phase_counter[4] ),
    .X(_257_));
 sg13g2_a21oi_1 _695_ (.A1(_062_),
    .A2(_257_),
    .Y(_258_),
    .B1(\neuron2.phase_counter[7] ));
 sg13g2_a21o_2 _696_ (.A2(_257_),
    .A1(_062_),
    .B1(\neuron2.phase_counter[7] ),
    .X(_259_));
 sg13g2_and2_1 _697_ (.A(net113),
    .B(net107),
    .X(_260_));
 sg13g2_nand2_1 _698_ (.Y(_261_),
    .A(net113),
    .B(net106));
 sg13g2_nor2_1 _699_ (.A(net111),
    .B(_261_),
    .Y(_262_));
 sg13g2_xnor2_1 _700_ (.Y(_263_),
    .A(net4),
    .B(_262_));
 sg13g2_a21oi_2 _701_ (.B1(_263_),
    .Y(_264_),
    .A2(_258_),
    .A1(net99));
 sg13g2_nand2_1 _702_ (.Y(_265_),
    .A(\neuron2.membrane_potential[0] ),
    .B(_264_));
 sg13g2_xnor2_1 _703_ (.Y(_266_),
    .A(\neuron2.membrane_potential[0] ),
    .B(_264_));
 sg13g2_nor2_1 _704_ (.A(_437_),
    .B(_046_),
    .Y(_267_));
 sg13g2_nor4_2 _705_ (.A(\neuron2.membrane_potential[6] ),
    .B(\neuron2.membrane_potential[7] ),
    .C(_251_),
    .Y(_268_),
    .D(_267_));
 sg13g2_inv_1 _706_ (.Y(_269_),
    .A(_268_));
 sg13g2_and2_1 _707_ (.A(_266_),
    .B(_269_),
    .X(_270_));
 sg13g2_xnor2_1 _708_ (.Y(_271_),
    .A(_266_),
    .B(_268_));
 sg13g2_nand2b_1 _709_ (.Y(_272_),
    .B(net48),
    .A_N(net130));
 sg13g2_o21ai_1 _710_ (.B1(_272_),
    .Y(_033_),
    .A1(_256_),
    .A2(_271_));
 sg13g2_nand3_1 _711_ (.B(net113),
    .C(net106),
    .A(net4),
    .Y(_273_));
 sg13g2_nand2_2 _712_ (.Y(_274_),
    .A(net112),
    .B(net107));
 sg13g2_a21oi_1 _713_ (.A1(net112),
    .A2(net107),
    .Y(_275_),
    .B1(net120));
 sg13g2_a21o_1 _714_ (.A2(net106),
    .A1(net112),
    .B1(net120),
    .X(_276_));
 sg13g2_nand3_1 _715_ (.B(net112),
    .C(net106),
    .A(net120),
    .Y(_277_));
 sg13g2_and4_1 _716_ (.A(net4),
    .B(_260_),
    .C(_276_),
    .D(_277_),
    .X(_278_));
 sg13g2_a22oi_1 _717_ (.Y(_279_),
    .B1(_276_),
    .B2(_277_),
    .A2(_260_),
    .A1(net4));
 sg13g2_o21ai_1 _718_ (.B1(_074_),
    .Y(_280_),
    .A1(_278_),
    .A2(_279_));
 sg13g2_a21oi_1 _719_ (.A1(net99),
    .A2(_258_),
    .Y(_281_),
    .B1(_095_));
 sg13g2_nand2_1 _720_ (.Y(_282_),
    .A(net6),
    .B(net106));
 sg13g2_or2_1 _721_ (.X(_283_),
    .B(_282_),
    .A(_097_));
 sg13g2_and3_1 _722_ (.X(_284_),
    .A(_280_),
    .B(_281_),
    .C(_283_));
 sg13g2_a21oi_2 _723_ (.B1(_283_),
    .Y(_285_),
    .A2(_281_),
    .A1(_280_));
 sg13g2_o21ai_1 _724_ (.B1(\neuron2.membrane_potential[1] ),
    .Y(_286_),
    .A1(_284_),
    .A2(_285_));
 sg13g2_nor3_1 _725_ (.A(\neuron2.membrane_potential[1] ),
    .B(_284_),
    .C(_285_),
    .Y(_287_));
 sg13g2_nor3_1 _726_ (.A(_046_),
    .B(_284_),
    .C(_285_),
    .Y(_288_));
 sg13g2_o21ai_1 _727_ (.B1(_046_),
    .Y(_289_),
    .A1(_284_),
    .A2(_285_));
 sg13g2_nor2b_1 _728_ (.A(_288_),
    .B_N(_289_),
    .Y(_290_));
 sg13g2_xnor2_1 _729_ (.Y(_291_),
    .A(_265_),
    .B(_290_));
 sg13g2_nand2_1 _730_ (.Y(_292_),
    .A(_270_),
    .B(_291_));
 sg13g2_o21ai_1 _731_ (.B1(_255_),
    .Y(_293_),
    .A1(_270_),
    .A2(_291_));
 sg13g2_nand2b_1 _732_ (.Y(_294_),
    .B(_292_),
    .A_N(_293_));
 sg13g2_o21ai_1 _733_ (.B1(_294_),
    .Y(_034_),
    .A1(_436_),
    .A2(net130));
 sg13g2_a21oi_1 _734_ (.A1(_266_),
    .A2(_291_),
    .Y(_295_),
    .B1(_268_));
 sg13g2_o21ai_1 _735_ (.B1(_286_),
    .Y(_296_),
    .A1(_265_),
    .A2(_287_));
 sg13g2_a21oi_1 _736_ (.A1(net113),
    .A2(net106),
    .Y(_297_),
    .B1(net118));
 sg13g2_nand3_1 _737_ (.B(net118),
    .C(net106),
    .A(net113),
    .Y(_298_));
 sg13g2_nor2b_1 _738_ (.A(_297_),
    .B_N(_298_),
    .Y(_299_));
 sg13g2_nand3_1 _739_ (.B(net6),
    .C(net106),
    .A(net120),
    .Y(_300_));
 sg13g2_xnor2_1 _740_ (.Y(_301_),
    .A(_299_),
    .B(_300_));
 sg13g2_nor2_1 _741_ (.A(_097_),
    .B(_301_),
    .Y(_302_));
 sg13g2_o21ai_1 _742_ (.B1(_277_),
    .Y(_303_),
    .A1(_273_),
    .A2(_275_));
 sg13g2_and2_1 _743_ (.A(net9),
    .B(net108),
    .X(_304_));
 sg13g2_nand2_2 _744_ (.Y(_305_),
    .A(net9),
    .B(net108));
 sg13g2_nand2_1 _745_ (.Y(_306_),
    .A(_053_),
    .B(_305_));
 sg13g2_nor2_1 _746_ (.A(_053_),
    .B(_305_),
    .Y(_307_));
 sg13g2_xnor2_1 _747_ (.Y(_308_),
    .A(net118),
    .B(_304_));
 sg13g2_xnor2_1 _748_ (.Y(_309_),
    .A(_303_),
    .B(_308_));
 sg13g2_nor2_1 _749_ (.A(_122_),
    .B(_123_),
    .Y(_310_));
 sg13g2_o21ai_1 _750_ (.B1(_310_),
    .Y(_311_),
    .A1(net111),
    .A2(_309_));
 sg13g2_a21oi_2 _751_ (.B1(_282_),
    .Y(_312_),
    .A2(_259_),
    .A1(net118));
 sg13g2_and3_1 _752_ (.X(_313_),
    .A(net118),
    .B(_259_),
    .C(_282_));
 sg13g2_o21ai_1 _753_ (.B1(_123_),
    .Y(_314_),
    .A1(_312_),
    .A2(_313_));
 sg13g2_and3_1 _754_ (.X(_315_),
    .A(_097_),
    .B(_311_),
    .C(_314_));
 sg13g2_o21ai_1 _755_ (.B1(_002_),
    .Y(_316_),
    .A1(_302_),
    .A2(_315_));
 sg13g2_nor3_1 _756_ (.A(_002_),
    .B(_302_),
    .C(_315_),
    .Y(_317_));
 sg13g2_or3_1 _757_ (.A(_002_),
    .B(_302_),
    .C(_315_),
    .X(_318_));
 sg13g2_nand2_1 _758_ (.Y(_319_),
    .A(_316_),
    .B(_318_));
 sg13g2_xnor2_1 _759_ (.Y(_320_),
    .A(_296_),
    .B(_319_));
 sg13g2_a21oi_1 _760_ (.A1(_295_),
    .A2(_320_),
    .Y(_321_),
    .B1(_256_));
 sg13g2_o21ai_1 _761_ (.B1(_321_),
    .Y(_322_),
    .A1(_295_),
    .A2(_320_));
 sg13g2_o21ai_1 _762_ (.B1(_322_),
    .Y(_035_),
    .A1(_437_),
    .A2(net130));
 sg13g2_a21oi_1 _763_ (.A1(_296_),
    .A2(_316_),
    .Y(_323_),
    .B1(_317_));
 sg13g2_nand3_1 _764_ (.B(net116),
    .C(net108),
    .A(net112),
    .Y(_324_));
 sg13g2_xor2_1 _765_ (.B(_274_),
    .A(net117),
    .X(_325_));
 sg13g2_o21ai_1 _766_ (.B1(_298_),
    .Y(_326_),
    .A1(_297_),
    .A2(_300_));
 sg13g2_nand2b_1 _767_ (.Y(_327_),
    .B(_326_),
    .A_N(_325_));
 sg13g2_nand2b_1 _768_ (.Y(_328_),
    .B(_325_),
    .A_N(_326_));
 sg13g2_a21o_1 _769_ (.A2(_328_),
    .A1(_327_),
    .B1(_097_),
    .X(_329_));
 sg13g2_a21oi_1 _770_ (.A1(_303_),
    .A2(_306_),
    .Y(_330_),
    .B1(_307_));
 sg13g2_nand2_2 _771_ (.Y(_331_),
    .A(net10),
    .B(net109));
 sg13g2_a21oi_1 _772_ (.A1(net10),
    .A2(net108),
    .Y(_332_),
    .B1(net116));
 sg13g2_nand3_1 _773_ (.B(net10),
    .C(net108),
    .A(net116),
    .Y(_333_));
 sg13g2_nor2b_1 _774_ (.A(_332_),
    .B_N(_333_),
    .Y(_334_));
 sg13g2_xnor2_1 _775_ (.Y(_335_),
    .A(_330_),
    .B(_334_));
 sg13g2_o21ai_1 _776_ (.B1(_141_),
    .Y(_336_),
    .A1(net110),
    .A2(_335_));
 sg13g2_and3_1 _777_ (.X(_337_),
    .A(net117),
    .B(_259_),
    .C(_261_));
 sg13g2_nand3_1 _778_ (.B(_259_),
    .C(_261_),
    .A(net117),
    .Y(_338_));
 sg13g2_a21oi_1 _779_ (.A1(net117),
    .A2(_259_),
    .Y(_339_),
    .B1(_261_));
 sg13g2_or3_1 _780_ (.A(_312_),
    .B(_337_),
    .C(_339_),
    .X(_340_));
 sg13g2_o21ai_1 _781_ (.B1(_312_),
    .Y(_341_),
    .A1(_337_),
    .A2(_339_));
 sg13g2_nand3_1 _782_ (.B(_340_),
    .C(_341_),
    .A(net99),
    .Y(_342_));
 sg13g2_nand3_1 _783_ (.B(_336_),
    .C(_342_),
    .A(_097_),
    .Y(_343_));
 sg13g2_and3_1 _784_ (.X(_344_),
    .A(\neuron2.membrane_potential[3] ),
    .B(_329_),
    .C(_343_));
 sg13g2_nand3_1 _785_ (.B(_329_),
    .C(_343_),
    .A(\neuron2.membrane_potential[3] ),
    .Y(_345_));
 sg13g2_a21oi_1 _786_ (.A1(_329_),
    .A2(_343_),
    .Y(_346_),
    .B1(\neuron2.membrane_potential[3] ));
 sg13g2_nor2_1 _787_ (.A(_344_),
    .B(_346_),
    .Y(_347_));
 sg13g2_xnor2_1 _788_ (.Y(_348_),
    .A(_323_),
    .B(_347_));
 sg13g2_o21ai_1 _789_ (.B1(_292_),
    .Y(_349_),
    .A1(_268_),
    .A2(_320_));
 sg13g2_nor2b_1 _790_ (.A(_348_),
    .B_N(_349_),
    .Y(_350_));
 sg13g2_xnor2_1 _791_ (.Y(_351_),
    .A(_348_),
    .B(_349_));
 sg13g2_nand2b_1 _792_ (.Y(_352_),
    .B(net58),
    .A_N(net130));
 sg13g2_o21ai_1 _793_ (.B1(_352_),
    .Y(_036_),
    .A1(_256_),
    .A2(_351_));
 sg13g2_nand2b_1 _794_ (.Y(_353_),
    .B(net32),
    .A_N(net130));
 sg13g2_o21ai_1 _795_ (.B1(_345_),
    .Y(_354_),
    .A1(_323_),
    .A2(_346_));
 sg13g2_xnor2_1 _796_ (.Y(_355_),
    .A(net115),
    .B(_304_));
 sg13g2_a21oi_1 _797_ (.A1(_324_),
    .A2(_327_),
    .Y(_356_),
    .B1(_355_));
 sg13g2_nand3_1 _798_ (.B(_327_),
    .C(_355_),
    .A(_324_),
    .Y(_357_));
 sg13g2_nand2b_1 _799_ (.Y(_358_),
    .B(_357_),
    .A_N(_356_));
 sg13g2_nand2_2 _800_ (.Y(_359_),
    .A(net11),
    .B(net109));
 sg13g2_and3_1 _801_ (.X(_360_),
    .A(net114),
    .B(net11),
    .C(net109));
 sg13g2_nand2b_1 _802_ (.Y(_361_),
    .B(_359_),
    .A_N(net114));
 sg13g2_nand2b_1 _803_ (.Y(_362_),
    .B(_361_),
    .A_N(_360_));
 sg13g2_o21ai_1 _804_ (.B1(_333_),
    .Y(_363_),
    .A1(_330_),
    .A2(_332_));
 sg13g2_xnor2_1 _805_ (.Y(_364_),
    .A(_362_),
    .B(_363_));
 sg13g2_o21ai_1 _806_ (.B1(_173_),
    .Y(_365_),
    .A1(net110),
    .A2(_364_));
 sg13g2_o21ai_1 _807_ (.B1(_338_),
    .Y(_366_),
    .A1(_312_),
    .A2(_339_));
 sg13g2_nand2_1 _808_ (.Y(_367_),
    .A(net115),
    .B(_259_));
 sg13g2_nor2b_1 _809_ (.A(_367_),
    .B_N(_274_),
    .Y(_368_));
 sg13g2_xnor2_1 _810_ (.Y(_369_),
    .A(_274_),
    .B(_367_));
 sg13g2_or2_1 _811_ (.X(_370_),
    .B(_369_),
    .A(_366_));
 sg13g2_a21oi_1 _812_ (.A1(_366_),
    .A2(_369_),
    .Y(_371_),
    .B1(_124_));
 sg13g2_a21oi_1 _813_ (.A1(_370_),
    .A2(_371_),
    .Y(_372_),
    .B1(net101));
 sg13g2_a22oi_1 _814_ (.Y(_373_),
    .B1(_365_),
    .B2(_372_),
    .A2(_358_),
    .A1(net100));
 sg13g2_and2_1 _815_ (.A(\neuron2.membrane_potential[4] ),
    .B(_373_),
    .X(_374_));
 sg13g2_xor2_1 _816_ (.B(_373_),
    .A(\neuron2.membrane_potential[4] ),
    .X(_375_));
 sg13g2_xnor2_1 _817_ (.Y(_376_),
    .A(_354_),
    .B(_375_));
 sg13g2_and2_1 _818_ (.A(_350_),
    .B(_376_),
    .X(_377_));
 sg13g2_o21ai_1 _819_ (.B1(_255_),
    .Y(_378_),
    .A1(_350_),
    .A2(_376_));
 sg13g2_o21ai_1 _820_ (.B1(_353_),
    .Y(_037_),
    .A1(_377_),
    .A2(_378_));
 sg13g2_nand2b_1 _821_ (.Y(_379_),
    .B(net33),
    .A_N(net130));
 sg13g2_a21o_1 _822_ (.A2(_375_),
    .A1(_354_),
    .B1(_374_),
    .X(_380_));
 sg13g2_nand2_1 _823_ (.Y(_381_),
    .A(net12),
    .B(net109));
 sg13g2_a21oi_1 _824_ (.A1(_361_),
    .A2(_363_),
    .Y(_382_),
    .B1(_360_));
 sg13g2_nor2_1 _825_ (.A(_381_),
    .B(_382_),
    .Y(_383_));
 sg13g2_a21oi_1 _826_ (.A1(_381_),
    .A2(_382_),
    .Y(_384_),
    .B1(net110));
 sg13g2_nand2b_1 _827_ (.Y(_385_),
    .B(_384_),
    .A_N(_383_));
 sg13g2_a21oi_1 _828_ (.A1(_366_),
    .A2(_369_),
    .Y(_386_),
    .B1(_368_));
 sg13g2_nor2_1 _829_ (.A(_304_),
    .B(_386_),
    .Y(_387_));
 sg13g2_xnor2_1 _830_ (.Y(_388_),
    .A(_305_),
    .B(_386_));
 sg13g2_a21oi_1 _831_ (.A1(net99),
    .A2(_388_),
    .Y(_389_),
    .B1(net100));
 sg13g2_a21oi_1 _832_ (.A1(net114),
    .A2(_304_),
    .Y(_390_),
    .B1(_356_));
 sg13g2_nor2_1 _833_ (.A(_331_),
    .B(_390_),
    .Y(_391_));
 sg13g2_xnor2_1 _834_ (.Y(_392_),
    .A(_331_),
    .B(_390_));
 sg13g2_a22oi_1 _835_ (.Y(_393_),
    .B1(_392_),
    .B2(net100),
    .A2(_389_),
    .A1(_385_));
 sg13g2_and2_1 _836_ (.A(\neuron2.membrane_potential[5] ),
    .B(_393_),
    .X(_394_));
 sg13g2_xor2_1 _837_ (.B(_393_),
    .A(\neuron2.membrane_potential[5] ),
    .X(_395_));
 sg13g2_xnor2_1 _838_ (.Y(_396_),
    .A(_380_),
    .B(_395_));
 sg13g2_and3_1 _839_ (.X(_397_),
    .A(_350_),
    .B(_376_),
    .C(_396_));
 sg13g2_o21ai_1 _840_ (.B1(_255_),
    .Y(_398_),
    .A1(_377_),
    .A2(_396_));
 sg13g2_o21ai_1 _841_ (.B1(_379_),
    .Y(_038_),
    .A1(_397_),
    .A2(_398_));
 sg13g2_a21oi_1 _842_ (.A1(_380_),
    .A2(_395_),
    .Y(_399_),
    .B1(_394_));
 sg13g2_nand2_1 _843_ (.Y(_400_),
    .A(net11),
    .B(_391_));
 sg13g2_mux2_1 _844_ (.A0(_359_),
    .A1(net11),
    .S(_391_),
    .X(_401_));
 sg13g2_inv_1 _845_ (.Y(_402_),
    .A(_401_));
 sg13g2_and2_1 _846_ (.A(_331_),
    .B(_387_),
    .X(_403_));
 sg13g2_xor2_1 _847_ (.B(_387_),
    .A(_331_),
    .X(_404_));
 sg13g2_a21oi_1 _848_ (.A1(net13),
    .A2(net109),
    .Y(_405_),
    .B1(_383_));
 sg13g2_and2_1 _849_ (.A(net13),
    .B(_383_),
    .X(_406_));
 sg13g2_nor3_1 _850_ (.A(net110),
    .B(_405_),
    .C(_406_),
    .Y(_407_));
 sg13g2_a221oi_1 _851_ (.B2(net99),
    .C1(_407_),
    .B1(_404_),
    .A1(net100),
    .Y(_408_),
    .A2(_402_));
 sg13g2_or2_1 _852_ (.X(_409_),
    .B(_408_),
    .A(_003_));
 sg13g2_xnor2_1 _853_ (.Y(_410_),
    .A(_003_),
    .B(_408_));
 sg13g2_xor2_1 _854_ (.B(_410_),
    .A(_399_),
    .X(_411_));
 sg13g2_nor2b_1 _855_ (.A(_411_),
    .B_N(_397_),
    .Y(_412_));
 sg13g2_xnor2_1 _856_ (.Y(_413_),
    .A(_397_),
    .B(_411_));
 sg13g2_nand2b_1 _857_ (.Y(_414_),
    .B(net52),
    .A_N(net128));
 sg13g2_o21ai_1 _858_ (.B1(_414_),
    .Y(_039_),
    .A1(_256_),
    .A2(_413_));
 sg13g2_nand2b_1 _859_ (.Y(_415_),
    .B(net56),
    .A_N(net128));
 sg13g2_o21ai_1 _860_ (.B1(_409_),
    .Y(_416_),
    .A1(_399_),
    .A2(_410_));
 sg13g2_o21ai_1 _861_ (.B1(net99),
    .Y(_417_),
    .A1(_359_),
    .A2(_403_));
 sg13g2_a21oi_1 _862_ (.A1(_359_),
    .A2(_403_),
    .Y(_418_),
    .B1(_417_));
 sg13g2_xor2_1 _863_ (.B(_400_),
    .A(_381_),
    .X(_419_));
 sg13g2_a221oi_1 _864_ (.B2(net100),
    .C1(_418_),
    .B1(_419_),
    .A1(_074_),
    .Y(_420_),
    .A2(_406_));
 sg13g2_xor2_1 _865_ (.B(_420_),
    .A(\neuron2.membrane_potential[7] ),
    .X(_421_));
 sg13g2_xnor2_1 _866_ (.Y(_422_),
    .A(_416_),
    .B(_421_));
 sg13g2_nor2_1 _867_ (.A(_412_),
    .B(_422_),
    .Y(_423_));
 sg13g2_a21o_1 _868_ (.A2(_422_),
    .A1(_412_),
    .B1(_256_),
    .X(_424_));
 sg13g2_o21ai_1 _869_ (.B1(_415_),
    .Y(_040_),
    .A1(_423_),
    .A2(_424_));
 sg13g2_o21ai_1 _870_ (.B1(_254_),
    .Y(_425_),
    .A1(net105),
    .A2(net128));
 sg13g2_inv_1 _871_ (.Y(_041_),
    .A(_425_));
 sg13g2_nor2_1 _872_ (.A(_250_),
    .B(_254_),
    .Y(_426_));
 sg13g2_nor2_1 _873_ (.A(net64),
    .B(_426_),
    .Y(_427_));
 sg13g2_a21oi_1 _874_ (.A1(net64),
    .A2(net128),
    .Y(_042_),
    .B1(_427_));
 sg13g2_xor2_1 _875_ (.B(net66),
    .A(net64),
    .X(_428_));
 sg13g2_o21ai_1 _876_ (.B1(_256_),
    .Y(_429_),
    .A1(net66),
    .A2(net129));
 sg13g2_a21oi_1 _877_ (.A1(_253_),
    .A2(_428_),
    .Y(_043_),
    .B1(net67));
 sg13g2_xnor2_1 _878_ (.Y(_430_),
    .A(_004_),
    .B(_249_));
 sg13g2_nor2b_1 _879_ (.A(net128),
    .B_N(net80),
    .Y(_431_));
 sg13g2_a21o_1 _880_ (.A2(_430_),
    .A1(_426_),
    .B1(_431_),
    .X(_044_));
 sg13g2_nand4_1 _881_ (.B(\neuron2.refractory_counter[2] ),
    .C(_004_),
    .A(_055_),
    .Y(_432_),
    .D(_249_));
 sg13g2_nand2_1 _882_ (.Y(_433_),
    .A(_252_),
    .B(_432_));
 sg13g2_nand3_1 _883_ (.B(net128),
    .C(_249_),
    .A(_004_),
    .Y(_434_));
 sg13g2_a22oi_1 _884_ (.Y(_435_),
    .B1(_434_),
    .B2(net40),
    .A2(_433_),
    .A1(net128));
 sg13g2_inv_1 _885_ (.Y(_045_),
    .A(net41));
 sg13g2_dfrbp_1 _886_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net124),
    .D(net29),
    .Q_N(_005_),
    .Q(\neuron2.phase_counter[0] ));
 sg13g2_dfrbp_1 _887_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net124),
    .D(net77),
    .Q_N(_459_),
    .Q(\neuron2.phase_counter[1] ));
 sg13g2_dfrbp_1 _888_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net124),
    .D(net45),
    .Q_N(_458_),
    .Q(\neuron2.phase_counter[2] ));
 sg13g2_dfrbp_1 _889_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net124),
    .D(net39),
    .Q_N(_457_),
    .Q(\neuron2.phase_counter[3] ));
 sg13g2_dfrbp_1 _890_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net124),
    .D(net55),
    .Q_N(_456_),
    .Q(\neuron2.phase_counter[4] ));
 sg13g2_dfrbp_1 _891_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net125),
    .D(_017_),
    .Q_N(_455_),
    .Q(\neuron2.phase_counter[5] ));
 sg13g2_dfrbp_1 _892_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net125),
    .D(net37),
    .Q_N(_454_),
    .Q(\neuron2.phase_counter[6] ));
 sg13g2_dfrbp_1 _893_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net125),
    .D(net43),
    .Q_N(_453_),
    .Q(\neuron2.phase_counter[7] ));
 sg13g2_dfrbp_1 _894_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net123),
    .D(net73),
    .Q_N(_452_),
    .Q(uio_out[0]));
 sg13g2_dfrbp_1 _895_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net123),
    .D(_021_),
    .Q_N(uio_out[1]),
    .Q(_006_));
 sg13g2_dfrbp_1 _896_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net123),
    .D(net61),
    .Q_N(_000_),
    .Q(uio_out[2]));
 sg13g2_dfrbp_1 _897_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net123),
    .D(net69),
    .Q_N(_451_),
    .Q(uio_out[3]));
 sg13g2_dfrbp_1 _898_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net121),
    .D(_024_),
    .Q_N(uio_out[4]),
    .Q(_007_));
 sg13g2_dfrbp_1 _899_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net121),
    .D(_025_),
    .Q_N(uio_out[5]),
    .Q(_008_));
 sg13g2_dfrbp_1 _900_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net121),
    .D(net83),
    .Q_N(_450_),
    .Q(uio_out[6]));
 sg13g2_dfrbp_1 _901_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net121),
    .D(_027_),
    .Q_N(_449_),
    .Q(uio_out[7]));
 sg13g2_dfrbp_1 _902_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net122),
    .D(_028_),
    .Q_N(_448_),
    .Q(\neuron1.spike ));
 sg13g2_dfrbp_1 _903_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net121),
    .D(net63),
    .Q_N(_447_),
    .Q(\neuron1.refractory_counter[0] ));
 sg13g2_dfrbp_1 _904_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net121),
    .D(_030_),
    .Q_N(_446_),
    .Q(\neuron1.refractory_counter[1] ));
 sg13g2_dfrbp_1 _905_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net121),
    .D(net79),
    .Q_N(_001_),
    .Q(\neuron1.refractory_counter[2] ));
 sg13g2_dfrbp_1 _906_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net121),
    .D(_032_),
    .Q_N(_445_),
    .Q(\neuron1.refractory_counter[3] ));
 sg13g2_dfrbp_1 _907_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net124),
    .D(net49),
    .Q_N(_444_),
    .Q(\neuron2.membrane_potential[0] ));
 sg13g2_dfrbp_1 _908_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net124),
    .D(_034_),
    .Q_N(\neuron2.membrane_potential[1] ),
    .Q(_009_));
 sg13g2_dfrbp_1 _909_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net124),
    .D(net51),
    .Q_N(_002_),
    .Q(\neuron2.membrane_potential[2] ));
 sg13g2_dfrbp_1 _910_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net125),
    .D(net59),
    .Q_N(_443_),
    .Q(\neuron2.membrane_potential[3] ));
 sg13g2_dfrbp_1 _911_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net125),
    .D(_037_),
    .Q_N(\neuron2.membrane_potential[4] ),
    .Q(_010_));
 sg13g2_dfrbp_1 _912_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net125),
    .D(_038_),
    .Q_N(\neuron2.membrane_potential[5] ),
    .Q(_011_));
 sg13g2_dfrbp_1 _913_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net122),
    .D(net53),
    .Q_N(_003_),
    .Q(\neuron2.membrane_potential[6] ));
 sg13g2_dfrbp_1 _914_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net122),
    .D(net57),
    .Q_N(_442_),
    .Q(\neuron2.membrane_potential[7] ));
 sg13g2_dfrbp_1 _915_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net122),
    .D(_041_),
    .Q_N(_441_),
    .Q(\neuron2.spike ));
 sg13g2_dfrbp_1 _916_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net122),
    .D(_042_),
    .Q_N(_440_),
    .Q(\neuron2.refractory_counter[0] ));
 sg13g2_dfrbp_1 _917_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net122),
    .D(_043_),
    .Q_N(_439_),
    .Q(\neuron2.refractory_counter[1] ));
 sg13g2_dfrbp_1 _918_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net122),
    .D(net81),
    .Q_N(_004_),
    .Q(\neuron2.refractory_counter[2] ));
 sg13g2_dfrbp_1 _919_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net122),
    .D(_045_),
    .Q_N(_438_),
    .Q(\neuron2.refractory_counter[3] ));
 sg13g2_tielo tt_um_lif_tk_15 (.L_LO(net15));
 sg13g2_tielo tt_um_lif_tk_16 (.L_LO(net16));
 sg13g2_tielo tt_um_lif_tk_17 (.L_LO(net17));
 sg13g2_tielo tt_um_lif_tk_18 (.L_LO(net18));
 sg13g2_tielo tt_um_lif_tk_19 (.L_LO(net19));
 sg13g2_tielo tt_um_lif_tk_20 (.L_LO(net20));
 sg13g2_tielo tt_um_lif_tk_21 (.L_LO(net21));
 sg13g2_tielo tt_um_lif_tk_22 (.L_LO(net22));
 sg13g2_tielo tt_um_lif_tk_23 (.L_LO(net23));
 sg13g2_tielo tt_um_lif_tk_24 (.L_LO(net24));
 sg13g2_tielo tt_um_lif_tk_25 (.L_LO(net25));
 sg13g2_tielo tt_um_lif_tk_26 (.L_LO(net26));
 sg13g2_tielo tt_um_lif_tk_27 (.L_LO(net27));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_1 _934_ (.A(net109),
    .X(uo_out[0]));
 sg13g2_buf_1 _935_ (.A(net102),
    .X(uo_out[1]));
 sg13g2_buf_4 fanout99 (.X(net99),
    .A(_123_));
 sg13g2_buf_2 fanout100 (.A(_096_),
    .X(net100));
 sg13g2_buf_2 fanout101 (.A(_096_),
    .X(net101));
 sg13g2_buf_2 fanout102 (.A(net105),
    .X(net102));
 sg13g2_buf_2 fanout103 (.A(net104),
    .X(net103));
 sg13g2_buf_1 fanout104 (.A(net105),
    .X(net104));
 sg13g2_buf_2 fanout105 (.A(net84),
    .X(net105));
 sg13g2_buf_2 fanout106 (.A(net107),
    .X(net106));
 sg13g2_buf_1 fanout107 (.A(net108),
    .X(net107));
 sg13g2_buf_2 fanout108 (.A(net109),
    .X(net108));
 sg13g2_buf_2 fanout109 (.A(net85),
    .X(net109));
 sg13g2_buf_2 fanout110 (.A(_075_),
    .X(net110));
 sg13g2_buf_1 fanout111 (.A(_075_),
    .X(net111));
 sg13g2_buf_2 fanout112 (.A(net8),
    .X(net112));
 sg13g2_buf_2 fanout113 (.A(net7),
    .X(net113));
 sg13g2_buf_2 fanout114 (.A(ui_in[7]),
    .X(net114));
 sg13g2_buf_2 fanout115 (.A(ui_in[7]),
    .X(net115));
 sg13g2_buf_2 fanout116 (.A(ui_in[6]),
    .X(net116));
 sg13g2_buf_2 fanout117 (.A(ui_in[6]),
    .X(net117));
 sg13g2_buf_2 fanout118 (.A(ui_in[5]),
    .X(net118));
 sg13g2_buf_1 fanout119 (.A(ui_in[5]),
    .X(net119));
 sg13g2_buf_2 fanout120 (.A(net5),
    .X(net120));
 sg13g2_buf_4 fanout121 (.X(net121),
    .A(net123));
 sg13g2_buf_4 fanout122 (.X(net122),
    .A(net123));
 sg13g2_buf_4 fanout123 (.X(net123),
    .A(rst_n));
 sg13g2_buf_4 fanout124 (.X(net124),
    .A(net125));
 sg13g2_buf_4 fanout125 (.X(net125),
    .A(rst_n));
 sg13g2_buf_2 fanout126 (.A(net127),
    .X(net126));
 sg13g2_buf_2 fanout127 (.A(net131),
    .X(net127));
 sg13g2_buf_2 fanout128 (.A(net129),
    .X(net128));
 sg13g2_buf_1 fanout129 (.A(net131),
    .X(net129));
 sg13g2_buf_2 fanout130 (.A(net131),
    .X(net130));
 sg13g2_buf_2 fanout131 (.A(ena),
    .X(net131));
 sg13g2_buf_2 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_2 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_2 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_buf_2 input6 (.A(uio_in[0]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(uio_in[1]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(uio_in[2]),
    .X(net8));
 sg13g2_buf_2 input9 (.A(uio_in[3]),
    .X(net9));
 sg13g2_buf_2 input10 (.A(uio_in[4]),
    .X(net10));
 sg13g2_buf_2 input11 (.A(uio_in[5]),
    .X(net11));
 sg13g2_buf_1 input12 (.A(uio_in[6]),
    .X(net12));
 sg13g2_buf_1 input13 (.A(uio_in[7]),
    .X(net13));
 sg13g2_tielo tt_um_lif_tk_14 (.L_LO(net14));
 sg13g2_buf_2 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sg13g2_buf_2 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sg13g2_buf_2 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sg13g2_buf_2 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sg13g2_buf_2 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sg13g2_buf_2 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sg13g2_buf_2 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sg13g2_buf_2 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_3_1__leaf_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_3_2__leaf_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_3_3__leaf_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_3_5__leaf_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_3_6__leaf_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_3_7__leaf_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(_005_),
    .X(net28));
 sg13g2_dlygate4sd3_1 hold2 (.A(_012_),
    .X(net29));
 sg13g2_dlygate4sd3_1 hold3 (.A(_007_),
    .X(net30));
 sg13g2_dlygate4sd3_1 hold4 (.A(_006_),
    .X(net31));
 sg13g2_dlygate4sd3_1 hold5 (.A(_010_),
    .X(net32));
 sg13g2_dlygate4sd3_1 hold6 (.A(_011_),
    .X(net33));
 sg13g2_dlygate4sd3_1 hold7 (.A(_008_),
    .X(net34));
 sg13g2_dlygate4sd3_1 hold8 (.A(_009_),
    .X(net35));
 sg13g2_dlygate4sd3_1 hold9 (.A(\neuron2.phase_counter[6] ),
    .X(net36));
 sg13g2_dlygate4sd3_1 hold10 (.A(_018_),
    .X(net37));
 sg13g2_dlygate4sd3_1 hold11 (.A(\neuron2.phase_counter[3] ),
    .X(net38));
 sg13g2_dlygate4sd3_1 hold12 (.A(_015_),
    .X(net39));
 sg13g2_dlygate4sd3_1 hold13 (.A(\neuron2.refractory_counter[3] ),
    .X(net40));
 sg13g2_dlygate4sd3_1 hold14 (.A(_435_),
    .X(net41));
 sg13g2_dlygate4sd3_1 hold15 (.A(\neuron2.phase_counter[7] ),
    .X(net42));
 sg13g2_dlygate4sd3_1 hold16 (.A(_019_),
    .X(net43));
 sg13g2_dlygate4sd3_1 hold17 (.A(\neuron2.phase_counter[2] ),
    .X(net44));
 sg13g2_dlygate4sd3_1 hold18 (.A(_014_),
    .X(net45));
 sg13g2_dlygate4sd3_1 hold19 (.A(\neuron1.refractory_counter[3] ),
    .X(net46));
 sg13g2_dlygate4sd3_1 hold20 (.A(_248_),
    .X(net47));
 sg13g2_dlygate4sd3_1 hold21 (.A(\neuron2.membrane_potential[0] ),
    .X(net48));
 sg13g2_dlygate4sd3_1 hold22 (.A(_033_),
    .X(net49));
 sg13g2_dlygate4sd3_1 hold23 (.A(\neuron2.membrane_potential[2] ),
    .X(net50));
 sg13g2_dlygate4sd3_1 hold24 (.A(_035_),
    .X(net51));
 sg13g2_dlygate4sd3_1 hold25 (.A(\neuron2.membrane_potential[6] ),
    .X(net52));
 sg13g2_dlygate4sd3_1 hold26 (.A(_039_),
    .X(net53));
 sg13g2_dlygate4sd3_1 hold27 (.A(\neuron2.phase_counter[4] ),
    .X(net54));
 sg13g2_dlygate4sd3_1 hold28 (.A(_016_),
    .X(net55));
 sg13g2_dlygate4sd3_1 hold29 (.A(\neuron2.membrane_potential[7] ),
    .X(net56));
 sg13g2_dlygate4sd3_1 hold30 (.A(_040_),
    .X(net57));
 sg13g2_dlygate4sd3_1 hold31 (.A(\neuron2.membrane_potential[3] ),
    .X(net58));
 sg13g2_dlygate4sd3_1 hold32 (.A(_036_),
    .X(net59));
 sg13g2_dlygate4sd3_1 hold33 (.A(uio_out[2]),
    .X(net60));
 sg13g2_dlygate4sd3_1 hold34 (.A(_022_),
    .X(net61));
 sg13g2_dlygate4sd3_1 hold35 (.A(\neuron1.refractory_counter[0] ),
    .X(net62));
 sg13g2_dlygate4sd3_1 hold36 (.A(_029_),
    .X(net63));
 sg13g2_dlygate4sd3_1 hold37 (.A(\neuron2.refractory_counter[0] ),
    .X(net64));
 sg13g2_dlygate4sd3_1 hold38 (.A(uio_out[7]),
    .X(net65));
 sg13g2_dlygate4sd3_1 hold39 (.A(\neuron2.refractory_counter[1] ),
    .X(net66));
 sg13g2_dlygate4sd3_1 hold40 (.A(_429_),
    .X(net67));
 sg13g2_dlygate4sd3_1 hold41 (.A(uio_out[3]),
    .X(net68));
 sg13g2_dlygate4sd3_1 hold42 (.A(_023_),
    .X(net69));
 sg13g2_dlygate4sd3_1 hold43 (.A(\neuron1.refractory_counter[1] ),
    .X(net70));
 sg13g2_dlygate4sd3_1 hold44 (.A(_242_),
    .X(net71));
 sg13g2_dlygate4sd3_1 hold45 (.A(uio_out[0]),
    .X(net72));
 sg13g2_dlygate4sd3_1 hold46 (.A(_020_),
    .X(net73));
 sg13g2_dlygate4sd3_1 hold47 (.A(\neuron2.phase_counter[5] ),
    .X(net74));
 sg13g2_dlygate4sd3_1 hold48 (.A(\neuron2.phase_counter[1] ),
    .X(net75));
 sg13g2_dlygate4sd3_1 hold49 (.A(_057_),
    .X(net76));
 sg13g2_dlygate4sd3_1 hold50 (.A(_013_),
    .X(net77));
 sg13g2_dlygate4sd3_1 hold51 (.A(\neuron1.refractory_counter[2] ),
    .X(net78));
 sg13g2_dlygate4sd3_1 hold52 (.A(_031_),
    .X(net79));
 sg13g2_dlygate4sd3_1 hold53 (.A(\neuron2.refractory_counter[2] ),
    .X(net80));
 sg13g2_dlygate4sd3_1 hold54 (.A(_044_),
    .X(net81));
 sg13g2_dlygate4sd3_1 hold55 (.A(uio_out[6]),
    .X(net82));
 sg13g2_dlygate4sd3_1 hold56 (.A(_026_),
    .X(net83));
 sg13g2_dlygate4sd3_1 hold57 (.A(\neuron2.spike ),
    .X(net84));
 sg13g2_dlygate4sd3_1 hold58 (.A(\neuron1.spike ),
    .X(net85));
 sg13g2_dlygate4sd3_1 hold59 (.A(\neuron2.refractory_counter[2] ),
    .X(net86));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_fill_2 FILLER_14_406 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_252 ();
 sg13g2_decap_8 FILLER_15_259 ();
 sg13g2_decap_8 FILLER_15_266 ();
 sg13g2_decap_8 FILLER_15_273 ();
 sg13g2_decap_8 FILLER_15_280 ();
 sg13g2_decap_8 FILLER_15_287 ();
 sg13g2_decap_8 FILLER_15_294 ();
 sg13g2_decap_8 FILLER_15_301 ();
 sg13g2_decap_8 FILLER_15_308 ();
 sg13g2_decap_8 FILLER_15_315 ();
 sg13g2_decap_8 FILLER_15_322 ();
 sg13g2_decap_8 FILLER_15_329 ();
 sg13g2_decap_8 FILLER_15_336 ();
 sg13g2_decap_8 FILLER_15_343 ();
 sg13g2_decap_8 FILLER_15_350 ();
 sg13g2_decap_8 FILLER_15_357 ();
 sg13g2_decap_8 FILLER_15_364 ();
 sg13g2_decap_8 FILLER_15_371 ();
 sg13g2_decap_8 FILLER_15_378 ();
 sg13g2_decap_8 FILLER_15_385 ();
 sg13g2_decap_8 FILLER_15_392 ();
 sg13g2_decap_8 FILLER_15_399 ();
 sg13g2_fill_2 FILLER_15_406 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_decap_8 FILLER_16_217 ();
 sg13g2_decap_8 FILLER_16_224 ();
 sg13g2_decap_8 FILLER_16_231 ();
 sg13g2_decap_8 FILLER_16_238 ();
 sg13g2_decap_8 FILLER_16_245 ();
 sg13g2_decap_8 FILLER_16_252 ();
 sg13g2_decap_8 FILLER_16_259 ();
 sg13g2_decap_8 FILLER_16_266 ();
 sg13g2_decap_8 FILLER_16_273 ();
 sg13g2_decap_8 FILLER_16_280 ();
 sg13g2_decap_8 FILLER_16_287 ();
 sg13g2_decap_8 FILLER_16_294 ();
 sg13g2_decap_8 FILLER_16_301 ();
 sg13g2_decap_8 FILLER_16_308 ();
 sg13g2_decap_8 FILLER_16_315 ();
 sg13g2_decap_8 FILLER_16_322 ();
 sg13g2_decap_8 FILLER_16_329 ();
 sg13g2_decap_8 FILLER_16_336 ();
 sg13g2_decap_8 FILLER_16_343 ();
 sg13g2_decap_8 FILLER_16_350 ();
 sg13g2_decap_8 FILLER_16_357 ();
 sg13g2_decap_8 FILLER_16_364 ();
 sg13g2_decap_8 FILLER_16_371 ();
 sg13g2_decap_8 FILLER_16_378 ();
 sg13g2_decap_8 FILLER_16_385 ();
 sg13g2_decap_8 FILLER_16_392 ();
 sg13g2_decap_8 FILLER_16_399 ();
 sg13g2_fill_2 FILLER_16_406 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_decap_8 FILLER_17_168 ();
 sg13g2_decap_8 FILLER_17_175 ();
 sg13g2_decap_8 FILLER_17_182 ();
 sg13g2_decap_8 FILLER_17_189 ();
 sg13g2_decap_8 FILLER_17_196 ();
 sg13g2_decap_8 FILLER_17_203 ();
 sg13g2_decap_8 FILLER_17_210 ();
 sg13g2_decap_8 FILLER_17_217 ();
 sg13g2_decap_8 FILLER_17_224 ();
 sg13g2_decap_8 FILLER_17_231 ();
 sg13g2_decap_8 FILLER_17_238 ();
 sg13g2_decap_8 FILLER_17_245 ();
 sg13g2_decap_8 FILLER_17_252 ();
 sg13g2_decap_8 FILLER_17_259 ();
 sg13g2_decap_8 FILLER_17_266 ();
 sg13g2_decap_8 FILLER_17_273 ();
 sg13g2_decap_8 FILLER_17_280 ();
 sg13g2_decap_8 FILLER_17_287 ();
 sg13g2_decap_8 FILLER_17_294 ();
 sg13g2_decap_8 FILLER_17_301 ();
 sg13g2_decap_8 FILLER_17_308 ();
 sg13g2_decap_8 FILLER_17_315 ();
 sg13g2_decap_8 FILLER_17_322 ();
 sg13g2_decap_8 FILLER_17_329 ();
 sg13g2_decap_8 FILLER_17_336 ();
 sg13g2_decap_8 FILLER_17_343 ();
 sg13g2_decap_8 FILLER_17_350 ();
 sg13g2_decap_8 FILLER_17_357 ();
 sg13g2_decap_8 FILLER_17_364 ();
 sg13g2_decap_8 FILLER_17_371 ();
 sg13g2_decap_8 FILLER_17_378 ();
 sg13g2_decap_8 FILLER_17_385 ();
 sg13g2_decap_8 FILLER_17_392 ();
 sg13g2_decap_8 FILLER_17_399 ();
 sg13g2_fill_2 FILLER_17_406 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_decap_8 FILLER_18_147 ();
 sg13g2_decap_8 FILLER_18_154 ();
 sg13g2_decap_8 FILLER_18_161 ();
 sg13g2_decap_8 FILLER_18_168 ();
 sg13g2_decap_8 FILLER_18_175 ();
 sg13g2_decap_8 FILLER_18_182 ();
 sg13g2_decap_8 FILLER_18_189 ();
 sg13g2_decap_8 FILLER_18_196 ();
 sg13g2_decap_8 FILLER_18_203 ();
 sg13g2_decap_8 FILLER_18_210 ();
 sg13g2_decap_8 FILLER_18_217 ();
 sg13g2_decap_8 FILLER_18_224 ();
 sg13g2_decap_8 FILLER_18_231 ();
 sg13g2_decap_8 FILLER_18_238 ();
 sg13g2_decap_8 FILLER_18_245 ();
 sg13g2_decap_8 FILLER_18_252 ();
 sg13g2_decap_8 FILLER_18_259 ();
 sg13g2_decap_8 FILLER_18_266 ();
 sg13g2_decap_8 FILLER_18_273 ();
 sg13g2_decap_8 FILLER_18_280 ();
 sg13g2_decap_8 FILLER_18_287 ();
 sg13g2_decap_8 FILLER_18_294 ();
 sg13g2_decap_8 FILLER_18_301 ();
 sg13g2_decap_8 FILLER_18_308 ();
 sg13g2_decap_8 FILLER_18_315 ();
 sg13g2_decap_8 FILLER_18_322 ();
 sg13g2_decap_8 FILLER_18_329 ();
 sg13g2_decap_8 FILLER_18_336 ();
 sg13g2_decap_8 FILLER_18_343 ();
 sg13g2_decap_8 FILLER_18_350 ();
 sg13g2_decap_8 FILLER_18_357 ();
 sg13g2_decap_8 FILLER_18_364 ();
 sg13g2_decap_8 FILLER_18_371 ();
 sg13g2_decap_8 FILLER_18_378 ();
 sg13g2_decap_8 FILLER_18_385 ();
 sg13g2_decap_8 FILLER_18_392 ();
 sg13g2_decap_8 FILLER_18_399 ();
 sg13g2_fill_2 FILLER_18_406 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_decap_8 FILLER_19_140 ();
 sg13g2_decap_8 FILLER_19_147 ();
 sg13g2_decap_8 FILLER_19_154 ();
 sg13g2_decap_8 FILLER_19_161 ();
 sg13g2_decap_8 FILLER_19_168 ();
 sg13g2_decap_8 FILLER_19_175 ();
 sg13g2_decap_8 FILLER_19_182 ();
 sg13g2_decap_8 FILLER_19_189 ();
 sg13g2_decap_8 FILLER_19_196 ();
 sg13g2_decap_8 FILLER_19_203 ();
 sg13g2_decap_8 FILLER_19_210 ();
 sg13g2_decap_8 FILLER_19_217 ();
 sg13g2_decap_8 FILLER_19_224 ();
 sg13g2_decap_8 FILLER_19_231 ();
 sg13g2_decap_8 FILLER_19_238 ();
 sg13g2_decap_8 FILLER_19_245 ();
 sg13g2_decap_8 FILLER_19_252 ();
 sg13g2_decap_8 FILLER_19_259 ();
 sg13g2_decap_8 FILLER_19_266 ();
 sg13g2_decap_8 FILLER_19_273 ();
 sg13g2_decap_8 FILLER_19_280 ();
 sg13g2_decap_8 FILLER_19_287 ();
 sg13g2_decap_8 FILLER_19_294 ();
 sg13g2_decap_8 FILLER_19_301 ();
 sg13g2_decap_8 FILLER_19_308 ();
 sg13g2_decap_8 FILLER_19_315 ();
 sg13g2_decap_8 FILLER_19_322 ();
 sg13g2_decap_8 FILLER_19_329 ();
 sg13g2_decap_8 FILLER_19_336 ();
 sg13g2_decap_8 FILLER_19_343 ();
 sg13g2_decap_8 FILLER_19_350 ();
 sg13g2_decap_8 FILLER_19_357 ();
 sg13g2_decap_8 FILLER_19_364 ();
 sg13g2_decap_8 FILLER_19_371 ();
 sg13g2_decap_8 FILLER_19_378 ();
 sg13g2_decap_8 FILLER_19_385 ();
 sg13g2_decap_8 FILLER_19_392 ();
 sg13g2_decap_8 FILLER_19_399 ();
 sg13g2_fill_2 FILLER_19_406 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_decap_8 FILLER_20_126 ();
 sg13g2_decap_8 FILLER_20_133 ();
 sg13g2_decap_8 FILLER_20_140 ();
 sg13g2_decap_8 FILLER_20_147 ();
 sg13g2_decap_8 FILLER_20_154 ();
 sg13g2_decap_8 FILLER_20_161 ();
 sg13g2_decap_8 FILLER_20_168 ();
 sg13g2_decap_8 FILLER_20_175 ();
 sg13g2_decap_8 FILLER_20_182 ();
 sg13g2_decap_8 FILLER_20_189 ();
 sg13g2_decap_8 FILLER_20_196 ();
 sg13g2_decap_8 FILLER_20_203 ();
 sg13g2_decap_8 FILLER_20_210 ();
 sg13g2_decap_8 FILLER_20_217 ();
 sg13g2_decap_8 FILLER_20_224 ();
 sg13g2_decap_8 FILLER_20_231 ();
 sg13g2_decap_8 FILLER_20_238 ();
 sg13g2_decap_8 FILLER_20_245 ();
 sg13g2_decap_8 FILLER_20_252 ();
 sg13g2_decap_8 FILLER_20_259 ();
 sg13g2_decap_8 FILLER_20_266 ();
 sg13g2_decap_8 FILLER_20_273 ();
 sg13g2_decap_8 FILLER_20_280 ();
 sg13g2_decap_8 FILLER_20_287 ();
 sg13g2_decap_8 FILLER_20_294 ();
 sg13g2_decap_8 FILLER_20_301 ();
 sg13g2_decap_8 FILLER_20_308 ();
 sg13g2_decap_8 FILLER_20_315 ();
 sg13g2_decap_8 FILLER_20_322 ();
 sg13g2_decap_8 FILLER_20_329 ();
 sg13g2_decap_8 FILLER_20_336 ();
 sg13g2_decap_8 FILLER_20_343 ();
 sg13g2_decap_8 FILLER_20_350 ();
 sg13g2_decap_8 FILLER_20_357 ();
 sg13g2_decap_8 FILLER_20_364 ();
 sg13g2_decap_8 FILLER_20_371 ();
 sg13g2_decap_8 FILLER_20_378 ();
 sg13g2_decap_8 FILLER_20_385 ();
 sg13g2_decap_8 FILLER_20_392 ();
 sg13g2_decap_8 FILLER_20_399 ();
 sg13g2_fill_2 FILLER_20_406 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_decap_8 FILLER_21_119 ();
 sg13g2_decap_8 FILLER_21_126 ();
 sg13g2_decap_8 FILLER_21_133 ();
 sg13g2_decap_8 FILLER_21_140 ();
 sg13g2_decap_8 FILLER_21_147 ();
 sg13g2_decap_8 FILLER_21_154 ();
 sg13g2_decap_8 FILLER_21_161 ();
 sg13g2_decap_8 FILLER_21_168 ();
 sg13g2_decap_8 FILLER_21_175 ();
 sg13g2_decap_8 FILLER_21_182 ();
 sg13g2_decap_8 FILLER_21_189 ();
 sg13g2_decap_8 FILLER_21_196 ();
 sg13g2_decap_8 FILLER_21_203 ();
 sg13g2_decap_8 FILLER_21_210 ();
 sg13g2_decap_8 FILLER_21_217 ();
 sg13g2_decap_8 FILLER_21_224 ();
 sg13g2_decap_8 FILLER_21_231 ();
 sg13g2_decap_8 FILLER_21_238 ();
 sg13g2_decap_8 FILLER_21_245 ();
 sg13g2_decap_8 FILLER_21_252 ();
 sg13g2_decap_8 FILLER_21_259 ();
 sg13g2_decap_8 FILLER_21_266 ();
 sg13g2_decap_8 FILLER_21_273 ();
 sg13g2_decap_8 FILLER_21_280 ();
 sg13g2_decap_8 FILLER_21_287 ();
 sg13g2_decap_8 FILLER_21_294 ();
 sg13g2_decap_8 FILLER_21_301 ();
 sg13g2_fill_1 FILLER_21_308 ();
 sg13g2_decap_8 FILLER_21_313 ();
 sg13g2_decap_8 FILLER_21_320 ();
 sg13g2_decap_8 FILLER_21_327 ();
 sg13g2_decap_8 FILLER_21_334 ();
 sg13g2_decap_8 FILLER_21_341 ();
 sg13g2_decap_8 FILLER_21_348 ();
 sg13g2_decap_8 FILLER_21_355 ();
 sg13g2_fill_1 FILLER_21_362 ();
 sg13g2_fill_2 FILLER_21_373 ();
 sg13g2_fill_1 FILLER_21_375 ();
 sg13g2_fill_2 FILLER_21_387 ();
 sg13g2_fill_1 FILLER_21_389 ();
 sg13g2_decap_8 FILLER_21_398 ();
 sg13g2_decap_4 FILLER_21_405 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_8 FILLER_22_105 ();
 sg13g2_decap_8 FILLER_22_112 ();
 sg13g2_decap_8 FILLER_22_119 ();
 sg13g2_decap_8 FILLER_22_126 ();
 sg13g2_decap_8 FILLER_22_133 ();
 sg13g2_decap_8 FILLER_22_140 ();
 sg13g2_decap_8 FILLER_22_147 ();
 sg13g2_decap_8 FILLER_22_154 ();
 sg13g2_decap_4 FILLER_22_161 ();
 sg13g2_fill_1 FILLER_22_165 ();
 sg13g2_decap_8 FILLER_22_171 ();
 sg13g2_decap_8 FILLER_22_178 ();
 sg13g2_decap_8 FILLER_22_185 ();
 sg13g2_decap_8 FILLER_22_192 ();
 sg13g2_decap_8 FILLER_22_209 ();
 sg13g2_decap_8 FILLER_22_216 ();
 sg13g2_decap_8 FILLER_22_223 ();
 sg13g2_decap_8 FILLER_22_230 ();
 sg13g2_fill_2 FILLER_22_237 ();
 sg13g2_decap_4 FILLER_22_269 ();
 sg13g2_decap_4 FILLER_22_299 ();
 sg13g2_decap_8 FILLER_22_333 ();
 sg13g2_decap_4 FILLER_22_340 ();
 sg13g2_decap_8 FILLER_22_400 ();
 sg13g2_fill_2 FILLER_22_407 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_98 ();
 sg13g2_decap_8 FILLER_23_105 ();
 sg13g2_decap_8 FILLER_23_112 ();
 sg13g2_decap_8 FILLER_23_119 ();
 sg13g2_decap_8 FILLER_23_126 ();
 sg13g2_decap_8 FILLER_23_133 ();
 sg13g2_decap_8 FILLER_23_140 ();
 sg13g2_decap_4 FILLER_23_147 ();
 sg13g2_fill_1 FILLER_23_151 ();
 sg13g2_fill_1 FILLER_23_185 ();
 sg13g2_decap_4 FILLER_23_264 ();
 sg13g2_fill_1 FILLER_23_277 ();
 sg13g2_fill_1 FILLER_23_365 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_decap_8 FILLER_24_98 ();
 sg13g2_decap_8 FILLER_24_105 ();
 sg13g2_decap_8 FILLER_24_112 ();
 sg13g2_decap_8 FILLER_24_119 ();
 sg13g2_decap_8 FILLER_24_126 ();
 sg13g2_decap_8 FILLER_24_133 ();
 sg13g2_decap_8 FILLER_24_140 ();
 sg13g2_fill_1 FILLER_24_147 ();
 sg13g2_decap_4 FILLER_24_191 ();
 sg13g2_fill_1 FILLER_24_227 ();
 sg13g2_fill_1 FILLER_24_250 ();
 sg13g2_fill_2 FILLER_24_261 ();
 sg13g2_fill_2 FILLER_24_277 ();
 sg13g2_fill_1 FILLER_24_295 ();
 sg13g2_fill_1 FILLER_24_324 ();
 sg13g2_fill_2 FILLER_24_350 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_8 FILLER_25_91 ();
 sg13g2_decap_8 FILLER_25_98 ();
 sg13g2_decap_8 FILLER_25_105 ();
 sg13g2_decap_8 FILLER_25_112 ();
 sg13g2_decap_8 FILLER_25_119 ();
 sg13g2_decap_8 FILLER_25_126 ();
 sg13g2_decap_4 FILLER_25_133 ();
 sg13g2_fill_2 FILLER_25_199 ();
 sg13g2_decap_4 FILLER_25_207 ();
 sg13g2_decap_4 FILLER_25_285 ();
 sg13g2_fill_1 FILLER_25_289 ();
 sg13g2_fill_1 FILLER_25_321 ();
 sg13g2_decap_4 FILLER_25_340 ();
 sg13g2_fill_1 FILLER_25_376 ();
 sg13g2_decap_4 FILLER_25_405 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_decap_8 FILLER_26_91 ();
 sg13g2_decap_8 FILLER_26_98 ();
 sg13g2_decap_8 FILLER_26_105 ();
 sg13g2_decap_8 FILLER_26_117 ();
 sg13g2_fill_2 FILLER_26_124 ();
 sg13g2_fill_1 FILLER_26_126 ();
 sg13g2_decap_8 FILLER_26_132 ();
 sg13g2_decap_8 FILLER_26_139 ();
 sg13g2_decap_4 FILLER_26_146 ();
 sg13g2_fill_2 FILLER_26_150 ();
 sg13g2_fill_1 FILLER_26_201 ();
 sg13g2_fill_2 FILLER_26_212 ();
 sg13g2_decap_4 FILLER_26_223 ();
 sg13g2_fill_2 FILLER_26_251 ();
 sg13g2_decap_4 FILLER_26_258 ();
 sg13g2_fill_1 FILLER_26_262 ();
 sg13g2_decap_4 FILLER_26_276 ();
 sg13g2_decap_8 FILLER_26_292 ();
 sg13g2_fill_1 FILLER_26_299 ();
 sg13g2_fill_2 FILLER_26_340 ();
 sg13g2_fill_1 FILLER_26_342 ();
 sg13g2_fill_1 FILLER_26_382 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_decap_8 FILLER_27_84 ();
 sg13g2_decap_8 FILLER_27_91 ();
 sg13g2_fill_1 FILLER_27_98 ();
 sg13g2_fill_2 FILLER_27_108 ();
 sg13g2_decap_4 FILLER_27_125 ();
 sg13g2_fill_2 FILLER_27_138 ();
 sg13g2_decap_8 FILLER_27_149 ();
 sg13g2_decap_4 FILLER_27_156 ();
 sg13g2_fill_1 FILLER_27_200 ();
 sg13g2_fill_2 FILLER_27_209 ();
 sg13g2_fill_2 FILLER_27_279 ();
 sg13g2_fill_1 FILLER_27_281 ();
 sg13g2_decap_8 FILLER_27_299 ();
 sg13g2_fill_2 FILLER_27_314 ();
 sg13g2_fill_1 FILLER_27_316 ();
 sg13g2_decap_8 FILLER_27_338 ();
 sg13g2_fill_2 FILLER_27_345 ();
 sg13g2_fill_1 FILLER_27_347 ();
 sg13g2_fill_1 FILLER_27_368 ();
 sg13g2_decap_4 FILLER_27_403 ();
 sg13g2_fill_2 FILLER_27_407 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_decap_4 FILLER_28_110 ();
 sg13g2_fill_2 FILLER_28_123 ();
 sg13g2_fill_1 FILLER_28_125 ();
 sg13g2_decap_4 FILLER_28_152 ();
 sg13g2_fill_2 FILLER_28_156 ();
 sg13g2_fill_2 FILLER_28_166 ();
 sg13g2_fill_2 FILLER_28_175 ();
 sg13g2_fill_1 FILLER_28_228 ();
 sg13g2_decap_8 FILLER_28_242 ();
 sg13g2_decap_8 FILLER_28_249 ();
 sg13g2_decap_4 FILLER_28_256 ();
 sg13g2_fill_1 FILLER_28_260 ();
 sg13g2_decap_8 FILLER_28_268 ();
 sg13g2_decap_4 FILLER_28_275 ();
 sg13g2_fill_2 FILLER_28_309 ();
 sg13g2_fill_1 FILLER_28_311 ();
 sg13g2_fill_2 FILLER_28_317 ();
 sg13g2_fill_2 FILLER_28_338 ();
 sg13g2_fill_1 FILLER_28_361 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_decap_8 FILLER_29_84 ();
 sg13g2_fill_2 FILLER_29_91 ();
 sg13g2_decap_4 FILLER_29_102 ();
 sg13g2_fill_1 FILLER_29_106 ();
 sg13g2_fill_2 FILLER_29_136 ();
 sg13g2_decap_8 FILLER_29_145 ();
 sg13g2_fill_1 FILLER_29_152 ();
 sg13g2_fill_2 FILLER_29_161 ();
 sg13g2_fill_1 FILLER_29_204 ();
 sg13g2_fill_2 FILLER_29_243 ();
 sg13g2_decap_4 FILLER_29_259 ();
 sg13g2_decap_4 FILLER_29_286 ();
 sg13g2_fill_2 FILLER_29_290 ();
 sg13g2_fill_1 FILLER_29_297 ();
 sg13g2_fill_1 FILLER_29_308 ();
 sg13g2_fill_2 FILLER_29_328 ();
 sg13g2_fill_1 FILLER_29_330 ();
 sg13g2_decap_4 FILLER_29_339 ();
 sg13g2_fill_2 FILLER_29_343 ();
 sg13g2_fill_2 FILLER_29_373 ();
 sg13g2_fill_1 FILLER_29_382 ();
 sg13g2_fill_2 FILLER_29_392 ();
 sg13g2_fill_1 FILLER_29_408 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_4 FILLER_30_70 ();
 sg13g2_fill_1 FILLER_30_74 ();
 sg13g2_fill_1 FILLER_30_104 ();
 sg13g2_fill_2 FILLER_30_162 ();
 sg13g2_fill_1 FILLER_30_164 ();
 sg13g2_fill_1 FILLER_30_170 ();
 sg13g2_fill_2 FILLER_30_227 ();
 sg13g2_fill_2 FILLER_30_244 ();
 sg13g2_fill_1 FILLER_30_256 ();
 sg13g2_fill_1 FILLER_30_262 ();
 sg13g2_decap_4 FILLER_30_282 ();
 sg13g2_fill_2 FILLER_30_286 ();
 sg13g2_fill_1 FILLER_30_315 ();
 sg13g2_fill_2 FILLER_30_348 ();
 sg13g2_decap_4 FILLER_30_360 ();
 sg13g2_fill_1 FILLER_30_364 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_decap_8 FILLER_31_84 ();
 sg13g2_decap_8 FILLER_31_91 ();
 sg13g2_decap_8 FILLER_31_98 ();
 sg13g2_fill_2 FILLER_31_105 ();
 sg13g2_fill_2 FILLER_31_123 ();
 sg13g2_fill_2 FILLER_31_138 ();
 sg13g2_decap_8 FILLER_31_145 ();
 sg13g2_fill_1 FILLER_31_152 ();
 sg13g2_fill_2 FILLER_31_178 ();
 sg13g2_fill_1 FILLER_31_180 ();
 sg13g2_decap_8 FILLER_31_202 ();
 sg13g2_decap_8 FILLER_31_209 ();
 sg13g2_fill_1 FILLER_31_232 ();
 sg13g2_fill_1 FILLER_31_238 ();
 sg13g2_fill_2 FILLER_31_254 ();
 sg13g2_decap_4 FILLER_31_261 ();
 sg13g2_fill_1 FILLER_31_265 ();
 sg13g2_fill_2 FILLER_31_275 ();
 sg13g2_fill_2 FILLER_31_282 ();
 sg13g2_decap_8 FILLER_31_289 ();
 sg13g2_fill_1 FILLER_31_296 ();
 sg13g2_fill_2 FILLER_31_303 ();
 sg13g2_fill_1 FILLER_31_305 ();
 sg13g2_fill_2 FILLER_31_314 ();
 sg13g2_decap_4 FILLER_31_320 ();
 sg13g2_decap_8 FILLER_31_329 ();
 sg13g2_decap_4 FILLER_31_336 ();
 sg13g2_fill_2 FILLER_31_340 ();
 sg13g2_fill_2 FILLER_31_359 ();
 sg13g2_fill_1 FILLER_31_376 ();
 sg13g2_fill_1 FILLER_31_382 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_4 FILLER_32_77 ();
 sg13g2_fill_2 FILLER_32_81 ();
 sg13g2_fill_2 FILLER_32_128 ();
 sg13g2_fill_1 FILLER_32_130 ();
 sg13g2_fill_2 FILLER_32_157 ();
 sg13g2_decap_8 FILLER_32_213 ();
 sg13g2_fill_2 FILLER_32_220 ();
 sg13g2_fill_2 FILLER_32_237 ();
 sg13g2_fill_1 FILLER_32_239 ();
 sg13g2_fill_2 FILLER_32_247 ();
 sg13g2_fill_2 FILLER_32_257 ();
 sg13g2_decap_4 FILLER_32_277 ();
 sg13g2_decap_8 FILLER_32_296 ();
 sg13g2_decap_8 FILLER_32_303 ();
 sg13g2_fill_2 FILLER_32_310 ();
 sg13g2_fill_1 FILLER_32_329 ();
 sg13g2_fill_2 FILLER_32_338 ();
 sg13g2_fill_1 FILLER_32_340 ();
 sg13g2_decap_4 FILLER_32_354 ();
 sg13g2_decap_4 FILLER_32_379 ();
 sg13g2_fill_1 FILLER_32_392 ();
 sg13g2_decap_8 FILLER_32_402 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_decap_8 FILLER_33_91 ();
 sg13g2_fill_1 FILLER_33_98 ();
 sg13g2_fill_2 FILLER_33_107 ();
 sg13g2_fill_2 FILLER_33_123 ();
 sg13g2_fill_1 FILLER_33_125 ();
 sg13g2_fill_1 FILLER_33_145 ();
 sg13g2_fill_2 FILLER_33_155 ();
 sg13g2_fill_1 FILLER_33_162 ();
 sg13g2_fill_2 FILLER_33_198 ();
 sg13g2_decap_8 FILLER_33_212 ();
 sg13g2_decap_8 FILLER_33_219 ();
 sg13g2_fill_1 FILLER_33_230 ();
 sg13g2_decap_4 FILLER_33_240 ();
 sg13g2_decap_8 FILLER_33_249 ();
 sg13g2_fill_1 FILLER_33_256 ();
 sg13g2_decap_4 FILLER_33_262 ();
 sg13g2_fill_1 FILLER_33_266 ();
 sg13g2_decap_8 FILLER_33_272 ();
 sg13g2_fill_1 FILLER_33_279 ();
 sg13g2_decap_8 FILLER_33_285 ();
 sg13g2_fill_1 FILLER_33_292 ();
 sg13g2_decap_4 FILLER_33_306 ();
 sg13g2_fill_1 FILLER_33_310 ();
 sg13g2_fill_2 FILLER_33_321 ();
 sg13g2_decap_8 FILLER_33_332 ();
 sg13g2_fill_2 FILLER_33_339 ();
 sg13g2_fill_1 FILLER_33_341 ();
 sg13g2_decap_8 FILLER_33_351 ();
 sg13g2_fill_1 FILLER_33_358 ();
 sg13g2_decap_4 FILLER_33_374 ();
 sg13g2_fill_1 FILLER_33_378 ();
 sg13g2_decap_8 FILLER_33_384 ();
 sg13g2_fill_2 FILLER_33_391 ();
 sg13g2_decap_8 FILLER_33_402 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_4 FILLER_34_84 ();
 sg13g2_fill_1 FILLER_34_114 ();
 sg13g2_fill_2 FILLER_34_130 ();
 sg13g2_fill_1 FILLER_34_150 ();
 sg13g2_fill_1 FILLER_34_182 ();
 sg13g2_decap_4 FILLER_34_191 ();
 sg13g2_fill_1 FILLER_34_195 ();
 sg13g2_decap_4 FILLER_34_210 ();
 sg13g2_fill_2 FILLER_34_214 ();
 sg13g2_fill_1 FILLER_34_237 ();
 sg13g2_fill_2 FILLER_34_246 ();
 sg13g2_fill_2 FILLER_34_256 ();
 sg13g2_fill_1 FILLER_34_258 ();
 sg13g2_fill_1 FILLER_34_266 ();
 sg13g2_fill_2 FILLER_34_284 ();
 sg13g2_fill_2 FILLER_34_326 ();
 sg13g2_fill_2 FILLER_34_344 ();
 sg13g2_fill_2 FILLER_34_360 ();
 sg13g2_decap_8 FILLER_34_380 ();
 sg13g2_decap_8 FILLER_34_387 ();
 sg13g2_decap_8 FILLER_34_394 ();
 sg13g2_decap_8 FILLER_34_401 ();
 sg13g2_fill_1 FILLER_34_408 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_4 FILLER_35_77 ();
 sg13g2_fill_1 FILLER_35_81 ();
 sg13g2_fill_1 FILLER_35_108 ();
 sg13g2_decap_4 FILLER_35_153 ();
 sg13g2_fill_1 FILLER_35_157 ();
 sg13g2_fill_2 FILLER_35_179 ();
 sg13g2_fill_1 FILLER_35_181 ();
 sg13g2_decap_8 FILLER_35_202 ();
 sg13g2_decap_4 FILLER_35_209 ();
 sg13g2_fill_1 FILLER_35_213 ();
 sg13g2_fill_2 FILLER_35_230 ();
 sg13g2_fill_1 FILLER_35_232 ();
 sg13g2_fill_2 FILLER_35_253 ();
 sg13g2_fill_1 FILLER_35_255 ();
 sg13g2_decap_8 FILLER_35_285 ();
 sg13g2_fill_2 FILLER_35_292 ();
 sg13g2_fill_1 FILLER_35_307 ();
 sg13g2_decap_4 FILLER_35_313 ();
 sg13g2_fill_2 FILLER_35_317 ();
 sg13g2_fill_1 FILLER_35_322 ();
 sg13g2_fill_1 FILLER_35_327 ();
 sg13g2_decap_8 FILLER_35_336 ();
 sg13g2_decap_4 FILLER_35_343 ();
 sg13g2_fill_2 FILLER_35_347 ();
 sg13g2_decap_8 FILLER_35_354 ();
 sg13g2_fill_2 FILLER_35_361 ();
 sg13g2_fill_1 FILLER_35_363 ();
 sg13g2_decap_8 FILLER_35_374 ();
 sg13g2_decap_8 FILLER_35_381 ();
 sg13g2_decap_8 FILLER_35_388 ();
 sg13g2_decap_8 FILLER_35_395 ();
 sg13g2_decap_8 FILLER_35_402 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_fill_2 FILLER_36_91 ();
 sg13g2_fill_2 FILLER_36_128 ();
 sg13g2_fill_2 FILLER_36_139 ();
 sg13g2_fill_1 FILLER_36_141 ();
 sg13g2_fill_2 FILLER_36_155 ();
 sg13g2_decap_8 FILLER_36_171 ();
 sg13g2_decap_8 FILLER_36_178 ();
 sg13g2_decap_8 FILLER_36_185 ();
 sg13g2_decap_4 FILLER_36_192 ();
 sg13g2_decap_4 FILLER_36_205 ();
 sg13g2_fill_1 FILLER_36_213 ();
 sg13g2_fill_2 FILLER_36_222 ();
 sg13g2_decap_8 FILLER_36_251 ();
 sg13g2_fill_1 FILLER_36_264 ();
 sg13g2_decap_8 FILLER_36_273 ();
 sg13g2_fill_1 FILLER_36_280 ();
 sg13g2_fill_1 FILLER_36_286 ();
 sg13g2_fill_2 FILLER_36_304 ();
 sg13g2_decap_4 FILLER_36_319 ();
 sg13g2_fill_2 FILLER_36_336 ();
 sg13g2_fill_1 FILLER_36_338 ();
 sg13g2_fill_2 FILLER_36_364 ();
 sg13g2_fill_1 FILLER_36_366 ();
 sg13g2_decap_8 FILLER_36_382 ();
 sg13g2_decap_8 FILLER_36_389 ();
 sg13g2_decap_8 FILLER_36_396 ();
 sg13g2_decap_4 FILLER_36_403 ();
 sg13g2_fill_2 FILLER_36_407 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_4 FILLER_37_77 ();
 sg13g2_fill_2 FILLER_37_81 ();
 sg13g2_fill_2 FILLER_37_109 ();
 sg13g2_fill_2 FILLER_37_149 ();
 sg13g2_decap_8 FILLER_37_195 ();
 sg13g2_fill_1 FILLER_37_202 ();
 sg13g2_fill_2 FILLER_37_224 ();
 sg13g2_fill_2 FILLER_37_286 ();
 sg13g2_fill_2 FILLER_37_293 ();
 sg13g2_fill_1 FILLER_37_295 ();
 sg13g2_fill_2 FILLER_37_316 ();
 sg13g2_decap_8 FILLER_37_367 ();
 sg13g2_decap_8 FILLER_37_374 ();
 sg13g2_decap_8 FILLER_37_381 ();
 sg13g2_decap_8 FILLER_37_388 ();
 sg13g2_decap_8 FILLER_37_395 ();
 sg13g2_decap_8 FILLER_37_402 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_4 FILLER_38_60 ();
 sg13g2_decap_4 FILLER_38_68 ();
 sg13g2_decap_4 FILLER_38_76 ();
 sg13g2_decap_4 FILLER_38_84 ();
 sg13g2_fill_1 FILLER_38_92 ();
 sg13g2_fill_1 FILLER_38_132 ();
 sg13g2_decap_4 FILLER_38_151 ();
 sg13g2_fill_2 FILLER_38_155 ();
 sg13g2_decap_4 FILLER_38_165 ();
 sg13g2_fill_1 FILLER_38_169 ();
 sg13g2_decap_4 FILLER_38_179 ();
 sg13g2_fill_1 FILLER_38_183 ();
 sg13g2_decap_4 FILLER_38_188 ();
 sg13g2_decap_4 FILLER_38_196 ();
 sg13g2_decap_4 FILLER_38_204 ();
 sg13g2_fill_2 FILLER_38_228 ();
 sg13g2_fill_1 FILLER_38_230 ();
 sg13g2_decap_8 FILLER_38_240 ();
 sg13g2_fill_1 FILLER_38_247 ();
 sg13g2_fill_2 FILLER_38_261 ();
 sg13g2_fill_1 FILLER_38_263 ();
 sg13g2_fill_2 FILLER_38_269 ();
 sg13g2_fill_1 FILLER_38_271 ();
 sg13g2_fill_1 FILLER_38_303 ();
 sg13g2_fill_2 FILLER_38_317 ();
 sg13g2_fill_1 FILLER_38_319 ();
 sg13g2_fill_1 FILLER_38_330 ();
 sg13g2_fill_2 FILLER_38_349 ();
 sg13g2_fill_1 FILLER_38_367 ();
 sg13g2_decap_8 FILLER_38_373 ();
 sg13g2_decap_8 FILLER_38_380 ();
 sg13g2_decap_8 FILLER_38_387 ();
 sg13g2_decap_8 FILLER_38_394 ();
 sg13g2_decap_8 FILLER_38_401 ();
 sg13g2_fill_1 FILLER_38_408 ();
 assign uio_oe[0] = net14;
 assign uio_oe[1] = net15;
 assign uio_oe[2] = net16;
 assign uio_oe[3] = net17;
 assign uio_oe[4] = net18;
 assign uio_oe[5] = net19;
 assign uio_oe[6] = net20;
 assign uio_oe[7] = net21;
 assign uo_out[2] = net22;
 assign uo_out[3] = net23;
 assign uo_out[4] = net24;
 assign uo_out[5] = net25;
 assign uo_out[6] = net26;
 assign uo_out[7] = net27;
endmodule
